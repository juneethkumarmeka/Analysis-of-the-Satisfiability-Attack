module basic_3000_30000_3500_25_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_2646,In_1527);
xor U1 (N_1,In_2980,In_2703);
or U2 (N_2,In_1792,In_2604);
and U3 (N_3,In_1200,In_2757);
or U4 (N_4,In_1075,In_2003);
nand U5 (N_5,In_132,In_906);
xnor U6 (N_6,In_2833,In_711);
and U7 (N_7,In_1327,In_2183);
nand U8 (N_8,In_2236,In_1514);
xor U9 (N_9,In_2205,In_2756);
nand U10 (N_10,In_257,In_2537);
and U11 (N_11,In_288,In_1165);
xor U12 (N_12,In_909,In_815);
or U13 (N_13,In_979,In_1612);
nor U14 (N_14,In_1584,In_541);
nor U15 (N_15,In_1754,In_141);
nand U16 (N_16,In_2777,In_1941);
and U17 (N_17,In_1014,In_1274);
nand U18 (N_18,In_1846,In_753);
xnor U19 (N_19,In_2953,In_1302);
nand U20 (N_20,In_360,In_76);
nor U21 (N_21,In_1541,In_2843);
nor U22 (N_22,In_39,In_1288);
nand U23 (N_23,In_1565,In_1083);
nor U24 (N_24,In_1537,In_876);
nand U25 (N_25,In_1155,In_210);
xnor U26 (N_26,In_649,In_1618);
xnor U27 (N_27,In_1556,In_2421);
and U28 (N_28,In_406,In_1539);
nand U29 (N_29,In_990,In_1477);
and U30 (N_30,In_608,In_1436);
xor U31 (N_31,In_1358,In_648);
or U32 (N_32,In_2311,In_2288);
xor U33 (N_33,In_2123,In_1210);
or U34 (N_34,In_681,In_2717);
or U35 (N_35,In_2344,In_184);
nor U36 (N_36,In_462,In_1986);
and U37 (N_37,In_1172,In_1797);
or U38 (N_38,In_757,In_2088);
or U39 (N_39,In_2232,In_2367);
or U40 (N_40,In_1933,In_236);
nor U41 (N_41,In_350,In_1608);
and U42 (N_42,In_584,In_2809);
or U43 (N_43,In_485,In_2971);
and U44 (N_44,In_2093,In_836);
nand U45 (N_45,In_2231,In_7);
xnor U46 (N_46,In_1446,In_2138);
nand U47 (N_47,In_1983,In_286);
or U48 (N_48,In_2171,In_1273);
or U49 (N_49,In_1790,In_1115);
nand U50 (N_50,In_583,In_2496);
xnor U51 (N_51,In_1648,In_1109);
nor U52 (N_52,In_358,In_1750);
xor U53 (N_53,In_2312,In_1837);
or U54 (N_54,In_915,In_1409);
xor U55 (N_55,In_827,In_2209);
nor U56 (N_56,In_1704,In_847);
nor U57 (N_57,In_1043,In_2921);
or U58 (N_58,In_606,In_1632);
or U59 (N_59,In_2359,In_49);
xnor U60 (N_60,In_460,In_2148);
nand U61 (N_61,In_2876,In_593);
nand U62 (N_62,In_264,In_1135);
xnor U63 (N_63,In_2340,In_1237);
xnor U64 (N_64,In_1830,In_1993);
nand U65 (N_65,In_1832,In_200);
nor U66 (N_66,In_2126,In_800);
nor U67 (N_67,In_919,In_2939);
nor U68 (N_68,In_722,In_1473);
nor U69 (N_69,In_837,In_1300);
xor U70 (N_70,In_225,In_659);
xnor U71 (N_71,In_1817,In_2742);
nor U72 (N_72,In_529,In_1851);
nor U73 (N_73,In_2070,In_653);
or U74 (N_74,In_1079,In_1478);
and U75 (N_75,In_2701,In_1948);
nor U76 (N_76,In_89,In_120);
xnor U77 (N_77,In_1679,In_2060);
and U78 (N_78,In_638,In_448);
or U79 (N_79,In_2861,In_2597);
nor U80 (N_80,In_1206,In_2897);
or U81 (N_81,In_280,In_2035);
xor U82 (N_82,In_1913,In_705);
and U83 (N_83,In_1201,In_2838);
nor U84 (N_84,In_1928,In_1470);
nand U85 (N_85,In_1720,In_521);
xnor U86 (N_86,In_715,In_609);
nor U87 (N_87,In_1334,In_586);
nand U88 (N_88,In_1108,In_1220);
nand U89 (N_89,In_1410,In_3);
nor U90 (N_90,In_1439,In_641);
nand U91 (N_91,In_1377,In_1449);
nand U92 (N_92,In_1569,In_2476);
xor U93 (N_93,In_1959,In_2101);
and U94 (N_94,In_1225,In_870);
nand U95 (N_95,In_374,In_2918);
nor U96 (N_96,In_1884,In_1329);
xnor U97 (N_97,In_773,In_2736);
nand U98 (N_98,In_552,In_1250);
or U99 (N_99,In_2135,In_390);
nor U100 (N_100,In_18,In_1758);
nor U101 (N_101,In_109,In_1634);
xnor U102 (N_102,In_871,In_183);
or U103 (N_103,In_1291,In_2002);
xor U104 (N_104,In_1550,In_1783);
xor U105 (N_105,In_1474,In_2022);
xnor U106 (N_106,In_1796,In_1886);
nor U107 (N_107,In_1232,In_2826);
and U108 (N_108,In_2629,In_1977);
nand U109 (N_109,In_1405,In_180);
nor U110 (N_110,In_2474,In_233);
and U111 (N_111,In_978,In_585);
or U112 (N_112,In_53,In_492);
or U113 (N_113,In_1203,In_1373);
and U114 (N_114,In_2361,In_304);
nand U115 (N_115,In_1150,In_381);
or U116 (N_116,In_2743,In_154);
xnor U117 (N_117,In_664,In_537);
nor U118 (N_118,In_2178,In_289);
xor U119 (N_119,In_400,In_2529);
xor U120 (N_120,In_1209,In_291);
nand U121 (N_121,In_307,In_2674);
or U122 (N_122,In_2572,In_311);
or U123 (N_123,In_656,In_54);
xor U124 (N_124,In_2976,In_1099);
xor U125 (N_125,In_2201,In_781);
nand U126 (N_126,In_1022,In_2341);
nor U127 (N_127,In_1320,In_153);
nor U128 (N_128,In_1169,In_762);
nor U129 (N_129,In_735,In_2793);
and U130 (N_130,In_113,In_1778);
and U131 (N_131,In_1205,In_2563);
and U132 (N_132,In_1416,In_1950);
nor U133 (N_133,In_1516,In_1581);
or U134 (N_134,In_260,In_103);
xnor U135 (N_135,In_2776,In_1147);
nor U136 (N_136,In_2654,In_2159);
xnor U137 (N_137,In_2274,In_1283);
nor U138 (N_138,In_118,In_738);
xor U139 (N_139,In_2914,In_1860);
nand U140 (N_140,In_1380,In_1735);
or U141 (N_141,In_646,In_69);
or U142 (N_142,In_241,In_2540);
xor U143 (N_143,In_1666,In_830);
nor U144 (N_144,In_918,In_21);
nand U145 (N_145,In_1806,In_614);
xnor U146 (N_146,In_2521,In_235);
nor U147 (N_147,In_2078,In_734);
nand U148 (N_148,In_563,In_1518);
xnor U149 (N_149,In_1064,In_96);
nand U150 (N_150,In_2439,In_904);
xor U151 (N_151,In_469,In_2010);
nand U152 (N_152,In_323,In_1231);
nor U153 (N_153,In_1143,In_65);
nand U154 (N_154,In_2794,In_926);
xor U155 (N_155,In_293,In_393);
xnor U156 (N_156,In_1167,In_1962);
xnor U157 (N_157,In_1825,In_1211);
xnor U158 (N_158,In_305,In_1642);
or U159 (N_159,In_556,In_2357);
and U160 (N_160,In_1828,In_2266);
nand U161 (N_161,In_631,In_453);
nor U162 (N_162,In_512,In_2734);
or U163 (N_163,In_553,In_1363);
and U164 (N_164,In_888,In_1719);
nand U165 (N_165,In_1271,In_2260);
and U166 (N_166,In_2940,In_2542);
and U167 (N_167,In_1713,In_2873);
xor U168 (N_168,In_1768,In_680);
or U169 (N_169,In_1515,In_254);
nor U170 (N_170,In_1114,In_1568);
nand U171 (N_171,In_1818,In_1492);
nor U172 (N_172,In_945,In_1392);
xnor U173 (N_173,In_2835,In_226);
xnor U174 (N_174,In_2589,In_1090);
xnor U175 (N_175,In_2422,In_1272);
xor U176 (N_176,In_2075,In_1062);
xor U177 (N_177,In_2056,In_1775);
nor U178 (N_178,In_2841,In_1965);
and U179 (N_179,In_1468,In_2272);
nor U180 (N_180,In_1630,In_295);
nand U181 (N_181,In_494,In_952);
or U182 (N_182,In_1918,In_1954);
nor U183 (N_183,In_48,In_2883);
or U184 (N_184,In_1265,In_1123);
nand U185 (N_185,In_2112,In_2225);
nor U186 (N_186,In_2983,In_1655);
nor U187 (N_187,In_2040,In_1289);
nand U188 (N_188,In_519,In_1803);
nor U189 (N_189,In_679,In_452);
xnor U190 (N_190,In_961,In_2160);
nor U191 (N_191,In_2658,In_2599);
and U192 (N_192,In_2220,In_2299);
and U193 (N_193,In_694,In_2251);
nor U194 (N_194,In_176,In_2402);
xnor U195 (N_195,In_1465,In_1684);
or U196 (N_196,In_2106,In_1802);
nand U197 (N_197,In_1957,In_1239);
xor U198 (N_198,In_2152,In_1985);
or U199 (N_199,In_2417,In_2552);
xnor U200 (N_200,In_1042,In_999);
and U201 (N_201,In_538,In_1512);
and U202 (N_202,In_473,In_1498);
or U203 (N_203,In_2189,In_1489);
nand U204 (N_204,In_1670,In_514);
or U205 (N_205,In_376,In_2096);
and U206 (N_206,In_2760,In_2238);
or U207 (N_207,In_2142,In_2615);
and U208 (N_208,In_2676,In_2023);
or U209 (N_209,In_2694,In_1738);
nand U210 (N_210,In_969,In_1972);
nand U211 (N_211,In_2191,In_838);
xor U212 (N_212,In_2398,In_1412);
nor U213 (N_213,In_768,In_2788);
or U214 (N_214,In_2036,In_240);
or U215 (N_215,In_1445,In_1773);
nand U216 (N_216,In_943,In_33);
nor U217 (N_217,In_1103,In_1030);
xor U218 (N_218,In_2371,In_205);
nand U219 (N_219,In_2234,In_855);
xnor U220 (N_220,In_691,In_1112);
xnor U221 (N_221,In_1736,In_145);
xor U222 (N_222,In_946,In_1127);
and U223 (N_223,In_951,In_1558);
xnor U224 (N_224,In_825,In_2771);
xor U225 (N_225,In_1301,In_309);
xnor U226 (N_226,In_2878,In_2305);
or U227 (N_227,In_2484,In_2591);
nor U228 (N_228,In_1906,In_2320);
and U229 (N_229,In_81,In_2194);
xnor U230 (N_230,In_1786,In_1572);
nor U231 (N_231,In_1129,In_1888);
nand U232 (N_232,In_1138,In_1900);
or U233 (N_233,In_2558,In_312);
and U234 (N_234,In_1069,In_1545);
nor U235 (N_235,In_2334,In_1943);
and U236 (N_236,In_2568,In_2192);
or U237 (N_237,In_1882,In_2764);
nor U238 (N_238,In_1945,In_630);
or U239 (N_239,In_2864,In_921);
xnor U240 (N_240,In_2202,In_1348);
xor U241 (N_241,In_2773,In_195);
nor U242 (N_242,In_139,In_51);
nand U243 (N_243,In_138,In_1314);
nor U244 (N_244,In_980,In_1659);
nand U245 (N_245,In_1092,In_2387);
or U246 (N_246,In_1893,In_1927);
xor U247 (N_247,In_2089,In_1868);
or U248 (N_248,In_1134,In_1344);
or U249 (N_249,In_1379,In_95);
nand U250 (N_250,In_1304,In_2098);
and U251 (N_251,In_1374,In_1493);
or U252 (N_252,In_1184,In_480);
nor U253 (N_253,In_1095,In_721);
nor U254 (N_254,In_2051,In_610);
nand U255 (N_255,In_2620,In_2718);
nor U256 (N_256,In_2170,In_2784);
xnor U257 (N_257,In_1607,In_8);
xnor U258 (N_258,In_808,In_643);
xor U259 (N_259,In_2923,In_2808);
nand U260 (N_260,In_334,In_156);
nor U261 (N_261,In_2968,In_2292);
nor U262 (N_262,In_2814,In_1491);
and U263 (N_263,In_2603,In_337);
and U264 (N_264,In_2375,In_2887);
xnor U265 (N_265,In_2011,In_2265);
nor U266 (N_266,In_2570,In_1524);
nand U267 (N_267,In_947,In_2627);
or U268 (N_268,In_1311,In_1430);
nand U269 (N_269,In_2043,In_1080);
and U270 (N_270,In_1873,In_821);
xnor U271 (N_271,In_2698,In_761);
or U272 (N_272,In_1819,In_395);
and U273 (N_273,In_1332,In_1251);
nor U274 (N_274,In_661,In_2435);
nor U275 (N_275,In_1345,In_190);
or U276 (N_276,In_1816,In_412);
xnor U277 (N_277,In_1907,In_1106);
xor U278 (N_278,In_1644,In_1234);
and U279 (N_279,In_955,In_2304);
and U280 (N_280,In_461,In_434);
xor U281 (N_281,In_2221,In_1598);
xor U282 (N_282,In_981,In_887);
or U283 (N_283,In_2210,In_1708);
nor U284 (N_284,In_1371,In_2198);
or U285 (N_285,In_532,In_881);
or U286 (N_286,In_2640,In_1450);
xnor U287 (N_287,In_1676,In_1898);
and U288 (N_288,In_1890,In_1215);
nand U289 (N_289,In_573,In_447);
nor U290 (N_290,In_2463,In_2522);
nor U291 (N_291,In_2016,In_2066);
and U292 (N_292,In_645,In_1742);
nand U293 (N_293,In_1551,In_2120);
nor U294 (N_294,In_2704,In_256);
nand U295 (N_295,In_404,In_1994);
nor U296 (N_296,In_1388,In_787);
nor U297 (N_297,In_2626,In_547);
and U298 (N_298,In_1864,In_2127);
and U299 (N_299,In_269,In_427);
and U300 (N_300,In_418,In_1519);
or U301 (N_301,In_2073,In_809);
nand U302 (N_302,In_2445,In_755);
xor U303 (N_303,In_1966,In_451);
or U304 (N_304,In_2867,In_2337);
and U305 (N_305,In_468,In_303);
and U306 (N_306,In_2740,In_2319);
nor U307 (N_307,In_474,In_351);
nor U308 (N_308,In_1964,In_581);
or U309 (N_309,In_28,In_2947);
xor U310 (N_310,In_2578,In_1255);
xor U311 (N_311,In_1511,In_930);
and U312 (N_312,In_1086,In_1457);
or U313 (N_313,In_1743,In_2748);
nor U314 (N_314,In_208,In_34);
or U315 (N_315,In_2103,In_2416);
nor U316 (N_316,In_594,In_2353);
and U317 (N_317,In_626,In_1590);
nor U318 (N_318,In_1940,In_2770);
or U319 (N_319,In_740,In_867);
nor U320 (N_320,In_1126,In_384);
and U321 (N_321,In_507,In_696);
and U322 (N_322,In_1880,In_84);
nand U323 (N_323,In_1001,In_939);
nor U324 (N_324,In_336,In_2431);
nor U325 (N_325,In_2048,In_1751);
nand U326 (N_326,In_1160,In_2928);
xnor U327 (N_327,In_2163,In_1012);
xnor U328 (N_328,In_2847,In_2107);
xnor U329 (N_329,In_565,In_900);
or U330 (N_330,In_2598,In_159);
nand U331 (N_331,In_315,In_1267);
and U332 (N_332,In_2638,In_2392);
and U333 (N_333,In_501,In_2839);
or U334 (N_334,In_1257,In_2269);
and U335 (N_335,In_1253,In_2042);
xor U336 (N_336,In_908,In_2677);
and U337 (N_337,In_826,In_1107);
nand U338 (N_338,In_2280,In_123);
and U339 (N_339,In_2630,In_1858);
xnor U340 (N_340,In_2019,In_2014);
or U341 (N_341,In_824,In_2915);
nand U342 (N_342,In_2328,In_729);
and U343 (N_343,In_1661,In_793);
nor U344 (N_344,In_758,In_2739);
or U345 (N_345,In_2336,In_328);
or U346 (N_346,In_1869,In_2896);
nand U347 (N_347,In_2506,In_903);
xor U348 (N_348,In_2574,In_2176);
or U349 (N_349,In_249,In_2696);
or U350 (N_350,In_987,In_2390);
or U351 (N_351,In_1694,In_2689);
or U352 (N_352,In_1722,In_1402);
xor U353 (N_353,In_1045,In_419);
xnor U354 (N_354,In_1047,In_2612);
nor U355 (N_355,In_2716,In_2486);
nor U356 (N_356,In_223,In_2936);
nor U357 (N_357,In_1259,In_2984);
nor U358 (N_358,In_267,In_2785);
or U359 (N_359,In_2779,In_2609);
nor U360 (N_360,In_2219,In_2741);
and U361 (N_361,In_1098,In_970);
nand U362 (N_362,In_739,In_2645);
nor U363 (N_363,In_318,In_2356);
nor U364 (N_364,In_684,In_2875);
nand U365 (N_365,In_25,In_1488);
nand U366 (N_366,In_2683,In_36);
xor U367 (N_367,In_1157,In_2081);
nand U368 (N_368,In_604,In_1595);
xor U369 (N_369,In_2182,In_378);
nand U370 (N_370,In_1531,In_1875);
xor U371 (N_371,In_963,In_2457);
xnor U372 (N_372,In_2263,In_2245);
or U373 (N_373,In_72,In_2715);
nor U374 (N_374,In_513,In_2907);
or U375 (N_375,In_2203,In_320);
nand U376 (N_376,In_1383,In_588);
xnor U377 (N_377,In_234,In_255);
and U378 (N_378,In_2283,In_278);
xor U379 (N_379,In_1024,In_2097);
or U380 (N_380,In_1417,In_2854);
nor U381 (N_381,In_441,In_1153);
xor U382 (N_382,In_1894,In_1261);
nor U383 (N_383,In_263,In_1101);
and U384 (N_384,In_807,In_2555);
and U385 (N_385,In_2149,In_329);
and U386 (N_386,In_1523,In_791);
or U387 (N_387,In_1480,In_2362);
xor U388 (N_388,In_471,In_428);
nand U389 (N_389,In_2721,In_1386);
xor U390 (N_390,In_1503,In_134);
nand U391 (N_391,In_2270,In_202);
nand U392 (N_392,In_43,In_1822);
nor U393 (N_393,In_2383,In_1823);
nor U394 (N_394,In_247,In_704);
and U395 (N_395,In_306,In_672);
nand U396 (N_396,In_2863,In_701);
or U397 (N_397,In_1501,In_2366);
nand U398 (N_398,In_1988,In_2026);
nand U399 (N_399,In_1370,In_1769);
nand U400 (N_400,In_292,In_1422);
nor U401 (N_401,In_1840,In_17);
and U402 (N_402,In_112,In_2514);
xnor U403 (N_403,In_968,In_1174);
nor U404 (N_404,In_1861,In_1441);
or U405 (N_405,In_844,In_2360);
or U406 (N_406,In_2850,In_1223);
xnor U407 (N_407,In_2027,In_2543);
or U408 (N_408,In_2333,In_94);
nand U409 (N_409,In_1507,In_2548);
nand U410 (N_410,In_2651,In_1040);
nor U411 (N_411,In_2637,In_2623);
or U412 (N_412,In_491,In_639);
nand U413 (N_413,In_2799,In_1308);
nand U414 (N_414,In_1168,In_2924);
xnor U415 (N_415,In_2140,In_651);
and U416 (N_416,In_2859,In_2471);
nor U417 (N_417,In_2158,In_1481);
or U418 (N_418,In_1831,In_107);
xor U419 (N_419,In_2146,In_1467);
or U420 (N_420,In_1159,In_2750);
or U421 (N_421,In_251,In_1820);
xor U422 (N_422,In_476,In_355);
xor U423 (N_423,In_1924,In_935);
xor U424 (N_424,In_1362,In_879);
nand U425 (N_425,In_1725,In_2571);
and U426 (N_426,In_1350,In_265);
nor U427 (N_427,In_566,In_228);
nor U428 (N_428,In_1285,In_1357);
and U429 (N_429,In_2485,In_1997);
nor U430 (N_430,In_1217,In_2943);
or U431 (N_431,In_1647,In_261);
nor U432 (N_432,In_2824,In_170);
or U433 (N_433,In_231,In_41);
xor U434 (N_434,In_1310,In_1182);
or U435 (N_435,In_1435,In_2214);
nor U436 (N_436,In_2,In_163);
or U437 (N_437,In_2338,In_271);
xnor U438 (N_438,In_2590,In_622);
xnor U439 (N_439,In_2546,In_2673);
and U440 (N_440,In_1510,In_2216);
and U441 (N_441,In_1675,In_803);
nor U442 (N_442,In_1863,In_2047);
or U443 (N_443,In_1020,In_340);
xor U444 (N_444,In_71,In_1398);
nor U445 (N_445,In_2468,In_1849);
or U446 (N_446,In_1599,In_2982);
and U447 (N_447,In_2483,In_1406);
nand U448 (N_448,In_1088,In_2979);
nor U449 (N_449,In_1872,In_702);
xor U450 (N_450,In_108,In_181);
and U451 (N_451,In_1987,In_923);
and U452 (N_452,In_819,In_1032);
and U453 (N_453,In_1408,In_863);
and U454 (N_454,In_1204,In_2823);
and U455 (N_455,In_354,In_607);
or U456 (N_456,In_2579,In_784);
xnor U457 (N_457,In_1755,In_1620);
nand U458 (N_458,In_932,In_2561);
and U459 (N_459,In_675,In_2156);
nor U460 (N_460,In_859,In_2478);
or U461 (N_461,In_1397,In_398);
xnor U462 (N_462,In_2562,In_1657);
nand U463 (N_463,In_423,In_2902);
and U464 (N_464,In_2470,In_1645);
nand U465 (N_465,In_1227,In_2157);
nor U466 (N_466,In_1932,In_1323);
nand U467 (N_467,In_203,In_2346);
nand U468 (N_468,In_1140,In_811);
and U469 (N_469,In_2420,In_2858);
or U470 (N_470,In_2168,In_222);
xor U471 (N_471,In_2706,In_1728);
nor U472 (N_472,In_1601,In_1015);
nor U473 (N_473,In_2807,In_411);
and U474 (N_474,In_1963,In_1367);
nor U475 (N_475,In_1782,In_4);
xnor U476 (N_476,In_1243,In_2941);
nor U477 (N_477,In_2925,In_1154);
nand U478 (N_478,In_1553,In_1235);
xnor U479 (N_479,In_2790,In_2301);
nand U480 (N_480,In_2802,In_1390);
and U481 (N_481,In_135,In_1682);
xnor U482 (N_482,In_2433,In_1685);
nand U483 (N_483,In_1784,In_2957);
xor U484 (N_484,In_2294,In_1198);
xnor U485 (N_485,In_2278,In_1151);
and U486 (N_486,In_2796,In_2992);
xnor U487 (N_487,In_2379,In_2394);
nand U488 (N_488,In_1447,In_835);
nand U489 (N_489,In_1303,In_1364);
or U490 (N_490,In_2735,In_2732);
nor U491 (N_491,In_1910,In_575);
or U492 (N_492,In_2049,In_1240);
or U493 (N_493,In_2512,In_2449);
nor U494 (N_494,In_1008,In_2937);
nand U495 (N_495,In_252,In_764);
and U496 (N_496,In_2104,In_227);
nor U497 (N_497,In_1164,In_796);
and U498 (N_498,In_1570,In_1804);
nor U499 (N_499,In_2600,In_1218);
or U500 (N_500,In_2472,In_862);
nand U501 (N_501,In_1887,In_2871);
nor U502 (N_502,In_326,In_2291);
or U503 (N_503,In_1381,In_2224);
or U504 (N_504,In_832,In_2009);
and U505 (N_505,In_2931,In_2964);
or U506 (N_506,In_2862,In_1800);
nor U507 (N_507,In_1176,In_1592);
nand U508 (N_508,In_232,In_2650);
nor U509 (N_509,In_339,In_143);
or U510 (N_510,In_1546,In_2634);
xor U511 (N_511,In_1411,In_542);
or U512 (N_512,In_726,In_1183);
nor U513 (N_513,In_770,In_394);
nand U514 (N_514,In_424,In_79);
nor U515 (N_515,In_857,In_1826);
xnor U516 (N_516,In_1433,In_2765);
or U517 (N_517,In_1680,In_99);
xnor U518 (N_518,In_2879,In_365);
xor U519 (N_519,In_1128,In_1815);
and U520 (N_520,In_2670,In_2324);
or U521 (N_521,In_1654,In_913);
nor U522 (N_522,In_322,In_177);
nand U523 (N_523,In_2493,In_366);
and U524 (N_524,In_788,In_1626);
and U525 (N_525,In_2147,In_1799);
or U526 (N_526,In_849,In_1018);
and U527 (N_527,In_2050,In_2230);
nand U528 (N_528,In_2830,In_2500);
or U529 (N_529,In_2045,In_155);
nand U530 (N_530,In_2702,In_55);
and U531 (N_531,In_2237,In_1663);
xor U532 (N_532,In_810,In_1499);
nor U533 (N_533,In_1835,In_2437);
nand U534 (N_534,In_1801,In_52);
nand U535 (N_535,In_1596,In_890);
nand U536 (N_536,In_1709,In_962);
nand U537 (N_537,In_524,In_2256);
and U538 (N_538,In_1420,In_1710);
or U539 (N_539,In_2697,In_2063);
or U540 (N_540,In_2744,In_642);
nor U541 (N_541,In_230,In_2836);
and U542 (N_542,In_2282,In_1221);
nor U543 (N_543,In_1980,In_2714);
nor U544 (N_544,In_2415,In_956);
and U545 (N_545,In_1418,In_1202);
or U546 (N_546,In_1337,In_1776);
nand U547 (N_547,In_727,In_536);
nor U548 (N_548,In_2226,In_85);
and U549 (N_549,In_1976,In_756);
or U550 (N_550,In_443,In_1934);
and U551 (N_551,In_1896,In_346);
nand U552 (N_552,In_1186,In_2378);
nand U553 (N_553,In_2001,In_475);
and U554 (N_554,In_1772,In_2213);
nor U555 (N_555,In_2761,In_335);
xnor U556 (N_556,In_2642,In_1286);
nor U557 (N_557,In_2526,In_218);
nor U558 (N_558,In_248,In_2122);
and U559 (N_559,In_2917,In_2668);
xnor U560 (N_560,In_582,In_1953);
and U561 (N_561,In_2723,In_2820);
or U562 (N_562,In_2293,In_928);
nor U563 (N_563,In_1321,In_1421);
or U564 (N_564,In_2241,In_719);
or U565 (N_565,In_144,In_2648);
and U566 (N_566,In_1692,In_1133);
or U567 (N_567,In_2091,In_2817);
or U568 (N_568,In_1027,In_490);
and U569 (N_569,In_1276,In_1629);
nand U570 (N_570,In_1385,In_2453);
xnor U571 (N_571,In_133,In_1212);
or U572 (N_572,In_2419,In_164);
nor U573 (N_573,In_1949,In_2448);
and U574 (N_574,In_2602,In_2946);
nor U575 (N_575,In_2504,In_345);
and U576 (N_576,In_93,In_2768);
nor U577 (N_577,In_2405,In_435);
nand U578 (N_578,In_2384,In_1387);
xor U579 (N_579,In_98,In_875);
nor U580 (N_580,In_668,In_1382);
xor U581 (N_581,In_2920,In_2533);
and U582 (N_582,In_2041,In_2977);
xor U583 (N_583,In_1827,In_2447);
nor U584 (N_584,In_450,In_518);
nand U585 (N_585,In_2587,In_1765);
xor U586 (N_586,In_2330,In_2207);
xor U587 (N_587,In_747,In_2679);
nand U588 (N_588,In_244,In_689);
xnor U589 (N_589,In_1999,In_2990);
nand U590 (N_590,In_2755,In_615);
or U591 (N_591,In_2682,In_1296);
and U592 (N_592,In_111,In_2046);
xnor U593 (N_593,In_670,In_1502);
and U594 (N_594,In_2206,In_1717);
xnor U595 (N_595,In_1698,In_42);
or U596 (N_596,In_2550,In_2899);
xnor U597 (N_597,In_699,In_1780);
and U598 (N_598,In_1313,In_924);
nor U599 (N_599,In_508,In_277);
nor U600 (N_600,In_455,In_569);
nand U601 (N_601,In_942,In_1944);
nand U602 (N_602,In_528,In_1879);
and U603 (N_603,In_2724,In_2223);
or U604 (N_604,In_1668,In_1559);
xor U605 (N_605,In_2380,In_1309);
or U606 (N_606,In_2647,In_2686);
nor U607 (N_607,In_2235,In_1041);
xnor U608 (N_608,In_2664,In_1677);
nor U609 (N_609,In_2994,In_2025);
or U610 (N_610,In_1936,In_2110);
or U611 (N_611,In_1189,In_1855);
and U612 (N_612,In_1617,In_841);
or U613 (N_613,In_776,In_2729);
nand U614 (N_614,In_983,In_1810);
and U615 (N_615,In_2052,In_812);
nand U616 (N_616,In_1611,In_914);
nand U617 (N_617,In_1403,In_2217);
xor U618 (N_618,In_677,In_1181);
or U619 (N_619,In_1305,In_1102);
or U620 (N_620,In_572,In_714);
xnor U621 (N_621,In_2154,In_2846);
xor U622 (N_622,In_331,In_1190);
xor U623 (N_623,In_2462,In_2385);
nand U624 (N_624,In_2296,In_1119);
or U625 (N_625,In_463,In_994);
and U626 (N_626,In_2618,In_284);
xor U627 (N_627,In_1967,In_363);
nor U628 (N_628,In_479,In_1627);
and U629 (N_629,In_717,In_2185);
nand U630 (N_630,In_907,In_432);
or U631 (N_631,In_1476,In_30);
or U632 (N_632,In_2388,In_2408);
xor U633 (N_633,In_666,In_813);
and U634 (N_634,In_1805,In_1646);
and U635 (N_635,In_613,In_338);
or U636 (N_636,In_1269,In_243);
nor U637 (N_637,In_1878,In_1490);
xnor U638 (N_638,In_2427,In_682);
nor U639 (N_639,In_2536,In_147);
and U640 (N_640,In_2490,In_467);
nor U641 (N_641,In_2720,In_958);
or U642 (N_642,In_1785,In_1016);
nor U643 (N_643,In_1958,In_1137);
or U644 (N_644,In_1636,In_1686);
nor U645 (N_645,In_578,In_67);
xnor U646 (N_646,In_1258,In_1066);
nand U647 (N_647,In_2745,In_2636);
xor U648 (N_648,In_1508,In_1346);
nand U649 (N_649,In_2869,In_2667);
nand U650 (N_650,In_2880,In_399);
and U651 (N_651,In_1315,In_1148);
and U652 (N_652,In_217,In_1033);
xnor U653 (N_653,In_2730,In_313);
or U654 (N_654,In_168,In_2196);
nor U655 (N_655,In_1173,In_2520);
nor U656 (N_656,In_1471,In_1586);
xnor U657 (N_657,In_530,In_874);
and U658 (N_658,In_1667,In_470);
nand U659 (N_659,In_2855,In_1633);
or U660 (N_660,In_2692,In_2944);
nand U661 (N_661,In_868,In_2988);
nor U662 (N_662,In_927,In_1564);
nand U663 (N_663,In_2407,In_1500);
nand U664 (N_664,In_2996,In_2436);
xnor U665 (N_665,In_349,In_2541);
or U666 (N_666,In_750,In_2798);
and U667 (N_667,In_1096,In_2444);
nand U668 (N_668,In_2124,In_2821);
and U669 (N_669,In_1693,In_2477);
and U670 (N_670,In_842,In_276);
nor U671 (N_671,In_356,In_493);
or U672 (N_672,In_1384,In_2938);
xor U673 (N_673,In_2297,In_2285);
and U674 (N_674,In_1991,In_1307);
xnor U675 (N_675,In_116,In_2510);
xor U676 (N_676,In_746,In_2929);
nor U677 (N_677,In_991,In_2967);
nand U678 (N_678,In_2894,In_70);
and U679 (N_679,In_2315,In_894);
or U680 (N_680,In_1881,In_2488);
or U681 (N_681,In_1049,In_1969);
or U682 (N_682,In_1744,In_74);
and U683 (N_683,In_1326,In_2945);
or U684 (N_684,In_2465,In_1319);
nand U685 (N_685,In_1850,In_840);
xor U686 (N_686,In_953,In_125);
and U687 (N_687,In_1787,In_669);
xor U688 (N_688,In_777,In_14);
xor U689 (N_689,In_1287,In_707);
nor U690 (N_690,In_1156,In_816);
nand U691 (N_691,In_1506,In_35);
or U692 (N_692,In_5,In_396);
or U693 (N_693,In_2464,In_1922);
or U694 (N_694,In_2635,In_2751);
or U695 (N_695,In_1774,In_86);
xor U696 (N_696,In_2661,In_1974);
nand U697 (N_697,In_272,In_1197);
nor U698 (N_698,In_526,In_1811);
nor U699 (N_699,In_567,In_710);
nand U700 (N_700,In_617,In_327);
nor U701 (N_701,In_2811,In_1533);
nor U702 (N_702,In_1901,In_2044);
nor U703 (N_703,In_1866,In_1625);
and U704 (N_704,In_1149,In_1455);
or U705 (N_705,In_2024,In_457);
or U706 (N_706,In_2169,In_62);
or U707 (N_707,In_2594,In_294);
or U708 (N_708,In_2617,In_2440);
nand U709 (N_709,In_674,In_1652);
nor U710 (N_710,In_2812,In_212);
nor U711 (N_711,In_1544,In_505);
nand U712 (N_712,In_897,In_430);
or U713 (N_713,In_2190,In_574);
nand U714 (N_714,In_2519,In_26);
nor U715 (N_715,In_2787,In_2071);
and U716 (N_716,In_774,In_2489);
and U717 (N_717,In_2874,In_1230);
and U718 (N_718,In_1971,In_2829);
nor U719 (N_719,In_2501,In_1853);
nor U720 (N_720,In_676,In_1268);
or U721 (N_721,In_517,In_1623);
nor U722 (N_722,In_1228,In_2396);
and U723 (N_723,In_1885,In_624);
and U724 (N_724,In_1573,In_1689);
nand U725 (N_725,In_1013,In_2655);
or U726 (N_726,In_2517,In_188);
or U727 (N_727,In_1393,In_1621);
and U728 (N_728,In_1973,In_216);
xor U729 (N_729,In_1748,In_2252);
nand U730 (N_730,In_1116,In_1376);
or U731 (N_731,In_2028,In_1624);
or U732 (N_732,In_2370,In_576);
nor U733 (N_733,In_1842,In_2165);
and U734 (N_734,In_1077,In_1360);
nor U735 (N_735,In_1530,In_2614);
xor U736 (N_736,In_2399,In_2261);
or U737 (N_737,In_2678,In_2675);
nor U738 (N_738,In_2860,In_1856);
nand U739 (N_739,In_1459,In_2004);
nand U740 (N_740,In_2067,In_2423);
or U741 (N_741,In_1280,In_2509);
and U742 (N_742,In_2508,In_214);
or U743 (N_743,In_2580,In_686);
and U744 (N_744,In_1029,In_368);
nand U745 (N_745,In_344,In_379);
nand U746 (N_746,In_1241,In_2058);
xor U747 (N_747,In_2215,In_1697);
or U748 (N_748,In_1368,In_797);
xor U749 (N_749,In_359,In_511);
or U750 (N_750,In_1930,In_1575);
nor U751 (N_751,In_2057,In_640);
nand U752 (N_752,In_1588,In_2400);
nand U753 (N_753,In_2619,In_2166);
xor U754 (N_754,In_2628,In_104);
and U755 (N_755,In_748,In_2348);
and U756 (N_756,In_1068,In_568);
nor U757 (N_757,In_865,In_2954);
and U758 (N_758,In_546,In_992);
nand U759 (N_759,In_1946,In_2167);
and U760 (N_760,In_1213,In_477);
nand U761 (N_761,In_332,In_2930);
xnor U762 (N_762,In_1087,In_2310);
or U763 (N_763,In_1061,In_766);
and U764 (N_764,In_798,In_2566);
xor U765 (N_765,In_1979,In_685);
nor U766 (N_766,In_2993,In_2459);
xor U767 (N_767,In_38,In_64);
or U768 (N_768,In_2708,In_1703);
or U769 (N_769,In_2204,In_499);
or U770 (N_770,In_2553,In_2528);
and U771 (N_771,In_219,In_603);
and U772 (N_772,In_2254,In_2195);
xor U773 (N_773,In_1690,In_1535);
nand U774 (N_774,In_1600,In_2480);
xor U775 (N_775,In_426,In_31);
nand U776 (N_776,In_1756,In_2547);
and U777 (N_777,In_92,In_416);
and U778 (N_778,In_2633,In_996);
or U779 (N_779,In_2418,In_1122);
xor U780 (N_780,In_2995,In_317);
xor U781 (N_781,In_2082,In_2560);
nor U782 (N_782,In_105,In_1369);
or U783 (N_783,In_2079,In_2395);
nand U784 (N_784,In_2118,In_2053);
xor U785 (N_785,In_1699,In_391);
or U786 (N_786,In_2376,In_373);
or U787 (N_787,In_1696,In_1807);
nand U788 (N_788,In_2725,In_2845);
or U789 (N_789,In_902,In_194);
xor U790 (N_790,In_2137,In_1005);
nor U791 (N_791,In_1081,In_2981);
nand U792 (N_792,In_2255,In_1023);
xnor U793 (N_793,In_131,In_442);
or U794 (N_794,In_2368,In_433);
nand U795 (N_795,In_829,In_1437);
nand U796 (N_796,In_509,In_1723);
nand U797 (N_797,In_550,In_2767);
nor U798 (N_798,In_2693,In_413);
xor U799 (N_799,In_2030,In_201);
nor U800 (N_800,In_948,In_801);
nor U801 (N_801,In_2085,In_2428);
nor U802 (N_802,In_510,In_1579);
and U803 (N_803,In_2239,In_2187);
and U804 (N_804,In_2389,In_1019);
nand U805 (N_805,In_976,In_1298);
or U806 (N_806,In_1920,In_2212);
or U807 (N_807,In_2660,In_1074);
and U808 (N_808,In_2895,In_2800);
and U809 (N_809,In_128,In_2128);
xor U810 (N_810,In_1472,In_2556);
nor U811 (N_811,In_2913,In_2332);
nor U812 (N_812,In_1740,In_2922);
nand U813 (N_813,In_500,In_281);
or U814 (N_814,In_2054,In_2949);
nand U815 (N_815,In_1113,In_938);
nor U816 (N_816,In_440,In_2527);
or U817 (N_817,In_1121,In_1821);
nor U818 (N_818,In_627,In_725);
nand U819 (N_819,In_2987,In_253);
nand U820 (N_820,In_1282,In_993);
and U821 (N_821,In_589,In_2262);
and U822 (N_822,In_407,In_2473);
nand U823 (N_823,In_497,In_2181);
nand U824 (N_824,In_1724,In_2401);
nor U825 (N_825,In_2782,In_2100);
and U826 (N_826,In_2381,In_1006);
nor U827 (N_827,In_839,In_2284);
and U828 (N_828,In_2386,In_287);
nor U829 (N_829,In_1711,In_1889);
or U830 (N_830,In_654,In_1316);
and U831 (N_831,In_1562,In_1025);
nor U832 (N_832,In_1054,In_693);
and U833 (N_833,In_806,In_564);
xnor U834 (N_834,In_1036,In_348);
or U835 (N_835,In_90,In_1110);
nor U836 (N_836,In_2074,In_2119);
xnor U837 (N_837,In_579,In_459);
nor U838 (N_838,In_2243,In_2935);
or U839 (N_839,In_660,In_2888);
or U840 (N_840,In_1779,In_2662);
nand U841 (N_841,In_101,In_80);
or U842 (N_842,In_760,In_2822);
nor U843 (N_843,In_1195,In_2352);
and U844 (N_844,In_445,In_1331);
or U845 (N_845,In_1706,In_713);
and U846 (N_846,In_1144,In_723);
nand U847 (N_847,In_2904,In_2731);
xnor U848 (N_848,In_2828,In_1877);
nand U849 (N_849,In_2061,In_965);
nor U850 (N_850,In_2503,In_1705);
nand U851 (N_851,In_1714,In_66);
or U852 (N_852,In_2966,In_1004);
or U853 (N_853,In_2424,In_2685);
xor U854 (N_854,In_1640,In_1059);
or U855 (N_855,In_759,In_856);
or U856 (N_856,In_1770,In_1529);
nand U857 (N_857,In_1741,In_197);
xnor U858 (N_858,In_302,In_1867);
nor U859 (N_859,In_1995,In_1895);
nand U860 (N_860,In_891,In_487);
and U861 (N_861,In_63,In_245);
nand U862 (N_862,In_2792,In_321);
nor U863 (N_863,In_732,In_1678);
nand U864 (N_864,In_117,In_751);
nand U865 (N_865,In_2733,In_173);
or U866 (N_866,In_2273,In_916);
nand U867 (N_867,In_24,In_1424);
and U868 (N_868,In_119,In_282);
and U869 (N_869,In_1549,In_2893);
nand U870 (N_870,In_1938,In_1606);
nand U871 (N_871,In_663,In_486);
nor U872 (N_872,In_2643,In_782);
nand U873 (N_873,In_2712,In_619);
nand U874 (N_874,In_1583,In_2583);
nand U875 (N_875,In_1760,In_1120);
xor U876 (N_876,In_597,In_905);
nand U877 (N_877,In_375,In_383);
nor U878 (N_878,In_2622,In_2898);
nand U879 (N_879,In_2034,In_2200);
nor U880 (N_880,In_1673,In_32);
or U881 (N_881,In_1852,In_1180);
and U882 (N_882,In_198,In_2518);
or U883 (N_883,In_559,In_10);
nor U884 (N_884,In_2271,In_1808);
and U885 (N_885,In_931,In_1214);
nor U886 (N_886,In_2644,In_804);
or U887 (N_887,In_2115,In_2511);
or U888 (N_888,In_1052,In_160);
nor U889 (N_889,In_1761,In_2911);
and U890 (N_890,In_2410,In_466);
nand U891 (N_891,In_2253,In_1238);
and U892 (N_892,In_2438,In_1638);
or U893 (N_893,In_985,In_1401);
xnor U894 (N_894,In_1207,In_623);
xnor U895 (N_895,In_61,In_2507);
nor U896 (N_896,In_1216,In_743);
xor U897 (N_897,In_1733,In_1605);
xor U898 (N_898,In_2709,In_1359);
or U899 (N_899,In_1580,In_2710);
nor U900 (N_900,In_1067,In_192);
or U901 (N_901,In_1970,In_1351);
xor U902 (N_902,In_481,In_545);
xnor U903 (N_903,In_1674,In_1124);
and U904 (N_904,In_250,In_2102);
nor U905 (N_905,In_1171,In_2355);
or U906 (N_906,In_2831,In_2007);
or U907 (N_907,In_370,In_535);
or U908 (N_908,In_1084,In_2851);
xor U909 (N_909,In_1961,In_1912);
nor U910 (N_910,In_2684,In_2246);
and U911 (N_911,In_1942,In_2707);
or U912 (N_912,In_1245,In_2582);
or U913 (N_913,In_1279,In_551);
xor U914 (N_914,In_1847,In_1794);
or U915 (N_915,In_2759,In_484);
xnor U916 (N_916,In_2564,In_1372);
or U917 (N_917,In_298,In_37);
or U918 (N_918,In_1727,In_920);
or U919 (N_919,In_2177,In_1248);
or U920 (N_920,In_2866,In_1297);
xnor U921 (N_921,In_1085,In_1294);
xor U922 (N_922,In_737,In_1496);
and U923 (N_923,In_211,In_2687);
and U924 (N_924,In_1484,In_2374);
nand U925 (N_925,In_562,In_1452);
and U926 (N_926,In_1577,In_2197);
xor U927 (N_927,In_2656,In_12);
or U928 (N_928,In_129,In_709);
and U929 (N_929,In_988,In_2461);
or U930 (N_930,In_2885,In_1395);
or U931 (N_931,In_2055,In_23);
or U932 (N_932,In_1904,In_290);
or U933 (N_933,In_2179,In_57);
nor U934 (N_934,In_1242,In_2145);
and U935 (N_935,In_446,In_274);
nor U936 (N_936,In_2013,In_2029);
xor U937 (N_937,In_864,In_802);
nor U938 (N_938,In_2882,In_893);
or U939 (N_939,In_972,In_658);
xor U940 (N_940,In_115,In_2916);
nor U941 (N_941,In_2298,In_2538);
nor U942 (N_942,In_2456,In_2927);
nor U943 (N_943,In_749,In_421);
nor U944 (N_944,In_1616,In_989);
or U945 (N_945,In_2012,In_2909);
nand U946 (N_946,In_1247,In_2786);
xor U947 (N_947,In_618,In_1026);
and U948 (N_948,In_2539,In_982);
or U949 (N_949,In_580,In_861);
xor U950 (N_950,In_1587,In_1843);
and U951 (N_951,In_688,In_1483);
nor U952 (N_952,In_1603,In_805);
or U953 (N_953,In_2377,In_1399);
or U954 (N_954,In_1649,In_786);
xnor U955 (N_955,In_2129,In_2889);
nand U956 (N_956,In_2631,In_2805);
xnor U957 (N_957,In_2713,In_377);
xnor U958 (N_958,In_543,In_2397);
and U959 (N_959,In_1613,In_2932);
nand U960 (N_960,In_706,In_2150);
or U961 (N_961,In_2441,In_1226);
or U962 (N_962,In_744,In_1505);
and U963 (N_963,In_794,In_1065);
and U964 (N_964,In_142,In_637);
and U965 (N_965,In_1643,In_590);
or U966 (N_966,In_778,In_388);
nor U967 (N_967,In_1593,In_2109);
or U968 (N_968,In_1125,In_2443);
nand U969 (N_969,In_1982,In_1051);
nand U970 (N_970,In_2775,In_382);
and U971 (N_971,In_77,In_238);
nand U972 (N_972,In_599,In_1017);
and U973 (N_973,In_157,In_2985);
nand U974 (N_974,In_692,In_1845);
or U975 (N_975,In_436,In_2884);
nor U976 (N_976,In_697,In_1342);
or U977 (N_977,In_2039,In_1463);
and U978 (N_978,In_199,In_683);
nor U979 (N_979,In_2738,In_2565);
xor U980 (N_980,In_1732,In_1229);
xnor U981 (N_981,In_229,In_1336);
nand U982 (N_982,In_984,In_2277);
or U983 (N_983,In_2172,In_9);
and U984 (N_984,In_2699,In_2242);
xor U985 (N_985,In_799,In_11);
and U986 (N_986,In_308,In_636);
nand U987 (N_987,In_152,In_1117);
or U988 (N_988,In_2065,In_1557);
nand U989 (N_989,In_2414,In_1007);
nor U990 (N_990,In_2752,In_2121);
and U991 (N_991,In_1841,In_1766);
and U992 (N_992,In_2323,In_941);
nor U993 (N_993,In_262,In_1702);
xor U994 (N_994,In_652,In_2373);
and U995 (N_995,In_1781,In_478);
and U996 (N_996,In_1306,In_2080);
nor U997 (N_997,In_58,In_2015);
nand U998 (N_998,In_1262,In_2267);
xnor U999 (N_999,In_1055,In_2942);
and U1000 (N_1000,In_2502,In_166);
and U1001 (N_1001,In_2700,In_534);
nor U1002 (N_1002,In_527,In_2132);
nand U1003 (N_1003,In_371,In_1555);
and U1004 (N_1004,In_790,In_2797);
xor U1005 (N_1005,In_973,In_174);
nand U1006 (N_1006,In_934,In_2890);
and U1007 (N_1007,In_964,In_2228);
nor U1008 (N_1008,In_140,In_1594);
and U1009 (N_1009,In_1978,In_873);
and U1010 (N_1010,In_1299,In_44);
nand U1011 (N_1011,In_1284,In_2300);
nand U1012 (N_1012,In_2090,In_2467);
or U1013 (N_1013,In_2962,In_1707);
xor U1014 (N_1014,In_1955,In_1665);
or U1015 (N_1015,In_2006,In_2426);
or U1016 (N_1016,In_2155,In_1266);
or U1017 (N_1017,In_1131,In_27);
or U1018 (N_1018,In_221,In_357);
xor U1019 (N_1019,In_2404,In_647);
nor U1020 (N_1020,In_121,In_409);
and U1021 (N_1021,In_1767,In_1547);
xor U1022 (N_1022,In_1419,In_1177);
and U1023 (N_1023,In_2813,In_733);
and U1024 (N_1024,In_88,In_1947);
nor U1025 (N_1025,In_937,In_591);
nor U1026 (N_1026,In_1060,In_525);
or U1027 (N_1027,In_1731,In_2064);
nand U1028 (N_1028,In_1219,In_596);
or U1029 (N_1029,In_2868,In_2313);
and U1030 (N_1030,In_2595,In_137);
and U1031 (N_1031,In_533,In_1839);
nand U1032 (N_1032,In_911,In_2632);
nor U1033 (N_1033,In_633,In_246);
nor U1034 (N_1034,In_950,In_2411);
nor U1035 (N_1035,In_2430,In_2763);
xnor U1036 (N_1036,In_2289,In_1793);
nor U1037 (N_1037,In_1662,In_1021);
nor U1038 (N_1038,In_1091,In_1829);
nand U1039 (N_1039,In_1911,In_2409);
xnor U1040 (N_1040,In_431,In_1897);
nand U1041 (N_1041,In_846,In_2577);
nor U1042 (N_1042,In_259,In_671);
and U1043 (N_1043,In_1175,In_1324);
or U1044 (N_1044,In_2451,In_2840);
or U1045 (N_1045,In_2335,In_1256);
or U1046 (N_1046,In_1528,In_1278);
nand U1047 (N_1047,In_858,In_2532);
nand U1048 (N_1048,In_1093,In_1366);
nor U1049 (N_1049,In_2321,In_629);
nor U1050 (N_1050,In_1482,In_1349);
xnor U1051 (N_1051,In_601,In_1464);
nand U1052 (N_1052,In_1078,In_892);
or U1053 (N_1053,In_736,In_151);
nor U1054 (N_1054,In_2276,In_2567);
nor U1055 (N_1055,In_971,In_2952);
nand U1056 (N_1056,In_102,In_1264);
nor U1057 (N_1057,In_1352,In_1290);
xor U1058 (N_1058,In_1522,In_1532);
and U1059 (N_1059,In_1915,In_2680);
xnor U1060 (N_1060,In_1726,In_165);
or U1061 (N_1061,In_1333,In_465);
and U1062 (N_1062,In_456,In_1141);
xor U1063 (N_1063,In_2554,In_828);
xor U1064 (N_1064,In_488,In_2857);
nand U1065 (N_1065,In_2008,In_2076);
nand U1066 (N_1066,In_59,In_850);
nand U1067 (N_1067,In_297,In_912);
or U1068 (N_1068,In_1139,In_2343);
and U1069 (N_1069,In_1073,In_1609);
nor U1070 (N_1070,In_78,In_114);
xnor U1071 (N_1071,In_1859,In_489);
nor U1072 (N_1072,In_967,In_1998);
or U1073 (N_1073,In_1739,In_402);
nor U1074 (N_1074,In_2575,In_215);
nand U1075 (N_1075,In_325,In_2613);
nand U1076 (N_1076,In_2327,In_1509);
or U1077 (N_1077,In_2747,In_1152);
nor U1078 (N_1078,In_818,In_1960);
and U1079 (N_1079,In_504,In_1361);
nor U1080 (N_1080,In_401,In_2758);
and U1081 (N_1081,In_2691,In_2413);
nor U1082 (N_1082,In_644,In_1683);
xor U1083 (N_1083,In_2726,In_352);
or U1084 (N_1084,In_2434,In_2286);
xor U1085 (N_1085,In_2136,In_823);
or U1086 (N_1086,In_986,In_1317);
nand U1087 (N_1087,In_1427,In_1597);
xor U1088 (N_1088,In_833,In_439);
nor U1089 (N_1089,In_522,In_2072);
nor U1090 (N_1090,In_2815,In_2188);
or U1091 (N_1091,In_213,In_2690);
and U1092 (N_1092,In_2069,In_498);
xor U1093 (N_1093,In_595,In_2659);
nand U1094 (N_1094,In_2032,In_1423);
and U1095 (N_1095,In_852,In_1479);
xor U1096 (N_1096,In_2727,In_1179);
xor U1097 (N_1097,In_2534,In_1070);
nor U1098 (N_1098,In_2314,In_544);
or U1099 (N_1099,In_2018,In_1876);
nand U1100 (N_1100,In_1631,In_621);
or U1101 (N_1101,In_2229,In_1142);
and U1102 (N_1102,In_1105,In_1729);
or U1103 (N_1103,In_1582,In_2974);
xor U1104 (N_1104,In_2345,In_1701);
nand U1105 (N_1105,In_1453,In_1865);
or U1106 (N_1106,In_2825,In_1391);
nor U1107 (N_1107,In_2455,In_772);
nand U1108 (N_1108,In_15,In_2113);
and U1109 (N_1109,In_2479,In_1561);
xnor U1110 (N_1110,In_1615,In_561);
and U1111 (N_1111,In_2865,In_2535);
nor U1112 (N_1112,In_2906,In_2672);
and U1113 (N_1113,In_2307,In_2250);
nor U1114 (N_1114,In_1542,In_2606);
nor U1115 (N_1115,In_1330,In_2588);
and U1116 (N_1116,In_1192,In_2804);
and U1117 (N_1117,In_1762,In_1870);
and U1118 (N_1118,In_780,In_678);
or U1119 (N_1119,In_1355,In_2870);
nand U1120 (N_1120,In_2222,In_301);
nand U1121 (N_1121,In_1292,In_2903);
xnor U1122 (N_1122,In_1737,In_2695);
or U1123 (N_1123,In_2342,In_869);
nor U1124 (N_1124,In_1341,In_843);
or U1125 (N_1125,In_1764,In_611);
nor U1126 (N_1126,In_2969,In_1037);
nor U1127 (N_1127,In_1076,In_592);
or U1128 (N_1128,In_625,In_2482);
and U1129 (N_1129,In_1132,In_1824);
or U1130 (N_1130,In_1789,In_1909);
or U1131 (N_1131,In_560,In_1935);
xnor U1132 (N_1132,In_1208,In_2934);
or U1133 (N_1133,In_2295,In_414);
and U1134 (N_1134,In_2099,In_1462);
and U1135 (N_1135,In_1328,In_2624);
and U1136 (N_1136,In_1671,In_2259);
nor U1137 (N_1137,In_429,In_1567);
and U1138 (N_1138,In_2834,In_2722);
or U1139 (N_1139,In_1354,In_2892);
or U1140 (N_1140,In_1899,In_877);
nand U1141 (N_1141,In_204,In_2481);
nand U1142 (N_1142,In_795,In_910);
and U1143 (N_1143,In_266,In_444);
nand U1144 (N_1144,In_1044,In_1653);
or U1145 (N_1145,In_343,In_2130);
or U1146 (N_1146,In_1788,In_2248);
and U1147 (N_1147,In_2806,In_2531);
nor U1148 (N_1148,In_2193,In_769);
or U1149 (N_1149,In_896,In_126);
xnor U1150 (N_1150,In_319,In_2021);
xnor U1151 (N_1151,In_1375,In_1146);
or U1152 (N_1152,In_995,In_1560);
and U1153 (N_1153,In_1908,In_2406);
or U1154 (N_1154,In_754,In_146);
xnor U1155 (N_1155,In_2143,In_2033);
nand U1156 (N_1156,In_2031,In_966);
xnor U1157 (N_1157,In_171,In_1089);
xor U1158 (N_1158,In_2791,In_1244);
and U1159 (N_1159,In_464,In_2803);
and U1160 (N_1160,In_273,In_2900);
and U1161 (N_1161,In_2322,In_1035);
or U1162 (N_1162,In_2601,In_1318);
and U1163 (N_1163,In_1660,In_834);
nand U1164 (N_1164,In_2681,In_1669);
xor U1165 (N_1165,In_1521,In_1996);
or U1166 (N_1166,In_1892,In_2525);
nor U1167 (N_1167,In_1130,In_1222);
or U1168 (N_1168,In_1639,In_929);
or U1169 (N_1169,In_2610,In_158);
xor U1170 (N_1170,In_2948,In_1554);
xnor U1171 (N_1171,In_880,In_1038);
nand U1172 (N_1172,In_2671,In_2973);
nand U1173 (N_1173,In_520,In_1681);
xnor U1174 (N_1174,In_1002,In_2268);
and U1175 (N_1175,In_122,In_2753);
xnor U1176 (N_1176,In_1046,In_1905);
nor U1177 (N_1177,In_458,In_1641);
nand U1178 (N_1178,In_417,In_2848);
nand U1179 (N_1179,In_2153,In_883);
nand U1180 (N_1180,In_1339,In_2569);
and U1181 (N_1181,In_1548,In_2037);
and U1182 (N_1182,In_1721,In_2005);
xnor U1183 (N_1183,In_1981,In_2881);
xor U1184 (N_1184,In_1414,In_1563);
nand U1185 (N_1185,In_1444,In_2652);
or U1186 (N_1186,In_2059,In_2559);
nor U1187 (N_1187,In_1428,In_1486);
nor U1188 (N_1188,In_2240,In_161);
nand U1189 (N_1189,In_2491,In_2832);
or U1190 (N_1190,In_1111,In_47);
nor U1191 (N_1191,In_752,In_2780);
nand U1192 (N_1192,In_959,In_1010);
and U1193 (N_1193,In_2494,In_2592);
nor U1194 (N_1194,In_2349,In_2769);
or U1195 (N_1195,In_1058,In_2997);
nor U1196 (N_1196,In_1448,In_2233);
nor U1197 (N_1197,In_2087,In_1538);
nand U1198 (N_1198,In_2853,In_2958);
nor U1199 (N_1199,In_1425,In_13);
and U1200 (N_1200,N_190,N_1096);
xor U1201 (N_1201,N_1105,N_79);
xor U1202 (N_1202,N_1186,In_196);
xnor U1203 (N_1203,In_2663,In_949);
or U1204 (N_1204,N_8,N_659);
xnor U1205 (N_1205,N_945,N_337);
or U1206 (N_1206,N_960,N_983);
and U1207 (N_1207,In_186,N_693);
nand U1208 (N_1208,N_146,N_1023);
nor U1209 (N_1209,In_1166,In_2111);
or U1210 (N_1210,In_2287,N_1199);
and U1211 (N_1211,N_1028,N_1181);
or U1212 (N_1212,N_631,N_541);
nor U1213 (N_1213,N_501,N_237);
xnor U1214 (N_1214,N_1165,N_923);
or U1215 (N_1215,N_788,N_707);
and U1216 (N_1216,N_17,In_554);
and U1217 (N_1217,In_2669,N_76);
or U1218 (N_1218,N_1106,In_1759);
or U1219 (N_1219,N_1018,In_2351);
or U1220 (N_1220,In_1404,N_151);
and U1221 (N_1221,N_331,N_360);
or U1222 (N_1222,N_1097,N_307);
xor U1223 (N_1223,N_534,N_253);
and U1224 (N_1224,N_56,N_1076);
nand U1225 (N_1225,N_235,In_2151);
nor U1226 (N_1226,N_830,In_516);
nor U1227 (N_1227,N_792,N_979);
nand U1228 (N_1228,N_464,In_1628);
xor U1229 (N_1229,N_1126,N_268);
nand U1230 (N_1230,N_1147,N_269);
and U1231 (N_1231,N_572,N_385);
nor U1232 (N_1232,N_343,In_2608);
or U1233 (N_1233,N_84,N_1170);
xor U1234 (N_1234,N_378,In_2326);
nor U1235 (N_1235,In_2666,In_1687);
nand U1236 (N_1236,N_611,N_581);
or U1237 (N_1237,N_548,In_300);
and U1238 (N_1238,N_388,N_1145);
and U1239 (N_1239,N_398,N_74);
and U1240 (N_1240,N_1090,In_1295);
or U1241 (N_1241,In_605,N_1166);
nor U1242 (N_1242,In_2746,In_1356);
xor U1243 (N_1243,In_1431,N_1152);
xnor U1244 (N_1244,N_699,N_95);
nand U1245 (N_1245,In_2281,N_556);
nand U1246 (N_1246,N_896,N_841);
and U1247 (N_1247,N_83,N_905);
nor U1248 (N_1248,N_472,N_1007);
or U1249 (N_1249,In_765,N_174);
nand U1250 (N_1250,N_758,N_374);
and U1251 (N_1251,N_951,N_1047);
nor U1252 (N_1252,In_2139,N_149);
and U1253 (N_1253,In_1700,N_1192);
nor U1254 (N_1254,In_1795,In_193);
xor U1255 (N_1255,N_932,In_2499);
xor U1256 (N_1256,In_974,N_32);
and U1257 (N_1257,N_117,N_296);
nand U1258 (N_1258,N_132,In_1552);
nand U1259 (N_1259,N_255,In_73);
xnor U1260 (N_1260,N_805,N_831);
xor U1261 (N_1261,In_1252,N_716);
xor U1262 (N_1262,N_958,N_94);
nor U1263 (N_1263,In_2458,N_516);
and U1264 (N_1264,N_802,In_2017);
nand U1265 (N_1265,In_1312,N_537);
or U1266 (N_1266,N_764,N_20);
nand U1267 (N_1267,N_1034,N_876);
and U1268 (N_1268,N_463,N_1098);
and U1269 (N_1269,N_785,N_260);
and U1270 (N_1270,N_383,N_929);
nor U1271 (N_1271,N_1189,N_419);
or U1272 (N_1272,N_955,In_1199);
and U1273 (N_1273,In_724,N_1087);
and U1274 (N_1274,N_6,In_1188);
nor U1275 (N_1275,In_673,N_1177);
and U1276 (N_1276,N_1021,N_523);
xor U1277 (N_1277,N_191,N_63);
nand U1278 (N_1278,In_1715,N_489);
nand U1279 (N_1279,N_925,N_288);
and U1280 (N_1280,N_1038,N_23);
nand U1281 (N_1281,N_1048,In_634);
nor U1282 (N_1282,N_50,N_382);
nand U1283 (N_1283,N_563,N_1154);
or U1284 (N_1284,In_1798,In_2257);
nor U1285 (N_1285,N_1141,In_1917);
nor U1286 (N_1286,In_2616,In_2737);
nand U1287 (N_1287,N_601,N_427);
xor U1288 (N_1288,In_1263,N_47);
xnor U1289 (N_1289,In_1325,In_690);
nand U1290 (N_1290,N_11,In_2382);
nor U1291 (N_1291,N_927,N_1000);
nor U1292 (N_1292,N_543,N_302);
nor U1293 (N_1293,In_1984,In_1485);
and U1294 (N_1294,N_811,N_970);
nor U1295 (N_1295,N_171,N_594);
xnor U1296 (N_1296,N_946,In_975);
nand U1297 (N_1297,In_1454,N_1053);
xnor U1298 (N_1298,N_597,In_2959);
xnor U1299 (N_1299,N_506,N_1131);
or U1300 (N_1300,N_1022,N_387);
or U1301 (N_1301,In_2505,N_647);
and U1302 (N_1302,N_717,N_100);
nand U1303 (N_1303,N_477,N_106);
and U1304 (N_1304,In_1610,N_613);
xnor U1305 (N_1305,In_2849,N_849);
nor U1306 (N_1306,N_234,N_466);
nand U1307 (N_1307,N_502,In_299);
and U1308 (N_1308,N_964,In_616);
nand U1309 (N_1309,In_1749,N_790);
nand U1310 (N_1310,N_229,N_565);
xor U1311 (N_1311,In_2576,N_1171);
nand U1312 (N_1312,N_912,N_692);
or U1313 (N_1313,N_257,N_13);
and U1314 (N_1314,In_922,N_418);
and U1315 (N_1315,N_737,In_2077);
xnor U1316 (N_1316,In_2515,N_380);
and U1317 (N_1317,N_999,N_756);
nand U1318 (N_1318,N_373,N_1117);
nand U1319 (N_1319,In_925,In_2173);
or U1320 (N_1320,In_2910,N_1020);
and U1321 (N_1321,N_1058,N_180);
and U1322 (N_1322,In_162,N_454);
xnor U1323 (N_1323,N_820,In_169);
nand U1324 (N_1324,N_800,N_650);
and U1325 (N_1325,N_924,In_2719);
xor U1326 (N_1326,N_163,In_179);
and U1327 (N_1327,In_2530,In_1277);
nor U1328 (N_1328,N_511,N_573);
xnor U1329 (N_1329,N_291,In_2339);
and U1330 (N_1330,N_584,In_1475);
nand U1331 (N_1331,In_333,N_495);
and U1332 (N_1332,In_2038,N_199);
nand U1333 (N_1333,N_452,N_987);
xnor U1334 (N_1334,N_747,In_789);
nor U1335 (N_1335,N_461,In_1461);
or U1336 (N_1336,In_2279,N_1081);
nand U1337 (N_1337,N_364,N_254);
and U1338 (N_1338,In_283,In_853);
or U1339 (N_1339,N_797,N_774);
nand U1340 (N_1340,N_80,N_474);
nand U1341 (N_1341,N_730,N_177);
or U1342 (N_1342,In_364,N_204);
xor U1343 (N_1343,N_705,N_167);
or U1344 (N_1344,N_834,N_408);
xor U1345 (N_1345,N_96,N_169);
nor U1346 (N_1346,In_1451,In_1857);
nor U1347 (N_1347,N_469,N_1066);
nor U1348 (N_1348,In_1,N_904);
and U1349 (N_1349,N_1185,In_1809);
or U1350 (N_1350,In_2961,N_216);
or U1351 (N_1351,N_1110,N_1135);
and U1352 (N_1352,N_524,In_1034);
nor U1353 (N_1353,N_354,N_604);
xnor U1354 (N_1354,In_2762,In_2131);
nand U1355 (N_1355,N_950,In_1635);
nor U1356 (N_1356,N_21,N_73);
nor U1357 (N_1357,N_455,In_1672);
nor U1358 (N_1358,N_1094,N_784);
nand U1359 (N_1359,In_698,N_685);
nand U1360 (N_1360,N_921,N_60);
nor U1361 (N_1361,N_101,N_826);
or U1362 (N_1362,In_2956,N_1102);
xnor U1363 (N_1363,N_324,In_957);
and U1364 (N_1364,N_1010,N_576);
xor U1365 (N_1365,N_1003,In_1874);
and U1366 (N_1366,N_1124,N_1085);
and U1367 (N_1367,N_356,In_1745);
or U1368 (N_1368,In_731,In_314);
nand U1369 (N_1369,N_297,In_2083);
and U1370 (N_1370,N_348,N_677);
or U1371 (N_1371,N_226,In_895);
nand U1372 (N_1372,N_298,N_326);
nand U1373 (N_1373,N_1006,In_712);
nor U1374 (N_1374,N_759,In_415);
or U1375 (N_1375,In_422,In_2545);
and U1376 (N_1376,N_943,N_14);
and U1377 (N_1377,In_2772,N_1155);
or U1378 (N_1378,N_603,N_507);
nand U1379 (N_1379,N_569,In_367);
xnor U1380 (N_1380,N_1035,N_24);
or U1381 (N_1381,N_224,N_1027);
nand U1382 (N_1382,N_103,In_185);
and U1383 (N_1383,In_2827,N_273);
nand U1384 (N_1384,N_210,N_963);
xnor U1385 (N_1385,N_672,N_989);
and U1386 (N_1386,N_9,N_892);
nand U1387 (N_1387,In_2593,In_860);
or U1388 (N_1388,N_532,N_895);
xor U1389 (N_1389,N_809,N_813);
nand U1390 (N_1390,In_1712,N_858);
xnor U1391 (N_1391,N_557,In_1513);
or U1392 (N_1392,N_230,N_1093);
xnor U1393 (N_1393,N_251,N_689);
nand U1394 (N_1394,In_2275,N_766);
nor U1395 (N_1395,N_487,N_10);
nand U1396 (N_1396,N_691,N_799);
xor U1397 (N_1397,In_178,In_1158);
or U1398 (N_1398,N_649,In_718);
nand U1399 (N_1399,N_314,N_564);
nor U1400 (N_1400,In_1057,N_186);
xnor U1401 (N_1401,N_726,N_856);
nor U1402 (N_1402,In_1576,N_862);
and U1403 (N_1403,N_882,N_351);
nand U1404 (N_1404,N_357,In_438);
and U1405 (N_1405,N_984,In_2317);
nand U1406 (N_1406,N_1129,N_308);
nand U1407 (N_1407,N_345,N_709);
nand U1408 (N_1408,In_936,N_675);
nand U1409 (N_1409,N_475,N_447);
xor U1410 (N_1410,N_467,N_212);
nor U1411 (N_1411,N_12,In_1838);
and U1412 (N_1412,N_25,N_803);
nor U1413 (N_1413,N_944,N_429);
nand U1414 (N_1414,N_330,N_1089);
or U1415 (N_1415,N_341,In_1254);
or U1416 (N_1416,N_918,In_1525);
and U1417 (N_1417,In_2258,N_838);
nand U1418 (N_1418,In_2108,In_1571);
xnor U1419 (N_1419,In_506,In_1429);
and U1420 (N_1420,N_962,In_1335);
and U1421 (N_1421,In_2810,N_740);
nor U1422 (N_1422,In_2364,In_632);
nor U1423 (N_1423,N_860,N_1008);
and U1424 (N_1424,In_2442,In_650);
nand U1425 (N_1425,N_1121,In_1118);
nor U1426 (N_1426,N_61,N_656);
nand U1427 (N_1427,N_46,N_484);
or U1428 (N_1428,In_1003,In_2308);
and U1429 (N_1429,N_424,In_1094);
nor U1430 (N_1430,N_591,N_696);
and U1431 (N_1431,N_715,In_1989);
and U1432 (N_1432,In_1591,N_325);
or U1433 (N_1433,N_844,In_1746);
and U1434 (N_1434,N_562,N_1108);
xor U1435 (N_1435,N_112,In_700);
nand U1436 (N_1436,In_1956,N_434);
nor U1437 (N_1437,N_899,N_1196);
xor U1438 (N_1438,N_301,N_1);
xnor U1439 (N_1439,In_708,N_570);
nand U1440 (N_1440,In_1163,N_335);
nor U1441 (N_1441,In_1540,N_1068);
and U1442 (N_1442,In_555,N_1041);
nand U1443 (N_1443,N_33,In_1365);
or U1444 (N_1444,N_43,In_136);
or U1445 (N_1445,N_901,N_561);
and U1446 (N_1446,N_36,N_519);
or U1447 (N_1447,N_814,N_19);
nand U1448 (N_1448,N_205,N_525);
nor U1449 (N_1449,N_843,In_1578);
and U1450 (N_1450,N_1140,In_2783);
or U1451 (N_1451,In_2549,N_402);
nand U1452 (N_1452,In_2350,In_2403);
and U1453 (N_1453,N_976,N_104);
xor U1454 (N_1454,In_2144,N_93);
and U1455 (N_1455,In_2856,N_1042);
nand U1456 (N_1456,In_362,N_616);
nand U1457 (N_1457,N_289,N_718);
nor U1458 (N_1458,In_2062,N_855);
or U1459 (N_1459,In_2365,N_623);
xnor U1460 (N_1460,N_85,N_609);
and U1461 (N_1461,In_1193,N_62);
and U1462 (N_1462,N_536,N_98);
xnor U1463 (N_1463,N_92,N_1161);
nor U1464 (N_1464,N_959,In_1072);
xnor U1465 (N_1465,N_818,N_735);
or U1466 (N_1466,N_883,N_1187);
or U1467 (N_1467,N_366,N_1079);
xor U1468 (N_1468,In_1249,In_872);
nand U1469 (N_1469,In_531,In_1187);
nand U1470 (N_1470,In_2795,In_82);
nor U1471 (N_1471,N_339,N_473);
or U1472 (N_1472,N_490,N_280);
and U1473 (N_1473,N_968,N_973);
nor U1474 (N_1474,N_866,In_845);
or U1475 (N_1475,In_1442,In_2711);
and U1476 (N_1476,In_2068,N_290);
nor U1477 (N_1477,N_796,In_110);
or U1478 (N_1478,N_86,In_347);
nand U1479 (N_1479,N_767,N_219);
or U1480 (N_1480,N_369,In_1650);
or U1481 (N_1481,In_1992,In_1161);
nor U1482 (N_1482,In_2688,N_198);
xor U1483 (N_1483,In_2393,N_721);
nor U1484 (N_1484,N_54,In_2891);
and U1485 (N_1485,In_2621,N_1073);
and U1486 (N_1486,In_1923,N_589);
nand U1487 (N_1487,In_1871,N_635);
and U1488 (N_1488,N_1045,N_122);
nor U1489 (N_1489,N_530,In_570);
nor U1490 (N_1490,N_1025,N_1030);
nand U1491 (N_1491,N_403,N_399);
xnor U1492 (N_1492,N_195,N_214);
and U1493 (N_1493,N_196,N_250);
or U1494 (N_1494,N_978,N_679);
or U1495 (N_1495,N_406,N_285);
xnor U1496 (N_1496,In_2789,N_593);
and U1497 (N_1497,In_817,In_182);
or U1498 (N_1498,N_275,N_152);
xor U1499 (N_1499,N_1056,N_173);
xnor U1500 (N_1500,In_2551,N_449);
or U1501 (N_1501,N_910,N_142);
or U1502 (N_1502,N_231,In_1460);
and U1503 (N_1503,N_465,N_162);
xnor U1504 (N_1504,N_1014,In_1191);
nand U1505 (N_1505,In_889,N_851);
nor U1506 (N_1506,In_730,N_684);
or U1507 (N_1507,N_145,N_450);
nor U1508 (N_1508,In_2363,In_1136);
nor U1509 (N_1509,N_607,N_201);
and U1510 (N_1510,In_1691,N_16);
nand U1511 (N_1511,N_1061,In_316);
or U1512 (N_1512,N_299,N_215);
and U1513 (N_1513,In_1688,N_857);
nand U1514 (N_1514,N_687,N_352);
nor U1515 (N_1515,N_937,N_41);
xor U1516 (N_1516,N_1064,In_612);
and U1517 (N_1517,N_405,N_668);
or U1518 (N_1518,In_2249,N_263);
or U1519 (N_1519,N_340,N_829);
nor U1520 (N_1520,In_1534,In_1543);
or U1521 (N_1521,N_441,N_165);
nor U1522 (N_1522,N_131,N_746);
and U1523 (N_1523,N_941,In_454);
and U1524 (N_1524,N_926,N_1088);
nor U1525 (N_1525,N_942,N_850);
xnor U1526 (N_1526,N_189,In_2978);
nand U1527 (N_1527,N_517,In_502);
or U1528 (N_1528,N_713,In_1604);
nand U1529 (N_1529,N_185,N_346);
and U1530 (N_1530,N_868,N_542);
xnor U1531 (N_1531,N_706,N_821);
and U1532 (N_1532,N_267,In_2965);
and U1533 (N_1533,N_153,N_854);
and U1534 (N_1534,N_200,In_2581);
xnor U1535 (N_1535,N_550,N_1142);
nand U1536 (N_1536,N_752,N_852);
or U1537 (N_1537,N_241,N_3);
and U1538 (N_1538,N_236,N_410);
and U1539 (N_1539,In_2141,In_779);
or U1540 (N_1540,N_956,In_1990);
nor U1541 (N_1541,N_1183,N_518);
or U1542 (N_1542,In_2625,In_207);
nand U1543 (N_1543,N_900,In_2801);
nor U1544 (N_1544,N_1149,N_197);
nand U1545 (N_1545,N_438,N_1114);
or U1546 (N_1546,N_126,N_1070);
and U1547 (N_1547,In_2544,In_83);
nand U1548 (N_1548,In_1275,In_600);
xor U1549 (N_1549,N_738,In_665);
nor U1550 (N_1550,N_396,N_266);
or U1551 (N_1551,In_1752,In_885);
nand U1552 (N_1552,N_252,In_2999);
nand U1553 (N_1553,N_712,N_342);
xnor U1554 (N_1554,In_866,N_897);
xnor U1555 (N_1555,N_318,In_224);
xor U1556 (N_1556,N_634,N_328);
nand U1557 (N_1557,N_313,N_459);
xnor U1558 (N_1558,N_66,In_2819);
and U1559 (N_1559,N_771,In_425);
and U1560 (N_1560,N_1162,N_361);
nand U1561 (N_1561,In_1347,N_1082);
nand U1562 (N_1562,N_5,In_1753);
or U1563 (N_1563,In_148,In_2347);
and U1564 (N_1564,N_920,In_602);
xor U1565 (N_1565,N_903,N_140);
nand U1566 (N_1566,N_401,N_247);
xnor U1567 (N_1567,N_560,In_657);
or U1568 (N_1568,In_483,In_1622);
nor U1569 (N_1569,N_610,N_754);
and U1570 (N_1570,N_57,In_695);
nor U1571 (N_1571,In_2369,N_283);
nor U1572 (N_1572,In_2095,N_977);
nor U1573 (N_1573,N_1063,In_1407);
xnor U1574 (N_1574,N_1055,In_2446);
or U1575 (N_1575,N_683,N_178);
xnor U1576 (N_1576,In_1340,N_615);
and U1577 (N_1577,N_1104,In_472);
nor U1578 (N_1578,In_175,In_783);
xor U1579 (N_1579,In_814,N_31);
nand U1580 (N_1580,N_724,N_1122);
and U1581 (N_1581,In_940,N_779);
nor U1582 (N_1582,In_29,N_786);
or U1583 (N_1583,In_2372,N_674);
and U1584 (N_1584,In_106,N_940);
or U1585 (N_1585,In_851,In_2309);
nand U1586 (N_1586,N_38,In_1097);
nor U1587 (N_1587,In_2318,In_2412);
or U1588 (N_1588,In_667,In_239);
xnor U1589 (N_1589,In_2264,N_551);
or U1590 (N_1590,In_2325,N_221);
xnor U1591 (N_1591,In_2774,In_687);
nor U1592 (N_1592,N_776,N_768);
and U1593 (N_1593,In_2454,N_22);
nor U1594 (N_1594,N_1116,N_393);
nand U1595 (N_1595,In_577,In_1695);
nor U1596 (N_1596,N_184,N_847);
xnor U1597 (N_1597,N_397,In_2586);
nand U1598 (N_1598,N_626,In_635);
and U1599 (N_1599,N_749,N_1011);
xnor U1600 (N_1600,N_1139,N_667);
and U1601 (N_1601,In_1185,In_2086);
or U1602 (N_1602,N_35,N_48);
nand U1603 (N_1603,N_547,N_77);
and U1604 (N_1604,N_608,N_1160);
nand U1605 (N_1605,N_1031,N_1167);
nand U1606 (N_1606,N_1072,In_1389);
and U1607 (N_1607,N_645,N_44);
or U1608 (N_1608,In_150,In_2877);
and U1609 (N_1609,N_933,N_479);
or U1610 (N_1610,N_426,N_871);
nor U1611 (N_1611,N_264,In_1777);
nor U1612 (N_1612,In_167,N_770);
or U1613 (N_1613,In_998,N_220);
nand U1614 (N_1614,In_2492,N_544);
or U1615 (N_1615,N_78,In_50);
xor U1616 (N_1616,In_220,N_1109);
nor U1617 (N_1617,N_540,N_138);
nor U1618 (N_1618,N_1153,N_954);
or U1619 (N_1619,N_761,N_931);
nor U1620 (N_1620,N_657,N_496);
xnor U1621 (N_1621,In_2125,N_121);
xor U1622 (N_1622,N_832,N_867);
and U1623 (N_1623,N_837,N_1156);
or U1624 (N_1624,N_701,In_1951);
and U1625 (N_1625,In_1718,N_890);
nor U1626 (N_1626,In_1394,N_510);
or U1627 (N_1627,In_1734,N_134);
or U1628 (N_1628,N_678,N_193);
nand U1629 (N_1629,N_842,In_2306);
xnor U1630 (N_1630,In_408,N_125);
nor U1631 (N_1631,In_2705,N_875);
or U1632 (N_1632,In_997,In_2872);
nand U1633 (N_1633,In_792,N_240);
xnor U1634 (N_1634,N_115,N_639);
and U1635 (N_1635,In_1771,N_908);
nor U1636 (N_1636,N_505,In_2105);
and U1637 (N_1637,N_1198,N_783);
nor U1638 (N_1638,N_894,N_187);
nand U1639 (N_1639,N_75,In_1602);
and U1640 (N_1640,N_279,N_760);
or U1641 (N_1641,N_492,N_972);
and U1642 (N_1642,N_26,N_1084);
nand U1643 (N_1643,N_966,N_1015);
and U1644 (N_1644,In_1487,In_515);
xnor U1645 (N_1645,N_981,N_315);
nor U1646 (N_1646,N_600,In_884);
and U1647 (N_1647,In_1614,N_332);
nor U1648 (N_1648,In_1791,N_88);
or U1649 (N_1649,In_1000,In_1224);
nand U1650 (N_1650,N_777,N_218);
or U1651 (N_1651,In_2247,In_2114);
xnor U1652 (N_1652,In_767,In_1854);
nor U1653 (N_1653,In_1469,N_1146);
nand U1654 (N_1654,In_854,N_130);
nor U1655 (N_1655,N_703,N_529);
nor U1656 (N_1656,N_884,In_1656);
or U1657 (N_1657,N_725,N_1113);
nand U1658 (N_1658,N_446,N_70);
xor U1659 (N_1659,In_1574,N_443);
and U1660 (N_1660,N_336,N_372);
or U1661 (N_1661,N_582,In_189);
nand U1662 (N_1662,N_1184,N_347);
and U1663 (N_1663,N_1046,N_1159);
nand U1664 (N_1664,N_213,N_723);
xor U1665 (N_1665,N_898,In_1260);
and U1666 (N_1666,N_836,In_495);
or U1667 (N_1667,N_500,In_2425);
nor U1668 (N_1668,N_498,N_128);
or U1669 (N_1669,N_793,N_585);
and U1670 (N_1670,N_935,In_539);
xnor U1671 (N_1671,In_540,N_986);
or U1672 (N_1672,N_521,In_1396);
nor U1673 (N_1673,In_2497,N_1069);
xnor U1674 (N_1674,In_2842,N_72);
xnor U1675 (N_1675,N_512,N_284);
nand U1676 (N_1676,N_526,N_147);
and U1677 (N_1677,In_1585,In_1937);
nand U1678 (N_1678,In_2329,N_514);
or U1679 (N_1679,N_433,N_625);
nand U1680 (N_1680,N_872,N_503);
nand U1681 (N_1681,In_1902,N_99);
or U1682 (N_1682,N_1009,N_488);
and U1683 (N_1683,In_2358,N_1158);
nand U1684 (N_1684,N_775,In_1925);
and U1685 (N_1685,N_349,In_2641);
nand U1686 (N_1686,In_420,In_258);
or U1687 (N_1687,In_1432,N_1037);
and U1688 (N_1688,N_1150,N_697);
or U1689 (N_1689,In_1050,N_312);
xor U1690 (N_1690,N_227,N_322);
nor U1691 (N_1691,N_1172,N_671);
nand U1692 (N_1692,N_1120,N_442);
or U1693 (N_1693,N_889,N_1119);
and U1694 (N_1694,In_2908,In_1619);
and U1695 (N_1695,N_1193,In_2975);
nand U1696 (N_1696,N_928,N_567);
nor U1697 (N_1697,N_772,In_342);
and U1698 (N_1698,In_403,N_137);
nand U1699 (N_1699,In_2303,In_2963);
and U1700 (N_1700,N_618,N_533);
xor U1701 (N_1701,N_590,In_1378);
nand U1702 (N_1702,N_991,N_116);
xnor U1703 (N_1703,N_1051,In_763);
nor U1704 (N_1704,N_531,N_359);
or U1705 (N_1705,N_636,N_861);
or U1706 (N_1706,In_1145,N_458);
xor U1707 (N_1707,N_245,N_554);
nor U1708 (N_1708,In_130,N_888);
and U1709 (N_1709,N_810,N_460);
nand U1710 (N_1710,N_2,In_1434);
or U1711 (N_1711,In_1975,N_1052);
nor U1712 (N_1712,N_468,N_546);
nor U1713 (N_1713,In_1322,N_739);
or U1714 (N_1714,N_580,N_176);
and U1715 (N_1715,In_206,N_421);
nor U1716 (N_1716,N_353,In_1053);
and U1717 (N_1717,N_967,N_108);
nor U1718 (N_1718,N_68,N_1144);
nor U1719 (N_1719,N_571,In_954);
nor U1720 (N_1720,In_716,N_435);
nor U1721 (N_1721,N_1137,N_18);
and U1722 (N_1722,In_2331,N_217);
nor U1723 (N_1723,In_1834,N_81);
and U1724 (N_1724,N_1169,N_136);
and U1725 (N_1725,N_259,N_1033);
xnor U1726 (N_1726,N_249,N_664);
or U1727 (N_1727,N_295,In_620);
xnor U1728 (N_1728,In_56,In_745);
or U1729 (N_1729,In_2605,N_670);
nor U1730 (N_1730,In_60,In_75);
xnor U1731 (N_1731,N_617,N_67);
or U1732 (N_1732,N_690,N_457);
nand U1733 (N_1733,N_381,N_305);
and U1734 (N_1734,N_961,N_815);
and U1735 (N_1735,In_1891,N_1191);
nor U1736 (N_1736,N_827,N_919);
and U1737 (N_1737,In_2513,N_261);
nor U1738 (N_1738,N_437,N_630);
xor U1739 (N_1739,In_703,In_2208);
or U1740 (N_1740,In_1566,N_819);
xnor U1741 (N_1741,N_744,N_1133);
or U1742 (N_1742,In_2161,N_845);
xnor U1743 (N_1743,N_612,N_1163);
nand U1744 (N_1744,N_82,N_965);
nor U1745 (N_1745,In_2844,In_187);
xnor U1746 (N_1746,N_64,In_1031);
xnor U1747 (N_1747,N_159,N_394);
or U1748 (N_1748,In_886,N_161);
nor U1749 (N_1749,N_111,N_90);
or U1750 (N_1750,N_276,N_669);
xnor U1751 (N_1751,In_557,In_330);
xnor U1752 (N_1752,N_1188,In_1862);
nor U1753 (N_1753,N_1083,N_114);
and U1754 (N_1754,N_620,N_881);
nand U1755 (N_1755,In_1495,N_1179);
and U1756 (N_1756,N_509,In_1178);
nand U1757 (N_1757,N_155,N_28);
and U1758 (N_1758,In_1170,In_1883);
nor U1759 (N_1759,In_1426,N_953);
or U1760 (N_1760,N_915,N_392);
or U1761 (N_1761,In_20,N_272);
and U1762 (N_1762,N_916,In_1048);
nor U1763 (N_1763,N_886,N_1178);
or U1764 (N_1764,In_785,N_470);
nand U1765 (N_1765,In_2316,N_300);
xor U1766 (N_1766,In_1903,In_503);
or U1767 (N_1767,N_990,N_528);
nand U1768 (N_1768,N_791,In_2429);
or U1769 (N_1769,In_279,N_181);
and U1770 (N_1770,N_596,In_2199);
nand U1771 (N_1771,N_878,N_440);
nand U1772 (N_1772,N_1175,In_2749);
or U1773 (N_1773,In_1009,N_278);
and U1774 (N_1774,N_110,N_436);
and U1775 (N_1775,N_370,N_1118);
or U1776 (N_1776,N_676,In_100);
or U1777 (N_1777,N_1100,N_39);
and U1778 (N_1778,N_807,N_1173);
and U1779 (N_1779,In_2665,In_268);
xnor U1780 (N_1780,In_45,N_365);
nor U1781 (N_1781,In_1343,N_545);
and U1782 (N_1782,N_102,In_1100);
nand U1783 (N_1783,N_1103,N_732);
xor U1784 (N_1784,N_258,In_2290);
and U1785 (N_1785,N_139,N_522);
and U1786 (N_1786,N_686,N_508);
xor U1787 (N_1787,In_1504,N_294);
xor U1788 (N_1788,In_2134,N_817);
and U1789 (N_1789,N_711,In_405);
or U1790 (N_1790,In_1497,N_164);
xnor U1791 (N_1791,N_780,In_449);
nor U1792 (N_1792,In_1747,In_310);
nand U1793 (N_1793,In_1968,N_798);
xnor U1794 (N_1794,N_579,N_913);
nor U1795 (N_1795,N_462,In_820);
nor U1796 (N_1796,N_384,N_309);
or U1797 (N_1797,In_0,N_407);
nand U1798 (N_1798,N_491,In_1763);
nor U1799 (N_1799,N_400,N_1127);
nor U1800 (N_1800,N_700,In_1353);
and U1801 (N_1801,N_306,In_741);
and U1802 (N_1802,N_1078,N_311);
nand U1803 (N_1803,N_207,N_1036);
and U1804 (N_1804,N_906,In_2886);
nor U1805 (N_1805,N_552,N_350);
or U1806 (N_1806,In_1716,N_499);
or U1807 (N_1807,In_369,In_2766);
nor U1808 (N_1808,N_624,N_632);
nand U1809 (N_1809,N_688,N_504);
or U1810 (N_1810,N_1101,In_2991);
xor U1811 (N_1811,In_1494,In_2649);
nor U1812 (N_1812,N_719,In_1757);
and U1813 (N_1813,N_566,N_1017);
xor U1814 (N_1814,N_824,N_65);
and U1815 (N_1815,N_614,In_1926);
or U1816 (N_1816,N_391,In_1952);
and U1817 (N_1817,N_476,N_368);
xnor U1818 (N_1818,In_1440,N_478);
nor U1819 (N_1819,N_1043,N_828);
xor U1820 (N_1820,N_271,N_769);
nand U1821 (N_1821,In_242,In_2596);
or U1822 (N_1822,N_1001,In_2950);
nand U1823 (N_1823,N_535,N_157);
or U1824 (N_1824,N_42,N_781);
xor U1825 (N_1825,N_568,In_1517);
nand U1826 (N_1826,N_794,N_595);
xnor U1827 (N_1827,N_710,N_606);
nor U1828 (N_1828,N_448,In_2778);
nor U1829 (N_1829,In_324,N_907);
or U1830 (N_1830,In_662,In_523);
and U1831 (N_1831,N_880,N_578);
or U1832 (N_1832,In_296,N_1012);
xor U1833 (N_1833,N_127,In_6);
xor U1834 (N_1834,N_708,In_97);
and U1835 (N_1835,In_2970,N_4);
and U1836 (N_1836,N_642,N_605);
nand U1837 (N_1837,N_423,N_1128);
and U1838 (N_1838,N_1054,In_1293);
xor U1839 (N_1839,N_113,N_124);
nand U1840 (N_1840,N_627,N_109);
nand U1841 (N_1841,N_120,N_773);
nor U1842 (N_1842,N_281,N_728);
nor U1843 (N_1843,N_859,N_395);
nand U1844 (N_1844,N_1195,N_154);
xnor U1845 (N_1845,In_341,In_237);
nand U1846 (N_1846,N_317,In_2754);
xor U1847 (N_1847,N_277,N_839);
nor U1848 (N_1848,N_985,N_1049);
and U1849 (N_1849,N_782,In_1196);
and U1850 (N_1850,In_387,N_485);
or U1851 (N_1851,N_1143,N_1176);
xnor U1852 (N_1852,N_939,N_952);
nand U1853 (N_1853,N_640,N_170);
xor U1854 (N_1854,N_980,N_864);
nand U1855 (N_1855,In_720,N_320);
nor U1856 (N_1856,In_2905,N_292);
xor U1857 (N_1857,N_246,N_202);
and U1858 (N_1858,N_869,N_53);
nand U1859 (N_1859,N_304,N_748);
nor U1860 (N_1860,N_975,N_144);
nand U1861 (N_1861,N_1180,N_1080);
nor U1862 (N_1862,N_1077,N_682);
and U1863 (N_1863,N_644,In_2495);
nor U1864 (N_1864,In_1104,N_574);
and U1865 (N_1865,N_49,In_397);
or U1866 (N_1866,N_638,N_575);
and U1867 (N_1867,In_1916,N_344);
nand U1868 (N_1868,In_1536,In_1848);
xnor U1869 (N_1869,N_673,In_2174);
nand U1870 (N_1870,In_2244,N_1115);
and U1871 (N_1871,N_729,N_1138);
xor U1872 (N_1872,In_46,N_1197);
nand U1873 (N_1873,N_922,In_40);
and U1874 (N_1874,N_1182,N_194);
xor U1875 (N_1875,N_135,In_1415);
nand U1876 (N_1876,In_124,N_808);
nor U1877 (N_1877,N_1002,In_1931);
or U1878 (N_1878,In_1836,N_577);
and U1879 (N_1879,In_1914,In_2020);
and U1880 (N_1880,N_1130,N_222);
nor U1881 (N_1881,N_168,N_422);
nand U1882 (N_1882,N_166,N_745);
nor U1883 (N_1883,N_806,N_321);
and U1884 (N_1884,N_714,N_1005);
xor U1885 (N_1885,N_822,In_1466);
and U1886 (N_1886,In_68,In_549);
or U1887 (N_1887,N_1092,In_2912);
xor U1888 (N_1888,In_1939,N_55);
xnor U1889 (N_1889,In_1039,N_762);
and U1890 (N_1890,N_1040,N_750);
and U1891 (N_1891,In_2487,N_1050);
xor U1892 (N_1892,N_948,N_274);
xor U1893 (N_1893,N_549,N_914);
nand U1894 (N_1894,In_771,In_2837);
nor U1895 (N_1895,N_1059,N_949);
xnor U1896 (N_1896,N_661,N_957);
nand U1897 (N_1897,N_389,In_878);
nor U1898 (N_1898,In_2227,N_282);
nor U1899 (N_1899,N_160,In_2186);
or U1900 (N_1900,N_209,N_1174);
or U1901 (N_1901,N_877,In_571);
or U1902 (N_1902,N_789,N_666);
nor U1903 (N_1903,In_410,In_1082);
nor U1904 (N_1904,In_16,N_902);
nand U1905 (N_1905,In_149,In_2781);
xor U1906 (N_1906,In_1063,N_34);
or U1907 (N_1907,In_275,N_646);
xnor U1908 (N_1908,N_727,In_2516);
nor U1909 (N_1909,In_191,N_1019);
and U1910 (N_1910,In_1071,In_2639);
and U1911 (N_1911,N_30,N_58);
nand U1912 (N_1912,N_319,N_27);
and U1913 (N_1913,N_538,In_898);
or U1914 (N_1914,In_1730,N_652);
nand U1915 (N_1915,N_150,N_239);
nand U1916 (N_1916,N_1065,In_2466);
or U1917 (N_1917,N_1032,In_19);
nand U1918 (N_1918,In_1236,N_643);
xor U1919 (N_1919,N_795,N_367);
and U1920 (N_1920,N_377,In_285);
nand U1921 (N_1921,N_105,In_2092);
or U1922 (N_1922,In_2933,N_1194);
nor U1923 (N_1923,N_853,In_2116);
xor U1924 (N_1924,N_262,In_1413);
xnor U1925 (N_1925,In_1589,N_879);
nor U1926 (N_1926,N_586,N_731);
nor U1927 (N_1927,In_1028,N_52);
nand U1928 (N_1928,N_119,In_1443);
xnor U1929 (N_1929,In_2354,In_2000);
or U1930 (N_1930,N_148,N_816);
or U1931 (N_1931,N_969,N_482);
or U1932 (N_1932,N_741,N_863);
and U1933 (N_1933,In_1658,N_665);
or U1934 (N_1934,N_0,In_2469);
or U1935 (N_1935,In_2498,N_734);
or U1936 (N_1936,N_29,In_848);
nand U1937 (N_1937,N_425,N_404);
nand U1938 (N_1938,In_977,N_223);
nor U1939 (N_1939,N_938,N_228);
nand U1940 (N_1940,In_1162,N_420);
or U1941 (N_1941,N_97,N_996);
or U1942 (N_1942,N_286,N_192);
or U1943 (N_1943,N_588,N_256);
or U1944 (N_1944,N_993,N_751);
or U1945 (N_1945,N_1016,N_763);
and U1946 (N_1946,N_974,N_371);
xnor U1947 (N_1947,N_662,N_823);
or U1948 (N_1948,In_1520,N_172);
nor U1949 (N_1949,In_1246,N_757);
or U1950 (N_1950,N_208,In_1919);
and U1951 (N_1951,In_2926,N_733);
and U1952 (N_1952,In_2585,N_515);
nor U1953 (N_1953,In_822,In_2960);
and U1954 (N_1954,N_175,In_901);
and U1955 (N_1955,N_248,N_1148);
nand U1956 (N_1956,In_2816,N_118);
xor U1957 (N_1957,N_412,N_835);
xor U1958 (N_1958,N_559,In_2818);
nand U1959 (N_1959,In_1338,In_1929);
or U1960 (N_1960,In_2133,N_107);
and U1961 (N_1961,N_694,N_801);
nor U1962 (N_1962,N_7,In_2919);
xnor U1963 (N_1963,In_2557,N_743);
nor U1964 (N_1964,In_2611,In_2951);
xnor U1965 (N_1965,N_480,In_742);
and U1966 (N_1966,In_1833,In_831);
or U1967 (N_1967,N_333,N_1004);
xor U1968 (N_1968,N_243,In_209);
nand U1969 (N_1969,In_558,N_494);
or U1970 (N_1970,In_172,N_1099);
xnor U1971 (N_1971,N_520,N_1060);
xor U1972 (N_1972,N_702,N_598);
nand U1973 (N_1973,In_372,N_493);
and U1974 (N_1974,In_1056,N_909);
nor U1975 (N_1975,N_334,N_37);
nand U1976 (N_1976,N_1075,In_2180);
and U1977 (N_1977,In_2302,In_2391);
and U1978 (N_1978,In_2972,N_481);
xnor U1979 (N_1979,In_2986,N_244);
nand U1980 (N_1980,N_753,N_720);
nand U1981 (N_1981,In_270,N_156);
xor U1982 (N_1982,In_2117,N_376);
or U1983 (N_1983,In_2584,N_695);
nand U1984 (N_1984,In_2184,N_287);
and U1985 (N_1985,N_1168,N_742);
nor U1986 (N_1986,N_755,N_583);
and U1987 (N_1987,N_602,N_998);
nor U1988 (N_1988,N_363,In_1813);
nor U1989 (N_1989,N_658,N_225);
nand U1990 (N_1990,N_409,In_2901);
and U1991 (N_1991,N_293,In_1438);
nand U1992 (N_1992,N_655,N_1112);
and U1993 (N_1993,N_471,N_1013);
xor U1994 (N_1994,N_1091,N_641);
xor U1995 (N_1995,N_848,N_513);
nor U1996 (N_1996,In_587,N_51);
nand U1997 (N_1997,N_680,In_2523);
nand U1998 (N_1998,N_622,N_1125);
nor U1999 (N_1999,N_439,N_873);
nor U2000 (N_2000,N_206,N_621);
xnor U2001 (N_2001,N_1074,N_390);
or U2002 (N_2002,N_539,N_123);
xor U2003 (N_2003,In_628,N_558);
nand U2004 (N_2004,In_380,N_182);
nor U2005 (N_2005,N_787,In_1400);
xnor U2006 (N_2006,In_598,N_1086);
or U2007 (N_2007,In_2524,N_486);
xor U2008 (N_2008,In_1637,N_415);
xnor U2009 (N_2009,N_663,In_2852);
nor U2010 (N_2010,N_453,N_310);
nor U2011 (N_2011,N_994,N_1062);
xor U2012 (N_2012,N_653,N_599);
nor U2013 (N_2013,N_386,In_917);
nand U2014 (N_2014,N_451,N_681);
nand U2015 (N_2015,N_812,N_628);
nor U2016 (N_2016,N_988,N_431);
nor U2017 (N_2017,In_385,N_232);
and U2018 (N_2018,N_1157,N_456);
nand U2019 (N_2019,In_2998,N_825);
nor U2020 (N_2020,N_444,N_804);
nor U2021 (N_2021,N_233,N_698);
nand U2022 (N_2022,N_1029,In_2460);
nor U2023 (N_2023,N_1095,N_651);
xnor U2024 (N_2024,In_91,N_417);
xnor U2025 (N_2025,N_497,N_40);
or U2026 (N_2026,In_2475,N_870);
nand U2027 (N_2027,N_995,In_437);
nand U2028 (N_2028,In_1011,In_1194);
or U2029 (N_2029,N_934,N_736);
nand U2030 (N_2030,N_411,N_893);
and U2031 (N_2031,In_1458,In_2657);
or U2032 (N_2032,N_188,N_887);
and U2033 (N_2033,N_587,N_45);
and U2034 (N_2034,N_430,N_947);
xnor U2035 (N_2035,N_379,N_133);
or U2036 (N_2036,In_1664,In_496);
and U2037 (N_2037,In_2728,N_619);
nand U2038 (N_2038,N_660,N_59);
and U2039 (N_2039,N_527,N_840);
nand U2040 (N_2040,N_917,N_428);
nand U2041 (N_2041,N_445,N_483);
xor U2042 (N_2042,In_1921,N_1071);
xnor U2043 (N_2043,N_143,N_327);
xnor U2044 (N_2044,N_1024,In_944);
nor U2045 (N_2045,N_1164,In_389);
nor U2046 (N_2046,In_353,N_885);
nor U2047 (N_2047,In_482,In_960);
and U2048 (N_2048,In_1814,N_414);
xor U2049 (N_2049,In_655,In_1456);
or U2050 (N_2050,In_2084,N_1107);
nand U2051 (N_2051,In_1844,N_87);
xnor U2052 (N_2052,N_358,N_633);
or U2053 (N_2053,In_2211,N_1136);
nor U2054 (N_2054,In_2450,N_1026);
nand U2055 (N_2055,N_69,N_316);
nand U2056 (N_2056,In_2162,N_329);
xnor U2057 (N_2057,N_179,In_1270);
and U2058 (N_2058,N_91,N_338);
nand U2059 (N_2059,In_2094,N_158);
nand U2060 (N_2060,In_728,N_911);
xor U2061 (N_2061,N_930,N_637);
and U2062 (N_2062,N_15,N_242);
or U2063 (N_2063,N_555,N_129);
xor U2064 (N_2064,N_1123,In_361);
nor U2065 (N_2065,N_1067,N_416);
or U2066 (N_2066,In_127,In_775);
nor U2067 (N_2067,N_1190,N_270);
xnor U2068 (N_2068,In_22,N_355);
and U2069 (N_2069,In_2432,In_392);
or U2070 (N_2070,In_2175,In_548);
and U2071 (N_2071,N_1132,N_648);
nand U2072 (N_2072,N_89,N_432);
nand U2073 (N_2073,N_303,N_765);
and U2074 (N_2074,N_183,N_141);
or U2075 (N_2075,N_1039,N_553);
nor U2076 (N_2076,In_1281,N_629);
xnor U2077 (N_2077,N_362,In_1651);
nand U2078 (N_2078,In_2607,N_704);
nand U2079 (N_2079,In_2653,N_211);
and U2080 (N_2080,N_203,N_1151);
nor U2081 (N_2081,N_1134,N_992);
or U2082 (N_2082,In_933,N_982);
and U2083 (N_2083,N_592,N_891);
nor U2084 (N_2084,N_997,N_846);
nor U2085 (N_2085,In_899,N_71);
nor U2086 (N_2086,N_874,In_2989);
or U2087 (N_2087,In_1526,In_2955);
nand U2088 (N_2088,In_2164,N_238);
nand U2089 (N_2089,N_865,In_2452);
nor U2090 (N_2090,N_375,In_386);
xor U2091 (N_2091,N_936,N_722);
and U2092 (N_2092,In_882,N_1057);
nand U2093 (N_2093,In_87,In_1233);
nor U2094 (N_2094,N_654,In_2573);
and U2095 (N_2095,N_323,N_1044);
xnor U2096 (N_2096,N_833,N_778);
and U2097 (N_2097,N_971,N_1111);
nand U2098 (N_2098,In_2218,N_413);
and U2099 (N_2099,In_1812,N_265);
nor U2100 (N_2100,N_60,In_1199);
and U2101 (N_2101,N_263,N_250);
or U2102 (N_2102,N_48,In_2358);
nor U2103 (N_2103,N_61,In_2576);
nand U2104 (N_2104,In_2608,N_895);
nand U2105 (N_2105,N_350,N_1145);
xnor U2106 (N_2106,In_2391,In_482);
and U2107 (N_2107,N_1175,N_973);
and U2108 (N_2108,N_58,In_2886);
nor U2109 (N_2109,N_88,In_1325);
nand U2110 (N_2110,N_512,In_1431);
xnor U2111 (N_2111,N_1112,N_1041);
nor U2112 (N_2112,In_372,In_1658);
xnor U2113 (N_2113,N_1091,N_474);
nand U2114 (N_2114,N_521,N_946);
or U2115 (N_2115,In_2108,N_516);
nor U2116 (N_2116,N_294,In_2524);
nor U2117 (N_2117,N_368,N_505);
and U2118 (N_2118,In_1798,N_104);
and U2119 (N_2119,N_139,N_751);
nand U2120 (N_2120,In_2774,N_167);
and U2121 (N_2121,N_496,N_313);
nand U2122 (N_2122,N_929,N_369);
and U2123 (N_2123,N_663,In_655);
nor U2124 (N_2124,N_664,N_423);
xnor U2125 (N_2125,N_955,N_163);
or U2126 (N_2126,In_2339,N_863);
nor U2127 (N_2127,N_262,In_616);
nor U2128 (N_2128,N_659,In_540);
xnor U2129 (N_2129,N_672,N_22);
nand U2130 (N_2130,In_1650,In_502);
nor U2131 (N_2131,In_185,In_1442);
nor U2132 (N_2132,N_225,N_1040);
nor U2133 (N_2133,N_1117,N_907);
and U2134 (N_2134,In_1874,N_1156);
nor U2135 (N_2135,N_284,N_428);
nand U2136 (N_2136,N_841,N_802);
xnor U2137 (N_2137,In_2611,In_632);
xnor U2138 (N_2138,In_239,In_2549);
nor U2139 (N_2139,N_810,N_634);
nor U2140 (N_2140,N_778,In_2762);
and U2141 (N_2141,In_1193,N_372);
or U2142 (N_2142,N_655,N_518);
nor U2143 (N_2143,N_797,N_1021);
nand U2144 (N_2144,N_1002,N_738);
and U2145 (N_2145,N_588,N_563);
or U2146 (N_2146,N_544,N_609);
or U2147 (N_2147,N_978,In_1246);
nor U2148 (N_2148,N_1118,In_2611);
xnor U2149 (N_2149,N_180,N_328);
nand U2150 (N_2150,N_248,N_553);
and U2151 (N_2151,In_2551,In_886);
and U2152 (N_2152,N_1062,In_2593);
or U2153 (N_2153,N_412,In_2926);
and U2154 (N_2154,In_100,In_1931);
nor U2155 (N_2155,N_39,In_1166);
xor U2156 (N_2156,N_51,N_45);
nand U2157 (N_2157,N_165,N_986);
nor U2158 (N_2158,In_2498,In_539);
and U2159 (N_2159,N_143,N_675);
nand U2160 (N_2160,N_1154,N_936);
and U2161 (N_2161,N_468,N_827);
nor U2162 (N_2162,In_2000,N_791);
xor U2163 (N_2163,N_680,In_1763);
or U2164 (N_2164,N_3,N_1109);
and U2165 (N_2165,N_702,In_172);
and U2166 (N_2166,N_131,N_723);
xnor U2167 (N_2167,In_1749,N_101);
xnor U2168 (N_2168,N_870,N_86);
nor U2169 (N_2169,N_501,In_1252);
nand U2170 (N_2170,N_644,N_1021);
and U2171 (N_2171,N_968,N_331);
or U2172 (N_2172,N_55,In_899);
nor U2173 (N_2173,In_333,N_429);
and U2174 (N_2174,N_115,In_2450);
or U2175 (N_2175,In_73,In_1347);
nand U2176 (N_2176,In_2530,N_735);
xor U2177 (N_2177,N_248,N_1117);
or U2178 (N_2178,N_1183,N_683);
and U2179 (N_2179,In_2959,N_214);
xnor U2180 (N_2180,N_660,N_560);
or U2181 (N_2181,N_327,N_916);
nor U2182 (N_2182,In_2475,N_427);
nand U2183 (N_2183,In_179,N_904);
nor U2184 (N_2184,N_304,N_815);
or U2185 (N_2185,N_246,N_902);
or U2186 (N_2186,N_910,N_345);
xnor U2187 (N_2187,In_2581,N_683);
or U2188 (N_2188,In_179,N_615);
and U2189 (N_2189,N_116,N_364);
xor U2190 (N_2190,N_928,N_100);
and U2191 (N_2191,N_640,N_886);
nor U2192 (N_2192,In_557,N_510);
nand U2193 (N_2193,N_1126,N_201);
nor U2194 (N_2194,In_0,In_1734);
nor U2195 (N_2195,In_1145,N_451);
nor U2196 (N_2196,N_889,N_408);
and U2197 (N_2197,N_434,N_472);
nand U2198 (N_2198,N_788,N_387);
or U2199 (N_2199,N_891,In_333);
nand U2200 (N_2200,In_496,In_2450);
or U2201 (N_2201,In_1158,In_1614);
or U2202 (N_2202,In_175,In_2593);
xnor U2203 (N_2203,In_1540,N_36);
nor U2204 (N_2204,In_1097,In_2363);
xor U2205 (N_2205,In_1443,N_946);
xor U2206 (N_2206,N_910,N_484);
xor U2207 (N_2207,N_656,In_687);
and U2208 (N_2208,N_912,In_196);
xor U2209 (N_2209,In_2458,In_540);
nor U2210 (N_2210,N_344,In_169);
and U2211 (N_2211,N_115,N_933);
xor U2212 (N_2212,N_548,N_320);
nand U2213 (N_2213,N_88,In_1688);
nand U2214 (N_2214,In_2621,N_199);
and U2215 (N_2215,N_560,In_364);
nor U2216 (N_2216,N_829,N_272);
xnor U2217 (N_2217,N_756,In_2766);
and U2218 (N_2218,N_1120,N_294);
or U2219 (N_2219,N_1069,N_668);
nor U2220 (N_2220,N_719,N_499);
and U2221 (N_2221,In_45,N_519);
xor U2222 (N_2222,N_563,N_367);
and U2223 (N_2223,N_1073,N_499);
nand U2224 (N_2224,N_651,N_865);
nand U2225 (N_2225,In_1353,N_458);
nand U2226 (N_2226,In_1178,N_484);
nand U2227 (N_2227,In_1883,N_332);
or U2228 (N_2228,N_148,N_939);
nand U2229 (N_2229,N_486,In_106);
and U2230 (N_2230,In_1813,N_882);
xor U2231 (N_2231,N_174,N_365);
xor U2232 (N_2232,N_990,N_996);
and U2233 (N_2233,N_473,N_1039);
xor U2234 (N_2234,N_443,N_298);
or U2235 (N_2235,N_404,In_1937);
nand U2236 (N_2236,N_138,N_1118);
xnor U2237 (N_2237,N_193,N_554);
xor U2238 (N_2238,In_2495,In_2891);
and U2239 (N_2239,N_54,In_554);
or U2240 (N_2240,N_47,N_1154);
nor U2241 (N_2241,N_87,N_302);
nand U2242 (N_2242,N_186,N_45);
nand U2243 (N_2243,In_1763,N_447);
or U2244 (N_2244,In_2905,In_600);
and U2245 (N_2245,N_1124,N_873);
nand U2246 (N_2246,In_1566,In_162);
nor U2247 (N_2247,In_1003,N_480);
xnor U2248 (N_2248,In_2092,N_13);
nor U2249 (N_2249,In_2856,N_445);
or U2250 (N_2250,N_1126,N_256);
or U2251 (N_2251,N_420,N_909);
and U2252 (N_2252,N_1115,N_374);
xor U2253 (N_2253,N_1148,In_2852);
and U2254 (N_2254,N_40,N_231);
xor U2255 (N_2255,N_1069,N_468);
and U2256 (N_2256,N_267,N_1116);
or U2257 (N_2257,N_90,N_108);
xnor U2258 (N_2258,In_820,N_426);
xor U2259 (N_2259,In_716,In_2038);
nand U2260 (N_2260,N_679,N_73);
xor U2261 (N_2261,In_1295,N_879);
xnor U2262 (N_2262,N_1073,N_876);
or U2263 (N_2263,N_422,N_373);
and U2264 (N_2264,In_1504,N_1022);
nand U2265 (N_2265,N_194,N_749);
nand U2266 (N_2266,In_2331,N_1111);
or U2267 (N_2267,In_814,In_2649);
xor U2268 (N_2268,N_939,In_75);
nor U2269 (N_2269,In_2038,In_1923);
or U2270 (N_2270,In_1833,N_454);
xor U2271 (N_2271,In_2442,N_492);
nand U2272 (N_2272,N_806,N_660);
or U2273 (N_2273,N_1145,N_23);
nor U2274 (N_2274,N_109,N_626);
xor U2275 (N_2275,N_914,N_323);
nand U2276 (N_2276,N_279,N_422);
xor U2277 (N_2277,In_1931,N_941);
or U2278 (N_2278,N_808,N_1158);
nand U2279 (N_2279,N_638,In_2584);
nand U2280 (N_2280,In_2403,In_712);
nand U2281 (N_2281,N_523,N_925);
and U2282 (N_2282,In_848,In_29);
xnor U2283 (N_2283,N_317,In_2905);
nand U2284 (N_2284,N_673,N_1177);
or U2285 (N_2285,In_1566,N_242);
or U2286 (N_2286,N_117,N_1139);
nor U2287 (N_2287,In_169,In_771);
and U2288 (N_2288,N_862,N_257);
xor U2289 (N_2289,In_1914,N_783);
xor U2290 (N_2290,N_369,N_516);
nand U2291 (N_2291,N_312,In_179);
and U2292 (N_2292,N_676,N_574);
nor U2293 (N_2293,N_276,In_2111);
and U2294 (N_2294,N_895,N_272);
nor U2295 (N_2295,N_1001,N_1095);
or U2296 (N_2296,N_911,In_2908);
or U2297 (N_2297,N_1053,N_738);
nand U2298 (N_2298,N_164,In_2586);
or U2299 (N_2299,N_1177,In_193);
or U2300 (N_2300,N_385,In_73);
nand U2301 (N_2301,N_663,N_783);
nand U2302 (N_2302,In_2549,In_1343);
or U2303 (N_2303,In_2326,N_434);
nand U2304 (N_2304,N_216,In_2819);
or U2305 (N_2305,In_792,N_1041);
nand U2306 (N_2306,In_1254,N_1046);
nand U2307 (N_2307,N_542,N_987);
nor U2308 (N_2308,N_529,N_66);
nand U2309 (N_2309,N_76,In_506);
xnor U2310 (N_2310,N_882,N_1051);
or U2311 (N_2311,In_2516,In_2513);
xnor U2312 (N_2312,In_2586,N_825);
nor U2313 (N_2313,N_11,N_4);
or U2314 (N_2314,N_206,N_951);
or U2315 (N_2315,N_658,In_2499);
xor U2316 (N_2316,N_314,N_456);
or U2317 (N_2317,In_2249,N_224);
xor U2318 (N_2318,In_1497,N_1096);
and U2319 (N_2319,N_1178,N_477);
or U2320 (N_2320,In_1340,N_828);
xor U2321 (N_2321,N_829,In_724);
nor U2322 (N_2322,In_2844,N_442);
nor U2323 (N_2323,In_820,In_408);
xor U2324 (N_2324,N_1199,N_103);
nand U2325 (N_2325,N_412,In_270);
nand U2326 (N_2326,In_1757,In_438);
nor U2327 (N_2327,In_1759,N_446);
xnor U2328 (N_2328,N_372,N_1154);
or U2329 (N_2329,N_250,In_178);
xnor U2330 (N_2330,In_2326,N_1044);
and U2331 (N_2331,N_398,In_1353);
xnor U2332 (N_2332,In_283,N_786);
nor U2333 (N_2333,N_906,N_998);
nand U2334 (N_2334,In_1540,N_745);
xor U2335 (N_2335,N_108,In_2516);
xor U2336 (N_2336,N_716,N_943);
nand U2337 (N_2337,N_912,In_342);
xor U2338 (N_2338,N_1163,N_82);
nand U2339 (N_2339,N_58,N_879);
nand U2340 (N_2340,In_2000,N_487);
and U2341 (N_2341,N_45,In_2639);
xor U2342 (N_2342,N_764,N_794);
and U2343 (N_2343,N_499,In_1281);
nand U2344 (N_2344,In_2038,N_556);
or U2345 (N_2345,N_346,N_382);
nor U2346 (N_2346,N_1075,N_336);
xor U2347 (N_2347,N_359,In_1249);
xor U2348 (N_2348,In_2611,N_657);
and U2349 (N_2349,In_2000,N_562);
nor U2350 (N_2350,N_119,N_681);
and U2351 (N_2351,N_863,In_2778);
xor U2352 (N_2352,N_591,N_941);
xor U2353 (N_2353,N_620,In_1520);
xor U2354 (N_2354,N_13,N_689);
nor U2355 (N_2355,N_75,In_1485);
xnor U2356 (N_2356,N_463,In_1585);
nor U2357 (N_2357,In_1378,In_2513);
xnor U2358 (N_2358,N_687,N_967);
or U2359 (N_2359,In_1914,N_95);
and U2360 (N_2360,N_88,N_498);
nor U2361 (N_2361,N_539,N_324);
nor U2362 (N_2362,In_1812,N_234);
or U2363 (N_2363,In_2068,N_738);
or U2364 (N_2364,In_731,N_1105);
nor U2365 (N_2365,N_789,In_2886);
xnor U2366 (N_2366,In_2608,N_852);
nor U2367 (N_2367,N_336,In_936);
or U2368 (N_2368,N_838,N_673);
xnor U2369 (N_2369,In_2108,N_347);
nand U2370 (N_2370,N_692,N_68);
or U2371 (N_2371,N_1081,In_2117);
and U2372 (N_2372,In_936,N_874);
or U2373 (N_2373,N_525,N_98);
nand U2374 (N_2374,In_1504,N_112);
or U2375 (N_2375,N_600,N_998);
and U2376 (N_2376,In_940,N_98);
and U2377 (N_2377,N_924,In_1034);
and U2378 (N_2378,N_396,N_786);
nand U2379 (N_2379,In_372,N_552);
and U2380 (N_2380,N_250,N_143);
nand U2381 (N_2381,In_149,In_2358);
and U2382 (N_2382,N_525,N_247);
nor U2383 (N_2383,N_1136,In_620);
and U2384 (N_2384,In_1322,N_1070);
and U2385 (N_2385,N_619,N_1052);
nand U2386 (N_2386,N_938,N_381);
and U2387 (N_2387,In_872,N_326);
and U2388 (N_2388,N_969,N_1199);
xor U2389 (N_2389,In_172,In_1194);
nor U2390 (N_2390,N_240,N_62);
xnor U2391 (N_2391,N_1039,N_1132);
nand U2392 (N_2392,N_534,In_2852);
xor U2393 (N_2393,N_732,In_367);
xor U2394 (N_2394,In_1000,In_2607);
nor U2395 (N_2395,In_1236,N_678);
nor U2396 (N_2396,In_2498,N_874);
nand U2397 (N_2397,N_400,N_1078);
nor U2398 (N_2398,N_496,N_564);
nor U2399 (N_2399,N_898,N_22);
nor U2400 (N_2400,N_1617,N_1382);
or U2401 (N_2401,N_1760,N_1290);
nor U2402 (N_2402,N_1842,N_2077);
nor U2403 (N_2403,N_2152,N_1609);
or U2404 (N_2404,N_1692,N_2323);
nor U2405 (N_2405,N_1424,N_1643);
xnor U2406 (N_2406,N_1254,N_1326);
and U2407 (N_2407,N_2266,N_1548);
nand U2408 (N_2408,N_2210,N_2366);
nor U2409 (N_2409,N_2288,N_1366);
and U2410 (N_2410,N_1377,N_1249);
and U2411 (N_2411,N_1257,N_1245);
nor U2412 (N_2412,N_1357,N_2377);
and U2413 (N_2413,N_1573,N_2016);
nand U2414 (N_2414,N_1576,N_1260);
nand U2415 (N_2415,N_1409,N_1822);
or U2416 (N_2416,N_1704,N_1740);
nor U2417 (N_2417,N_1426,N_1989);
nor U2418 (N_2418,N_1845,N_2125);
nand U2419 (N_2419,N_1949,N_1721);
and U2420 (N_2420,N_1264,N_1475);
xor U2421 (N_2421,N_1946,N_2304);
or U2422 (N_2422,N_1579,N_2151);
xnor U2423 (N_2423,N_2342,N_1966);
xnor U2424 (N_2424,N_1283,N_1227);
or U2425 (N_2425,N_1272,N_1574);
and U2426 (N_2426,N_1994,N_1469);
xnor U2427 (N_2427,N_2061,N_1807);
xnor U2428 (N_2428,N_2078,N_2254);
nor U2429 (N_2429,N_1504,N_1559);
nor U2430 (N_2430,N_1282,N_2352);
nor U2431 (N_2431,N_1291,N_1995);
xor U2432 (N_2432,N_1316,N_1820);
nor U2433 (N_2433,N_2319,N_1857);
and U2434 (N_2434,N_1432,N_2073);
xor U2435 (N_2435,N_1870,N_2388);
and U2436 (N_2436,N_1892,N_1325);
nor U2437 (N_2437,N_2126,N_2317);
nand U2438 (N_2438,N_1418,N_1869);
nand U2439 (N_2439,N_1557,N_1205);
and U2440 (N_2440,N_1905,N_2264);
xor U2441 (N_2441,N_2386,N_2167);
xnor U2442 (N_2442,N_1259,N_1278);
nand U2443 (N_2443,N_1729,N_2337);
nand U2444 (N_2444,N_1275,N_1390);
xor U2445 (N_2445,N_2108,N_1303);
or U2446 (N_2446,N_2112,N_1737);
nand U2447 (N_2447,N_2148,N_1751);
and U2448 (N_2448,N_1431,N_1441);
nand U2449 (N_2449,N_2267,N_2208);
and U2450 (N_2450,N_2199,N_2391);
or U2451 (N_2451,N_1517,N_1956);
and U2452 (N_2452,N_2168,N_2291);
or U2453 (N_2453,N_2284,N_2081);
xnor U2454 (N_2454,N_1376,N_1626);
and U2455 (N_2455,N_1543,N_2235);
or U2456 (N_2456,N_2049,N_1637);
and U2457 (N_2457,N_2072,N_2348);
xnor U2458 (N_2458,N_1450,N_2233);
nor U2459 (N_2459,N_1670,N_1440);
nand U2460 (N_2460,N_2101,N_2054);
nand U2461 (N_2461,N_1246,N_1705);
and U2462 (N_2462,N_1638,N_2369);
xnor U2463 (N_2463,N_2368,N_1403);
xor U2464 (N_2464,N_1556,N_1420);
and U2465 (N_2465,N_2378,N_2028);
and U2466 (N_2466,N_1320,N_2023);
or U2467 (N_2467,N_1887,N_2040);
nor U2468 (N_2468,N_1301,N_1314);
nand U2469 (N_2469,N_1250,N_1329);
or U2470 (N_2470,N_2055,N_1564);
xnor U2471 (N_2471,N_1738,N_1458);
xor U2472 (N_2472,N_1970,N_1470);
nand U2473 (N_2473,N_2156,N_2035);
nand U2474 (N_2474,N_1448,N_1660);
nand U2475 (N_2475,N_2362,N_1319);
nand U2476 (N_2476,N_1306,N_1658);
and U2477 (N_2477,N_1761,N_2026);
nand U2478 (N_2478,N_1287,N_1715);
or U2479 (N_2479,N_2292,N_1951);
xor U2480 (N_2480,N_1948,N_1790);
xor U2481 (N_2481,N_1647,N_2012);
nand U2482 (N_2482,N_1388,N_1953);
xnor U2483 (N_2483,N_2294,N_2225);
nor U2484 (N_2484,N_1210,N_1687);
or U2485 (N_2485,N_1594,N_1498);
xnor U2486 (N_2486,N_2153,N_1874);
nand U2487 (N_2487,N_2336,N_1219);
xnor U2488 (N_2488,N_1554,N_1566);
nor U2489 (N_2489,N_2129,N_1629);
or U2490 (N_2490,N_1520,N_2221);
nor U2491 (N_2491,N_1233,N_2331);
nor U2492 (N_2492,N_1456,N_2371);
nor U2493 (N_2493,N_1493,N_2066);
and U2494 (N_2494,N_2296,N_1367);
nand U2495 (N_2495,N_1302,N_1960);
and U2496 (N_2496,N_1497,N_2370);
nand U2497 (N_2497,N_2176,N_2321);
and U2498 (N_2498,N_2015,N_2350);
nor U2499 (N_2499,N_1269,N_1865);
and U2500 (N_2500,N_2003,N_1500);
and U2501 (N_2501,N_1894,N_1622);
and U2502 (N_2502,N_1932,N_2027);
or U2503 (N_2503,N_2107,N_1963);
or U2504 (N_2504,N_1603,N_2216);
nor U2505 (N_2505,N_1982,N_1919);
nor U2506 (N_2506,N_1238,N_2299);
or U2507 (N_2507,N_2102,N_1755);
or U2508 (N_2508,N_2230,N_1639);
or U2509 (N_2509,N_2359,N_1881);
or U2510 (N_2510,N_1453,N_1502);
and U2511 (N_2511,N_1425,N_1665);
or U2512 (N_2512,N_2259,N_1797);
nand U2513 (N_2513,N_1336,N_1397);
nor U2514 (N_2514,N_2140,N_1833);
and U2515 (N_2515,N_1363,N_1296);
and U2516 (N_2516,N_2393,N_1856);
and U2517 (N_2517,N_2154,N_2051);
xor U2518 (N_2518,N_1411,N_2241);
xnor U2519 (N_2519,N_1372,N_2121);
and U2520 (N_2520,N_1795,N_1774);
nand U2521 (N_2521,N_1351,N_2089);
and U2522 (N_2522,N_1890,N_2227);
nand U2523 (N_2523,N_1612,N_2379);
or U2524 (N_2524,N_2374,N_1754);
nand U2525 (N_2525,N_1310,N_2137);
nor U2526 (N_2526,N_1240,N_1234);
xnor U2527 (N_2527,N_2250,N_1602);
and U2528 (N_2528,N_1863,N_1699);
and U2529 (N_2529,N_1414,N_1800);
or U2530 (N_2530,N_1746,N_2287);
xnor U2531 (N_2531,N_1987,N_2269);
nand U2532 (N_2532,N_1364,N_1619);
nor U2533 (N_2533,N_1630,N_1584);
or U2534 (N_2534,N_2302,N_1752);
xnor U2535 (N_2535,N_2138,N_2247);
or U2536 (N_2536,N_1975,N_1567);
nand U2537 (N_2537,N_2273,N_1945);
nor U2538 (N_2538,N_1930,N_2279);
nor U2539 (N_2539,N_2004,N_1582);
and U2540 (N_2540,N_1389,N_1950);
nor U2541 (N_2541,N_2071,N_2117);
xor U2542 (N_2542,N_1861,N_1385);
xnor U2543 (N_2543,N_2160,N_1811);
nor U2544 (N_2544,N_1258,N_1914);
xor U2545 (N_2545,N_1312,N_1819);
nand U2546 (N_2546,N_1702,N_1806);
nand U2547 (N_2547,N_1479,N_2118);
nand U2548 (N_2548,N_2310,N_2064);
and U2549 (N_2549,N_1247,N_2324);
nand U2550 (N_2550,N_1777,N_1483);
or U2551 (N_2551,N_2180,N_1361);
and U2552 (N_2552,N_1736,N_1540);
xor U2553 (N_2553,N_1748,N_1600);
xor U2554 (N_2554,N_1972,N_2084);
or U2555 (N_2555,N_1443,N_2022);
xor U2556 (N_2556,N_2276,N_1663);
or U2557 (N_2557,N_1749,N_1328);
and U2558 (N_2558,N_1262,N_1346);
or U2559 (N_2559,N_1625,N_1508);
and U2560 (N_2560,N_2146,N_2209);
xnor U2561 (N_2561,N_2007,N_1697);
and U2562 (N_2562,N_1590,N_1506);
nand U2563 (N_2563,N_1877,N_1267);
or U2564 (N_2564,N_1532,N_1848);
or U2565 (N_2565,N_1786,N_1775);
nor U2566 (N_2566,N_1354,N_1536);
or U2567 (N_2567,N_2345,N_1709);
nor U2568 (N_2568,N_2372,N_1779);
nor U2569 (N_2569,N_2075,N_1534);
nand U2570 (N_2570,N_1862,N_2270);
or U2571 (N_2571,N_1356,N_1438);
nor U2572 (N_2572,N_1313,N_2177);
or U2573 (N_2573,N_1488,N_2063);
xnor U2574 (N_2574,N_1350,N_2231);
and U2575 (N_2575,N_1521,N_1668);
nor U2576 (N_2576,N_1967,N_2364);
nand U2577 (N_2577,N_2019,N_1788);
and U2578 (N_2578,N_1391,N_1591);
and U2579 (N_2579,N_1792,N_2303);
nor U2580 (N_2580,N_2262,N_1642);
xor U2581 (N_2581,N_1941,N_2173);
nor U2582 (N_2582,N_1286,N_1631);
nor U2583 (N_2583,N_1201,N_1791);
and U2584 (N_2584,N_1375,N_1846);
xor U2585 (N_2585,N_1449,N_1731);
xor U2586 (N_2586,N_2339,N_2002);
nor U2587 (N_2587,N_1365,N_2358);
nor U2588 (N_2588,N_2001,N_1598);
xor U2589 (N_2589,N_1990,N_1206);
nor U2590 (N_2590,N_1942,N_2340);
nor U2591 (N_2591,N_2045,N_1937);
nand U2592 (N_2592,N_1596,N_2005);
xnor U2593 (N_2593,N_1527,N_1929);
nor U2594 (N_2594,N_1383,N_2316);
or U2595 (N_2595,N_1974,N_1789);
xnor U2596 (N_2596,N_1802,N_1537);
xnor U2597 (N_2597,N_2215,N_1624);
nand U2598 (N_2598,N_1778,N_1655);
xnor U2599 (N_2599,N_1879,N_1433);
and U2600 (N_2600,N_1243,N_1682);
nand U2601 (N_2601,N_1969,N_2275);
nand U2602 (N_2602,N_1374,N_1916);
nand U2603 (N_2603,N_1962,N_1444);
nand U2604 (N_2604,N_1782,N_2282);
nor U2605 (N_2605,N_1711,N_1384);
nor U2606 (N_2606,N_1991,N_1379);
or U2607 (N_2607,N_1880,N_1327);
xnor U2608 (N_2608,N_1265,N_1378);
or U2609 (N_2609,N_2399,N_2166);
nor U2610 (N_2610,N_2312,N_1701);
xnor U2611 (N_2611,N_1222,N_2020);
and U2612 (N_2612,N_1439,N_1553);
nor U2613 (N_2613,N_1864,N_1466);
and U2614 (N_2614,N_1766,N_1964);
nor U2615 (N_2615,N_1331,N_2205);
and U2616 (N_2616,N_2238,N_1853);
and U2617 (N_2617,N_2122,N_2236);
nor U2618 (N_2618,N_2283,N_2039);
nand U2619 (N_2619,N_1211,N_1836);
or U2620 (N_2620,N_2357,N_1614);
or U2621 (N_2621,N_1271,N_1252);
xnor U2622 (N_2622,N_2243,N_1958);
or U2623 (N_2623,N_1938,N_2328);
or U2624 (N_2624,N_1649,N_1297);
or U2625 (N_2625,N_1280,N_1578);
xor U2626 (N_2626,N_1451,N_1232);
nand U2627 (N_2627,N_2006,N_2162);
or U2628 (N_2628,N_1362,N_1539);
nand U2629 (N_2629,N_1417,N_1509);
nand U2630 (N_2630,N_1756,N_2031);
nand U2631 (N_2631,N_1834,N_1940);
nand U2632 (N_2632,N_2212,N_1773);
nand U2633 (N_2633,N_1753,N_2387);
nor U2634 (N_2634,N_2344,N_2320);
nor U2635 (N_2635,N_1640,N_2131);
xor U2636 (N_2636,N_1744,N_2097);
or U2637 (N_2637,N_1353,N_2080);
nor U2638 (N_2638,N_1851,N_2327);
xnor U2639 (N_2639,N_1656,N_1764);
nand U2640 (N_2640,N_2274,N_2206);
or U2641 (N_2641,N_1318,N_1435);
nand U2642 (N_2642,N_2315,N_1955);
nand U2643 (N_2643,N_1648,N_1231);
xnor U2644 (N_2644,N_1634,N_2029);
xnor U2645 (N_2645,N_2234,N_2392);
and U2646 (N_2646,N_1422,N_1847);
and U2647 (N_2647,N_1671,N_2143);
nand U2648 (N_2648,N_2087,N_2201);
nand U2649 (N_2649,N_1814,N_1273);
or U2650 (N_2650,N_2334,N_1436);
nor U2651 (N_2651,N_2010,N_1657);
and U2652 (N_2652,N_1810,N_1413);
or U2653 (N_2653,N_2157,N_1781);
or U2654 (N_2654,N_2314,N_1454);
xnor U2655 (N_2655,N_2088,N_1825);
or U2656 (N_2656,N_2298,N_1519);
nor U2657 (N_2657,N_1583,N_1550);
xor U2658 (N_2658,N_2009,N_1524);
xor U2659 (N_2659,N_2018,N_1959);
nor U2660 (N_2660,N_1783,N_2311);
xnor U2661 (N_2661,N_1636,N_1279);
nand U2662 (N_2662,N_1920,N_1867);
nor U2663 (N_2663,N_1855,N_1799);
or U2664 (N_2664,N_1985,N_1381);
nand U2665 (N_2665,N_2318,N_2197);
or U2666 (N_2666,N_2104,N_1912);
xor U2667 (N_2667,N_1393,N_1398);
or U2668 (N_2668,N_1935,N_2091);
xnor U2669 (N_2669,N_2326,N_1632);
nor U2670 (N_2670,N_2183,N_1486);
xnor U2671 (N_2671,N_1213,N_2343);
xor U2672 (N_2672,N_1821,N_2149);
or U2673 (N_2673,N_2204,N_2036);
and U2674 (N_2674,N_2113,N_2115);
or U2675 (N_2675,N_2185,N_2067);
nor U2676 (N_2676,N_1722,N_1703);
nor U2677 (N_2677,N_2008,N_1401);
or U2678 (N_2678,N_1859,N_1976);
or U2679 (N_2679,N_2365,N_1404);
and U2680 (N_2680,N_1549,N_2188);
nor U2681 (N_2681,N_2278,N_1577);
nor U2682 (N_2682,N_1575,N_2301);
or U2683 (N_2683,N_1804,N_1568);
nand U2684 (N_2684,N_1535,N_1973);
and U2685 (N_2685,N_1679,N_1465);
and U2686 (N_2686,N_1307,N_1248);
xor U2687 (N_2687,N_1416,N_1918);
nand U2688 (N_2688,N_2082,N_1511);
or U2689 (N_2689,N_1597,N_1459);
or U2690 (N_2690,N_2214,N_1212);
and U2691 (N_2691,N_2226,N_1294);
and U2692 (N_2692,N_1452,N_1505);
nor U2693 (N_2693,N_1717,N_2281);
xor U2694 (N_2694,N_1496,N_1680);
nor U2695 (N_2695,N_1882,N_1552);
and U2696 (N_2696,N_1368,N_2286);
nand U2697 (N_2697,N_1876,N_1669);
xor U2698 (N_2698,N_1803,N_1491);
nand U2699 (N_2699,N_1798,N_1606);
or U2700 (N_2700,N_2277,N_2128);
xnor U2701 (N_2701,N_1889,N_1933);
nand U2702 (N_2702,N_2062,N_2179);
xor U2703 (N_2703,N_1993,N_2145);
nand U2704 (N_2704,N_1652,N_1544);
xnor U2705 (N_2705,N_1263,N_1979);
nor U2706 (N_2706,N_1898,N_2330);
xnor U2707 (N_2707,N_2114,N_1739);
and U2708 (N_2708,N_1678,N_1471);
or U2709 (N_2709,N_1747,N_2136);
nor U2710 (N_2710,N_1208,N_2060);
xor U2711 (N_2711,N_2014,N_2300);
xnor U2712 (N_2712,N_1224,N_1545);
nor U2713 (N_2713,N_1487,N_1745);
and U2714 (N_2714,N_1662,N_2033);
nand U2715 (N_2715,N_1694,N_1695);
or U2716 (N_2716,N_1239,N_1570);
or U2717 (N_2717,N_1408,N_1369);
xor U2718 (N_2718,N_1827,N_2085);
nor U2719 (N_2719,N_1529,N_1884);
or U2720 (N_2720,N_1317,N_1909);
xor U2721 (N_2721,N_1743,N_2134);
and U2722 (N_2722,N_1342,N_2181);
and U2723 (N_2723,N_1724,N_2347);
or U2724 (N_2724,N_1666,N_1683);
nor U2725 (N_2725,N_2164,N_2200);
or U2726 (N_2726,N_1651,N_1592);
and U2727 (N_2727,N_2186,N_1844);
and U2728 (N_2728,N_1984,N_2351);
xnor U2729 (N_2729,N_1883,N_2397);
and U2730 (N_2730,N_1895,N_2398);
or U2731 (N_2731,N_1244,N_1400);
nor U2732 (N_2732,N_1341,N_1832);
and U2733 (N_2733,N_1473,N_2335);
nor U2734 (N_2734,N_1801,N_2217);
nor U2735 (N_2735,N_1727,N_1220);
nand U2736 (N_2736,N_2220,N_2240);
or U2737 (N_2737,N_1677,N_1292);
and U2738 (N_2738,N_1978,N_2174);
or U2739 (N_2739,N_2141,N_1253);
nor U2740 (N_2740,N_1664,N_2184);
nor U2741 (N_2741,N_1893,N_1478);
and U2742 (N_2742,N_2195,N_1593);
and U2743 (N_2743,N_1757,N_2132);
and U2744 (N_2744,N_1809,N_1586);
xor U2745 (N_2745,N_1712,N_1971);
nand U2746 (N_2746,N_1481,N_2041);
nand U2747 (N_2747,N_1808,N_2069);
nor U2748 (N_2748,N_2322,N_1530);
xor U2749 (N_2749,N_1707,N_2159);
or U2750 (N_2750,N_2079,N_2383);
and U2751 (N_2751,N_1225,N_2382);
or U2752 (N_2752,N_1896,N_2305);
and U2753 (N_2753,N_1907,N_1293);
nand U2754 (N_2754,N_1300,N_1407);
nor U2755 (N_2755,N_2395,N_1688);
nand U2756 (N_2756,N_1512,N_1434);
and U2757 (N_2757,N_2248,N_1623);
nand U2758 (N_2758,N_1295,N_1394);
nand U2759 (N_2759,N_1395,N_1276);
xor U2760 (N_2760,N_1437,N_1667);
or U2761 (N_2761,N_1285,N_1464);
nand U2762 (N_2762,N_1785,N_1348);
nand U2763 (N_2763,N_1759,N_1337);
nor U2764 (N_2764,N_1514,N_2139);
xnor U2765 (N_2765,N_1924,N_1805);
or U2766 (N_2766,N_1968,N_1528);
xor U2767 (N_2767,N_2182,N_1691);
nand U2768 (N_2768,N_1462,N_1392);
nor U2769 (N_2769,N_1558,N_1742);
nor U2770 (N_2770,N_1713,N_2268);
xnor U2771 (N_2771,N_2098,N_1216);
or U2772 (N_2772,N_2384,N_1607);
or U2773 (N_2773,N_1321,N_1762);
or U2774 (N_2774,N_1936,N_1828);
and U2775 (N_2775,N_2218,N_1463);
and U2776 (N_2776,N_2308,N_1467);
xor U2777 (N_2777,N_1347,N_1446);
and U2778 (N_2778,N_2057,N_1965);
xnor U2779 (N_2779,N_2239,N_1226);
nand U2780 (N_2780,N_1230,N_1719);
or U2781 (N_2781,N_2171,N_2237);
or U2782 (N_2782,N_1983,N_1787);
xor U2783 (N_2783,N_2325,N_1371);
nand U2784 (N_2784,N_1686,N_1599);
nand U2785 (N_2785,N_1281,N_2047);
and U2786 (N_2786,N_1402,N_1674);
xnor U2787 (N_2787,N_1838,N_1732);
nand U2788 (N_2788,N_1455,N_1311);
xor U2789 (N_2789,N_1538,N_2123);
nand U2790 (N_2790,N_1406,N_1335);
nor U2791 (N_2791,N_2349,N_2090);
nor U2792 (N_2792,N_1274,N_1480);
or U2793 (N_2793,N_2193,N_1405);
nand U2794 (N_2794,N_1830,N_1813);
and U2795 (N_2795,N_1235,N_1772);
nand U2796 (N_2796,N_1555,N_1943);
xor U2797 (N_2797,N_1997,N_1917);
nor U2798 (N_2798,N_1360,N_1412);
or U2799 (N_2799,N_1266,N_2133);
or U2800 (N_2800,N_2030,N_2261);
xor U2801 (N_2801,N_1661,N_2255);
and U2802 (N_2802,N_1345,N_1581);
or U2803 (N_2803,N_1977,N_2251);
and U2804 (N_2804,N_1340,N_1650);
and U2805 (N_2805,N_1507,N_2394);
nor U2806 (N_2806,N_2058,N_1728);
nor U2807 (N_2807,N_1299,N_2376);
xor U2808 (N_2808,N_1430,N_1981);
nor U2809 (N_2809,N_2068,N_1826);
and U2810 (N_2810,N_1868,N_1733);
xor U2811 (N_2811,N_2313,N_2094);
or U2812 (N_2812,N_1698,N_1992);
nor U2813 (N_2813,N_1849,N_1644);
nor U2814 (N_2814,N_2190,N_1840);
nor U2815 (N_2815,N_1839,N_2295);
xor U2816 (N_2816,N_1492,N_1816);
nor U2817 (N_2817,N_1604,N_2375);
nand U2818 (N_2818,N_1872,N_2307);
and U2819 (N_2819,N_1223,N_2025);
nor U2820 (N_2820,N_1305,N_1309);
xnor U2821 (N_2821,N_2390,N_2135);
or U2822 (N_2822,N_1672,N_1888);
and U2823 (N_2823,N_1858,N_1427);
or U2824 (N_2824,N_2096,N_1899);
nand U2825 (N_2825,N_2252,N_1349);
nand U2826 (N_2826,N_1901,N_1533);
and U2827 (N_2827,N_1428,N_1690);
nor U2828 (N_2828,N_1871,N_1229);
and U2829 (N_2829,N_1551,N_1886);
and U2830 (N_2830,N_2203,N_1676);
or U2831 (N_2831,N_2207,N_1468);
nor U2832 (N_2832,N_1714,N_2170);
xnor U2833 (N_2833,N_2367,N_1289);
and U2834 (N_2834,N_2172,N_2341);
and U2835 (N_2835,N_1415,N_1202);
nor U2836 (N_2836,N_1716,N_2165);
or U2837 (N_2837,N_1461,N_1457);
and U2838 (N_2838,N_1780,N_1998);
and U2839 (N_2839,N_2095,N_1957);
and U2840 (N_2840,N_1215,N_1768);
and U2841 (N_2841,N_1910,N_1261);
nor U2842 (N_2842,N_2070,N_2155);
nand U2843 (N_2843,N_1387,N_1322);
nand U2844 (N_2844,N_2163,N_1522);
nand U2845 (N_2845,N_1494,N_1525);
nand U2846 (N_2846,N_1835,N_1706);
xnor U2847 (N_2847,N_1939,N_1902);
and U2848 (N_2848,N_1380,N_1344);
nand U2849 (N_2849,N_1547,N_2147);
or U2850 (N_2850,N_1684,N_1818);
and U2851 (N_2851,N_1646,N_1516);
nand U2852 (N_2852,N_1352,N_1944);
nand U2853 (N_2853,N_2038,N_2285);
and U2854 (N_2854,N_2191,N_2293);
xor U2855 (N_2855,N_2272,N_2361);
xor U2856 (N_2856,N_1204,N_1618);
and U2857 (N_2857,N_1718,N_1355);
and U2858 (N_2858,N_1815,N_2158);
nand U2859 (N_2859,N_2329,N_1251);
xor U2860 (N_2860,N_1284,N_1723);
nor U2861 (N_2861,N_2109,N_2385);
nor U2862 (N_2862,N_1784,N_1495);
nand U2863 (N_2863,N_2034,N_1693);
nand U2864 (N_2864,N_1445,N_2202);
and U2865 (N_2865,N_2024,N_1654);
or U2866 (N_2866,N_2249,N_2048);
nand U2867 (N_2867,N_1343,N_1515);
nor U2868 (N_2868,N_1423,N_1866);
and U2869 (N_2869,N_1214,N_1635);
or U2870 (N_2870,N_1645,N_1460);
nand U2871 (N_2871,N_2013,N_2144);
xnor U2872 (N_2872,N_2150,N_1926);
nand U2873 (N_2873,N_2333,N_1850);
and U2874 (N_2874,N_1358,N_1675);
nand U2875 (N_2875,N_1334,N_1763);
and U2876 (N_2876,N_1589,N_1370);
or U2877 (N_2877,N_2021,N_1332);
nand U2878 (N_2878,N_1900,N_1616);
nor U2879 (N_2879,N_1580,N_2059);
xnor U2880 (N_2880,N_1277,N_2142);
nand U2881 (N_2881,N_1986,N_2271);
nand U2882 (N_2882,N_2256,N_1906);
and U2883 (N_2883,N_1854,N_1241);
nor U2884 (N_2884,N_1560,N_1922);
xnor U2885 (N_2885,N_1298,N_2119);
and U2886 (N_2886,N_1518,N_1200);
and U2887 (N_2887,N_1817,N_2092);
nand U2888 (N_2888,N_1904,N_1308);
xnor U2889 (N_2889,N_2360,N_1324);
and U2890 (N_2890,N_1288,N_1710);
nand U2891 (N_2891,N_1831,N_2189);
nor U2892 (N_2892,N_1585,N_2222);
nand U2893 (N_2893,N_1562,N_1477);
and U2894 (N_2894,N_2263,N_1999);
nor U2895 (N_2895,N_1796,N_1841);
nor U2896 (N_2896,N_2187,N_1776);
nand U2897 (N_2897,N_2338,N_2198);
nor U2898 (N_2898,N_1860,N_1256);
and U2899 (N_2899,N_2050,N_1653);
and U2900 (N_2900,N_1221,N_2194);
or U2901 (N_2901,N_1875,N_1934);
nand U2902 (N_2902,N_1961,N_1615);
and U2903 (N_2903,N_1765,N_2083);
nor U2904 (N_2904,N_1330,N_2053);
xnor U2905 (N_2905,N_2232,N_1741);
nand U2906 (N_2906,N_1700,N_1829);
or U2907 (N_2907,N_2346,N_1563);
and U2908 (N_2908,N_2065,N_1421);
or U2909 (N_2909,N_1911,N_1696);
xnor U2910 (N_2910,N_1315,N_1476);
nor U2911 (N_2911,N_2074,N_2192);
and U2912 (N_2912,N_1236,N_2127);
xor U2913 (N_2913,N_1595,N_1611);
and U2914 (N_2914,N_1484,N_2116);
nor U2915 (N_2915,N_1228,N_2178);
xor U2916 (N_2916,N_2130,N_1891);
nor U2917 (N_2917,N_2169,N_1952);
xnor U2918 (N_2918,N_2052,N_1217);
xnor U2919 (N_2919,N_2043,N_1499);
nor U2920 (N_2920,N_1338,N_1837);
and U2921 (N_2921,N_1339,N_2253);
or U2922 (N_2922,N_1769,N_1927);
nand U2923 (N_2923,N_2389,N_1954);
nor U2924 (N_2924,N_1531,N_2076);
and U2925 (N_2925,N_1750,N_1843);
or U2926 (N_2926,N_1237,N_1897);
xor U2927 (N_2927,N_2120,N_1542);
nor U2928 (N_2928,N_2244,N_2258);
nor U2929 (N_2929,N_2161,N_2242);
nor U2930 (N_2930,N_2260,N_1523);
or U2931 (N_2931,N_1947,N_2103);
or U2932 (N_2932,N_1996,N_1613);
nor U2933 (N_2933,N_1605,N_2332);
nand U2934 (N_2934,N_2044,N_2046);
nor U2935 (N_2935,N_1903,N_1601);
or U2936 (N_2936,N_2246,N_1323);
nor U2937 (N_2937,N_2363,N_1429);
or U2938 (N_2938,N_1610,N_1561);
nand U2939 (N_2939,N_1673,N_1482);
xor U2940 (N_2940,N_1878,N_1503);
and U2941 (N_2941,N_1396,N_1885);
nand U2942 (N_2942,N_2228,N_2086);
nor U2943 (N_2943,N_1726,N_2355);
nor U2944 (N_2944,N_1633,N_1242);
nand U2945 (N_2945,N_2100,N_1685);
nand U2946 (N_2946,N_1410,N_2111);
and U2947 (N_2947,N_1824,N_1620);
xnor U2948 (N_2948,N_1373,N_2224);
or U2949 (N_2949,N_2124,N_2110);
xnor U2950 (N_2950,N_2354,N_1255);
and U2951 (N_2951,N_2017,N_1442);
nand U2952 (N_2952,N_2056,N_2373);
nand U2953 (N_2953,N_2011,N_1734);
nor U2954 (N_2954,N_1565,N_1913);
xnor U2955 (N_2955,N_2229,N_2196);
xnor U2956 (N_2956,N_1268,N_1587);
nand U2957 (N_2957,N_1915,N_1681);
xnor U2958 (N_2958,N_1720,N_2032);
or U2959 (N_2959,N_1931,N_2213);
nand U2960 (N_2960,N_1513,N_1203);
or U2961 (N_2961,N_1770,N_2037);
nor U2962 (N_2962,N_1725,N_2000);
nand U2963 (N_2963,N_1209,N_2219);
xor U2964 (N_2964,N_1474,N_1333);
xnor U2965 (N_2965,N_2380,N_1925);
and U2966 (N_2966,N_1735,N_1852);
xnor U2967 (N_2967,N_1359,N_1386);
nand U2968 (N_2968,N_1689,N_2309);
nand U2969 (N_2969,N_2381,N_2106);
or U2970 (N_2970,N_2353,N_2290);
or U2971 (N_2971,N_1546,N_1304);
or U2972 (N_2972,N_1621,N_1928);
xnor U2973 (N_2973,N_1988,N_1572);
nand U2974 (N_2974,N_1823,N_2257);
nand U2975 (N_2975,N_1489,N_1708);
nor U2976 (N_2976,N_1571,N_2297);
nand U2977 (N_2977,N_1526,N_1588);
nor U2978 (N_2978,N_1628,N_1771);
and U2979 (N_2979,N_1641,N_1793);
nor U2980 (N_2980,N_1730,N_2356);
or U2981 (N_2981,N_2105,N_1472);
nand U2982 (N_2982,N_1419,N_1541);
nor U2983 (N_2983,N_2093,N_1980);
or U2984 (N_2984,N_1270,N_2211);
nand U2985 (N_2985,N_1218,N_1659);
and U2986 (N_2986,N_2245,N_1627);
nand U2987 (N_2987,N_2099,N_1510);
nor U2988 (N_2988,N_2223,N_1608);
and U2989 (N_2989,N_1569,N_2306);
nor U2990 (N_2990,N_1921,N_1490);
nor U2991 (N_2991,N_1399,N_1794);
and U2992 (N_2992,N_1767,N_1908);
nor U2993 (N_2993,N_1447,N_2280);
or U2994 (N_2994,N_2042,N_1207);
xor U2995 (N_2995,N_1923,N_2265);
or U2996 (N_2996,N_2175,N_2289);
nor U2997 (N_2997,N_1485,N_2396);
or U2998 (N_2998,N_1873,N_1501);
nand U2999 (N_2999,N_1812,N_1758);
nor U3000 (N_3000,N_1981,N_1219);
xor U3001 (N_3001,N_1295,N_1257);
and U3002 (N_3002,N_2265,N_1721);
or U3003 (N_3003,N_1776,N_1493);
nand U3004 (N_3004,N_2283,N_1204);
and U3005 (N_3005,N_1481,N_1461);
or U3006 (N_3006,N_2042,N_1942);
nor U3007 (N_3007,N_2111,N_2328);
and U3008 (N_3008,N_1270,N_1622);
nand U3009 (N_3009,N_1561,N_2224);
nand U3010 (N_3010,N_1604,N_1431);
or U3011 (N_3011,N_2078,N_2201);
nor U3012 (N_3012,N_1622,N_1637);
nand U3013 (N_3013,N_2289,N_1984);
nand U3014 (N_3014,N_2270,N_2127);
and U3015 (N_3015,N_1256,N_2378);
or U3016 (N_3016,N_1517,N_1402);
nand U3017 (N_3017,N_1583,N_1671);
nand U3018 (N_3018,N_1597,N_1757);
or U3019 (N_3019,N_2086,N_1760);
xor U3020 (N_3020,N_2128,N_1577);
xnor U3021 (N_3021,N_2031,N_2382);
xor U3022 (N_3022,N_1705,N_1384);
nand U3023 (N_3023,N_1824,N_1593);
or U3024 (N_3024,N_1992,N_1819);
and U3025 (N_3025,N_1362,N_1383);
and U3026 (N_3026,N_1301,N_1874);
nor U3027 (N_3027,N_1871,N_1632);
nor U3028 (N_3028,N_1607,N_1558);
or U3029 (N_3029,N_1734,N_2144);
xnor U3030 (N_3030,N_2312,N_1368);
or U3031 (N_3031,N_1484,N_2279);
nor U3032 (N_3032,N_1553,N_1793);
or U3033 (N_3033,N_1551,N_2303);
or U3034 (N_3034,N_1947,N_1828);
nor U3035 (N_3035,N_1391,N_2060);
xor U3036 (N_3036,N_1615,N_2326);
xor U3037 (N_3037,N_1397,N_2375);
nor U3038 (N_3038,N_1770,N_1923);
xnor U3039 (N_3039,N_2062,N_1214);
nor U3040 (N_3040,N_1685,N_2069);
and U3041 (N_3041,N_1333,N_1611);
nor U3042 (N_3042,N_2052,N_1697);
nor U3043 (N_3043,N_2392,N_1779);
xor U3044 (N_3044,N_1232,N_2325);
and U3045 (N_3045,N_1578,N_2017);
xnor U3046 (N_3046,N_2168,N_1757);
and U3047 (N_3047,N_1987,N_1672);
or U3048 (N_3048,N_1605,N_1816);
xnor U3049 (N_3049,N_1714,N_1561);
and U3050 (N_3050,N_1599,N_1915);
or U3051 (N_3051,N_1223,N_1622);
or U3052 (N_3052,N_1450,N_2349);
xnor U3053 (N_3053,N_2328,N_1266);
or U3054 (N_3054,N_1657,N_1909);
and U3055 (N_3055,N_1547,N_1680);
or U3056 (N_3056,N_1548,N_1423);
nor U3057 (N_3057,N_2036,N_1904);
nand U3058 (N_3058,N_1536,N_1631);
xnor U3059 (N_3059,N_1372,N_1392);
xor U3060 (N_3060,N_1422,N_1746);
or U3061 (N_3061,N_1356,N_1958);
nand U3062 (N_3062,N_1604,N_2129);
and U3063 (N_3063,N_2188,N_1830);
nor U3064 (N_3064,N_2239,N_1650);
or U3065 (N_3065,N_1251,N_1456);
nand U3066 (N_3066,N_2068,N_2377);
or U3067 (N_3067,N_2331,N_1839);
nor U3068 (N_3068,N_1863,N_1599);
nor U3069 (N_3069,N_1292,N_1610);
or U3070 (N_3070,N_1304,N_1741);
nand U3071 (N_3071,N_1365,N_1437);
or U3072 (N_3072,N_1255,N_2037);
and U3073 (N_3073,N_2019,N_1427);
nand U3074 (N_3074,N_1449,N_1336);
nand U3075 (N_3075,N_1317,N_2306);
nor U3076 (N_3076,N_1595,N_2220);
or U3077 (N_3077,N_1417,N_1900);
nand U3078 (N_3078,N_1891,N_2121);
xor U3079 (N_3079,N_2180,N_1930);
xnor U3080 (N_3080,N_1634,N_2106);
nor U3081 (N_3081,N_2106,N_1849);
and U3082 (N_3082,N_2288,N_1646);
and U3083 (N_3083,N_2107,N_1630);
nor U3084 (N_3084,N_2268,N_2207);
nand U3085 (N_3085,N_1350,N_1588);
or U3086 (N_3086,N_1543,N_1250);
nand U3087 (N_3087,N_2014,N_1927);
xnor U3088 (N_3088,N_2154,N_2017);
xnor U3089 (N_3089,N_1576,N_1470);
xor U3090 (N_3090,N_1227,N_2202);
xor U3091 (N_3091,N_1765,N_2338);
and U3092 (N_3092,N_1371,N_1624);
nand U3093 (N_3093,N_2254,N_1202);
xnor U3094 (N_3094,N_1493,N_1408);
nor U3095 (N_3095,N_1342,N_1785);
and U3096 (N_3096,N_1379,N_2363);
and U3097 (N_3097,N_2312,N_2171);
and U3098 (N_3098,N_1846,N_1442);
and U3099 (N_3099,N_1279,N_1348);
nand U3100 (N_3100,N_1587,N_1779);
xnor U3101 (N_3101,N_2186,N_1434);
and U3102 (N_3102,N_2365,N_1415);
nor U3103 (N_3103,N_2313,N_1820);
nand U3104 (N_3104,N_2200,N_1655);
nor U3105 (N_3105,N_1581,N_2363);
nor U3106 (N_3106,N_1775,N_1271);
nor U3107 (N_3107,N_1273,N_1915);
and U3108 (N_3108,N_1971,N_1374);
or U3109 (N_3109,N_1711,N_1947);
nor U3110 (N_3110,N_2292,N_2238);
xnor U3111 (N_3111,N_1578,N_1508);
xor U3112 (N_3112,N_1975,N_2008);
or U3113 (N_3113,N_1894,N_2027);
nand U3114 (N_3114,N_1840,N_1374);
xnor U3115 (N_3115,N_1815,N_2255);
and U3116 (N_3116,N_1499,N_2396);
xor U3117 (N_3117,N_1770,N_1548);
and U3118 (N_3118,N_1644,N_1898);
nor U3119 (N_3119,N_2006,N_1650);
nor U3120 (N_3120,N_2362,N_1302);
nor U3121 (N_3121,N_1587,N_1496);
nand U3122 (N_3122,N_2395,N_2130);
nand U3123 (N_3123,N_1517,N_2084);
or U3124 (N_3124,N_2177,N_2192);
xnor U3125 (N_3125,N_1605,N_2395);
and U3126 (N_3126,N_2023,N_1355);
and U3127 (N_3127,N_1452,N_2259);
nor U3128 (N_3128,N_1782,N_1206);
xor U3129 (N_3129,N_1451,N_1411);
nand U3130 (N_3130,N_1650,N_2081);
nand U3131 (N_3131,N_1269,N_2372);
xnor U3132 (N_3132,N_1285,N_1632);
or U3133 (N_3133,N_2220,N_2074);
or U3134 (N_3134,N_2280,N_1229);
nand U3135 (N_3135,N_1610,N_2307);
and U3136 (N_3136,N_2167,N_1734);
xor U3137 (N_3137,N_1848,N_1577);
nand U3138 (N_3138,N_2360,N_1876);
xor U3139 (N_3139,N_1585,N_2287);
nand U3140 (N_3140,N_1927,N_1779);
and U3141 (N_3141,N_1654,N_1557);
and U3142 (N_3142,N_2074,N_2254);
xnor U3143 (N_3143,N_2148,N_1965);
xnor U3144 (N_3144,N_2343,N_1467);
xnor U3145 (N_3145,N_2121,N_1440);
nand U3146 (N_3146,N_2022,N_1668);
and U3147 (N_3147,N_1731,N_1260);
or U3148 (N_3148,N_2308,N_2315);
or U3149 (N_3149,N_1636,N_1314);
or U3150 (N_3150,N_1575,N_1474);
and U3151 (N_3151,N_1503,N_1441);
xnor U3152 (N_3152,N_2300,N_2391);
nand U3153 (N_3153,N_1474,N_2087);
xnor U3154 (N_3154,N_1225,N_1209);
nor U3155 (N_3155,N_1424,N_1816);
nor U3156 (N_3156,N_1205,N_2284);
xnor U3157 (N_3157,N_1780,N_2374);
nand U3158 (N_3158,N_2168,N_2363);
and U3159 (N_3159,N_1730,N_1467);
nand U3160 (N_3160,N_2395,N_1877);
nor U3161 (N_3161,N_1507,N_2137);
nand U3162 (N_3162,N_1641,N_2071);
xnor U3163 (N_3163,N_2047,N_1768);
or U3164 (N_3164,N_2166,N_2392);
and U3165 (N_3165,N_1346,N_1778);
xnor U3166 (N_3166,N_1513,N_1698);
nand U3167 (N_3167,N_2005,N_2164);
nor U3168 (N_3168,N_1432,N_1765);
nand U3169 (N_3169,N_1247,N_2113);
or U3170 (N_3170,N_1851,N_1626);
nand U3171 (N_3171,N_1686,N_2126);
nor U3172 (N_3172,N_2358,N_1665);
nor U3173 (N_3173,N_2020,N_1662);
nor U3174 (N_3174,N_1691,N_1515);
nor U3175 (N_3175,N_2141,N_2230);
xnor U3176 (N_3176,N_2225,N_2351);
xnor U3177 (N_3177,N_1487,N_1321);
nor U3178 (N_3178,N_2373,N_2135);
nor U3179 (N_3179,N_2280,N_1248);
or U3180 (N_3180,N_2119,N_1996);
nand U3181 (N_3181,N_1912,N_1865);
xor U3182 (N_3182,N_2153,N_1587);
nand U3183 (N_3183,N_1762,N_2337);
or U3184 (N_3184,N_1214,N_1524);
and U3185 (N_3185,N_1875,N_1538);
nand U3186 (N_3186,N_2071,N_1311);
xnor U3187 (N_3187,N_1488,N_1840);
or U3188 (N_3188,N_2365,N_1990);
nand U3189 (N_3189,N_2269,N_2165);
and U3190 (N_3190,N_1478,N_1915);
xor U3191 (N_3191,N_1517,N_2229);
and U3192 (N_3192,N_1211,N_1660);
nand U3193 (N_3193,N_1970,N_1688);
nor U3194 (N_3194,N_2076,N_1410);
nand U3195 (N_3195,N_2329,N_2269);
or U3196 (N_3196,N_1378,N_1365);
xnor U3197 (N_3197,N_1293,N_1753);
nor U3198 (N_3198,N_2213,N_1637);
or U3199 (N_3199,N_1357,N_1682);
or U3200 (N_3200,N_2373,N_1522);
xnor U3201 (N_3201,N_1322,N_1720);
and U3202 (N_3202,N_1927,N_2302);
or U3203 (N_3203,N_2303,N_1582);
or U3204 (N_3204,N_2018,N_1945);
nor U3205 (N_3205,N_1553,N_1612);
or U3206 (N_3206,N_1310,N_1981);
or U3207 (N_3207,N_1206,N_1444);
nor U3208 (N_3208,N_1806,N_1260);
nand U3209 (N_3209,N_1814,N_1258);
nor U3210 (N_3210,N_1784,N_2061);
nand U3211 (N_3211,N_2092,N_2340);
and U3212 (N_3212,N_2093,N_2014);
nor U3213 (N_3213,N_2118,N_1493);
xnor U3214 (N_3214,N_2138,N_2381);
xnor U3215 (N_3215,N_1468,N_1579);
or U3216 (N_3216,N_1756,N_1898);
and U3217 (N_3217,N_1573,N_1996);
nand U3218 (N_3218,N_1825,N_1601);
nor U3219 (N_3219,N_2028,N_1303);
nor U3220 (N_3220,N_2250,N_1448);
xor U3221 (N_3221,N_1204,N_1733);
xor U3222 (N_3222,N_1734,N_2267);
xnor U3223 (N_3223,N_2356,N_2308);
xnor U3224 (N_3224,N_2086,N_2333);
nor U3225 (N_3225,N_1383,N_1813);
nor U3226 (N_3226,N_1565,N_2153);
nand U3227 (N_3227,N_1651,N_1752);
or U3228 (N_3228,N_2359,N_1649);
nor U3229 (N_3229,N_1934,N_1976);
nand U3230 (N_3230,N_1728,N_2270);
and U3231 (N_3231,N_1222,N_2231);
nand U3232 (N_3232,N_1665,N_2207);
and U3233 (N_3233,N_1452,N_2235);
and U3234 (N_3234,N_2275,N_1315);
xnor U3235 (N_3235,N_2017,N_1996);
nor U3236 (N_3236,N_1579,N_1900);
and U3237 (N_3237,N_1293,N_2281);
or U3238 (N_3238,N_2080,N_1844);
xor U3239 (N_3239,N_2163,N_2239);
or U3240 (N_3240,N_1603,N_1723);
nor U3241 (N_3241,N_1541,N_1531);
nor U3242 (N_3242,N_1465,N_1690);
nand U3243 (N_3243,N_1816,N_2254);
or U3244 (N_3244,N_2179,N_1777);
xor U3245 (N_3245,N_1893,N_1854);
or U3246 (N_3246,N_1544,N_1683);
xor U3247 (N_3247,N_1656,N_1497);
or U3248 (N_3248,N_1855,N_1295);
and U3249 (N_3249,N_1265,N_2321);
nand U3250 (N_3250,N_2190,N_1873);
or U3251 (N_3251,N_1326,N_1707);
and U3252 (N_3252,N_1902,N_2243);
or U3253 (N_3253,N_1784,N_1470);
or U3254 (N_3254,N_1851,N_2218);
xnor U3255 (N_3255,N_2293,N_2300);
and U3256 (N_3256,N_1296,N_1994);
nand U3257 (N_3257,N_1856,N_1488);
or U3258 (N_3258,N_1546,N_2115);
nor U3259 (N_3259,N_1520,N_1817);
nand U3260 (N_3260,N_1769,N_1857);
and U3261 (N_3261,N_1637,N_1901);
xor U3262 (N_3262,N_2345,N_1322);
nand U3263 (N_3263,N_2009,N_1483);
or U3264 (N_3264,N_1207,N_1960);
and U3265 (N_3265,N_1720,N_1306);
nand U3266 (N_3266,N_1735,N_1455);
or U3267 (N_3267,N_1811,N_1409);
nor U3268 (N_3268,N_1745,N_1414);
or U3269 (N_3269,N_2262,N_2069);
xnor U3270 (N_3270,N_2321,N_1440);
nor U3271 (N_3271,N_1533,N_1289);
and U3272 (N_3272,N_1266,N_1843);
and U3273 (N_3273,N_2243,N_1323);
xnor U3274 (N_3274,N_1392,N_1959);
nor U3275 (N_3275,N_1518,N_1847);
or U3276 (N_3276,N_1742,N_1808);
xor U3277 (N_3277,N_1206,N_1637);
nor U3278 (N_3278,N_1264,N_2322);
nand U3279 (N_3279,N_1325,N_1498);
nand U3280 (N_3280,N_2163,N_1686);
xnor U3281 (N_3281,N_2156,N_1997);
or U3282 (N_3282,N_1234,N_2371);
or U3283 (N_3283,N_2393,N_2358);
nand U3284 (N_3284,N_2320,N_2296);
or U3285 (N_3285,N_1394,N_1796);
xnor U3286 (N_3286,N_1802,N_2018);
xnor U3287 (N_3287,N_2088,N_1489);
and U3288 (N_3288,N_2369,N_1724);
and U3289 (N_3289,N_2172,N_2278);
nand U3290 (N_3290,N_1955,N_1526);
nor U3291 (N_3291,N_1224,N_2009);
or U3292 (N_3292,N_1254,N_1928);
xor U3293 (N_3293,N_2184,N_1376);
xor U3294 (N_3294,N_1789,N_1689);
or U3295 (N_3295,N_1735,N_1959);
xor U3296 (N_3296,N_1969,N_2133);
nand U3297 (N_3297,N_1797,N_2074);
nor U3298 (N_3298,N_1808,N_2044);
xnor U3299 (N_3299,N_1413,N_1597);
nand U3300 (N_3300,N_1508,N_1835);
nor U3301 (N_3301,N_1489,N_1985);
or U3302 (N_3302,N_1324,N_2170);
nand U3303 (N_3303,N_2270,N_2353);
and U3304 (N_3304,N_1881,N_1535);
or U3305 (N_3305,N_1985,N_2371);
nand U3306 (N_3306,N_1510,N_1344);
xnor U3307 (N_3307,N_2376,N_1755);
and U3308 (N_3308,N_2233,N_2101);
and U3309 (N_3309,N_1747,N_1914);
nor U3310 (N_3310,N_1767,N_1950);
nand U3311 (N_3311,N_2212,N_1619);
or U3312 (N_3312,N_1606,N_2092);
nor U3313 (N_3313,N_1282,N_1585);
xor U3314 (N_3314,N_1547,N_1495);
xor U3315 (N_3315,N_1764,N_1733);
xnor U3316 (N_3316,N_1226,N_1383);
xor U3317 (N_3317,N_2259,N_1416);
nor U3318 (N_3318,N_1813,N_2080);
nand U3319 (N_3319,N_1428,N_2102);
nand U3320 (N_3320,N_1395,N_1578);
and U3321 (N_3321,N_1524,N_1323);
xnor U3322 (N_3322,N_1560,N_1259);
or U3323 (N_3323,N_2056,N_1755);
nor U3324 (N_3324,N_2340,N_2349);
nor U3325 (N_3325,N_2241,N_2384);
xnor U3326 (N_3326,N_1725,N_1663);
or U3327 (N_3327,N_1240,N_1872);
nor U3328 (N_3328,N_1288,N_2009);
xnor U3329 (N_3329,N_2322,N_1298);
nand U3330 (N_3330,N_2342,N_2219);
or U3331 (N_3331,N_1845,N_1915);
xnor U3332 (N_3332,N_2057,N_2393);
nor U3333 (N_3333,N_1790,N_2173);
and U3334 (N_3334,N_1300,N_1260);
xnor U3335 (N_3335,N_2052,N_1281);
xor U3336 (N_3336,N_1399,N_1798);
nor U3337 (N_3337,N_2236,N_1920);
nor U3338 (N_3338,N_1453,N_1338);
or U3339 (N_3339,N_1301,N_1884);
and U3340 (N_3340,N_1940,N_2323);
nor U3341 (N_3341,N_1797,N_1524);
xnor U3342 (N_3342,N_2227,N_2320);
or U3343 (N_3343,N_1232,N_1952);
xor U3344 (N_3344,N_1638,N_2097);
or U3345 (N_3345,N_1634,N_2197);
nand U3346 (N_3346,N_2259,N_2393);
xnor U3347 (N_3347,N_1616,N_1941);
and U3348 (N_3348,N_1393,N_1467);
nor U3349 (N_3349,N_1376,N_1875);
nor U3350 (N_3350,N_2107,N_2347);
and U3351 (N_3351,N_2121,N_2335);
and U3352 (N_3352,N_2300,N_1888);
nor U3353 (N_3353,N_1516,N_1871);
nor U3354 (N_3354,N_1917,N_2389);
or U3355 (N_3355,N_2040,N_1431);
nor U3356 (N_3356,N_2260,N_1614);
xnor U3357 (N_3357,N_2214,N_1822);
nor U3358 (N_3358,N_1755,N_1264);
and U3359 (N_3359,N_1478,N_1583);
or U3360 (N_3360,N_1329,N_1634);
or U3361 (N_3361,N_2324,N_2131);
nand U3362 (N_3362,N_1730,N_1643);
or U3363 (N_3363,N_2152,N_2042);
or U3364 (N_3364,N_1918,N_1493);
nor U3365 (N_3365,N_1381,N_1569);
xnor U3366 (N_3366,N_2278,N_1916);
nand U3367 (N_3367,N_1392,N_1350);
xnor U3368 (N_3368,N_1616,N_2314);
or U3369 (N_3369,N_2337,N_1765);
xnor U3370 (N_3370,N_1623,N_1859);
nor U3371 (N_3371,N_1716,N_1514);
nor U3372 (N_3372,N_1287,N_1625);
xor U3373 (N_3373,N_1671,N_1923);
nor U3374 (N_3374,N_1851,N_2262);
and U3375 (N_3375,N_2112,N_1977);
xor U3376 (N_3376,N_1561,N_1993);
nor U3377 (N_3377,N_1425,N_2244);
nor U3378 (N_3378,N_1227,N_1311);
and U3379 (N_3379,N_1417,N_2108);
xor U3380 (N_3380,N_1282,N_1960);
and U3381 (N_3381,N_1689,N_2220);
nor U3382 (N_3382,N_1862,N_1898);
and U3383 (N_3383,N_1245,N_1541);
and U3384 (N_3384,N_1918,N_2105);
xor U3385 (N_3385,N_1516,N_2150);
nand U3386 (N_3386,N_1991,N_1561);
nor U3387 (N_3387,N_1221,N_1214);
nor U3388 (N_3388,N_1620,N_1483);
nor U3389 (N_3389,N_2312,N_1589);
xor U3390 (N_3390,N_1911,N_1441);
and U3391 (N_3391,N_2077,N_1996);
nor U3392 (N_3392,N_1589,N_1795);
nand U3393 (N_3393,N_2043,N_1412);
nand U3394 (N_3394,N_1901,N_1387);
nor U3395 (N_3395,N_1642,N_1615);
nand U3396 (N_3396,N_1272,N_1822);
xnor U3397 (N_3397,N_1406,N_2034);
xnor U3398 (N_3398,N_2185,N_1227);
nand U3399 (N_3399,N_2107,N_1345);
xnor U3400 (N_3400,N_1338,N_2227);
and U3401 (N_3401,N_1804,N_1559);
or U3402 (N_3402,N_1544,N_1676);
nand U3403 (N_3403,N_1785,N_1364);
nor U3404 (N_3404,N_1878,N_1398);
nand U3405 (N_3405,N_1514,N_1201);
xor U3406 (N_3406,N_1637,N_1274);
xnor U3407 (N_3407,N_2215,N_1833);
nor U3408 (N_3408,N_2360,N_1473);
or U3409 (N_3409,N_1317,N_1307);
nand U3410 (N_3410,N_1949,N_2092);
nor U3411 (N_3411,N_2362,N_1258);
nor U3412 (N_3412,N_2366,N_1564);
nor U3413 (N_3413,N_1438,N_1907);
nor U3414 (N_3414,N_1514,N_2390);
nand U3415 (N_3415,N_1755,N_1407);
nor U3416 (N_3416,N_2377,N_1491);
nor U3417 (N_3417,N_1535,N_1855);
and U3418 (N_3418,N_1305,N_2262);
nand U3419 (N_3419,N_1700,N_2335);
nor U3420 (N_3420,N_2216,N_1253);
and U3421 (N_3421,N_2286,N_1643);
nand U3422 (N_3422,N_1646,N_1893);
nor U3423 (N_3423,N_1803,N_1558);
nand U3424 (N_3424,N_1333,N_1890);
nand U3425 (N_3425,N_1470,N_2212);
nand U3426 (N_3426,N_1209,N_2188);
xnor U3427 (N_3427,N_2160,N_1496);
xnor U3428 (N_3428,N_2326,N_2104);
nand U3429 (N_3429,N_1776,N_2135);
nand U3430 (N_3430,N_2047,N_1835);
and U3431 (N_3431,N_1776,N_2281);
or U3432 (N_3432,N_1523,N_2351);
and U3433 (N_3433,N_2262,N_1258);
and U3434 (N_3434,N_1849,N_1845);
and U3435 (N_3435,N_1445,N_2315);
nand U3436 (N_3436,N_2341,N_1443);
xor U3437 (N_3437,N_1678,N_1637);
xor U3438 (N_3438,N_1479,N_1408);
xor U3439 (N_3439,N_1563,N_2360);
or U3440 (N_3440,N_1511,N_1335);
and U3441 (N_3441,N_1332,N_1445);
or U3442 (N_3442,N_1691,N_2081);
xnor U3443 (N_3443,N_1658,N_1729);
or U3444 (N_3444,N_1404,N_2017);
xor U3445 (N_3445,N_1417,N_1419);
nand U3446 (N_3446,N_1681,N_1205);
and U3447 (N_3447,N_1462,N_1636);
and U3448 (N_3448,N_1405,N_1625);
nor U3449 (N_3449,N_1778,N_1835);
xnor U3450 (N_3450,N_1997,N_1643);
nand U3451 (N_3451,N_2207,N_2309);
nand U3452 (N_3452,N_1860,N_1282);
xor U3453 (N_3453,N_1687,N_1829);
and U3454 (N_3454,N_2178,N_1387);
xor U3455 (N_3455,N_1796,N_1566);
xnor U3456 (N_3456,N_1347,N_2208);
xnor U3457 (N_3457,N_2355,N_1538);
xor U3458 (N_3458,N_2223,N_2188);
xnor U3459 (N_3459,N_1549,N_2025);
nand U3460 (N_3460,N_1579,N_2131);
nor U3461 (N_3461,N_1259,N_1200);
nand U3462 (N_3462,N_1361,N_1422);
nor U3463 (N_3463,N_1698,N_1215);
nor U3464 (N_3464,N_1625,N_1481);
or U3465 (N_3465,N_2329,N_1988);
and U3466 (N_3466,N_1996,N_1847);
and U3467 (N_3467,N_1984,N_1223);
xor U3468 (N_3468,N_2159,N_1614);
xor U3469 (N_3469,N_1558,N_1762);
and U3470 (N_3470,N_1914,N_1430);
nor U3471 (N_3471,N_1785,N_2275);
and U3472 (N_3472,N_1496,N_2089);
or U3473 (N_3473,N_1597,N_1294);
and U3474 (N_3474,N_1207,N_2056);
xnor U3475 (N_3475,N_2231,N_2094);
xnor U3476 (N_3476,N_1670,N_1706);
nor U3477 (N_3477,N_1964,N_1351);
nand U3478 (N_3478,N_1206,N_1665);
xor U3479 (N_3479,N_1206,N_1274);
nor U3480 (N_3480,N_1420,N_1433);
xnor U3481 (N_3481,N_1659,N_1687);
and U3482 (N_3482,N_1498,N_1849);
and U3483 (N_3483,N_1505,N_1521);
nor U3484 (N_3484,N_2268,N_1440);
and U3485 (N_3485,N_2355,N_1997);
or U3486 (N_3486,N_1552,N_2072);
nand U3487 (N_3487,N_1273,N_1694);
xnor U3488 (N_3488,N_1820,N_1348);
or U3489 (N_3489,N_2243,N_1760);
nand U3490 (N_3490,N_1985,N_1393);
xor U3491 (N_3491,N_2161,N_1342);
and U3492 (N_3492,N_1269,N_2133);
and U3493 (N_3493,N_2300,N_1378);
xnor U3494 (N_3494,N_1741,N_1992);
or U3495 (N_3495,N_2374,N_2265);
xnor U3496 (N_3496,N_2074,N_2361);
nand U3497 (N_3497,N_2157,N_2395);
or U3498 (N_3498,N_1269,N_2076);
nand U3499 (N_3499,N_1622,N_1431);
nand U3500 (N_3500,N_1303,N_1800);
xor U3501 (N_3501,N_1383,N_1693);
nand U3502 (N_3502,N_1365,N_2125);
or U3503 (N_3503,N_1943,N_1857);
nor U3504 (N_3504,N_1788,N_1224);
or U3505 (N_3505,N_1340,N_1296);
nand U3506 (N_3506,N_1979,N_1540);
or U3507 (N_3507,N_2084,N_1833);
nor U3508 (N_3508,N_1749,N_1348);
and U3509 (N_3509,N_1573,N_2126);
or U3510 (N_3510,N_1664,N_1365);
xor U3511 (N_3511,N_1206,N_2153);
and U3512 (N_3512,N_1827,N_1283);
or U3513 (N_3513,N_1642,N_1766);
nand U3514 (N_3514,N_1318,N_1254);
and U3515 (N_3515,N_1438,N_2019);
xor U3516 (N_3516,N_1205,N_1352);
nand U3517 (N_3517,N_1383,N_1663);
nand U3518 (N_3518,N_2313,N_2349);
and U3519 (N_3519,N_2028,N_1844);
or U3520 (N_3520,N_1617,N_2297);
and U3521 (N_3521,N_2068,N_2204);
xnor U3522 (N_3522,N_2183,N_1260);
nand U3523 (N_3523,N_1952,N_1807);
xor U3524 (N_3524,N_1220,N_1257);
nand U3525 (N_3525,N_1455,N_1742);
or U3526 (N_3526,N_2001,N_1648);
xor U3527 (N_3527,N_1977,N_2370);
nand U3528 (N_3528,N_2304,N_1763);
nand U3529 (N_3529,N_1733,N_1569);
or U3530 (N_3530,N_1824,N_1759);
nand U3531 (N_3531,N_2165,N_2121);
xor U3532 (N_3532,N_1378,N_1811);
nand U3533 (N_3533,N_1480,N_1471);
nand U3534 (N_3534,N_2230,N_1251);
or U3535 (N_3535,N_2053,N_1272);
and U3536 (N_3536,N_1833,N_2089);
xnor U3537 (N_3537,N_1844,N_1888);
and U3538 (N_3538,N_1932,N_1304);
and U3539 (N_3539,N_2158,N_2364);
nand U3540 (N_3540,N_1527,N_1983);
nand U3541 (N_3541,N_2275,N_1258);
and U3542 (N_3542,N_1702,N_1343);
nand U3543 (N_3543,N_2149,N_1989);
xnor U3544 (N_3544,N_1461,N_1592);
xnor U3545 (N_3545,N_2309,N_1919);
xnor U3546 (N_3546,N_1373,N_1696);
xor U3547 (N_3547,N_2214,N_1277);
nand U3548 (N_3548,N_1492,N_2076);
xor U3549 (N_3549,N_1966,N_1703);
nand U3550 (N_3550,N_2371,N_2210);
nor U3551 (N_3551,N_2052,N_1234);
xnor U3552 (N_3552,N_1877,N_1695);
and U3553 (N_3553,N_1949,N_1446);
nand U3554 (N_3554,N_1317,N_1481);
and U3555 (N_3555,N_1332,N_1651);
or U3556 (N_3556,N_1235,N_2368);
xor U3557 (N_3557,N_2029,N_1315);
and U3558 (N_3558,N_1739,N_1281);
xnor U3559 (N_3559,N_1876,N_1501);
xnor U3560 (N_3560,N_2030,N_2226);
nor U3561 (N_3561,N_2207,N_1840);
and U3562 (N_3562,N_1621,N_2190);
and U3563 (N_3563,N_1802,N_2109);
nor U3564 (N_3564,N_1497,N_2395);
or U3565 (N_3565,N_1460,N_2166);
nor U3566 (N_3566,N_2217,N_2165);
or U3567 (N_3567,N_1929,N_1349);
xnor U3568 (N_3568,N_2133,N_1455);
xnor U3569 (N_3569,N_1773,N_1845);
nor U3570 (N_3570,N_1641,N_1646);
or U3571 (N_3571,N_1679,N_1934);
and U3572 (N_3572,N_1406,N_1579);
nand U3573 (N_3573,N_1614,N_1765);
nand U3574 (N_3574,N_1217,N_1397);
xnor U3575 (N_3575,N_1662,N_2171);
nor U3576 (N_3576,N_2283,N_2212);
or U3577 (N_3577,N_1915,N_1426);
nor U3578 (N_3578,N_2046,N_1400);
xnor U3579 (N_3579,N_1610,N_2273);
nand U3580 (N_3580,N_1550,N_1581);
and U3581 (N_3581,N_1703,N_2306);
xnor U3582 (N_3582,N_2383,N_1917);
nor U3583 (N_3583,N_2067,N_2105);
nand U3584 (N_3584,N_2374,N_1544);
nor U3585 (N_3585,N_2369,N_1428);
nor U3586 (N_3586,N_2105,N_1291);
xnor U3587 (N_3587,N_1911,N_2399);
nor U3588 (N_3588,N_1315,N_2113);
or U3589 (N_3589,N_1572,N_1905);
nand U3590 (N_3590,N_1733,N_1806);
nor U3591 (N_3591,N_2285,N_1852);
and U3592 (N_3592,N_1848,N_1285);
nor U3593 (N_3593,N_2345,N_1498);
xor U3594 (N_3594,N_1980,N_1451);
nor U3595 (N_3595,N_1469,N_2281);
xor U3596 (N_3596,N_1211,N_1514);
nor U3597 (N_3597,N_2178,N_1383);
and U3598 (N_3598,N_1400,N_1230);
nand U3599 (N_3599,N_1297,N_2306);
nor U3600 (N_3600,N_2645,N_2706);
and U3601 (N_3601,N_3086,N_2690);
or U3602 (N_3602,N_3576,N_2964);
and U3603 (N_3603,N_2939,N_2979);
nand U3604 (N_3604,N_3052,N_3208);
xor U3605 (N_3605,N_3130,N_3202);
and U3606 (N_3606,N_2998,N_2551);
and U3607 (N_3607,N_2944,N_2684);
nor U3608 (N_3608,N_2489,N_2624);
and U3609 (N_3609,N_3294,N_2679);
nand U3610 (N_3610,N_3488,N_3393);
xnor U3611 (N_3611,N_2416,N_3232);
nor U3612 (N_3612,N_3074,N_2921);
and U3613 (N_3613,N_2932,N_2935);
or U3614 (N_3614,N_2815,N_3476);
nor U3615 (N_3615,N_2731,N_2747);
or U3616 (N_3616,N_2984,N_2759);
or U3617 (N_3617,N_2665,N_2777);
nand U3618 (N_3618,N_2894,N_3186);
nand U3619 (N_3619,N_2622,N_2514);
nor U3620 (N_3620,N_3429,N_3566);
or U3621 (N_3621,N_2830,N_3088);
xnor U3622 (N_3622,N_3360,N_3077);
xnor U3623 (N_3623,N_3594,N_2403);
xnor U3624 (N_3624,N_3326,N_2440);
and U3625 (N_3625,N_2556,N_3554);
nand U3626 (N_3626,N_2816,N_3501);
and U3627 (N_3627,N_2620,N_2574);
or U3628 (N_3628,N_2621,N_2917);
xnor U3629 (N_3629,N_3376,N_3427);
nor U3630 (N_3630,N_3398,N_2829);
nand U3631 (N_3631,N_3569,N_3544);
nor U3632 (N_3632,N_2421,N_2609);
nand U3633 (N_3633,N_2908,N_3371);
or U3634 (N_3634,N_2450,N_3322);
or U3635 (N_3635,N_3076,N_2886);
xor U3636 (N_3636,N_3201,N_2693);
xnor U3637 (N_3637,N_2584,N_2615);
or U3638 (N_3638,N_2666,N_3384);
nand U3639 (N_3639,N_2866,N_2737);
or U3640 (N_3640,N_3518,N_2763);
or U3641 (N_3641,N_3587,N_3014);
or U3642 (N_3642,N_3206,N_2632);
nand U3643 (N_3643,N_2843,N_3457);
or U3644 (N_3644,N_3215,N_2862);
nor U3645 (N_3645,N_3281,N_3072);
and U3646 (N_3646,N_3034,N_3510);
and U3647 (N_3647,N_3081,N_2951);
xor U3648 (N_3648,N_3579,N_2740);
nor U3649 (N_3649,N_2918,N_3597);
and U3650 (N_3650,N_2723,N_2812);
xor U3651 (N_3651,N_2837,N_2699);
or U3652 (N_3652,N_3433,N_3486);
or U3653 (N_3653,N_3599,N_2750);
or U3654 (N_3654,N_3291,N_3330);
or U3655 (N_3655,N_2545,N_2681);
or U3656 (N_3656,N_2425,N_3289);
nor U3657 (N_3657,N_3496,N_3254);
or U3658 (N_3658,N_2923,N_2488);
nor U3659 (N_3659,N_3042,N_3351);
and U3660 (N_3660,N_3468,N_3099);
nor U3661 (N_3661,N_3151,N_2503);
xor U3662 (N_3662,N_2582,N_3475);
nand U3663 (N_3663,N_2871,N_3144);
xor U3664 (N_3664,N_2818,N_2457);
xor U3665 (N_3665,N_3466,N_3142);
or U3666 (N_3666,N_2664,N_2994);
and U3667 (N_3667,N_3116,N_3036);
xor U3668 (N_3668,N_3128,N_2557);
nor U3669 (N_3669,N_3019,N_3020);
nor U3670 (N_3670,N_2965,N_3137);
or U3671 (N_3671,N_3157,N_3032);
xor U3672 (N_3672,N_2641,N_3540);
and U3673 (N_3673,N_3120,N_3568);
nor U3674 (N_3674,N_2889,N_3063);
nor U3675 (N_3675,N_3354,N_3258);
nor U3676 (N_3676,N_3346,N_2771);
and U3677 (N_3677,N_2870,N_3284);
nor U3678 (N_3678,N_3191,N_3494);
nand U3679 (N_3679,N_3175,N_3064);
or U3680 (N_3680,N_3382,N_3506);
xor U3681 (N_3681,N_2784,N_3065);
or U3682 (N_3682,N_2728,N_2509);
xnor U3683 (N_3683,N_3010,N_2607);
nand U3684 (N_3684,N_3362,N_3165);
nor U3685 (N_3685,N_2546,N_2774);
and U3686 (N_3686,N_2564,N_2490);
and U3687 (N_3687,N_2717,N_2492);
or U3688 (N_3688,N_3403,N_3100);
nor U3689 (N_3689,N_2821,N_2419);
or U3690 (N_3690,N_3453,N_2937);
nor U3691 (N_3691,N_3452,N_3177);
or U3692 (N_3692,N_2482,N_3256);
nor U3693 (N_3693,N_3105,N_2903);
nand U3694 (N_3694,N_3567,N_2630);
or U3695 (N_3695,N_2558,N_3425);
nand U3696 (N_3696,N_2594,N_3173);
or U3697 (N_3697,N_3017,N_3269);
and U3698 (N_3698,N_3359,N_3564);
nand U3699 (N_3699,N_2807,N_3514);
and U3700 (N_3700,N_2603,N_2980);
xnor U3701 (N_3701,N_2924,N_2649);
nor U3702 (N_3702,N_2726,N_2606);
nand U3703 (N_3703,N_3111,N_3369);
and U3704 (N_3704,N_2888,N_3027);
nand U3705 (N_3705,N_2700,N_2709);
and U3706 (N_3706,N_2860,N_2651);
and U3707 (N_3707,N_2424,N_2695);
nand U3708 (N_3708,N_2877,N_3218);
xor U3709 (N_3709,N_2741,N_3214);
xor U3710 (N_3710,N_2989,N_3549);
nand U3711 (N_3711,N_2461,N_3419);
xor U3712 (N_3712,N_3227,N_3463);
or U3713 (N_3713,N_3489,N_2780);
xor U3714 (N_3714,N_2782,N_2480);
xor U3715 (N_3715,N_2477,N_3178);
nand U3716 (N_3716,N_2563,N_3041);
and U3717 (N_3717,N_3069,N_2955);
nand U3718 (N_3718,N_2864,N_3230);
nand U3719 (N_3719,N_3029,N_3589);
or U3720 (N_3720,N_2495,N_3181);
nor U3721 (N_3721,N_3028,N_2811);
nand U3722 (N_3722,N_3220,N_2813);
and U3723 (N_3723,N_2978,N_3091);
or U3724 (N_3724,N_3524,N_2902);
nand U3725 (N_3725,N_3412,N_2662);
and U3726 (N_3726,N_3307,N_2948);
or U3727 (N_3727,N_2855,N_3535);
and U3728 (N_3728,N_2547,N_2643);
and U3729 (N_3729,N_2909,N_2688);
nand U3730 (N_3730,N_2460,N_3328);
nor U3731 (N_3731,N_3305,N_2972);
nor U3732 (N_3732,N_2869,N_2443);
xnor U3733 (N_3733,N_3509,N_3456);
and U3734 (N_3734,N_3199,N_3500);
xnor U3735 (N_3735,N_3370,N_3443);
nand U3736 (N_3736,N_3237,N_2960);
and U3737 (N_3737,N_3394,N_3377);
nand U3738 (N_3738,N_3592,N_3113);
or U3739 (N_3739,N_2861,N_3595);
nand U3740 (N_3740,N_3149,N_3536);
nor U3741 (N_3741,N_2840,N_3431);
nor U3742 (N_3742,N_3161,N_3591);
and U3743 (N_3743,N_2444,N_2498);
or U3744 (N_3744,N_3451,N_2687);
and U3745 (N_3745,N_2768,N_2596);
or U3746 (N_3746,N_2507,N_2744);
nand U3747 (N_3747,N_3092,N_3304);
nor U3748 (N_3748,N_2578,N_2758);
nor U3749 (N_3749,N_3170,N_3079);
or U3750 (N_3750,N_3001,N_2954);
and U3751 (N_3751,N_2928,N_2749);
nand U3752 (N_3752,N_3297,N_2966);
xnor U3753 (N_3753,N_2846,N_2483);
xnor U3754 (N_3754,N_2707,N_3174);
or U3755 (N_3755,N_2623,N_2540);
nor U3756 (N_3756,N_3273,N_3096);
or U3757 (N_3757,N_3048,N_3156);
nor U3758 (N_3758,N_2704,N_2531);
and U3759 (N_3759,N_2472,N_2510);
xor U3760 (N_3760,N_3152,N_2549);
and U3761 (N_3761,N_2802,N_2486);
or U3762 (N_3762,N_2414,N_2764);
and U3763 (N_3763,N_3411,N_3288);
or U3764 (N_3764,N_2720,N_2478);
xnor U3765 (N_3765,N_2865,N_3071);
or U3766 (N_3766,N_3490,N_3391);
or U3767 (N_3767,N_3439,N_2828);
xor U3768 (N_3768,N_3428,N_2942);
nand U3769 (N_3769,N_2947,N_2656);
nand U3770 (N_3770,N_3271,N_2445);
or U3771 (N_3771,N_3553,N_2775);
or U3772 (N_3772,N_3250,N_3310);
nand U3773 (N_3773,N_2439,N_3037);
or U3774 (N_3774,N_2613,N_3233);
and U3775 (N_3775,N_2660,N_2742);
nand U3776 (N_3776,N_2827,N_3303);
xnor U3777 (N_3777,N_2867,N_2449);
nand U3778 (N_3778,N_3499,N_3583);
nor U3779 (N_3779,N_3355,N_2801);
nor U3780 (N_3780,N_3213,N_3538);
nor U3781 (N_3781,N_2400,N_2804);
xnor U3782 (N_3782,N_3415,N_2823);
or U3783 (N_3783,N_2410,N_3319);
nor U3784 (N_3784,N_2705,N_3184);
xnor U3785 (N_3785,N_3316,N_3542);
and U3786 (N_3786,N_2712,N_3332);
and U3787 (N_3787,N_3450,N_2868);
nand U3788 (N_3788,N_3240,N_2408);
and U3789 (N_3789,N_3241,N_2970);
or U3790 (N_3790,N_3163,N_3015);
and U3791 (N_3791,N_3030,N_2961);
xor U3792 (N_3792,N_3057,N_2575);
and U3793 (N_3793,N_2646,N_3033);
and U3794 (N_3794,N_3141,N_3278);
or U3795 (N_3795,N_3314,N_3083);
nand U3796 (N_3796,N_3372,N_2916);
nor U3797 (N_3797,N_3378,N_2891);
nor U3798 (N_3798,N_3302,N_2438);
or U3799 (N_3799,N_2958,N_3194);
xnor U3800 (N_3800,N_2698,N_2415);
nor U3801 (N_3801,N_2748,N_3123);
xor U3802 (N_3802,N_2999,N_3352);
or U3803 (N_3803,N_2733,N_2661);
and U3804 (N_3804,N_2967,N_2422);
and U3805 (N_3805,N_3570,N_3508);
xnor U3806 (N_3806,N_3051,N_3262);
xor U3807 (N_3807,N_2962,N_3530);
xor U3808 (N_3808,N_3502,N_2428);
nor U3809 (N_3809,N_2929,N_3270);
and U3810 (N_3810,N_2859,N_2466);
xor U3811 (N_3811,N_3136,N_2919);
or U3812 (N_3812,N_2675,N_3059);
xnor U3813 (N_3813,N_3541,N_3021);
and U3814 (N_3814,N_2853,N_2655);
nor U3815 (N_3815,N_2659,N_2587);
nor U3816 (N_3816,N_3217,N_2423);
nand U3817 (N_3817,N_3343,N_2647);
nor U3818 (N_3818,N_3062,N_2756);
nor U3819 (N_3819,N_2590,N_2734);
and U3820 (N_3820,N_3402,N_2875);
and U3821 (N_3821,N_2691,N_3045);
or U3822 (N_3822,N_2455,N_3460);
xor U3823 (N_3823,N_3388,N_2579);
nor U3824 (N_3824,N_2442,N_2934);
and U3825 (N_3825,N_2599,N_2931);
xnor U3826 (N_3826,N_3498,N_3375);
nand U3827 (N_3827,N_2475,N_3462);
nand U3828 (N_3828,N_3590,N_2897);
nor U3829 (N_3829,N_3066,N_2678);
nor U3830 (N_3830,N_2710,N_3164);
nand U3831 (N_3831,N_2792,N_2560);
or U3832 (N_3832,N_3018,N_3287);
nor U3833 (N_3833,N_2516,N_3108);
nor U3834 (N_3834,N_3110,N_2793);
or U3835 (N_3835,N_2494,N_3012);
xnor U3836 (N_3836,N_3275,N_2533);
nand U3837 (N_3837,N_3242,N_3293);
or U3838 (N_3838,N_2773,N_2508);
nor U3839 (N_3839,N_3171,N_2990);
nand U3840 (N_3840,N_3285,N_3195);
or U3841 (N_3841,N_2500,N_3395);
nand U3842 (N_3842,N_3449,N_2639);
nand U3843 (N_3843,N_2676,N_3121);
xnor U3844 (N_3844,N_3147,N_2436);
nand U3845 (N_3845,N_3166,N_2765);
nand U3846 (N_3846,N_2476,N_2406);
or U3847 (N_3847,N_2640,N_3264);
nor U3848 (N_3848,N_2798,N_2404);
nand U3849 (N_3849,N_3219,N_2454);
or U3850 (N_3850,N_2588,N_3356);
xnor U3851 (N_3851,N_3272,N_3532);
or U3852 (N_3852,N_3228,N_3454);
nand U3853 (N_3853,N_3521,N_2799);
xor U3854 (N_3854,N_3537,N_3068);
xor U3855 (N_3855,N_3248,N_2402);
and U3856 (N_3856,N_2993,N_3574);
xnor U3857 (N_3857,N_3117,N_2506);
nand U3858 (N_3858,N_3090,N_3131);
xor U3859 (N_3859,N_3257,N_3323);
xor U3860 (N_3860,N_3246,N_3389);
nand U3861 (N_3861,N_3252,N_3448);
nand U3862 (N_3862,N_2692,N_2435);
or U3863 (N_3863,N_3085,N_2568);
nand U3864 (N_3864,N_3479,N_3338);
nand U3865 (N_3865,N_3279,N_3480);
nor U3866 (N_3866,N_3469,N_2434);
xor U3867 (N_3867,N_2890,N_2790);
nor U3868 (N_3868,N_3047,N_3094);
nor U3869 (N_3869,N_3575,N_2608);
or U3870 (N_3870,N_2496,N_2635);
xnor U3871 (N_3871,N_3158,N_2851);
or U3872 (N_3872,N_2760,N_3512);
or U3873 (N_3873,N_3588,N_3515);
and U3874 (N_3874,N_2576,N_2987);
nand U3875 (N_3875,N_3404,N_3317);
nor U3876 (N_3876,N_2626,N_2803);
nor U3877 (N_3877,N_2601,N_2854);
or U3878 (N_3878,N_3561,N_2631);
or U3879 (N_3879,N_3473,N_3421);
or U3880 (N_3880,N_3482,N_3109);
or U3881 (N_3881,N_3301,N_2776);
or U3882 (N_3882,N_2432,N_2633);
nor U3883 (N_3883,N_2513,N_3337);
or U3884 (N_3884,N_2910,N_2783);
nor U3885 (N_3885,N_3078,N_3331);
nand U3886 (N_3886,N_2766,N_3523);
and U3887 (N_3887,N_3299,N_2441);
xnor U3888 (N_3888,N_3358,N_3552);
or U3889 (N_3889,N_3003,N_2473);
and U3890 (N_3890,N_3245,N_3408);
and U3891 (N_3891,N_2612,N_2767);
or U3892 (N_3892,N_3527,N_3060);
xor U3893 (N_3893,N_3207,N_2992);
nor U3894 (N_3894,N_2686,N_2976);
nand U3895 (N_3895,N_2674,N_2856);
nand U3896 (N_3896,N_3212,N_3209);
nand U3897 (N_3897,N_3286,N_3320);
nand U3898 (N_3898,N_3432,N_2627);
nor U3899 (N_3899,N_3190,N_2570);
and U3900 (N_3900,N_2462,N_2893);
nand U3901 (N_3901,N_2447,N_2810);
or U3902 (N_3902,N_3283,N_2673);
xnor U3903 (N_3903,N_3417,N_2788);
and U3904 (N_3904,N_2880,N_3183);
nor U3905 (N_3905,N_2927,N_3438);
xor U3906 (N_3906,N_3519,N_3004);
or U3907 (N_3907,N_3361,N_3216);
and U3908 (N_3908,N_2484,N_3268);
nor U3909 (N_3909,N_3545,N_3298);
and U3910 (N_3910,N_3344,N_2427);
and U3911 (N_3911,N_3089,N_3347);
nand U3912 (N_3912,N_2562,N_2718);
xor U3913 (N_3913,N_3464,N_3087);
or U3914 (N_3914,N_3381,N_3407);
and U3915 (N_3915,N_2420,N_2725);
and U3916 (N_3916,N_2650,N_3016);
xor U3917 (N_3917,N_3026,N_2940);
xnor U3918 (N_3918,N_2878,N_2833);
or U3919 (N_3919,N_3374,N_3075);
and U3920 (N_3920,N_2431,N_2795);
and U3921 (N_3921,N_3380,N_2952);
xnor U3922 (N_3922,N_3477,N_2504);
xnor U3923 (N_3923,N_3290,N_3023);
or U3924 (N_3924,N_3483,N_3097);
and U3925 (N_3925,N_2571,N_3396);
or U3926 (N_3926,N_2922,N_3148);
xnor U3927 (N_3927,N_2913,N_3253);
xor U3928 (N_3928,N_3572,N_2754);
and U3929 (N_3929,N_3334,N_3410);
nor U3930 (N_3930,N_3373,N_3321);
xor U3931 (N_3931,N_2644,N_2702);
nor U3932 (N_3932,N_2629,N_3481);
and U3933 (N_3933,N_2604,N_2835);
and U3934 (N_3934,N_3160,N_2806);
nor U3935 (N_3935,N_2453,N_2413);
nor U3936 (N_3936,N_3363,N_3470);
xnor U3937 (N_3937,N_3584,N_2511);
or U3938 (N_3938,N_2523,N_3390);
and U3939 (N_3939,N_2505,N_2914);
and U3940 (N_3940,N_3211,N_3366);
nor U3941 (N_3941,N_2518,N_3399);
xnor U3942 (N_3942,N_2470,N_2525);
and U3943 (N_3943,N_3556,N_2452);
xnor U3944 (N_3944,N_3102,N_2501);
or U3945 (N_3945,N_2642,N_2719);
or U3946 (N_3946,N_3467,N_3577);
nand U3947 (N_3947,N_3169,N_3555);
or U3948 (N_3948,N_3424,N_3571);
xor U3949 (N_3949,N_2479,N_2682);
and U3950 (N_3950,N_3365,N_2986);
xor U3951 (N_3951,N_2493,N_3005);
and U3952 (N_3952,N_2834,N_3259);
nor U3953 (N_3953,N_2600,N_3277);
xnor U3954 (N_3954,N_3188,N_3441);
or U3955 (N_3955,N_2899,N_2527);
or U3956 (N_3956,N_2538,N_3367);
and U3957 (N_3957,N_3397,N_3383);
nor U3958 (N_3958,N_3533,N_2822);
and U3959 (N_3959,N_3180,N_2554);
nor U3960 (N_3960,N_2945,N_2657);
xor U3961 (N_3961,N_3311,N_3444);
xnor U3962 (N_3962,N_2592,N_3251);
nand U3963 (N_3963,N_2654,N_3392);
and U3964 (N_3964,N_3098,N_2915);
nand U3965 (N_3965,N_3414,N_3560);
and U3966 (N_3966,N_3229,N_3458);
xnor U3967 (N_3967,N_2925,N_2819);
xnor U3968 (N_3968,N_3073,N_3582);
and U3969 (N_3969,N_3282,N_3276);
nor U3970 (N_3970,N_3104,N_3009);
xor U3971 (N_3971,N_2667,N_2991);
or U3972 (N_3972,N_2529,N_3324);
or U3973 (N_3973,N_2985,N_2845);
nand U3974 (N_3974,N_2573,N_2949);
and U3975 (N_3975,N_2729,N_2714);
or U3976 (N_3976,N_3422,N_2971);
nor U3977 (N_3977,N_2789,N_3006);
xnor U3978 (N_3978,N_2652,N_2904);
and U3979 (N_3979,N_2614,N_2738);
nor U3980 (N_3980,N_2743,N_2543);
and U3981 (N_3981,N_3061,N_2745);
nor U3982 (N_3982,N_3058,N_3082);
or U3983 (N_3983,N_2561,N_3562);
nor U3984 (N_3984,N_2672,N_2786);
nor U3985 (N_3985,N_3146,N_2975);
and U3986 (N_3986,N_2814,N_3013);
nor U3987 (N_3987,N_3497,N_2581);
or U3988 (N_3988,N_2724,N_2872);
nand U3989 (N_3989,N_2732,N_2959);
xor U3990 (N_3990,N_3124,N_2553);
or U3991 (N_3991,N_2826,N_3247);
nand U3992 (N_3992,N_3416,N_2446);
nand U3993 (N_3993,N_2580,N_3127);
and U3994 (N_3994,N_3487,N_2566);
nand U3995 (N_3995,N_3106,N_3231);
nor U3996 (N_3996,N_3260,N_2694);
nor U3997 (N_3997,N_2882,N_3516);
xor U3998 (N_3998,N_2938,N_3011);
xnor U3999 (N_3999,N_2685,N_3405);
and U4000 (N_4000,N_2739,N_3505);
xnor U4001 (N_4001,N_2471,N_2418);
nand U4002 (N_4002,N_3565,N_2499);
xor U4003 (N_4003,N_2524,N_3134);
nor U4004 (N_4004,N_2838,N_3308);
or U4005 (N_4005,N_2648,N_2973);
and U4006 (N_4006,N_3126,N_2794);
nor U4007 (N_4007,N_3187,N_3563);
nor U4008 (N_4008,N_2634,N_3244);
nor U4009 (N_4009,N_2831,N_2817);
and U4010 (N_4010,N_2669,N_2953);
nor U4011 (N_4011,N_2583,N_3546);
xnor U4012 (N_4012,N_3197,N_3484);
nor U4013 (N_4013,N_2873,N_2497);
xnor U4014 (N_4014,N_3135,N_3493);
nor U4015 (N_4015,N_3526,N_2863);
and U4016 (N_4016,N_3239,N_2805);
nor U4017 (N_4017,N_2437,N_3593);
and U4018 (N_4018,N_3353,N_3379);
nor U4019 (N_4019,N_2746,N_2521);
or U4020 (N_4020,N_3312,N_2933);
or U4021 (N_4021,N_2487,N_3038);
and U4022 (N_4022,N_3243,N_3296);
xnor U4023 (N_4023,N_3053,N_2848);
and U4024 (N_4024,N_2946,N_3333);
xor U4025 (N_4025,N_2433,N_2901);
or U4026 (N_4026,N_3295,N_2956);
and U4027 (N_4027,N_3035,N_2548);
xnor U4028 (N_4028,N_2544,N_3315);
and U4029 (N_4029,N_3543,N_3387);
nand U4030 (N_4030,N_2820,N_2930);
and U4031 (N_4031,N_3436,N_3226);
nor U4032 (N_4032,N_3409,N_3386);
and U4033 (N_4033,N_2824,N_2520);
nor U4034 (N_4034,N_2589,N_2950);
nor U4035 (N_4035,N_2565,N_2905);
nor U4036 (N_4036,N_3522,N_3551);
and U4037 (N_4037,N_3155,N_2997);
and U4038 (N_4038,N_3235,N_2519);
xnor U4039 (N_4039,N_2658,N_3557);
or U4040 (N_4040,N_3309,N_2572);
xor U4041 (N_4041,N_3531,N_2892);
nand U4042 (N_4042,N_3204,N_2638);
nor U4043 (N_4043,N_2761,N_2577);
or U4044 (N_4044,N_3313,N_2456);
xor U4045 (N_4045,N_3492,N_3598);
or U4046 (N_4046,N_3573,N_2405);
nand U4047 (N_4047,N_3129,N_3140);
xor U4048 (N_4048,N_3507,N_3054);
and U4049 (N_4049,N_2491,N_2617);
and U4050 (N_4050,N_2844,N_2464);
or U4051 (N_4051,N_2458,N_2598);
or U4052 (N_4052,N_3385,N_3084);
xnor U4053 (N_4053,N_3031,N_2515);
nor U4054 (N_4054,N_2762,N_3223);
or U4055 (N_4055,N_3503,N_2781);
or U4056 (N_4056,N_2809,N_2883);
or U4057 (N_4057,N_3525,N_3093);
and U4058 (N_4058,N_3154,N_2593);
nor U4059 (N_4059,N_3472,N_3274);
nand U4060 (N_4060,N_3118,N_3025);
nand U4061 (N_4061,N_2481,N_2534);
xor U4062 (N_4062,N_2896,N_3044);
nor U4063 (N_4063,N_3133,N_3517);
or U4064 (N_4064,N_2982,N_2683);
nor U4065 (N_4065,N_2969,N_3349);
xnor U4066 (N_4066,N_2605,N_3095);
nor U4067 (N_4067,N_2907,N_3143);
xnor U4068 (N_4068,N_3039,N_3406);
nand U4069 (N_4069,N_2800,N_2757);
nor U4070 (N_4070,N_3168,N_3357);
nor U4071 (N_4071,N_2730,N_2858);
or U4072 (N_4072,N_2895,N_2668);
nor U4073 (N_4073,N_3504,N_2701);
and U4074 (N_4074,N_2996,N_2736);
and U4075 (N_4075,N_2451,N_3446);
nand U4076 (N_4076,N_3203,N_2787);
and U4077 (N_4077,N_3132,N_2528);
and U4078 (N_4078,N_3585,N_3280);
xnor U4079 (N_4079,N_3342,N_2751);
nand U4080 (N_4080,N_3008,N_2841);
or U4081 (N_4081,N_2411,N_2469);
nor U4082 (N_4082,N_2552,N_3114);
nor U4083 (N_4083,N_3236,N_2537);
xnor U4084 (N_4084,N_2716,N_3049);
nand U4085 (N_4085,N_3067,N_3368);
nand U4086 (N_4086,N_2791,N_2463);
or U4087 (N_4087,N_2769,N_2625);
or U4088 (N_4088,N_3461,N_3265);
xnor U4089 (N_4089,N_3261,N_3150);
and U4090 (N_4090,N_2968,N_3167);
or U4091 (N_4091,N_3101,N_2708);
nand U4092 (N_4092,N_3196,N_2619);
nor U4093 (N_4093,N_3455,N_3002);
xnor U4094 (N_4094,N_3182,N_2770);
and U4095 (N_4095,N_3263,N_3238);
nand U4096 (N_4096,N_2539,N_3300);
nor U4097 (N_4097,N_2839,N_2628);
nand U4098 (N_4098,N_2522,N_3547);
xnor U4099 (N_4099,N_2876,N_2850);
xor U4100 (N_4100,N_3198,N_2879);
or U4101 (N_4101,N_3267,N_3266);
and U4102 (N_4102,N_3024,N_3056);
nor U4103 (N_4103,N_3578,N_2417);
or U4104 (N_4104,N_3210,N_3176);
nand U4105 (N_4105,N_2689,N_2637);
nor U4106 (N_4106,N_3440,N_3070);
and U4107 (N_4107,N_2459,N_3192);
and U4108 (N_4108,N_2906,N_2852);
nor U4109 (N_4109,N_3445,N_2735);
or U4110 (N_4110,N_3306,N_2517);
nor U4111 (N_4111,N_2727,N_2755);
nand U4112 (N_4112,N_2722,N_2920);
nor U4113 (N_4113,N_2530,N_2785);
and U4114 (N_4114,N_3055,N_2474);
and U4115 (N_4115,N_3046,N_2526);
nand U4116 (N_4116,N_3345,N_2911);
and U4117 (N_4117,N_3558,N_2429);
or U4118 (N_4118,N_3350,N_2825);
nand U4119 (N_4119,N_3596,N_3529);
nand U4120 (N_4120,N_2796,N_2541);
xor U4121 (N_4121,N_2943,N_2857);
nand U4122 (N_4122,N_3292,N_2616);
or U4123 (N_4123,N_2536,N_3520);
nor U4124 (N_4124,N_2610,N_2842);
or U4125 (N_4125,N_2430,N_2941);
nor U4126 (N_4126,N_2963,N_2532);
nor U4127 (N_4127,N_2671,N_3107);
or U4128 (N_4128,N_3528,N_3435);
or U4129 (N_4129,N_3586,N_2926);
and U4130 (N_4130,N_2898,N_3162);
and U4131 (N_4131,N_2680,N_3474);
or U4132 (N_4132,N_2715,N_2808);
nand U4133 (N_4133,N_2772,N_2836);
nand U4134 (N_4134,N_3138,N_2797);
nand U4135 (N_4135,N_2988,N_3511);
nor U4136 (N_4136,N_2401,N_3491);
or U4137 (N_4137,N_2512,N_2881);
nand U4138 (N_4138,N_3185,N_3413);
or U4139 (N_4139,N_2957,N_3513);
or U4140 (N_4140,N_3112,N_2713);
nand U4141 (N_4141,N_3103,N_3539);
nand U4142 (N_4142,N_3534,N_3348);
nand U4143 (N_4143,N_3224,N_3495);
nand U4144 (N_4144,N_3153,N_2535);
nand U4145 (N_4145,N_3115,N_3364);
nor U4146 (N_4146,N_2602,N_3040);
nor U4147 (N_4147,N_2555,N_2465);
nand U4148 (N_4148,N_3022,N_3418);
xor U4149 (N_4149,N_3423,N_3119);
nand U4150 (N_4150,N_3122,N_3430);
and U4151 (N_4151,N_3179,N_3255);
and U4152 (N_4152,N_3341,N_2595);
and U4153 (N_4153,N_2778,N_2977);
and U4154 (N_4154,N_2618,N_3318);
nand U4155 (N_4155,N_2779,N_3420);
nand U4156 (N_4156,N_2752,N_3327);
nor U4157 (N_4157,N_2653,N_2981);
or U4158 (N_4158,N_2697,N_3325);
and U4159 (N_4159,N_3401,N_2567);
nand U4160 (N_4160,N_2832,N_2542);
xnor U4161 (N_4161,N_3548,N_3459);
nand U4162 (N_4162,N_3478,N_3249);
xnor U4163 (N_4163,N_2696,N_2677);
nor U4164 (N_4164,N_3221,N_2887);
nand U4165 (N_4165,N_2407,N_2636);
or U4166 (N_4166,N_2597,N_2711);
and U4167 (N_4167,N_2847,N_3172);
or U4168 (N_4168,N_3335,N_3200);
nor U4169 (N_4169,N_3447,N_3234);
nor U4170 (N_4170,N_2409,N_2426);
and U4171 (N_4171,N_3339,N_2983);
nor U4172 (N_4172,N_2569,N_3465);
xor U4173 (N_4173,N_2995,N_3193);
and U4174 (N_4174,N_3581,N_3050);
nand U4175 (N_4175,N_3125,N_3580);
nand U4176 (N_4176,N_2663,N_2703);
nand U4177 (N_4177,N_3400,N_3139);
nand U4178 (N_4178,N_2936,N_3434);
nor U4179 (N_4179,N_3159,N_2900);
or U4180 (N_4180,N_3559,N_2591);
nand U4181 (N_4181,N_3225,N_2670);
nand U4182 (N_4182,N_3329,N_3000);
nand U4183 (N_4183,N_2721,N_2753);
xnor U4184 (N_4184,N_3437,N_2974);
nand U4185 (N_4185,N_2550,N_3007);
or U4186 (N_4186,N_2559,N_3340);
nand U4187 (N_4187,N_2874,N_2885);
nor U4188 (N_4188,N_3043,N_3189);
or U4189 (N_4189,N_2485,N_2412);
xor U4190 (N_4190,N_3485,N_2912);
or U4191 (N_4191,N_3442,N_2611);
nor U4192 (N_4192,N_2849,N_2884);
nand U4193 (N_4193,N_2585,N_3426);
or U4194 (N_4194,N_2586,N_3080);
xor U4195 (N_4195,N_3336,N_2502);
or U4196 (N_4196,N_3145,N_2448);
nand U4197 (N_4197,N_3550,N_3471);
and U4198 (N_4198,N_3222,N_2468);
nor U4199 (N_4199,N_3205,N_2467);
nand U4200 (N_4200,N_3466,N_2410);
or U4201 (N_4201,N_3443,N_3028);
nor U4202 (N_4202,N_2508,N_3355);
xor U4203 (N_4203,N_2581,N_2667);
nor U4204 (N_4204,N_2654,N_2516);
and U4205 (N_4205,N_3543,N_3359);
nor U4206 (N_4206,N_2615,N_3468);
or U4207 (N_4207,N_3541,N_3288);
xor U4208 (N_4208,N_2808,N_2885);
or U4209 (N_4209,N_3344,N_2566);
nor U4210 (N_4210,N_3316,N_2817);
nand U4211 (N_4211,N_3083,N_3368);
nor U4212 (N_4212,N_3118,N_2554);
nand U4213 (N_4213,N_2771,N_2707);
and U4214 (N_4214,N_3516,N_2878);
nand U4215 (N_4215,N_2923,N_2597);
or U4216 (N_4216,N_3030,N_2948);
nand U4217 (N_4217,N_3439,N_3199);
xnor U4218 (N_4218,N_3391,N_2539);
or U4219 (N_4219,N_2972,N_2413);
nand U4220 (N_4220,N_3221,N_2546);
xor U4221 (N_4221,N_3254,N_3559);
nand U4222 (N_4222,N_3475,N_2799);
nor U4223 (N_4223,N_2700,N_2601);
and U4224 (N_4224,N_2777,N_2572);
or U4225 (N_4225,N_2975,N_2693);
or U4226 (N_4226,N_2640,N_3281);
xor U4227 (N_4227,N_3402,N_2923);
nand U4228 (N_4228,N_3069,N_2906);
nor U4229 (N_4229,N_2828,N_3102);
or U4230 (N_4230,N_2529,N_2749);
or U4231 (N_4231,N_2434,N_3212);
or U4232 (N_4232,N_3003,N_2628);
nor U4233 (N_4233,N_2938,N_3028);
or U4234 (N_4234,N_2761,N_3567);
xnor U4235 (N_4235,N_3134,N_3274);
and U4236 (N_4236,N_3541,N_2660);
and U4237 (N_4237,N_2905,N_2601);
xor U4238 (N_4238,N_2618,N_2620);
nand U4239 (N_4239,N_3048,N_2867);
xor U4240 (N_4240,N_2715,N_3087);
and U4241 (N_4241,N_3057,N_3594);
and U4242 (N_4242,N_2822,N_3341);
xnor U4243 (N_4243,N_2687,N_2995);
nand U4244 (N_4244,N_2611,N_2977);
nor U4245 (N_4245,N_3072,N_2607);
xor U4246 (N_4246,N_2639,N_2627);
and U4247 (N_4247,N_2566,N_2953);
nand U4248 (N_4248,N_3396,N_3446);
xnor U4249 (N_4249,N_2584,N_3395);
nand U4250 (N_4250,N_2952,N_2803);
xor U4251 (N_4251,N_2438,N_3071);
and U4252 (N_4252,N_3394,N_2974);
nor U4253 (N_4253,N_2467,N_2553);
xor U4254 (N_4254,N_3205,N_3311);
xnor U4255 (N_4255,N_3471,N_2637);
xnor U4256 (N_4256,N_2437,N_3077);
nand U4257 (N_4257,N_2727,N_2990);
xor U4258 (N_4258,N_3075,N_2564);
xor U4259 (N_4259,N_2720,N_3119);
nand U4260 (N_4260,N_2578,N_2934);
or U4261 (N_4261,N_2717,N_2475);
and U4262 (N_4262,N_3462,N_3353);
xor U4263 (N_4263,N_2961,N_2606);
xor U4264 (N_4264,N_3485,N_2717);
xnor U4265 (N_4265,N_2583,N_2957);
xnor U4266 (N_4266,N_3426,N_3445);
or U4267 (N_4267,N_3512,N_3024);
and U4268 (N_4268,N_2400,N_2430);
xor U4269 (N_4269,N_3536,N_2869);
nor U4270 (N_4270,N_3179,N_2831);
and U4271 (N_4271,N_2896,N_2626);
xor U4272 (N_4272,N_3297,N_2781);
nand U4273 (N_4273,N_2829,N_3339);
and U4274 (N_4274,N_3376,N_3101);
nor U4275 (N_4275,N_3034,N_2792);
nand U4276 (N_4276,N_3230,N_2787);
xor U4277 (N_4277,N_3204,N_3009);
or U4278 (N_4278,N_2525,N_2655);
nor U4279 (N_4279,N_3256,N_2593);
nand U4280 (N_4280,N_3594,N_2765);
xnor U4281 (N_4281,N_2583,N_3430);
nor U4282 (N_4282,N_3061,N_2750);
xor U4283 (N_4283,N_3397,N_3169);
and U4284 (N_4284,N_3068,N_3317);
nor U4285 (N_4285,N_3082,N_2964);
nor U4286 (N_4286,N_2909,N_3314);
nand U4287 (N_4287,N_3249,N_2428);
and U4288 (N_4288,N_2697,N_3283);
nand U4289 (N_4289,N_3455,N_3512);
or U4290 (N_4290,N_3547,N_3003);
nand U4291 (N_4291,N_3308,N_3403);
nand U4292 (N_4292,N_2896,N_2464);
nand U4293 (N_4293,N_2986,N_2709);
nor U4294 (N_4294,N_2669,N_2606);
and U4295 (N_4295,N_2706,N_2755);
xor U4296 (N_4296,N_3301,N_2763);
and U4297 (N_4297,N_3363,N_2499);
nor U4298 (N_4298,N_3504,N_2830);
xnor U4299 (N_4299,N_2978,N_2700);
or U4300 (N_4300,N_2646,N_2752);
and U4301 (N_4301,N_2526,N_2840);
and U4302 (N_4302,N_2674,N_2759);
nor U4303 (N_4303,N_2712,N_2713);
and U4304 (N_4304,N_2915,N_2669);
nand U4305 (N_4305,N_2408,N_2725);
and U4306 (N_4306,N_3253,N_3451);
and U4307 (N_4307,N_3599,N_3211);
nor U4308 (N_4308,N_3005,N_2717);
and U4309 (N_4309,N_3175,N_2773);
xor U4310 (N_4310,N_2692,N_2781);
or U4311 (N_4311,N_2797,N_3355);
nor U4312 (N_4312,N_2731,N_3526);
xor U4313 (N_4313,N_3568,N_3300);
and U4314 (N_4314,N_2448,N_3010);
nand U4315 (N_4315,N_3532,N_3000);
nor U4316 (N_4316,N_2770,N_2819);
xor U4317 (N_4317,N_2473,N_2436);
nor U4318 (N_4318,N_2641,N_3290);
nand U4319 (N_4319,N_2648,N_2546);
nand U4320 (N_4320,N_3000,N_2610);
or U4321 (N_4321,N_3478,N_2628);
and U4322 (N_4322,N_3241,N_3579);
or U4323 (N_4323,N_3464,N_3540);
xor U4324 (N_4324,N_3074,N_2407);
nand U4325 (N_4325,N_2820,N_3562);
xnor U4326 (N_4326,N_2570,N_2433);
nand U4327 (N_4327,N_3414,N_2987);
xnor U4328 (N_4328,N_2456,N_3005);
nand U4329 (N_4329,N_3215,N_3008);
or U4330 (N_4330,N_3386,N_3161);
xor U4331 (N_4331,N_2414,N_2873);
xor U4332 (N_4332,N_2599,N_3564);
nor U4333 (N_4333,N_2902,N_2791);
xor U4334 (N_4334,N_2657,N_2881);
and U4335 (N_4335,N_2767,N_2610);
nor U4336 (N_4336,N_2901,N_2425);
and U4337 (N_4337,N_3310,N_2968);
nor U4338 (N_4338,N_2559,N_3032);
or U4339 (N_4339,N_2884,N_3591);
nor U4340 (N_4340,N_2429,N_3137);
xor U4341 (N_4341,N_2466,N_2700);
or U4342 (N_4342,N_3069,N_3112);
nand U4343 (N_4343,N_2885,N_3596);
xnor U4344 (N_4344,N_3265,N_2497);
nand U4345 (N_4345,N_3267,N_2917);
or U4346 (N_4346,N_2645,N_3382);
nor U4347 (N_4347,N_3534,N_3017);
or U4348 (N_4348,N_3357,N_2920);
or U4349 (N_4349,N_2536,N_2737);
nand U4350 (N_4350,N_2676,N_2859);
or U4351 (N_4351,N_2856,N_2789);
or U4352 (N_4352,N_3310,N_3349);
xor U4353 (N_4353,N_2581,N_3427);
and U4354 (N_4354,N_3281,N_3237);
or U4355 (N_4355,N_3597,N_2420);
and U4356 (N_4356,N_3441,N_2822);
xor U4357 (N_4357,N_2762,N_2518);
nand U4358 (N_4358,N_3386,N_2941);
or U4359 (N_4359,N_2470,N_3571);
and U4360 (N_4360,N_3529,N_3410);
or U4361 (N_4361,N_3476,N_3251);
xor U4362 (N_4362,N_3382,N_3195);
or U4363 (N_4363,N_2731,N_2468);
and U4364 (N_4364,N_3025,N_3273);
nand U4365 (N_4365,N_3093,N_2815);
and U4366 (N_4366,N_2745,N_3323);
nand U4367 (N_4367,N_2672,N_3255);
nor U4368 (N_4368,N_2437,N_2889);
xor U4369 (N_4369,N_2644,N_2958);
or U4370 (N_4370,N_2846,N_3455);
and U4371 (N_4371,N_2583,N_2892);
nand U4372 (N_4372,N_2921,N_3135);
nor U4373 (N_4373,N_2623,N_2696);
or U4374 (N_4374,N_2734,N_2947);
nor U4375 (N_4375,N_2951,N_3308);
or U4376 (N_4376,N_3357,N_3021);
or U4377 (N_4377,N_2818,N_2973);
or U4378 (N_4378,N_2819,N_3410);
or U4379 (N_4379,N_2896,N_2786);
or U4380 (N_4380,N_2907,N_2453);
xnor U4381 (N_4381,N_3026,N_3212);
or U4382 (N_4382,N_3386,N_2511);
nand U4383 (N_4383,N_2570,N_3050);
or U4384 (N_4384,N_2998,N_2751);
nor U4385 (N_4385,N_3010,N_3284);
or U4386 (N_4386,N_3368,N_2966);
xnor U4387 (N_4387,N_2550,N_2978);
or U4388 (N_4388,N_2401,N_2807);
and U4389 (N_4389,N_3036,N_3542);
nor U4390 (N_4390,N_3015,N_2647);
nand U4391 (N_4391,N_3514,N_2962);
nand U4392 (N_4392,N_2622,N_2922);
nand U4393 (N_4393,N_2815,N_3372);
or U4394 (N_4394,N_3055,N_2494);
and U4395 (N_4395,N_2888,N_2663);
xor U4396 (N_4396,N_2715,N_2800);
or U4397 (N_4397,N_3157,N_2935);
nand U4398 (N_4398,N_2604,N_2745);
and U4399 (N_4399,N_3329,N_2586);
and U4400 (N_4400,N_3541,N_3295);
xor U4401 (N_4401,N_3449,N_2832);
or U4402 (N_4402,N_3298,N_3180);
and U4403 (N_4403,N_2671,N_3399);
xnor U4404 (N_4404,N_3555,N_3317);
and U4405 (N_4405,N_3269,N_3414);
or U4406 (N_4406,N_3335,N_2711);
and U4407 (N_4407,N_3005,N_3427);
or U4408 (N_4408,N_3489,N_2619);
nor U4409 (N_4409,N_2539,N_3047);
nand U4410 (N_4410,N_2934,N_3167);
xnor U4411 (N_4411,N_3292,N_3222);
nand U4412 (N_4412,N_3560,N_3453);
xor U4413 (N_4413,N_2892,N_2503);
or U4414 (N_4414,N_3138,N_2871);
or U4415 (N_4415,N_2752,N_2640);
nand U4416 (N_4416,N_3192,N_2733);
xor U4417 (N_4417,N_2712,N_3263);
or U4418 (N_4418,N_2547,N_2692);
or U4419 (N_4419,N_2486,N_3253);
nor U4420 (N_4420,N_2917,N_2926);
or U4421 (N_4421,N_3436,N_3241);
nand U4422 (N_4422,N_3031,N_3095);
or U4423 (N_4423,N_2860,N_3476);
and U4424 (N_4424,N_3543,N_3457);
nor U4425 (N_4425,N_2923,N_2931);
nor U4426 (N_4426,N_3157,N_3397);
nor U4427 (N_4427,N_3148,N_2541);
nand U4428 (N_4428,N_3567,N_2564);
or U4429 (N_4429,N_2754,N_2702);
and U4430 (N_4430,N_2754,N_2871);
and U4431 (N_4431,N_3257,N_3391);
or U4432 (N_4432,N_3285,N_2552);
nor U4433 (N_4433,N_3567,N_3450);
xnor U4434 (N_4434,N_3099,N_2429);
and U4435 (N_4435,N_3122,N_2434);
and U4436 (N_4436,N_2557,N_3330);
and U4437 (N_4437,N_2557,N_3422);
or U4438 (N_4438,N_3581,N_3152);
xor U4439 (N_4439,N_3032,N_3049);
and U4440 (N_4440,N_2649,N_3275);
or U4441 (N_4441,N_2888,N_2902);
and U4442 (N_4442,N_2611,N_3413);
nand U4443 (N_4443,N_2742,N_3411);
nor U4444 (N_4444,N_3024,N_2640);
xnor U4445 (N_4445,N_3178,N_3427);
or U4446 (N_4446,N_2498,N_2757);
xnor U4447 (N_4447,N_3467,N_2761);
and U4448 (N_4448,N_2404,N_3113);
xnor U4449 (N_4449,N_2533,N_2853);
nand U4450 (N_4450,N_2770,N_3115);
nor U4451 (N_4451,N_3108,N_2856);
nand U4452 (N_4452,N_3372,N_3143);
and U4453 (N_4453,N_3479,N_2921);
nor U4454 (N_4454,N_2915,N_2476);
xor U4455 (N_4455,N_2606,N_2492);
nand U4456 (N_4456,N_3572,N_3524);
nor U4457 (N_4457,N_3597,N_3401);
nor U4458 (N_4458,N_2594,N_3055);
xor U4459 (N_4459,N_3234,N_2533);
or U4460 (N_4460,N_3108,N_2688);
xor U4461 (N_4461,N_3434,N_3492);
and U4462 (N_4462,N_3534,N_3180);
nand U4463 (N_4463,N_3571,N_2999);
xnor U4464 (N_4464,N_3020,N_3326);
nor U4465 (N_4465,N_3124,N_3549);
nand U4466 (N_4466,N_3142,N_2470);
nand U4467 (N_4467,N_3525,N_3435);
nand U4468 (N_4468,N_3257,N_2713);
nor U4469 (N_4469,N_3198,N_2901);
nand U4470 (N_4470,N_2879,N_3537);
nand U4471 (N_4471,N_3220,N_3309);
nand U4472 (N_4472,N_2702,N_2452);
or U4473 (N_4473,N_3573,N_3528);
xnor U4474 (N_4474,N_2553,N_2533);
nor U4475 (N_4475,N_2416,N_2762);
xor U4476 (N_4476,N_3554,N_2802);
nand U4477 (N_4477,N_2490,N_3082);
or U4478 (N_4478,N_3152,N_2658);
and U4479 (N_4479,N_2721,N_3302);
and U4480 (N_4480,N_3312,N_2811);
and U4481 (N_4481,N_3058,N_2565);
xnor U4482 (N_4482,N_2608,N_3396);
or U4483 (N_4483,N_3364,N_3007);
nor U4484 (N_4484,N_3188,N_3478);
nand U4485 (N_4485,N_3220,N_3054);
nor U4486 (N_4486,N_3301,N_2770);
or U4487 (N_4487,N_2439,N_2850);
nand U4488 (N_4488,N_3530,N_3351);
xor U4489 (N_4489,N_2976,N_2401);
xnor U4490 (N_4490,N_3244,N_3003);
nor U4491 (N_4491,N_2646,N_2877);
and U4492 (N_4492,N_3569,N_3048);
xnor U4493 (N_4493,N_3032,N_2762);
nand U4494 (N_4494,N_3023,N_2417);
or U4495 (N_4495,N_3072,N_2487);
nor U4496 (N_4496,N_2927,N_2414);
xor U4497 (N_4497,N_2596,N_2691);
nand U4498 (N_4498,N_2883,N_2768);
nor U4499 (N_4499,N_3170,N_3127);
nor U4500 (N_4500,N_3549,N_3151);
nor U4501 (N_4501,N_3170,N_2538);
nor U4502 (N_4502,N_3215,N_3366);
and U4503 (N_4503,N_3313,N_2824);
and U4504 (N_4504,N_3287,N_2525);
nand U4505 (N_4505,N_3513,N_3571);
and U4506 (N_4506,N_3191,N_3227);
nand U4507 (N_4507,N_3005,N_2454);
and U4508 (N_4508,N_2876,N_2450);
and U4509 (N_4509,N_2554,N_2607);
or U4510 (N_4510,N_2976,N_3055);
and U4511 (N_4511,N_3484,N_2675);
and U4512 (N_4512,N_3267,N_3169);
nor U4513 (N_4513,N_3508,N_2457);
and U4514 (N_4514,N_2981,N_3120);
xor U4515 (N_4515,N_3119,N_2658);
nor U4516 (N_4516,N_2442,N_2902);
and U4517 (N_4517,N_3142,N_3157);
xor U4518 (N_4518,N_2429,N_2968);
nand U4519 (N_4519,N_2679,N_3246);
and U4520 (N_4520,N_2590,N_3380);
nand U4521 (N_4521,N_3016,N_2581);
xnor U4522 (N_4522,N_2431,N_3486);
xnor U4523 (N_4523,N_3158,N_2653);
nand U4524 (N_4524,N_2895,N_2603);
or U4525 (N_4525,N_3562,N_3586);
and U4526 (N_4526,N_2973,N_3198);
nand U4527 (N_4527,N_2706,N_2416);
or U4528 (N_4528,N_3406,N_3494);
xor U4529 (N_4529,N_2475,N_2897);
and U4530 (N_4530,N_3361,N_3271);
and U4531 (N_4531,N_2646,N_2694);
nand U4532 (N_4532,N_3315,N_3019);
xor U4533 (N_4533,N_2457,N_2661);
or U4534 (N_4534,N_2631,N_3441);
nand U4535 (N_4535,N_2591,N_2479);
and U4536 (N_4536,N_2972,N_3105);
nand U4537 (N_4537,N_3110,N_2727);
nand U4538 (N_4538,N_2426,N_3371);
or U4539 (N_4539,N_3284,N_2456);
nand U4540 (N_4540,N_2680,N_2843);
or U4541 (N_4541,N_3203,N_2641);
nand U4542 (N_4542,N_2698,N_3533);
nand U4543 (N_4543,N_3103,N_2941);
or U4544 (N_4544,N_2579,N_3142);
xor U4545 (N_4545,N_2984,N_3354);
or U4546 (N_4546,N_2841,N_3230);
nand U4547 (N_4547,N_2740,N_2694);
or U4548 (N_4548,N_2412,N_2583);
nor U4549 (N_4549,N_2872,N_2977);
nand U4550 (N_4550,N_2843,N_2998);
or U4551 (N_4551,N_2883,N_3063);
or U4552 (N_4552,N_2427,N_2433);
and U4553 (N_4553,N_3167,N_3042);
nor U4554 (N_4554,N_3013,N_2792);
nor U4555 (N_4555,N_3120,N_2546);
nor U4556 (N_4556,N_3561,N_3047);
xor U4557 (N_4557,N_2535,N_3267);
and U4558 (N_4558,N_2595,N_3219);
nand U4559 (N_4559,N_3325,N_2631);
and U4560 (N_4560,N_3078,N_3234);
xor U4561 (N_4561,N_3010,N_3428);
and U4562 (N_4562,N_2582,N_3334);
nand U4563 (N_4563,N_3581,N_3373);
and U4564 (N_4564,N_2908,N_2460);
nand U4565 (N_4565,N_3082,N_3501);
and U4566 (N_4566,N_3233,N_2584);
nand U4567 (N_4567,N_2553,N_2441);
and U4568 (N_4568,N_2507,N_3128);
nand U4569 (N_4569,N_2494,N_3548);
nor U4570 (N_4570,N_3598,N_3012);
or U4571 (N_4571,N_3436,N_2453);
xor U4572 (N_4572,N_3191,N_3266);
nand U4573 (N_4573,N_3560,N_3128);
and U4574 (N_4574,N_2428,N_3529);
xor U4575 (N_4575,N_2608,N_2802);
nor U4576 (N_4576,N_2440,N_3317);
and U4577 (N_4577,N_3408,N_3558);
or U4578 (N_4578,N_3490,N_3199);
or U4579 (N_4579,N_2651,N_2786);
nand U4580 (N_4580,N_3298,N_3166);
or U4581 (N_4581,N_3146,N_2757);
and U4582 (N_4582,N_3573,N_2850);
xor U4583 (N_4583,N_2663,N_2746);
or U4584 (N_4584,N_3489,N_3267);
or U4585 (N_4585,N_2831,N_2978);
or U4586 (N_4586,N_3581,N_2951);
nor U4587 (N_4587,N_2885,N_3262);
or U4588 (N_4588,N_2860,N_3031);
nor U4589 (N_4589,N_2981,N_2788);
nor U4590 (N_4590,N_3520,N_3175);
and U4591 (N_4591,N_3571,N_3483);
or U4592 (N_4592,N_3159,N_3152);
nor U4593 (N_4593,N_2599,N_3446);
nand U4594 (N_4594,N_3326,N_2893);
nor U4595 (N_4595,N_2928,N_2805);
nor U4596 (N_4596,N_3482,N_2948);
nor U4597 (N_4597,N_3264,N_3270);
xnor U4598 (N_4598,N_3305,N_3078);
xor U4599 (N_4599,N_2569,N_2736);
nor U4600 (N_4600,N_2647,N_3200);
or U4601 (N_4601,N_2907,N_3478);
or U4602 (N_4602,N_2773,N_3122);
nand U4603 (N_4603,N_3458,N_3010);
nand U4604 (N_4604,N_2583,N_3053);
nor U4605 (N_4605,N_2590,N_2638);
or U4606 (N_4606,N_3474,N_3491);
or U4607 (N_4607,N_2571,N_2937);
nor U4608 (N_4608,N_2522,N_3100);
xnor U4609 (N_4609,N_2810,N_3066);
nor U4610 (N_4610,N_2609,N_3118);
and U4611 (N_4611,N_3598,N_3221);
or U4612 (N_4612,N_2464,N_3184);
nand U4613 (N_4613,N_2751,N_3077);
nor U4614 (N_4614,N_2790,N_3228);
and U4615 (N_4615,N_3100,N_2884);
xnor U4616 (N_4616,N_3426,N_3019);
nor U4617 (N_4617,N_3380,N_2752);
xnor U4618 (N_4618,N_2525,N_3517);
nor U4619 (N_4619,N_2936,N_2480);
nand U4620 (N_4620,N_3574,N_2598);
or U4621 (N_4621,N_3456,N_2961);
xor U4622 (N_4622,N_2864,N_2568);
nor U4623 (N_4623,N_3354,N_3127);
nor U4624 (N_4624,N_2832,N_3205);
nor U4625 (N_4625,N_2645,N_3431);
nor U4626 (N_4626,N_2732,N_3063);
xor U4627 (N_4627,N_3365,N_3036);
and U4628 (N_4628,N_3578,N_3090);
xor U4629 (N_4629,N_3307,N_2522);
nor U4630 (N_4630,N_3113,N_3170);
nor U4631 (N_4631,N_3598,N_3074);
nor U4632 (N_4632,N_2657,N_2693);
xnor U4633 (N_4633,N_2482,N_3559);
nand U4634 (N_4634,N_2545,N_3411);
nor U4635 (N_4635,N_3004,N_3039);
or U4636 (N_4636,N_3047,N_2588);
and U4637 (N_4637,N_2701,N_2877);
or U4638 (N_4638,N_2570,N_3094);
nor U4639 (N_4639,N_2417,N_2527);
nor U4640 (N_4640,N_2789,N_3498);
nand U4641 (N_4641,N_2796,N_2631);
nor U4642 (N_4642,N_2991,N_2904);
and U4643 (N_4643,N_2697,N_2733);
or U4644 (N_4644,N_3452,N_3083);
and U4645 (N_4645,N_2850,N_3131);
nor U4646 (N_4646,N_3599,N_2666);
xor U4647 (N_4647,N_3324,N_2833);
xor U4648 (N_4648,N_2805,N_2839);
xor U4649 (N_4649,N_2440,N_2906);
or U4650 (N_4650,N_3073,N_2893);
and U4651 (N_4651,N_2544,N_2505);
or U4652 (N_4652,N_2415,N_2489);
or U4653 (N_4653,N_2451,N_3478);
nand U4654 (N_4654,N_2666,N_2400);
nand U4655 (N_4655,N_2482,N_3123);
nand U4656 (N_4656,N_3522,N_2911);
or U4657 (N_4657,N_2402,N_2938);
nor U4658 (N_4658,N_2933,N_2567);
or U4659 (N_4659,N_3298,N_2505);
or U4660 (N_4660,N_3400,N_3010);
or U4661 (N_4661,N_2830,N_3116);
and U4662 (N_4662,N_3490,N_2695);
nor U4663 (N_4663,N_2574,N_3149);
nand U4664 (N_4664,N_2449,N_2579);
nor U4665 (N_4665,N_2617,N_3243);
or U4666 (N_4666,N_2793,N_3508);
nand U4667 (N_4667,N_2429,N_3516);
or U4668 (N_4668,N_2945,N_3515);
or U4669 (N_4669,N_3506,N_3323);
xor U4670 (N_4670,N_2884,N_2811);
nand U4671 (N_4671,N_3415,N_3211);
nor U4672 (N_4672,N_3436,N_3268);
and U4673 (N_4673,N_2433,N_3001);
xnor U4674 (N_4674,N_2643,N_3598);
xnor U4675 (N_4675,N_3047,N_3212);
or U4676 (N_4676,N_3041,N_3255);
and U4677 (N_4677,N_3145,N_2836);
or U4678 (N_4678,N_3446,N_3076);
or U4679 (N_4679,N_2798,N_3245);
or U4680 (N_4680,N_3236,N_2568);
or U4681 (N_4681,N_3141,N_3230);
or U4682 (N_4682,N_2919,N_2724);
nand U4683 (N_4683,N_2418,N_3138);
xnor U4684 (N_4684,N_3555,N_2450);
xnor U4685 (N_4685,N_2744,N_2654);
xnor U4686 (N_4686,N_3222,N_3235);
and U4687 (N_4687,N_2743,N_2727);
and U4688 (N_4688,N_3111,N_3286);
and U4689 (N_4689,N_3106,N_3166);
and U4690 (N_4690,N_3142,N_3276);
nor U4691 (N_4691,N_3563,N_3045);
xor U4692 (N_4692,N_2542,N_3471);
nand U4693 (N_4693,N_3540,N_3243);
or U4694 (N_4694,N_2953,N_2845);
and U4695 (N_4695,N_2705,N_3095);
or U4696 (N_4696,N_2909,N_3213);
nor U4697 (N_4697,N_2885,N_2469);
xor U4698 (N_4698,N_2503,N_3181);
xor U4699 (N_4699,N_3550,N_2969);
and U4700 (N_4700,N_2567,N_3352);
nor U4701 (N_4701,N_3442,N_3203);
and U4702 (N_4702,N_2607,N_2581);
nor U4703 (N_4703,N_3498,N_3222);
or U4704 (N_4704,N_2919,N_3013);
nand U4705 (N_4705,N_3409,N_3385);
or U4706 (N_4706,N_3521,N_3165);
and U4707 (N_4707,N_3134,N_2675);
nand U4708 (N_4708,N_2791,N_3244);
nor U4709 (N_4709,N_2874,N_2681);
and U4710 (N_4710,N_3183,N_2830);
nor U4711 (N_4711,N_3591,N_2619);
or U4712 (N_4712,N_2590,N_2828);
or U4713 (N_4713,N_3033,N_2631);
nand U4714 (N_4714,N_2786,N_2479);
or U4715 (N_4715,N_2695,N_3147);
nor U4716 (N_4716,N_2418,N_2689);
nor U4717 (N_4717,N_3029,N_3587);
or U4718 (N_4718,N_2938,N_2929);
xor U4719 (N_4719,N_3459,N_2852);
and U4720 (N_4720,N_3352,N_3334);
nor U4721 (N_4721,N_3286,N_2671);
or U4722 (N_4722,N_3226,N_3140);
nor U4723 (N_4723,N_3003,N_2778);
nand U4724 (N_4724,N_3113,N_3385);
and U4725 (N_4725,N_3060,N_2873);
or U4726 (N_4726,N_3066,N_2687);
or U4727 (N_4727,N_3582,N_2615);
or U4728 (N_4728,N_3223,N_2767);
nand U4729 (N_4729,N_2776,N_2807);
nor U4730 (N_4730,N_2847,N_2898);
xor U4731 (N_4731,N_2732,N_2650);
nor U4732 (N_4732,N_3167,N_2961);
xnor U4733 (N_4733,N_3387,N_3260);
nand U4734 (N_4734,N_2736,N_2877);
xnor U4735 (N_4735,N_2937,N_3444);
or U4736 (N_4736,N_2463,N_2609);
or U4737 (N_4737,N_3151,N_3389);
or U4738 (N_4738,N_2581,N_2786);
xor U4739 (N_4739,N_2972,N_2649);
xnor U4740 (N_4740,N_2610,N_2886);
or U4741 (N_4741,N_2648,N_2400);
and U4742 (N_4742,N_3435,N_3080);
nor U4743 (N_4743,N_2524,N_2425);
or U4744 (N_4744,N_2540,N_3273);
and U4745 (N_4745,N_3505,N_2806);
nand U4746 (N_4746,N_2750,N_2843);
and U4747 (N_4747,N_3255,N_3325);
nand U4748 (N_4748,N_3235,N_2831);
nor U4749 (N_4749,N_2511,N_2925);
xnor U4750 (N_4750,N_3415,N_3353);
xnor U4751 (N_4751,N_3465,N_3060);
nor U4752 (N_4752,N_2745,N_3531);
nor U4753 (N_4753,N_3431,N_2910);
and U4754 (N_4754,N_3285,N_2655);
xnor U4755 (N_4755,N_2950,N_3367);
xnor U4756 (N_4756,N_2528,N_2917);
or U4757 (N_4757,N_2841,N_3024);
nand U4758 (N_4758,N_2754,N_2626);
xor U4759 (N_4759,N_3344,N_2761);
nor U4760 (N_4760,N_2530,N_3292);
nor U4761 (N_4761,N_2479,N_2805);
or U4762 (N_4762,N_3396,N_3072);
or U4763 (N_4763,N_2832,N_3451);
xor U4764 (N_4764,N_2594,N_2758);
nor U4765 (N_4765,N_2531,N_3010);
xnor U4766 (N_4766,N_2938,N_2852);
nor U4767 (N_4767,N_3376,N_2527);
nor U4768 (N_4768,N_3188,N_3336);
or U4769 (N_4769,N_2545,N_3566);
and U4770 (N_4770,N_3408,N_2412);
and U4771 (N_4771,N_2501,N_3481);
nor U4772 (N_4772,N_3147,N_2748);
or U4773 (N_4773,N_3541,N_3373);
xnor U4774 (N_4774,N_2579,N_2498);
xnor U4775 (N_4775,N_2583,N_3382);
xnor U4776 (N_4776,N_3212,N_2693);
nor U4777 (N_4777,N_2442,N_2641);
nand U4778 (N_4778,N_3320,N_2528);
and U4779 (N_4779,N_2738,N_3378);
xor U4780 (N_4780,N_3029,N_2472);
and U4781 (N_4781,N_3065,N_3517);
or U4782 (N_4782,N_2556,N_3450);
nor U4783 (N_4783,N_3321,N_2415);
xor U4784 (N_4784,N_2479,N_3574);
xnor U4785 (N_4785,N_3203,N_3574);
nand U4786 (N_4786,N_3223,N_3137);
or U4787 (N_4787,N_2721,N_2728);
nand U4788 (N_4788,N_3564,N_2840);
xnor U4789 (N_4789,N_2980,N_2931);
nor U4790 (N_4790,N_3429,N_2513);
or U4791 (N_4791,N_3454,N_3583);
nand U4792 (N_4792,N_2933,N_3193);
xor U4793 (N_4793,N_3475,N_3092);
xnor U4794 (N_4794,N_3164,N_2482);
nor U4795 (N_4795,N_3009,N_2941);
xnor U4796 (N_4796,N_2761,N_2537);
nor U4797 (N_4797,N_2463,N_2789);
nand U4798 (N_4798,N_3253,N_2883);
xnor U4799 (N_4799,N_3566,N_2473);
nand U4800 (N_4800,N_3858,N_4439);
nand U4801 (N_4801,N_4553,N_4698);
xor U4802 (N_4802,N_4373,N_4455);
or U4803 (N_4803,N_4481,N_4342);
xnor U4804 (N_4804,N_4382,N_3674);
or U4805 (N_4805,N_4551,N_4337);
and U4806 (N_4806,N_4119,N_3912);
and U4807 (N_4807,N_4503,N_4179);
nor U4808 (N_4808,N_4605,N_4304);
xor U4809 (N_4809,N_4130,N_4302);
nand U4810 (N_4810,N_4197,N_4482);
and U4811 (N_4811,N_4762,N_4193);
xnor U4812 (N_4812,N_4157,N_4068);
and U4813 (N_4813,N_3751,N_4377);
nand U4814 (N_4814,N_4617,N_4225);
and U4815 (N_4815,N_4165,N_4160);
nand U4816 (N_4816,N_4451,N_4094);
and U4817 (N_4817,N_4779,N_4743);
xor U4818 (N_4818,N_3722,N_3744);
or U4819 (N_4819,N_4100,N_4274);
or U4820 (N_4820,N_4109,N_3915);
nand U4821 (N_4821,N_3843,N_3705);
xor U4822 (N_4822,N_3974,N_4674);
xnor U4823 (N_4823,N_4376,N_4404);
xor U4824 (N_4824,N_4453,N_3787);
or U4825 (N_4825,N_4209,N_3738);
nor U4826 (N_4826,N_4387,N_4391);
and U4827 (N_4827,N_4520,N_4671);
nand U4828 (N_4828,N_4266,N_4516);
xor U4829 (N_4829,N_3792,N_4026);
and U4830 (N_4830,N_3921,N_3856);
nor U4831 (N_4831,N_4147,N_4688);
nand U4832 (N_4832,N_3965,N_3621);
or U4833 (N_4833,N_4349,N_3770);
or U4834 (N_4834,N_4704,N_4000);
or U4835 (N_4835,N_3944,N_4564);
or U4836 (N_4836,N_4500,N_3958);
nand U4837 (N_4837,N_4378,N_4465);
and U4838 (N_4838,N_4610,N_4246);
nor U4839 (N_4839,N_3716,N_3654);
nand U4840 (N_4840,N_4150,N_3760);
nor U4841 (N_4841,N_4466,N_4051);
or U4842 (N_4842,N_4033,N_4399);
and U4843 (N_4843,N_4129,N_4265);
xor U4844 (N_4844,N_3901,N_4393);
or U4845 (N_4845,N_4189,N_4488);
nand U4846 (N_4846,N_3872,N_4400);
xnor U4847 (N_4847,N_4372,N_4662);
and U4848 (N_4848,N_4788,N_3839);
nand U4849 (N_4849,N_4708,N_3933);
nand U4850 (N_4850,N_4449,N_4594);
nor U4851 (N_4851,N_4028,N_3752);
nor U4852 (N_4852,N_4543,N_3956);
and U4853 (N_4853,N_3694,N_3859);
xnor U4854 (N_4854,N_4243,N_4355);
and U4855 (N_4855,N_3922,N_3880);
nor U4856 (N_4856,N_4043,N_4116);
xor U4857 (N_4857,N_4559,N_4340);
or U4858 (N_4858,N_3885,N_3703);
nor U4859 (N_4859,N_3689,N_4050);
xor U4860 (N_4860,N_3765,N_4023);
xor U4861 (N_4861,N_4227,N_3690);
or U4862 (N_4862,N_4663,N_3785);
nand U4863 (N_4863,N_4714,N_3747);
or U4864 (N_4864,N_3647,N_4418);
xor U4865 (N_4865,N_4600,N_3819);
nor U4866 (N_4866,N_4240,N_3896);
or U4867 (N_4867,N_4245,N_3851);
and U4868 (N_4868,N_3935,N_4398);
nor U4869 (N_4869,N_4421,N_4767);
nor U4870 (N_4870,N_4134,N_4030);
nor U4871 (N_4871,N_4271,N_4595);
or U4872 (N_4872,N_4303,N_4352);
xor U4873 (N_4873,N_3619,N_4408);
or U4874 (N_4874,N_4626,N_4327);
xnor U4875 (N_4875,N_3946,N_3725);
or U4876 (N_4876,N_4707,N_4711);
or U4877 (N_4877,N_4506,N_3838);
and U4878 (N_4878,N_4095,N_4347);
xor U4879 (N_4879,N_4277,N_4394);
xnor U4880 (N_4880,N_4385,N_3848);
nand U4881 (N_4881,N_4734,N_4728);
and U4882 (N_4882,N_3604,N_4690);
and U4883 (N_4883,N_4363,N_3772);
nand U4884 (N_4884,N_4141,N_4320);
or U4885 (N_4885,N_4776,N_3650);
and U4886 (N_4886,N_4736,N_4383);
or U4887 (N_4887,N_4729,N_4463);
xor U4888 (N_4888,N_3952,N_4461);
and U4889 (N_4889,N_4508,N_3937);
nor U4890 (N_4890,N_3841,N_3957);
and U4891 (N_4891,N_4745,N_4735);
or U4892 (N_4892,N_3825,N_3989);
nor U4893 (N_4893,N_3750,N_4331);
and U4894 (N_4894,N_4174,N_4066);
xor U4895 (N_4895,N_4003,N_4231);
nor U4896 (N_4896,N_4200,N_4081);
or U4897 (N_4897,N_3749,N_3671);
nor U4898 (N_4898,N_3633,N_4162);
nor U4899 (N_4899,N_4298,N_3798);
xor U4900 (N_4900,N_4625,N_4341);
and U4901 (N_4901,N_3846,N_4317);
xor U4902 (N_4902,N_4115,N_4038);
and U4903 (N_4903,N_4470,N_4550);
or U4904 (N_4904,N_3834,N_4422);
or U4905 (N_4905,N_3620,N_3913);
nor U4906 (N_4906,N_3822,N_3774);
xnor U4907 (N_4907,N_3823,N_4701);
nor U4908 (N_4908,N_4517,N_3998);
and U4909 (N_4909,N_3876,N_4702);
nand U4910 (N_4910,N_4353,N_4732);
or U4911 (N_4911,N_4281,N_4042);
and U4912 (N_4912,N_4526,N_3763);
nand U4913 (N_4913,N_4326,N_3803);
xor U4914 (N_4914,N_4673,N_3666);
nand U4915 (N_4915,N_4612,N_3636);
xnor U4916 (N_4916,N_4345,N_4253);
nand U4917 (N_4917,N_4211,N_4187);
xor U4918 (N_4918,N_4096,N_3977);
and U4919 (N_4919,N_4754,N_4417);
or U4920 (N_4920,N_3693,N_4343);
nand U4921 (N_4921,N_3735,N_4135);
nor U4922 (N_4922,N_4017,N_4318);
nand U4923 (N_4923,N_4772,N_4644);
xnor U4924 (N_4924,N_3649,N_3610);
nor U4925 (N_4925,N_4660,N_3826);
nor U4926 (N_4926,N_4228,N_4777);
and U4927 (N_4927,N_4218,N_4713);
nand U4928 (N_4928,N_4206,N_4339);
nand U4929 (N_4929,N_4446,N_3852);
xnor U4930 (N_4930,N_4616,N_4560);
nor U4931 (N_4931,N_4098,N_3854);
or U4932 (N_4932,N_4155,N_4739);
and U4933 (N_4933,N_4783,N_3925);
nand U4934 (N_4934,N_4726,N_4367);
xor U4935 (N_4935,N_4636,N_3987);
and U4936 (N_4936,N_3831,N_3845);
nand U4937 (N_4937,N_4024,N_3991);
nand U4938 (N_4938,N_4618,N_4272);
nor U4939 (N_4939,N_3714,N_4438);
nor U4940 (N_4940,N_3948,N_4267);
or U4941 (N_4941,N_4061,N_4537);
nand U4942 (N_4942,N_3736,N_4715);
and U4943 (N_4943,N_4556,N_3753);
nand U4944 (N_4944,N_4678,N_4686);
and U4945 (N_4945,N_4493,N_4679);
and U4946 (N_4946,N_4477,N_3691);
xnor U4947 (N_4947,N_4368,N_4709);
nor U4948 (N_4948,N_4668,N_4501);
nor U4949 (N_4949,N_3655,N_4593);
and U4950 (N_4950,N_4216,N_4031);
nand U4951 (N_4951,N_4259,N_3951);
nor U4952 (N_4952,N_4585,N_4138);
nor U4953 (N_4953,N_3985,N_4260);
xnor U4954 (N_4954,N_3833,N_4648);
xor U4955 (N_4955,N_4603,N_3943);
nor U4956 (N_4956,N_3615,N_3969);
nor U4957 (N_4957,N_4101,N_4442);
and U4958 (N_4958,N_3942,N_4620);
or U4959 (N_4959,N_4299,N_3962);
and U4960 (N_4960,N_4167,N_4676);
nor U4961 (N_4961,N_4143,N_4787);
nor U4962 (N_4962,N_3889,N_3869);
and U4963 (N_4963,N_3993,N_4044);
xnor U4964 (N_4964,N_3603,N_4108);
xor U4965 (N_4965,N_4063,N_4490);
and U4966 (N_4966,N_3642,N_4006);
nand U4967 (N_4967,N_4464,N_4164);
xnor U4968 (N_4968,N_4062,N_4548);
xor U4969 (N_4969,N_4346,N_3618);
or U4970 (N_4970,N_4703,N_4474);
xor U4971 (N_4971,N_3811,N_3908);
and U4972 (N_4972,N_4250,N_4215);
nand U4973 (N_4973,N_3984,N_4622);
nand U4974 (N_4974,N_3609,N_3635);
xnor U4975 (N_4975,N_4639,N_3634);
or U4976 (N_4976,N_4110,N_4624);
and U4977 (N_4977,N_3656,N_3886);
and U4978 (N_4978,N_3664,N_3967);
and U4979 (N_4979,N_4746,N_4191);
nor U4980 (N_4980,N_4531,N_4627);
or U4981 (N_4981,N_3737,N_4074);
nor U4982 (N_4982,N_4512,N_4423);
and U4983 (N_4983,N_4136,N_4573);
xor U4984 (N_4984,N_3730,N_4675);
nand U4985 (N_4985,N_4669,N_3662);
nor U4986 (N_4986,N_4224,N_3806);
or U4987 (N_4987,N_4547,N_4275);
xnor U4988 (N_4988,N_4381,N_3623);
or U4989 (N_4989,N_3867,N_4263);
xnor U4990 (N_4990,N_3931,N_4397);
nor U4991 (N_4991,N_4070,N_3874);
and U4992 (N_4992,N_4236,N_3924);
nor U4993 (N_4993,N_4757,N_3676);
and U4994 (N_4994,N_3805,N_4264);
and U4995 (N_4995,N_4780,N_4609);
xor U4996 (N_4996,N_3727,N_3849);
or U4997 (N_4997,N_3732,N_3776);
or U4998 (N_4998,N_3812,N_4571);
nand U4999 (N_4999,N_3853,N_3726);
nand U5000 (N_5000,N_4518,N_3653);
nor U5001 (N_5001,N_4276,N_4117);
or U5002 (N_5002,N_4409,N_4049);
and U5003 (N_5003,N_4297,N_3778);
nor U5004 (N_5004,N_4196,N_4120);
or U5005 (N_5005,N_3679,N_4007);
and U5006 (N_5006,N_4720,N_3626);
xnor U5007 (N_5007,N_4557,N_4034);
nor U5008 (N_5008,N_4410,N_4795);
nand U5009 (N_5009,N_4414,N_4572);
and U5010 (N_5010,N_4311,N_3746);
nand U5011 (N_5011,N_4080,N_4148);
or U5012 (N_5012,N_4005,N_4581);
nor U5013 (N_5013,N_4667,N_4306);
nand U5014 (N_5014,N_4613,N_3923);
and U5015 (N_5015,N_3608,N_4507);
and U5016 (N_5016,N_4380,N_4471);
xnor U5017 (N_5017,N_4085,N_3895);
nand U5018 (N_5018,N_3968,N_4717);
nor U5019 (N_5019,N_4476,N_4468);
and U5020 (N_5020,N_4473,N_3761);
nor U5021 (N_5021,N_4226,N_4203);
or U5022 (N_5022,N_3651,N_3938);
xnor U5023 (N_5023,N_3961,N_4601);
nand U5024 (N_5024,N_3959,N_4020);
xnor U5025 (N_5025,N_4151,N_4219);
or U5026 (N_5026,N_4480,N_3978);
or U5027 (N_5027,N_4533,N_4322);
nand U5028 (N_5028,N_4121,N_4775);
and U5029 (N_5029,N_4527,N_4596);
and U5030 (N_5030,N_3904,N_4048);
xor U5031 (N_5031,N_4666,N_4727);
nand U5032 (N_5032,N_3818,N_4694);
xnor U5033 (N_5033,N_4047,N_3794);
and U5034 (N_5034,N_3971,N_3791);
nand U5035 (N_5035,N_4587,N_3729);
nor U5036 (N_5036,N_3641,N_4770);
or U5037 (N_5037,N_4640,N_4021);
or U5038 (N_5038,N_4213,N_4152);
or U5039 (N_5039,N_3638,N_4499);
nand U5040 (N_5040,N_3769,N_4032);
or U5041 (N_5041,N_4172,N_4205);
xnor U5042 (N_5042,N_4334,N_4107);
xnor U5043 (N_5043,N_4724,N_3683);
nor U5044 (N_5044,N_4035,N_4190);
nand U5045 (N_5045,N_3809,N_4638);
and U5046 (N_5046,N_3710,N_3780);
and U5047 (N_5047,N_3646,N_3622);
nand U5048 (N_5048,N_4362,N_3930);
or U5049 (N_5049,N_4126,N_4697);
nor U5050 (N_5050,N_3926,N_3865);
and U5051 (N_5051,N_4577,N_4356);
or U5052 (N_5052,N_4255,N_4554);
nor U5053 (N_5053,N_4008,N_4123);
or U5054 (N_5054,N_3972,N_4186);
xor U5055 (N_5055,N_3900,N_4221);
nand U5056 (N_5056,N_4037,N_4099);
and U5057 (N_5057,N_4544,N_4329);
nor U5058 (N_5058,N_4045,N_3884);
nor U5059 (N_5059,N_4183,N_3600);
xor U5060 (N_5060,N_4722,N_3860);
xor U5061 (N_5061,N_4436,N_4432);
or U5062 (N_5062,N_3907,N_3652);
nor U5063 (N_5063,N_3684,N_4539);
nor U5064 (N_5064,N_4350,N_4784);
nor U5065 (N_5065,N_4307,N_4296);
or U5066 (N_5066,N_4723,N_4124);
nor U5067 (N_5067,N_4525,N_4153);
and U5068 (N_5068,N_4486,N_4693);
nand U5069 (N_5069,N_3829,N_4106);
nor U5070 (N_5070,N_3940,N_4046);
or U5071 (N_5071,N_4791,N_4628);
nor U5072 (N_5072,N_3768,N_4055);
nor U5073 (N_5073,N_4405,N_4357);
nand U5074 (N_5074,N_3767,N_4485);
xor U5075 (N_5075,N_3741,N_4194);
xnor U5076 (N_5076,N_4336,N_4755);
xor U5077 (N_5077,N_3709,N_4498);
or U5078 (N_5078,N_4684,N_3918);
or U5079 (N_5079,N_3892,N_4168);
nor U5080 (N_5080,N_3932,N_4472);
nor U5081 (N_5081,N_4606,N_3832);
and U5082 (N_5082,N_3677,N_4672);
and U5083 (N_5083,N_4567,N_3947);
or U5084 (N_5084,N_4721,N_3973);
nand U5085 (N_5085,N_4075,N_4309);
xor U5086 (N_5086,N_3706,N_4608);
nand U5087 (N_5087,N_3643,N_4237);
or U5088 (N_5088,N_4204,N_4534);
or U5089 (N_5089,N_4575,N_4744);
nand U5090 (N_5090,N_4132,N_4103);
xor U5091 (N_5091,N_4437,N_4576);
and U5092 (N_5092,N_4330,N_4665);
or U5093 (N_5093,N_4786,N_4258);
xnor U5094 (N_5094,N_3715,N_3721);
nand U5095 (N_5095,N_3999,N_4386);
and U5096 (N_5096,N_4725,N_4649);
nor U5097 (N_5097,N_3807,N_3857);
nand U5098 (N_5098,N_4022,N_3866);
nor U5099 (N_5099,N_3740,N_3996);
nor U5100 (N_5100,N_3673,N_3879);
or U5101 (N_5101,N_3963,N_4053);
nor U5102 (N_5102,N_4484,N_4435);
or U5103 (N_5103,N_4333,N_3628);
nand U5104 (N_5104,N_3840,N_4097);
xnor U5105 (N_5105,N_4328,N_4630);
xor U5106 (N_5106,N_3888,N_3745);
nor U5107 (N_5107,N_3612,N_3790);
nand U5108 (N_5108,N_4647,N_4392);
nor U5109 (N_5109,N_4344,N_4450);
nor U5110 (N_5110,N_3797,N_4681);
or U5111 (N_5111,N_4558,N_4521);
xor U5112 (N_5112,N_4419,N_3862);
or U5113 (N_5113,N_3698,N_3617);
nor U5114 (N_5114,N_4467,N_3927);
or U5115 (N_5115,N_4010,N_3708);
and U5116 (N_5116,N_4360,N_3661);
xor U5117 (N_5117,N_4395,N_4538);
nand U5118 (N_5118,N_3775,N_4166);
nor U5119 (N_5119,N_4175,N_3658);
nor U5120 (N_5120,N_4761,N_3827);
nand U5121 (N_5121,N_4092,N_4441);
nand U5122 (N_5122,N_4323,N_4443);
or U5123 (N_5123,N_4156,N_4069);
nor U5124 (N_5124,N_4479,N_4748);
nand U5125 (N_5125,N_4511,N_4768);
or U5126 (N_5126,N_3637,N_3629);
xor U5127 (N_5127,N_3648,N_3875);
nor U5128 (N_5128,N_4712,N_4396);
or U5129 (N_5129,N_4651,N_3868);
or U5130 (N_5130,N_4128,N_4431);
and U5131 (N_5131,N_4753,N_4234);
nand U5132 (N_5132,N_4113,N_4154);
and U5133 (N_5133,N_4615,N_4781);
or U5134 (N_5134,N_3699,N_4661);
and U5135 (N_5135,N_4285,N_4036);
and U5136 (N_5136,N_4492,N_3916);
xor U5137 (N_5137,N_4579,N_4384);
nand U5138 (N_5138,N_3645,N_4737);
nand U5139 (N_5139,N_3981,N_4241);
or U5140 (N_5140,N_4086,N_4532);
xor U5141 (N_5141,N_4652,N_3631);
nand U5142 (N_5142,N_4689,N_3665);
and U5143 (N_5143,N_3669,N_4146);
or U5144 (N_5144,N_4590,N_4161);
or U5145 (N_5145,N_4706,N_3960);
or U5146 (N_5146,N_4426,N_4294);
xnor U5147 (N_5147,N_4140,N_3801);
nand U5148 (N_5148,N_4114,N_4252);
and U5149 (N_5149,N_3607,N_4248);
nor U5150 (N_5150,N_3611,N_4429);
xnor U5151 (N_5151,N_4586,N_3898);
or U5152 (N_5152,N_4562,N_4730);
nor U5153 (N_5153,N_4509,N_3817);
nand U5154 (N_5154,N_4619,N_4176);
and U5155 (N_5155,N_3660,N_4052);
and U5156 (N_5156,N_4778,N_4082);
nand U5157 (N_5157,N_4057,N_4589);
or U5158 (N_5158,N_3863,N_3979);
xnor U5159 (N_5159,N_3894,N_4015);
and U5160 (N_5160,N_3897,N_4188);
xnor U5161 (N_5161,N_4771,N_3687);
xnor U5162 (N_5162,N_3632,N_4522);
nor U5163 (N_5163,N_3864,N_4535);
or U5164 (N_5164,N_4133,N_3835);
and U5165 (N_5165,N_4278,N_4580);
xor U5166 (N_5166,N_4591,N_3704);
or U5167 (N_5167,N_4524,N_4584);
nor U5168 (N_5168,N_3605,N_3670);
nand U5169 (N_5169,N_3847,N_4270);
nand U5170 (N_5170,N_4144,N_4301);
nor U5171 (N_5171,N_4089,N_3992);
or U5172 (N_5172,N_4599,N_3734);
xor U5173 (N_5173,N_3711,N_4653);
nor U5174 (N_5174,N_3887,N_4321);
or U5175 (N_5175,N_4390,N_4561);
nor U5176 (N_5176,N_4290,N_3782);
xnor U5177 (N_5177,N_4705,N_4242);
or U5178 (N_5178,N_4799,N_4181);
xor U5179 (N_5179,N_4621,N_4741);
or U5180 (N_5180,N_4013,N_4529);
and U5181 (N_5181,N_3954,N_4406);
nand U5182 (N_5182,N_4502,N_4632);
and U5183 (N_5183,N_4412,N_3850);
nand U5184 (N_5184,N_4566,N_4454);
or U5185 (N_5185,N_4578,N_4122);
nand U5186 (N_5186,N_3893,N_4401);
xnor U5187 (N_5187,N_4659,N_3828);
nand U5188 (N_5188,N_4180,N_4093);
or U5189 (N_5189,N_4379,N_4459);
nor U5190 (N_5190,N_3675,N_4235);
xor U5191 (N_5191,N_4489,N_4305);
or U5192 (N_5192,N_3905,N_3697);
xnor U5193 (N_5193,N_4084,N_4088);
and U5194 (N_5194,N_3657,N_3804);
xor U5195 (N_5195,N_4232,N_4315);
or U5196 (N_5196,N_3728,N_4288);
or U5197 (N_5197,N_4491,N_3821);
xnor U5198 (N_5198,N_4268,N_3781);
or U5199 (N_5199,N_3983,N_4658);
xor U5200 (N_5200,N_4425,N_4765);
and U5201 (N_5201,N_4677,N_4029);
nand U5202 (N_5202,N_4497,N_4794);
xor U5203 (N_5203,N_3994,N_3627);
and U5204 (N_5204,N_4764,N_4261);
nand U5205 (N_5205,N_4541,N_4588);
and U5206 (N_5206,N_3995,N_4763);
or U5207 (N_5207,N_4067,N_3920);
nor U5208 (N_5208,N_4293,N_3903);
nand U5209 (N_5209,N_4475,N_4760);
xnor U5210 (N_5210,N_4016,N_4254);
nand U5211 (N_5211,N_3997,N_4112);
nor U5212 (N_5212,N_3755,N_3719);
nor U5213 (N_5213,N_4568,N_4249);
and U5214 (N_5214,N_4256,N_4790);
nand U5215 (N_5215,N_4719,N_3601);
or U5216 (N_5216,N_4087,N_4338);
xor U5217 (N_5217,N_4145,N_3795);
or U5218 (N_5218,N_3639,N_4312);
nor U5219 (N_5219,N_4065,N_4319);
nand U5220 (N_5220,N_4583,N_4528);
xnor U5221 (N_5221,N_4054,N_3970);
nand U5222 (N_5222,N_4182,N_4105);
and U5223 (N_5223,N_3739,N_4510);
xor U5224 (N_5224,N_4483,N_4629);
xor U5225 (N_5225,N_4371,N_4078);
xor U5226 (N_5226,N_4230,N_3723);
or U5227 (N_5227,N_4223,N_4462);
xnor U5228 (N_5228,N_3717,N_4504);
nand U5229 (N_5229,N_4286,N_3917);
xnor U5230 (N_5230,N_3982,N_4403);
nor U5231 (N_5231,N_4635,N_3702);
nand U5232 (N_5232,N_4782,N_4604);
or U5233 (N_5233,N_3881,N_4797);
or U5234 (N_5234,N_3659,N_4792);
xnor U5235 (N_5235,N_4375,N_3748);
nor U5236 (N_5236,N_3883,N_3815);
or U5237 (N_5237,N_3799,N_4072);
and U5238 (N_5238,N_4348,N_4798);
nand U5239 (N_5239,N_4494,N_4420);
nor U5240 (N_5240,N_4059,N_4351);
and U5241 (N_5241,N_4633,N_4514);
or U5242 (N_5242,N_4752,N_3796);
xnor U5243 (N_5243,N_3990,N_4262);
or U5244 (N_5244,N_4565,N_3914);
nor U5245 (N_5245,N_4139,N_3733);
and U5246 (N_5246,N_4716,N_4212);
xnor U5247 (N_5247,N_3945,N_3686);
nand U5248 (N_5248,N_4657,N_4738);
and U5249 (N_5249,N_4447,N_3678);
or U5250 (N_5250,N_4416,N_3837);
xor U5251 (N_5251,N_4536,N_4102);
or U5252 (N_5252,N_4424,N_3764);
or U5253 (N_5253,N_4027,N_3939);
xnor U5254 (N_5254,N_3929,N_3890);
nand U5255 (N_5255,N_4592,N_4004);
nand U5256 (N_5256,N_4201,N_4774);
xor U5257 (N_5257,N_4430,N_4118);
or U5258 (N_5258,N_4199,N_4643);
nor U5259 (N_5259,N_4014,N_3616);
or U5260 (N_5260,N_3783,N_4750);
xor U5261 (N_5261,N_4064,N_4407);
and U5262 (N_5262,N_4018,N_4598);
nor U5263 (N_5263,N_4220,N_4040);
or U5264 (N_5264,N_3640,N_4295);
nand U5265 (N_5265,N_4523,N_3682);
nand U5266 (N_5266,N_3724,N_4056);
xnor U5267 (N_5267,N_3680,N_4244);
nor U5268 (N_5268,N_3919,N_4184);
xnor U5269 (N_5269,N_4308,N_4171);
and U5270 (N_5270,N_3758,N_4513);
or U5271 (N_5271,N_4680,N_4041);
nand U5272 (N_5272,N_4279,N_4469);
nand U5273 (N_5273,N_3754,N_3773);
and U5274 (N_5274,N_4170,N_4125);
nor U5275 (N_5275,N_3988,N_3743);
nand U5276 (N_5276,N_3842,N_4354);
nand U5277 (N_5277,N_4793,N_3789);
nor U5278 (N_5278,N_3955,N_4691);
or U5279 (N_5279,N_3800,N_4332);
or U5280 (N_5280,N_4570,N_3802);
nand U5281 (N_5281,N_4433,N_3786);
or U5282 (N_5282,N_4359,N_4602);
and U5283 (N_5283,N_4300,N_3667);
or U5284 (N_5284,N_4198,N_4545);
nand U5285 (N_5285,N_3696,N_3756);
or U5286 (N_5286,N_4325,N_4158);
or U5287 (N_5287,N_4549,N_3891);
or U5288 (N_5288,N_4361,N_4682);
xnor U5289 (N_5289,N_4530,N_3663);
nand U5290 (N_5290,N_4458,N_3814);
nor U5291 (N_5291,N_4460,N_4009);
or U5292 (N_5292,N_4289,N_4519);
nor U5293 (N_5293,N_4335,N_4656);
xnor U5294 (N_5294,N_3855,N_3882);
nor U5295 (N_5295,N_4169,N_4019);
xnor U5296 (N_5296,N_4444,N_4185);
and U5297 (N_5297,N_3784,N_4273);
and U5298 (N_5298,N_3625,N_4369);
nand U5299 (N_5299,N_4239,N_4077);
xor U5300 (N_5300,N_4785,N_4364);
and U5301 (N_5301,N_3810,N_4552);
and U5302 (N_5302,N_4071,N_3613);
or U5303 (N_5303,N_4001,N_4411);
or U5304 (N_5304,N_4413,N_4733);
xnor U5305 (N_5305,N_3788,N_4699);
nor U5306 (N_5306,N_3808,N_3602);
nor U5307 (N_5307,N_4747,N_4083);
nor U5308 (N_5308,N_3976,N_3759);
and U5309 (N_5309,N_3681,N_4457);
or U5310 (N_5310,N_4111,N_4655);
and U5311 (N_5311,N_4751,N_4011);
or U5312 (N_5312,N_4637,N_4104);
nor U5313 (N_5313,N_4440,N_4208);
or U5314 (N_5314,N_3731,N_4058);
or U5315 (N_5315,N_3777,N_4796);
or U5316 (N_5316,N_4607,N_4456);
or U5317 (N_5317,N_4773,N_3707);
or U5318 (N_5318,N_4149,N_4076);
nand U5319 (N_5319,N_4641,N_4324);
nor U5320 (N_5320,N_4445,N_4310);
or U5321 (N_5321,N_3910,N_4291);
xnor U5322 (N_5322,N_4611,N_3861);
nand U5323 (N_5323,N_3830,N_3975);
and U5324 (N_5324,N_3824,N_4683);
or U5325 (N_5325,N_3949,N_4687);
and U5326 (N_5326,N_3986,N_4448);
xnor U5327 (N_5327,N_3964,N_3873);
xor U5328 (N_5328,N_4654,N_4495);
and U5329 (N_5329,N_4238,N_4650);
nor U5330 (N_5330,N_3701,N_3757);
nor U5331 (N_5331,N_3771,N_3630);
xor U5332 (N_5332,N_3685,N_3624);
or U5333 (N_5333,N_4284,N_4428);
xor U5334 (N_5334,N_4374,N_3793);
nor U5335 (N_5335,N_4251,N_4269);
nor U5336 (N_5336,N_4137,N_3668);
nor U5337 (N_5337,N_4173,N_4766);
nor U5338 (N_5338,N_3688,N_3934);
nand U5339 (N_5339,N_4389,N_3779);
nand U5340 (N_5340,N_3928,N_3902);
xor U5341 (N_5341,N_4692,N_4233);
nor U5342 (N_5342,N_4487,N_4670);
or U5343 (N_5343,N_4758,N_3936);
xnor U5344 (N_5344,N_4452,N_3700);
nor U5345 (N_5345,N_3836,N_4740);
xor U5346 (N_5346,N_4002,N_4217);
nand U5347 (N_5347,N_4710,N_4642);
xor U5348 (N_5348,N_4247,N_4090);
and U5349 (N_5349,N_4214,N_4177);
nand U5350 (N_5350,N_4555,N_4388);
or U5351 (N_5351,N_3911,N_4316);
and U5352 (N_5352,N_4478,N_4012);
nor U5353 (N_5353,N_4073,N_4614);
and U5354 (N_5354,N_4569,N_4415);
or U5355 (N_5355,N_4314,N_3909);
or U5356 (N_5356,N_4646,N_3712);
or U5357 (N_5357,N_4142,N_3644);
xor U5358 (N_5358,N_4039,N_4163);
xor U5359 (N_5359,N_3813,N_3950);
nand U5360 (N_5360,N_4178,N_4131);
or U5361 (N_5361,N_4313,N_4210);
xor U5362 (N_5362,N_4366,N_4546);
or U5363 (N_5363,N_3966,N_4623);
xor U5364 (N_5364,N_4695,N_4434);
nand U5365 (N_5365,N_4718,N_4685);
and U5366 (N_5366,N_4505,N_4515);
xor U5367 (N_5367,N_4091,N_4287);
or U5368 (N_5368,N_3672,N_4542);
nand U5369 (N_5369,N_4292,N_4222);
or U5370 (N_5370,N_3870,N_4563);
nand U5371 (N_5371,N_4427,N_3844);
nor U5372 (N_5372,N_4079,N_4645);
and U5373 (N_5373,N_3820,N_3720);
xnor U5374 (N_5374,N_3953,N_4574);
xnor U5375 (N_5375,N_3906,N_3606);
xnor U5376 (N_5376,N_3614,N_4365);
nor U5377 (N_5377,N_3941,N_3762);
xnor U5378 (N_5378,N_3980,N_4370);
nand U5379 (N_5379,N_3695,N_4540);
nand U5380 (N_5380,N_3692,N_4696);
and U5381 (N_5381,N_3816,N_4025);
or U5382 (N_5382,N_4664,N_4496);
or U5383 (N_5383,N_4582,N_4159);
or U5384 (N_5384,N_3713,N_4127);
or U5385 (N_5385,N_4192,N_4756);
nand U5386 (N_5386,N_4257,N_3878);
or U5387 (N_5387,N_4634,N_4769);
or U5388 (N_5388,N_4700,N_4207);
xor U5389 (N_5389,N_3899,N_3742);
nand U5390 (N_5390,N_4742,N_4229);
nand U5391 (N_5391,N_4731,N_4195);
or U5392 (N_5392,N_4759,N_4202);
or U5393 (N_5393,N_4631,N_4280);
and U5394 (N_5394,N_3877,N_4597);
xnor U5395 (N_5395,N_4749,N_3871);
nand U5396 (N_5396,N_4282,N_3766);
nor U5397 (N_5397,N_4358,N_4402);
nand U5398 (N_5398,N_4789,N_4060);
nor U5399 (N_5399,N_3718,N_4283);
nand U5400 (N_5400,N_3969,N_3923);
and U5401 (N_5401,N_4479,N_4070);
or U5402 (N_5402,N_4608,N_3627);
and U5403 (N_5403,N_3993,N_4781);
nor U5404 (N_5404,N_4198,N_4021);
and U5405 (N_5405,N_3663,N_4568);
nor U5406 (N_5406,N_4736,N_4269);
and U5407 (N_5407,N_4522,N_4216);
and U5408 (N_5408,N_3905,N_4408);
nand U5409 (N_5409,N_3891,N_4689);
nor U5410 (N_5410,N_4445,N_3796);
nor U5411 (N_5411,N_4652,N_3774);
or U5412 (N_5412,N_4147,N_3632);
or U5413 (N_5413,N_4054,N_4124);
nor U5414 (N_5414,N_4683,N_3631);
nand U5415 (N_5415,N_3700,N_4732);
nand U5416 (N_5416,N_3870,N_4352);
xnor U5417 (N_5417,N_3678,N_4637);
nand U5418 (N_5418,N_4104,N_4500);
nor U5419 (N_5419,N_4765,N_4539);
nand U5420 (N_5420,N_4549,N_3732);
xor U5421 (N_5421,N_3632,N_4024);
nor U5422 (N_5422,N_4505,N_3691);
and U5423 (N_5423,N_4418,N_4040);
or U5424 (N_5424,N_4678,N_4784);
xnor U5425 (N_5425,N_4123,N_4323);
xor U5426 (N_5426,N_3914,N_4016);
nand U5427 (N_5427,N_3704,N_4133);
nand U5428 (N_5428,N_3978,N_4319);
xnor U5429 (N_5429,N_4011,N_4222);
nor U5430 (N_5430,N_3799,N_4775);
xnor U5431 (N_5431,N_4210,N_3685);
and U5432 (N_5432,N_3879,N_4565);
nor U5433 (N_5433,N_4752,N_3994);
or U5434 (N_5434,N_3624,N_4282);
nor U5435 (N_5435,N_3909,N_4723);
nor U5436 (N_5436,N_4423,N_4197);
nand U5437 (N_5437,N_3797,N_4397);
xnor U5438 (N_5438,N_4520,N_4076);
and U5439 (N_5439,N_4795,N_3633);
and U5440 (N_5440,N_4196,N_4459);
xnor U5441 (N_5441,N_4600,N_4066);
and U5442 (N_5442,N_3942,N_4776);
or U5443 (N_5443,N_4646,N_4331);
or U5444 (N_5444,N_3862,N_3789);
or U5445 (N_5445,N_4257,N_4699);
nand U5446 (N_5446,N_4699,N_4366);
and U5447 (N_5447,N_4707,N_4562);
nand U5448 (N_5448,N_4524,N_4043);
and U5449 (N_5449,N_4617,N_4063);
or U5450 (N_5450,N_4249,N_3919);
and U5451 (N_5451,N_4298,N_4467);
nor U5452 (N_5452,N_4344,N_4404);
xor U5453 (N_5453,N_4693,N_3739);
nor U5454 (N_5454,N_3974,N_4507);
or U5455 (N_5455,N_3622,N_4368);
xor U5456 (N_5456,N_3610,N_3940);
nand U5457 (N_5457,N_4135,N_4399);
and U5458 (N_5458,N_4651,N_4445);
nor U5459 (N_5459,N_4614,N_3897);
xnor U5460 (N_5460,N_4445,N_3966);
or U5461 (N_5461,N_4338,N_4544);
or U5462 (N_5462,N_4164,N_3974);
xor U5463 (N_5463,N_4023,N_4571);
xnor U5464 (N_5464,N_3645,N_4129);
nand U5465 (N_5465,N_4456,N_4002);
nor U5466 (N_5466,N_4752,N_3672);
nand U5467 (N_5467,N_4664,N_4208);
nor U5468 (N_5468,N_4358,N_3954);
nor U5469 (N_5469,N_4488,N_3838);
nand U5470 (N_5470,N_4086,N_4706);
xnor U5471 (N_5471,N_3680,N_3929);
nand U5472 (N_5472,N_3673,N_4477);
xnor U5473 (N_5473,N_4494,N_4625);
nand U5474 (N_5474,N_4281,N_3756);
nand U5475 (N_5475,N_4281,N_4462);
nand U5476 (N_5476,N_4139,N_4491);
nand U5477 (N_5477,N_3739,N_4525);
xnor U5478 (N_5478,N_4022,N_4061);
or U5479 (N_5479,N_4084,N_4201);
nand U5480 (N_5480,N_3784,N_4645);
nor U5481 (N_5481,N_3701,N_4571);
nor U5482 (N_5482,N_4314,N_4679);
nor U5483 (N_5483,N_3902,N_3653);
xor U5484 (N_5484,N_4445,N_3905);
or U5485 (N_5485,N_4307,N_3708);
nor U5486 (N_5486,N_4159,N_3948);
or U5487 (N_5487,N_3957,N_4441);
or U5488 (N_5488,N_3837,N_3678);
or U5489 (N_5489,N_3963,N_3858);
nor U5490 (N_5490,N_3696,N_4571);
xor U5491 (N_5491,N_4504,N_4702);
or U5492 (N_5492,N_4235,N_4447);
nor U5493 (N_5493,N_3795,N_4611);
nand U5494 (N_5494,N_3654,N_4650);
nand U5495 (N_5495,N_4237,N_4067);
or U5496 (N_5496,N_4125,N_4690);
nor U5497 (N_5497,N_4745,N_4553);
xnor U5498 (N_5498,N_4007,N_3611);
xnor U5499 (N_5499,N_4305,N_3844);
nand U5500 (N_5500,N_3652,N_4651);
or U5501 (N_5501,N_4785,N_3924);
or U5502 (N_5502,N_4044,N_4563);
xor U5503 (N_5503,N_4395,N_4381);
xor U5504 (N_5504,N_3663,N_3705);
xor U5505 (N_5505,N_4412,N_4554);
xnor U5506 (N_5506,N_4160,N_3965);
xor U5507 (N_5507,N_3634,N_4626);
xor U5508 (N_5508,N_4671,N_4659);
or U5509 (N_5509,N_3993,N_4480);
nand U5510 (N_5510,N_4690,N_4217);
and U5511 (N_5511,N_4384,N_4666);
xnor U5512 (N_5512,N_4023,N_3994);
or U5513 (N_5513,N_3776,N_3762);
xor U5514 (N_5514,N_3811,N_3883);
or U5515 (N_5515,N_3784,N_4321);
xnor U5516 (N_5516,N_4457,N_3721);
nand U5517 (N_5517,N_4212,N_3699);
or U5518 (N_5518,N_4026,N_4609);
xor U5519 (N_5519,N_3973,N_3881);
or U5520 (N_5520,N_4023,N_3769);
or U5521 (N_5521,N_3956,N_4039);
or U5522 (N_5522,N_3679,N_4265);
or U5523 (N_5523,N_4028,N_4444);
xnor U5524 (N_5524,N_4141,N_3675);
and U5525 (N_5525,N_3673,N_4422);
nand U5526 (N_5526,N_3850,N_4770);
and U5527 (N_5527,N_3994,N_3687);
nand U5528 (N_5528,N_4458,N_4732);
and U5529 (N_5529,N_4487,N_3636);
nor U5530 (N_5530,N_4692,N_3977);
nand U5531 (N_5531,N_3649,N_4386);
or U5532 (N_5532,N_3649,N_4347);
xnor U5533 (N_5533,N_3799,N_3894);
and U5534 (N_5534,N_4615,N_4138);
nand U5535 (N_5535,N_4737,N_4377);
xor U5536 (N_5536,N_3715,N_4709);
xnor U5537 (N_5537,N_4003,N_4136);
nor U5538 (N_5538,N_4586,N_4495);
or U5539 (N_5539,N_4376,N_4117);
xnor U5540 (N_5540,N_4551,N_3611);
or U5541 (N_5541,N_4714,N_4557);
or U5542 (N_5542,N_3918,N_4655);
and U5543 (N_5543,N_3977,N_4216);
nand U5544 (N_5544,N_4635,N_4064);
xor U5545 (N_5545,N_4196,N_3621);
or U5546 (N_5546,N_3908,N_4516);
and U5547 (N_5547,N_4309,N_3808);
and U5548 (N_5548,N_4417,N_3945);
nor U5549 (N_5549,N_3682,N_4339);
or U5550 (N_5550,N_4742,N_4717);
nand U5551 (N_5551,N_3615,N_4421);
nor U5552 (N_5552,N_4161,N_4606);
xor U5553 (N_5553,N_3785,N_4183);
and U5554 (N_5554,N_4183,N_4699);
xnor U5555 (N_5555,N_3776,N_4376);
xnor U5556 (N_5556,N_4324,N_4614);
nand U5557 (N_5557,N_4681,N_4380);
or U5558 (N_5558,N_4442,N_3619);
or U5559 (N_5559,N_4262,N_4053);
nor U5560 (N_5560,N_4364,N_4061);
nand U5561 (N_5561,N_4427,N_4758);
xor U5562 (N_5562,N_4793,N_4115);
nor U5563 (N_5563,N_4538,N_4761);
or U5564 (N_5564,N_3623,N_3844);
nor U5565 (N_5565,N_4417,N_4295);
xor U5566 (N_5566,N_4066,N_4736);
nand U5567 (N_5567,N_4475,N_4014);
nand U5568 (N_5568,N_4038,N_4168);
nand U5569 (N_5569,N_4634,N_4732);
xnor U5570 (N_5570,N_4019,N_4163);
or U5571 (N_5571,N_3747,N_4354);
or U5572 (N_5572,N_4625,N_3936);
and U5573 (N_5573,N_4358,N_4282);
nand U5574 (N_5574,N_4401,N_4627);
nand U5575 (N_5575,N_4679,N_3826);
or U5576 (N_5576,N_3894,N_4746);
and U5577 (N_5577,N_4076,N_4392);
and U5578 (N_5578,N_3962,N_4130);
nand U5579 (N_5579,N_3720,N_4583);
nor U5580 (N_5580,N_4420,N_4406);
nand U5581 (N_5581,N_4216,N_3828);
or U5582 (N_5582,N_4619,N_4546);
or U5583 (N_5583,N_3616,N_4665);
nand U5584 (N_5584,N_4611,N_4205);
nor U5585 (N_5585,N_4450,N_4092);
nor U5586 (N_5586,N_4617,N_4098);
nand U5587 (N_5587,N_4047,N_4580);
or U5588 (N_5588,N_3969,N_4368);
and U5589 (N_5589,N_4559,N_3925);
and U5590 (N_5590,N_4559,N_3708);
nand U5591 (N_5591,N_4615,N_4169);
nand U5592 (N_5592,N_4699,N_4671);
and U5593 (N_5593,N_3969,N_4042);
or U5594 (N_5594,N_4391,N_4761);
and U5595 (N_5595,N_3980,N_4434);
or U5596 (N_5596,N_3932,N_4044);
nor U5597 (N_5597,N_3739,N_4376);
and U5598 (N_5598,N_4141,N_4208);
nand U5599 (N_5599,N_4531,N_3818);
and U5600 (N_5600,N_4453,N_3641);
and U5601 (N_5601,N_4548,N_4118);
nor U5602 (N_5602,N_3639,N_3618);
and U5603 (N_5603,N_3993,N_3717);
xor U5604 (N_5604,N_3987,N_4292);
nand U5605 (N_5605,N_4550,N_3843);
and U5606 (N_5606,N_4424,N_3978);
or U5607 (N_5607,N_4303,N_3775);
nand U5608 (N_5608,N_3770,N_4555);
nand U5609 (N_5609,N_3796,N_3919);
xnor U5610 (N_5610,N_3812,N_4143);
nand U5611 (N_5611,N_4365,N_3755);
nor U5612 (N_5612,N_3790,N_3604);
xor U5613 (N_5613,N_3790,N_4412);
or U5614 (N_5614,N_4534,N_4359);
xor U5615 (N_5615,N_4255,N_4722);
or U5616 (N_5616,N_4339,N_4417);
or U5617 (N_5617,N_3623,N_4725);
xnor U5618 (N_5618,N_3661,N_4128);
nand U5619 (N_5619,N_4229,N_4534);
and U5620 (N_5620,N_3794,N_4436);
nand U5621 (N_5621,N_3636,N_3851);
nand U5622 (N_5622,N_4188,N_4286);
and U5623 (N_5623,N_4304,N_3721);
nor U5624 (N_5624,N_4199,N_4218);
nor U5625 (N_5625,N_4198,N_4664);
nor U5626 (N_5626,N_4040,N_4328);
or U5627 (N_5627,N_3749,N_4587);
xnor U5628 (N_5628,N_3654,N_4633);
nand U5629 (N_5629,N_3689,N_4110);
and U5630 (N_5630,N_4504,N_4349);
xnor U5631 (N_5631,N_4295,N_3764);
nor U5632 (N_5632,N_3792,N_3880);
or U5633 (N_5633,N_4619,N_4298);
or U5634 (N_5634,N_3827,N_4785);
and U5635 (N_5635,N_3917,N_3726);
or U5636 (N_5636,N_4010,N_4099);
xor U5637 (N_5637,N_3758,N_4428);
xor U5638 (N_5638,N_4078,N_3793);
xnor U5639 (N_5639,N_4652,N_4568);
and U5640 (N_5640,N_3824,N_3635);
nand U5641 (N_5641,N_4303,N_4585);
nand U5642 (N_5642,N_4010,N_4752);
nor U5643 (N_5643,N_4528,N_3933);
nand U5644 (N_5644,N_3992,N_3834);
xor U5645 (N_5645,N_4394,N_4037);
nand U5646 (N_5646,N_4704,N_4387);
or U5647 (N_5647,N_4309,N_4371);
or U5648 (N_5648,N_3773,N_4575);
or U5649 (N_5649,N_4035,N_4532);
nand U5650 (N_5650,N_4377,N_3782);
and U5651 (N_5651,N_3726,N_4166);
or U5652 (N_5652,N_4138,N_4455);
xor U5653 (N_5653,N_3950,N_4223);
or U5654 (N_5654,N_3876,N_4299);
nand U5655 (N_5655,N_4678,N_4421);
and U5656 (N_5656,N_4128,N_4760);
and U5657 (N_5657,N_4400,N_3691);
xnor U5658 (N_5658,N_3835,N_4297);
nand U5659 (N_5659,N_3898,N_3914);
nand U5660 (N_5660,N_4397,N_3669);
nand U5661 (N_5661,N_4388,N_4110);
nand U5662 (N_5662,N_3907,N_3615);
or U5663 (N_5663,N_4397,N_3932);
and U5664 (N_5664,N_4366,N_4080);
nor U5665 (N_5665,N_3640,N_4396);
or U5666 (N_5666,N_3602,N_4325);
nand U5667 (N_5667,N_4629,N_3736);
nand U5668 (N_5668,N_3876,N_4019);
or U5669 (N_5669,N_3706,N_3955);
or U5670 (N_5670,N_3774,N_4605);
xor U5671 (N_5671,N_3708,N_4362);
and U5672 (N_5672,N_3944,N_4465);
and U5673 (N_5673,N_3862,N_3717);
nand U5674 (N_5674,N_4755,N_4164);
and U5675 (N_5675,N_3909,N_4322);
nand U5676 (N_5676,N_4089,N_3777);
nor U5677 (N_5677,N_3603,N_4134);
xor U5678 (N_5678,N_3797,N_4135);
nor U5679 (N_5679,N_4131,N_4237);
or U5680 (N_5680,N_4330,N_4732);
xnor U5681 (N_5681,N_4116,N_4433);
xnor U5682 (N_5682,N_4255,N_3631);
nor U5683 (N_5683,N_3649,N_3681);
or U5684 (N_5684,N_4314,N_4695);
and U5685 (N_5685,N_4769,N_4313);
and U5686 (N_5686,N_4014,N_4689);
and U5687 (N_5687,N_4446,N_4787);
nor U5688 (N_5688,N_4021,N_3966);
and U5689 (N_5689,N_3744,N_4468);
or U5690 (N_5690,N_4322,N_4157);
nand U5691 (N_5691,N_3832,N_4361);
xnor U5692 (N_5692,N_4417,N_4757);
nand U5693 (N_5693,N_4264,N_4200);
or U5694 (N_5694,N_4563,N_4295);
xnor U5695 (N_5695,N_4649,N_4556);
nand U5696 (N_5696,N_4581,N_4729);
xor U5697 (N_5697,N_3974,N_3759);
nand U5698 (N_5698,N_4442,N_4298);
nand U5699 (N_5699,N_4272,N_4451);
or U5700 (N_5700,N_4291,N_3948);
nor U5701 (N_5701,N_4514,N_3749);
xor U5702 (N_5702,N_4658,N_4298);
or U5703 (N_5703,N_3752,N_3792);
or U5704 (N_5704,N_4673,N_3814);
nor U5705 (N_5705,N_4527,N_4544);
xor U5706 (N_5706,N_4434,N_4175);
xnor U5707 (N_5707,N_4729,N_4220);
nand U5708 (N_5708,N_4440,N_4658);
nor U5709 (N_5709,N_3829,N_4371);
or U5710 (N_5710,N_4542,N_3882);
nand U5711 (N_5711,N_4261,N_4287);
nor U5712 (N_5712,N_4577,N_4256);
nand U5713 (N_5713,N_3639,N_3992);
xnor U5714 (N_5714,N_3684,N_3876);
and U5715 (N_5715,N_4287,N_4729);
xor U5716 (N_5716,N_4402,N_3795);
and U5717 (N_5717,N_4193,N_4230);
or U5718 (N_5718,N_4626,N_3713);
or U5719 (N_5719,N_4177,N_4668);
nor U5720 (N_5720,N_4533,N_4505);
and U5721 (N_5721,N_4108,N_4506);
xor U5722 (N_5722,N_4751,N_4651);
xnor U5723 (N_5723,N_4282,N_4024);
or U5724 (N_5724,N_3699,N_4725);
and U5725 (N_5725,N_4026,N_4557);
xor U5726 (N_5726,N_3698,N_3811);
and U5727 (N_5727,N_3670,N_4404);
or U5728 (N_5728,N_3646,N_4706);
nor U5729 (N_5729,N_4108,N_4427);
xor U5730 (N_5730,N_4685,N_4536);
xor U5731 (N_5731,N_3818,N_4481);
and U5732 (N_5732,N_4086,N_4224);
nand U5733 (N_5733,N_3918,N_3782);
nor U5734 (N_5734,N_4758,N_3746);
nor U5735 (N_5735,N_4532,N_4624);
xor U5736 (N_5736,N_4203,N_4263);
or U5737 (N_5737,N_4339,N_3662);
nand U5738 (N_5738,N_4122,N_3714);
or U5739 (N_5739,N_4203,N_4416);
nand U5740 (N_5740,N_3606,N_4017);
nor U5741 (N_5741,N_4794,N_4270);
xnor U5742 (N_5742,N_3871,N_4152);
xnor U5743 (N_5743,N_3678,N_3963);
nor U5744 (N_5744,N_4270,N_4510);
xnor U5745 (N_5745,N_4477,N_4355);
nor U5746 (N_5746,N_4761,N_4625);
nor U5747 (N_5747,N_3685,N_3888);
or U5748 (N_5748,N_4113,N_4525);
nand U5749 (N_5749,N_4110,N_4783);
and U5750 (N_5750,N_3808,N_3896);
nor U5751 (N_5751,N_3960,N_4675);
xnor U5752 (N_5752,N_4454,N_3695);
nand U5753 (N_5753,N_4458,N_4143);
or U5754 (N_5754,N_3833,N_3944);
or U5755 (N_5755,N_4517,N_4035);
and U5756 (N_5756,N_4576,N_3963);
nor U5757 (N_5757,N_4324,N_4677);
nor U5758 (N_5758,N_4072,N_4508);
and U5759 (N_5759,N_4384,N_3947);
or U5760 (N_5760,N_3623,N_4478);
or U5761 (N_5761,N_3849,N_4421);
xor U5762 (N_5762,N_4488,N_4579);
and U5763 (N_5763,N_3885,N_4667);
xor U5764 (N_5764,N_4648,N_3736);
and U5765 (N_5765,N_4420,N_4309);
and U5766 (N_5766,N_4624,N_4616);
xnor U5767 (N_5767,N_3910,N_3621);
xnor U5768 (N_5768,N_4595,N_4536);
xor U5769 (N_5769,N_4006,N_4648);
xor U5770 (N_5770,N_4230,N_4595);
nand U5771 (N_5771,N_4583,N_4735);
nand U5772 (N_5772,N_4462,N_3806);
nand U5773 (N_5773,N_4526,N_4670);
and U5774 (N_5774,N_4075,N_3877);
nand U5775 (N_5775,N_4483,N_4549);
xor U5776 (N_5776,N_3806,N_4735);
and U5777 (N_5777,N_3894,N_4195);
and U5778 (N_5778,N_4543,N_4547);
or U5779 (N_5779,N_4313,N_4173);
nand U5780 (N_5780,N_3634,N_4419);
nand U5781 (N_5781,N_4735,N_4442);
and U5782 (N_5782,N_3692,N_4624);
or U5783 (N_5783,N_3973,N_3928);
nor U5784 (N_5784,N_4194,N_4342);
nor U5785 (N_5785,N_4187,N_4756);
nand U5786 (N_5786,N_4240,N_4400);
nand U5787 (N_5787,N_3847,N_3617);
nor U5788 (N_5788,N_4033,N_3945);
and U5789 (N_5789,N_3804,N_4471);
xnor U5790 (N_5790,N_3970,N_3663);
or U5791 (N_5791,N_4147,N_4464);
nand U5792 (N_5792,N_3954,N_4673);
nor U5793 (N_5793,N_3830,N_3992);
nand U5794 (N_5794,N_4775,N_4297);
or U5795 (N_5795,N_3991,N_4240);
and U5796 (N_5796,N_4427,N_4144);
or U5797 (N_5797,N_3860,N_4182);
or U5798 (N_5798,N_3975,N_3931);
and U5799 (N_5799,N_4442,N_4276);
xor U5800 (N_5800,N_3628,N_3878);
nor U5801 (N_5801,N_3612,N_4199);
nor U5802 (N_5802,N_4450,N_4071);
xor U5803 (N_5803,N_4682,N_4072);
or U5804 (N_5804,N_4533,N_3613);
xor U5805 (N_5805,N_3880,N_3864);
nor U5806 (N_5806,N_4016,N_4534);
or U5807 (N_5807,N_4182,N_3717);
and U5808 (N_5808,N_4580,N_4162);
nand U5809 (N_5809,N_4131,N_4597);
nand U5810 (N_5810,N_4339,N_4471);
or U5811 (N_5811,N_4386,N_3644);
xnor U5812 (N_5812,N_4578,N_4507);
nand U5813 (N_5813,N_3973,N_3683);
nand U5814 (N_5814,N_4265,N_4494);
and U5815 (N_5815,N_4329,N_4388);
or U5816 (N_5816,N_4121,N_4306);
nor U5817 (N_5817,N_4580,N_3810);
or U5818 (N_5818,N_4650,N_3704);
and U5819 (N_5819,N_4300,N_4124);
or U5820 (N_5820,N_4476,N_4680);
xor U5821 (N_5821,N_4094,N_4466);
xnor U5822 (N_5822,N_4371,N_4043);
nor U5823 (N_5823,N_4215,N_4009);
and U5824 (N_5824,N_3979,N_3734);
nand U5825 (N_5825,N_3663,N_4041);
or U5826 (N_5826,N_4617,N_4732);
or U5827 (N_5827,N_4327,N_4190);
xnor U5828 (N_5828,N_4206,N_4762);
nor U5829 (N_5829,N_4189,N_3919);
nor U5830 (N_5830,N_4052,N_3673);
or U5831 (N_5831,N_4272,N_3612);
nand U5832 (N_5832,N_4685,N_4000);
xor U5833 (N_5833,N_4468,N_4457);
or U5834 (N_5834,N_4331,N_3883);
and U5835 (N_5835,N_3928,N_4779);
and U5836 (N_5836,N_3992,N_3699);
or U5837 (N_5837,N_3936,N_3980);
xnor U5838 (N_5838,N_4209,N_4290);
nor U5839 (N_5839,N_4449,N_4310);
nand U5840 (N_5840,N_3755,N_4410);
nand U5841 (N_5841,N_3975,N_4716);
and U5842 (N_5842,N_3624,N_4248);
or U5843 (N_5843,N_4624,N_4191);
nand U5844 (N_5844,N_4686,N_4070);
nand U5845 (N_5845,N_4542,N_3781);
nand U5846 (N_5846,N_4340,N_4262);
or U5847 (N_5847,N_4065,N_4769);
xor U5848 (N_5848,N_3701,N_3651);
nor U5849 (N_5849,N_3810,N_4431);
nor U5850 (N_5850,N_3704,N_3604);
nand U5851 (N_5851,N_4677,N_4755);
or U5852 (N_5852,N_3683,N_4283);
nand U5853 (N_5853,N_4237,N_3938);
nor U5854 (N_5854,N_4581,N_3991);
nand U5855 (N_5855,N_4541,N_4375);
xnor U5856 (N_5856,N_3768,N_3986);
xnor U5857 (N_5857,N_4518,N_4211);
or U5858 (N_5858,N_4794,N_4269);
or U5859 (N_5859,N_3729,N_3993);
nor U5860 (N_5860,N_3762,N_4484);
or U5861 (N_5861,N_3801,N_3772);
or U5862 (N_5862,N_4720,N_3986);
nand U5863 (N_5863,N_3624,N_3873);
and U5864 (N_5864,N_4242,N_4256);
and U5865 (N_5865,N_4703,N_3602);
nand U5866 (N_5866,N_4755,N_4113);
nand U5867 (N_5867,N_4739,N_4092);
and U5868 (N_5868,N_4334,N_4063);
and U5869 (N_5869,N_3664,N_4529);
or U5870 (N_5870,N_3689,N_3916);
xor U5871 (N_5871,N_3774,N_3671);
nor U5872 (N_5872,N_4411,N_4047);
or U5873 (N_5873,N_3747,N_4064);
xor U5874 (N_5874,N_4516,N_3628);
or U5875 (N_5875,N_4106,N_4175);
nand U5876 (N_5876,N_4396,N_3831);
and U5877 (N_5877,N_4361,N_4330);
xnor U5878 (N_5878,N_4764,N_3773);
nand U5879 (N_5879,N_4329,N_3658);
nor U5880 (N_5880,N_4079,N_4736);
or U5881 (N_5881,N_4424,N_4437);
or U5882 (N_5882,N_4135,N_3811);
xnor U5883 (N_5883,N_4451,N_4052);
nor U5884 (N_5884,N_4749,N_4406);
nand U5885 (N_5885,N_4770,N_3921);
and U5886 (N_5886,N_3637,N_4674);
and U5887 (N_5887,N_4355,N_4070);
nand U5888 (N_5888,N_4751,N_4044);
and U5889 (N_5889,N_3918,N_4084);
xor U5890 (N_5890,N_3876,N_3878);
or U5891 (N_5891,N_3970,N_4484);
nor U5892 (N_5892,N_4510,N_4190);
nor U5893 (N_5893,N_4223,N_4690);
and U5894 (N_5894,N_3674,N_4476);
or U5895 (N_5895,N_3915,N_4559);
xor U5896 (N_5896,N_4062,N_3770);
xnor U5897 (N_5897,N_4539,N_4719);
or U5898 (N_5898,N_4397,N_3764);
nor U5899 (N_5899,N_4579,N_3721);
nand U5900 (N_5900,N_4616,N_3772);
nor U5901 (N_5901,N_3606,N_3887);
xor U5902 (N_5902,N_4207,N_4493);
nor U5903 (N_5903,N_4092,N_4511);
xnor U5904 (N_5904,N_4283,N_3854);
nand U5905 (N_5905,N_4660,N_4746);
or U5906 (N_5906,N_3821,N_3901);
xnor U5907 (N_5907,N_4212,N_4792);
xor U5908 (N_5908,N_4121,N_4225);
nand U5909 (N_5909,N_4114,N_4016);
or U5910 (N_5910,N_4374,N_3927);
and U5911 (N_5911,N_4566,N_4061);
nand U5912 (N_5912,N_4404,N_4446);
and U5913 (N_5913,N_4522,N_3707);
or U5914 (N_5914,N_4659,N_4197);
or U5915 (N_5915,N_4542,N_4599);
and U5916 (N_5916,N_4180,N_4536);
or U5917 (N_5917,N_4351,N_4630);
nor U5918 (N_5918,N_3622,N_4324);
xnor U5919 (N_5919,N_4684,N_4290);
nand U5920 (N_5920,N_4625,N_4683);
xor U5921 (N_5921,N_4556,N_4342);
xnor U5922 (N_5922,N_4081,N_4744);
nor U5923 (N_5923,N_3787,N_3783);
nand U5924 (N_5924,N_4408,N_4692);
and U5925 (N_5925,N_3626,N_4272);
nor U5926 (N_5926,N_4649,N_3708);
and U5927 (N_5927,N_4680,N_4577);
xor U5928 (N_5928,N_4787,N_4530);
or U5929 (N_5929,N_3739,N_3608);
nand U5930 (N_5930,N_4545,N_4587);
and U5931 (N_5931,N_3741,N_4119);
nand U5932 (N_5932,N_4282,N_4286);
xnor U5933 (N_5933,N_4586,N_4050);
xnor U5934 (N_5934,N_4667,N_4501);
nand U5935 (N_5935,N_4372,N_4382);
xor U5936 (N_5936,N_3914,N_4336);
and U5937 (N_5937,N_4357,N_3704);
or U5938 (N_5938,N_4599,N_4406);
or U5939 (N_5939,N_4576,N_4757);
nor U5940 (N_5940,N_4643,N_4763);
nand U5941 (N_5941,N_4576,N_4027);
or U5942 (N_5942,N_3707,N_3755);
xor U5943 (N_5943,N_4241,N_3797);
nand U5944 (N_5944,N_3824,N_4679);
or U5945 (N_5945,N_3642,N_3745);
and U5946 (N_5946,N_4252,N_3989);
nor U5947 (N_5947,N_4352,N_4374);
nand U5948 (N_5948,N_4044,N_3961);
nor U5949 (N_5949,N_4304,N_4078);
nand U5950 (N_5950,N_4507,N_4291);
or U5951 (N_5951,N_4353,N_4121);
xnor U5952 (N_5952,N_4194,N_3941);
nand U5953 (N_5953,N_3645,N_3942);
nand U5954 (N_5954,N_4597,N_4155);
nor U5955 (N_5955,N_4380,N_3668);
xor U5956 (N_5956,N_3797,N_3961);
and U5957 (N_5957,N_4453,N_3657);
or U5958 (N_5958,N_4195,N_4144);
or U5959 (N_5959,N_3917,N_4501);
or U5960 (N_5960,N_3607,N_4452);
nor U5961 (N_5961,N_4257,N_4045);
xnor U5962 (N_5962,N_4576,N_3983);
xnor U5963 (N_5963,N_4446,N_3685);
or U5964 (N_5964,N_4512,N_4631);
nand U5965 (N_5965,N_3771,N_4053);
and U5966 (N_5966,N_4778,N_3871);
nand U5967 (N_5967,N_4265,N_4071);
nor U5968 (N_5968,N_3606,N_4054);
nor U5969 (N_5969,N_4595,N_4550);
and U5970 (N_5970,N_4488,N_4526);
or U5971 (N_5971,N_4764,N_3611);
or U5972 (N_5972,N_3752,N_3946);
xnor U5973 (N_5973,N_4427,N_4512);
or U5974 (N_5974,N_3885,N_4583);
and U5975 (N_5975,N_3959,N_4555);
nand U5976 (N_5976,N_4262,N_4207);
nor U5977 (N_5977,N_3930,N_4624);
or U5978 (N_5978,N_4395,N_3701);
xnor U5979 (N_5979,N_4572,N_3727);
nand U5980 (N_5980,N_3841,N_4368);
nor U5981 (N_5981,N_4647,N_4237);
and U5982 (N_5982,N_4687,N_4749);
and U5983 (N_5983,N_3614,N_3877);
and U5984 (N_5984,N_3877,N_4590);
or U5985 (N_5985,N_3648,N_4197);
xor U5986 (N_5986,N_4136,N_3827);
nor U5987 (N_5987,N_4198,N_4210);
or U5988 (N_5988,N_4602,N_4734);
or U5989 (N_5989,N_4196,N_4370);
nand U5990 (N_5990,N_4633,N_4022);
nor U5991 (N_5991,N_3856,N_4156);
nor U5992 (N_5992,N_3841,N_4634);
or U5993 (N_5993,N_3795,N_4280);
or U5994 (N_5994,N_3683,N_4199);
xor U5995 (N_5995,N_4092,N_4001);
nor U5996 (N_5996,N_4598,N_4661);
and U5997 (N_5997,N_4095,N_4256);
and U5998 (N_5998,N_4752,N_4040);
nand U5999 (N_5999,N_4028,N_4529);
or U6000 (N_6000,N_5589,N_5818);
and U6001 (N_6001,N_5267,N_4813);
or U6002 (N_6002,N_5629,N_5316);
xnor U6003 (N_6003,N_5324,N_5740);
xnor U6004 (N_6004,N_5081,N_5386);
nor U6005 (N_6005,N_5605,N_5608);
or U6006 (N_6006,N_5652,N_5349);
nor U6007 (N_6007,N_4982,N_5735);
xor U6008 (N_6008,N_5283,N_5343);
nor U6009 (N_6009,N_5725,N_4820);
or U6010 (N_6010,N_4938,N_5213);
and U6011 (N_6011,N_5557,N_5759);
nor U6012 (N_6012,N_5295,N_5761);
nand U6013 (N_6013,N_5160,N_5001);
nor U6014 (N_6014,N_5253,N_5974);
xnor U6015 (N_6015,N_5126,N_5808);
xnor U6016 (N_6016,N_5799,N_5143);
nor U6017 (N_6017,N_5811,N_5565);
nand U6018 (N_6018,N_5127,N_5035);
and U6019 (N_6019,N_5642,N_5959);
and U6020 (N_6020,N_5902,N_5226);
nand U6021 (N_6021,N_5996,N_5678);
and U6022 (N_6022,N_5699,N_5390);
and U6023 (N_6023,N_4847,N_5745);
and U6024 (N_6024,N_5979,N_4921);
nor U6025 (N_6025,N_5185,N_5013);
nand U6026 (N_6026,N_5111,N_4880);
and U6027 (N_6027,N_5654,N_5675);
and U6028 (N_6028,N_5406,N_5950);
nor U6029 (N_6029,N_5792,N_5003);
nor U6030 (N_6030,N_4931,N_5869);
xor U6031 (N_6031,N_5716,N_5870);
nor U6032 (N_6032,N_4856,N_4935);
and U6033 (N_6033,N_4869,N_5090);
nor U6034 (N_6034,N_4929,N_5362);
and U6035 (N_6035,N_5899,N_4802);
nand U6036 (N_6036,N_5278,N_5795);
and U6037 (N_6037,N_5914,N_5169);
and U6038 (N_6038,N_5783,N_5655);
and U6039 (N_6039,N_5232,N_5167);
nand U6040 (N_6040,N_5038,N_5796);
xor U6041 (N_6041,N_4867,N_5002);
xor U6042 (N_6042,N_5322,N_4848);
xor U6043 (N_6043,N_4837,N_5918);
nand U6044 (N_6044,N_5022,N_5115);
and U6045 (N_6045,N_5692,N_5906);
or U6046 (N_6046,N_4834,N_5104);
xnor U6047 (N_6047,N_5216,N_5643);
nor U6048 (N_6048,N_4971,N_5339);
nand U6049 (N_6049,N_5769,N_5261);
and U6050 (N_6050,N_5572,N_4927);
or U6051 (N_6051,N_5314,N_5434);
xnor U6052 (N_6052,N_5384,N_5068);
nand U6053 (N_6053,N_5426,N_5802);
xor U6054 (N_6054,N_5351,N_5919);
nand U6055 (N_6055,N_5884,N_5530);
and U6056 (N_6056,N_5536,N_5435);
xor U6057 (N_6057,N_5177,N_4955);
nor U6058 (N_6058,N_5487,N_5703);
and U6059 (N_6059,N_5566,N_5989);
and U6060 (N_6060,N_4859,N_5052);
nand U6061 (N_6061,N_5952,N_5192);
nor U6062 (N_6062,N_5024,N_5453);
nand U6063 (N_6063,N_5449,N_5303);
nand U6064 (N_6064,N_5910,N_5864);
nor U6065 (N_6065,N_4868,N_5866);
or U6066 (N_6066,N_5455,N_5405);
nand U6067 (N_6067,N_5586,N_5971);
and U6068 (N_6068,N_5999,N_5903);
nor U6069 (N_6069,N_4969,N_5410);
or U6070 (N_6070,N_5420,N_4894);
and U6071 (N_6071,N_5970,N_5542);
or U6072 (N_6072,N_5496,N_5008);
xor U6073 (N_6073,N_5293,N_5086);
nor U6074 (N_6074,N_4887,N_5797);
nand U6075 (N_6075,N_4806,N_5562);
nor U6076 (N_6076,N_5116,N_5300);
or U6077 (N_6077,N_5590,N_5354);
or U6078 (N_6078,N_5569,N_5584);
xnor U6079 (N_6079,N_5737,N_5581);
xor U6080 (N_6080,N_5229,N_5306);
nor U6081 (N_6081,N_5645,N_5066);
or U6082 (N_6082,N_5345,N_5934);
and U6083 (N_6083,N_5443,N_5875);
nor U6084 (N_6084,N_5025,N_5028);
or U6085 (N_6085,N_5534,N_5555);
nor U6086 (N_6086,N_5129,N_5271);
or U6087 (N_6087,N_5431,N_4947);
and U6088 (N_6088,N_4832,N_5578);
nor U6089 (N_6089,N_5892,N_4904);
nand U6090 (N_6090,N_4956,N_5401);
nand U6091 (N_6091,N_5720,N_5809);
and U6092 (N_6092,N_4844,N_4899);
or U6093 (N_6093,N_5398,N_5612);
nor U6094 (N_6094,N_4811,N_5516);
nand U6095 (N_6095,N_5347,N_5098);
or U6096 (N_6096,N_5641,N_5011);
nand U6097 (N_6097,N_5459,N_5913);
or U6098 (N_6098,N_5844,N_5871);
nor U6099 (N_6099,N_5452,N_5742);
xnor U6100 (N_6100,N_5299,N_5123);
xor U6101 (N_6101,N_5489,N_5576);
nor U6102 (N_6102,N_5393,N_5446);
or U6103 (N_6103,N_4974,N_5812);
xnor U6104 (N_6104,N_5364,N_5760);
nor U6105 (N_6105,N_5616,N_5805);
nand U6106 (N_6106,N_5515,N_4817);
or U6107 (N_6107,N_5658,N_5858);
or U6108 (N_6108,N_5718,N_5266);
and U6109 (N_6109,N_5631,N_5574);
or U6110 (N_6110,N_5281,N_5845);
nor U6111 (N_6111,N_5419,N_4916);
nand U6112 (N_6112,N_5311,N_5307);
nor U6113 (N_6113,N_5456,N_4901);
xnor U6114 (N_6114,N_5156,N_5243);
nand U6115 (N_6115,N_5724,N_5147);
nand U6116 (N_6116,N_5776,N_5150);
and U6117 (N_6117,N_5888,N_5772);
nor U6118 (N_6118,N_5548,N_4959);
or U6119 (N_6119,N_5212,N_5747);
xnor U6120 (N_6120,N_5075,N_5492);
or U6121 (N_6121,N_5089,N_4997);
or U6122 (N_6122,N_4895,N_5834);
or U6123 (N_6123,N_5611,N_5210);
nand U6124 (N_6124,N_5626,N_5882);
and U6125 (N_6125,N_5744,N_5943);
and U6126 (N_6126,N_5662,N_5620);
and U6127 (N_6127,N_5319,N_5920);
nand U6128 (N_6128,N_4906,N_4851);
nor U6129 (N_6129,N_4908,N_5695);
and U6130 (N_6130,N_5831,N_5137);
or U6131 (N_6131,N_4865,N_4841);
nor U6132 (N_6132,N_4958,N_5828);
and U6133 (N_6133,N_5621,N_5255);
nand U6134 (N_6134,N_4885,N_5694);
and U6135 (N_6135,N_5606,N_5832);
and U6136 (N_6136,N_5738,N_4824);
xnor U6137 (N_6137,N_5817,N_5535);
nor U6138 (N_6138,N_5335,N_5579);
xor U6139 (N_6139,N_5121,N_4888);
and U6140 (N_6140,N_5385,N_5117);
or U6141 (N_6141,N_4877,N_5248);
or U6142 (N_6142,N_5264,N_5750);
nor U6143 (N_6143,N_5976,N_5768);
and U6144 (N_6144,N_5173,N_5027);
nor U6145 (N_6145,N_4976,N_4989);
and U6146 (N_6146,N_5545,N_5225);
nor U6147 (N_6147,N_5998,N_5342);
or U6148 (N_6148,N_5184,N_5191);
xnor U6149 (N_6149,N_5045,N_5704);
or U6150 (N_6150,N_5285,N_5915);
nand U6151 (N_6151,N_5337,N_5269);
nand U6152 (N_6152,N_5897,N_5767);
xnor U6153 (N_6153,N_4900,N_5290);
nand U6154 (N_6154,N_5208,N_5119);
nand U6155 (N_6155,N_5949,N_5848);
or U6156 (N_6156,N_5830,N_5042);
or U6157 (N_6157,N_4858,N_5272);
or U6158 (N_6158,N_5023,N_5188);
or U6159 (N_6159,N_5244,N_4953);
nand U6160 (N_6160,N_5790,N_5930);
and U6161 (N_6161,N_5701,N_5541);
nand U6162 (N_6162,N_5540,N_5057);
xnor U6163 (N_6163,N_5228,N_5366);
nand U6164 (N_6164,N_5961,N_4804);
nand U6165 (N_6165,N_5263,N_4928);
and U6166 (N_6166,N_4998,N_5682);
and U6167 (N_6167,N_5741,N_5344);
or U6168 (N_6168,N_5883,N_5528);
xnor U6169 (N_6169,N_5529,N_5093);
nand U6170 (N_6170,N_5085,N_5617);
nand U6171 (N_6171,N_4903,N_5885);
and U6172 (N_6172,N_5757,N_5539);
nand U6173 (N_6173,N_5220,N_5646);
nand U6174 (N_6174,N_5670,N_5180);
or U6175 (N_6175,N_5174,N_5224);
xor U6176 (N_6176,N_5702,N_5242);
nand U6177 (N_6177,N_5622,N_5779);
or U6178 (N_6178,N_5135,N_4860);
xor U6179 (N_6179,N_5592,N_4828);
nor U6180 (N_6180,N_5838,N_5781);
nand U6181 (N_6181,N_4807,N_5441);
or U6182 (N_6182,N_5069,N_5407);
xor U6183 (N_6183,N_5958,N_5793);
xnor U6184 (N_6184,N_5689,N_4829);
nand U6185 (N_6185,N_5500,N_5754);
nand U6186 (N_6186,N_5547,N_5907);
nand U6187 (N_6187,N_5018,N_5485);
nor U6188 (N_6188,N_5153,N_5030);
nand U6189 (N_6189,N_4826,N_5333);
and U6190 (N_6190,N_5105,N_5901);
xor U6191 (N_6191,N_5777,N_4984);
nand U6192 (N_6192,N_5713,N_5580);
or U6193 (N_6193,N_5651,N_5610);
and U6194 (N_6194,N_5604,N_5032);
and U6195 (N_6195,N_5043,N_5341);
and U6196 (N_6196,N_4833,N_4979);
or U6197 (N_6197,N_5439,N_4972);
and U6198 (N_6198,N_5292,N_5323);
or U6199 (N_6199,N_5992,N_5421);
or U6200 (N_6200,N_5062,N_5103);
or U6201 (N_6201,N_4946,N_5039);
xnor U6202 (N_6202,N_5661,N_5050);
nand U6203 (N_6203,N_5071,N_5088);
nand U6204 (N_6204,N_5935,N_5107);
nor U6205 (N_6205,N_5917,N_5861);
nor U6206 (N_6206,N_5029,N_5204);
nor U6207 (N_6207,N_5317,N_5131);
and U6208 (N_6208,N_5236,N_5582);
or U6209 (N_6209,N_5411,N_5879);
xnor U6210 (N_6210,N_5332,N_4852);
nor U6211 (N_6211,N_5739,N_5964);
xnor U6212 (N_6212,N_5721,N_5775);
or U6213 (N_6213,N_5521,N_5233);
xor U6214 (N_6214,N_5392,N_5647);
nor U6215 (N_6215,N_5980,N_5549);
nand U6216 (N_6216,N_5245,N_5644);
xor U6217 (N_6217,N_4812,N_4914);
nor U6218 (N_6218,N_5820,N_5904);
nand U6219 (N_6219,N_5656,N_5438);
xnor U6220 (N_6220,N_4891,N_5862);
xor U6221 (N_6221,N_5559,N_5479);
xor U6222 (N_6222,N_5480,N_5923);
nor U6223 (N_6223,N_5822,N_5618);
xnor U6224 (N_6224,N_5440,N_5004);
nand U6225 (N_6225,N_5826,N_5097);
nand U6226 (N_6226,N_5158,N_5451);
nor U6227 (N_6227,N_5183,N_5983);
xnor U6228 (N_6228,N_4840,N_5764);
nand U6229 (N_6229,N_5601,N_5433);
and U6230 (N_6230,N_5491,N_5170);
nand U6231 (N_6231,N_4855,N_5598);
and U6232 (N_6232,N_5051,N_5214);
nor U6233 (N_6233,N_5395,N_5360);
nor U6234 (N_6234,N_5396,N_5939);
or U6235 (N_6235,N_5462,N_5554);
xnor U6236 (N_6236,N_5370,N_4944);
and U6237 (N_6237,N_5046,N_5460);
and U6238 (N_6238,N_5298,N_5712);
nor U6239 (N_6239,N_5009,N_5436);
nor U6240 (N_6240,N_5798,N_5168);
nor U6241 (N_6241,N_5490,N_5524);
nand U6242 (N_6242,N_5077,N_4910);
xnor U6243 (N_6243,N_5803,N_5374);
or U6244 (N_6244,N_5222,N_5931);
xnor U6245 (N_6245,N_4950,N_4988);
or U6246 (N_6246,N_5065,N_5274);
nand U6247 (N_6247,N_5673,N_4814);
or U6248 (N_6248,N_5669,N_4823);
nor U6249 (N_6249,N_5685,N_5938);
or U6250 (N_6250,N_5425,N_5305);
nor U6251 (N_6251,N_5719,N_5997);
nand U6252 (N_6252,N_5201,N_5369);
nand U6253 (N_6253,N_5154,N_4861);
nand U6254 (N_6254,N_5273,N_5017);
xnor U6255 (N_6255,N_5313,N_5734);
nand U6256 (N_6256,N_5859,N_5648);
or U6257 (N_6257,N_4986,N_5680);
nand U6258 (N_6258,N_5593,N_5036);
nand U6259 (N_6259,N_5786,N_5928);
nand U6260 (N_6260,N_4967,N_4992);
nand U6261 (N_6261,N_5890,N_4965);
nand U6262 (N_6262,N_5849,N_5752);
or U6263 (N_6263,N_5607,N_5763);
nor U6264 (N_6264,N_5857,N_5816);
nor U6265 (N_6265,N_5758,N_5991);
and U6266 (N_6266,N_5955,N_5973);
xor U6267 (N_6267,N_5778,N_5927);
xnor U6268 (N_6268,N_4919,N_5762);
xnor U6269 (N_6269,N_5603,N_4839);
or U6270 (N_6270,N_5368,N_5940);
and U6271 (N_6271,N_5302,N_5304);
nor U6272 (N_6272,N_5765,N_5159);
nor U6273 (N_6273,N_5157,N_5241);
and U6274 (N_6274,N_5109,N_5498);
nand U6275 (N_6275,N_5988,N_4960);
nor U6276 (N_6276,N_5504,N_4827);
nor U6277 (N_6277,N_5427,N_4857);
nor U6278 (N_6278,N_5697,N_4896);
nor U6279 (N_6279,N_5723,N_5289);
or U6280 (N_6280,N_5755,N_4892);
nor U6281 (N_6281,N_4925,N_5409);
xor U6282 (N_6282,N_5962,N_5731);
xnor U6283 (N_6283,N_5707,N_5061);
nand U6284 (N_6284,N_5259,N_5275);
xnor U6285 (N_6285,N_5891,N_5600);
nand U6286 (N_6286,N_5037,N_5625);
and U6287 (N_6287,N_5389,N_5921);
nor U6288 (N_6288,N_5710,N_5476);
xor U6289 (N_6289,N_5136,N_5058);
xnor U6290 (N_6290,N_5470,N_5133);
and U6291 (N_6291,N_5074,N_5729);
nand U6292 (N_6292,N_4945,N_4970);
or U6293 (N_6293,N_5246,N_5230);
and U6294 (N_6294,N_4878,N_4917);
and U6295 (N_6295,N_5717,N_5072);
or U6296 (N_6296,N_5815,N_4991);
nor U6297 (N_6297,N_5358,N_5079);
nor U6298 (N_6298,N_5987,N_5014);
xor U6299 (N_6299,N_5020,N_5691);
nor U6300 (N_6300,N_5193,N_5583);
and U6301 (N_6301,N_5749,N_5444);
or U6302 (N_6302,N_5387,N_5215);
xnor U6303 (N_6303,N_5800,N_5457);
nand U6304 (N_6304,N_5101,N_5855);
nor U6305 (N_6305,N_5394,N_5262);
or U6306 (N_6306,N_5481,N_5563);
and U6307 (N_6307,N_5801,N_5546);
or U6308 (N_6308,N_5375,N_5895);
or U6309 (N_6309,N_5199,N_5698);
or U6310 (N_6310,N_5746,N_5296);
or U6311 (N_6311,N_5836,N_5334);
and U6312 (N_6312,N_5108,N_5972);
xnor U6313 (N_6313,N_4949,N_4873);
and U6314 (N_6314,N_5966,N_5474);
nor U6315 (N_6315,N_5376,N_5841);
and U6316 (N_6316,N_5055,N_5340);
nor U6317 (N_6317,N_5310,N_5247);
xor U6318 (N_6318,N_5969,N_4845);
nor U6319 (N_6319,N_5929,N_5488);
nor U6320 (N_6320,N_4875,N_5522);
nand U6321 (N_6321,N_5482,N_5422);
or U6322 (N_6322,N_5688,N_5006);
or U6323 (N_6323,N_5889,N_4831);
and U6324 (N_6324,N_5993,N_5696);
nor U6325 (N_6325,N_5679,N_5591);
nor U6326 (N_6326,N_5019,N_5363);
nand U6327 (N_6327,N_5780,N_5330);
xnor U6328 (N_6328,N_5627,N_5346);
xor U6329 (N_6329,N_5251,N_5381);
and U6330 (N_6330,N_5207,N_4810);
nand U6331 (N_6331,N_5209,N_5837);
or U6332 (N_6332,N_5198,N_4881);
xnor U6333 (N_6333,N_5359,N_5770);
xor U6334 (N_6334,N_5700,N_5315);
nor U6335 (N_6335,N_5833,N_5840);
or U6336 (N_6336,N_5736,N_4893);
nor U6337 (N_6337,N_4815,N_5078);
nand U6338 (N_6338,N_5469,N_5711);
or U6339 (N_6339,N_5948,N_5677);
nand U6340 (N_6340,N_5595,N_5909);
and U6341 (N_6341,N_5788,N_5258);
and U6342 (N_6342,N_4999,N_5846);
and U6343 (N_6343,N_4801,N_5968);
nand U6344 (N_6344,N_5674,N_5965);
or U6345 (N_6345,N_5428,N_5571);
nand U6346 (N_6346,N_5171,N_5120);
and U6347 (N_6347,N_5356,N_5829);
xnor U6348 (N_6348,N_5076,N_5348);
or U6349 (N_6349,N_4994,N_4890);
and U6350 (N_6350,N_4836,N_4907);
xnor U6351 (N_6351,N_5860,N_5839);
and U6352 (N_6352,N_5223,N_5059);
nand U6353 (N_6353,N_5640,N_5663);
xor U6354 (N_6354,N_5570,N_5458);
and U6355 (N_6355,N_5596,N_5944);
and U6356 (N_6356,N_5995,N_5163);
or U6357 (N_6357,N_5878,N_5100);
and U6358 (N_6358,N_5986,N_4913);
and U6359 (N_6359,N_5186,N_5912);
or U6360 (N_6360,N_5690,N_4943);
or U6361 (N_6361,N_5175,N_5942);
nand U6362 (N_6362,N_5807,N_4968);
and U6363 (N_6363,N_5063,N_4822);
xor U6364 (N_6364,N_5021,N_5774);
xnor U6365 (N_6365,N_5981,N_5309);
and U6366 (N_6366,N_4934,N_5517);
nand U6367 (N_6367,N_5865,N_5561);
and U6368 (N_6368,N_4951,N_5047);
or U6369 (N_6369,N_4862,N_5331);
xor U6370 (N_6370,N_5187,N_5250);
nor U6371 (N_6371,N_4985,N_5937);
and U6372 (N_6372,N_5519,N_4948);
and U6373 (N_6373,N_5577,N_5464);
nand U6374 (N_6374,N_5709,N_5146);
nor U6375 (N_6375,N_5877,N_4952);
nor U6376 (N_6376,N_5134,N_5318);
or U6377 (N_6377,N_5666,N_4830);
and U6378 (N_6378,N_5178,N_5497);
xor U6379 (N_6379,N_4838,N_4909);
and U6380 (N_6380,N_5665,N_5714);
nand U6381 (N_6381,N_5414,N_5372);
nor U6382 (N_6382,N_5835,N_5615);
nor U6383 (N_6383,N_5286,N_5585);
or U6384 (N_6384,N_5400,N_5636);
nand U6385 (N_6385,N_5445,N_5373);
nor U6386 (N_6386,N_5182,N_5091);
or U6387 (N_6387,N_4864,N_5196);
or U6388 (N_6388,N_5867,N_5667);
or U6389 (N_6389,N_5484,N_4966);
nor U6390 (N_6390,N_5659,N_5785);
or U6391 (N_6391,N_5412,N_5454);
or U6392 (N_6392,N_5325,N_5507);
nor U6393 (N_6393,N_5234,N_5613);
nor U6394 (N_6394,N_5568,N_5288);
xor U6395 (N_6395,N_5383,N_5657);
and U6396 (N_6396,N_5794,N_4942);
or U6397 (N_6397,N_5722,N_4898);
xnor U6398 (N_6398,N_5513,N_5377);
or U6399 (N_6399,N_5053,N_5113);
nand U6400 (N_6400,N_5260,N_5102);
or U6401 (N_6401,N_5531,N_5112);
nand U6402 (N_6402,N_5321,N_5005);
xnor U6403 (N_6403,N_4964,N_5827);
and U6404 (N_6404,N_5511,N_5437);
or U6405 (N_6405,N_5573,N_5994);
xnor U6406 (N_6406,N_4850,N_5868);
xor U6407 (N_6407,N_5417,N_5353);
or U6408 (N_6408,N_5893,N_5189);
nor U6409 (N_6409,N_5277,N_5672);
xor U6410 (N_6410,N_4883,N_5916);
or U6411 (N_6411,N_4940,N_5056);
xor U6412 (N_6412,N_5064,N_5211);
xor U6413 (N_6413,N_5371,N_5532);
nor U6414 (N_6414,N_5130,N_4854);
xor U6415 (N_6415,N_5520,N_4911);
or U6416 (N_6416,N_5905,N_5034);
or U6417 (N_6417,N_5284,N_5985);
and U6418 (N_6418,N_5361,N_5537);
nor U6419 (N_6419,N_5525,N_5543);
and U6420 (N_6420,N_5467,N_5338);
or U6421 (N_6421,N_4871,N_5896);
or U6422 (N_6422,N_5326,N_4937);
and U6423 (N_6423,N_5843,N_5784);
nor U6424 (N_6424,N_5813,N_5280);
nand U6425 (N_6425,N_4897,N_5587);
or U6426 (N_6426,N_5588,N_5379);
nor U6427 (N_6427,N_5894,N_5430);
and U6428 (N_6428,N_5924,N_5967);
xor U6429 (N_6429,N_5461,N_4803);
nand U6430 (N_6430,N_5686,N_5205);
or U6431 (N_6431,N_5416,N_5082);
nand U6432 (N_6432,N_4983,N_5791);
and U6433 (N_6433,N_5041,N_5087);
or U6434 (N_6434,N_5473,N_5898);
nor U6435 (N_6435,N_5523,N_4889);
or U6436 (N_6436,N_5477,N_5953);
or U6437 (N_6437,N_5096,N_5506);
nor U6438 (N_6438,N_5294,N_5140);
or U6439 (N_6439,N_5502,N_4961);
nand U6440 (N_6440,N_4809,N_5402);
or U6441 (N_6441,N_5558,N_4863);
and U6442 (N_6442,N_5650,N_4819);
xor U6443 (N_6443,N_5668,N_4843);
xor U6444 (N_6444,N_4926,N_5544);
xor U6445 (N_6445,N_4842,N_5202);
xor U6446 (N_6446,N_5031,N_5681);
or U6447 (N_6447,N_4912,N_5162);
and U6448 (N_6448,N_5388,N_5408);
or U6449 (N_6449,N_5044,N_5854);
and U6450 (N_6450,N_4874,N_5556);
nand U6451 (N_6451,N_5609,N_5179);
and U6452 (N_6452,N_4924,N_5297);
and U6453 (N_6453,N_4962,N_5465);
or U6454 (N_6454,N_5448,N_5329);
nand U6455 (N_6455,N_5925,N_5638);
xor U6456 (N_6456,N_4884,N_5887);
nor U6457 (N_6457,N_4954,N_5602);
nand U6458 (N_6458,N_5810,N_5128);
and U6459 (N_6459,N_4973,N_5429);
xor U6460 (N_6460,N_5947,N_5984);
and U6461 (N_6461,N_5415,N_5705);
or U6462 (N_6462,N_5463,N_5693);
or U6463 (N_6463,N_5886,N_5132);
xor U6464 (N_6464,N_5756,N_5872);
or U6465 (N_6465,N_5527,N_5922);
and U6466 (N_6466,N_4963,N_5282);
and U6467 (N_6467,N_5468,N_5936);
nor U6468 (N_6468,N_4886,N_5526);
nor U6469 (N_6469,N_5092,N_5628);
xor U6470 (N_6470,N_5821,N_5851);
and U6471 (N_6471,N_4918,N_5708);
xnor U6472 (N_6472,N_5350,N_5141);
and U6473 (N_6473,N_5145,N_5880);
or U6474 (N_6474,N_5594,N_4816);
xor U6475 (N_6475,N_5010,N_5637);
nor U6476 (N_6476,N_5687,N_5378);
or U6477 (N_6477,N_4805,N_5856);
and U6478 (N_6478,N_5466,N_5118);
nand U6479 (N_6479,N_5291,N_4882);
or U6480 (N_6480,N_5122,N_5726);
xnor U6481 (N_6481,N_5080,N_5503);
xnor U6482 (N_6482,N_4872,N_5683);
xor U6483 (N_6483,N_5099,N_5960);
and U6484 (N_6484,N_5982,N_5256);
nor U6485 (N_6485,N_5597,N_5823);
and U6486 (N_6486,N_5478,N_5847);
or U6487 (N_6487,N_5505,N_5493);
and U6488 (N_6488,N_4821,N_4853);
nor U6489 (N_6489,N_5161,N_5040);
or U6490 (N_6490,N_5125,N_5287);
xnor U6491 (N_6491,N_5941,N_5083);
xor U6492 (N_6492,N_5730,N_5308);
nor U6493 (N_6493,N_5951,N_5252);
nand U6494 (N_6494,N_5630,N_4975);
xor U6495 (N_6495,N_5152,N_5900);
xnor U6496 (N_6496,N_5782,N_5552);
xor U6497 (N_6497,N_5853,N_5494);
nand U6498 (N_6498,N_5945,N_4987);
nand U6499 (N_6499,N_4990,N_5560);
nor U6500 (N_6500,N_5876,N_5926);
or U6501 (N_6501,N_5975,N_4922);
xor U6502 (N_6502,N_5475,N_5094);
or U6503 (N_6503,N_5235,N_5254);
and U6504 (N_6504,N_5575,N_4846);
and U6505 (N_6505,N_5472,N_5789);
or U6506 (N_6506,N_5397,N_5471);
nor U6507 (N_6507,N_5450,N_5257);
nor U6508 (N_6508,N_4993,N_4835);
and U6509 (N_6509,N_5442,N_5911);
nor U6510 (N_6510,N_5265,N_5268);
xnor U6511 (N_6511,N_5151,N_5728);
and U6512 (N_6512,N_5514,N_5512);
and U6513 (N_6513,N_5144,N_5624);
or U6514 (N_6514,N_5195,N_4920);
or U6515 (N_6515,N_5424,N_5227);
xnor U6516 (N_6516,N_5142,N_5564);
nand U6517 (N_6517,N_5567,N_5312);
or U6518 (N_6518,N_5946,N_4957);
nor U6519 (N_6519,N_5165,N_5956);
xnor U6520 (N_6520,N_5824,N_5881);
and U6521 (N_6521,N_5049,N_5773);
or U6522 (N_6522,N_5733,N_5495);
nor U6523 (N_6523,N_5933,N_4800);
xnor U6524 (N_6524,N_5016,N_4879);
nor U6525 (N_6525,N_5367,N_5301);
nand U6526 (N_6526,N_5743,N_5753);
nand U6527 (N_6527,N_5200,N_5033);
and U6528 (N_6528,N_5181,N_5518);
xor U6529 (N_6529,N_4978,N_5218);
or U6530 (N_6530,N_5908,N_5060);
nand U6531 (N_6531,N_5380,N_5635);
xor U6532 (N_6532,N_5501,N_5619);
nand U6533 (N_6533,N_5715,N_5404);
nor U6534 (N_6534,N_5320,N_5070);
and U6535 (N_6535,N_5852,N_4939);
xor U6536 (N_6536,N_5676,N_5599);
nand U6537 (N_6537,N_4981,N_5197);
xor U6538 (N_6538,N_5007,N_5054);
nor U6539 (N_6539,N_5418,N_5932);
or U6540 (N_6540,N_5176,N_5653);
nor U6541 (N_6541,N_5432,N_5486);
or U6542 (N_6542,N_5787,N_5114);
or U6543 (N_6543,N_5873,N_5155);
xor U6544 (N_6544,N_4905,N_5508);
xnor U6545 (N_6545,N_5874,N_4977);
xor U6546 (N_6546,N_4866,N_4980);
xnor U6547 (N_6547,N_4941,N_5550);
and U6548 (N_6548,N_5766,N_5825);
or U6549 (N_6549,N_5957,N_5623);
nor U6550 (N_6550,N_5327,N_5553);
and U6551 (N_6551,N_5249,N_4932);
and U6552 (N_6552,N_5221,N_4915);
or U6553 (N_6553,N_5012,N_5954);
nand U6554 (N_6554,N_4930,N_5510);
or U6555 (N_6555,N_5382,N_5138);
and U6556 (N_6556,N_5639,N_5026);
and U6557 (N_6557,N_5203,N_5357);
xor U6558 (N_6558,N_5649,N_4870);
nand U6559 (N_6559,N_5819,N_5206);
xnor U6560 (N_6560,N_5978,N_5842);
xnor U6561 (N_6561,N_5067,N_5660);
or U6562 (N_6562,N_5237,N_4902);
nor U6563 (N_6563,N_5706,N_4825);
or U6564 (N_6564,N_5538,N_5352);
and U6565 (N_6565,N_5084,N_5279);
nand U6566 (N_6566,N_5509,N_5139);
or U6567 (N_6567,N_5751,N_5551);
nor U6568 (N_6568,N_5399,N_5231);
and U6569 (N_6569,N_5684,N_5166);
and U6570 (N_6570,N_5664,N_5963);
or U6571 (N_6571,N_5217,N_5172);
and U6572 (N_6572,N_5124,N_4996);
nor U6573 (N_6573,N_5106,N_5423);
nand U6574 (N_6574,N_5447,N_5219);
xor U6575 (N_6575,N_5190,N_5148);
xnor U6576 (N_6576,N_4936,N_5015);
xnor U6577 (N_6577,N_5240,N_5149);
or U6578 (N_6578,N_4923,N_5633);
nor U6579 (N_6579,N_5073,N_5977);
nand U6580 (N_6580,N_5814,N_5806);
xnor U6581 (N_6581,N_4849,N_5095);
and U6582 (N_6582,N_5336,N_5850);
or U6583 (N_6583,N_5355,N_4995);
nor U6584 (N_6584,N_4876,N_5110);
nor U6585 (N_6585,N_5391,N_5727);
xor U6586 (N_6586,N_5732,N_5614);
and U6587 (N_6587,N_5238,N_5771);
nor U6588 (N_6588,N_5164,N_5270);
nand U6589 (N_6589,N_5634,N_4933);
nor U6590 (N_6590,N_5671,N_5863);
and U6591 (N_6591,N_5000,N_5990);
and U6592 (N_6592,N_5328,N_5533);
or U6593 (N_6593,N_5048,N_4808);
xnor U6594 (N_6594,N_5483,N_4818);
nand U6595 (N_6595,N_5804,N_5632);
xnor U6596 (N_6596,N_5365,N_5239);
nor U6597 (N_6597,N_5748,N_5413);
and U6598 (N_6598,N_5403,N_5276);
and U6599 (N_6599,N_5194,N_5499);
nor U6600 (N_6600,N_4854,N_5732);
nand U6601 (N_6601,N_4840,N_4870);
nand U6602 (N_6602,N_5074,N_5009);
nand U6603 (N_6603,N_5012,N_5720);
nand U6604 (N_6604,N_5192,N_5697);
nor U6605 (N_6605,N_5627,N_4946);
or U6606 (N_6606,N_5939,N_5427);
nand U6607 (N_6607,N_5633,N_5747);
and U6608 (N_6608,N_5529,N_5858);
nor U6609 (N_6609,N_5409,N_5669);
nor U6610 (N_6610,N_5097,N_5437);
xor U6611 (N_6611,N_4829,N_5070);
or U6612 (N_6612,N_5094,N_5551);
xor U6613 (N_6613,N_5909,N_5346);
or U6614 (N_6614,N_5714,N_5076);
and U6615 (N_6615,N_5579,N_5998);
or U6616 (N_6616,N_5939,N_5730);
xnor U6617 (N_6617,N_5416,N_5247);
or U6618 (N_6618,N_5837,N_5502);
xor U6619 (N_6619,N_5041,N_5560);
nor U6620 (N_6620,N_5002,N_5160);
and U6621 (N_6621,N_4932,N_5653);
nand U6622 (N_6622,N_5862,N_5753);
nor U6623 (N_6623,N_4876,N_5670);
xnor U6624 (N_6624,N_5231,N_5107);
and U6625 (N_6625,N_5820,N_5149);
and U6626 (N_6626,N_5936,N_5265);
nand U6627 (N_6627,N_5263,N_4809);
nor U6628 (N_6628,N_5156,N_5870);
and U6629 (N_6629,N_5598,N_5760);
xnor U6630 (N_6630,N_5489,N_5433);
and U6631 (N_6631,N_5647,N_5200);
xor U6632 (N_6632,N_4996,N_5232);
and U6633 (N_6633,N_5316,N_5375);
and U6634 (N_6634,N_5915,N_5977);
nor U6635 (N_6635,N_5578,N_5155);
xnor U6636 (N_6636,N_5716,N_4808);
xnor U6637 (N_6637,N_5884,N_5078);
and U6638 (N_6638,N_4896,N_5945);
and U6639 (N_6639,N_4814,N_5434);
nand U6640 (N_6640,N_4822,N_5789);
nor U6641 (N_6641,N_5853,N_5093);
nor U6642 (N_6642,N_5344,N_5908);
nand U6643 (N_6643,N_5570,N_4933);
nand U6644 (N_6644,N_5826,N_4933);
nor U6645 (N_6645,N_4993,N_5427);
or U6646 (N_6646,N_5234,N_5495);
nor U6647 (N_6647,N_4841,N_5029);
or U6648 (N_6648,N_5957,N_5757);
nand U6649 (N_6649,N_5349,N_5501);
xnor U6650 (N_6650,N_5064,N_5200);
and U6651 (N_6651,N_5035,N_5562);
xor U6652 (N_6652,N_5431,N_5396);
or U6653 (N_6653,N_4893,N_5830);
or U6654 (N_6654,N_5433,N_5157);
nor U6655 (N_6655,N_5266,N_5077);
or U6656 (N_6656,N_5962,N_5258);
xnor U6657 (N_6657,N_5198,N_5200);
nand U6658 (N_6658,N_5218,N_5909);
nor U6659 (N_6659,N_5809,N_5588);
or U6660 (N_6660,N_5226,N_5727);
or U6661 (N_6661,N_4824,N_5870);
or U6662 (N_6662,N_4967,N_5055);
or U6663 (N_6663,N_5657,N_5742);
nor U6664 (N_6664,N_5903,N_5989);
or U6665 (N_6665,N_5805,N_5989);
and U6666 (N_6666,N_5694,N_5648);
xnor U6667 (N_6667,N_5041,N_5144);
or U6668 (N_6668,N_5534,N_5566);
nand U6669 (N_6669,N_5155,N_5497);
nand U6670 (N_6670,N_5583,N_5027);
xor U6671 (N_6671,N_4967,N_5205);
nand U6672 (N_6672,N_5995,N_4928);
nand U6673 (N_6673,N_5158,N_5733);
or U6674 (N_6674,N_5212,N_5050);
nor U6675 (N_6675,N_5692,N_4902);
or U6676 (N_6676,N_4996,N_5893);
nor U6677 (N_6677,N_5315,N_5348);
and U6678 (N_6678,N_5819,N_5601);
nor U6679 (N_6679,N_5339,N_5611);
and U6680 (N_6680,N_5323,N_5441);
and U6681 (N_6681,N_5581,N_5357);
and U6682 (N_6682,N_5386,N_4980);
or U6683 (N_6683,N_5518,N_5304);
nor U6684 (N_6684,N_4893,N_5221);
or U6685 (N_6685,N_5999,N_4845);
nand U6686 (N_6686,N_5222,N_4990);
nand U6687 (N_6687,N_5200,N_5766);
and U6688 (N_6688,N_5535,N_5633);
and U6689 (N_6689,N_5214,N_4864);
and U6690 (N_6690,N_5272,N_5916);
and U6691 (N_6691,N_5314,N_4962);
or U6692 (N_6692,N_5764,N_5280);
nor U6693 (N_6693,N_5841,N_5136);
nand U6694 (N_6694,N_4898,N_5181);
nand U6695 (N_6695,N_4840,N_5892);
xnor U6696 (N_6696,N_5585,N_4805);
nor U6697 (N_6697,N_4914,N_5236);
nor U6698 (N_6698,N_4984,N_5373);
nand U6699 (N_6699,N_5127,N_5222);
nand U6700 (N_6700,N_5448,N_5767);
nand U6701 (N_6701,N_5606,N_5062);
and U6702 (N_6702,N_5375,N_4893);
xor U6703 (N_6703,N_4899,N_5144);
nor U6704 (N_6704,N_5655,N_5546);
and U6705 (N_6705,N_4952,N_5135);
xor U6706 (N_6706,N_4924,N_5825);
or U6707 (N_6707,N_5178,N_5524);
nor U6708 (N_6708,N_5037,N_5477);
nor U6709 (N_6709,N_5823,N_5425);
xor U6710 (N_6710,N_5668,N_5861);
and U6711 (N_6711,N_5937,N_4850);
and U6712 (N_6712,N_5631,N_5927);
and U6713 (N_6713,N_5733,N_5182);
or U6714 (N_6714,N_4967,N_5910);
and U6715 (N_6715,N_5805,N_5280);
xnor U6716 (N_6716,N_5761,N_5167);
nand U6717 (N_6717,N_5642,N_4940);
or U6718 (N_6718,N_5964,N_5026);
xnor U6719 (N_6719,N_4880,N_5843);
nor U6720 (N_6720,N_5153,N_5426);
and U6721 (N_6721,N_5014,N_5631);
and U6722 (N_6722,N_5967,N_5084);
or U6723 (N_6723,N_4963,N_5250);
and U6724 (N_6724,N_5905,N_5980);
nand U6725 (N_6725,N_5078,N_5532);
nand U6726 (N_6726,N_4912,N_5033);
nand U6727 (N_6727,N_4878,N_5723);
nor U6728 (N_6728,N_5503,N_5734);
nor U6729 (N_6729,N_4952,N_5126);
nand U6730 (N_6730,N_5378,N_5515);
nand U6731 (N_6731,N_4965,N_5518);
and U6732 (N_6732,N_5869,N_5630);
nand U6733 (N_6733,N_5726,N_5431);
or U6734 (N_6734,N_5806,N_5444);
and U6735 (N_6735,N_5440,N_5056);
or U6736 (N_6736,N_5689,N_5951);
nand U6737 (N_6737,N_4825,N_4849);
xor U6738 (N_6738,N_5480,N_5004);
or U6739 (N_6739,N_5575,N_5659);
or U6740 (N_6740,N_5045,N_5524);
xnor U6741 (N_6741,N_5852,N_5575);
nor U6742 (N_6742,N_5920,N_5980);
and U6743 (N_6743,N_5396,N_5932);
and U6744 (N_6744,N_4896,N_5622);
nand U6745 (N_6745,N_5929,N_4959);
nor U6746 (N_6746,N_5096,N_5614);
nor U6747 (N_6747,N_5932,N_5411);
xor U6748 (N_6748,N_5412,N_5880);
or U6749 (N_6749,N_4946,N_5010);
and U6750 (N_6750,N_5886,N_5202);
xnor U6751 (N_6751,N_4956,N_5320);
and U6752 (N_6752,N_5939,N_5824);
nand U6753 (N_6753,N_4835,N_5507);
xnor U6754 (N_6754,N_4861,N_4873);
xnor U6755 (N_6755,N_5395,N_5652);
nor U6756 (N_6756,N_5548,N_5144);
or U6757 (N_6757,N_5270,N_5601);
and U6758 (N_6758,N_4947,N_5669);
and U6759 (N_6759,N_5884,N_4970);
nand U6760 (N_6760,N_5842,N_5043);
xor U6761 (N_6761,N_5051,N_5128);
xnor U6762 (N_6762,N_5443,N_5915);
xnor U6763 (N_6763,N_5982,N_5770);
or U6764 (N_6764,N_5231,N_5009);
and U6765 (N_6765,N_5010,N_5476);
xor U6766 (N_6766,N_5956,N_5755);
nor U6767 (N_6767,N_4897,N_5571);
nor U6768 (N_6768,N_5577,N_4885);
nor U6769 (N_6769,N_5299,N_5534);
nor U6770 (N_6770,N_4996,N_5033);
nor U6771 (N_6771,N_4956,N_5502);
nor U6772 (N_6772,N_4993,N_5223);
nand U6773 (N_6773,N_5283,N_5634);
nor U6774 (N_6774,N_5758,N_5036);
and U6775 (N_6775,N_4833,N_5760);
or U6776 (N_6776,N_5495,N_5642);
xnor U6777 (N_6777,N_5366,N_4801);
or U6778 (N_6778,N_5817,N_5836);
or U6779 (N_6779,N_5914,N_5577);
nor U6780 (N_6780,N_5373,N_5497);
and U6781 (N_6781,N_5849,N_5537);
or U6782 (N_6782,N_5773,N_5162);
nor U6783 (N_6783,N_5977,N_5371);
or U6784 (N_6784,N_5835,N_4992);
nand U6785 (N_6785,N_4902,N_5751);
and U6786 (N_6786,N_5312,N_4982);
xnor U6787 (N_6787,N_5698,N_5137);
nor U6788 (N_6788,N_5386,N_4992);
nand U6789 (N_6789,N_5057,N_5795);
xor U6790 (N_6790,N_5530,N_5287);
nand U6791 (N_6791,N_5732,N_5547);
xor U6792 (N_6792,N_5632,N_5398);
nand U6793 (N_6793,N_5517,N_5430);
or U6794 (N_6794,N_4881,N_5316);
or U6795 (N_6795,N_4907,N_5137);
xor U6796 (N_6796,N_5077,N_5067);
nor U6797 (N_6797,N_5669,N_5718);
nor U6798 (N_6798,N_5342,N_5639);
or U6799 (N_6799,N_5011,N_5035);
or U6800 (N_6800,N_5896,N_5701);
and U6801 (N_6801,N_5329,N_4906);
nor U6802 (N_6802,N_5052,N_5235);
nor U6803 (N_6803,N_5279,N_5581);
xnor U6804 (N_6804,N_5627,N_5757);
nor U6805 (N_6805,N_5183,N_5520);
and U6806 (N_6806,N_5744,N_5498);
and U6807 (N_6807,N_5055,N_5343);
nor U6808 (N_6808,N_5351,N_5437);
nand U6809 (N_6809,N_5956,N_5725);
or U6810 (N_6810,N_5201,N_5807);
or U6811 (N_6811,N_5657,N_5994);
or U6812 (N_6812,N_5271,N_5632);
nor U6813 (N_6813,N_5158,N_5995);
nand U6814 (N_6814,N_5366,N_4888);
nor U6815 (N_6815,N_5993,N_5152);
nand U6816 (N_6816,N_5954,N_5648);
and U6817 (N_6817,N_5378,N_5287);
or U6818 (N_6818,N_5703,N_5511);
xor U6819 (N_6819,N_5680,N_5433);
and U6820 (N_6820,N_5834,N_5432);
nor U6821 (N_6821,N_5479,N_5590);
nand U6822 (N_6822,N_5325,N_5656);
xor U6823 (N_6823,N_4983,N_4813);
or U6824 (N_6824,N_5084,N_5077);
nand U6825 (N_6825,N_5894,N_5474);
and U6826 (N_6826,N_5353,N_5107);
and U6827 (N_6827,N_4885,N_4946);
and U6828 (N_6828,N_4826,N_4940);
or U6829 (N_6829,N_4939,N_5229);
nand U6830 (N_6830,N_5093,N_5648);
nand U6831 (N_6831,N_5935,N_5581);
xnor U6832 (N_6832,N_5475,N_5232);
xnor U6833 (N_6833,N_5817,N_5971);
nor U6834 (N_6834,N_5372,N_5145);
xor U6835 (N_6835,N_4889,N_5103);
nor U6836 (N_6836,N_5999,N_5447);
and U6837 (N_6837,N_5328,N_5297);
or U6838 (N_6838,N_5846,N_5214);
nand U6839 (N_6839,N_5307,N_5999);
xnor U6840 (N_6840,N_5399,N_5533);
nand U6841 (N_6841,N_5953,N_5175);
or U6842 (N_6842,N_4895,N_5751);
nand U6843 (N_6843,N_5398,N_5350);
nor U6844 (N_6844,N_4822,N_4908);
and U6845 (N_6845,N_5690,N_5370);
xnor U6846 (N_6846,N_5489,N_5284);
nor U6847 (N_6847,N_4901,N_5829);
and U6848 (N_6848,N_4866,N_5430);
or U6849 (N_6849,N_4967,N_5801);
nand U6850 (N_6850,N_5245,N_5069);
or U6851 (N_6851,N_5732,N_5313);
or U6852 (N_6852,N_5904,N_5751);
or U6853 (N_6853,N_5915,N_5517);
xnor U6854 (N_6854,N_4810,N_5423);
or U6855 (N_6855,N_5652,N_5379);
or U6856 (N_6856,N_5429,N_4915);
nor U6857 (N_6857,N_5389,N_5228);
and U6858 (N_6858,N_5773,N_4943);
nand U6859 (N_6859,N_5258,N_5544);
and U6860 (N_6860,N_5861,N_5478);
nor U6861 (N_6861,N_5016,N_5565);
and U6862 (N_6862,N_5028,N_5620);
nand U6863 (N_6863,N_5649,N_4940);
nand U6864 (N_6864,N_5199,N_5172);
nand U6865 (N_6865,N_5642,N_5313);
xor U6866 (N_6866,N_5051,N_5527);
xnor U6867 (N_6867,N_5214,N_5107);
xor U6868 (N_6868,N_5831,N_5242);
nand U6869 (N_6869,N_5541,N_5914);
or U6870 (N_6870,N_5437,N_5084);
xor U6871 (N_6871,N_5252,N_5780);
or U6872 (N_6872,N_5039,N_5842);
nor U6873 (N_6873,N_5087,N_5030);
and U6874 (N_6874,N_4824,N_5816);
nand U6875 (N_6875,N_5296,N_4947);
xor U6876 (N_6876,N_5126,N_5663);
xnor U6877 (N_6877,N_5871,N_5576);
xor U6878 (N_6878,N_5584,N_5415);
and U6879 (N_6879,N_5896,N_5717);
nor U6880 (N_6880,N_4843,N_5030);
or U6881 (N_6881,N_5158,N_5588);
nor U6882 (N_6882,N_5293,N_5995);
xor U6883 (N_6883,N_5254,N_5409);
nor U6884 (N_6884,N_5789,N_5865);
or U6885 (N_6885,N_5990,N_5980);
and U6886 (N_6886,N_5891,N_5059);
and U6887 (N_6887,N_5210,N_5265);
nand U6888 (N_6888,N_4891,N_5348);
or U6889 (N_6889,N_5864,N_5308);
xor U6890 (N_6890,N_4955,N_5723);
and U6891 (N_6891,N_5940,N_5475);
nor U6892 (N_6892,N_5676,N_5969);
nor U6893 (N_6893,N_5808,N_5221);
nor U6894 (N_6894,N_5347,N_5670);
nor U6895 (N_6895,N_5176,N_5705);
or U6896 (N_6896,N_5193,N_5763);
and U6897 (N_6897,N_5154,N_5253);
nand U6898 (N_6898,N_4950,N_5333);
xor U6899 (N_6899,N_5344,N_4848);
nand U6900 (N_6900,N_5462,N_5534);
or U6901 (N_6901,N_4846,N_5686);
nand U6902 (N_6902,N_5158,N_5040);
and U6903 (N_6903,N_5478,N_4874);
xnor U6904 (N_6904,N_5697,N_5949);
xor U6905 (N_6905,N_5531,N_5129);
or U6906 (N_6906,N_5065,N_5880);
nand U6907 (N_6907,N_4980,N_5236);
and U6908 (N_6908,N_5395,N_4886);
xnor U6909 (N_6909,N_5002,N_5397);
nand U6910 (N_6910,N_4966,N_5931);
nand U6911 (N_6911,N_4973,N_5900);
nand U6912 (N_6912,N_5478,N_5326);
nor U6913 (N_6913,N_5315,N_4937);
xnor U6914 (N_6914,N_5257,N_5479);
and U6915 (N_6915,N_5714,N_5145);
or U6916 (N_6916,N_4825,N_5604);
or U6917 (N_6917,N_5635,N_4932);
xnor U6918 (N_6918,N_5807,N_5868);
or U6919 (N_6919,N_5906,N_5072);
nand U6920 (N_6920,N_5615,N_5945);
nand U6921 (N_6921,N_5372,N_5079);
or U6922 (N_6922,N_5177,N_5232);
nand U6923 (N_6923,N_5305,N_5499);
nor U6924 (N_6924,N_5517,N_5937);
and U6925 (N_6925,N_4989,N_5067);
xor U6926 (N_6926,N_5509,N_5860);
nor U6927 (N_6927,N_4932,N_5584);
and U6928 (N_6928,N_5733,N_5917);
nand U6929 (N_6929,N_5568,N_5551);
or U6930 (N_6930,N_5634,N_5818);
nor U6931 (N_6931,N_5553,N_5339);
nand U6932 (N_6932,N_5381,N_5207);
or U6933 (N_6933,N_5199,N_4866);
or U6934 (N_6934,N_5208,N_5733);
or U6935 (N_6935,N_5058,N_5218);
and U6936 (N_6936,N_4905,N_5540);
xor U6937 (N_6937,N_4988,N_5414);
nor U6938 (N_6938,N_4879,N_5189);
xnor U6939 (N_6939,N_5875,N_5207);
and U6940 (N_6940,N_5572,N_5728);
and U6941 (N_6941,N_5405,N_4901);
nand U6942 (N_6942,N_5194,N_5067);
and U6943 (N_6943,N_5617,N_5780);
nand U6944 (N_6944,N_5687,N_4823);
nor U6945 (N_6945,N_5484,N_5320);
nor U6946 (N_6946,N_4807,N_5518);
nor U6947 (N_6947,N_5893,N_5684);
nand U6948 (N_6948,N_5252,N_5461);
nand U6949 (N_6949,N_5989,N_5274);
nand U6950 (N_6950,N_5420,N_5823);
xnor U6951 (N_6951,N_5295,N_5550);
xnor U6952 (N_6952,N_4940,N_5112);
nand U6953 (N_6953,N_5109,N_5644);
nor U6954 (N_6954,N_5559,N_5779);
nand U6955 (N_6955,N_4899,N_5508);
nand U6956 (N_6956,N_4961,N_5440);
nor U6957 (N_6957,N_5026,N_5515);
nor U6958 (N_6958,N_4887,N_5799);
or U6959 (N_6959,N_4897,N_5263);
xnor U6960 (N_6960,N_4882,N_5210);
and U6961 (N_6961,N_5067,N_5899);
xnor U6962 (N_6962,N_5839,N_4995);
or U6963 (N_6963,N_5451,N_5173);
nor U6964 (N_6964,N_5899,N_4931);
or U6965 (N_6965,N_4880,N_5299);
nor U6966 (N_6966,N_5473,N_5409);
xor U6967 (N_6967,N_5259,N_5946);
nand U6968 (N_6968,N_5054,N_5827);
nand U6969 (N_6969,N_5435,N_5786);
xor U6970 (N_6970,N_4817,N_5856);
nor U6971 (N_6971,N_5903,N_5474);
nand U6972 (N_6972,N_5917,N_5047);
nor U6973 (N_6973,N_5945,N_5214);
and U6974 (N_6974,N_5867,N_5330);
or U6975 (N_6975,N_5125,N_5346);
and U6976 (N_6976,N_5668,N_5680);
nor U6977 (N_6977,N_5295,N_5331);
nand U6978 (N_6978,N_5442,N_5551);
or U6979 (N_6979,N_5145,N_5678);
nor U6980 (N_6980,N_4835,N_5962);
xor U6981 (N_6981,N_5762,N_5712);
nor U6982 (N_6982,N_5324,N_5024);
and U6983 (N_6983,N_5346,N_5107);
nand U6984 (N_6984,N_5871,N_5853);
nor U6985 (N_6985,N_4935,N_5286);
and U6986 (N_6986,N_5960,N_5401);
and U6987 (N_6987,N_5440,N_5288);
nor U6988 (N_6988,N_5124,N_4855);
xnor U6989 (N_6989,N_5470,N_5024);
nand U6990 (N_6990,N_5432,N_5981);
nand U6991 (N_6991,N_5622,N_4960);
xor U6992 (N_6992,N_5956,N_5671);
xor U6993 (N_6993,N_5300,N_5514);
xnor U6994 (N_6994,N_5317,N_5542);
and U6995 (N_6995,N_4989,N_5752);
and U6996 (N_6996,N_5559,N_5308);
and U6997 (N_6997,N_5623,N_5776);
and U6998 (N_6998,N_5942,N_5933);
and U6999 (N_6999,N_5685,N_5185);
xnor U7000 (N_7000,N_5557,N_5484);
or U7001 (N_7001,N_5238,N_5463);
and U7002 (N_7002,N_5792,N_5464);
nor U7003 (N_7003,N_5858,N_5789);
and U7004 (N_7004,N_4942,N_4867);
or U7005 (N_7005,N_5173,N_5213);
and U7006 (N_7006,N_5051,N_5004);
nor U7007 (N_7007,N_5072,N_5918);
and U7008 (N_7008,N_5409,N_4927);
nand U7009 (N_7009,N_5121,N_5124);
or U7010 (N_7010,N_5694,N_5309);
nand U7011 (N_7011,N_5350,N_5828);
and U7012 (N_7012,N_5620,N_5148);
nor U7013 (N_7013,N_4955,N_5542);
nor U7014 (N_7014,N_5022,N_5279);
nor U7015 (N_7015,N_5546,N_5489);
and U7016 (N_7016,N_5891,N_5408);
and U7017 (N_7017,N_5056,N_5684);
nand U7018 (N_7018,N_5471,N_5900);
and U7019 (N_7019,N_5820,N_5893);
or U7020 (N_7020,N_5819,N_5397);
nor U7021 (N_7021,N_4919,N_5808);
nand U7022 (N_7022,N_5218,N_5513);
nand U7023 (N_7023,N_5273,N_5617);
or U7024 (N_7024,N_5469,N_5328);
nor U7025 (N_7025,N_5687,N_4800);
nor U7026 (N_7026,N_5489,N_5455);
nor U7027 (N_7027,N_5042,N_5047);
xnor U7028 (N_7028,N_5155,N_5422);
or U7029 (N_7029,N_5596,N_5860);
nor U7030 (N_7030,N_5860,N_5311);
or U7031 (N_7031,N_5285,N_5245);
and U7032 (N_7032,N_5816,N_5688);
and U7033 (N_7033,N_4946,N_5841);
xor U7034 (N_7034,N_5314,N_5348);
and U7035 (N_7035,N_5027,N_5360);
nor U7036 (N_7036,N_5622,N_5512);
or U7037 (N_7037,N_5564,N_5754);
and U7038 (N_7038,N_5661,N_4990);
nand U7039 (N_7039,N_4818,N_5302);
xnor U7040 (N_7040,N_5443,N_5776);
xnor U7041 (N_7041,N_5870,N_4821);
or U7042 (N_7042,N_5411,N_4912);
xnor U7043 (N_7043,N_5998,N_5260);
or U7044 (N_7044,N_5365,N_4899);
xor U7045 (N_7045,N_5879,N_5590);
nand U7046 (N_7046,N_4886,N_5843);
nor U7047 (N_7047,N_5763,N_5468);
or U7048 (N_7048,N_4878,N_5093);
or U7049 (N_7049,N_5922,N_5004);
or U7050 (N_7050,N_5179,N_5680);
nor U7051 (N_7051,N_5798,N_5628);
or U7052 (N_7052,N_5748,N_4928);
or U7053 (N_7053,N_4932,N_5411);
xor U7054 (N_7054,N_5681,N_5880);
or U7055 (N_7055,N_5980,N_5013);
or U7056 (N_7056,N_4882,N_5886);
nor U7057 (N_7057,N_5735,N_5984);
xnor U7058 (N_7058,N_5782,N_5699);
or U7059 (N_7059,N_5844,N_4954);
nand U7060 (N_7060,N_5277,N_5004);
or U7061 (N_7061,N_4848,N_5673);
nand U7062 (N_7062,N_5115,N_4989);
nor U7063 (N_7063,N_5533,N_4830);
nand U7064 (N_7064,N_5553,N_5890);
or U7065 (N_7065,N_5934,N_5450);
xnor U7066 (N_7066,N_5654,N_5164);
xor U7067 (N_7067,N_5599,N_5035);
or U7068 (N_7068,N_5029,N_5752);
xor U7069 (N_7069,N_5427,N_5536);
or U7070 (N_7070,N_4933,N_5030);
and U7071 (N_7071,N_4841,N_5595);
or U7072 (N_7072,N_5387,N_5624);
xnor U7073 (N_7073,N_4859,N_4863);
nor U7074 (N_7074,N_5728,N_5551);
nand U7075 (N_7075,N_5964,N_4950);
nand U7076 (N_7076,N_5542,N_5843);
or U7077 (N_7077,N_5062,N_5386);
or U7078 (N_7078,N_5304,N_4871);
nand U7079 (N_7079,N_5031,N_5623);
nor U7080 (N_7080,N_5818,N_5611);
nor U7081 (N_7081,N_5585,N_4842);
or U7082 (N_7082,N_5590,N_5853);
xor U7083 (N_7083,N_5689,N_5035);
nand U7084 (N_7084,N_5302,N_5871);
nand U7085 (N_7085,N_5510,N_5985);
nor U7086 (N_7086,N_5477,N_5276);
and U7087 (N_7087,N_4821,N_5938);
nor U7088 (N_7088,N_5588,N_5787);
xor U7089 (N_7089,N_5181,N_5003);
or U7090 (N_7090,N_5594,N_5962);
nor U7091 (N_7091,N_4991,N_5832);
nor U7092 (N_7092,N_5863,N_5007);
and U7093 (N_7093,N_5741,N_5816);
and U7094 (N_7094,N_5716,N_5140);
xor U7095 (N_7095,N_5249,N_5393);
or U7096 (N_7096,N_5818,N_5692);
or U7097 (N_7097,N_5201,N_5706);
nor U7098 (N_7098,N_5214,N_5372);
xor U7099 (N_7099,N_5066,N_5130);
nand U7100 (N_7100,N_5511,N_5394);
or U7101 (N_7101,N_5260,N_5247);
and U7102 (N_7102,N_5981,N_4971);
nor U7103 (N_7103,N_5932,N_5458);
and U7104 (N_7104,N_5960,N_4924);
and U7105 (N_7105,N_5818,N_5329);
nor U7106 (N_7106,N_5431,N_5374);
and U7107 (N_7107,N_5484,N_5255);
nand U7108 (N_7108,N_5024,N_5591);
or U7109 (N_7109,N_5679,N_4809);
nor U7110 (N_7110,N_5505,N_4960);
xnor U7111 (N_7111,N_5470,N_5475);
nor U7112 (N_7112,N_5690,N_5534);
xor U7113 (N_7113,N_5867,N_5309);
and U7114 (N_7114,N_4861,N_5992);
nand U7115 (N_7115,N_4883,N_5481);
and U7116 (N_7116,N_5467,N_4867);
xor U7117 (N_7117,N_5286,N_5087);
xnor U7118 (N_7118,N_5168,N_5200);
nor U7119 (N_7119,N_5708,N_5955);
nand U7120 (N_7120,N_5810,N_5005);
and U7121 (N_7121,N_4825,N_5901);
nor U7122 (N_7122,N_5020,N_5534);
nand U7123 (N_7123,N_4832,N_5280);
or U7124 (N_7124,N_5202,N_5125);
nor U7125 (N_7125,N_5099,N_5323);
xor U7126 (N_7126,N_5243,N_5363);
nand U7127 (N_7127,N_5812,N_5462);
nand U7128 (N_7128,N_4894,N_5564);
nand U7129 (N_7129,N_4917,N_5538);
xor U7130 (N_7130,N_5349,N_5995);
and U7131 (N_7131,N_5661,N_4878);
xor U7132 (N_7132,N_5797,N_5780);
nor U7133 (N_7133,N_5718,N_4889);
nand U7134 (N_7134,N_5514,N_5778);
xor U7135 (N_7135,N_5091,N_5301);
and U7136 (N_7136,N_5338,N_5384);
xnor U7137 (N_7137,N_5272,N_5325);
xor U7138 (N_7138,N_5387,N_5556);
or U7139 (N_7139,N_5333,N_5025);
and U7140 (N_7140,N_5587,N_5660);
xnor U7141 (N_7141,N_5764,N_5390);
nand U7142 (N_7142,N_5472,N_5818);
or U7143 (N_7143,N_4990,N_5226);
nand U7144 (N_7144,N_5579,N_5747);
or U7145 (N_7145,N_5207,N_5549);
nand U7146 (N_7146,N_5241,N_5900);
nand U7147 (N_7147,N_4844,N_5460);
and U7148 (N_7148,N_5782,N_5259);
xor U7149 (N_7149,N_5070,N_4814);
or U7150 (N_7150,N_5736,N_5077);
nor U7151 (N_7151,N_5437,N_5340);
and U7152 (N_7152,N_5839,N_5399);
xnor U7153 (N_7153,N_5455,N_5116);
or U7154 (N_7154,N_5859,N_5015);
and U7155 (N_7155,N_5704,N_5982);
nand U7156 (N_7156,N_5962,N_5921);
or U7157 (N_7157,N_5012,N_5721);
nand U7158 (N_7158,N_5055,N_5148);
nand U7159 (N_7159,N_5707,N_5182);
and U7160 (N_7160,N_5937,N_5940);
xor U7161 (N_7161,N_5431,N_5451);
xor U7162 (N_7162,N_5421,N_5695);
nor U7163 (N_7163,N_5586,N_5604);
or U7164 (N_7164,N_5352,N_4913);
xnor U7165 (N_7165,N_5155,N_5697);
or U7166 (N_7166,N_4921,N_5014);
and U7167 (N_7167,N_5979,N_5709);
nand U7168 (N_7168,N_5237,N_5748);
or U7169 (N_7169,N_4921,N_4864);
nor U7170 (N_7170,N_5110,N_5552);
and U7171 (N_7171,N_5112,N_5535);
xnor U7172 (N_7172,N_5973,N_5068);
or U7173 (N_7173,N_5659,N_5465);
or U7174 (N_7174,N_5890,N_5739);
or U7175 (N_7175,N_5052,N_4824);
or U7176 (N_7176,N_5103,N_5460);
nand U7177 (N_7177,N_5906,N_5049);
and U7178 (N_7178,N_5115,N_5747);
nor U7179 (N_7179,N_5637,N_5260);
nand U7180 (N_7180,N_4855,N_5039);
nor U7181 (N_7181,N_5642,N_5260);
nor U7182 (N_7182,N_5079,N_5690);
and U7183 (N_7183,N_5285,N_4977);
nor U7184 (N_7184,N_4819,N_5533);
nor U7185 (N_7185,N_5158,N_5425);
and U7186 (N_7186,N_4967,N_4859);
nor U7187 (N_7187,N_5106,N_4835);
nand U7188 (N_7188,N_5383,N_5500);
and U7189 (N_7189,N_5379,N_5513);
xor U7190 (N_7190,N_5611,N_5955);
or U7191 (N_7191,N_5951,N_5008);
and U7192 (N_7192,N_5117,N_5057);
and U7193 (N_7193,N_5632,N_5241);
nand U7194 (N_7194,N_5483,N_5339);
and U7195 (N_7195,N_5514,N_5919);
xor U7196 (N_7196,N_5746,N_5154);
or U7197 (N_7197,N_5450,N_5522);
xor U7198 (N_7198,N_5956,N_4811);
xnor U7199 (N_7199,N_5987,N_4951);
and U7200 (N_7200,N_6422,N_6444);
nand U7201 (N_7201,N_7131,N_6036);
and U7202 (N_7202,N_6851,N_6742);
or U7203 (N_7203,N_6349,N_6842);
nand U7204 (N_7204,N_6386,N_6876);
nor U7205 (N_7205,N_6594,N_6301);
xor U7206 (N_7206,N_6912,N_6617);
nand U7207 (N_7207,N_6189,N_6153);
or U7208 (N_7208,N_6062,N_6995);
xor U7209 (N_7209,N_6275,N_6928);
nand U7210 (N_7210,N_6103,N_6091);
nor U7211 (N_7211,N_6320,N_7152);
or U7212 (N_7212,N_6493,N_6272);
nor U7213 (N_7213,N_6824,N_7033);
or U7214 (N_7214,N_6451,N_6508);
xor U7215 (N_7215,N_6407,N_7104);
nand U7216 (N_7216,N_7074,N_6013);
nor U7217 (N_7217,N_6828,N_6981);
or U7218 (N_7218,N_6843,N_6185);
and U7219 (N_7219,N_6055,N_6672);
nand U7220 (N_7220,N_6001,N_6381);
nor U7221 (N_7221,N_6316,N_7170);
nor U7222 (N_7222,N_6504,N_6171);
or U7223 (N_7223,N_6243,N_6741);
nand U7224 (N_7224,N_6433,N_6633);
or U7225 (N_7225,N_7044,N_7123);
and U7226 (N_7226,N_6092,N_7120);
xnor U7227 (N_7227,N_7012,N_6994);
xnor U7228 (N_7228,N_6781,N_6966);
or U7229 (N_7229,N_6247,N_7070);
nand U7230 (N_7230,N_6748,N_6608);
xnor U7231 (N_7231,N_6277,N_6464);
nor U7232 (N_7232,N_6454,N_6478);
and U7233 (N_7233,N_6979,N_7112);
nand U7234 (N_7234,N_6144,N_6197);
and U7235 (N_7235,N_7197,N_7137);
nand U7236 (N_7236,N_7018,N_7179);
and U7237 (N_7237,N_6329,N_7061);
or U7238 (N_7238,N_6399,N_6941);
and U7239 (N_7239,N_6899,N_6612);
or U7240 (N_7240,N_6836,N_6701);
and U7241 (N_7241,N_7181,N_6921);
nand U7242 (N_7242,N_6235,N_6116);
or U7243 (N_7243,N_6064,N_6098);
and U7244 (N_7244,N_6840,N_6990);
or U7245 (N_7245,N_6854,N_6203);
and U7246 (N_7246,N_6948,N_6778);
or U7247 (N_7247,N_6218,N_7083);
or U7248 (N_7248,N_6459,N_6711);
or U7249 (N_7249,N_6592,N_6527);
or U7250 (N_7250,N_6727,N_7023);
and U7251 (N_7251,N_6968,N_6883);
nand U7252 (N_7252,N_6517,N_6667);
or U7253 (N_7253,N_6202,N_6580);
and U7254 (N_7254,N_6264,N_6702);
xor U7255 (N_7255,N_6246,N_6986);
or U7256 (N_7256,N_6518,N_6686);
or U7257 (N_7257,N_6101,N_7186);
or U7258 (N_7258,N_6368,N_6113);
or U7259 (N_7259,N_6880,N_6031);
nand U7260 (N_7260,N_6654,N_6249);
or U7261 (N_7261,N_7065,N_6201);
and U7262 (N_7262,N_6513,N_6957);
and U7263 (N_7263,N_6437,N_6790);
nor U7264 (N_7264,N_6128,N_6998);
and U7265 (N_7265,N_6176,N_7085);
nor U7266 (N_7266,N_6578,N_6678);
nand U7267 (N_7267,N_7160,N_6895);
nand U7268 (N_7268,N_6210,N_6314);
or U7269 (N_7269,N_6465,N_6814);
or U7270 (N_7270,N_6687,N_6147);
and U7271 (N_7271,N_6328,N_6042);
and U7272 (N_7272,N_6310,N_6457);
and U7273 (N_7273,N_6446,N_6567);
nor U7274 (N_7274,N_6354,N_6233);
or U7275 (N_7275,N_6306,N_6412);
or U7276 (N_7276,N_7121,N_6124);
or U7277 (N_7277,N_6769,N_6273);
or U7278 (N_7278,N_6905,N_6351);
and U7279 (N_7279,N_6281,N_7095);
nand U7280 (N_7280,N_6122,N_6510);
and U7281 (N_7281,N_6058,N_6041);
nor U7282 (N_7282,N_6779,N_6269);
and U7283 (N_7283,N_6174,N_7084);
and U7284 (N_7284,N_7029,N_6123);
and U7285 (N_7285,N_6010,N_6544);
nand U7286 (N_7286,N_6333,N_6516);
nand U7287 (N_7287,N_6522,N_6619);
nor U7288 (N_7288,N_6056,N_6117);
nand U7289 (N_7289,N_7056,N_6557);
and U7290 (N_7290,N_6776,N_6016);
or U7291 (N_7291,N_6724,N_6323);
nor U7292 (N_7292,N_6024,N_6733);
or U7293 (N_7293,N_7184,N_6983);
and U7294 (N_7294,N_6216,N_6401);
nand U7295 (N_7295,N_7149,N_6213);
or U7296 (N_7296,N_6258,N_7043);
and U7297 (N_7297,N_6436,N_6652);
or U7298 (N_7298,N_6052,N_6474);
xnor U7299 (N_7299,N_7047,N_6632);
nor U7300 (N_7300,N_6028,N_6607);
xor U7301 (N_7301,N_6536,N_6429);
xor U7302 (N_7302,N_6127,N_7117);
nand U7303 (N_7303,N_6388,N_7193);
nand U7304 (N_7304,N_6560,N_7159);
nor U7305 (N_7305,N_6735,N_6975);
and U7306 (N_7306,N_6494,N_6573);
or U7307 (N_7307,N_6805,N_6085);
nor U7308 (N_7308,N_6974,N_6390);
nor U7309 (N_7309,N_7192,N_6749);
nand U7310 (N_7310,N_6938,N_6581);
xor U7311 (N_7311,N_6045,N_6468);
xor U7312 (N_7312,N_7093,N_6878);
or U7313 (N_7313,N_7060,N_6224);
and U7314 (N_7314,N_6331,N_7140);
nor U7315 (N_7315,N_7180,N_6409);
nor U7316 (N_7316,N_6146,N_7054);
nor U7317 (N_7317,N_7068,N_6196);
and U7318 (N_7318,N_7031,N_7183);
nand U7319 (N_7319,N_6673,N_6019);
and U7320 (N_7320,N_6708,N_6078);
and U7321 (N_7321,N_6487,N_7053);
nor U7322 (N_7322,N_6298,N_6115);
nand U7323 (N_7323,N_6783,N_7147);
nor U7324 (N_7324,N_6547,N_6897);
xor U7325 (N_7325,N_6151,N_7036);
and U7326 (N_7326,N_6138,N_7004);
nor U7327 (N_7327,N_6473,N_6102);
nor U7328 (N_7328,N_6661,N_6743);
nor U7329 (N_7329,N_6162,N_7167);
nand U7330 (N_7330,N_6130,N_6793);
nand U7331 (N_7331,N_6336,N_6671);
nor U7332 (N_7332,N_6448,N_6432);
xnor U7333 (N_7333,N_6097,N_6466);
nor U7334 (N_7334,N_6035,N_7046);
xor U7335 (N_7335,N_6345,N_7002);
nor U7336 (N_7336,N_6060,N_6898);
and U7337 (N_7337,N_6295,N_6768);
xnor U7338 (N_7338,N_7113,N_6713);
xor U7339 (N_7339,N_6942,N_7037);
nand U7340 (N_7340,N_6395,N_7088);
xnor U7341 (N_7341,N_6148,N_6199);
or U7342 (N_7342,N_6903,N_6657);
and U7343 (N_7343,N_6022,N_6077);
and U7344 (N_7344,N_6435,N_7163);
nor U7345 (N_7345,N_6591,N_6606);
nor U7346 (N_7346,N_6579,N_6152);
nand U7347 (N_7347,N_6809,N_7017);
and U7348 (N_7348,N_6523,N_7020);
nand U7349 (N_7349,N_6865,N_6441);
nand U7350 (N_7350,N_6166,N_6009);
and U7351 (N_7351,N_6566,N_6112);
xor U7352 (N_7352,N_6070,N_6373);
xnor U7353 (N_7353,N_6369,N_7116);
or U7354 (N_7354,N_7196,N_6620);
nor U7355 (N_7355,N_6495,N_6861);
nand U7356 (N_7356,N_6204,N_6274);
nor U7357 (N_7357,N_6629,N_7075);
nand U7358 (N_7358,N_6181,N_6018);
xor U7359 (N_7359,N_6260,N_6406);
nand U7360 (N_7360,N_6556,N_6255);
or U7361 (N_7361,N_6154,N_7114);
xor U7362 (N_7362,N_7059,N_6421);
nand U7363 (N_7363,N_6521,N_6683);
nor U7364 (N_7364,N_6926,N_6625);
nand U7365 (N_7365,N_6073,N_6384);
xor U7366 (N_7366,N_6830,N_7127);
nand U7367 (N_7367,N_6428,N_7158);
or U7368 (N_7368,N_7190,N_6392);
nand U7369 (N_7369,N_6884,N_6665);
nand U7370 (N_7370,N_6643,N_6961);
or U7371 (N_7371,N_6832,N_6215);
and U7372 (N_7372,N_7150,N_6284);
nor U7373 (N_7373,N_7154,N_6826);
xnor U7374 (N_7374,N_6820,N_6136);
or U7375 (N_7375,N_6304,N_6554);
or U7376 (N_7376,N_7051,N_6370);
and U7377 (N_7377,N_7132,N_6935);
nor U7378 (N_7378,N_6256,N_7134);
nand U7379 (N_7379,N_6096,N_6038);
xor U7380 (N_7380,N_6584,N_6653);
and U7381 (N_7381,N_6924,N_6909);
or U7382 (N_7382,N_6332,N_6853);
nor U7383 (N_7383,N_6956,N_6712);
xor U7384 (N_7384,N_6866,N_6195);
xnor U7385 (N_7385,N_6729,N_6798);
xor U7386 (N_7386,N_6261,N_6358);
xor U7387 (N_7387,N_7019,N_6722);
nor U7388 (N_7388,N_6469,N_6416);
nand U7389 (N_7389,N_6142,N_6699);
nand U7390 (N_7390,N_6426,N_6500);
and U7391 (N_7391,N_6794,N_6543);
and U7392 (N_7392,N_6186,N_6491);
or U7393 (N_7393,N_6126,N_6582);
or U7394 (N_7394,N_6890,N_6476);
xor U7395 (N_7395,N_6574,N_6925);
xnor U7396 (N_7396,N_6453,N_6172);
xor U7397 (N_7397,N_6593,N_6503);
xor U7398 (N_7398,N_6691,N_6973);
xnor U7399 (N_7399,N_6291,N_6475);
nor U7400 (N_7400,N_6161,N_7042);
and U7401 (N_7401,N_6636,N_6044);
and U7402 (N_7402,N_6221,N_6006);
or U7403 (N_7403,N_6936,N_6850);
xor U7404 (N_7404,N_6312,N_6755);
xor U7405 (N_7405,N_6685,N_6847);
or U7406 (N_7406,N_6764,N_6682);
nor U7407 (N_7407,N_6962,N_7010);
nand U7408 (N_7408,N_6537,N_6819);
nand U7409 (N_7409,N_6463,N_6051);
and U7410 (N_7410,N_7141,N_6859);
nor U7411 (N_7411,N_6303,N_6848);
or U7412 (N_7412,N_7143,N_6738);
or U7413 (N_7413,N_6757,N_6697);
xor U7414 (N_7414,N_6046,N_6940);
and U7415 (N_7415,N_6911,N_6797);
xor U7416 (N_7416,N_6397,N_6095);
xor U7417 (N_7417,N_6572,N_7130);
or U7418 (N_7418,N_6963,N_6139);
xor U7419 (N_7419,N_6262,N_6311);
nand U7420 (N_7420,N_7125,N_6109);
and U7421 (N_7421,N_6869,N_6761);
nand U7422 (N_7422,N_6945,N_6470);
or U7423 (N_7423,N_6834,N_6565);
xor U7424 (N_7424,N_6377,N_6561);
and U7425 (N_7425,N_6693,N_6057);
xor U7426 (N_7426,N_7021,N_6075);
nand U7427 (N_7427,N_6084,N_6539);
or U7428 (N_7428,N_7066,N_6932);
and U7429 (N_7429,N_6319,N_6484);
nand U7430 (N_7430,N_6003,N_6969);
xor U7431 (N_7431,N_6588,N_6913);
nor U7432 (N_7432,N_7138,N_7173);
nor U7433 (N_7433,N_6879,N_6656);
nand U7434 (N_7434,N_6119,N_6135);
nand U7435 (N_7435,N_6835,N_6944);
nor U7436 (N_7436,N_6257,N_6511);
and U7437 (N_7437,N_7005,N_6296);
and U7438 (N_7438,N_7055,N_6613);
xor U7439 (N_7439,N_6007,N_6694);
nor U7440 (N_7440,N_6447,N_6049);
or U7441 (N_7441,N_6339,N_6456);
nor U7442 (N_7442,N_6745,N_7162);
nor U7443 (N_7443,N_6756,N_6791);
or U7444 (N_7444,N_6692,N_6106);
nor U7445 (N_7445,N_6223,N_6417);
nand U7446 (N_7446,N_7091,N_7009);
or U7447 (N_7447,N_6970,N_6307);
nand U7448 (N_7448,N_7040,N_6040);
or U7449 (N_7449,N_6398,N_6187);
or U7450 (N_7450,N_6371,N_6927);
and U7451 (N_7451,N_6562,N_6150);
and U7452 (N_7452,N_6750,N_6770);
nand U7453 (N_7453,N_6603,N_6061);
or U7454 (N_7454,N_6767,N_6870);
or U7455 (N_7455,N_6918,N_6167);
and U7456 (N_7456,N_6266,N_7006);
nand U7457 (N_7457,N_6496,N_6991);
or U7458 (N_7458,N_6618,N_6967);
nor U7459 (N_7459,N_6731,N_6964);
and U7460 (N_7460,N_7100,N_6270);
xnor U7461 (N_7461,N_6568,N_6011);
or U7462 (N_7462,N_6093,N_6226);
nor U7463 (N_7463,N_6728,N_6361);
or U7464 (N_7464,N_6334,N_7097);
and U7465 (N_7465,N_6048,N_6411);
and U7466 (N_7466,N_7049,N_7098);
nand U7467 (N_7467,N_6133,N_6839);
and U7468 (N_7468,N_6740,N_6340);
and U7469 (N_7469,N_7000,N_6483);
xor U7470 (N_7470,N_6739,N_7057);
xnor U7471 (N_7471,N_7030,N_7025);
nor U7472 (N_7472,N_6670,N_6610);
or U7473 (N_7473,N_7191,N_6989);
nand U7474 (N_7474,N_6442,N_6378);
and U7475 (N_7475,N_6472,N_6467);
nor U7476 (N_7476,N_6540,N_6631);
or U7477 (N_7477,N_6951,N_7078);
xor U7478 (N_7478,N_6232,N_6773);
nand U7479 (N_7479,N_6954,N_7032);
and U7480 (N_7480,N_6279,N_6730);
nand U7481 (N_7481,N_6424,N_7014);
and U7482 (N_7482,N_6071,N_6775);
or U7483 (N_7483,N_6772,N_6714);
nor U7484 (N_7484,N_6276,N_6183);
or U7485 (N_7485,N_6357,N_7166);
or U7486 (N_7486,N_6532,N_6887);
and U7487 (N_7487,N_6004,N_6282);
nand U7488 (N_7488,N_6359,N_6716);
nand U7489 (N_7489,N_6507,N_6259);
and U7490 (N_7490,N_6821,N_6317);
xnor U7491 (N_7491,N_6910,N_6977);
xnor U7492 (N_7492,N_6251,N_6346);
or U7493 (N_7493,N_6118,N_7153);
nand U7494 (N_7494,N_6882,N_6054);
and U7495 (N_7495,N_6434,N_6627);
nand U7496 (N_7496,N_6747,N_6953);
nand U7497 (N_7497,N_7109,N_6015);
or U7498 (N_7498,N_6512,N_6400);
or U7499 (N_7499,N_6173,N_7108);
or U7500 (N_7500,N_6647,N_6245);
and U7501 (N_7501,N_6025,N_6929);
nor U7502 (N_7502,N_6486,N_7148);
or U7503 (N_7503,N_6032,N_6877);
and U7504 (N_7504,N_6389,N_6121);
nand U7505 (N_7505,N_6156,N_6703);
nand U7506 (N_7506,N_6595,N_6611);
nand U7507 (N_7507,N_6047,N_6219);
nand U7508 (N_7508,N_6355,N_6342);
nand U7509 (N_7509,N_6250,N_6017);
or U7510 (N_7510,N_6885,N_6445);
nor U7511 (N_7511,N_6053,N_6391);
nand U7512 (N_7512,N_7102,N_7022);
nand U7513 (N_7513,N_6583,N_6005);
nor U7514 (N_7514,N_6080,N_6800);
or U7515 (N_7515,N_6450,N_6165);
or U7516 (N_7516,N_6709,N_6947);
nand U7517 (N_7517,N_6815,N_6002);
and U7518 (N_7518,N_6037,N_6083);
or U7519 (N_7519,N_6230,N_6157);
nand U7520 (N_7520,N_7146,N_6293);
nand U7521 (N_7521,N_6972,N_6363);
or U7522 (N_7522,N_6253,N_6132);
nand U7523 (N_7523,N_6405,N_6829);
nand U7524 (N_7524,N_6987,N_6072);
and U7525 (N_7525,N_6430,N_6922);
nor U7526 (N_7526,N_6177,N_7129);
xnor U7527 (N_7527,N_6680,N_6825);
and U7528 (N_7528,N_7174,N_6271);
and U7529 (N_7529,N_6178,N_6525);
nor U7530 (N_7530,N_6980,N_6376);
or U7531 (N_7531,N_6640,N_6352);
nand U7532 (N_7532,N_6637,N_7105);
nor U7533 (N_7533,N_6471,N_6863);
nor U7534 (N_7534,N_6971,N_6033);
nor U7535 (N_7535,N_6318,N_6344);
nor U7536 (N_7536,N_6324,N_6894);
xnor U7537 (N_7537,N_6217,N_6753);
or U7538 (N_7538,N_6190,N_6404);
nand U7539 (N_7539,N_6238,N_6094);
and U7540 (N_7540,N_6958,N_6020);
and U7541 (N_7541,N_6191,N_6188);
or U7542 (N_7542,N_6758,N_6237);
nor U7543 (N_7543,N_6244,N_6563);
or U7544 (N_7544,N_6184,N_6485);
nor U7545 (N_7545,N_7011,N_6000);
nor U7546 (N_7546,N_6548,N_6065);
nor U7547 (N_7547,N_6916,N_6628);
xor U7548 (N_7548,N_6182,N_6804);
and U7549 (N_7549,N_6666,N_6646);
nor U7550 (N_7550,N_6600,N_6641);
nor U7551 (N_7551,N_6802,N_7099);
or U7552 (N_7552,N_7168,N_6228);
nor U7553 (N_7553,N_6597,N_6659);
nand U7554 (N_7554,N_6626,N_6949);
and U7555 (N_7555,N_6481,N_6695);
xor U7556 (N_7556,N_6066,N_7124);
and U7557 (N_7557,N_6789,N_6414);
xnor U7558 (N_7558,N_6831,N_6734);
or U7559 (N_7559,N_6497,N_6908);
nor U7560 (N_7560,N_6658,N_6871);
or U7561 (N_7561,N_7089,N_6131);
xor U7562 (N_7562,N_6639,N_6978);
nor U7563 (N_7563,N_6596,N_6089);
xnor U7564 (N_7564,N_6982,N_6423);
nor U7565 (N_7565,N_6589,N_6933);
xor U7566 (N_7566,N_6872,N_6891);
or U7567 (N_7567,N_6205,N_6689);
xor U7568 (N_7568,N_6531,N_6993);
and U7569 (N_7569,N_6315,N_6787);
and U7570 (N_7570,N_6519,N_7079);
and U7571 (N_7571,N_7077,N_6305);
xnor U7572 (N_7572,N_6140,N_6645);
nand U7573 (N_7573,N_6746,N_6413);
xnor U7574 (N_7574,N_6239,N_6766);
xor U7575 (N_7575,N_6438,N_7151);
xnor U7576 (N_7576,N_6192,N_6137);
xnor U7577 (N_7577,N_6943,N_6515);
xor U7578 (N_7578,N_6586,N_6785);
or U7579 (N_7579,N_6427,N_6759);
nor U7580 (N_7580,N_6559,N_6396);
nor U7581 (N_7581,N_6867,N_6719);
or U7582 (N_7582,N_6914,N_6375);
or U7583 (N_7583,N_6030,N_6208);
nand U7584 (N_7584,N_7072,N_6159);
nor U7585 (N_7585,N_6648,N_7024);
or U7586 (N_7586,N_6535,N_7171);
or U7587 (N_7587,N_6452,N_7144);
nor U7588 (N_7588,N_6415,N_6664);
or U7589 (N_7589,N_6598,N_6919);
or U7590 (N_7590,N_6059,N_6668);
xor U7591 (N_7591,N_6777,N_6360);
xor U7592 (N_7592,N_6571,N_6679);
nor U7593 (N_7593,N_6546,N_7076);
nor U7594 (N_7594,N_6341,N_7090);
and U7595 (N_7595,N_6149,N_7145);
and U7596 (N_7596,N_6207,N_7107);
and U7597 (N_7597,N_6267,N_7087);
and U7598 (N_7598,N_6505,N_6630);
xnor U7599 (N_7599,N_6616,N_6550);
nand U7600 (N_7600,N_6858,N_6886);
nor U7601 (N_7601,N_6214,N_6601);
nor U7602 (N_7602,N_6299,N_6621);
or U7603 (N_7603,N_6420,N_6960);
and U7604 (N_7604,N_7195,N_6372);
nand U7605 (N_7605,N_7165,N_7086);
or U7606 (N_7606,N_6380,N_6988);
and U7607 (N_7607,N_6801,N_6286);
xor U7608 (N_7608,N_6599,N_6367);
and U7609 (N_7609,N_7001,N_6726);
nor U7610 (N_7610,N_6717,N_6997);
xnor U7611 (N_7611,N_6076,N_6087);
and U7612 (N_7612,N_7187,N_6393);
or U7613 (N_7613,N_6252,N_6439);
or U7614 (N_7614,N_6827,N_7039);
nand U7615 (N_7615,N_6488,N_6164);
nand U7616 (N_7616,N_7198,N_6294);
and U7617 (N_7617,N_6337,N_6043);
nor U7618 (N_7618,N_6227,N_7136);
nor U7619 (N_7619,N_6220,N_6774);
or U7620 (N_7620,N_6461,N_6996);
nand U7621 (N_7621,N_6602,N_6180);
xnor U7622 (N_7622,N_6552,N_6736);
nor U7623 (N_7623,N_6212,N_6034);
nor U7624 (N_7624,N_6283,N_6855);
and U7625 (N_7625,N_6482,N_6737);
nor U7626 (N_7626,N_7062,N_6690);
xnor U7627 (N_7627,N_6309,N_6169);
and U7628 (N_7628,N_7041,N_6240);
nor U7629 (N_7629,N_7157,N_6462);
and U7630 (N_7630,N_6330,N_6923);
or U7631 (N_7631,N_6873,N_6479);
or U7632 (N_7632,N_6575,N_6538);
xor U7633 (N_7633,N_6822,N_6338);
nand U7634 (N_7634,N_7182,N_6385);
nor U7635 (N_7635,N_6526,N_6108);
and U7636 (N_7636,N_7045,N_6343);
or U7637 (N_7637,N_6782,N_6350);
nor U7638 (N_7638,N_6506,N_6129);
nor U7639 (N_7639,N_6322,N_6881);
xor U7640 (N_7640,N_6353,N_6431);
nand U7641 (N_7641,N_6460,N_7063);
nand U7642 (N_7642,N_7155,N_6784);
nand U7643 (N_7643,N_6965,N_6026);
or U7644 (N_7644,N_6795,N_6934);
or U7645 (N_7645,N_6752,N_6651);
or U7646 (N_7646,N_6955,N_6817);
or U7647 (N_7647,N_6528,N_6570);
nand U7648 (N_7648,N_6930,N_6676);
xor U7649 (N_7649,N_6104,N_7164);
nand U7650 (N_7650,N_7064,N_6248);
and U7651 (N_7651,N_6107,N_6732);
or U7652 (N_7652,N_6638,N_6175);
or U7653 (N_7653,N_6263,N_6348);
and U7654 (N_7654,N_6120,N_6896);
xnor U7655 (N_7655,N_6321,N_7135);
nor U7656 (N_7656,N_6624,N_6143);
xor U7657 (N_7657,N_6014,N_6039);
or U7658 (N_7658,N_6168,N_6145);
xor U7659 (N_7659,N_6862,N_6950);
or U7660 (N_7660,N_6892,N_6549);
and U7661 (N_7661,N_6242,N_6590);
xor U7662 (N_7662,N_6362,N_7052);
nand U7663 (N_7663,N_6684,N_6302);
and U7664 (N_7664,N_7015,N_6771);
nand U7665 (N_7665,N_6762,N_6287);
or U7666 (N_7666,N_6707,N_6806);
xor U7667 (N_7667,N_6786,N_6520);
xor U7668 (N_7668,N_6408,N_6674);
or U7669 (N_7669,N_6833,N_7034);
or U7670 (N_7670,N_6999,N_6799);
nand U7671 (N_7671,N_6347,N_6803);
nand U7672 (N_7672,N_6440,N_6265);
nor U7673 (N_7673,N_6300,N_6939);
nand U7674 (N_7674,N_6696,N_6356);
xor U7675 (N_7675,N_6125,N_6290);
or U7676 (N_7676,N_7177,N_6788);
nor U7677 (N_7677,N_7139,N_6327);
nand U7678 (N_7678,N_6236,N_6234);
or U7679 (N_7679,N_6141,N_6751);
xor U7680 (N_7680,N_7126,N_6655);
and U7681 (N_7681,N_6816,N_7008);
or U7682 (N_7682,N_6615,N_7185);
nand U7683 (N_7683,N_6023,N_6838);
or U7684 (N_7684,N_7081,N_7103);
nor U7685 (N_7685,N_6514,N_6681);
xnor U7686 (N_7686,N_6533,N_6292);
nor U7687 (N_7687,N_7073,N_6326);
or U7688 (N_7688,N_7161,N_6365);
and U7689 (N_7689,N_6710,N_6379);
or U7690 (N_7690,N_6099,N_6489);
nand U7691 (N_7691,N_6383,N_6170);
xnor U7692 (N_7692,N_6985,N_6364);
nor U7693 (N_7693,N_6622,N_6082);
xnor U7694 (N_7694,N_6642,N_6335);
or U7695 (N_7695,N_6846,N_6754);
and U7696 (N_7696,N_7050,N_6366);
or U7697 (N_7697,N_7118,N_6864);
or U7698 (N_7698,N_6792,N_6609);
and U7699 (N_7699,N_7194,N_6050);
xnor U7700 (N_7700,N_7172,N_6067);
xnor U7701 (N_7701,N_7035,N_7013);
and U7702 (N_7702,N_6325,N_6875);
xor U7703 (N_7703,N_7038,N_6425);
nor U7704 (N_7704,N_6160,N_6946);
or U7705 (N_7705,N_6410,N_6976);
xor U7706 (N_7706,N_6564,N_6198);
or U7707 (N_7707,N_6499,N_6577);
and U7708 (N_7708,N_6663,N_6984);
nand U7709 (N_7709,N_6553,N_6086);
and U7710 (N_7710,N_6081,N_6718);
nand U7711 (N_7711,N_6194,N_6623);
xor U7712 (N_7712,N_6818,N_7027);
nand U7713 (N_7713,N_7101,N_6289);
nand U7714 (N_7714,N_6992,N_6915);
nor U7715 (N_7715,N_7106,N_6551);
xnor U7716 (N_7716,N_6675,N_6254);
nor U7717 (N_7717,N_6837,N_6874);
nand U7718 (N_7718,N_6209,N_6480);
and U7719 (N_7719,N_7067,N_7071);
nand U7720 (N_7720,N_6931,N_6725);
nand U7721 (N_7721,N_6394,N_6900);
or U7722 (N_7722,N_6545,N_6587);
nor U7723 (N_7723,N_6229,N_6576);
nor U7724 (N_7724,N_6660,N_6111);
and U7725 (N_7725,N_6849,N_7119);
and U7726 (N_7726,N_6952,N_7092);
nor U7727 (N_7727,N_6715,N_7028);
nand U7728 (N_7728,N_6644,N_6313);
or U7729 (N_7729,N_7156,N_6158);
and U7730 (N_7730,N_6604,N_6268);
and U7731 (N_7731,N_6860,N_7176);
and U7732 (N_7732,N_6524,N_6542);
and U7733 (N_7733,N_6297,N_6029);
nor U7734 (N_7734,N_6856,N_6907);
nand U7735 (N_7735,N_6534,N_6477);
xor U7736 (N_7736,N_6280,N_6231);
and U7737 (N_7737,N_6490,N_7115);
or U7738 (N_7738,N_7082,N_6222);
xnor U7739 (N_7739,N_6419,N_6796);
xnor U7740 (N_7740,N_6455,N_6649);
and U7741 (N_7741,N_6114,N_6845);
xor U7742 (N_7742,N_6698,N_6241);
xnor U7743 (N_7743,N_6721,N_6634);
xnor U7744 (N_7744,N_7016,N_6068);
nand U7745 (N_7745,N_6206,N_6211);
or U7746 (N_7746,N_6012,N_6288);
or U7747 (N_7747,N_6901,N_6959);
nand U7748 (N_7748,N_6823,N_6090);
nor U7749 (N_7749,N_7094,N_6449);
and U7750 (N_7750,N_6134,N_6852);
nor U7751 (N_7751,N_6720,N_6179);
or U7752 (N_7752,N_7175,N_6677);
nor U7753 (N_7753,N_6458,N_6723);
xnor U7754 (N_7754,N_7133,N_7069);
nand U7755 (N_7755,N_7110,N_6889);
or U7756 (N_7756,N_7169,N_6705);
or U7757 (N_7757,N_6308,N_6700);
nand U7758 (N_7758,N_6509,N_6225);
or U7759 (N_7759,N_7188,N_6555);
and U7760 (N_7760,N_7058,N_6063);
and U7761 (N_7761,N_6635,N_6069);
nor U7762 (N_7762,N_6920,N_6811);
and U7763 (N_7763,N_6027,N_6763);
and U7764 (N_7764,N_6402,N_6917);
and U7765 (N_7765,N_6857,N_6558);
nor U7766 (N_7766,N_6902,N_6807);
xnor U7767 (N_7767,N_6100,N_7178);
and U7768 (N_7768,N_6808,N_7026);
or U7769 (N_7769,N_6704,N_7048);
and U7770 (N_7770,N_6403,N_7007);
xnor U7771 (N_7771,N_6008,N_6669);
xnor U7772 (N_7772,N_6812,N_6844);
nor U7773 (N_7773,N_6706,N_6105);
xor U7774 (N_7774,N_6780,N_6021);
and U7775 (N_7775,N_7096,N_6906);
and U7776 (N_7776,N_6418,N_6662);
xnor U7777 (N_7777,N_6585,N_6278);
and U7778 (N_7778,N_7080,N_6569);
or U7779 (N_7779,N_6088,N_6163);
or U7780 (N_7780,N_6285,N_6893);
nor U7781 (N_7781,N_6605,N_6387);
nor U7782 (N_7782,N_6813,N_7142);
nor U7783 (N_7783,N_7128,N_6529);
or U7784 (N_7784,N_6744,N_6110);
and U7785 (N_7785,N_6688,N_6492);
or U7786 (N_7786,N_6888,N_7199);
nor U7787 (N_7787,N_6760,N_6841);
and U7788 (N_7788,N_7111,N_6498);
or U7789 (N_7789,N_6443,N_6155);
xnor U7790 (N_7790,N_6904,N_6868);
xor U7791 (N_7791,N_6810,N_6074);
nor U7792 (N_7792,N_6937,N_6374);
nand U7793 (N_7793,N_6079,N_6200);
nor U7794 (N_7794,N_6541,N_6193);
nand U7795 (N_7795,N_6502,N_6530);
nor U7796 (N_7796,N_6501,N_7189);
and U7797 (N_7797,N_7122,N_6382);
nor U7798 (N_7798,N_6650,N_6614);
nor U7799 (N_7799,N_7003,N_6765);
nand U7800 (N_7800,N_7056,N_6109);
xnor U7801 (N_7801,N_6486,N_6621);
and U7802 (N_7802,N_6845,N_6899);
or U7803 (N_7803,N_7063,N_6506);
or U7804 (N_7804,N_6503,N_6161);
xor U7805 (N_7805,N_6552,N_6350);
or U7806 (N_7806,N_6405,N_6813);
or U7807 (N_7807,N_7129,N_7066);
nor U7808 (N_7808,N_6768,N_6861);
or U7809 (N_7809,N_7024,N_6191);
or U7810 (N_7810,N_6191,N_6380);
nand U7811 (N_7811,N_7083,N_6312);
xor U7812 (N_7812,N_6607,N_6850);
nor U7813 (N_7813,N_7125,N_6919);
nand U7814 (N_7814,N_6413,N_6183);
nand U7815 (N_7815,N_6551,N_6691);
nor U7816 (N_7816,N_6538,N_7006);
nor U7817 (N_7817,N_6401,N_6218);
xnor U7818 (N_7818,N_6831,N_6238);
nand U7819 (N_7819,N_6114,N_6141);
nor U7820 (N_7820,N_6880,N_6771);
nand U7821 (N_7821,N_6877,N_6855);
xor U7822 (N_7822,N_6562,N_7091);
nand U7823 (N_7823,N_6914,N_7167);
nand U7824 (N_7824,N_6843,N_6299);
nor U7825 (N_7825,N_6820,N_6525);
and U7826 (N_7826,N_6388,N_6057);
nand U7827 (N_7827,N_7104,N_6216);
nand U7828 (N_7828,N_7087,N_6569);
xnor U7829 (N_7829,N_6872,N_6098);
nand U7830 (N_7830,N_6636,N_7086);
nand U7831 (N_7831,N_6138,N_6293);
nor U7832 (N_7832,N_6185,N_6596);
or U7833 (N_7833,N_6200,N_6344);
nand U7834 (N_7834,N_6536,N_6542);
and U7835 (N_7835,N_6318,N_7133);
or U7836 (N_7836,N_6985,N_6185);
nand U7837 (N_7837,N_6328,N_6945);
nand U7838 (N_7838,N_6885,N_6946);
xor U7839 (N_7839,N_6150,N_7035);
nand U7840 (N_7840,N_6754,N_6073);
nand U7841 (N_7841,N_6525,N_6735);
xnor U7842 (N_7842,N_6692,N_6196);
and U7843 (N_7843,N_6036,N_6875);
xnor U7844 (N_7844,N_6606,N_6720);
and U7845 (N_7845,N_6562,N_6240);
or U7846 (N_7846,N_6591,N_6137);
nand U7847 (N_7847,N_7193,N_6953);
xnor U7848 (N_7848,N_6057,N_7165);
nor U7849 (N_7849,N_6028,N_6094);
xor U7850 (N_7850,N_6603,N_6809);
or U7851 (N_7851,N_6886,N_6393);
and U7852 (N_7852,N_6187,N_6005);
nor U7853 (N_7853,N_6595,N_6861);
and U7854 (N_7854,N_6270,N_6100);
nand U7855 (N_7855,N_6707,N_7179);
nand U7856 (N_7856,N_7065,N_6791);
nand U7857 (N_7857,N_6889,N_6611);
or U7858 (N_7858,N_7002,N_6041);
xnor U7859 (N_7859,N_6578,N_7141);
and U7860 (N_7860,N_6413,N_6978);
and U7861 (N_7861,N_6829,N_6308);
and U7862 (N_7862,N_6257,N_6706);
and U7863 (N_7863,N_6292,N_6389);
and U7864 (N_7864,N_6517,N_6191);
nor U7865 (N_7865,N_6326,N_6181);
xor U7866 (N_7866,N_7154,N_6430);
nor U7867 (N_7867,N_6595,N_6893);
xor U7868 (N_7868,N_7039,N_6113);
nor U7869 (N_7869,N_6540,N_6902);
and U7870 (N_7870,N_6152,N_7025);
or U7871 (N_7871,N_6508,N_6318);
nor U7872 (N_7872,N_6683,N_7159);
and U7873 (N_7873,N_6814,N_6523);
nor U7874 (N_7874,N_7043,N_6786);
nand U7875 (N_7875,N_6176,N_6052);
nand U7876 (N_7876,N_6632,N_6637);
xor U7877 (N_7877,N_7109,N_6482);
nand U7878 (N_7878,N_6319,N_6659);
nand U7879 (N_7879,N_6164,N_7052);
and U7880 (N_7880,N_7091,N_7130);
and U7881 (N_7881,N_6261,N_6847);
and U7882 (N_7882,N_6364,N_6594);
xor U7883 (N_7883,N_6392,N_7125);
xor U7884 (N_7884,N_6066,N_6710);
xor U7885 (N_7885,N_6500,N_6435);
nand U7886 (N_7886,N_6135,N_6625);
and U7887 (N_7887,N_7001,N_6562);
or U7888 (N_7888,N_6272,N_6053);
nor U7889 (N_7889,N_6906,N_6426);
xnor U7890 (N_7890,N_6975,N_6783);
nand U7891 (N_7891,N_6479,N_7164);
or U7892 (N_7892,N_6403,N_6578);
xor U7893 (N_7893,N_6521,N_6846);
nor U7894 (N_7894,N_6615,N_7000);
nand U7895 (N_7895,N_6172,N_6904);
and U7896 (N_7896,N_7094,N_6578);
nor U7897 (N_7897,N_6267,N_6598);
or U7898 (N_7898,N_6197,N_6801);
and U7899 (N_7899,N_7193,N_6991);
or U7900 (N_7900,N_6326,N_6388);
and U7901 (N_7901,N_6575,N_6779);
xnor U7902 (N_7902,N_6861,N_6451);
nor U7903 (N_7903,N_6598,N_6248);
or U7904 (N_7904,N_6533,N_7199);
or U7905 (N_7905,N_6915,N_7011);
xnor U7906 (N_7906,N_6908,N_7131);
xnor U7907 (N_7907,N_6140,N_6604);
or U7908 (N_7908,N_6314,N_6827);
nor U7909 (N_7909,N_6780,N_6641);
or U7910 (N_7910,N_6500,N_6258);
and U7911 (N_7911,N_6233,N_7045);
and U7912 (N_7912,N_6218,N_6329);
and U7913 (N_7913,N_6087,N_6465);
nand U7914 (N_7914,N_7191,N_7067);
and U7915 (N_7915,N_6343,N_6218);
nor U7916 (N_7916,N_6956,N_6944);
or U7917 (N_7917,N_6544,N_6845);
nor U7918 (N_7918,N_6189,N_6805);
nand U7919 (N_7919,N_6340,N_6457);
and U7920 (N_7920,N_6245,N_6775);
nor U7921 (N_7921,N_6111,N_6606);
xnor U7922 (N_7922,N_6115,N_7004);
nand U7923 (N_7923,N_6916,N_6001);
and U7924 (N_7924,N_6919,N_6952);
xor U7925 (N_7925,N_6705,N_7060);
nor U7926 (N_7926,N_6469,N_6115);
and U7927 (N_7927,N_6875,N_6356);
nand U7928 (N_7928,N_6200,N_6902);
or U7929 (N_7929,N_6529,N_7058);
or U7930 (N_7930,N_6812,N_6841);
nand U7931 (N_7931,N_6601,N_6394);
or U7932 (N_7932,N_7078,N_6437);
nand U7933 (N_7933,N_7100,N_6093);
and U7934 (N_7934,N_6537,N_6264);
xor U7935 (N_7935,N_6611,N_6665);
nand U7936 (N_7936,N_6666,N_6500);
nor U7937 (N_7937,N_6989,N_6453);
nand U7938 (N_7938,N_6324,N_6397);
xnor U7939 (N_7939,N_6738,N_6602);
and U7940 (N_7940,N_6819,N_6767);
nor U7941 (N_7941,N_6093,N_6005);
or U7942 (N_7942,N_7046,N_6786);
or U7943 (N_7943,N_6931,N_6811);
xor U7944 (N_7944,N_6012,N_6028);
or U7945 (N_7945,N_6171,N_6547);
or U7946 (N_7946,N_6749,N_6386);
nand U7947 (N_7947,N_6185,N_6530);
nor U7948 (N_7948,N_6197,N_6697);
and U7949 (N_7949,N_6403,N_6547);
nor U7950 (N_7950,N_6346,N_7168);
nor U7951 (N_7951,N_6743,N_6544);
and U7952 (N_7952,N_7124,N_6533);
nand U7953 (N_7953,N_6557,N_6546);
or U7954 (N_7954,N_7141,N_6590);
or U7955 (N_7955,N_6075,N_6256);
xor U7956 (N_7956,N_7183,N_6067);
or U7957 (N_7957,N_6342,N_6190);
xor U7958 (N_7958,N_6613,N_6250);
and U7959 (N_7959,N_7094,N_6265);
nand U7960 (N_7960,N_6004,N_6342);
or U7961 (N_7961,N_6451,N_6037);
nor U7962 (N_7962,N_6705,N_6266);
nor U7963 (N_7963,N_7047,N_6684);
or U7964 (N_7964,N_6199,N_6379);
xor U7965 (N_7965,N_6786,N_6928);
nand U7966 (N_7966,N_6764,N_6986);
xor U7967 (N_7967,N_7078,N_6942);
xor U7968 (N_7968,N_7088,N_6794);
nand U7969 (N_7969,N_6687,N_6709);
xor U7970 (N_7970,N_6898,N_6901);
or U7971 (N_7971,N_6627,N_7149);
nand U7972 (N_7972,N_6754,N_6436);
nor U7973 (N_7973,N_7150,N_6292);
nand U7974 (N_7974,N_6290,N_6664);
and U7975 (N_7975,N_6167,N_7166);
nand U7976 (N_7976,N_6217,N_6870);
nor U7977 (N_7977,N_6016,N_6859);
nand U7978 (N_7978,N_7144,N_7051);
nand U7979 (N_7979,N_6720,N_6028);
nor U7980 (N_7980,N_6752,N_6123);
and U7981 (N_7981,N_6399,N_6858);
or U7982 (N_7982,N_7193,N_6637);
xor U7983 (N_7983,N_6189,N_7149);
and U7984 (N_7984,N_6323,N_6717);
nand U7985 (N_7985,N_7178,N_6408);
nor U7986 (N_7986,N_6642,N_6173);
nand U7987 (N_7987,N_6141,N_6085);
nand U7988 (N_7988,N_6783,N_6966);
or U7989 (N_7989,N_6236,N_6903);
nor U7990 (N_7990,N_6459,N_6046);
nand U7991 (N_7991,N_6590,N_6250);
nor U7992 (N_7992,N_6702,N_7006);
nor U7993 (N_7993,N_7091,N_7027);
nor U7994 (N_7994,N_6491,N_6627);
and U7995 (N_7995,N_7071,N_6980);
and U7996 (N_7996,N_6369,N_6404);
xnor U7997 (N_7997,N_6117,N_6378);
or U7998 (N_7998,N_6425,N_6796);
and U7999 (N_7999,N_6234,N_6572);
nand U8000 (N_8000,N_6528,N_6559);
xnor U8001 (N_8001,N_6175,N_6183);
xnor U8002 (N_8002,N_7116,N_7097);
or U8003 (N_8003,N_6490,N_6693);
or U8004 (N_8004,N_6999,N_7124);
or U8005 (N_8005,N_7102,N_6825);
xor U8006 (N_8006,N_6944,N_6322);
nand U8007 (N_8007,N_6016,N_6248);
and U8008 (N_8008,N_7162,N_7041);
nor U8009 (N_8009,N_6657,N_7004);
nor U8010 (N_8010,N_6949,N_6395);
xor U8011 (N_8011,N_6829,N_6289);
nor U8012 (N_8012,N_6477,N_6242);
xnor U8013 (N_8013,N_6448,N_6204);
nor U8014 (N_8014,N_6779,N_6337);
and U8015 (N_8015,N_6771,N_6955);
nand U8016 (N_8016,N_7114,N_6527);
nor U8017 (N_8017,N_6890,N_6844);
nor U8018 (N_8018,N_6688,N_6839);
or U8019 (N_8019,N_6193,N_6862);
nand U8020 (N_8020,N_6087,N_6999);
nor U8021 (N_8021,N_6538,N_6123);
or U8022 (N_8022,N_6323,N_7149);
or U8023 (N_8023,N_6404,N_6560);
xnor U8024 (N_8024,N_7049,N_6811);
nor U8025 (N_8025,N_6309,N_6433);
and U8026 (N_8026,N_6903,N_6723);
or U8027 (N_8027,N_6305,N_7061);
or U8028 (N_8028,N_6283,N_6844);
xnor U8029 (N_8029,N_7178,N_7040);
or U8030 (N_8030,N_6761,N_6743);
nor U8031 (N_8031,N_7098,N_6249);
xnor U8032 (N_8032,N_6643,N_6115);
and U8033 (N_8033,N_6730,N_7154);
or U8034 (N_8034,N_6182,N_7040);
nand U8035 (N_8035,N_7090,N_7097);
or U8036 (N_8036,N_7043,N_6262);
and U8037 (N_8037,N_6411,N_6384);
nor U8038 (N_8038,N_6612,N_7057);
or U8039 (N_8039,N_6313,N_6206);
or U8040 (N_8040,N_7000,N_6864);
or U8041 (N_8041,N_6584,N_6459);
or U8042 (N_8042,N_6240,N_6852);
nand U8043 (N_8043,N_6596,N_6028);
and U8044 (N_8044,N_6606,N_6618);
nor U8045 (N_8045,N_6944,N_6631);
nor U8046 (N_8046,N_6061,N_6325);
nand U8047 (N_8047,N_6786,N_6853);
and U8048 (N_8048,N_6310,N_6845);
xnor U8049 (N_8049,N_6645,N_7150);
and U8050 (N_8050,N_6383,N_6487);
or U8051 (N_8051,N_7084,N_6547);
nor U8052 (N_8052,N_6086,N_6982);
nor U8053 (N_8053,N_6243,N_6965);
nand U8054 (N_8054,N_6007,N_6628);
or U8055 (N_8055,N_7010,N_6548);
nand U8056 (N_8056,N_6203,N_6421);
nand U8057 (N_8057,N_6181,N_6677);
xor U8058 (N_8058,N_6940,N_6291);
or U8059 (N_8059,N_7000,N_6932);
nor U8060 (N_8060,N_6104,N_6119);
nand U8061 (N_8061,N_6154,N_6890);
or U8062 (N_8062,N_6710,N_7063);
and U8063 (N_8063,N_6121,N_7054);
nand U8064 (N_8064,N_6069,N_6490);
nor U8065 (N_8065,N_6000,N_6382);
nand U8066 (N_8066,N_7006,N_6659);
and U8067 (N_8067,N_6082,N_6328);
nand U8068 (N_8068,N_6469,N_6134);
or U8069 (N_8069,N_7131,N_6204);
nand U8070 (N_8070,N_6442,N_6292);
nor U8071 (N_8071,N_6569,N_7142);
and U8072 (N_8072,N_6205,N_7031);
or U8073 (N_8073,N_6677,N_6241);
nand U8074 (N_8074,N_6653,N_6756);
nor U8075 (N_8075,N_6310,N_7007);
and U8076 (N_8076,N_6588,N_6342);
xnor U8077 (N_8077,N_6205,N_6654);
or U8078 (N_8078,N_6114,N_6208);
nor U8079 (N_8079,N_6934,N_6545);
and U8080 (N_8080,N_6541,N_6133);
and U8081 (N_8081,N_6414,N_7084);
xor U8082 (N_8082,N_6559,N_6312);
and U8083 (N_8083,N_6890,N_6989);
nor U8084 (N_8084,N_6846,N_6814);
or U8085 (N_8085,N_6712,N_6013);
and U8086 (N_8086,N_6764,N_6125);
and U8087 (N_8087,N_6716,N_6501);
nor U8088 (N_8088,N_6245,N_6884);
nor U8089 (N_8089,N_6252,N_6451);
and U8090 (N_8090,N_6317,N_6125);
nand U8091 (N_8091,N_7106,N_6709);
or U8092 (N_8092,N_6627,N_6270);
nand U8093 (N_8093,N_6773,N_6992);
and U8094 (N_8094,N_6935,N_6825);
nand U8095 (N_8095,N_6690,N_7021);
and U8096 (N_8096,N_6281,N_6257);
nor U8097 (N_8097,N_6773,N_6336);
nor U8098 (N_8098,N_6184,N_6590);
xnor U8099 (N_8099,N_6232,N_7191);
or U8100 (N_8100,N_6405,N_6056);
xor U8101 (N_8101,N_6693,N_6704);
xor U8102 (N_8102,N_7045,N_6478);
and U8103 (N_8103,N_7035,N_6891);
nand U8104 (N_8104,N_6478,N_6359);
nor U8105 (N_8105,N_6497,N_6167);
xor U8106 (N_8106,N_6283,N_6400);
or U8107 (N_8107,N_6223,N_7030);
nor U8108 (N_8108,N_6878,N_6074);
nor U8109 (N_8109,N_6008,N_6509);
or U8110 (N_8110,N_6997,N_6807);
xnor U8111 (N_8111,N_6155,N_6103);
and U8112 (N_8112,N_6012,N_6465);
nand U8113 (N_8113,N_6794,N_6370);
xor U8114 (N_8114,N_6259,N_6605);
and U8115 (N_8115,N_6558,N_6131);
xor U8116 (N_8116,N_6774,N_7003);
and U8117 (N_8117,N_6860,N_6556);
or U8118 (N_8118,N_7027,N_7147);
and U8119 (N_8119,N_6856,N_7082);
or U8120 (N_8120,N_6308,N_6917);
xor U8121 (N_8121,N_6746,N_6332);
xor U8122 (N_8122,N_7107,N_6918);
and U8123 (N_8123,N_6682,N_6958);
nor U8124 (N_8124,N_6970,N_7170);
or U8125 (N_8125,N_7188,N_6138);
or U8126 (N_8126,N_6008,N_6595);
or U8127 (N_8127,N_6560,N_6237);
xnor U8128 (N_8128,N_7153,N_6880);
or U8129 (N_8129,N_6876,N_6711);
or U8130 (N_8130,N_6005,N_6204);
xor U8131 (N_8131,N_7099,N_7041);
and U8132 (N_8132,N_6890,N_7139);
nor U8133 (N_8133,N_6314,N_7138);
and U8134 (N_8134,N_6160,N_6363);
nor U8135 (N_8135,N_6926,N_7150);
nand U8136 (N_8136,N_6587,N_6498);
or U8137 (N_8137,N_6487,N_6885);
xor U8138 (N_8138,N_6964,N_6085);
xnor U8139 (N_8139,N_6526,N_7039);
nand U8140 (N_8140,N_6562,N_6151);
or U8141 (N_8141,N_6646,N_6373);
nand U8142 (N_8142,N_6635,N_6510);
and U8143 (N_8143,N_6754,N_6555);
xnor U8144 (N_8144,N_7017,N_6258);
or U8145 (N_8145,N_6920,N_7184);
nor U8146 (N_8146,N_6164,N_6847);
nand U8147 (N_8147,N_6548,N_6863);
xnor U8148 (N_8148,N_6879,N_6460);
or U8149 (N_8149,N_6684,N_6851);
nand U8150 (N_8150,N_7065,N_6051);
nand U8151 (N_8151,N_6295,N_6756);
xnor U8152 (N_8152,N_6022,N_7125);
or U8153 (N_8153,N_6193,N_6927);
nand U8154 (N_8154,N_6716,N_6736);
nor U8155 (N_8155,N_6874,N_6771);
nand U8156 (N_8156,N_7000,N_6290);
xor U8157 (N_8157,N_7120,N_6171);
xnor U8158 (N_8158,N_6901,N_6979);
nor U8159 (N_8159,N_6992,N_7137);
or U8160 (N_8160,N_6843,N_6914);
nor U8161 (N_8161,N_6369,N_6111);
nor U8162 (N_8162,N_6105,N_6024);
or U8163 (N_8163,N_6059,N_6008);
nand U8164 (N_8164,N_6495,N_6248);
nand U8165 (N_8165,N_7038,N_6888);
nand U8166 (N_8166,N_6350,N_6070);
or U8167 (N_8167,N_6016,N_6387);
or U8168 (N_8168,N_7140,N_6326);
nor U8169 (N_8169,N_6346,N_6378);
nand U8170 (N_8170,N_6822,N_6618);
nand U8171 (N_8171,N_6989,N_7105);
nand U8172 (N_8172,N_6255,N_7132);
or U8173 (N_8173,N_6624,N_7078);
nand U8174 (N_8174,N_6553,N_6026);
and U8175 (N_8175,N_6163,N_6093);
nand U8176 (N_8176,N_6057,N_6826);
nand U8177 (N_8177,N_6157,N_6208);
xor U8178 (N_8178,N_6891,N_6940);
xnor U8179 (N_8179,N_6709,N_6746);
and U8180 (N_8180,N_6738,N_6991);
or U8181 (N_8181,N_6905,N_6699);
and U8182 (N_8182,N_6372,N_6108);
or U8183 (N_8183,N_6657,N_6230);
nand U8184 (N_8184,N_6542,N_6223);
or U8185 (N_8185,N_6376,N_6844);
nor U8186 (N_8186,N_6796,N_7165);
xnor U8187 (N_8187,N_6346,N_6668);
xnor U8188 (N_8188,N_6568,N_6375);
xnor U8189 (N_8189,N_6164,N_6501);
nor U8190 (N_8190,N_7100,N_7049);
xnor U8191 (N_8191,N_6333,N_6460);
or U8192 (N_8192,N_7071,N_6556);
or U8193 (N_8193,N_6414,N_6869);
nand U8194 (N_8194,N_6501,N_6181);
nand U8195 (N_8195,N_6395,N_6268);
nand U8196 (N_8196,N_6395,N_6292);
nand U8197 (N_8197,N_6319,N_6622);
nand U8198 (N_8198,N_6772,N_6251);
and U8199 (N_8199,N_6759,N_6483);
nor U8200 (N_8200,N_6176,N_6570);
or U8201 (N_8201,N_6100,N_6813);
or U8202 (N_8202,N_7045,N_6220);
and U8203 (N_8203,N_6260,N_6455);
xnor U8204 (N_8204,N_7145,N_6063);
xnor U8205 (N_8205,N_6275,N_6612);
or U8206 (N_8206,N_6391,N_6403);
nor U8207 (N_8207,N_6991,N_6378);
nand U8208 (N_8208,N_6327,N_6972);
nand U8209 (N_8209,N_7050,N_6003);
nand U8210 (N_8210,N_6870,N_7031);
nand U8211 (N_8211,N_6445,N_7110);
nor U8212 (N_8212,N_6103,N_7041);
or U8213 (N_8213,N_6081,N_6955);
or U8214 (N_8214,N_6452,N_6662);
xnor U8215 (N_8215,N_6947,N_6340);
or U8216 (N_8216,N_6892,N_6327);
and U8217 (N_8217,N_7151,N_6125);
nor U8218 (N_8218,N_6736,N_6215);
nand U8219 (N_8219,N_6553,N_6994);
nor U8220 (N_8220,N_7054,N_7133);
or U8221 (N_8221,N_6059,N_7002);
xor U8222 (N_8222,N_6718,N_6703);
and U8223 (N_8223,N_6781,N_7152);
xor U8224 (N_8224,N_6505,N_6474);
nand U8225 (N_8225,N_6390,N_6210);
nand U8226 (N_8226,N_6494,N_6955);
or U8227 (N_8227,N_6373,N_6695);
xor U8228 (N_8228,N_7111,N_6973);
nor U8229 (N_8229,N_6966,N_7180);
nand U8230 (N_8230,N_7106,N_6106);
and U8231 (N_8231,N_6117,N_6347);
nand U8232 (N_8232,N_6384,N_6689);
or U8233 (N_8233,N_6032,N_6462);
or U8234 (N_8234,N_6433,N_6965);
nand U8235 (N_8235,N_6394,N_6450);
nor U8236 (N_8236,N_6297,N_6952);
nor U8237 (N_8237,N_6895,N_7111);
or U8238 (N_8238,N_7174,N_7108);
nand U8239 (N_8239,N_7052,N_6917);
and U8240 (N_8240,N_6080,N_6550);
and U8241 (N_8241,N_6871,N_6572);
or U8242 (N_8242,N_6679,N_7142);
nand U8243 (N_8243,N_6122,N_6850);
xor U8244 (N_8244,N_6862,N_6777);
nand U8245 (N_8245,N_6360,N_6064);
nor U8246 (N_8246,N_6745,N_6874);
nand U8247 (N_8247,N_6765,N_6284);
xor U8248 (N_8248,N_6798,N_6548);
xor U8249 (N_8249,N_6215,N_6792);
or U8250 (N_8250,N_6867,N_6304);
nand U8251 (N_8251,N_6439,N_6518);
nor U8252 (N_8252,N_7168,N_6532);
nor U8253 (N_8253,N_6248,N_6229);
and U8254 (N_8254,N_6491,N_7156);
and U8255 (N_8255,N_6478,N_6633);
or U8256 (N_8256,N_7172,N_7094);
and U8257 (N_8257,N_6528,N_6429);
nor U8258 (N_8258,N_6440,N_6509);
and U8259 (N_8259,N_6656,N_6591);
nor U8260 (N_8260,N_6672,N_6415);
nor U8261 (N_8261,N_6833,N_6901);
xor U8262 (N_8262,N_6962,N_6877);
or U8263 (N_8263,N_6028,N_6984);
nor U8264 (N_8264,N_6574,N_6638);
nor U8265 (N_8265,N_6451,N_6407);
xor U8266 (N_8266,N_7101,N_6564);
and U8267 (N_8267,N_6684,N_6007);
xnor U8268 (N_8268,N_6126,N_6811);
and U8269 (N_8269,N_6683,N_6119);
nor U8270 (N_8270,N_6889,N_7157);
and U8271 (N_8271,N_6995,N_6212);
nor U8272 (N_8272,N_7156,N_6321);
nand U8273 (N_8273,N_7178,N_7137);
xnor U8274 (N_8274,N_6658,N_7152);
or U8275 (N_8275,N_6148,N_6593);
nand U8276 (N_8276,N_6034,N_6937);
xor U8277 (N_8277,N_6958,N_7069);
nor U8278 (N_8278,N_6460,N_6880);
nor U8279 (N_8279,N_7199,N_6499);
nor U8280 (N_8280,N_6436,N_6955);
nor U8281 (N_8281,N_6150,N_6942);
nand U8282 (N_8282,N_6711,N_6260);
nor U8283 (N_8283,N_6632,N_6389);
nor U8284 (N_8284,N_6582,N_6439);
or U8285 (N_8285,N_6548,N_7162);
nand U8286 (N_8286,N_6642,N_6961);
or U8287 (N_8287,N_6646,N_6902);
xnor U8288 (N_8288,N_6149,N_6635);
nor U8289 (N_8289,N_6262,N_6832);
nor U8290 (N_8290,N_7104,N_7020);
and U8291 (N_8291,N_6358,N_6250);
nor U8292 (N_8292,N_6653,N_6514);
or U8293 (N_8293,N_6597,N_6463);
nand U8294 (N_8294,N_6787,N_6183);
nor U8295 (N_8295,N_6114,N_6561);
xnor U8296 (N_8296,N_6830,N_6239);
or U8297 (N_8297,N_6908,N_6940);
nor U8298 (N_8298,N_6009,N_6051);
and U8299 (N_8299,N_6141,N_7095);
or U8300 (N_8300,N_6449,N_6150);
xor U8301 (N_8301,N_6016,N_6701);
nor U8302 (N_8302,N_6111,N_6151);
or U8303 (N_8303,N_6635,N_6143);
nand U8304 (N_8304,N_6686,N_7135);
nand U8305 (N_8305,N_7169,N_6939);
nand U8306 (N_8306,N_6409,N_6381);
nand U8307 (N_8307,N_7085,N_6339);
xnor U8308 (N_8308,N_6104,N_6135);
xor U8309 (N_8309,N_6102,N_6199);
or U8310 (N_8310,N_6383,N_6035);
xnor U8311 (N_8311,N_6221,N_7006);
xor U8312 (N_8312,N_6647,N_6608);
nand U8313 (N_8313,N_6004,N_7161);
nand U8314 (N_8314,N_6561,N_7176);
nor U8315 (N_8315,N_6279,N_6872);
or U8316 (N_8316,N_6681,N_6705);
and U8317 (N_8317,N_7122,N_6434);
xor U8318 (N_8318,N_6913,N_6832);
or U8319 (N_8319,N_6096,N_6277);
or U8320 (N_8320,N_6283,N_6998);
nor U8321 (N_8321,N_6097,N_6195);
and U8322 (N_8322,N_6143,N_6638);
nor U8323 (N_8323,N_6233,N_7128);
xnor U8324 (N_8324,N_6433,N_6119);
xor U8325 (N_8325,N_6702,N_6360);
and U8326 (N_8326,N_7096,N_6887);
and U8327 (N_8327,N_6634,N_6984);
xor U8328 (N_8328,N_6542,N_7168);
and U8329 (N_8329,N_6289,N_6871);
and U8330 (N_8330,N_6502,N_6682);
xnor U8331 (N_8331,N_6572,N_6376);
xor U8332 (N_8332,N_7025,N_7107);
and U8333 (N_8333,N_6163,N_6304);
nor U8334 (N_8334,N_6586,N_7058);
nor U8335 (N_8335,N_6623,N_6539);
nor U8336 (N_8336,N_6955,N_6208);
and U8337 (N_8337,N_6636,N_6104);
nor U8338 (N_8338,N_6948,N_7156);
and U8339 (N_8339,N_6538,N_6687);
and U8340 (N_8340,N_6560,N_7112);
and U8341 (N_8341,N_6599,N_6103);
and U8342 (N_8342,N_6470,N_6440);
and U8343 (N_8343,N_7182,N_6892);
or U8344 (N_8344,N_6727,N_6930);
or U8345 (N_8345,N_6074,N_6280);
xnor U8346 (N_8346,N_6738,N_6037);
xnor U8347 (N_8347,N_6941,N_6139);
nand U8348 (N_8348,N_6629,N_6033);
nor U8349 (N_8349,N_6749,N_7043);
nand U8350 (N_8350,N_6604,N_6798);
nand U8351 (N_8351,N_6732,N_6121);
nor U8352 (N_8352,N_6979,N_6747);
xor U8353 (N_8353,N_6516,N_6386);
and U8354 (N_8354,N_6522,N_6591);
or U8355 (N_8355,N_7109,N_6635);
and U8356 (N_8356,N_6876,N_7115);
or U8357 (N_8357,N_6153,N_6248);
or U8358 (N_8358,N_7022,N_6349);
and U8359 (N_8359,N_6034,N_6493);
or U8360 (N_8360,N_6119,N_6207);
or U8361 (N_8361,N_6463,N_6167);
and U8362 (N_8362,N_6994,N_6498);
and U8363 (N_8363,N_6688,N_6372);
xnor U8364 (N_8364,N_6220,N_6704);
and U8365 (N_8365,N_6179,N_6524);
nand U8366 (N_8366,N_7117,N_6813);
and U8367 (N_8367,N_6838,N_7185);
and U8368 (N_8368,N_6454,N_7168);
xor U8369 (N_8369,N_6533,N_6833);
and U8370 (N_8370,N_6119,N_6459);
or U8371 (N_8371,N_6994,N_6270);
or U8372 (N_8372,N_6805,N_6065);
or U8373 (N_8373,N_6228,N_6888);
nand U8374 (N_8374,N_6082,N_6578);
and U8375 (N_8375,N_6491,N_6220);
and U8376 (N_8376,N_6106,N_7153);
and U8377 (N_8377,N_7082,N_6602);
nor U8378 (N_8378,N_6063,N_6640);
nor U8379 (N_8379,N_6671,N_6737);
nor U8380 (N_8380,N_6885,N_6983);
nand U8381 (N_8381,N_6692,N_7046);
and U8382 (N_8382,N_6097,N_6098);
and U8383 (N_8383,N_6744,N_6421);
xnor U8384 (N_8384,N_6226,N_7072);
and U8385 (N_8385,N_6345,N_6625);
and U8386 (N_8386,N_6580,N_6577);
and U8387 (N_8387,N_7119,N_6735);
or U8388 (N_8388,N_6320,N_6058);
and U8389 (N_8389,N_7120,N_6264);
nand U8390 (N_8390,N_6429,N_6362);
or U8391 (N_8391,N_6441,N_6345);
nor U8392 (N_8392,N_6702,N_6157);
or U8393 (N_8393,N_6404,N_6744);
or U8394 (N_8394,N_6545,N_6974);
or U8395 (N_8395,N_6265,N_7067);
xnor U8396 (N_8396,N_6876,N_6407);
nand U8397 (N_8397,N_7141,N_6320);
xnor U8398 (N_8398,N_6829,N_6165);
nand U8399 (N_8399,N_6037,N_6481);
and U8400 (N_8400,N_8010,N_7243);
xor U8401 (N_8401,N_7852,N_7233);
and U8402 (N_8402,N_7334,N_7426);
xnor U8403 (N_8403,N_8351,N_7476);
nor U8404 (N_8404,N_7752,N_7326);
nor U8405 (N_8405,N_7818,N_8395);
nand U8406 (N_8406,N_7435,N_7646);
xor U8407 (N_8407,N_8250,N_7890);
and U8408 (N_8408,N_7493,N_8264);
and U8409 (N_8409,N_8149,N_7430);
and U8410 (N_8410,N_8150,N_8223);
or U8411 (N_8411,N_7912,N_8139);
nor U8412 (N_8412,N_8002,N_8204);
nor U8413 (N_8413,N_7443,N_8369);
xnor U8414 (N_8414,N_8336,N_8231);
or U8415 (N_8415,N_7397,N_8287);
or U8416 (N_8416,N_7717,N_8328);
and U8417 (N_8417,N_7952,N_7774);
or U8418 (N_8418,N_8116,N_8020);
nor U8419 (N_8419,N_7679,N_8105);
or U8420 (N_8420,N_8366,N_7645);
and U8421 (N_8421,N_8153,N_7737);
nand U8422 (N_8422,N_8217,N_7368);
xor U8423 (N_8423,N_8271,N_7467);
xnor U8424 (N_8424,N_8243,N_7214);
xor U8425 (N_8425,N_8234,N_7631);
xor U8426 (N_8426,N_7223,N_8205);
nand U8427 (N_8427,N_7358,N_8145);
xnor U8428 (N_8428,N_7515,N_7591);
nor U8429 (N_8429,N_7868,N_7968);
nor U8430 (N_8430,N_7580,N_7786);
nand U8431 (N_8431,N_7880,N_7558);
and U8432 (N_8432,N_8021,N_7290);
and U8433 (N_8433,N_8170,N_8327);
nand U8434 (N_8434,N_7224,N_7696);
or U8435 (N_8435,N_7510,N_7815);
and U8436 (N_8436,N_7716,N_7583);
xor U8437 (N_8437,N_8094,N_8214);
and U8438 (N_8438,N_7913,N_7727);
xnor U8439 (N_8439,N_7825,N_8381);
nand U8440 (N_8440,N_8106,N_7616);
and U8441 (N_8441,N_8386,N_7548);
or U8442 (N_8442,N_7437,N_7947);
nor U8443 (N_8443,N_7915,N_7925);
nor U8444 (N_8444,N_7980,N_7639);
nor U8445 (N_8445,N_7340,N_7565);
nand U8446 (N_8446,N_8087,N_7544);
nor U8447 (N_8447,N_8143,N_7338);
nand U8448 (N_8448,N_7377,N_7601);
or U8449 (N_8449,N_8064,N_7799);
nor U8450 (N_8450,N_7981,N_7628);
or U8451 (N_8451,N_7267,N_8163);
and U8452 (N_8452,N_7919,N_7485);
or U8453 (N_8453,N_7746,N_7330);
or U8454 (N_8454,N_8356,N_7826);
nor U8455 (N_8455,N_8158,N_8229);
nor U8456 (N_8456,N_7865,N_7835);
nand U8457 (N_8457,N_8342,N_7574);
nand U8458 (N_8458,N_8061,N_7230);
nand U8459 (N_8459,N_7823,N_7794);
or U8460 (N_8460,N_7775,N_8049);
nor U8461 (N_8461,N_7692,N_8279);
xnor U8462 (N_8462,N_8341,N_7235);
or U8463 (N_8463,N_7674,N_8398);
nor U8464 (N_8464,N_7201,N_7779);
xor U8465 (N_8465,N_7448,N_8011);
nand U8466 (N_8466,N_7964,N_7948);
xor U8467 (N_8467,N_8117,N_8194);
xor U8468 (N_8468,N_8102,N_7719);
xor U8469 (N_8469,N_8046,N_7380);
nor U8470 (N_8470,N_7879,N_7318);
nand U8471 (N_8471,N_8058,N_7513);
nor U8472 (N_8472,N_7521,N_8224);
or U8473 (N_8473,N_8345,N_7602);
and U8474 (N_8474,N_7975,N_7830);
xor U8475 (N_8475,N_8173,N_8278);
or U8476 (N_8476,N_8182,N_7519);
nor U8477 (N_8477,N_7906,N_7221);
nand U8478 (N_8478,N_8232,N_8384);
nand U8479 (N_8479,N_7884,N_7986);
nor U8480 (N_8480,N_8206,N_7232);
and U8481 (N_8481,N_8000,N_7654);
or U8482 (N_8482,N_8344,N_7572);
nor U8483 (N_8483,N_7262,N_8005);
nand U8484 (N_8484,N_7741,N_7404);
xnor U8485 (N_8485,N_7655,N_7999);
nor U8486 (N_8486,N_7609,N_7263);
nand U8487 (N_8487,N_8315,N_8247);
or U8488 (N_8488,N_8188,N_7789);
and U8489 (N_8489,N_7596,N_8080);
nand U8490 (N_8490,N_7252,N_8245);
nand U8491 (N_8491,N_8195,N_7522);
or U8492 (N_8492,N_8372,N_8165);
and U8493 (N_8493,N_7342,N_7311);
nand U8494 (N_8494,N_8131,N_7759);
nand U8495 (N_8495,N_8036,N_7400);
and U8496 (N_8496,N_8193,N_7289);
nand U8497 (N_8497,N_8374,N_7240);
nand U8498 (N_8498,N_7712,N_7374);
and U8499 (N_8499,N_8083,N_8317);
xnor U8500 (N_8500,N_8082,N_7914);
xnor U8501 (N_8501,N_8110,N_8026);
nor U8502 (N_8502,N_7264,N_7846);
nor U8503 (N_8503,N_7579,N_7511);
nor U8504 (N_8504,N_7216,N_7754);
and U8505 (N_8505,N_8004,N_7926);
nor U8506 (N_8506,N_8112,N_8295);
xnor U8507 (N_8507,N_7545,N_7390);
nor U8508 (N_8508,N_7406,N_8385);
and U8509 (N_8509,N_7635,N_8177);
nand U8510 (N_8510,N_7969,N_7415);
xnor U8511 (N_8511,N_7734,N_7402);
and U8512 (N_8512,N_8147,N_7346);
nor U8513 (N_8513,N_7901,N_8034);
nor U8514 (N_8514,N_7417,N_7623);
xor U8515 (N_8515,N_7489,N_7977);
nor U8516 (N_8516,N_7575,N_7652);
and U8517 (N_8517,N_7502,N_7452);
and U8518 (N_8518,N_8033,N_7682);
xor U8519 (N_8519,N_8009,N_7576);
or U8520 (N_8520,N_7855,N_7806);
nor U8521 (N_8521,N_8339,N_8056);
nand U8522 (N_8522,N_8044,N_7463);
xor U8523 (N_8523,N_7568,N_8126);
nor U8524 (N_8524,N_8246,N_7651);
nor U8525 (N_8525,N_7753,N_8062);
xor U8526 (N_8526,N_7863,N_8274);
nand U8527 (N_8527,N_7496,N_7858);
or U8528 (N_8528,N_8099,N_7625);
and U8529 (N_8529,N_8207,N_7584);
or U8530 (N_8530,N_7622,N_7333);
and U8531 (N_8531,N_7530,N_7399);
and U8532 (N_8532,N_7962,N_7644);
or U8533 (N_8533,N_8171,N_7720);
nand U8534 (N_8534,N_7634,N_7503);
or U8535 (N_8535,N_8164,N_7791);
xor U8536 (N_8536,N_7617,N_7805);
xnor U8537 (N_8537,N_7817,N_7389);
or U8538 (N_8538,N_7292,N_8200);
and U8539 (N_8539,N_7797,N_8294);
nor U8540 (N_8540,N_8226,N_7424);
and U8541 (N_8541,N_7988,N_8065);
nor U8542 (N_8542,N_7219,N_8363);
nor U8543 (N_8543,N_8378,N_8118);
xnor U8544 (N_8544,N_7942,N_8151);
or U8545 (N_8545,N_7577,N_7270);
and U8546 (N_8546,N_8268,N_8031);
nor U8547 (N_8547,N_7328,N_7730);
nand U8548 (N_8548,N_8137,N_7239);
nand U8549 (N_8549,N_7638,N_8035);
xnor U8550 (N_8550,N_7840,N_7362);
xnor U8551 (N_8551,N_7319,N_7889);
xor U8552 (N_8552,N_8290,N_8197);
nor U8553 (N_8553,N_7668,N_7705);
and U8554 (N_8554,N_7841,N_7641);
or U8555 (N_8555,N_7520,N_7896);
nand U8556 (N_8556,N_7765,N_7850);
and U8557 (N_8557,N_7288,N_8376);
nand U8558 (N_8558,N_7353,N_8390);
xor U8559 (N_8559,N_7704,N_8007);
nor U8560 (N_8560,N_7633,N_8267);
or U8561 (N_8561,N_7920,N_8396);
or U8562 (N_8562,N_8138,N_8051);
xor U8563 (N_8563,N_8357,N_8047);
xor U8564 (N_8564,N_8189,N_7409);
nand U8565 (N_8565,N_7516,N_7708);
and U8566 (N_8566,N_8367,N_8235);
or U8567 (N_8567,N_7959,N_7935);
xor U8568 (N_8568,N_8387,N_8054);
nand U8569 (N_8569,N_8330,N_8359);
nand U8570 (N_8570,N_7853,N_7238);
and U8571 (N_8571,N_8043,N_7647);
nand U8572 (N_8572,N_7588,N_7283);
and U8573 (N_8573,N_7801,N_8069);
nor U8574 (N_8574,N_8142,N_7861);
nand U8575 (N_8575,N_7847,N_7594);
or U8576 (N_8576,N_8215,N_7939);
nor U8577 (N_8577,N_7302,N_7608);
nor U8578 (N_8578,N_7563,N_7788);
nor U8579 (N_8579,N_7732,N_7341);
or U8580 (N_8580,N_7758,N_8314);
nand U8581 (N_8581,N_7885,N_7802);
and U8582 (N_8582,N_7698,N_7251);
or U8583 (N_8583,N_8218,N_8275);
or U8584 (N_8584,N_8155,N_7686);
nand U8585 (N_8585,N_7369,N_8018);
xor U8586 (N_8586,N_7688,N_8208);
or U8587 (N_8587,N_8255,N_8300);
xor U8588 (N_8588,N_7281,N_7465);
and U8589 (N_8589,N_7945,N_7294);
or U8590 (N_8590,N_7856,N_7398);
and U8591 (N_8591,N_8213,N_8113);
and U8592 (N_8592,N_7665,N_7446);
and U8593 (N_8593,N_8115,N_7763);
or U8594 (N_8594,N_8225,N_8209);
and U8595 (N_8595,N_7304,N_7836);
or U8596 (N_8596,N_7848,N_8391);
or U8597 (N_8597,N_8329,N_7549);
and U8598 (N_8598,N_7337,N_7748);
xor U8599 (N_8599,N_8183,N_8146);
and U8600 (N_8600,N_7613,N_8172);
nand U8601 (N_8601,N_7672,N_7370);
nor U8602 (N_8602,N_7313,N_8338);
or U8603 (N_8603,N_8281,N_7764);
or U8604 (N_8604,N_7923,N_7383);
nor U8605 (N_8605,N_7680,N_7535);
xor U8606 (N_8606,N_7257,N_8248);
or U8607 (N_8607,N_7250,N_7691);
and U8608 (N_8608,N_7276,N_7882);
or U8609 (N_8609,N_7322,N_7551);
nor U8610 (N_8610,N_7570,N_7436);
nor U8611 (N_8611,N_7490,N_7391);
or U8612 (N_8612,N_7445,N_7562);
or U8613 (N_8613,N_7444,N_7990);
and U8614 (N_8614,N_7771,N_8097);
nand U8615 (N_8615,N_7961,N_7637);
xor U8616 (N_8616,N_7933,N_7321);
xnor U8617 (N_8617,N_7954,N_7903);
or U8618 (N_8618,N_8192,N_7298);
or U8619 (N_8619,N_8124,N_7751);
or U8620 (N_8620,N_7327,N_8201);
nor U8621 (N_8621,N_7643,N_7666);
and U8622 (N_8622,N_7247,N_7357);
xnor U8623 (N_8623,N_7245,N_8060);
nand U8624 (N_8624,N_7405,N_7301);
nor U8625 (N_8625,N_7905,N_8236);
nor U8626 (N_8626,N_8364,N_7600);
xor U8627 (N_8627,N_7208,N_7458);
or U8628 (N_8628,N_7743,N_7331);
and U8629 (N_8629,N_7894,N_7769);
xor U8630 (N_8630,N_7978,N_7897);
and U8631 (N_8631,N_7524,N_7658);
nand U8632 (N_8632,N_8276,N_8070);
nor U8633 (N_8633,N_7735,N_7315);
nand U8634 (N_8634,N_7620,N_7468);
and U8635 (N_8635,N_7356,N_7814);
and U8636 (N_8636,N_8098,N_8383);
or U8637 (N_8637,N_8257,N_7891);
or U8638 (N_8638,N_8100,N_7411);
xor U8639 (N_8639,N_7663,N_8256);
nand U8640 (N_8640,N_7268,N_8240);
nand U8641 (N_8641,N_8340,N_7982);
nand U8642 (N_8642,N_7603,N_7669);
and U8643 (N_8643,N_8350,N_7590);
xor U8644 (N_8644,N_7685,N_8399);
xnor U8645 (N_8645,N_7929,N_8190);
xor U8646 (N_8646,N_7953,N_7361);
nor U8647 (N_8647,N_8230,N_7222);
or U8648 (N_8648,N_7757,N_7494);
and U8649 (N_8649,N_8263,N_7483);
and U8650 (N_8650,N_8128,N_7261);
or U8651 (N_8651,N_8296,N_7550);
nor U8652 (N_8652,N_7248,N_7928);
nand U8653 (N_8653,N_8349,N_7569);
or U8654 (N_8654,N_7957,N_8397);
nor U8655 (N_8655,N_8178,N_7809);
or U8656 (N_8656,N_7607,N_8371);
nand U8657 (N_8657,N_8361,N_7626);
nor U8658 (N_8658,N_7832,N_7320);
or U8659 (N_8659,N_7828,N_7396);
or U8660 (N_8660,N_7225,N_7970);
and U8661 (N_8661,N_8119,N_8085);
or U8662 (N_8662,N_7495,N_7534);
and U8663 (N_8663,N_7618,N_7408);
nor U8664 (N_8664,N_8253,N_7422);
or U8665 (N_8665,N_7994,N_7944);
nor U8666 (N_8666,N_8310,N_7295);
nand U8667 (N_8667,N_7695,N_7810);
or U8668 (N_8668,N_8039,N_7941);
xnor U8669 (N_8669,N_7375,N_8244);
nor U8670 (N_8670,N_7792,N_7481);
or U8671 (N_8671,N_7546,N_7296);
xor U8672 (N_8672,N_8067,N_8259);
or U8673 (N_8673,N_8301,N_7715);
xnor U8674 (N_8674,N_8211,N_8157);
nor U8675 (N_8675,N_7462,N_8283);
xor U8676 (N_8676,N_7833,N_7785);
nand U8677 (N_8677,N_8377,N_7803);
nor U8678 (N_8678,N_8107,N_8071);
or U8679 (N_8679,N_7820,N_7724);
nor U8680 (N_8680,N_8125,N_7456);
and U8681 (N_8681,N_7517,N_8161);
nand U8682 (N_8682,N_7242,N_7536);
nand U8683 (N_8683,N_7471,N_7934);
nand U8684 (N_8684,N_7438,N_7845);
nor U8685 (N_8685,N_7813,N_7203);
nand U8686 (N_8686,N_7450,N_7429);
and U8687 (N_8687,N_7431,N_7834);
nor U8688 (N_8688,N_7960,N_8203);
nand U8689 (N_8689,N_7946,N_7611);
nor U8690 (N_8690,N_7653,N_7610);
nor U8691 (N_8691,N_8261,N_7816);
and U8692 (N_8692,N_8166,N_7269);
nand U8693 (N_8693,N_7425,N_8319);
nand U8694 (N_8694,N_7869,N_8104);
xor U8695 (N_8695,N_8121,N_7469);
xor U8696 (N_8696,N_7472,N_7434);
nor U8697 (N_8697,N_7713,N_7742);
xor U8698 (N_8698,N_7681,N_8003);
and U8699 (N_8699,N_8133,N_7323);
nand U8700 (N_8700,N_8072,N_8324);
or U8701 (N_8701,N_8288,N_7640);
and U8702 (N_8702,N_7287,N_7305);
and U8703 (N_8703,N_7624,N_7683);
xnor U8704 (N_8704,N_7236,N_8265);
and U8705 (N_8705,N_7540,N_8012);
or U8706 (N_8706,N_7687,N_7943);
xor U8707 (N_8707,N_7360,N_7403);
nand U8708 (N_8708,N_7231,N_7266);
xor U8709 (N_8709,N_7526,N_8152);
and U8710 (N_8710,N_7433,N_7987);
nor U8711 (N_8711,N_7755,N_7529);
xor U8712 (N_8712,N_7227,N_7523);
and U8713 (N_8713,N_7366,N_7985);
nand U8714 (N_8714,N_7206,N_7862);
nand U8715 (N_8715,N_8140,N_7386);
xor U8716 (N_8716,N_8291,N_7505);
and U8717 (N_8717,N_7207,N_8318);
nor U8718 (N_8718,N_7782,N_7260);
and U8719 (N_8719,N_7684,N_7678);
nor U8720 (N_8720,N_8202,N_7703);
and U8721 (N_8721,N_7614,N_7778);
nor U8722 (N_8722,N_8284,N_8368);
and U8723 (N_8723,N_7350,N_7297);
and U8724 (N_8724,N_7280,N_7739);
or U8725 (N_8725,N_7992,N_8022);
nand U8726 (N_8726,N_7395,N_7776);
nor U8727 (N_8727,N_8136,N_7597);
xor U8728 (N_8728,N_7899,N_7363);
nor U8729 (N_8729,N_8285,N_7870);
and U8730 (N_8730,N_7420,N_8365);
xnor U8731 (N_8731,N_8347,N_7381);
and U8732 (N_8732,N_8302,N_7228);
xnor U8733 (N_8733,N_8095,N_7694);
nor U8734 (N_8734,N_7744,N_7258);
and U8735 (N_8735,N_7916,N_7722);
nor U8736 (N_8736,N_8008,N_8216);
or U8737 (N_8737,N_7689,N_7930);
and U8738 (N_8738,N_8375,N_7486);
xor U8739 (N_8739,N_7586,N_7325);
and U8740 (N_8740,N_7547,N_7723);
or U8741 (N_8741,N_7567,N_7388);
nor U8742 (N_8742,N_7604,N_7533);
or U8743 (N_8743,N_8059,N_7555);
xnor U8744 (N_8744,N_8027,N_7419);
nand U8745 (N_8745,N_8389,N_8233);
xnor U8746 (N_8746,N_7619,N_7949);
and U8747 (N_8747,N_8186,N_8114);
nor U8748 (N_8748,N_7538,N_8331);
or U8749 (N_8749,N_7854,N_7210);
nand U8750 (N_8750,N_7507,N_7477);
xnor U8751 (N_8751,N_7950,N_8266);
and U8752 (N_8752,N_7780,N_8025);
or U8753 (N_8753,N_7273,N_7367);
nor U8754 (N_8754,N_7667,N_8185);
nand U8755 (N_8755,N_7531,N_8334);
or U8756 (N_8756,N_7385,N_7461);
and U8757 (N_8757,N_7349,N_8196);
and U8758 (N_8758,N_8111,N_7253);
nor U8759 (N_8759,N_7917,N_7976);
xnor U8760 (N_8760,N_7525,N_7829);
nor U8761 (N_8761,N_8014,N_7632);
xnor U8762 (N_8762,N_7621,N_8293);
nor U8763 (N_8763,N_7636,N_7589);
xnor U8764 (N_8764,N_7859,N_7344);
nor U8765 (N_8765,N_7401,N_7895);
xor U8766 (N_8766,N_7766,N_8077);
nor U8767 (N_8767,N_8320,N_7491);
xor U8768 (N_8768,N_7509,N_7747);
nor U8769 (N_8769,N_7745,N_8352);
or U8770 (N_8770,N_7413,N_7571);
nor U8771 (N_8771,N_8198,N_7956);
xnor U8772 (N_8772,N_7598,N_8045);
or U8773 (N_8773,N_7314,N_7442);
nor U8774 (N_8774,N_8313,N_7767);
nor U8775 (N_8775,N_8132,N_8063);
and U8776 (N_8776,N_7343,N_7875);
nor U8777 (N_8777,N_7989,N_7729);
or U8778 (N_8778,N_8237,N_8262);
xor U8779 (N_8779,N_8015,N_7592);
or U8780 (N_8780,N_8006,N_8289);
xor U8781 (N_8781,N_8286,N_7501);
and U8782 (N_8782,N_7254,N_7808);
and U8783 (N_8783,N_7372,N_7499);
nand U8784 (N_8784,N_8129,N_8148);
nor U8785 (N_8785,N_7966,N_7482);
nor U8786 (N_8786,N_7335,N_7587);
or U8787 (N_8787,N_7909,N_8316);
and U8788 (N_8788,N_7710,N_7936);
xor U8789 (N_8789,N_8308,N_7303);
nor U8790 (N_8790,N_8239,N_7428);
xor U8791 (N_8791,N_7821,N_8057);
nand U8792 (N_8792,N_7466,N_7421);
nor U8793 (N_8793,N_7872,N_8272);
nand U8794 (N_8794,N_7721,N_7451);
xnor U8795 (N_8795,N_7373,N_7497);
xnor U8796 (N_8796,N_7874,N_7241);
and U8797 (N_8797,N_7336,N_8013);
xnor U8798 (N_8798,N_7204,N_8269);
or U8799 (N_8799,N_8079,N_7709);
and U8800 (N_8800,N_7365,N_8354);
or U8801 (N_8801,N_7927,N_7642);
or U8802 (N_8802,N_8030,N_7881);
and U8803 (N_8803,N_8122,N_7293);
or U8804 (N_8804,N_7447,N_7807);
nand U8805 (N_8805,N_7931,N_7310);
and U8806 (N_8806,N_7857,N_8362);
or U8807 (N_8807,N_7736,N_7693);
nand U8808 (N_8808,N_7453,N_7629);
nand U8809 (N_8809,N_7898,N_7998);
and U8810 (N_8810,N_7887,N_7279);
or U8811 (N_8811,N_8024,N_8028);
and U8812 (N_8812,N_7518,N_7819);
nor U8813 (N_8813,N_7768,N_7627);
xor U8814 (N_8814,N_8093,N_7811);
or U8815 (N_8815,N_7282,N_8219);
xor U8816 (N_8816,N_7393,N_8311);
or U8817 (N_8817,N_8181,N_7997);
or U8818 (N_8818,N_8144,N_7756);
nor U8819 (N_8819,N_8084,N_7348);
or U8820 (N_8820,N_7559,N_7416);
xor U8821 (N_8821,N_8304,N_8388);
xor U8822 (N_8822,N_8017,N_7205);
xnor U8823 (N_8823,N_7392,N_8029);
nand U8824 (N_8824,N_8041,N_8199);
and U8825 (N_8825,N_8305,N_8343);
and U8826 (N_8826,N_7714,N_7760);
or U8827 (N_8827,N_7886,N_7275);
nand U8828 (N_8828,N_7749,N_7921);
or U8829 (N_8829,N_7506,N_7837);
or U8830 (N_8830,N_7867,N_7527);
and U8831 (N_8831,N_7700,N_7843);
xnor U8832 (N_8832,N_7211,N_7324);
or U8833 (N_8833,N_7552,N_8086);
nor U8834 (N_8834,N_7226,N_8220);
and U8835 (N_8835,N_8123,N_8078);
and U8836 (N_8836,N_7220,N_7384);
and U8837 (N_8837,N_8076,N_7484);
and U8838 (N_8838,N_8169,N_7812);
or U8839 (N_8839,N_7470,N_8242);
xnor U8840 (N_8840,N_7561,N_7697);
nor U8841 (N_8841,N_7371,N_7532);
nor U8842 (N_8842,N_7824,N_7878);
and U8843 (N_8843,N_7439,N_7351);
xnor U8844 (N_8844,N_7539,N_7364);
and U8845 (N_8845,N_8162,N_7475);
and U8846 (N_8846,N_7528,N_8325);
nand U8847 (N_8847,N_7657,N_8038);
and U8848 (N_8848,N_7670,N_7378);
and U8849 (N_8849,N_7738,N_7938);
or U8850 (N_8850,N_7479,N_8221);
nor U8851 (N_8851,N_8252,N_7514);
or U8852 (N_8852,N_8088,N_7649);
or U8853 (N_8853,N_7432,N_7234);
nand U8854 (N_8854,N_7460,N_8273);
and U8855 (N_8855,N_7725,N_7795);
nor U8856 (N_8856,N_7410,N_7873);
nand U8857 (N_8857,N_7664,N_7412);
and U8858 (N_8858,N_7578,N_7553);
and U8859 (N_8859,N_7973,N_7309);
nand U8860 (N_8860,N_8109,N_7783);
nor U8861 (N_8861,N_7822,N_7537);
nor U8862 (N_8862,N_8241,N_7904);
and U8863 (N_8863,N_7307,N_7512);
nand U8864 (N_8864,N_7844,N_8074);
and U8865 (N_8865,N_8360,N_7347);
or U8866 (N_8866,N_8127,N_7849);
xor U8867 (N_8867,N_7265,N_7541);
and U8868 (N_8868,N_7676,N_7556);
or U8869 (N_8869,N_7418,N_7379);
nor U8870 (N_8870,N_7864,N_7492);
nor U8871 (N_8871,N_7441,N_7557);
xor U8872 (N_8872,N_7474,N_7459);
nor U8873 (N_8873,N_7299,N_8306);
nor U8874 (N_8874,N_7427,N_8108);
nor U8875 (N_8875,N_8050,N_8096);
and U8876 (N_8876,N_7661,N_7237);
nor U8877 (N_8877,N_7595,N_8092);
nor U8878 (N_8878,N_7213,N_7259);
nor U8879 (N_8879,N_8270,N_7414);
xor U8880 (N_8880,N_8392,N_7306);
or U8881 (N_8881,N_7246,N_7498);
or U8882 (N_8882,N_8023,N_8073);
xor U8883 (N_8883,N_7718,N_7731);
nor U8884 (N_8884,N_8089,N_8382);
xnor U8885 (N_8885,N_8156,N_8141);
xor U8886 (N_8886,N_8333,N_8380);
nand U8887 (N_8887,N_7773,N_8348);
or U8888 (N_8888,N_8321,N_8249);
or U8889 (N_8889,N_7787,N_7937);
or U8890 (N_8890,N_8309,N_8212);
and U8891 (N_8891,N_7671,N_7883);
and U8892 (N_8892,N_7770,N_7740);
or U8893 (N_8893,N_8322,N_7272);
nor U8894 (N_8894,N_7300,N_7877);
or U8895 (N_8895,N_7394,N_8101);
and U8896 (N_8896,N_7793,N_7317);
and U8897 (N_8897,N_7979,N_7838);
or U8898 (N_8898,N_7728,N_7593);
nor U8899 (N_8899,N_8191,N_7871);
and U8900 (N_8900,N_8258,N_7967);
nand U8901 (N_8901,N_8167,N_7726);
nand U8902 (N_8902,N_7984,N_7706);
xnor U8903 (N_8903,N_8210,N_7648);
nor U8904 (N_8904,N_7339,N_7454);
nor U8905 (N_8905,N_7908,N_8066);
nand U8906 (N_8906,N_7605,N_7542);
xnor U8907 (N_8907,N_8134,N_7229);
nor U8908 (N_8908,N_7893,N_8227);
and U8909 (N_8909,N_8052,N_7345);
nand U8910 (N_8910,N_7478,N_7971);
and U8911 (N_8911,N_7932,N_8251);
nand U8912 (N_8912,N_8135,N_7352);
xnor U8913 (N_8913,N_7662,N_8332);
nor U8914 (N_8914,N_7464,N_8394);
xor U8915 (N_8915,N_7761,N_7831);
nand U8916 (N_8916,N_7993,N_8053);
xor U8917 (N_8917,N_8016,N_7940);
nor U8918 (N_8918,N_7630,N_7271);
or U8919 (N_8919,N_8075,N_7355);
nor U8920 (N_8920,N_7991,N_7200);
xnor U8921 (N_8921,N_7504,N_7907);
and U8922 (N_8922,N_7488,N_7573);
nand U8923 (N_8923,N_8298,N_7291);
xnor U8924 (N_8924,N_7308,N_7202);
and U8925 (N_8925,N_8175,N_7274);
nor U8926 (N_8926,N_7286,N_8393);
or U8927 (N_8927,N_7209,N_7900);
or U8928 (N_8928,N_8154,N_8358);
or U8929 (N_8929,N_7440,N_7800);
nand U8930 (N_8930,N_8335,N_7781);
and U8931 (N_8931,N_8346,N_8184);
and U8932 (N_8932,N_7543,N_7554);
or U8933 (N_8933,N_7382,N_7918);
or U8934 (N_8934,N_8042,N_7455);
xnor U8935 (N_8935,N_7284,N_7612);
nand U8936 (N_8936,N_7839,N_7866);
nor U8937 (N_8937,N_8282,N_7423);
xor U8938 (N_8938,N_7958,N_8297);
or U8939 (N_8939,N_8159,N_7332);
or U8940 (N_8940,N_8120,N_7707);
xnor U8941 (N_8941,N_7701,N_7711);
nand U8942 (N_8942,N_7564,N_7762);
xor U8943 (N_8943,N_8355,N_8055);
and U8944 (N_8944,N_8337,N_7965);
or U8945 (N_8945,N_7256,N_8130);
or U8946 (N_8946,N_7312,N_7508);
and U8947 (N_8947,N_8222,N_7615);
xnor U8948 (N_8948,N_7359,N_7702);
xnor U8949 (N_8949,N_8379,N_7972);
xnor U8950 (N_8950,N_8103,N_7860);
or U8951 (N_8951,N_7656,N_8370);
nor U8952 (N_8952,N_7804,N_8019);
nand U8953 (N_8953,N_7215,N_7902);
or U8954 (N_8954,N_7582,N_8179);
nand U8955 (N_8955,N_7376,N_8323);
or U8956 (N_8956,N_7278,N_7772);
or U8957 (N_8957,N_7750,N_7249);
or U8958 (N_8958,N_7566,N_8040);
or U8959 (N_8959,N_8091,N_7677);
xnor U8960 (N_8960,N_8353,N_8187);
xor U8961 (N_8961,N_7983,N_7212);
nor U8962 (N_8962,N_7244,N_8307);
xnor U8963 (N_8963,N_8312,N_7218);
nand U8964 (N_8964,N_7690,N_7487);
and U8965 (N_8965,N_7354,N_7842);
nand U8966 (N_8966,N_8174,N_7888);
nand U8967 (N_8967,N_7650,N_8037);
nor U8968 (N_8968,N_7996,N_7995);
or U8969 (N_8969,N_7892,N_7285);
nand U8970 (N_8970,N_7798,N_7316);
nor U8971 (N_8971,N_7581,N_7473);
xnor U8972 (N_8972,N_7777,N_7790);
xor U8973 (N_8973,N_7480,N_8303);
and U8974 (N_8974,N_7606,N_8168);
nor U8975 (N_8975,N_8068,N_7827);
nor U8976 (N_8976,N_7449,N_8292);
xnor U8977 (N_8977,N_7673,N_7876);
and U8978 (N_8978,N_7407,N_8228);
and U8979 (N_8979,N_7911,N_7500);
and U8980 (N_8980,N_7329,N_7955);
or U8981 (N_8981,N_8373,N_7974);
xnor U8982 (N_8982,N_7560,N_7255);
xnor U8983 (N_8983,N_8326,N_7922);
or U8984 (N_8984,N_7910,N_7675);
nor U8985 (N_8985,N_7796,N_7733);
and U8986 (N_8986,N_8081,N_8180);
or U8987 (N_8987,N_7699,N_7277);
nor U8988 (N_8988,N_7851,N_8299);
xor U8989 (N_8989,N_7585,N_7963);
nand U8990 (N_8990,N_7659,N_7217);
xor U8991 (N_8991,N_7599,N_8048);
and U8992 (N_8992,N_8277,N_7924);
or U8993 (N_8993,N_7660,N_8001);
xnor U8994 (N_8994,N_8032,N_7951);
xor U8995 (N_8995,N_8280,N_7387);
nand U8996 (N_8996,N_8260,N_8176);
xor U8997 (N_8997,N_8238,N_7457);
nor U8998 (N_8998,N_8254,N_7784);
and U8999 (N_8999,N_8090,N_8160);
nor U9000 (N_9000,N_8222,N_7283);
nor U9001 (N_9001,N_7425,N_7607);
and U9002 (N_9002,N_7607,N_7228);
nand U9003 (N_9003,N_7787,N_7254);
and U9004 (N_9004,N_7914,N_7830);
and U9005 (N_9005,N_8390,N_8266);
and U9006 (N_9006,N_7660,N_8328);
nor U9007 (N_9007,N_7991,N_8024);
xnor U9008 (N_9008,N_7718,N_7535);
and U9009 (N_9009,N_7827,N_7941);
nand U9010 (N_9010,N_7597,N_8355);
nor U9011 (N_9011,N_7301,N_7756);
nand U9012 (N_9012,N_7289,N_8297);
xnor U9013 (N_9013,N_7859,N_7685);
nand U9014 (N_9014,N_8274,N_7412);
nand U9015 (N_9015,N_7342,N_8217);
nand U9016 (N_9016,N_7811,N_7844);
nand U9017 (N_9017,N_7565,N_7419);
or U9018 (N_9018,N_8164,N_7485);
xor U9019 (N_9019,N_7777,N_7721);
nor U9020 (N_9020,N_7500,N_7212);
or U9021 (N_9021,N_7267,N_7971);
nor U9022 (N_9022,N_7443,N_7302);
xor U9023 (N_9023,N_8291,N_7305);
nand U9024 (N_9024,N_8247,N_7835);
and U9025 (N_9025,N_7845,N_7740);
nor U9026 (N_9026,N_7542,N_7251);
and U9027 (N_9027,N_7868,N_7393);
nand U9028 (N_9028,N_7743,N_8165);
xor U9029 (N_9029,N_8171,N_7792);
nand U9030 (N_9030,N_7715,N_8026);
and U9031 (N_9031,N_7909,N_7784);
and U9032 (N_9032,N_7359,N_8328);
nor U9033 (N_9033,N_7652,N_7591);
nand U9034 (N_9034,N_7564,N_7937);
or U9035 (N_9035,N_7314,N_8041);
nand U9036 (N_9036,N_7378,N_7458);
nor U9037 (N_9037,N_7670,N_7436);
and U9038 (N_9038,N_7461,N_7956);
or U9039 (N_9039,N_8308,N_7615);
nor U9040 (N_9040,N_7660,N_7690);
and U9041 (N_9041,N_8354,N_7390);
nor U9042 (N_9042,N_7475,N_8152);
xor U9043 (N_9043,N_7902,N_7418);
nor U9044 (N_9044,N_8105,N_7335);
xor U9045 (N_9045,N_7921,N_7730);
and U9046 (N_9046,N_7441,N_8178);
and U9047 (N_9047,N_8148,N_7974);
and U9048 (N_9048,N_8058,N_7885);
and U9049 (N_9049,N_8127,N_7562);
nand U9050 (N_9050,N_8099,N_7363);
and U9051 (N_9051,N_7887,N_7695);
or U9052 (N_9052,N_8244,N_7477);
xor U9053 (N_9053,N_8123,N_8353);
nor U9054 (N_9054,N_7992,N_8378);
nand U9055 (N_9055,N_8175,N_7573);
nor U9056 (N_9056,N_8159,N_7703);
xnor U9057 (N_9057,N_7785,N_7484);
and U9058 (N_9058,N_7352,N_7788);
nand U9059 (N_9059,N_7623,N_8385);
and U9060 (N_9060,N_7980,N_7796);
and U9061 (N_9061,N_8323,N_7229);
nand U9062 (N_9062,N_8332,N_8384);
and U9063 (N_9063,N_7543,N_7204);
nand U9064 (N_9064,N_7849,N_7310);
nor U9065 (N_9065,N_7367,N_7641);
or U9066 (N_9066,N_7829,N_7583);
nor U9067 (N_9067,N_8081,N_8046);
or U9068 (N_9068,N_8356,N_8303);
or U9069 (N_9069,N_8214,N_7785);
or U9070 (N_9070,N_7634,N_8192);
nor U9071 (N_9071,N_8145,N_7988);
nand U9072 (N_9072,N_8387,N_7876);
nor U9073 (N_9073,N_7334,N_7870);
and U9074 (N_9074,N_8157,N_7325);
nand U9075 (N_9075,N_7604,N_8374);
nand U9076 (N_9076,N_7429,N_8397);
nor U9077 (N_9077,N_7881,N_7245);
nor U9078 (N_9078,N_8200,N_7447);
xnor U9079 (N_9079,N_8080,N_7370);
nor U9080 (N_9080,N_8330,N_8333);
nand U9081 (N_9081,N_7775,N_7225);
and U9082 (N_9082,N_8133,N_8169);
nor U9083 (N_9083,N_7785,N_8226);
or U9084 (N_9084,N_7266,N_7623);
xor U9085 (N_9085,N_7888,N_7339);
nor U9086 (N_9086,N_8287,N_7772);
xnor U9087 (N_9087,N_7859,N_7752);
nor U9088 (N_9088,N_8133,N_8062);
nand U9089 (N_9089,N_8099,N_7972);
nand U9090 (N_9090,N_7996,N_7294);
and U9091 (N_9091,N_7825,N_8266);
nand U9092 (N_9092,N_7937,N_7365);
and U9093 (N_9093,N_7372,N_8377);
xor U9094 (N_9094,N_7877,N_8208);
and U9095 (N_9095,N_7594,N_7932);
nor U9096 (N_9096,N_8344,N_8213);
and U9097 (N_9097,N_7642,N_7863);
nor U9098 (N_9098,N_7895,N_7658);
or U9099 (N_9099,N_8381,N_7268);
and U9100 (N_9100,N_7435,N_7574);
or U9101 (N_9101,N_7549,N_8266);
and U9102 (N_9102,N_7743,N_8347);
and U9103 (N_9103,N_7366,N_8120);
nor U9104 (N_9104,N_7962,N_7636);
nor U9105 (N_9105,N_8308,N_7405);
or U9106 (N_9106,N_7702,N_8141);
and U9107 (N_9107,N_7333,N_7585);
and U9108 (N_9108,N_8002,N_8074);
nand U9109 (N_9109,N_7494,N_7266);
nand U9110 (N_9110,N_8140,N_7442);
nand U9111 (N_9111,N_7384,N_7357);
nand U9112 (N_9112,N_7357,N_8247);
nor U9113 (N_9113,N_8189,N_7620);
and U9114 (N_9114,N_7691,N_8201);
nand U9115 (N_9115,N_8040,N_8395);
nand U9116 (N_9116,N_7923,N_8171);
nand U9117 (N_9117,N_8045,N_7223);
or U9118 (N_9118,N_8076,N_7940);
or U9119 (N_9119,N_8271,N_7254);
nor U9120 (N_9120,N_7323,N_8276);
nor U9121 (N_9121,N_7381,N_7719);
nand U9122 (N_9122,N_8031,N_7677);
and U9123 (N_9123,N_7285,N_8205);
nand U9124 (N_9124,N_8260,N_7803);
and U9125 (N_9125,N_7832,N_7368);
and U9126 (N_9126,N_7536,N_7727);
xnor U9127 (N_9127,N_8160,N_7304);
xnor U9128 (N_9128,N_7547,N_8040);
xor U9129 (N_9129,N_7364,N_7986);
or U9130 (N_9130,N_7411,N_7433);
nand U9131 (N_9131,N_8053,N_8198);
xor U9132 (N_9132,N_7403,N_8337);
and U9133 (N_9133,N_7501,N_8176);
or U9134 (N_9134,N_7782,N_8200);
xor U9135 (N_9135,N_7459,N_7945);
nor U9136 (N_9136,N_8056,N_7947);
and U9137 (N_9137,N_8102,N_7800);
nor U9138 (N_9138,N_8220,N_8122);
nor U9139 (N_9139,N_7281,N_8354);
and U9140 (N_9140,N_7822,N_7459);
or U9141 (N_9141,N_8365,N_7632);
and U9142 (N_9142,N_7834,N_7668);
and U9143 (N_9143,N_8365,N_7236);
or U9144 (N_9144,N_7608,N_7622);
xor U9145 (N_9145,N_8014,N_7459);
xor U9146 (N_9146,N_7645,N_7737);
nand U9147 (N_9147,N_8286,N_7958);
nand U9148 (N_9148,N_7379,N_7244);
nor U9149 (N_9149,N_8138,N_8266);
nor U9150 (N_9150,N_8241,N_7884);
and U9151 (N_9151,N_7896,N_8327);
xnor U9152 (N_9152,N_8103,N_7448);
or U9153 (N_9153,N_7382,N_7446);
or U9154 (N_9154,N_8326,N_7702);
or U9155 (N_9155,N_8059,N_8229);
and U9156 (N_9156,N_8251,N_7516);
or U9157 (N_9157,N_7403,N_7742);
xnor U9158 (N_9158,N_7794,N_7453);
nand U9159 (N_9159,N_7355,N_8001);
xor U9160 (N_9160,N_8293,N_7783);
and U9161 (N_9161,N_7739,N_8027);
nand U9162 (N_9162,N_7584,N_7227);
and U9163 (N_9163,N_7352,N_8150);
nor U9164 (N_9164,N_7809,N_7841);
nor U9165 (N_9165,N_8188,N_8093);
or U9166 (N_9166,N_8205,N_8275);
nor U9167 (N_9167,N_7809,N_7800);
xnor U9168 (N_9168,N_7380,N_7621);
nand U9169 (N_9169,N_7237,N_8059);
and U9170 (N_9170,N_7595,N_7341);
nor U9171 (N_9171,N_7507,N_7789);
nor U9172 (N_9172,N_8212,N_7209);
and U9173 (N_9173,N_7359,N_7937);
nand U9174 (N_9174,N_7275,N_7679);
nor U9175 (N_9175,N_7949,N_8026);
and U9176 (N_9176,N_7957,N_8153);
xnor U9177 (N_9177,N_8191,N_7629);
and U9178 (N_9178,N_7609,N_7539);
nand U9179 (N_9179,N_8023,N_7695);
xnor U9180 (N_9180,N_7950,N_8061);
and U9181 (N_9181,N_7470,N_8308);
nor U9182 (N_9182,N_7566,N_8096);
nor U9183 (N_9183,N_7297,N_7639);
or U9184 (N_9184,N_7263,N_7660);
and U9185 (N_9185,N_7721,N_8031);
or U9186 (N_9186,N_8119,N_7685);
and U9187 (N_9187,N_7900,N_7880);
and U9188 (N_9188,N_8272,N_7529);
or U9189 (N_9189,N_7262,N_8253);
xnor U9190 (N_9190,N_7479,N_7787);
nor U9191 (N_9191,N_8267,N_8159);
nor U9192 (N_9192,N_7288,N_7659);
nand U9193 (N_9193,N_7846,N_7230);
nand U9194 (N_9194,N_8360,N_7626);
and U9195 (N_9195,N_7648,N_7207);
or U9196 (N_9196,N_7908,N_7305);
xnor U9197 (N_9197,N_7735,N_8361);
or U9198 (N_9198,N_7590,N_7730);
xor U9199 (N_9199,N_7649,N_7769);
and U9200 (N_9200,N_7318,N_8243);
xnor U9201 (N_9201,N_7763,N_8270);
or U9202 (N_9202,N_8397,N_7471);
nor U9203 (N_9203,N_7881,N_7607);
xnor U9204 (N_9204,N_8334,N_8188);
nand U9205 (N_9205,N_7549,N_8280);
or U9206 (N_9206,N_7559,N_7701);
nand U9207 (N_9207,N_8057,N_8352);
xor U9208 (N_9208,N_7271,N_7382);
xor U9209 (N_9209,N_8056,N_8024);
or U9210 (N_9210,N_8313,N_7718);
nor U9211 (N_9211,N_8041,N_7919);
nand U9212 (N_9212,N_7698,N_7879);
or U9213 (N_9213,N_7662,N_8092);
nand U9214 (N_9214,N_7455,N_8155);
or U9215 (N_9215,N_7964,N_7755);
nand U9216 (N_9216,N_8143,N_8022);
xnor U9217 (N_9217,N_7522,N_7686);
nand U9218 (N_9218,N_7525,N_7647);
and U9219 (N_9219,N_7722,N_7890);
nor U9220 (N_9220,N_8207,N_8096);
or U9221 (N_9221,N_7911,N_8069);
xnor U9222 (N_9222,N_8375,N_7601);
xor U9223 (N_9223,N_7428,N_7396);
nor U9224 (N_9224,N_8384,N_7850);
nand U9225 (N_9225,N_7733,N_8148);
nand U9226 (N_9226,N_7351,N_7757);
xnor U9227 (N_9227,N_7414,N_8106);
nand U9228 (N_9228,N_7882,N_7657);
and U9229 (N_9229,N_7325,N_7778);
nand U9230 (N_9230,N_7777,N_7379);
or U9231 (N_9231,N_7835,N_7819);
or U9232 (N_9232,N_7353,N_8239);
and U9233 (N_9233,N_8338,N_7901);
xor U9234 (N_9234,N_7880,N_8333);
or U9235 (N_9235,N_7400,N_7275);
xor U9236 (N_9236,N_8300,N_7749);
nor U9237 (N_9237,N_8226,N_7443);
and U9238 (N_9238,N_7299,N_7499);
and U9239 (N_9239,N_7466,N_7778);
and U9240 (N_9240,N_8071,N_7553);
and U9241 (N_9241,N_7402,N_7627);
nor U9242 (N_9242,N_7683,N_8183);
nand U9243 (N_9243,N_7634,N_7853);
or U9244 (N_9244,N_8114,N_7322);
nand U9245 (N_9245,N_8398,N_7241);
and U9246 (N_9246,N_7891,N_7879);
nor U9247 (N_9247,N_8050,N_8042);
and U9248 (N_9248,N_7786,N_7328);
and U9249 (N_9249,N_7879,N_7997);
xnor U9250 (N_9250,N_7598,N_7747);
or U9251 (N_9251,N_7247,N_7396);
or U9252 (N_9252,N_7907,N_7920);
nand U9253 (N_9253,N_8251,N_7879);
and U9254 (N_9254,N_7449,N_7247);
and U9255 (N_9255,N_7350,N_7994);
and U9256 (N_9256,N_7517,N_7898);
nand U9257 (N_9257,N_7820,N_7663);
or U9258 (N_9258,N_7634,N_8326);
nor U9259 (N_9259,N_7579,N_7841);
or U9260 (N_9260,N_7889,N_7413);
xor U9261 (N_9261,N_7239,N_8304);
xnor U9262 (N_9262,N_7904,N_7734);
or U9263 (N_9263,N_8337,N_8193);
xor U9264 (N_9264,N_7433,N_7595);
xor U9265 (N_9265,N_7334,N_8216);
and U9266 (N_9266,N_7330,N_7824);
nand U9267 (N_9267,N_7716,N_8390);
and U9268 (N_9268,N_7246,N_7614);
xnor U9269 (N_9269,N_7765,N_7257);
xor U9270 (N_9270,N_7280,N_7534);
nand U9271 (N_9271,N_7837,N_7858);
nor U9272 (N_9272,N_7277,N_7594);
or U9273 (N_9273,N_8183,N_7664);
and U9274 (N_9274,N_7240,N_7535);
or U9275 (N_9275,N_8213,N_7797);
or U9276 (N_9276,N_7380,N_8081);
nor U9277 (N_9277,N_7901,N_7943);
nand U9278 (N_9278,N_8135,N_7444);
nand U9279 (N_9279,N_8135,N_8235);
nand U9280 (N_9280,N_8145,N_8053);
nand U9281 (N_9281,N_7319,N_7449);
nand U9282 (N_9282,N_7657,N_7517);
and U9283 (N_9283,N_7840,N_8056);
nand U9284 (N_9284,N_7590,N_7530);
nand U9285 (N_9285,N_7975,N_8110);
nor U9286 (N_9286,N_8184,N_7835);
nor U9287 (N_9287,N_7291,N_7276);
or U9288 (N_9288,N_8199,N_8201);
nor U9289 (N_9289,N_7948,N_7714);
xor U9290 (N_9290,N_8048,N_8275);
and U9291 (N_9291,N_8264,N_7573);
and U9292 (N_9292,N_7360,N_7242);
nand U9293 (N_9293,N_7639,N_7915);
nor U9294 (N_9294,N_8102,N_8195);
nor U9295 (N_9295,N_7919,N_8300);
nand U9296 (N_9296,N_7381,N_7236);
nor U9297 (N_9297,N_7651,N_8315);
xor U9298 (N_9298,N_8207,N_7983);
and U9299 (N_9299,N_7898,N_8012);
xor U9300 (N_9300,N_7845,N_8170);
and U9301 (N_9301,N_7794,N_7737);
or U9302 (N_9302,N_7957,N_8200);
nor U9303 (N_9303,N_7337,N_7206);
xnor U9304 (N_9304,N_7248,N_7796);
xor U9305 (N_9305,N_7228,N_7797);
nor U9306 (N_9306,N_8351,N_8281);
or U9307 (N_9307,N_8029,N_7900);
or U9308 (N_9308,N_8374,N_7698);
nor U9309 (N_9309,N_8149,N_8148);
nand U9310 (N_9310,N_8095,N_8318);
or U9311 (N_9311,N_7846,N_8297);
and U9312 (N_9312,N_7587,N_8334);
nor U9313 (N_9313,N_8375,N_8017);
xor U9314 (N_9314,N_7802,N_7485);
nand U9315 (N_9315,N_8318,N_8029);
xnor U9316 (N_9316,N_7434,N_7806);
xnor U9317 (N_9317,N_7678,N_8011);
xnor U9318 (N_9318,N_8368,N_7899);
and U9319 (N_9319,N_8029,N_7442);
xor U9320 (N_9320,N_7538,N_7665);
xnor U9321 (N_9321,N_7340,N_8223);
or U9322 (N_9322,N_8360,N_7526);
and U9323 (N_9323,N_7925,N_8042);
nand U9324 (N_9324,N_7998,N_7908);
nor U9325 (N_9325,N_7215,N_7547);
nor U9326 (N_9326,N_7324,N_7600);
xor U9327 (N_9327,N_7576,N_7634);
and U9328 (N_9328,N_7455,N_7638);
and U9329 (N_9329,N_7514,N_8159);
and U9330 (N_9330,N_7881,N_7893);
nand U9331 (N_9331,N_7829,N_7369);
nand U9332 (N_9332,N_7243,N_8054);
and U9333 (N_9333,N_7925,N_8136);
or U9334 (N_9334,N_7429,N_7334);
xor U9335 (N_9335,N_8134,N_7643);
xor U9336 (N_9336,N_8142,N_7566);
nand U9337 (N_9337,N_8099,N_8318);
nor U9338 (N_9338,N_8188,N_7855);
and U9339 (N_9339,N_7640,N_7217);
or U9340 (N_9340,N_7880,N_7688);
nor U9341 (N_9341,N_8003,N_7485);
xnor U9342 (N_9342,N_7538,N_8369);
xor U9343 (N_9343,N_7904,N_7207);
and U9344 (N_9344,N_7676,N_8006);
nand U9345 (N_9345,N_7392,N_7491);
xor U9346 (N_9346,N_7893,N_7322);
or U9347 (N_9347,N_7331,N_7688);
nor U9348 (N_9348,N_8019,N_8342);
or U9349 (N_9349,N_8236,N_7295);
nor U9350 (N_9350,N_8125,N_8282);
and U9351 (N_9351,N_8388,N_7503);
xnor U9352 (N_9352,N_7289,N_7843);
and U9353 (N_9353,N_7414,N_8095);
nor U9354 (N_9354,N_7889,N_8366);
nand U9355 (N_9355,N_7846,N_7991);
nor U9356 (N_9356,N_8200,N_8256);
nor U9357 (N_9357,N_7420,N_8158);
or U9358 (N_9358,N_7814,N_8227);
and U9359 (N_9359,N_7438,N_7424);
or U9360 (N_9360,N_8295,N_8048);
or U9361 (N_9361,N_7739,N_7975);
nand U9362 (N_9362,N_7722,N_7793);
nand U9363 (N_9363,N_8067,N_8268);
or U9364 (N_9364,N_7570,N_8273);
xor U9365 (N_9365,N_7714,N_8266);
xnor U9366 (N_9366,N_8099,N_7385);
and U9367 (N_9367,N_7721,N_7516);
nor U9368 (N_9368,N_7972,N_7439);
nand U9369 (N_9369,N_7759,N_7603);
nor U9370 (N_9370,N_7438,N_7550);
and U9371 (N_9371,N_8263,N_7784);
and U9372 (N_9372,N_7424,N_7749);
xnor U9373 (N_9373,N_8228,N_8200);
or U9374 (N_9374,N_7915,N_7926);
xnor U9375 (N_9375,N_8258,N_8280);
or U9376 (N_9376,N_7505,N_7723);
or U9377 (N_9377,N_8200,N_7562);
nand U9378 (N_9378,N_7381,N_7307);
or U9379 (N_9379,N_7828,N_8082);
xor U9380 (N_9380,N_7529,N_8179);
or U9381 (N_9381,N_8047,N_7903);
nor U9382 (N_9382,N_7696,N_7908);
nor U9383 (N_9383,N_7910,N_7444);
nor U9384 (N_9384,N_8092,N_7898);
and U9385 (N_9385,N_7998,N_7850);
or U9386 (N_9386,N_8208,N_8137);
nand U9387 (N_9387,N_7259,N_7376);
xor U9388 (N_9388,N_7733,N_8212);
or U9389 (N_9389,N_7566,N_7370);
or U9390 (N_9390,N_8335,N_7480);
xor U9391 (N_9391,N_8397,N_7277);
and U9392 (N_9392,N_7315,N_8286);
nand U9393 (N_9393,N_8184,N_7867);
xor U9394 (N_9394,N_8022,N_7315);
or U9395 (N_9395,N_8377,N_8313);
or U9396 (N_9396,N_8255,N_7864);
xnor U9397 (N_9397,N_7962,N_8245);
xor U9398 (N_9398,N_7487,N_7333);
or U9399 (N_9399,N_8248,N_7730);
nand U9400 (N_9400,N_7437,N_7727);
nor U9401 (N_9401,N_7406,N_8039);
nand U9402 (N_9402,N_8089,N_7990);
or U9403 (N_9403,N_7869,N_8213);
xor U9404 (N_9404,N_7459,N_7856);
nand U9405 (N_9405,N_7797,N_7311);
xor U9406 (N_9406,N_7818,N_7425);
xnor U9407 (N_9407,N_7911,N_8154);
xor U9408 (N_9408,N_7236,N_8057);
xor U9409 (N_9409,N_7766,N_7315);
or U9410 (N_9410,N_7858,N_8356);
or U9411 (N_9411,N_8249,N_7270);
nor U9412 (N_9412,N_7717,N_7366);
xor U9413 (N_9413,N_8072,N_8215);
nand U9414 (N_9414,N_8227,N_8081);
or U9415 (N_9415,N_7352,N_7350);
or U9416 (N_9416,N_7228,N_8044);
nand U9417 (N_9417,N_7578,N_7574);
nor U9418 (N_9418,N_8294,N_7336);
nand U9419 (N_9419,N_8238,N_7867);
or U9420 (N_9420,N_8206,N_7812);
nor U9421 (N_9421,N_8354,N_7949);
xnor U9422 (N_9422,N_8346,N_8198);
nand U9423 (N_9423,N_7294,N_8068);
xor U9424 (N_9424,N_8247,N_7580);
nand U9425 (N_9425,N_7943,N_7703);
nor U9426 (N_9426,N_7382,N_7508);
nor U9427 (N_9427,N_7241,N_7218);
nand U9428 (N_9428,N_7740,N_7646);
nand U9429 (N_9429,N_7746,N_7222);
nor U9430 (N_9430,N_8022,N_8247);
nor U9431 (N_9431,N_7761,N_8345);
or U9432 (N_9432,N_7723,N_8237);
or U9433 (N_9433,N_8002,N_7978);
nand U9434 (N_9434,N_7784,N_7630);
and U9435 (N_9435,N_7346,N_8323);
xnor U9436 (N_9436,N_7432,N_7347);
or U9437 (N_9437,N_8225,N_7312);
nor U9438 (N_9438,N_7264,N_8230);
nor U9439 (N_9439,N_7257,N_7460);
nand U9440 (N_9440,N_7676,N_7455);
and U9441 (N_9441,N_7773,N_8063);
xor U9442 (N_9442,N_7422,N_7419);
or U9443 (N_9443,N_8176,N_7687);
or U9444 (N_9444,N_8119,N_7881);
nor U9445 (N_9445,N_7908,N_7335);
and U9446 (N_9446,N_8324,N_7571);
nor U9447 (N_9447,N_7982,N_7224);
and U9448 (N_9448,N_7247,N_7759);
nand U9449 (N_9449,N_8001,N_7711);
xnor U9450 (N_9450,N_8021,N_8077);
nand U9451 (N_9451,N_8294,N_7772);
nand U9452 (N_9452,N_7442,N_7202);
nand U9453 (N_9453,N_7212,N_8268);
xnor U9454 (N_9454,N_8365,N_8081);
nor U9455 (N_9455,N_7322,N_7859);
xnor U9456 (N_9456,N_7995,N_8343);
or U9457 (N_9457,N_7307,N_7301);
nand U9458 (N_9458,N_8268,N_7283);
nor U9459 (N_9459,N_7301,N_7773);
or U9460 (N_9460,N_7622,N_8299);
nand U9461 (N_9461,N_7861,N_7712);
nand U9462 (N_9462,N_7776,N_7374);
nor U9463 (N_9463,N_7421,N_8160);
nor U9464 (N_9464,N_8050,N_7881);
nor U9465 (N_9465,N_7858,N_7699);
xor U9466 (N_9466,N_8397,N_7758);
nor U9467 (N_9467,N_7698,N_8020);
nand U9468 (N_9468,N_7494,N_7302);
xnor U9469 (N_9469,N_8071,N_7989);
nand U9470 (N_9470,N_7299,N_7289);
or U9471 (N_9471,N_7762,N_7750);
nand U9472 (N_9472,N_7886,N_7474);
nand U9473 (N_9473,N_7743,N_8012);
and U9474 (N_9474,N_8264,N_7289);
or U9475 (N_9475,N_8254,N_7918);
nand U9476 (N_9476,N_7345,N_7669);
xor U9477 (N_9477,N_7434,N_8366);
and U9478 (N_9478,N_8040,N_7541);
xnor U9479 (N_9479,N_7820,N_7384);
nand U9480 (N_9480,N_8334,N_7415);
and U9481 (N_9481,N_8076,N_7629);
nand U9482 (N_9482,N_8235,N_7829);
nand U9483 (N_9483,N_8095,N_7536);
and U9484 (N_9484,N_7714,N_7613);
and U9485 (N_9485,N_7801,N_7504);
nor U9486 (N_9486,N_7466,N_7300);
nand U9487 (N_9487,N_7470,N_8132);
nand U9488 (N_9488,N_7275,N_8362);
nor U9489 (N_9489,N_8084,N_7351);
nor U9490 (N_9490,N_8095,N_7750);
or U9491 (N_9491,N_7552,N_7643);
nand U9492 (N_9492,N_7978,N_7617);
or U9493 (N_9493,N_7389,N_7927);
xnor U9494 (N_9494,N_8334,N_8362);
xor U9495 (N_9495,N_7929,N_7995);
or U9496 (N_9496,N_8364,N_8337);
nand U9497 (N_9497,N_7299,N_8350);
xor U9498 (N_9498,N_7311,N_7723);
or U9499 (N_9499,N_7302,N_7325);
or U9500 (N_9500,N_7755,N_8307);
nand U9501 (N_9501,N_7351,N_8060);
nand U9502 (N_9502,N_7999,N_8130);
nor U9503 (N_9503,N_8248,N_7562);
or U9504 (N_9504,N_7975,N_8199);
or U9505 (N_9505,N_7535,N_8034);
nor U9506 (N_9506,N_8127,N_7625);
and U9507 (N_9507,N_7848,N_8279);
nand U9508 (N_9508,N_7476,N_8101);
or U9509 (N_9509,N_7378,N_7829);
or U9510 (N_9510,N_8117,N_8338);
xnor U9511 (N_9511,N_7326,N_8003);
and U9512 (N_9512,N_7818,N_7431);
nor U9513 (N_9513,N_7363,N_8012);
xor U9514 (N_9514,N_8395,N_7420);
nor U9515 (N_9515,N_7984,N_7939);
xnor U9516 (N_9516,N_7681,N_8193);
and U9517 (N_9517,N_7558,N_7312);
or U9518 (N_9518,N_7557,N_7831);
and U9519 (N_9519,N_8104,N_7652);
nand U9520 (N_9520,N_8022,N_8136);
and U9521 (N_9521,N_7657,N_7270);
xor U9522 (N_9522,N_7562,N_7833);
and U9523 (N_9523,N_7379,N_8393);
nor U9524 (N_9524,N_7773,N_7358);
nand U9525 (N_9525,N_8024,N_7808);
xnor U9526 (N_9526,N_7827,N_8296);
nand U9527 (N_9527,N_7489,N_8066);
nand U9528 (N_9528,N_8204,N_7920);
and U9529 (N_9529,N_7837,N_7320);
xnor U9530 (N_9530,N_7652,N_7803);
xor U9531 (N_9531,N_7956,N_8225);
and U9532 (N_9532,N_7643,N_7694);
and U9533 (N_9533,N_7685,N_8293);
xnor U9534 (N_9534,N_7955,N_7607);
or U9535 (N_9535,N_7566,N_7985);
nor U9536 (N_9536,N_7516,N_7647);
or U9537 (N_9537,N_7430,N_7995);
xnor U9538 (N_9538,N_7363,N_7995);
xnor U9539 (N_9539,N_7246,N_8330);
xnor U9540 (N_9540,N_8283,N_7384);
nor U9541 (N_9541,N_7980,N_7234);
or U9542 (N_9542,N_7627,N_7309);
xnor U9543 (N_9543,N_7279,N_7862);
xor U9544 (N_9544,N_8110,N_8016);
or U9545 (N_9545,N_7782,N_7292);
or U9546 (N_9546,N_8359,N_8196);
and U9547 (N_9547,N_7558,N_8365);
nand U9548 (N_9548,N_8270,N_7643);
or U9549 (N_9549,N_7438,N_7839);
nor U9550 (N_9550,N_8191,N_7522);
nor U9551 (N_9551,N_7551,N_7330);
xor U9552 (N_9552,N_8334,N_7413);
nand U9553 (N_9553,N_7305,N_7348);
and U9554 (N_9554,N_8060,N_8046);
nor U9555 (N_9555,N_7976,N_7483);
and U9556 (N_9556,N_7926,N_7830);
nand U9557 (N_9557,N_7485,N_7380);
nand U9558 (N_9558,N_7685,N_7233);
xnor U9559 (N_9559,N_8304,N_7234);
xor U9560 (N_9560,N_7494,N_7542);
or U9561 (N_9561,N_8302,N_7374);
or U9562 (N_9562,N_7678,N_7430);
nor U9563 (N_9563,N_7742,N_8188);
or U9564 (N_9564,N_8303,N_7727);
and U9565 (N_9565,N_7530,N_7278);
nor U9566 (N_9566,N_8271,N_8113);
nand U9567 (N_9567,N_7918,N_7659);
nor U9568 (N_9568,N_8239,N_8382);
or U9569 (N_9569,N_7380,N_8104);
and U9570 (N_9570,N_7553,N_7619);
and U9571 (N_9571,N_7275,N_7217);
nand U9572 (N_9572,N_7301,N_8032);
nand U9573 (N_9573,N_8338,N_7469);
nor U9574 (N_9574,N_7647,N_8015);
or U9575 (N_9575,N_7627,N_7587);
nand U9576 (N_9576,N_8212,N_7826);
and U9577 (N_9577,N_7684,N_7524);
or U9578 (N_9578,N_7247,N_7501);
and U9579 (N_9579,N_7678,N_7278);
nand U9580 (N_9580,N_7685,N_7380);
and U9581 (N_9581,N_7311,N_7320);
nand U9582 (N_9582,N_8234,N_8253);
nor U9583 (N_9583,N_7337,N_7789);
nor U9584 (N_9584,N_8198,N_7802);
or U9585 (N_9585,N_7231,N_7645);
xor U9586 (N_9586,N_8377,N_8354);
nand U9587 (N_9587,N_7270,N_8075);
nand U9588 (N_9588,N_8230,N_8111);
xnor U9589 (N_9589,N_7466,N_8249);
or U9590 (N_9590,N_7853,N_7559);
or U9591 (N_9591,N_7956,N_7581);
nor U9592 (N_9592,N_7658,N_7622);
or U9593 (N_9593,N_8342,N_8308);
nor U9594 (N_9594,N_7248,N_7410);
and U9595 (N_9595,N_8327,N_8041);
nand U9596 (N_9596,N_7269,N_8138);
nand U9597 (N_9597,N_8073,N_7973);
nand U9598 (N_9598,N_8158,N_7369);
and U9599 (N_9599,N_8150,N_7600);
xor U9600 (N_9600,N_9477,N_8502);
or U9601 (N_9601,N_9047,N_9017);
or U9602 (N_9602,N_8719,N_8601);
or U9603 (N_9603,N_9157,N_8498);
nand U9604 (N_9604,N_9331,N_9392);
nor U9605 (N_9605,N_8709,N_8699);
xnor U9606 (N_9606,N_8729,N_9596);
nand U9607 (N_9607,N_8744,N_9574);
xnor U9608 (N_9608,N_9373,N_9554);
or U9609 (N_9609,N_8424,N_8901);
nor U9610 (N_9610,N_9352,N_8926);
and U9611 (N_9611,N_8478,N_9351);
or U9612 (N_9612,N_9390,N_9181);
xor U9613 (N_9613,N_9290,N_9315);
or U9614 (N_9614,N_9182,N_8983);
nor U9615 (N_9615,N_8669,N_8837);
nor U9616 (N_9616,N_8470,N_8619);
or U9617 (N_9617,N_8847,N_9243);
nor U9618 (N_9618,N_9457,N_9590);
xnor U9619 (N_9619,N_8716,N_9503);
or U9620 (N_9620,N_8516,N_8783);
nand U9621 (N_9621,N_9086,N_8609);
or U9622 (N_9622,N_8540,N_8757);
xor U9623 (N_9623,N_9480,N_9211);
nand U9624 (N_9624,N_9591,N_9174);
or U9625 (N_9625,N_8950,N_9512);
xor U9626 (N_9626,N_9472,N_8706);
or U9627 (N_9627,N_9179,N_8923);
xor U9628 (N_9628,N_9024,N_9319);
or U9629 (N_9629,N_9432,N_9012);
nor U9630 (N_9630,N_9430,N_8506);
nor U9631 (N_9631,N_8772,N_8414);
or U9632 (N_9632,N_8727,N_9049);
xor U9633 (N_9633,N_9587,N_8491);
and U9634 (N_9634,N_9402,N_9113);
and U9635 (N_9635,N_8530,N_8425);
xor U9636 (N_9636,N_8446,N_9494);
and U9637 (N_9637,N_8452,N_8936);
or U9638 (N_9638,N_9345,N_9001);
nor U9639 (N_9639,N_9454,N_9306);
nor U9640 (N_9640,N_8830,N_9483);
nand U9641 (N_9641,N_8542,N_8415);
or U9642 (N_9642,N_9560,N_9010);
nand U9643 (N_9643,N_8918,N_9418);
and U9644 (N_9644,N_9118,N_8982);
or U9645 (N_9645,N_8739,N_9581);
and U9646 (N_9646,N_8802,N_9028);
nand U9647 (N_9647,N_9405,N_9014);
nor U9648 (N_9648,N_9215,N_9470);
and U9649 (N_9649,N_9038,N_8900);
and U9650 (N_9650,N_8872,N_9170);
nor U9651 (N_9651,N_8660,N_9117);
nand U9652 (N_9652,N_9052,N_9207);
or U9653 (N_9653,N_9521,N_9252);
or U9654 (N_9654,N_9260,N_9226);
xor U9655 (N_9655,N_9556,N_9023);
or U9656 (N_9656,N_8490,N_9530);
and U9657 (N_9657,N_8819,N_8766);
and U9658 (N_9658,N_9068,N_9225);
and U9659 (N_9659,N_8643,N_9486);
nor U9660 (N_9660,N_8677,N_8980);
nand U9661 (N_9661,N_9496,N_9362);
and U9662 (N_9662,N_9350,N_8707);
or U9663 (N_9663,N_9079,N_9022);
nand U9664 (N_9664,N_8433,N_8764);
and U9665 (N_9665,N_8467,N_9167);
and U9666 (N_9666,N_8856,N_8788);
or U9667 (N_9667,N_9297,N_9070);
nand U9668 (N_9668,N_8972,N_8913);
and U9669 (N_9669,N_9407,N_8815);
nor U9670 (N_9670,N_8921,N_9111);
nand U9671 (N_9671,N_9580,N_9206);
xnor U9672 (N_9672,N_9365,N_8678);
nand U9673 (N_9673,N_8708,N_9193);
or U9674 (N_9674,N_9506,N_8653);
or U9675 (N_9675,N_8496,N_8906);
xnor U9676 (N_9676,N_9160,N_8547);
nor U9677 (N_9677,N_9371,N_9221);
nand U9678 (N_9678,N_8529,N_8474);
and U9679 (N_9679,N_8756,N_8705);
xor U9680 (N_9680,N_9162,N_8537);
xnor U9681 (N_9681,N_8561,N_8544);
nand U9682 (N_9682,N_8578,N_8689);
or U9683 (N_9683,N_9540,N_9437);
xor U9684 (N_9684,N_8483,N_8700);
nor U9685 (N_9685,N_9481,N_8748);
xnor U9686 (N_9686,N_9239,N_9305);
or U9687 (N_9687,N_9148,N_9577);
nand U9688 (N_9688,N_8551,N_9576);
xor U9689 (N_9689,N_9594,N_9338);
and U9690 (N_9690,N_9375,N_9125);
nor U9691 (N_9691,N_9080,N_8785);
xor U9692 (N_9692,N_8817,N_8541);
or U9693 (N_9693,N_8994,N_9381);
xnor U9694 (N_9694,N_8697,N_9075);
nand U9695 (N_9695,N_8987,N_8468);
nand U9696 (N_9696,N_9468,N_8975);
nand U9697 (N_9697,N_9466,N_9191);
or U9698 (N_9698,N_9364,N_8687);
xnor U9699 (N_9699,N_9000,N_9188);
or U9700 (N_9700,N_9573,N_8948);
and U9701 (N_9701,N_8686,N_9458);
xnor U9702 (N_9702,N_9161,N_8639);
or U9703 (N_9703,N_9097,N_9508);
and U9704 (N_9704,N_9220,N_9547);
or U9705 (N_9705,N_8615,N_8621);
xor U9706 (N_9706,N_9471,N_9548);
nor U9707 (N_9707,N_9124,N_8622);
or U9708 (N_9708,N_9115,N_8656);
nand U9709 (N_9709,N_8512,N_8665);
nor U9710 (N_9710,N_8489,N_8888);
xnor U9711 (N_9711,N_8846,N_9387);
nor U9712 (N_9712,N_8447,N_9398);
nand U9713 (N_9713,N_9469,N_8455);
xnor U9714 (N_9714,N_9278,N_8886);
nand U9715 (N_9715,N_8967,N_9077);
and U9716 (N_9716,N_9196,N_9213);
and U9717 (N_9717,N_8796,N_8976);
and U9718 (N_9718,N_9438,N_8422);
nand U9719 (N_9719,N_8614,N_8481);
nand U9720 (N_9720,N_8563,N_9133);
or U9721 (N_9721,N_9083,N_8778);
nand U9722 (N_9722,N_8903,N_9569);
and U9723 (N_9723,N_8620,N_9138);
nor U9724 (N_9724,N_8857,N_9489);
nand U9725 (N_9725,N_9178,N_9484);
or U9726 (N_9726,N_8443,N_9465);
xnor U9727 (N_9727,N_9516,N_9265);
nor U9728 (N_9728,N_9116,N_8878);
nand U9729 (N_9729,N_9456,N_9055);
or U9730 (N_9730,N_9443,N_9441);
or U9731 (N_9731,N_8775,N_9327);
or U9732 (N_9732,N_8768,N_8560);
and U9733 (N_9733,N_8771,N_8457);
nand U9734 (N_9734,N_9183,N_9132);
nand U9735 (N_9735,N_8947,N_9250);
xor U9736 (N_9736,N_9410,N_8645);
or U9737 (N_9737,N_9229,N_9254);
and U9738 (N_9738,N_9292,N_8995);
nor U9739 (N_9739,N_9499,N_8713);
xnor U9740 (N_9740,N_8835,N_8532);
nor U9741 (N_9741,N_8717,N_9413);
nor U9742 (N_9742,N_9522,N_9435);
nor U9743 (N_9743,N_9434,N_8673);
or U9744 (N_9744,N_9289,N_8877);
and U9745 (N_9745,N_9180,N_8962);
nand U9746 (N_9746,N_8984,N_8895);
and U9747 (N_9747,N_8465,N_9598);
nor U9748 (N_9748,N_8576,N_9277);
and U9749 (N_9749,N_9201,N_9171);
or U9750 (N_9750,N_8851,N_8864);
xor U9751 (N_9751,N_9427,N_9450);
nor U9752 (N_9752,N_9241,N_9420);
nor U9753 (N_9753,N_8957,N_8734);
nor U9754 (N_9754,N_8822,N_8504);
or U9755 (N_9755,N_9359,N_9421);
nand U9756 (N_9756,N_9110,N_8434);
nor U9757 (N_9757,N_9426,N_8832);
nor U9758 (N_9758,N_8992,N_9126);
nand U9759 (N_9759,N_8943,N_8435);
nor U9760 (N_9760,N_8676,N_9262);
nor U9761 (N_9761,N_8482,N_8998);
nand U9762 (N_9762,N_9357,N_9411);
nor U9763 (N_9763,N_8798,N_8632);
or U9764 (N_9764,N_8945,N_8604);
nor U9765 (N_9765,N_8445,N_8550);
or U9766 (N_9766,N_8965,N_8492);
nand U9767 (N_9767,N_8476,N_8630);
or U9768 (N_9768,N_9342,N_8685);
nor U9769 (N_9769,N_8911,N_9005);
nor U9770 (N_9770,N_8733,N_8955);
nor U9771 (N_9771,N_9224,N_8963);
nand U9772 (N_9772,N_9151,N_8602);
or U9773 (N_9773,N_9247,N_9310);
nor U9774 (N_9774,N_8456,N_8993);
nand U9775 (N_9775,N_9417,N_8843);
nand U9776 (N_9776,N_9562,N_9280);
xnor U9777 (N_9777,N_8937,N_9212);
nor U9778 (N_9778,N_9321,N_9041);
nand U9779 (N_9779,N_8809,N_8419);
nand U9780 (N_9780,N_8556,N_8932);
nand U9781 (N_9781,N_8858,N_9461);
nor U9782 (N_9782,N_9004,N_8960);
and U9783 (N_9783,N_9425,N_8666);
nand U9784 (N_9784,N_8789,N_9016);
nand U9785 (N_9785,N_8631,N_8519);
xor U9786 (N_9786,N_9475,N_8839);
or U9787 (N_9787,N_8825,N_8511);
or U9788 (N_9788,N_9048,N_8428);
nand U9789 (N_9789,N_8774,N_8919);
and U9790 (N_9790,N_8517,N_9449);
nand U9791 (N_9791,N_9159,N_8812);
and U9792 (N_9792,N_8701,N_9520);
nand U9793 (N_9793,N_8411,N_9296);
xor U9794 (N_9794,N_9042,N_9524);
and U9795 (N_9795,N_9197,N_9533);
nand U9796 (N_9796,N_8915,N_8905);
xnor U9797 (N_9797,N_8930,N_9380);
nand U9798 (N_9798,N_8741,N_8611);
and U9799 (N_9799,N_9071,N_9195);
xor U9800 (N_9800,N_9451,N_9036);
xor U9801 (N_9801,N_8480,N_9199);
nand U9802 (N_9802,N_8855,N_8964);
or U9803 (N_9803,N_9204,N_8641);
nand U9804 (N_9804,N_8494,N_8968);
nor U9805 (N_9805,N_9487,N_9491);
or U9806 (N_9806,N_8410,N_8587);
nand U9807 (N_9807,N_8724,N_9234);
nor U9808 (N_9808,N_8479,N_8786);
and U9809 (N_9809,N_9332,N_9130);
xnor U9810 (N_9810,N_9172,N_9184);
nor U9811 (N_9811,N_8626,N_8881);
xnor U9812 (N_9812,N_8600,N_8471);
nand U9813 (N_9813,N_8583,N_9102);
and U9814 (N_9814,N_9388,N_8728);
nand U9815 (N_9815,N_9511,N_8533);
xor U9816 (N_9816,N_8703,N_8637);
nand U9817 (N_9817,N_9498,N_8953);
nand U9818 (N_9818,N_9176,N_8460);
and U9819 (N_9819,N_8554,N_9139);
nand U9820 (N_9820,N_8674,N_9377);
xor U9821 (N_9821,N_8890,N_9222);
or U9822 (N_9822,N_9538,N_9216);
xor U9823 (N_9823,N_9145,N_9066);
and U9824 (N_9824,N_9433,N_9085);
nand U9825 (N_9825,N_9136,N_9103);
and U9826 (N_9826,N_9009,N_9309);
and U9827 (N_9827,N_9549,N_8859);
nand U9828 (N_9828,N_9579,N_8842);
and U9829 (N_9829,N_9492,N_8401);
nor U9830 (N_9830,N_8528,N_8657);
and U9831 (N_9831,N_8836,N_8612);
nand U9832 (N_9832,N_8940,N_8579);
and U9833 (N_9833,N_9393,N_9593);
and U9834 (N_9834,N_8966,N_9561);
or U9835 (N_9835,N_8990,N_8679);
nand U9836 (N_9836,N_9505,N_8951);
nor U9837 (N_9837,N_9372,N_9541);
or U9838 (N_9838,N_8499,N_9249);
nand U9839 (N_9839,N_8613,N_9099);
xor U9840 (N_9840,N_8523,N_9109);
or U9841 (N_9841,N_9589,N_8811);
xor U9842 (N_9842,N_8509,N_8608);
and U9843 (N_9843,N_9572,N_9553);
xnor U9844 (N_9844,N_8912,N_8751);
xnor U9845 (N_9845,N_8698,N_9253);
and U9846 (N_9846,N_9007,N_9464);
nor U9847 (N_9847,N_9476,N_9436);
nand U9848 (N_9848,N_9311,N_9033);
nand U9849 (N_9849,N_9527,N_8749);
nor U9850 (N_9850,N_9389,N_8553);
nand U9851 (N_9851,N_9269,N_9382);
or U9852 (N_9852,N_8816,N_8754);
nand U9853 (N_9853,N_9385,N_8454);
xor U9854 (N_9854,N_9045,N_8437);
nand U9855 (N_9855,N_9173,N_8803);
and U9856 (N_9856,N_8814,N_8603);
or U9857 (N_9857,N_9208,N_9051);
nor U9858 (N_9858,N_9584,N_9266);
xnor U9859 (N_9859,N_8670,N_9163);
xnor U9860 (N_9860,N_9270,N_8423);
nor U9861 (N_9861,N_9044,N_8833);
nand U9862 (N_9862,N_8444,N_8904);
xor U9863 (N_9863,N_8784,N_9513);
and U9864 (N_9864,N_9166,N_8552);
nand U9865 (N_9865,N_9013,N_8776);
nand U9866 (N_9866,N_9585,N_9150);
nor U9867 (N_9867,N_9061,N_9008);
or U9868 (N_9868,N_8868,N_9233);
xor U9869 (N_9869,N_8758,N_9299);
xor U9870 (N_9870,N_9106,N_8664);
or U9871 (N_9871,N_8651,N_8638);
or U9872 (N_9872,N_9261,N_9539);
nand U9873 (N_9873,N_8834,N_9356);
nor U9874 (N_9874,N_9142,N_8412);
nor U9875 (N_9875,N_8647,N_9123);
xor U9876 (N_9876,N_8969,N_9129);
nor U9877 (N_9877,N_8400,N_8873);
nor U9878 (N_9878,N_8896,N_9232);
nand U9879 (N_9879,N_8773,N_8623);
xor U9880 (N_9880,N_9019,N_8720);
nand U9881 (N_9881,N_8941,N_8485);
nand U9882 (N_9882,N_8743,N_9240);
xor U9883 (N_9883,N_9406,N_8746);
and U9884 (N_9884,N_9228,N_9490);
or U9885 (N_9885,N_9531,N_8655);
or U9886 (N_9886,N_9089,N_9281);
and U9887 (N_9887,N_8879,N_9276);
or U9888 (N_9888,N_9543,N_9107);
nand U9889 (N_9889,N_8979,N_9399);
or U9890 (N_9890,N_8642,N_9015);
or U9891 (N_9891,N_9187,N_9040);
nand U9892 (N_9892,N_9237,N_8497);
and U9893 (N_9893,N_9330,N_8871);
nor U9894 (N_9894,N_9235,N_8763);
and U9895 (N_9895,N_9114,N_8954);
xnor U9896 (N_9896,N_8870,N_9488);
and U9897 (N_9897,N_8634,N_8790);
xnor U9898 (N_9898,N_9128,N_9302);
or U9899 (N_9899,N_9343,N_9446);
or U9900 (N_9900,N_8605,N_8958);
and U9901 (N_9901,N_8688,N_9067);
xor U9902 (N_9902,N_8824,N_9282);
or U9903 (N_9903,N_9037,N_9460);
and U9904 (N_9904,N_9018,N_8750);
nand U9905 (N_9905,N_9186,N_9072);
xor U9906 (N_9906,N_9416,N_9273);
and U9907 (N_9907,N_8761,N_9101);
and U9908 (N_9908,N_9242,N_8577);
or U9909 (N_9909,N_9528,N_9246);
nand U9910 (N_9910,N_9096,N_9011);
nand U9911 (N_9911,N_8569,N_8978);
nor U9912 (N_9912,N_9412,N_9519);
and U9913 (N_9913,N_8505,N_9339);
or U9914 (N_9914,N_9069,N_9003);
and U9915 (N_9915,N_8416,N_8874);
and U9916 (N_9916,N_8715,N_9029);
nor U9917 (N_9917,N_8770,N_9092);
nor U9918 (N_9918,N_8795,N_8907);
and U9919 (N_9919,N_8791,N_9526);
or U9920 (N_9920,N_8559,N_9076);
nor U9921 (N_9921,N_8767,N_9177);
nand U9922 (N_9922,N_8885,N_9104);
xor U9923 (N_9923,N_9473,N_8531);
or U9924 (N_9924,N_8828,N_9131);
nand U9925 (N_9925,N_8555,N_8797);
xnor U9926 (N_9926,N_9156,N_9043);
nor U9927 (N_9927,N_9419,N_8925);
and U9928 (N_9928,N_8418,N_8929);
nand U9929 (N_9929,N_9564,N_9027);
nand U9930 (N_9930,N_8617,N_8762);
and U9931 (N_9931,N_8760,N_9578);
nand U9932 (N_9932,N_9358,N_9317);
nand U9933 (N_9933,N_8672,N_9555);
or U9934 (N_9934,N_8780,N_8794);
xnor U9935 (N_9935,N_8813,N_9062);
nand U9936 (N_9936,N_9403,N_9320);
nor U9937 (N_9937,N_8404,N_9158);
xnor U9938 (N_9938,N_9053,N_9284);
or U9939 (N_9939,N_9544,N_8782);
and U9940 (N_9940,N_9346,N_8882);
xor U9941 (N_9941,N_9303,N_8826);
and U9942 (N_9942,N_8752,N_8440);
nand U9943 (N_9943,N_9349,N_9251);
nor U9944 (N_9944,N_8821,N_9341);
or U9945 (N_9945,N_8829,N_8894);
xnor U9946 (N_9946,N_8690,N_8723);
nand U9947 (N_9947,N_9428,N_9384);
nor U9948 (N_9948,N_9408,N_8799);
or U9949 (N_9949,N_8736,N_8801);
xor U9950 (N_9950,N_9312,N_9328);
or U9951 (N_9951,N_8648,N_8472);
xor U9952 (N_9952,N_8714,N_9236);
nand U9953 (N_9953,N_8683,N_9353);
nand U9954 (N_9954,N_8938,N_8596);
xor U9955 (N_9955,N_8702,N_9091);
nand U9956 (N_9956,N_9583,N_9227);
nand U9957 (N_9957,N_9453,N_8513);
or U9958 (N_9958,N_8680,N_9588);
or U9959 (N_9959,N_8586,N_8942);
nor U9960 (N_9960,N_8624,N_9294);
and U9961 (N_9961,N_8807,N_9064);
and U9962 (N_9962,N_9209,N_8726);
or U9963 (N_9963,N_8538,N_8571);
and U9964 (N_9964,N_8845,N_9223);
xor U9965 (N_9965,N_9571,N_9198);
xnor U9966 (N_9966,N_9546,N_9065);
or U9967 (N_9967,N_9073,N_9448);
xnor U9968 (N_9968,N_9344,N_9194);
nor U9969 (N_9969,N_8590,N_8853);
nor U9970 (N_9970,N_9256,N_8747);
nand U9971 (N_9971,N_9295,N_8500);
nor U9972 (N_9972,N_8407,N_8974);
xor U9973 (N_9973,N_8607,N_9482);
nor U9974 (N_9974,N_8566,N_8889);
or U9975 (N_9975,N_9597,N_8759);
or U9976 (N_9976,N_8922,N_8408);
xor U9977 (N_9977,N_9169,N_9268);
nor U9978 (N_9978,N_9322,N_9401);
xor U9979 (N_9979,N_9378,N_8486);
or U9980 (N_9980,N_8536,N_8503);
and U9981 (N_9981,N_8573,N_8406);
nand U9982 (N_9982,N_9523,N_8989);
xnor U9983 (N_9983,N_8469,N_8927);
nor U9984 (N_9984,N_9248,N_8875);
and U9985 (N_9985,N_8652,N_9210);
nand U9986 (N_9986,N_9030,N_8891);
xnor U9987 (N_9987,N_8755,N_9267);
nand U9988 (N_9988,N_9165,N_9127);
or U9989 (N_9989,N_8463,N_9143);
and U9990 (N_9990,N_8898,N_8722);
nor U9991 (N_9991,N_9415,N_8704);
and U9992 (N_9992,N_8935,N_8931);
and U9993 (N_9993,N_9542,N_8887);
nor U9994 (N_9994,N_8737,N_9386);
nand U9995 (N_9995,N_8961,N_8884);
nand U9996 (N_9996,N_9545,N_8769);
nor U9997 (N_9997,N_8451,N_8597);
or U9998 (N_9998,N_9324,N_9271);
xor U9999 (N_9999,N_9367,N_8777);
and U10000 (N_10000,N_9535,N_8682);
and U10001 (N_10001,N_9383,N_9440);
or U10002 (N_10002,N_9200,N_8949);
xnor U10003 (N_10003,N_9087,N_9463);
nor U10004 (N_10004,N_8663,N_9366);
and U10005 (N_10005,N_8668,N_9502);
nand U10006 (N_10006,N_9063,N_9259);
xor U10007 (N_10007,N_8908,N_8477);
and U10008 (N_10008,N_9485,N_8650);
nor U10009 (N_10009,N_9034,N_9431);
or U10010 (N_10010,N_9122,N_9155);
nand U10011 (N_10011,N_8838,N_8458);
or U10012 (N_10012,N_9455,N_8997);
and U10013 (N_10013,N_8787,N_8920);
nand U10014 (N_10014,N_8712,N_9154);
nand U10015 (N_10015,N_8501,N_9557);
nand U10016 (N_10016,N_8403,N_9374);
xnor U10017 (N_10017,N_9105,N_9190);
xor U10018 (N_10018,N_9340,N_9120);
xor U10019 (N_10019,N_8409,N_8426);
and U10020 (N_10020,N_8522,N_8996);
nand U10021 (N_10021,N_9031,N_8661);
xnor U10022 (N_10022,N_8986,N_9060);
xnor U10023 (N_10023,N_9057,N_9323);
xnor U10024 (N_10024,N_9192,N_8618);
nand U10025 (N_10025,N_8515,N_9094);
nand U10026 (N_10026,N_9032,N_9500);
nand U10027 (N_10027,N_8779,N_8565);
nor U10028 (N_10028,N_9474,N_9424);
or U10029 (N_10029,N_9285,N_9025);
or U10030 (N_10030,N_9283,N_9098);
or U10031 (N_10031,N_9462,N_9536);
nand U10032 (N_10032,N_8939,N_8850);
or U10033 (N_10033,N_9230,N_9509);
nor U10034 (N_10034,N_8731,N_8909);
nand U10035 (N_10035,N_8484,N_9559);
or U10036 (N_10036,N_9495,N_8545);
and U10037 (N_10037,N_9257,N_9334);
nand U10038 (N_10038,N_9361,N_8981);
or U10039 (N_10039,N_8453,N_8848);
or U10040 (N_10040,N_8421,N_8633);
or U10041 (N_10041,N_9404,N_8459);
or U10042 (N_10042,N_9026,N_8820);
or U10043 (N_10043,N_8487,N_8721);
xnor U10044 (N_10044,N_9429,N_9175);
xor U10045 (N_10045,N_8438,N_8442);
xnor U10046 (N_10046,N_9575,N_8575);
or U10047 (N_10047,N_8781,N_9035);
nand U10048 (N_10048,N_8629,N_8402);
nand U10049 (N_10049,N_8933,N_8543);
nor U10050 (N_10050,N_8589,N_9144);
nor U10051 (N_10051,N_8946,N_8861);
xnor U10052 (N_10052,N_9141,N_8549);
or U10053 (N_10053,N_8892,N_8675);
nand U10054 (N_10054,N_9376,N_9279);
and U10055 (N_10055,N_9558,N_8521);
nand U10056 (N_10056,N_9510,N_8827);
nor U10057 (N_10057,N_8991,N_9082);
nand U10058 (N_10058,N_9287,N_8585);
nand U10059 (N_10059,N_9255,N_8448);
nand U10060 (N_10060,N_8581,N_8902);
xor U10061 (N_10061,N_8588,N_9565);
or U10062 (N_10062,N_9301,N_8854);
or U10063 (N_10063,N_9336,N_8636);
and U10064 (N_10064,N_8718,N_9363);
nor U10065 (N_10065,N_8567,N_9263);
and U10066 (N_10066,N_8985,N_9217);
nor U10067 (N_10067,N_9370,N_9369);
or U10068 (N_10068,N_8740,N_8971);
or U10069 (N_10069,N_8808,N_8649);
or U10070 (N_10070,N_9409,N_9056);
or U10071 (N_10071,N_9050,N_9313);
nor U10072 (N_10072,N_9397,N_8507);
nand U10073 (N_10073,N_8792,N_8449);
xnor U10074 (N_10074,N_8765,N_8534);
or U10075 (N_10075,N_9368,N_9314);
nand U10076 (N_10076,N_8535,N_8635);
and U10077 (N_10077,N_8849,N_9395);
nand U10078 (N_10078,N_9391,N_8671);
xor U10079 (N_10079,N_8973,N_8644);
and U10080 (N_10080,N_8897,N_8732);
xnor U10081 (N_10081,N_8510,N_9264);
nor U10082 (N_10082,N_8970,N_8562);
nand U10083 (N_10083,N_8738,N_9203);
xnor U10084 (N_10084,N_9134,N_9423);
xor U10085 (N_10085,N_8831,N_8610);
or U10086 (N_10086,N_8711,N_8606);
xor U10087 (N_10087,N_8742,N_8710);
nand U10088 (N_10088,N_8546,N_8594);
nand U10089 (N_10089,N_9478,N_9189);
and U10090 (N_10090,N_9396,N_9467);
xor U10091 (N_10091,N_8667,N_9238);
xor U10092 (N_10092,N_8681,N_9231);
xor U10093 (N_10093,N_9566,N_8493);
or U10094 (N_10094,N_8430,N_8863);
or U10095 (N_10095,N_9006,N_8753);
nor U10096 (N_10096,N_9518,N_9245);
nand U10097 (N_10097,N_8952,N_8417);
or U10098 (N_10098,N_9515,N_8805);
or U10099 (N_10099,N_8439,N_9379);
and U10100 (N_10100,N_8413,N_9595);
or U10101 (N_10101,N_8508,N_8917);
and U10102 (N_10102,N_9152,N_9459);
or U10103 (N_10103,N_9586,N_9149);
and U10104 (N_10104,N_9112,N_8495);
nand U10105 (N_10105,N_8988,N_8595);
nand U10106 (N_10106,N_8466,N_9298);
nand U10107 (N_10107,N_8431,N_9507);
xnor U10108 (N_10108,N_9074,N_9293);
nor U10109 (N_10109,N_8514,N_8916);
nand U10110 (N_10110,N_8924,N_8880);
xnor U10111 (N_10111,N_8899,N_8841);
or U10112 (N_10112,N_9307,N_9185);
xnor U10113 (N_10113,N_9078,N_9354);
nand U10114 (N_10114,N_8564,N_9355);
nor U10115 (N_10115,N_8745,N_9291);
and U10116 (N_10116,N_8910,N_9550);
and U10117 (N_10117,N_9529,N_8628);
nor U10118 (N_10118,N_8658,N_8818);
nand U10119 (N_10119,N_8548,N_9318);
xor U10120 (N_10120,N_8473,N_9517);
xnor U10121 (N_10121,N_9568,N_8580);
and U10122 (N_10122,N_9202,N_9275);
and U10123 (N_10123,N_8944,N_9348);
or U10124 (N_10124,N_9537,N_8570);
and U10125 (N_10125,N_8572,N_9563);
nand U10126 (N_10126,N_8462,N_8696);
or U10127 (N_10127,N_9258,N_9447);
or U10128 (N_10128,N_8860,N_9444);
nor U10129 (N_10129,N_8525,N_8592);
nand U10130 (N_10130,N_8810,N_8793);
and U10131 (N_10131,N_9108,N_9081);
xor U10132 (N_10132,N_9272,N_9214);
xnor U10133 (N_10133,N_9135,N_8804);
and U10134 (N_10134,N_8852,N_8869);
nor U10135 (N_10135,N_8488,N_8693);
or U10136 (N_10136,N_8557,N_8640);
and U10137 (N_10137,N_9329,N_8934);
nor U10138 (N_10138,N_9552,N_8526);
and U10139 (N_10139,N_9534,N_9439);
nand U10140 (N_10140,N_8800,N_9414);
nor U10141 (N_10141,N_8999,N_8518);
and U10142 (N_10142,N_8977,N_8691);
xnor U10143 (N_10143,N_8865,N_9445);
and U10144 (N_10144,N_9337,N_8616);
nand U10145 (N_10145,N_8876,N_9599);
xor U10146 (N_10146,N_9218,N_9501);
and U10147 (N_10147,N_9205,N_8558);
or U10148 (N_10148,N_9140,N_8432);
nand U10149 (N_10149,N_9100,N_9121);
xnor U10150 (N_10150,N_9452,N_9326);
xnor U10151 (N_10151,N_8866,N_8627);
and U10152 (N_10152,N_8598,N_9308);
nor U10153 (N_10153,N_9567,N_9347);
and U10154 (N_10154,N_8735,N_8461);
or U10155 (N_10155,N_8646,N_8694);
or U10156 (N_10156,N_9316,N_9093);
xnor U10157 (N_10157,N_9335,N_9504);
and U10158 (N_10158,N_9532,N_8527);
xor U10159 (N_10159,N_8914,N_8956);
or U10160 (N_10160,N_8654,N_8684);
and U10161 (N_10161,N_9137,N_9059);
or U10162 (N_10162,N_8840,N_8582);
or U10163 (N_10163,N_8883,N_8464);
or U10164 (N_10164,N_9095,N_9153);
xnor U10165 (N_10165,N_8893,N_8405);
or U10166 (N_10166,N_8475,N_9582);
or U10167 (N_10167,N_8420,N_9360);
nor U10168 (N_10168,N_9525,N_8441);
xor U10169 (N_10169,N_8450,N_9058);
nor U10170 (N_10170,N_8844,N_9333);
xnor U10171 (N_10171,N_9497,N_8591);
and U10172 (N_10172,N_9479,N_8568);
xor U10173 (N_10173,N_8574,N_8695);
nor U10174 (N_10174,N_9147,N_9442);
xnor U10175 (N_10175,N_8862,N_9020);
xor U10176 (N_10176,N_9084,N_9090);
nand U10177 (N_10177,N_8625,N_9002);
nor U10178 (N_10178,N_9288,N_8806);
nand U10179 (N_10179,N_9286,N_8520);
and U10180 (N_10180,N_8539,N_9274);
nor U10181 (N_10181,N_9422,N_9021);
nor U10182 (N_10182,N_9570,N_8823);
nor U10183 (N_10183,N_9304,N_9164);
xnor U10184 (N_10184,N_8725,N_9088);
nor U10185 (N_10185,N_8593,N_8524);
and U10186 (N_10186,N_9394,N_8730);
xor U10187 (N_10187,N_8429,N_9244);
nand U10188 (N_10188,N_9325,N_9551);
nand U10189 (N_10189,N_9146,N_9168);
nor U10190 (N_10190,N_8436,N_9039);
nand U10191 (N_10191,N_8659,N_8584);
and U10192 (N_10192,N_8928,N_9119);
and U10193 (N_10193,N_9400,N_8599);
xnor U10194 (N_10194,N_9219,N_9300);
nand U10195 (N_10195,N_8692,N_8959);
and U10196 (N_10196,N_8867,N_9046);
nand U10197 (N_10197,N_8662,N_9592);
or U10198 (N_10198,N_9054,N_8427);
xor U10199 (N_10199,N_9514,N_9493);
nand U10200 (N_10200,N_9517,N_8482);
and U10201 (N_10201,N_8442,N_8678);
nand U10202 (N_10202,N_8523,N_9005);
nor U10203 (N_10203,N_8702,N_8662);
xor U10204 (N_10204,N_8441,N_9052);
nand U10205 (N_10205,N_9102,N_8953);
nor U10206 (N_10206,N_8838,N_8682);
nand U10207 (N_10207,N_8405,N_8611);
xor U10208 (N_10208,N_9363,N_8586);
xnor U10209 (N_10209,N_8795,N_8589);
xnor U10210 (N_10210,N_8786,N_9261);
nor U10211 (N_10211,N_9431,N_9328);
xor U10212 (N_10212,N_9373,N_8904);
xor U10213 (N_10213,N_8556,N_8477);
nand U10214 (N_10214,N_9529,N_8880);
nor U10215 (N_10215,N_9121,N_8961);
nor U10216 (N_10216,N_9537,N_8473);
or U10217 (N_10217,N_8565,N_8881);
or U10218 (N_10218,N_8428,N_8975);
nand U10219 (N_10219,N_9342,N_9416);
nor U10220 (N_10220,N_9207,N_8529);
or U10221 (N_10221,N_9099,N_9173);
nand U10222 (N_10222,N_9496,N_8507);
and U10223 (N_10223,N_9390,N_8895);
xnor U10224 (N_10224,N_9533,N_9296);
xnor U10225 (N_10225,N_9470,N_9482);
or U10226 (N_10226,N_8809,N_9242);
xnor U10227 (N_10227,N_8432,N_9107);
xnor U10228 (N_10228,N_9311,N_8582);
xnor U10229 (N_10229,N_8842,N_8755);
or U10230 (N_10230,N_9021,N_9573);
nor U10231 (N_10231,N_9186,N_9329);
xnor U10232 (N_10232,N_9341,N_8892);
or U10233 (N_10233,N_9245,N_9412);
nor U10234 (N_10234,N_8990,N_8735);
xor U10235 (N_10235,N_8516,N_8533);
or U10236 (N_10236,N_8916,N_8550);
or U10237 (N_10237,N_8435,N_9166);
xor U10238 (N_10238,N_8587,N_9199);
or U10239 (N_10239,N_8436,N_8649);
nand U10240 (N_10240,N_8690,N_8468);
xnor U10241 (N_10241,N_8454,N_8580);
and U10242 (N_10242,N_9501,N_8720);
nor U10243 (N_10243,N_9383,N_8554);
nand U10244 (N_10244,N_9032,N_9051);
xor U10245 (N_10245,N_9205,N_9302);
or U10246 (N_10246,N_9481,N_9127);
nor U10247 (N_10247,N_8769,N_8928);
nand U10248 (N_10248,N_8632,N_8832);
nor U10249 (N_10249,N_8686,N_9133);
nor U10250 (N_10250,N_9107,N_9013);
or U10251 (N_10251,N_9533,N_9026);
and U10252 (N_10252,N_9041,N_8410);
and U10253 (N_10253,N_9486,N_9207);
xnor U10254 (N_10254,N_9078,N_8414);
nor U10255 (N_10255,N_8904,N_9052);
and U10256 (N_10256,N_8838,N_9356);
or U10257 (N_10257,N_9089,N_9270);
nor U10258 (N_10258,N_8472,N_9118);
nand U10259 (N_10259,N_9118,N_8441);
or U10260 (N_10260,N_8886,N_8780);
nand U10261 (N_10261,N_8757,N_8502);
nor U10262 (N_10262,N_9290,N_8662);
nand U10263 (N_10263,N_8943,N_9193);
and U10264 (N_10264,N_9425,N_9269);
and U10265 (N_10265,N_9120,N_9586);
nand U10266 (N_10266,N_8543,N_9315);
and U10267 (N_10267,N_8527,N_8781);
nor U10268 (N_10268,N_9586,N_8410);
xnor U10269 (N_10269,N_9350,N_9567);
and U10270 (N_10270,N_9384,N_8799);
xnor U10271 (N_10271,N_9452,N_9166);
or U10272 (N_10272,N_9302,N_8946);
nor U10273 (N_10273,N_9222,N_9421);
or U10274 (N_10274,N_8534,N_8989);
nor U10275 (N_10275,N_9252,N_9387);
or U10276 (N_10276,N_8583,N_9438);
or U10277 (N_10277,N_9316,N_9514);
xor U10278 (N_10278,N_8822,N_9249);
nor U10279 (N_10279,N_9512,N_8407);
or U10280 (N_10280,N_8679,N_9544);
nor U10281 (N_10281,N_8805,N_8969);
nand U10282 (N_10282,N_8834,N_9049);
nand U10283 (N_10283,N_9345,N_9140);
xnor U10284 (N_10284,N_8662,N_9175);
and U10285 (N_10285,N_8744,N_9377);
or U10286 (N_10286,N_8783,N_8835);
or U10287 (N_10287,N_9321,N_8602);
and U10288 (N_10288,N_8521,N_8550);
nand U10289 (N_10289,N_8993,N_8690);
and U10290 (N_10290,N_9131,N_9397);
nor U10291 (N_10291,N_8766,N_8455);
and U10292 (N_10292,N_9545,N_8605);
or U10293 (N_10293,N_8508,N_9227);
or U10294 (N_10294,N_9403,N_8425);
or U10295 (N_10295,N_8665,N_8605);
xnor U10296 (N_10296,N_9556,N_9036);
and U10297 (N_10297,N_8986,N_9386);
nor U10298 (N_10298,N_8707,N_9017);
nor U10299 (N_10299,N_8609,N_9323);
and U10300 (N_10300,N_8905,N_8474);
or U10301 (N_10301,N_8503,N_8993);
and U10302 (N_10302,N_8800,N_8511);
or U10303 (N_10303,N_8852,N_8826);
or U10304 (N_10304,N_8711,N_8928);
nand U10305 (N_10305,N_9018,N_9569);
and U10306 (N_10306,N_9525,N_9142);
and U10307 (N_10307,N_8679,N_8587);
nand U10308 (N_10308,N_8935,N_8649);
nor U10309 (N_10309,N_8690,N_8703);
nand U10310 (N_10310,N_9039,N_8877);
xnor U10311 (N_10311,N_9446,N_8681);
or U10312 (N_10312,N_8600,N_9128);
xor U10313 (N_10313,N_8451,N_9441);
xor U10314 (N_10314,N_8680,N_9472);
xnor U10315 (N_10315,N_9324,N_8610);
and U10316 (N_10316,N_9358,N_8887);
and U10317 (N_10317,N_9298,N_9327);
or U10318 (N_10318,N_9324,N_9386);
nor U10319 (N_10319,N_9520,N_9025);
nor U10320 (N_10320,N_9123,N_8668);
and U10321 (N_10321,N_8712,N_9449);
nor U10322 (N_10322,N_8652,N_9118);
xor U10323 (N_10323,N_9018,N_8997);
and U10324 (N_10324,N_9485,N_9588);
nor U10325 (N_10325,N_9141,N_9396);
or U10326 (N_10326,N_8711,N_9073);
or U10327 (N_10327,N_9016,N_9350);
xor U10328 (N_10328,N_8595,N_8763);
xor U10329 (N_10329,N_9423,N_8716);
nand U10330 (N_10330,N_8648,N_9349);
and U10331 (N_10331,N_8735,N_9580);
nand U10332 (N_10332,N_9393,N_9391);
and U10333 (N_10333,N_8485,N_9051);
nor U10334 (N_10334,N_8546,N_8627);
xor U10335 (N_10335,N_9072,N_8808);
and U10336 (N_10336,N_8537,N_8616);
and U10337 (N_10337,N_8554,N_9253);
nand U10338 (N_10338,N_8608,N_9545);
and U10339 (N_10339,N_8820,N_8760);
nand U10340 (N_10340,N_9129,N_9114);
nand U10341 (N_10341,N_8488,N_8946);
nor U10342 (N_10342,N_9491,N_9394);
and U10343 (N_10343,N_9034,N_8452);
and U10344 (N_10344,N_9484,N_8938);
nor U10345 (N_10345,N_8541,N_8901);
or U10346 (N_10346,N_9398,N_8771);
or U10347 (N_10347,N_8560,N_9244);
or U10348 (N_10348,N_8512,N_8997);
xor U10349 (N_10349,N_9459,N_9302);
or U10350 (N_10350,N_8939,N_9164);
or U10351 (N_10351,N_8694,N_8762);
nand U10352 (N_10352,N_8611,N_9170);
xnor U10353 (N_10353,N_8924,N_8830);
and U10354 (N_10354,N_8469,N_9163);
and U10355 (N_10355,N_8730,N_8946);
nor U10356 (N_10356,N_9489,N_8747);
and U10357 (N_10357,N_9311,N_8421);
or U10358 (N_10358,N_9108,N_9009);
nand U10359 (N_10359,N_9442,N_8476);
xnor U10360 (N_10360,N_9110,N_9449);
and U10361 (N_10361,N_8949,N_8715);
xor U10362 (N_10362,N_9442,N_8953);
xnor U10363 (N_10363,N_8628,N_9092);
or U10364 (N_10364,N_8640,N_9096);
and U10365 (N_10365,N_8941,N_8599);
or U10366 (N_10366,N_8756,N_9182);
or U10367 (N_10367,N_9220,N_8431);
nor U10368 (N_10368,N_9320,N_9101);
xor U10369 (N_10369,N_8409,N_9390);
or U10370 (N_10370,N_8741,N_9141);
or U10371 (N_10371,N_9561,N_9583);
nor U10372 (N_10372,N_8966,N_9104);
and U10373 (N_10373,N_8813,N_9598);
or U10374 (N_10374,N_8654,N_8648);
nand U10375 (N_10375,N_8759,N_8456);
nand U10376 (N_10376,N_9549,N_8744);
and U10377 (N_10377,N_8881,N_9512);
nand U10378 (N_10378,N_8612,N_8702);
and U10379 (N_10379,N_8788,N_8939);
or U10380 (N_10380,N_9525,N_8834);
and U10381 (N_10381,N_8413,N_8667);
nor U10382 (N_10382,N_8816,N_9559);
nor U10383 (N_10383,N_8462,N_9106);
xnor U10384 (N_10384,N_8650,N_8847);
xnor U10385 (N_10385,N_9531,N_9409);
xnor U10386 (N_10386,N_8624,N_8508);
or U10387 (N_10387,N_8781,N_9530);
and U10388 (N_10388,N_8597,N_8760);
xor U10389 (N_10389,N_9343,N_8499);
nand U10390 (N_10390,N_9018,N_9217);
xor U10391 (N_10391,N_8871,N_9516);
or U10392 (N_10392,N_8491,N_8606);
nand U10393 (N_10393,N_9443,N_8739);
xor U10394 (N_10394,N_9401,N_9001);
or U10395 (N_10395,N_9504,N_9459);
nand U10396 (N_10396,N_9418,N_9429);
xnor U10397 (N_10397,N_8679,N_8460);
and U10398 (N_10398,N_9351,N_9147);
nor U10399 (N_10399,N_8432,N_9591);
nand U10400 (N_10400,N_9529,N_8809);
nor U10401 (N_10401,N_8543,N_9525);
nand U10402 (N_10402,N_9133,N_9152);
or U10403 (N_10403,N_8479,N_9502);
xor U10404 (N_10404,N_9312,N_8706);
xor U10405 (N_10405,N_9241,N_8527);
xor U10406 (N_10406,N_9083,N_9148);
or U10407 (N_10407,N_8414,N_9551);
and U10408 (N_10408,N_9566,N_9441);
nor U10409 (N_10409,N_9366,N_8948);
nand U10410 (N_10410,N_8974,N_9469);
xnor U10411 (N_10411,N_8760,N_8835);
nor U10412 (N_10412,N_9430,N_9277);
xor U10413 (N_10413,N_9094,N_9496);
or U10414 (N_10414,N_8789,N_8568);
and U10415 (N_10415,N_9043,N_9312);
and U10416 (N_10416,N_9325,N_8451);
nor U10417 (N_10417,N_8517,N_9423);
nor U10418 (N_10418,N_8681,N_9498);
and U10419 (N_10419,N_8650,N_9401);
nand U10420 (N_10420,N_8720,N_9059);
nor U10421 (N_10421,N_9506,N_8672);
xor U10422 (N_10422,N_8457,N_9308);
xnor U10423 (N_10423,N_9288,N_9311);
nor U10424 (N_10424,N_8540,N_8528);
nor U10425 (N_10425,N_8533,N_9367);
and U10426 (N_10426,N_9355,N_8785);
xnor U10427 (N_10427,N_8460,N_9063);
or U10428 (N_10428,N_8734,N_8768);
and U10429 (N_10429,N_9161,N_9159);
or U10430 (N_10430,N_8737,N_8965);
and U10431 (N_10431,N_9589,N_8849);
xor U10432 (N_10432,N_9044,N_8910);
nand U10433 (N_10433,N_8835,N_8737);
and U10434 (N_10434,N_9277,N_9018);
and U10435 (N_10435,N_9495,N_8449);
and U10436 (N_10436,N_8475,N_8847);
xor U10437 (N_10437,N_9238,N_9149);
nor U10438 (N_10438,N_9483,N_9226);
or U10439 (N_10439,N_9462,N_9246);
and U10440 (N_10440,N_9333,N_9373);
or U10441 (N_10441,N_9315,N_9347);
nand U10442 (N_10442,N_9178,N_9387);
xnor U10443 (N_10443,N_8802,N_8510);
nand U10444 (N_10444,N_8620,N_9050);
xor U10445 (N_10445,N_8471,N_9203);
and U10446 (N_10446,N_8649,N_8546);
nand U10447 (N_10447,N_8641,N_8962);
xnor U10448 (N_10448,N_9214,N_8846);
nor U10449 (N_10449,N_9264,N_9254);
and U10450 (N_10450,N_9518,N_9028);
nand U10451 (N_10451,N_8607,N_8956);
and U10452 (N_10452,N_9002,N_9143);
nand U10453 (N_10453,N_9087,N_9197);
or U10454 (N_10454,N_9360,N_9452);
or U10455 (N_10455,N_9063,N_9369);
nor U10456 (N_10456,N_9070,N_9325);
nor U10457 (N_10457,N_8502,N_9139);
nor U10458 (N_10458,N_8664,N_8935);
xnor U10459 (N_10459,N_9023,N_8903);
nor U10460 (N_10460,N_8668,N_8991);
and U10461 (N_10461,N_8862,N_8489);
xor U10462 (N_10462,N_8708,N_8986);
or U10463 (N_10463,N_9490,N_9154);
and U10464 (N_10464,N_8530,N_8775);
nand U10465 (N_10465,N_8793,N_9536);
nor U10466 (N_10466,N_9589,N_9257);
nand U10467 (N_10467,N_9297,N_9035);
nand U10468 (N_10468,N_8958,N_9365);
and U10469 (N_10469,N_9079,N_9423);
nand U10470 (N_10470,N_9506,N_8436);
xor U10471 (N_10471,N_9221,N_8999);
or U10472 (N_10472,N_9173,N_9565);
and U10473 (N_10473,N_9580,N_8514);
and U10474 (N_10474,N_8710,N_9073);
xor U10475 (N_10475,N_8407,N_9457);
nand U10476 (N_10476,N_9555,N_8755);
and U10477 (N_10477,N_9408,N_8625);
nand U10478 (N_10478,N_9112,N_9366);
or U10479 (N_10479,N_9521,N_9526);
nand U10480 (N_10480,N_9260,N_9575);
nand U10481 (N_10481,N_9191,N_8793);
xor U10482 (N_10482,N_9319,N_9400);
and U10483 (N_10483,N_9060,N_8629);
nand U10484 (N_10484,N_8402,N_8923);
and U10485 (N_10485,N_9105,N_8903);
and U10486 (N_10486,N_9018,N_9469);
or U10487 (N_10487,N_8415,N_8509);
and U10488 (N_10488,N_9511,N_8604);
or U10489 (N_10489,N_9518,N_9550);
nand U10490 (N_10490,N_9585,N_9332);
nand U10491 (N_10491,N_8932,N_8914);
nor U10492 (N_10492,N_9049,N_8619);
xnor U10493 (N_10493,N_8647,N_9011);
nor U10494 (N_10494,N_8885,N_8877);
or U10495 (N_10495,N_8436,N_9193);
nor U10496 (N_10496,N_8923,N_9457);
nor U10497 (N_10497,N_8743,N_8525);
nor U10498 (N_10498,N_8708,N_8523);
or U10499 (N_10499,N_9151,N_8675);
nor U10500 (N_10500,N_9357,N_9132);
nor U10501 (N_10501,N_9232,N_8801);
nor U10502 (N_10502,N_8883,N_9351);
xor U10503 (N_10503,N_8645,N_8942);
nor U10504 (N_10504,N_9054,N_8441);
nor U10505 (N_10505,N_8619,N_8585);
or U10506 (N_10506,N_8928,N_8677);
or U10507 (N_10507,N_9511,N_9453);
or U10508 (N_10508,N_8479,N_8735);
and U10509 (N_10509,N_9043,N_8990);
or U10510 (N_10510,N_9505,N_9430);
nand U10511 (N_10511,N_8751,N_8404);
or U10512 (N_10512,N_8643,N_8543);
nand U10513 (N_10513,N_9029,N_9521);
xnor U10514 (N_10514,N_8455,N_8674);
xor U10515 (N_10515,N_9571,N_8435);
or U10516 (N_10516,N_8537,N_8881);
or U10517 (N_10517,N_8792,N_9399);
xnor U10518 (N_10518,N_9271,N_8568);
nor U10519 (N_10519,N_8718,N_8748);
nand U10520 (N_10520,N_8474,N_9498);
xnor U10521 (N_10521,N_9334,N_8680);
nand U10522 (N_10522,N_9177,N_9294);
xor U10523 (N_10523,N_8800,N_9490);
and U10524 (N_10524,N_8687,N_9118);
nor U10525 (N_10525,N_9320,N_8641);
nand U10526 (N_10526,N_9215,N_9197);
and U10527 (N_10527,N_8481,N_9415);
nand U10528 (N_10528,N_8446,N_9183);
nand U10529 (N_10529,N_8798,N_9007);
or U10530 (N_10530,N_8747,N_8787);
and U10531 (N_10531,N_9207,N_8847);
nand U10532 (N_10532,N_8662,N_8712);
xor U10533 (N_10533,N_8854,N_9526);
and U10534 (N_10534,N_9268,N_9263);
nand U10535 (N_10535,N_8806,N_9081);
nand U10536 (N_10536,N_8567,N_8895);
or U10537 (N_10537,N_8810,N_9140);
or U10538 (N_10538,N_9376,N_9039);
nor U10539 (N_10539,N_9258,N_9269);
and U10540 (N_10540,N_9084,N_9211);
and U10541 (N_10541,N_9078,N_8579);
xor U10542 (N_10542,N_8593,N_9314);
nand U10543 (N_10543,N_8946,N_8896);
nand U10544 (N_10544,N_8777,N_8659);
and U10545 (N_10545,N_9289,N_8863);
and U10546 (N_10546,N_9022,N_9569);
or U10547 (N_10547,N_8523,N_9143);
xnor U10548 (N_10548,N_9464,N_8961);
or U10549 (N_10549,N_9458,N_9192);
xnor U10550 (N_10550,N_8901,N_8520);
nand U10551 (N_10551,N_9494,N_9251);
nor U10552 (N_10552,N_8869,N_9565);
and U10553 (N_10553,N_8880,N_8662);
and U10554 (N_10554,N_8431,N_8804);
xor U10555 (N_10555,N_8457,N_8815);
xor U10556 (N_10556,N_9113,N_8651);
nand U10557 (N_10557,N_9002,N_8563);
nand U10558 (N_10558,N_8894,N_8625);
nor U10559 (N_10559,N_9505,N_8961);
nand U10560 (N_10560,N_8880,N_8781);
nand U10561 (N_10561,N_8994,N_8920);
or U10562 (N_10562,N_8486,N_9385);
xor U10563 (N_10563,N_9463,N_9224);
and U10564 (N_10564,N_9354,N_9431);
nor U10565 (N_10565,N_8545,N_8602);
xor U10566 (N_10566,N_8515,N_9438);
xor U10567 (N_10567,N_9002,N_8885);
nand U10568 (N_10568,N_9183,N_9437);
xor U10569 (N_10569,N_9213,N_9403);
xnor U10570 (N_10570,N_9596,N_8900);
or U10571 (N_10571,N_8966,N_9202);
nand U10572 (N_10572,N_8858,N_8610);
or U10573 (N_10573,N_9143,N_8472);
nand U10574 (N_10574,N_9114,N_9500);
and U10575 (N_10575,N_9206,N_8467);
nand U10576 (N_10576,N_8565,N_8930);
nor U10577 (N_10577,N_9587,N_8923);
nor U10578 (N_10578,N_8915,N_9273);
nor U10579 (N_10579,N_9120,N_9307);
nand U10580 (N_10580,N_9218,N_9499);
xor U10581 (N_10581,N_8617,N_8584);
nand U10582 (N_10582,N_9046,N_9457);
and U10583 (N_10583,N_8421,N_8460);
nor U10584 (N_10584,N_9597,N_9465);
nand U10585 (N_10585,N_8964,N_8888);
nand U10586 (N_10586,N_9248,N_9343);
nor U10587 (N_10587,N_9233,N_8669);
and U10588 (N_10588,N_8762,N_8936);
or U10589 (N_10589,N_8707,N_8740);
nor U10590 (N_10590,N_8475,N_9445);
xnor U10591 (N_10591,N_8622,N_9167);
and U10592 (N_10592,N_9182,N_9149);
xnor U10593 (N_10593,N_9010,N_9119);
nand U10594 (N_10594,N_8608,N_9346);
or U10595 (N_10595,N_9124,N_9100);
nand U10596 (N_10596,N_8799,N_8672);
nor U10597 (N_10597,N_8985,N_9583);
nor U10598 (N_10598,N_8895,N_8623);
xnor U10599 (N_10599,N_9337,N_8965);
xor U10600 (N_10600,N_8747,N_8517);
nand U10601 (N_10601,N_8721,N_9588);
or U10602 (N_10602,N_9536,N_9378);
or U10603 (N_10603,N_8800,N_9027);
nand U10604 (N_10604,N_8506,N_8461);
and U10605 (N_10605,N_9447,N_8729);
nand U10606 (N_10606,N_8404,N_9022);
nor U10607 (N_10607,N_8647,N_8667);
and U10608 (N_10608,N_9457,N_8552);
and U10609 (N_10609,N_9169,N_9015);
nand U10610 (N_10610,N_8857,N_9449);
and U10611 (N_10611,N_9332,N_8516);
or U10612 (N_10612,N_8863,N_8762);
or U10613 (N_10613,N_8775,N_9121);
or U10614 (N_10614,N_9148,N_8564);
xor U10615 (N_10615,N_8517,N_8742);
nor U10616 (N_10616,N_9518,N_9525);
and U10617 (N_10617,N_9193,N_8852);
nor U10618 (N_10618,N_8910,N_9124);
and U10619 (N_10619,N_8968,N_9455);
xor U10620 (N_10620,N_9379,N_9466);
xnor U10621 (N_10621,N_8695,N_9016);
nand U10622 (N_10622,N_9442,N_8850);
nand U10623 (N_10623,N_9032,N_8978);
xor U10624 (N_10624,N_9116,N_9488);
nand U10625 (N_10625,N_8700,N_9504);
nor U10626 (N_10626,N_9512,N_8490);
nand U10627 (N_10627,N_8690,N_9346);
nand U10628 (N_10628,N_8950,N_9425);
or U10629 (N_10629,N_8811,N_8501);
xnor U10630 (N_10630,N_9303,N_8937);
xnor U10631 (N_10631,N_9572,N_9374);
xnor U10632 (N_10632,N_8470,N_9559);
xnor U10633 (N_10633,N_8956,N_8826);
xnor U10634 (N_10634,N_9446,N_9018);
or U10635 (N_10635,N_8724,N_8614);
nand U10636 (N_10636,N_9399,N_9428);
nand U10637 (N_10637,N_9387,N_8648);
or U10638 (N_10638,N_8735,N_9404);
nand U10639 (N_10639,N_8686,N_9491);
nor U10640 (N_10640,N_9120,N_8878);
or U10641 (N_10641,N_9471,N_9338);
and U10642 (N_10642,N_9582,N_9158);
nor U10643 (N_10643,N_9544,N_9355);
xnor U10644 (N_10644,N_9298,N_9005);
nor U10645 (N_10645,N_8738,N_9048);
nor U10646 (N_10646,N_8833,N_8508);
or U10647 (N_10647,N_8416,N_8484);
or U10648 (N_10648,N_8796,N_9161);
nand U10649 (N_10649,N_9439,N_9434);
or U10650 (N_10650,N_9112,N_9388);
nor U10651 (N_10651,N_9185,N_9315);
and U10652 (N_10652,N_8514,N_8772);
xor U10653 (N_10653,N_8954,N_8889);
xnor U10654 (N_10654,N_8635,N_8529);
xor U10655 (N_10655,N_8633,N_9239);
and U10656 (N_10656,N_8792,N_9187);
and U10657 (N_10657,N_8948,N_8870);
nand U10658 (N_10658,N_8688,N_9278);
and U10659 (N_10659,N_8724,N_8998);
nor U10660 (N_10660,N_8450,N_9009);
or U10661 (N_10661,N_8515,N_8454);
xnor U10662 (N_10662,N_8894,N_8493);
nor U10663 (N_10663,N_9013,N_8857);
or U10664 (N_10664,N_8971,N_8429);
nand U10665 (N_10665,N_8657,N_8532);
xor U10666 (N_10666,N_9492,N_8483);
and U10667 (N_10667,N_9250,N_9038);
nand U10668 (N_10668,N_8904,N_8702);
nor U10669 (N_10669,N_9345,N_9594);
nand U10670 (N_10670,N_9405,N_8649);
xnor U10671 (N_10671,N_9058,N_8877);
or U10672 (N_10672,N_9264,N_8838);
and U10673 (N_10673,N_9275,N_8794);
nand U10674 (N_10674,N_9581,N_9185);
nand U10675 (N_10675,N_8767,N_9376);
nand U10676 (N_10676,N_9160,N_9287);
nand U10677 (N_10677,N_8692,N_8835);
nor U10678 (N_10678,N_9177,N_9363);
nor U10679 (N_10679,N_9585,N_9291);
nor U10680 (N_10680,N_8781,N_9295);
or U10681 (N_10681,N_9375,N_8525);
xor U10682 (N_10682,N_9556,N_8782);
and U10683 (N_10683,N_8659,N_8990);
and U10684 (N_10684,N_8735,N_8450);
and U10685 (N_10685,N_9416,N_9122);
nand U10686 (N_10686,N_8516,N_8433);
and U10687 (N_10687,N_8829,N_8535);
nand U10688 (N_10688,N_9035,N_9005);
nand U10689 (N_10689,N_9462,N_8578);
nor U10690 (N_10690,N_8586,N_9488);
or U10691 (N_10691,N_8922,N_8652);
nor U10692 (N_10692,N_8565,N_9252);
xor U10693 (N_10693,N_9103,N_8951);
nand U10694 (N_10694,N_8999,N_9120);
nand U10695 (N_10695,N_8868,N_8405);
xor U10696 (N_10696,N_8766,N_8786);
and U10697 (N_10697,N_8713,N_9054);
or U10698 (N_10698,N_9106,N_9071);
or U10699 (N_10699,N_9280,N_8588);
and U10700 (N_10700,N_8737,N_8868);
nor U10701 (N_10701,N_9246,N_8894);
nand U10702 (N_10702,N_9087,N_8498);
or U10703 (N_10703,N_9135,N_8499);
xor U10704 (N_10704,N_8629,N_9308);
and U10705 (N_10705,N_9556,N_8682);
xor U10706 (N_10706,N_9219,N_9097);
nor U10707 (N_10707,N_9320,N_9301);
and U10708 (N_10708,N_8616,N_9179);
and U10709 (N_10709,N_9487,N_8883);
or U10710 (N_10710,N_8968,N_8587);
nand U10711 (N_10711,N_8704,N_8856);
xnor U10712 (N_10712,N_8641,N_8405);
or U10713 (N_10713,N_9369,N_9484);
nor U10714 (N_10714,N_8599,N_8677);
nand U10715 (N_10715,N_8906,N_8840);
and U10716 (N_10716,N_8865,N_9062);
and U10717 (N_10717,N_8868,N_8974);
nor U10718 (N_10718,N_9529,N_8669);
or U10719 (N_10719,N_8549,N_9332);
nand U10720 (N_10720,N_8657,N_8839);
nor U10721 (N_10721,N_8841,N_9030);
or U10722 (N_10722,N_9526,N_8682);
xnor U10723 (N_10723,N_9224,N_8571);
nor U10724 (N_10724,N_9383,N_9410);
nor U10725 (N_10725,N_9343,N_9166);
nand U10726 (N_10726,N_8694,N_8710);
or U10727 (N_10727,N_9286,N_9027);
nand U10728 (N_10728,N_8867,N_8912);
nand U10729 (N_10729,N_9397,N_8413);
nor U10730 (N_10730,N_9322,N_9409);
or U10731 (N_10731,N_8720,N_8550);
or U10732 (N_10732,N_9501,N_9072);
and U10733 (N_10733,N_8765,N_8492);
nor U10734 (N_10734,N_8978,N_8903);
and U10735 (N_10735,N_8563,N_8548);
or U10736 (N_10736,N_9032,N_9341);
or U10737 (N_10737,N_9215,N_8801);
and U10738 (N_10738,N_9505,N_8850);
or U10739 (N_10739,N_9533,N_9145);
xor U10740 (N_10740,N_9277,N_8550);
and U10741 (N_10741,N_8578,N_8932);
nor U10742 (N_10742,N_8743,N_8409);
xnor U10743 (N_10743,N_9550,N_9591);
and U10744 (N_10744,N_9051,N_9353);
nor U10745 (N_10745,N_8946,N_9390);
xnor U10746 (N_10746,N_8533,N_8683);
nand U10747 (N_10747,N_8788,N_8687);
nor U10748 (N_10748,N_8880,N_9412);
or U10749 (N_10749,N_9221,N_8425);
nand U10750 (N_10750,N_9132,N_8894);
xor U10751 (N_10751,N_8639,N_8448);
or U10752 (N_10752,N_8413,N_8966);
and U10753 (N_10753,N_8524,N_9055);
and U10754 (N_10754,N_9432,N_8491);
or U10755 (N_10755,N_9010,N_9058);
nor U10756 (N_10756,N_8903,N_9504);
xor U10757 (N_10757,N_8826,N_9331);
and U10758 (N_10758,N_8905,N_9491);
or U10759 (N_10759,N_8736,N_9023);
or U10760 (N_10760,N_9172,N_8499);
nand U10761 (N_10761,N_8491,N_8753);
xnor U10762 (N_10762,N_8471,N_8957);
nand U10763 (N_10763,N_8519,N_9591);
nor U10764 (N_10764,N_9171,N_9054);
and U10765 (N_10765,N_9029,N_9231);
or U10766 (N_10766,N_9005,N_8560);
or U10767 (N_10767,N_8668,N_8479);
nor U10768 (N_10768,N_8960,N_8770);
nor U10769 (N_10769,N_9156,N_8876);
and U10770 (N_10770,N_9195,N_8499);
nand U10771 (N_10771,N_9124,N_8817);
nand U10772 (N_10772,N_9188,N_9468);
xor U10773 (N_10773,N_9438,N_8513);
and U10774 (N_10774,N_9124,N_9177);
nand U10775 (N_10775,N_9460,N_9188);
xor U10776 (N_10776,N_8896,N_9410);
or U10777 (N_10777,N_8705,N_8521);
or U10778 (N_10778,N_9516,N_9565);
and U10779 (N_10779,N_8514,N_8444);
and U10780 (N_10780,N_9171,N_8659);
xnor U10781 (N_10781,N_9259,N_8896);
nand U10782 (N_10782,N_9010,N_8910);
or U10783 (N_10783,N_8604,N_9009);
and U10784 (N_10784,N_8836,N_9100);
nor U10785 (N_10785,N_9121,N_9052);
nand U10786 (N_10786,N_8925,N_8481);
and U10787 (N_10787,N_8505,N_9087);
xor U10788 (N_10788,N_8489,N_8812);
xor U10789 (N_10789,N_9442,N_8761);
nand U10790 (N_10790,N_8441,N_9173);
nor U10791 (N_10791,N_9168,N_9511);
nand U10792 (N_10792,N_9066,N_9011);
or U10793 (N_10793,N_9244,N_9191);
or U10794 (N_10794,N_8755,N_9158);
or U10795 (N_10795,N_8805,N_8524);
and U10796 (N_10796,N_8915,N_8770);
and U10797 (N_10797,N_9194,N_8799);
nand U10798 (N_10798,N_9495,N_9259);
and U10799 (N_10799,N_8977,N_9541);
nand U10800 (N_10800,N_9760,N_9827);
xor U10801 (N_10801,N_10455,N_10593);
or U10802 (N_10802,N_10077,N_10498);
or U10803 (N_10803,N_10645,N_10008);
or U10804 (N_10804,N_10493,N_9955);
xor U10805 (N_10805,N_10391,N_9998);
and U10806 (N_10806,N_10512,N_10641);
or U10807 (N_10807,N_9796,N_10579);
or U10808 (N_10808,N_9606,N_9873);
or U10809 (N_10809,N_10612,N_9954);
or U10810 (N_10810,N_9874,N_9708);
nand U10811 (N_10811,N_9701,N_10603);
or U10812 (N_10812,N_10383,N_9979);
xor U10813 (N_10813,N_10095,N_10470);
nor U10814 (N_10814,N_10447,N_9944);
and U10815 (N_10815,N_10779,N_10179);
and U10816 (N_10816,N_10683,N_9913);
nor U10817 (N_10817,N_10009,N_10476);
nor U10818 (N_10818,N_10350,N_9650);
xor U10819 (N_10819,N_10673,N_10195);
or U10820 (N_10820,N_10301,N_10378);
nand U10821 (N_10821,N_10047,N_10634);
or U10822 (N_10822,N_10463,N_10467);
nand U10823 (N_10823,N_9725,N_9920);
and U10824 (N_10824,N_10252,N_10775);
and U10825 (N_10825,N_9731,N_10002);
and U10826 (N_10826,N_10701,N_10028);
nor U10827 (N_10827,N_9993,N_10040);
and U10828 (N_10828,N_10293,N_10668);
xor U10829 (N_10829,N_9627,N_10187);
or U10830 (N_10830,N_10550,N_9681);
or U10831 (N_10831,N_10073,N_10286);
nor U10832 (N_10832,N_9909,N_9939);
and U10833 (N_10833,N_10652,N_9855);
nand U10834 (N_10834,N_10653,N_9914);
and U10835 (N_10835,N_10680,N_9921);
nor U10836 (N_10836,N_10048,N_10235);
and U10837 (N_10837,N_9859,N_10222);
xor U10838 (N_10838,N_9798,N_10395);
or U10839 (N_10839,N_10224,N_10108);
xor U10840 (N_10840,N_10168,N_10537);
nand U10841 (N_10841,N_10750,N_9750);
xor U10842 (N_10842,N_10400,N_9770);
or U10843 (N_10843,N_9865,N_10558);
and U10844 (N_10844,N_10074,N_10704);
and U10845 (N_10845,N_10128,N_9857);
nor U10846 (N_10846,N_10500,N_10282);
or U10847 (N_10847,N_9705,N_9884);
and U10848 (N_10848,N_9973,N_10297);
and U10849 (N_10849,N_9947,N_10748);
nor U10850 (N_10850,N_10239,N_9726);
nand U10851 (N_10851,N_10072,N_9782);
and U10852 (N_10852,N_10709,N_9600);
nor U10853 (N_10853,N_9890,N_10106);
xor U10854 (N_10854,N_9604,N_9626);
or U10855 (N_10855,N_10244,N_10430);
and U10856 (N_10856,N_10032,N_10180);
xnor U10857 (N_10857,N_9736,N_10515);
and U10858 (N_10858,N_10021,N_10271);
and U10859 (N_10859,N_10156,N_10015);
or U10860 (N_10860,N_10436,N_9856);
nor U10861 (N_10861,N_10481,N_10361);
xnor U10862 (N_10862,N_9641,N_9815);
nand U10863 (N_10863,N_9635,N_10379);
or U10864 (N_10864,N_10534,N_9935);
or U10865 (N_10865,N_9823,N_10377);
nor U10866 (N_10866,N_9622,N_10206);
nor U10867 (N_10867,N_9964,N_10042);
xor U10868 (N_10868,N_10572,N_9612);
or U10869 (N_10869,N_10787,N_10631);
or U10870 (N_10870,N_10205,N_10563);
xnor U10871 (N_10871,N_10650,N_10718);
nor U10872 (N_10872,N_9863,N_10132);
nor U10873 (N_10873,N_10099,N_10774);
or U10874 (N_10874,N_9717,N_10365);
xnor U10875 (N_10875,N_10676,N_10554);
and U10876 (N_10876,N_9832,N_9679);
xnor U10877 (N_10877,N_10675,N_9610);
nor U10878 (N_10878,N_10635,N_9965);
xnor U10879 (N_10879,N_9729,N_10525);
nor U10880 (N_10880,N_10309,N_9879);
nand U10881 (N_10881,N_9766,N_10729);
nor U10882 (N_10882,N_10671,N_10405);
and U10883 (N_10883,N_10279,N_10576);
and U10884 (N_10884,N_10722,N_10566);
or U10885 (N_10885,N_10666,N_9942);
or U10886 (N_10886,N_10411,N_9742);
or U10887 (N_10887,N_9642,N_9945);
and U10888 (N_10888,N_10351,N_10169);
and U10889 (N_10889,N_9958,N_10011);
nor U10890 (N_10890,N_10343,N_10607);
nor U10891 (N_10891,N_9763,N_9999);
and U10892 (N_10892,N_9769,N_10597);
or U10893 (N_10893,N_10109,N_10139);
nand U10894 (N_10894,N_9905,N_10198);
and U10895 (N_10895,N_9715,N_10479);
and U10896 (N_10896,N_10535,N_10575);
and U10897 (N_10897,N_9783,N_9828);
xor U10898 (N_10898,N_10267,N_10539);
nand U10899 (N_10899,N_10532,N_9845);
and U10900 (N_10900,N_10465,N_9632);
nand U10901 (N_10901,N_9806,N_9931);
nor U10902 (N_10902,N_9847,N_9849);
and U10903 (N_10903,N_10204,N_10080);
xnor U10904 (N_10904,N_9946,N_10321);
and U10905 (N_10905,N_10357,N_9688);
or U10906 (N_10906,N_9899,N_9601);
nor U10907 (N_10907,N_9959,N_10258);
nand U10908 (N_10908,N_10273,N_10217);
nor U10909 (N_10909,N_9672,N_10513);
nand U10910 (N_10910,N_10790,N_9619);
and U10911 (N_10911,N_9932,N_10543);
xnor U10912 (N_10912,N_10574,N_9603);
xor U10913 (N_10913,N_10484,N_10150);
or U10914 (N_10914,N_10363,N_10308);
xor U10915 (N_10915,N_10017,N_10210);
nor U10916 (N_10916,N_10211,N_9869);
nor U10917 (N_10917,N_9804,N_10158);
and U10918 (N_10918,N_9822,N_10096);
or U10919 (N_10919,N_9704,N_10278);
and U10920 (N_10920,N_10514,N_10731);
nand U10921 (N_10921,N_9860,N_10107);
nor U10922 (N_10922,N_10589,N_10232);
or U10923 (N_10923,N_10637,N_9677);
nand U10924 (N_10924,N_10414,N_10538);
nor U10925 (N_10925,N_10386,N_9748);
xor U10926 (N_10926,N_10632,N_10753);
nor U10927 (N_10927,N_10622,N_10702);
nor U10928 (N_10928,N_10795,N_10112);
xor U10929 (N_10929,N_9901,N_10705);
nor U10930 (N_10930,N_10591,N_9900);
nand U10931 (N_10931,N_9903,N_10236);
and U10932 (N_10932,N_9662,N_10711);
nand U10933 (N_10933,N_10345,N_9614);
or U10934 (N_10934,N_10006,N_9838);
xor U10935 (N_10935,N_9911,N_10707);
nand U10936 (N_10936,N_10049,N_9776);
xor U10937 (N_10937,N_10508,N_9992);
nor U10938 (N_10938,N_10230,N_10243);
nor U10939 (N_10939,N_9734,N_10636);
or U10940 (N_10940,N_9950,N_10428);
nand U10941 (N_10941,N_10171,N_10600);
or U10942 (N_10942,N_10333,N_9961);
or U10943 (N_10943,N_9738,N_10613);
xor U10944 (N_10944,N_9780,N_10728);
nand U10945 (N_10945,N_10004,N_10005);
and U10946 (N_10946,N_9941,N_10388);
nand U10947 (N_10947,N_10218,N_10261);
nor U10948 (N_10948,N_10220,N_10577);
nor U10949 (N_10949,N_10340,N_10736);
or U10950 (N_10950,N_10324,N_10334);
nor U10951 (N_10951,N_10520,N_10466);
nor U10952 (N_10952,N_9840,N_10755);
nand U10953 (N_10953,N_10689,N_10415);
and U10954 (N_10954,N_10570,N_10254);
or U10955 (N_10955,N_9972,N_10121);
xor U10956 (N_10956,N_10473,N_10366);
and U10957 (N_10957,N_10253,N_10773);
nand U10958 (N_10958,N_10167,N_9669);
nand U10959 (N_10959,N_10506,N_10797);
and U10960 (N_10960,N_10488,N_9803);
xnor U10961 (N_10961,N_10085,N_10541);
or U10962 (N_10962,N_9975,N_9674);
nand U10963 (N_10963,N_10569,N_9970);
nand U10964 (N_10964,N_9943,N_10578);
and U10965 (N_10965,N_9687,N_10056);
and U10966 (N_10966,N_10076,N_10449);
nand U10967 (N_10967,N_10427,N_10276);
or U10968 (N_10968,N_9892,N_10407);
nor U10969 (N_10969,N_10289,N_10588);
nand U10970 (N_10970,N_10014,N_9661);
nand U10971 (N_10971,N_9930,N_10231);
xor U10972 (N_10972,N_10397,N_10010);
nand U10973 (N_10973,N_9984,N_9707);
nand U10974 (N_10974,N_10184,N_10051);
nor U10975 (N_10975,N_9639,N_10348);
nor U10976 (N_10976,N_10522,N_10586);
nor U10977 (N_10977,N_9850,N_9628);
or U10978 (N_10978,N_10759,N_9648);
xor U10979 (N_10979,N_9685,N_10125);
nor U10980 (N_10980,N_10209,N_10780);
nand U10981 (N_10981,N_10502,N_9985);
nor U10982 (N_10982,N_9673,N_9756);
and U10983 (N_10983,N_9989,N_10640);
nand U10984 (N_10984,N_10275,N_10528);
nor U10985 (N_10985,N_9956,N_9741);
xor U10986 (N_10986,N_9667,N_10749);
nor U10987 (N_10987,N_10472,N_10703);
nand U10988 (N_10988,N_10142,N_9907);
nand U10989 (N_10989,N_10082,N_9787);
or U10990 (N_10990,N_10442,N_9781);
xnor U10991 (N_10991,N_10492,N_10130);
and U10992 (N_10992,N_9933,N_10688);
and U10993 (N_10993,N_10098,N_9711);
and U10994 (N_10994,N_10192,N_10262);
nor U10995 (N_10995,N_10068,N_9646);
nor U10996 (N_10996,N_10331,N_9665);
nand U10997 (N_10997,N_10445,N_10059);
or U10998 (N_10998,N_10604,N_10583);
xor U10999 (N_10999,N_9758,N_10092);
nand U11000 (N_11000,N_10227,N_10486);
xnor U11001 (N_11001,N_9929,N_10527);
xor U11002 (N_11002,N_10374,N_9620);
nor U11003 (N_11003,N_9875,N_10186);
or U11004 (N_11004,N_10505,N_10043);
or U11005 (N_11005,N_9802,N_10660);
or U11006 (N_11006,N_9724,N_10406);
nor U11007 (N_11007,N_10560,N_10070);
nand U11008 (N_11008,N_9668,N_10446);
or U11009 (N_11009,N_10299,N_9615);
nor U11010 (N_11010,N_10246,N_10745);
and U11011 (N_11011,N_10475,N_10786);
or U11012 (N_11012,N_10398,N_10369);
and U11013 (N_11013,N_10131,N_10263);
or U11014 (N_11014,N_9767,N_10295);
or U11015 (N_11015,N_9799,N_10744);
and U11016 (N_11016,N_9871,N_10237);
xor U11017 (N_11017,N_10071,N_10437);
nand U11018 (N_11018,N_10152,N_9728);
nand U11019 (N_11019,N_10376,N_9652);
and U11020 (N_11020,N_9866,N_10644);
or U11021 (N_11021,N_10027,N_10385);
or U11022 (N_11022,N_10638,N_9656);
or U11023 (N_11023,N_10402,N_10422);
nor U11024 (N_11024,N_10684,N_9689);
nor U11025 (N_11025,N_9957,N_9877);
nor U11026 (N_11026,N_10435,N_10306);
or U11027 (N_11027,N_9841,N_9691);
or U11028 (N_11028,N_9740,N_10260);
nand U11029 (N_11029,N_9744,N_10228);
nor U11030 (N_11030,N_10274,N_10434);
nand U11031 (N_11031,N_9727,N_9761);
xor U11032 (N_11032,N_9629,N_10384);
nand U11033 (N_11033,N_10245,N_10618);
xnor U11034 (N_11034,N_10240,N_9962);
nand U11035 (N_11035,N_9819,N_10421);
xnor U11036 (N_11036,N_10598,N_10368);
and U11037 (N_11037,N_10328,N_10332);
nor U11038 (N_11038,N_10457,N_10359);
nor U11039 (N_11039,N_10677,N_9700);
or U11040 (N_11040,N_10019,N_10630);
or U11041 (N_11041,N_10234,N_10764);
nor U11042 (N_11042,N_10412,N_10494);
xnor U11043 (N_11043,N_9658,N_10174);
nand U11044 (N_11044,N_9808,N_10061);
nor U11045 (N_11045,N_10667,N_10143);
nor U11046 (N_11046,N_10410,N_10033);
nand U11047 (N_11047,N_10685,N_10471);
xnor U11048 (N_11048,N_10547,N_9854);
and U11049 (N_11049,N_10164,N_10225);
xor U11050 (N_11050,N_10444,N_10392);
nor U11051 (N_11051,N_9853,N_10138);
xnor U11052 (N_11052,N_9926,N_9784);
and U11053 (N_11053,N_10307,N_10100);
or U11054 (N_11054,N_9988,N_9925);
xor U11055 (N_11055,N_9852,N_9671);
or U11056 (N_11056,N_9963,N_9928);
and U11057 (N_11057,N_9816,N_10255);
and U11058 (N_11058,N_10501,N_10113);
or U11059 (N_11059,N_10381,N_10163);
and U11060 (N_11060,N_10140,N_10611);
nor U11061 (N_11061,N_9897,N_10247);
nand U11062 (N_11062,N_10432,N_10456);
or U11063 (N_11063,N_9683,N_10567);
nand U11064 (N_11064,N_10298,N_10416);
nand U11065 (N_11065,N_10248,N_10425);
xnor U11066 (N_11066,N_9699,N_9846);
or U11067 (N_11067,N_10123,N_10585);
nand U11068 (N_11068,N_9790,N_10341);
nor U11069 (N_11069,N_10188,N_10356);
nor U11070 (N_11070,N_10283,N_10511);
nor U11071 (N_11071,N_10018,N_10022);
or U11072 (N_11072,N_10438,N_10453);
or U11073 (N_11073,N_10788,N_10555);
nor U11074 (N_11074,N_9638,N_10347);
nor U11075 (N_11075,N_10686,N_9762);
or U11076 (N_11076,N_9966,N_10418);
nand U11077 (N_11077,N_10281,N_10609);
nor U11078 (N_11078,N_9991,N_9953);
nand U11079 (N_11079,N_10367,N_10656);
xnor U11080 (N_11080,N_9664,N_10647);
nor U11081 (N_11081,N_9647,N_9809);
and U11082 (N_11082,N_10706,N_9971);
nor U11083 (N_11083,N_10497,N_9753);
and U11084 (N_11084,N_9616,N_10672);
and U11085 (N_11085,N_10291,N_9800);
or U11086 (N_11086,N_10290,N_9660);
nor U11087 (N_11087,N_10238,N_10571);
and U11088 (N_11088,N_10208,N_10001);
xnor U11089 (N_11089,N_10399,N_9714);
or U11090 (N_11090,N_10046,N_9980);
xnor U11091 (N_11091,N_9952,N_10215);
nor U11092 (N_11092,N_10531,N_10304);
nand U11093 (N_11093,N_10251,N_10662);
nor U11094 (N_11094,N_10323,N_10646);
nor U11095 (N_11095,N_9654,N_9630);
or U11096 (N_11096,N_9645,N_10117);
and U11097 (N_11097,N_10768,N_10122);
or U11098 (N_11098,N_10483,N_10317);
nor U11099 (N_11099,N_9906,N_9653);
xnor U11100 (N_11100,N_10789,N_10777);
nand U11101 (N_11101,N_10272,N_10480);
or U11102 (N_11102,N_10110,N_9675);
xor U11103 (N_11103,N_10765,N_9842);
nor U11104 (N_11104,N_9960,N_10296);
nand U11105 (N_11105,N_10135,N_9663);
or U11106 (N_11106,N_9657,N_9613);
nor U11107 (N_11107,N_9825,N_9651);
nor U11108 (N_11108,N_10408,N_10714);
nor U11109 (N_11109,N_9730,N_10661);
nand U11110 (N_11110,N_10717,N_10794);
xor U11111 (N_11111,N_10189,N_10573);
nor U11112 (N_11112,N_10423,N_10545);
nor U11113 (N_11113,N_10148,N_9938);
xor U11114 (N_11114,N_9636,N_10770);
and U11115 (N_11115,N_10477,N_10389);
and U11116 (N_11116,N_9775,N_9792);
or U11117 (N_11117,N_10605,N_10325);
nand U11118 (N_11118,N_10249,N_9861);
xor U11119 (N_11119,N_10507,N_10358);
nor U11120 (N_11120,N_10312,N_10199);
nand U11121 (N_11121,N_9888,N_10322);
nand U11122 (N_11122,N_10330,N_10568);
nor U11123 (N_11123,N_10373,N_10758);
nand U11124 (N_11124,N_10337,N_9940);
nand U11125 (N_11125,N_10045,N_10126);
and U11126 (N_11126,N_10104,N_9719);
nand U11127 (N_11127,N_10037,N_10201);
or U11128 (N_11128,N_10387,N_9995);
and U11129 (N_11129,N_10695,N_9755);
and U11130 (N_11130,N_9818,N_10594);
xnor U11131 (N_11131,N_10458,N_10757);
nor U11132 (N_11132,N_9829,N_10499);
or U11133 (N_11133,N_10708,N_10173);
nand U11134 (N_11134,N_10746,N_9634);
nand U11135 (N_11135,N_10221,N_10503);
and U11136 (N_11136,N_10285,N_9895);
and U11137 (N_11137,N_9805,N_10691);
xnor U11138 (N_11138,N_9835,N_10025);
or U11139 (N_11139,N_10185,N_9607);
nor U11140 (N_11140,N_10791,N_9710);
or U11141 (N_11141,N_10101,N_10681);
and U11142 (N_11142,N_10270,N_10546);
nand U11143 (N_11143,N_10735,N_10516);
xnor U11144 (N_11144,N_9735,N_9713);
or U11145 (N_11145,N_10069,N_10733);
nor U11146 (N_11146,N_10065,N_10734);
nor U11147 (N_11147,N_9718,N_10763);
nand U11148 (N_11148,N_9848,N_9749);
xor U11149 (N_11149,N_10687,N_9703);
nor U11150 (N_11150,N_10741,N_9982);
and U11151 (N_11151,N_9678,N_9969);
and U11152 (N_11152,N_10521,N_10219);
and U11153 (N_11153,N_10154,N_10654);
nand U11154 (N_11154,N_10342,N_10581);
nand U11155 (N_11155,N_9870,N_9759);
xor U11156 (N_11156,N_10000,N_10592);
nor U11157 (N_11157,N_10256,N_9771);
nor U11158 (N_11158,N_9886,N_10259);
or U11159 (N_11159,N_9722,N_10196);
or U11160 (N_11160,N_10740,N_10643);
nand U11161 (N_11161,N_10426,N_10338);
or U11162 (N_11162,N_10057,N_10553);
nand U11163 (N_11163,N_10782,N_10084);
xor U11164 (N_11164,N_10316,N_10266);
or U11165 (N_11165,N_10772,N_10716);
and U11166 (N_11166,N_10738,N_9659);
and U11167 (N_11167,N_9797,N_9986);
and U11168 (N_11168,N_10264,N_9893);
nor U11169 (N_11169,N_9751,N_10030);
xor U11170 (N_11170,N_10796,N_9981);
and U11171 (N_11171,N_9680,N_10079);
nor U11172 (N_11172,N_10055,N_10093);
nand U11173 (N_11173,N_9983,N_9793);
nand U11174 (N_11174,N_9623,N_10181);
nand U11175 (N_11175,N_10743,N_10404);
nor U11176 (N_11176,N_10439,N_10336);
nand U11177 (N_11177,N_10754,N_9608);
and U11178 (N_11178,N_9976,N_9994);
or U11179 (N_11179,N_10007,N_9813);
xor U11180 (N_11180,N_10364,N_10360);
or U11181 (N_11181,N_10119,N_10146);
or U11182 (N_11182,N_10719,N_9774);
nor U11183 (N_11183,N_9885,N_10690);
and U11184 (N_11184,N_10064,N_10495);
nor U11185 (N_11185,N_10401,N_9752);
or U11186 (N_11186,N_10088,N_9898);
nor U11187 (N_11187,N_10133,N_9811);
or U11188 (N_11188,N_10023,N_10747);
nor U11189 (N_11189,N_10212,N_9904);
nor U11190 (N_11190,N_10627,N_10781);
nand U11191 (N_11191,N_10024,N_9891);
nor U11192 (N_11192,N_10223,N_10619);
nor U11193 (N_11193,N_10087,N_10161);
and U11194 (N_11194,N_10536,N_10769);
xnor U11195 (N_11195,N_10176,N_9788);
and U11196 (N_11196,N_10648,N_10417);
and U11197 (N_11197,N_10626,N_10191);
nand U11198 (N_11198,N_10320,N_10081);
nor U11199 (N_11199,N_9670,N_10207);
nand U11200 (N_11200,N_10303,N_9785);
or U11201 (N_11201,N_10792,N_10105);
xor U11202 (N_11202,N_10726,N_10052);
and U11203 (N_11203,N_9910,N_9611);
or U11204 (N_11204,N_10120,N_9821);
xor U11205 (N_11205,N_10614,N_10284);
nand U11206 (N_11206,N_10111,N_9912);
nor U11207 (N_11207,N_10776,N_10461);
and U11208 (N_11208,N_10698,N_10443);
and U11209 (N_11209,N_10038,N_9894);
and U11210 (N_11210,N_10440,N_10431);
and U11211 (N_11211,N_10633,N_10710);
nor U11212 (N_11212,N_10041,N_10396);
and U11213 (N_11213,N_10766,N_9990);
nand U11214 (N_11214,N_10382,N_10250);
nor U11215 (N_11215,N_9789,N_9794);
nor U11216 (N_11216,N_10075,N_10193);
nand U11217 (N_11217,N_10696,N_10058);
and U11218 (N_11218,N_10433,N_10663);
nand U11219 (N_11219,N_10557,N_10487);
nor U11220 (N_11220,N_9830,N_10615);
and U11221 (N_11221,N_10370,N_9814);
xor U11222 (N_11222,N_9666,N_9618);
nand U11223 (N_11223,N_10393,N_10664);
nor U11224 (N_11224,N_10756,N_10767);
or U11225 (N_11225,N_10580,N_9737);
nand U11226 (N_11226,N_10134,N_10362);
nand U11227 (N_11227,N_10490,N_10682);
nand U11228 (N_11228,N_10564,N_9694);
and U11229 (N_11229,N_9876,N_10172);
or U11230 (N_11230,N_10327,N_10371);
or U11231 (N_11231,N_10784,N_10464);
nor U11232 (N_11232,N_10468,N_10737);
nand U11233 (N_11233,N_10160,N_10229);
or U11234 (N_11234,N_9836,N_9949);
nor U11235 (N_11235,N_10799,N_10420);
xnor U11236 (N_11236,N_9915,N_10778);
nor U11237 (N_11237,N_10020,N_10147);
or U11238 (N_11238,N_10489,N_10269);
nand U11239 (N_11239,N_9765,N_10524);
and U11240 (N_11240,N_9918,N_10151);
or U11241 (N_11241,N_9698,N_10762);
or U11242 (N_11242,N_10102,N_10116);
nand U11243 (N_11243,N_9851,N_10268);
and U11244 (N_11244,N_9878,N_10413);
nand U11245 (N_11245,N_10561,N_9795);
or U11246 (N_11246,N_10202,N_10451);
and U11247 (N_11247,N_10649,N_10265);
nor U11248 (N_11248,N_10091,N_9643);
and U11249 (N_11249,N_9937,N_10403);
nor U11250 (N_11250,N_9732,N_9917);
or U11251 (N_11251,N_10277,N_10610);
xor U11252 (N_11252,N_9902,N_9690);
and U11253 (N_11253,N_9609,N_9896);
and U11254 (N_11254,N_10694,N_10424);
nand U11255 (N_11255,N_9831,N_10699);
and U11256 (N_11256,N_9702,N_10485);
nor U11257 (N_11257,N_9916,N_10089);
and U11258 (N_11258,N_9843,N_9754);
or U11259 (N_11259,N_9709,N_10036);
xor U11260 (N_11260,N_9936,N_10732);
xnor U11261 (N_11261,N_10136,N_10353);
or U11262 (N_11262,N_9772,N_10329);
nor U11263 (N_11263,N_10302,N_10459);
or U11264 (N_11264,N_9768,N_10016);
nand U11265 (N_11265,N_9605,N_10669);
or U11266 (N_11266,N_10582,N_10542);
or U11267 (N_11267,N_10454,N_10355);
or U11268 (N_11268,N_10044,N_10294);
or U11269 (N_11269,N_9881,N_9839);
nand U11270 (N_11270,N_10165,N_10628);
xnor U11271 (N_11271,N_10751,N_9872);
nand U11272 (N_11272,N_10530,N_10183);
or U11273 (N_11273,N_10203,N_10039);
or U11274 (N_11274,N_10197,N_10599);
or U11275 (N_11275,N_10601,N_9934);
xor U11276 (N_11276,N_10793,N_10724);
and U11277 (N_11277,N_10354,N_10639);
xor U11278 (N_11278,N_10620,N_10310);
nor U11279 (N_11279,N_10190,N_9745);
xnor U11280 (N_11280,N_10606,N_9697);
or U11281 (N_11281,N_10300,N_9621);
xnor U11282 (N_11282,N_10450,N_10114);
or U11283 (N_11283,N_9706,N_10013);
nor U11284 (N_11284,N_10034,N_9834);
nand U11285 (N_11285,N_10390,N_10149);
and U11286 (N_11286,N_10642,N_9977);
and U11287 (N_11287,N_10448,N_9720);
nor U11288 (N_11288,N_9997,N_10692);
nor U11289 (N_11289,N_10651,N_10474);
nand U11290 (N_11290,N_10533,N_9692);
and U11291 (N_11291,N_9743,N_10162);
nor U11292 (N_11292,N_9987,N_10145);
nor U11293 (N_11293,N_10752,N_9649);
nor U11294 (N_11294,N_10452,N_10725);
or U11295 (N_11295,N_10352,N_10409);
xor U11296 (N_11296,N_10509,N_10129);
and U11297 (N_11297,N_10170,N_9746);
xor U11298 (N_11298,N_9862,N_10659);
nand U11299 (N_11299,N_9824,N_10177);
and U11300 (N_11300,N_9625,N_10697);
nor U11301 (N_11301,N_10144,N_10761);
or U11302 (N_11302,N_10380,N_9889);
or U11303 (N_11303,N_10658,N_10318);
or U11304 (N_11304,N_9773,N_9757);
nand U11305 (N_11305,N_9807,N_9624);
and U11306 (N_11306,N_10621,N_9602);
nand U11307 (N_11307,N_10529,N_10315);
and U11308 (N_11308,N_10720,N_9637);
nor U11309 (N_11309,N_10241,N_9721);
and U11310 (N_11310,N_10311,N_9858);
and U11311 (N_11311,N_10257,N_10054);
nand U11312 (N_11312,N_10175,N_10617);
or U11313 (N_11313,N_10590,N_10103);
nor U11314 (N_11314,N_10124,N_10157);
xor U11315 (N_11315,N_10624,N_10549);
or U11316 (N_11316,N_10394,N_10097);
nor U11317 (N_11317,N_9833,N_10504);
xnor U11318 (N_11318,N_10584,N_9922);
xnor U11319 (N_11319,N_10623,N_9974);
or U11320 (N_11320,N_10742,N_10608);
nor U11321 (N_11321,N_9676,N_9844);
and U11322 (N_11322,N_9908,N_9712);
or U11323 (N_11323,N_9864,N_10200);
xnor U11324 (N_11324,N_10288,N_10478);
or U11325 (N_11325,N_10678,N_10115);
nor U11326 (N_11326,N_10596,N_10616);
and U11327 (N_11327,N_10066,N_10771);
nor U11328 (N_11328,N_10326,N_10319);
and U11329 (N_11329,N_9967,N_9655);
or U11330 (N_11330,N_10242,N_10216);
nor U11331 (N_11331,N_9801,N_10213);
xor U11332 (N_11332,N_10785,N_10565);
or U11333 (N_11333,N_9968,N_10141);
nor U11334 (N_11334,N_10625,N_9948);
or U11335 (N_11335,N_10665,N_10556);
or U11336 (N_11336,N_10657,N_10469);
or U11337 (N_11337,N_9786,N_10182);
nand U11338 (N_11338,N_10491,N_10035);
nor U11339 (N_11339,N_10339,N_10783);
or U11340 (N_11340,N_10372,N_9867);
nor U11341 (N_11341,N_10510,N_9686);
and U11342 (N_11342,N_10552,N_10441);
nand U11343 (N_11343,N_9777,N_10559);
and U11344 (N_11344,N_10214,N_9927);
xor U11345 (N_11345,N_9951,N_10517);
and U11346 (N_11346,N_10346,N_10287);
or U11347 (N_11347,N_9779,N_9716);
nand U11348 (N_11348,N_10166,N_9693);
nand U11349 (N_11349,N_10194,N_10562);
xnor U11350 (N_11350,N_10137,N_10602);
nand U11351 (N_11351,N_10280,N_10305);
xor U11352 (N_11352,N_9778,N_9633);
and U11353 (N_11353,N_10153,N_9640);
xnor U11354 (N_11354,N_9723,N_10050);
nand U11355 (N_11355,N_10798,N_10693);
and U11356 (N_11356,N_10062,N_10727);
or U11357 (N_11357,N_9923,N_9747);
and U11358 (N_11358,N_10460,N_10712);
xnor U11359 (N_11359,N_10063,N_10715);
nor U11360 (N_11360,N_10226,N_10730);
nor U11361 (N_11361,N_9868,N_10655);
xnor U11362 (N_11362,N_10349,N_10518);
nand U11363 (N_11363,N_10078,N_9791);
nand U11364 (N_11364,N_9924,N_10094);
xnor U11365 (N_11365,N_10587,N_9919);
xor U11366 (N_11366,N_10540,N_10526);
nand U11367 (N_11367,N_10523,N_9739);
nand U11368 (N_11368,N_9817,N_9810);
and U11369 (N_11369,N_10674,N_10003);
and U11370 (N_11370,N_9631,N_10083);
and U11371 (N_11371,N_10548,N_9820);
xnor U11372 (N_11372,N_10723,N_10713);
xnor U11373 (N_11373,N_10127,N_10012);
and U11374 (N_11374,N_10551,N_9733);
and U11375 (N_11375,N_10544,N_10760);
xnor U11376 (N_11376,N_9812,N_10721);
and U11377 (N_11377,N_10629,N_9978);
nand U11378 (N_11378,N_10314,N_10178);
or U11379 (N_11379,N_9883,N_10233);
nand U11380 (N_11380,N_10679,N_9996);
nor U11381 (N_11381,N_10090,N_10496);
or U11382 (N_11382,N_10053,N_9617);
nand U11383 (N_11383,N_10519,N_10595);
and U11384 (N_11384,N_9764,N_10026);
and U11385 (N_11385,N_9684,N_10155);
and U11386 (N_11386,N_10086,N_9695);
xnor U11387 (N_11387,N_10031,N_9882);
and U11388 (N_11388,N_10462,N_10060);
xor U11389 (N_11389,N_10159,N_10700);
xnor U11390 (N_11390,N_10335,N_9880);
nand U11391 (N_11391,N_9887,N_9682);
nor U11392 (N_11392,N_10067,N_10313);
xnor U11393 (N_11393,N_9826,N_10029);
nand U11394 (N_11394,N_10292,N_10429);
and U11395 (N_11395,N_10670,N_10375);
nor U11396 (N_11396,N_10739,N_10482);
or U11397 (N_11397,N_10419,N_10118);
nand U11398 (N_11398,N_9837,N_9644);
nand U11399 (N_11399,N_10344,N_9696);
nor U11400 (N_11400,N_10668,N_9924);
xnor U11401 (N_11401,N_10385,N_10270);
and U11402 (N_11402,N_9761,N_10561);
nor U11403 (N_11403,N_9701,N_10713);
nor U11404 (N_11404,N_9697,N_10776);
or U11405 (N_11405,N_10478,N_9707);
nand U11406 (N_11406,N_10187,N_10206);
and U11407 (N_11407,N_10559,N_10702);
nand U11408 (N_11408,N_9858,N_10682);
and U11409 (N_11409,N_10198,N_9873);
nand U11410 (N_11410,N_9895,N_9617);
xnor U11411 (N_11411,N_10761,N_10626);
and U11412 (N_11412,N_10639,N_10706);
nor U11413 (N_11413,N_10363,N_10524);
xnor U11414 (N_11414,N_10426,N_9979);
xor U11415 (N_11415,N_10772,N_10529);
nand U11416 (N_11416,N_9899,N_10060);
and U11417 (N_11417,N_10177,N_10481);
and U11418 (N_11418,N_10214,N_10296);
nand U11419 (N_11419,N_9753,N_10080);
nand U11420 (N_11420,N_10480,N_10131);
nor U11421 (N_11421,N_9905,N_10257);
and U11422 (N_11422,N_10750,N_10352);
or U11423 (N_11423,N_10399,N_10688);
or U11424 (N_11424,N_10376,N_10409);
and U11425 (N_11425,N_9675,N_9742);
xor U11426 (N_11426,N_9752,N_10062);
and U11427 (N_11427,N_9948,N_9713);
nor U11428 (N_11428,N_9654,N_10363);
xnor U11429 (N_11429,N_10202,N_10146);
xnor U11430 (N_11430,N_10304,N_10590);
nor U11431 (N_11431,N_10284,N_10424);
nor U11432 (N_11432,N_10754,N_9639);
nor U11433 (N_11433,N_10106,N_10259);
nor U11434 (N_11434,N_10297,N_10181);
nand U11435 (N_11435,N_10334,N_9948);
and U11436 (N_11436,N_10569,N_9966);
nand U11437 (N_11437,N_10234,N_9891);
and U11438 (N_11438,N_9888,N_9820);
and U11439 (N_11439,N_10392,N_10312);
and U11440 (N_11440,N_10346,N_9983);
nor U11441 (N_11441,N_10139,N_10163);
or U11442 (N_11442,N_9774,N_10285);
and U11443 (N_11443,N_10314,N_9737);
nor U11444 (N_11444,N_10017,N_10270);
and U11445 (N_11445,N_10444,N_9753);
or U11446 (N_11446,N_9717,N_10416);
nor U11447 (N_11447,N_9778,N_9689);
xnor U11448 (N_11448,N_9793,N_9756);
or U11449 (N_11449,N_9614,N_10015);
and U11450 (N_11450,N_10406,N_10737);
and U11451 (N_11451,N_10361,N_9824);
xnor U11452 (N_11452,N_10185,N_10225);
and U11453 (N_11453,N_9679,N_10780);
xnor U11454 (N_11454,N_10343,N_9639);
and U11455 (N_11455,N_10652,N_9702);
or U11456 (N_11456,N_10583,N_10183);
nand U11457 (N_11457,N_10494,N_9760);
and U11458 (N_11458,N_10120,N_10527);
or U11459 (N_11459,N_9851,N_10616);
nor U11460 (N_11460,N_10607,N_10226);
and U11461 (N_11461,N_9924,N_10595);
nor U11462 (N_11462,N_10505,N_10032);
xnor U11463 (N_11463,N_10215,N_10660);
or U11464 (N_11464,N_9607,N_10139);
and U11465 (N_11465,N_10369,N_10419);
or U11466 (N_11466,N_9730,N_10079);
and U11467 (N_11467,N_10495,N_9986);
and U11468 (N_11468,N_10169,N_9705);
xnor U11469 (N_11469,N_10507,N_10253);
or U11470 (N_11470,N_9882,N_10648);
xnor U11471 (N_11471,N_10034,N_10739);
xor U11472 (N_11472,N_9677,N_9777);
nor U11473 (N_11473,N_10164,N_9962);
xor U11474 (N_11474,N_10684,N_10516);
nand U11475 (N_11475,N_10304,N_9947);
nand U11476 (N_11476,N_10393,N_10470);
nand U11477 (N_11477,N_10716,N_10391);
and U11478 (N_11478,N_9993,N_9986);
and U11479 (N_11479,N_10090,N_10546);
nand U11480 (N_11480,N_10645,N_9994);
nor U11481 (N_11481,N_10374,N_10601);
nand U11482 (N_11482,N_10686,N_9988);
nor U11483 (N_11483,N_10709,N_10331);
nand U11484 (N_11484,N_10269,N_10783);
nand U11485 (N_11485,N_9872,N_10008);
or U11486 (N_11486,N_10382,N_10211);
or U11487 (N_11487,N_10250,N_10601);
and U11488 (N_11488,N_9842,N_10211);
or U11489 (N_11489,N_10639,N_9725);
or U11490 (N_11490,N_9948,N_10563);
xor U11491 (N_11491,N_10401,N_10506);
and U11492 (N_11492,N_10195,N_10598);
and U11493 (N_11493,N_10278,N_9929);
nor U11494 (N_11494,N_10494,N_10164);
nand U11495 (N_11495,N_10647,N_9940);
xnor U11496 (N_11496,N_10770,N_10657);
xor U11497 (N_11497,N_9650,N_10721);
or U11498 (N_11498,N_9779,N_10606);
and U11499 (N_11499,N_10081,N_10299);
xor U11500 (N_11500,N_10636,N_10306);
or U11501 (N_11501,N_9886,N_10494);
and U11502 (N_11502,N_9978,N_9606);
nor U11503 (N_11503,N_10270,N_10222);
and U11504 (N_11504,N_10232,N_10703);
or U11505 (N_11505,N_9694,N_9943);
and U11506 (N_11506,N_9810,N_10175);
nor U11507 (N_11507,N_10497,N_9650);
nor U11508 (N_11508,N_9627,N_10076);
and U11509 (N_11509,N_10643,N_9892);
and U11510 (N_11510,N_10515,N_10110);
nor U11511 (N_11511,N_10459,N_10026);
nor U11512 (N_11512,N_10149,N_9811);
nand U11513 (N_11513,N_10031,N_10456);
and U11514 (N_11514,N_9892,N_10281);
nand U11515 (N_11515,N_10604,N_10662);
xnor U11516 (N_11516,N_10072,N_9692);
or U11517 (N_11517,N_9689,N_10215);
nand U11518 (N_11518,N_10330,N_10087);
or U11519 (N_11519,N_10098,N_10464);
xor U11520 (N_11520,N_10276,N_10046);
nor U11521 (N_11521,N_9986,N_10021);
nor U11522 (N_11522,N_9993,N_9760);
or U11523 (N_11523,N_9719,N_9926);
or U11524 (N_11524,N_10560,N_10026);
xnor U11525 (N_11525,N_10502,N_10155);
nand U11526 (N_11526,N_10499,N_10648);
nor U11527 (N_11527,N_10029,N_10427);
nand U11528 (N_11528,N_10523,N_10564);
or U11529 (N_11529,N_10313,N_10175);
nor U11530 (N_11530,N_10449,N_9733);
xnor U11531 (N_11531,N_10136,N_10652);
nor U11532 (N_11532,N_9653,N_10549);
xnor U11533 (N_11533,N_10457,N_9852);
nand U11534 (N_11534,N_10321,N_10758);
nand U11535 (N_11535,N_9996,N_10095);
nor U11536 (N_11536,N_10641,N_10503);
nor U11537 (N_11537,N_9633,N_10738);
nor U11538 (N_11538,N_10606,N_10198);
nand U11539 (N_11539,N_10385,N_10485);
xor U11540 (N_11540,N_10698,N_10284);
nor U11541 (N_11541,N_10197,N_9993);
nor U11542 (N_11542,N_10274,N_10012);
xor U11543 (N_11543,N_10360,N_10745);
and U11544 (N_11544,N_10510,N_10709);
nand U11545 (N_11545,N_10509,N_10578);
xnor U11546 (N_11546,N_9728,N_10035);
or U11547 (N_11547,N_9882,N_10392);
nand U11548 (N_11548,N_9952,N_10036);
nor U11549 (N_11549,N_10550,N_10447);
nor U11550 (N_11550,N_9607,N_10518);
or U11551 (N_11551,N_9975,N_10352);
nor U11552 (N_11552,N_9894,N_9801);
or U11553 (N_11553,N_9973,N_9766);
and U11554 (N_11554,N_10531,N_10599);
xnor U11555 (N_11555,N_10155,N_10723);
nand U11556 (N_11556,N_10561,N_10330);
nor U11557 (N_11557,N_10513,N_9944);
nand U11558 (N_11558,N_10031,N_10087);
nand U11559 (N_11559,N_10191,N_10274);
and U11560 (N_11560,N_10705,N_10435);
nand U11561 (N_11561,N_9769,N_10339);
xor U11562 (N_11562,N_10348,N_10063);
xnor U11563 (N_11563,N_10180,N_10475);
xnor U11564 (N_11564,N_9609,N_10289);
and U11565 (N_11565,N_10729,N_10065);
and U11566 (N_11566,N_9703,N_10781);
nor U11567 (N_11567,N_9623,N_10543);
nor U11568 (N_11568,N_10146,N_10262);
nand U11569 (N_11569,N_10586,N_9777);
and U11570 (N_11570,N_10754,N_10253);
and U11571 (N_11571,N_9667,N_9896);
xnor U11572 (N_11572,N_9618,N_10153);
nand U11573 (N_11573,N_10509,N_9920);
nor U11574 (N_11574,N_10703,N_10714);
nand U11575 (N_11575,N_10028,N_10360);
nand U11576 (N_11576,N_9621,N_10429);
nand U11577 (N_11577,N_10147,N_10176);
xnor U11578 (N_11578,N_10225,N_10090);
nor U11579 (N_11579,N_10473,N_9847);
or U11580 (N_11580,N_9877,N_10141);
and U11581 (N_11581,N_10453,N_9859);
nor U11582 (N_11582,N_9751,N_10169);
and U11583 (N_11583,N_10185,N_10692);
or U11584 (N_11584,N_9691,N_9802);
or U11585 (N_11585,N_10138,N_10206);
and U11586 (N_11586,N_9680,N_10765);
or U11587 (N_11587,N_10215,N_10395);
xor U11588 (N_11588,N_10509,N_9913);
xnor U11589 (N_11589,N_10496,N_9856);
nand U11590 (N_11590,N_10419,N_10459);
xor U11591 (N_11591,N_10381,N_10185);
nand U11592 (N_11592,N_9916,N_10094);
and U11593 (N_11593,N_10396,N_10002);
nor U11594 (N_11594,N_10576,N_10603);
nor U11595 (N_11595,N_10282,N_9684);
nand U11596 (N_11596,N_10304,N_10617);
or U11597 (N_11597,N_10562,N_10345);
xnor U11598 (N_11598,N_10424,N_10124);
nand U11599 (N_11599,N_10139,N_10100);
nand U11600 (N_11600,N_10099,N_10710);
nand U11601 (N_11601,N_9738,N_10477);
and U11602 (N_11602,N_10625,N_10661);
or U11603 (N_11603,N_10523,N_9763);
xnor U11604 (N_11604,N_10105,N_9764);
xnor U11605 (N_11605,N_9863,N_10729);
nor U11606 (N_11606,N_10705,N_9708);
or U11607 (N_11607,N_9957,N_9918);
nor U11608 (N_11608,N_9706,N_10353);
nor U11609 (N_11609,N_10146,N_10329);
nor U11610 (N_11610,N_9680,N_9763);
nand U11611 (N_11611,N_10216,N_9640);
or U11612 (N_11612,N_10565,N_10182);
xor U11613 (N_11613,N_10342,N_10763);
nor U11614 (N_11614,N_10498,N_10696);
nor U11615 (N_11615,N_10123,N_9815);
or U11616 (N_11616,N_10139,N_10702);
nor U11617 (N_11617,N_9651,N_10230);
xor U11618 (N_11618,N_10394,N_9739);
and U11619 (N_11619,N_10280,N_9735);
xor U11620 (N_11620,N_10359,N_9662);
or U11621 (N_11621,N_10475,N_10170);
and U11622 (N_11622,N_10202,N_10585);
nor U11623 (N_11623,N_10180,N_10438);
or U11624 (N_11624,N_9645,N_10493);
or U11625 (N_11625,N_9902,N_10463);
xnor U11626 (N_11626,N_9681,N_10759);
and U11627 (N_11627,N_9700,N_10371);
xor U11628 (N_11628,N_9905,N_10204);
and U11629 (N_11629,N_10751,N_10381);
and U11630 (N_11630,N_9874,N_9962);
and U11631 (N_11631,N_10123,N_10279);
nand U11632 (N_11632,N_10741,N_9790);
nand U11633 (N_11633,N_10448,N_10038);
xnor U11634 (N_11634,N_9902,N_9882);
nand U11635 (N_11635,N_10196,N_10749);
or U11636 (N_11636,N_10165,N_10222);
and U11637 (N_11637,N_9660,N_9954);
nor U11638 (N_11638,N_10509,N_10345);
and U11639 (N_11639,N_9909,N_10633);
or U11640 (N_11640,N_10591,N_10266);
nor U11641 (N_11641,N_10523,N_9803);
nand U11642 (N_11642,N_10530,N_10787);
xnor U11643 (N_11643,N_9653,N_9661);
xnor U11644 (N_11644,N_10473,N_10754);
nor U11645 (N_11645,N_9636,N_10137);
nor U11646 (N_11646,N_10478,N_9651);
xor U11647 (N_11647,N_10096,N_9987);
or U11648 (N_11648,N_9958,N_10479);
or U11649 (N_11649,N_10592,N_10539);
or U11650 (N_11650,N_10151,N_9976);
and U11651 (N_11651,N_10035,N_10010);
or U11652 (N_11652,N_10040,N_10630);
nor U11653 (N_11653,N_10001,N_9700);
nor U11654 (N_11654,N_10612,N_10703);
or U11655 (N_11655,N_9909,N_10711);
nand U11656 (N_11656,N_9865,N_9843);
xor U11657 (N_11657,N_9708,N_10502);
nand U11658 (N_11658,N_9678,N_10768);
or U11659 (N_11659,N_9755,N_10072);
xnor U11660 (N_11660,N_10208,N_9662);
nor U11661 (N_11661,N_10770,N_9894);
and U11662 (N_11662,N_9977,N_10195);
xnor U11663 (N_11663,N_9744,N_9604);
nand U11664 (N_11664,N_9658,N_10100);
nand U11665 (N_11665,N_10615,N_10351);
and U11666 (N_11666,N_10711,N_10585);
nand U11667 (N_11667,N_9653,N_9800);
nor U11668 (N_11668,N_9853,N_9780);
and U11669 (N_11669,N_10171,N_10213);
and U11670 (N_11670,N_10193,N_10502);
nand U11671 (N_11671,N_10381,N_10412);
nor U11672 (N_11672,N_10569,N_9879);
and U11673 (N_11673,N_9858,N_9635);
or U11674 (N_11674,N_9675,N_10623);
nand U11675 (N_11675,N_10789,N_9668);
and U11676 (N_11676,N_10426,N_9998);
or U11677 (N_11677,N_10662,N_10587);
xor U11678 (N_11678,N_9866,N_9999);
nand U11679 (N_11679,N_9660,N_10726);
xnor U11680 (N_11680,N_10050,N_10454);
and U11681 (N_11681,N_10681,N_10589);
and U11682 (N_11682,N_9859,N_10739);
nand U11683 (N_11683,N_10375,N_10044);
nand U11684 (N_11684,N_9605,N_10407);
nand U11685 (N_11685,N_10003,N_9917);
or U11686 (N_11686,N_10562,N_10408);
or U11687 (N_11687,N_9897,N_10785);
or U11688 (N_11688,N_9749,N_10092);
and U11689 (N_11689,N_9655,N_9676);
xor U11690 (N_11690,N_10482,N_9804);
or U11691 (N_11691,N_10034,N_10770);
xor U11692 (N_11692,N_10742,N_9703);
xor U11693 (N_11693,N_9982,N_9669);
or U11694 (N_11694,N_9849,N_9963);
nor U11695 (N_11695,N_9793,N_9740);
xor U11696 (N_11696,N_9996,N_10425);
nor U11697 (N_11697,N_9871,N_9684);
or U11698 (N_11698,N_10354,N_10723);
or U11699 (N_11699,N_10734,N_9647);
nor U11700 (N_11700,N_10090,N_10713);
xnor U11701 (N_11701,N_10151,N_10772);
nor U11702 (N_11702,N_10372,N_10000);
nand U11703 (N_11703,N_10689,N_10469);
nand U11704 (N_11704,N_10574,N_10215);
and U11705 (N_11705,N_10770,N_10605);
nor U11706 (N_11706,N_9877,N_10384);
nor U11707 (N_11707,N_9980,N_10702);
nor U11708 (N_11708,N_9889,N_9987);
or U11709 (N_11709,N_10155,N_10599);
xnor U11710 (N_11710,N_10670,N_9903);
nand U11711 (N_11711,N_10606,N_10117);
nand U11712 (N_11712,N_10569,N_10085);
xnor U11713 (N_11713,N_9814,N_10312);
nor U11714 (N_11714,N_10501,N_10306);
nor U11715 (N_11715,N_10086,N_10205);
xnor U11716 (N_11716,N_10098,N_9973);
and U11717 (N_11717,N_9625,N_10419);
nand U11718 (N_11718,N_10514,N_10348);
or U11719 (N_11719,N_10526,N_9631);
or U11720 (N_11720,N_10371,N_10472);
and U11721 (N_11721,N_10564,N_10546);
nand U11722 (N_11722,N_10675,N_10236);
or U11723 (N_11723,N_9896,N_9602);
and U11724 (N_11724,N_10790,N_10284);
and U11725 (N_11725,N_10629,N_10376);
xnor U11726 (N_11726,N_10617,N_10019);
xor U11727 (N_11727,N_9827,N_10247);
nor U11728 (N_11728,N_10148,N_10456);
nand U11729 (N_11729,N_10184,N_10009);
and U11730 (N_11730,N_10607,N_10465);
nand U11731 (N_11731,N_10554,N_10510);
and U11732 (N_11732,N_10529,N_10338);
nand U11733 (N_11733,N_10529,N_10394);
nand U11734 (N_11734,N_10443,N_10779);
and U11735 (N_11735,N_9989,N_10279);
and U11736 (N_11736,N_10136,N_9909);
xor U11737 (N_11737,N_10734,N_9752);
nand U11738 (N_11738,N_9734,N_9684);
or U11739 (N_11739,N_10161,N_10180);
nor U11740 (N_11740,N_10399,N_10762);
nand U11741 (N_11741,N_9812,N_10305);
xor U11742 (N_11742,N_9873,N_9705);
nor U11743 (N_11743,N_9621,N_10108);
xor U11744 (N_11744,N_10694,N_10149);
nand U11745 (N_11745,N_10772,N_10161);
nor U11746 (N_11746,N_10323,N_9774);
nor U11747 (N_11747,N_9819,N_9912);
or U11748 (N_11748,N_10132,N_10246);
nor U11749 (N_11749,N_10363,N_9611);
xor U11750 (N_11750,N_10308,N_10765);
nand U11751 (N_11751,N_10356,N_10418);
nor U11752 (N_11752,N_10613,N_10516);
nor U11753 (N_11753,N_10032,N_10745);
nor U11754 (N_11754,N_10196,N_10752);
nand U11755 (N_11755,N_10176,N_9873);
and U11756 (N_11756,N_10028,N_10100);
or U11757 (N_11757,N_9671,N_9883);
nand U11758 (N_11758,N_10410,N_9644);
nor U11759 (N_11759,N_10771,N_9991);
xnor U11760 (N_11760,N_10763,N_10117);
xnor U11761 (N_11761,N_9694,N_9675);
or U11762 (N_11762,N_9665,N_10722);
or U11763 (N_11763,N_10079,N_9895);
nand U11764 (N_11764,N_9954,N_10774);
and U11765 (N_11765,N_10136,N_10254);
xor U11766 (N_11766,N_10445,N_10565);
xor U11767 (N_11767,N_9817,N_10420);
and U11768 (N_11768,N_9659,N_9736);
and U11769 (N_11769,N_10206,N_10181);
or U11770 (N_11770,N_10044,N_10549);
or U11771 (N_11771,N_10165,N_9924);
nor U11772 (N_11772,N_10177,N_10199);
nand U11773 (N_11773,N_10268,N_9631);
and U11774 (N_11774,N_10460,N_10604);
or U11775 (N_11775,N_10537,N_9966);
xnor U11776 (N_11776,N_9842,N_10213);
xor U11777 (N_11777,N_9880,N_10639);
xnor U11778 (N_11778,N_9727,N_9816);
nand U11779 (N_11779,N_10280,N_10647);
nand U11780 (N_11780,N_9675,N_10268);
or U11781 (N_11781,N_10576,N_10056);
xor U11782 (N_11782,N_10642,N_10238);
and U11783 (N_11783,N_10781,N_9875);
or U11784 (N_11784,N_10428,N_9871);
nor U11785 (N_11785,N_10054,N_10387);
nor U11786 (N_11786,N_9740,N_10556);
or U11787 (N_11787,N_10011,N_10095);
xor U11788 (N_11788,N_9865,N_9926);
and U11789 (N_11789,N_10345,N_10560);
nand U11790 (N_11790,N_9915,N_9907);
xnor U11791 (N_11791,N_10413,N_9770);
nand U11792 (N_11792,N_10546,N_10649);
and U11793 (N_11793,N_9952,N_10558);
nor U11794 (N_11794,N_10617,N_9683);
nor U11795 (N_11795,N_10623,N_9656);
nand U11796 (N_11796,N_9842,N_10728);
or U11797 (N_11797,N_9723,N_10491);
nor U11798 (N_11798,N_9789,N_10783);
and U11799 (N_11799,N_10487,N_10390);
xnor U11800 (N_11800,N_9858,N_9853);
nand U11801 (N_11801,N_10126,N_10693);
nand U11802 (N_11802,N_10225,N_10428);
or U11803 (N_11803,N_9782,N_10730);
xnor U11804 (N_11804,N_10457,N_10070);
or U11805 (N_11805,N_9965,N_10309);
or U11806 (N_11806,N_9728,N_10421);
and U11807 (N_11807,N_10794,N_10478);
and U11808 (N_11808,N_10767,N_10261);
nor U11809 (N_11809,N_10593,N_10358);
nor U11810 (N_11810,N_10279,N_10623);
xnor U11811 (N_11811,N_10712,N_10024);
xor U11812 (N_11812,N_10458,N_9752);
nor U11813 (N_11813,N_10201,N_10374);
xor U11814 (N_11814,N_10127,N_10029);
nor U11815 (N_11815,N_9676,N_9922);
or U11816 (N_11816,N_10416,N_10492);
xor U11817 (N_11817,N_10596,N_10565);
xor U11818 (N_11818,N_10258,N_10660);
or U11819 (N_11819,N_10473,N_10262);
or U11820 (N_11820,N_10775,N_10267);
and U11821 (N_11821,N_10712,N_10019);
xnor U11822 (N_11822,N_10083,N_10453);
nor U11823 (N_11823,N_10042,N_10436);
or U11824 (N_11824,N_10536,N_10724);
nor U11825 (N_11825,N_9876,N_10010);
or U11826 (N_11826,N_10347,N_9767);
or U11827 (N_11827,N_10605,N_10199);
nor U11828 (N_11828,N_9751,N_10687);
nor U11829 (N_11829,N_9872,N_9808);
xor U11830 (N_11830,N_10004,N_10127);
and U11831 (N_11831,N_9881,N_10548);
nand U11832 (N_11832,N_10034,N_10446);
xor U11833 (N_11833,N_10493,N_10364);
nand U11834 (N_11834,N_9903,N_10115);
nand U11835 (N_11835,N_10163,N_10480);
xnor U11836 (N_11836,N_9804,N_10507);
and U11837 (N_11837,N_10458,N_9836);
xor U11838 (N_11838,N_9767,N_9823);
xnor U11839 (N_11839,N_10469,N_10072);
and U11840 (N_11840,N_9776,N_10718);
nor U11841 (N_11841,N_10260,N_10337);
xor U11842 (N_11842,N_9639,N_10543);
or U11843 (N_11843,N_10419,N_9825);
nor U11844 (N_11844,N_9751,N_10675);
xnor U11845 (N_11845,N_10748,N_9795);
xnor U11846 (N_11846,N_10304,N_10518);
or U11847 (N_11847,N_10530,N_9694);
xnor U11848 (N_11848,N_9975,N_10393);
and U11849 (N_11849,N_9781,N_10073);
or U11850 (N_11850,N_9619,N_10117);
or U11851 (N_11851,N_9643,N_10261);
nand U11852 (N_11852,N_10323,N_10346);
and U11853 (N_11853,N_10186,N_10452);
or U11854 (N_11854,N_9878,N_10321);
nor U11855 (N_11855,N_10562,N_10264);
nor U11856 (N_11856,N_9939,N_10539);
nor U11857 (N_11857,N_10514,N_9645);
nor U11858 (N_11858,N_9792,N_10154);
nor U11859 (N_11859,N_10691,N_10334);
and U11860 (N_11860,N_10678,N_9940);
nand U11861 (N_11861,N_9904,N_10742);
or U11862 (N_11862,N_9679,N_9755);
nand U11863 (N_11863,N_10203,N_9641);
and U11864 (N_11864,N_10521,N_10610);
or U11865 (N_11865,N_10442,N_10702);
nor U11866 (N_11866,N_9921,N_10095);
nor U11867 (N_11867,N_9604,N_10263);
nor U11868 (N_11868,N_9673,N_10074);
and U11869 (N_11869,N_10004,N_9964);
nor U11870 (N_11870,N_10626,N_10431);
xnor U11871 (N_11871,N_10796,N_10173);
and U11872 (N_11872,N_10738,N_10015);
or U11873 (N_11873,N_10525,N_10159);
and U11874 (N_11874,N_10145,N_10008);
nor U11875 (N_11875,N_10736,N_10557);
nor U11876 (N_11876,N_10755,N_10001);
nand U11877 (N_11877,N_10226,N_9799);
or U11878 (N_11878,N_9720,N_10579);
nand U11879 (N_11879,N_9746,N_10563);
xnor U11880 (N_11880,N_10665,N_10653);
nand U11881 (N_11881,N_9804,N_10333);
or U11882 (N_11882,N_9663,N_9902);
nor U11883 (N_11883,N_10381,N_10176);
nor U11884 (N_11884,N_10520,N_10434);
nor U11885 (N_11885,N_10258,N_10295);
nand U11886 (N_11886,N_10128,N_9984);
nor U11887 (N_11887,N_10693,N_10141);
xnor U11888 (N_11888,N_10791,N_10749);
nor U11889 (N_11889,N_10110,N_9974);
or U11890 (N_11890,N_10599,N_10487);
nor U11891 (N_11891,N_10136,N_10587);
nand U11892 (N_11892,N_10406,N_10114);
xnor U11893 (N_11893,N_10578,N_9690);
nand U11894 (N_11894,N_10743,N_9674);
nor U11895 (N_11895,N_9703,N_10158);
or U11896 (N_11896,N_10305,N_10324);
nor U11897 (N_11897,N_10254,N_10194);
nand U11898 (N_11898,N_10681,N_9944);
xor U11899 (N_11899,N_10494,N_10525);
nor U11900 (N_11900,N_10102,N_10288);
xor U11901 (N_11901,N_10546,N_9983);
and U11902 (N_11902,N_10054,N_10661);
and U11903 (N_11903,N_10250,N_10732);
nand U11904 (N_11904,N_10157,N_9778);
nor U11905 (N_11905,N_10189,N_9939);
or U11906 (N_11906,N_10468,N_9684);
nor U11907 (N_11907,N_10102,N_9748);
and U11908 (N_11908,N_10634,N_10205);
xor U11909 (N_11909,N_10770,N_10402);
nand U11910 (N_11910,N_10479,N_10336);
nand U11911 (N_11911,N_10212,N_10757);
nor U11912 (N_11912,N_10020,N_10787);
and U11913 (N_11913,N_10763,N_9864);
and U11914 (N_11914,N_10361,N_10520);
xor U11915 (N_11915,N_10781,N_10545);
nor U11916 (N_11916,N_10453,N_10107);
or U11917 (N_11917,N_9717,N_10414);
nand U11918 (N_11918,N_9636,N_9798);
xnor U11919 (N_11919,N_9692,N_10565);
or U11920 (N_11920,N_9969,N_10097);
or U11921 (N_11921,N_10593,N_10013);
xnor U11922 (N_11922,N_10466,N_9988);
or U11923 (N_11923,N_10773,N_10353);
xnor U11924 (N_11924,N_9923,N_9928);
nor U11925 (N_11925,N_10154,N_10556);
or U11926 (N_11926,N_9783,N_9925);
xnor U11927 (N_11927,N_10252,N_10675);
nor U11928 (N_11928,N_10719,N_9648);
nor U11929 (N_11929,N_10737,N_10021);
xnor U11930 (N_11930,N_9841,N_10697);
and U11931 (N_11931,N_10168,N_9670);
and U11932 (N_11932,N_10196,N_9865);
nor U11933 (N_11933,N_10305,N_10303);
nor U11934 (N_11934,N_10762,N_9901);
nor U11935 (N_11935,N_9623,N_9822);
nand U11936 (N_11936,N_10068,N_10415);
nor U11937 (N_11937,N_10441,N_10427);
and U11938 (N_11938,N_9934,N_10508);
and U11939 (N_11939,N_10606,N_10321);
or U11940 (N_11940,N_10428,N_10029);
nand U11941 (N_11941,N_10334,N_9814);
and U11942 (N_11942,N_10729,N_10650);
nor U11943 (N_11943,N_9673,N_10694);
nor U11944 (N_11944,N_10716,N_10367);
nor U11945 (N_11945,N_9965,N_10424);
xnor U11946 (N_11946,N_10562,N_10149);
nand U11947 (N_11947,N_9816,N_10694);
xnor U11948 (N_11948,N_10560,N_10734);
xnor U11949 (N_11949,N_10625,N_9703);
nand U11950 (N_11950,N_10051,N_10431);
or U11951 (N_11951,N_9977,N_10483);
nand U11952 (N_11952,N_10356,N_10467);
or U11953 (N_11953,N_10598,N_10716);
nand U11954 (N_11954,N_10462,N_9865);
nand U11955 (N_11955,N_10463,N_10014);
or U11956 (N_11956,N_9838,N_10335);
and U11957 (N_11957,N_10024,N_9978);
xor U11958 (N_11958,N_9946,N_10209);
xnor U11959 (N_11959,N_10081,N_10158);
or U11960 (N_11960,N_9636,N_9793);
or U11961 (N_11961,N_9804,N_10348);
and U11962 (N_11962,N_9961,N_10693);
nand U11963 (N_11963,N_10452,N_10216);
xnor U11964 (N_11964,N_10145,N_10291);
xnor U11965 (N_11965,N_10378,N_10446);
nor U11966 (N_11966,N_10273,N_9830);
and U11967 (N_11967,N_10051,N_9638);
xor U11968 (N_11968,N_10478,N_10258);
and U11969 (N_11969,N_10524,N_10319);
xnor U11970 (N_11970,N_10080,N_10709);
xor U11971 (N_11971,N_10296,N_10050);
nand U11972 (N_11972,N_10622,N_10755);
nor U11973 (N_11973,N_10681,N_10635);
xor U11974 (N_11974,N_9924,N_10764);
or U11975 (N_11975,N_9928,N_10101);
nand U11976 (N_11976,N_10725,N_10252);
or U11977 (N_11977,N_10046,N_10581);
nor U11978 (N_11978,N_10105,N_10638);
xor U11979 (N_11979,N_9772,N_10646);
or U11980 (N_11980,N_10373,N_10238);
or U11981 (N_11981,N_10012,N_10548);
xor U11982 (N_11982,N_10417,N_10445);
nand U11983 (N_11983,N_9997,N_10738);
xnor U11984 (N_11984,N_10758,N_9614);
xnor U11985 (N_11985,N_10209,N_10293);
nand U11986 (N_11986,N_9851,N_10374);
and U11987 (N_11987,N_10260,N_10552);
and U11988 (N_11988,N_9706,N_9606);
or U11989 (N_11989,N_10335,N_10000);
and U11990 (N_11990,N_10050,N_10073);
or U11991 (N_11991,N_9766,N_9626);
and U11992 (N_11992,N_10333,N_10177);
or U11993 (N_11993,N_10015,N_10467);
nor U11994 (N_11994,N_10601,N_10075);
nand U11995 (N_11995,N_10000,N_9699);
and U11996 (N_11996,N_9963,N_10045);
xor U11997 (N_11997,N_10536,N_10500);
and U11998 (N_11998,N_10682,N_10756);
or U11999 (N_11999,N_10125,N_10719);
xor U12000 (N_12000,N_10817,N_11205);
and U12001 (N_12001,N_11839,N_11798);
xor U12002 (N_12002,N_11570,N_11632);
nand U12003 (N_12003,N_10918,N_10962);
or U12004 (N_12004,N_11065,N_11012);
and U12005 (N_12005,N_10982,N_11173);
or U12006 (N_12006,N_11085,N_10986);
nand U12007 (N_12007,N_11329,N_11309);
and U12008 (N_12008,N_11738,N_10909);
and U12009 (N_12009,N_11735,N_10979);
and U12010 (N_12010,N_10854,N_11061);
or U12011 (N_12011,N_11700,N_11635);
nand U12012 (N_12012,N_10885,N_11862);
nand U12013 (N_12013,N_11097,N_11230);
nor U12014 (N_12014,N_11807,N_11281);
nor U12015 (N_12015,N_11927,N_11656);
xor U12016 (N_12016,N_11528,N_11702);
or U12017 (N_12017,N_11695,N_11156);
and U12018 (N_12018,N_11289,N_11530);
xnor U12019 (N_12019,N_11201,N_11945);
nor U12020 (N_12020,N_11286,N_11578);
and U12021 (N_12021,N_11521,N_10893);
xor U12022 (N_12022,N_11339,N_11613);
nand U12023 (N_12023,N_11092,N_11791);
xnor U12024 (N_12024,N_11179,N_11002);
xor U12025 (N_12025,N_11623,N_11463);
nor U12026 (N_12026,N_11744,N_11140);
xnor U12027 (N_12027,N_11482,N_11010);
and U12028 (N_12028,N_11222,N_10999);
nand U12029 (N_12029,N_11626,N_11192);
nor U12030 (N_12030,N_11703,N_11291);
and U12031 (N_12031,N_11874,N_11535);
and U12032 (N_12032,N_11020,N_11911);
or U12033 (N_12033,N_10911,N_11612);
and U12034 (N_12034,N_11225,N_11048);
and U12035 (N_12035,N_11557,N_11942);
nand U12036 (N_12036,N_11228,N_10894);
or U12037 (N_12037,N_11729,N_11507);
nor U12038 (N_12038,N_11915,N_11479);
or U12039 (N_12039,N_11433,N_11963);
nand U12040 (N_12040,N_11089,N_11494);
nand U12041 (N_12041,N_11549,N_11907);
and U12042 (N_12042,N_11403,N_11891);
and U12043 (N_12043,N_11981,N_11055);
and U12044 (N_12044,N_10801,N_11502);
nand U12045 (N_12045,N_11475,N_11155);
and U12046 (N_12046,N_10876,N_10832);
and U12047 (N_12047,N_11468,N_10877);
xnor U12048 (N_12048,N_10919,N_11847);
or U12049 (N_12049,N_11239,N_11816);
xnor U12050 (N_12050,N_11529,N_10936);
nand U12051 (N_12051,N_11202,N_11860);
nor U12052 (N_12052,N_11288,N_10819);
nor U12053 (N_12053,N_11064,N_11759);
nor U12054 (N_12054,N_10816,N_11653);
nand U12055 (N_12055,N_11313,N_11478);
xnor U12056 (N_12056,N_11982,N_11168);
xor U12057 (N_12057,N_11211,N_11389);
nor U12058 (N_12058,N_11914,N_11689);
nor U12059 (N_12059,N_11636,N_10961);
nand U12060 (N_12060,N_11258,N_11131);
or U12061 (N_12061,N_11721,N_11280);
nor U12062 (N_12062,N_11849,N_11894);
and U12063 (N_12063,N_11762,N_11351);
and U12064 (N_12064,N_10944,N_11216);
and U12065 (N_12065,N_11101,N_11671);
nand U12066 (N_12066,N_11873,N_11818);
or U12067 (N_12067,N_11354,N_11797);
and U12068 (N_12068,N_11279,N_11925);
nor U12069 (N_12069,N_11633,N_10950);
xor U12070 (N_12070,N_11018,N_11769);
and U12071 (N_12071,N_11739,N_11506);
or U12072 (N_12072,N_10866,N_10825);
nand U12073 (N_12073,N_11990,N_10987);
and U12074 (N_12074,N_11728,N_11439);
or U12075 (N_12075,N_11262,N_10855);
nor U12076 (N_12076,N_10957,N_11268);
or U12077 (N_12077,N_11509,N_11863);
nor U12078 (N_12078,N_11464,N_11447);
nor U12079 (N_12079,N_11067,N_11522);
nand U12080 (N_12080,N_11640,N_11926);
xor U12081 (N_12081,N_10803,N_11964);
or U12082 (N_12082,N_11298,N_11774);
nand U12083 (N_12083,N_10867,N_11814);
or U12084 (N_12084,N_11095,N_11986);
nor U12085 (N_12085,N_11074,N_11758);
or U12086 (N_12086,N_11295,N_11954);
nand U12087 (N_12087,N_11181,N_11629);
or U12088 (N_12088,N_10847,N_11081);
nand U12089 (N_12089,N_11670,N_11078);
and U12090 (N_12090,N_10827,N_10949);
nand U12091 (N_12091,N_11121,N_11487);
xor U12092 (N_12092,N_11462,N_11719);
nor U12093 (N_12093,N_11287,N_11978);
nand U12094 (N_12094,N_10996,N_10839);
or U12095 (N_12095,N_11372,N_11550);
and U12096 (N_12096,N_11962,N_11944);
nand U12097 (N_12097,N_11851,N_10973);
nor U12098 (N_12098,N_11691,N_11826);
xor U12099 (N_12099,N_11659,N_11142);
xor U12100 (N_12100,N_11855,N_11501);
or U12101 (N_12101,N_10889,N_11842);
or U12102 (N_12102,N_11822,N_11946);
nor U12103 (N_12103,N_10964,N_11902);
and U12104 (N_12104,N_10835,N_11548);
xor U12105 (N_12105,N_11740,N_10872);
xor U12106 (N_12106,N_11000,N_11705);
nor U12107 (N_12107,N_11932,N_11731);
or U12108 (N_12108,N_11401,N_11254);
nor U12109 (N_12109,N_11238,N_11310);
and U12110 (N_12110,N_11830,N_11340);
xor U12111 (N_12111,N_11157,N_11264);
or U12112 (N_12112,N_10956,N_10887);
xnor U12113 (N_12113,N_11321,N_11330);
nor U12114 (N_12114,N_11765,N_11450);
and U12115 (N_12115,N_11203,N_11100);
xnor U12116 (N_12116,N_11060,N_11772);
nand U12117 (N_12117,N_11315,N_11032);
nand U12118 (N_12118,N_11196,N_11920);
or U12119 (N_12119,N_11404,N_10963);
nand U12120 (N_12120,N_11616,N_11579);
and U12121 (N_12121,N_11465,N_11887);
or U12122 (N_12122,N_11153,N_11525);
nor U12123 (N_12123,N_11805,N_11122);
or U12124 (N_12124,N_11422,N_11424);
or U12125 (N_12125,N_11253,N_10981);
nor U12126 (N_12126,N_11474,N_11793);
nor U12127 (N_12127,N_11107,N_11045);
or U12128 (N_12128,N_10969,N_11518);
or U12129 (N_12129,N_11341,N_11252);
or U12130 (N_12130,N_11250,N_11910);
or U12131 (N_12131,N_11186,N_11743);
nor U12132 (N_12132,N_11593,N_11130);
nor U12133 (N_12133,N_11349,N_11049);
xor U12134 (N_12134,N_11792,N_11106);
and U12135 (N_12135,N_11188,N_11471);
xnor U12136 (N_12136,N_11180,N_11421);
xnor U12137 (N_12137,N_11104,N_11195);
or U12138 (N_12138,N_11893,N_11362);
xnor U12139 (N_12139,N_11413,N_10846);
or U12140 (N_12140,N_10899,N_11678);
nand U12141 (N_12141,N_11650,N_11795);
nand U12142 (N_12142,N_11854,N_11609);
nor U12143 (N_12143,N_11835,N_11714);
nand U12144 (N_12144,N_11485,N_11241);
xor U12145 (N_12145,N_11643,N_11311);
nand U12146 (N_12146,N_10988,N_11878);
nand U12147 (N_12147,N_11226,N_11290);
xnor U12148 (N_12148,N_11392,N_11076);
and U12149 (N_12149,N_11388,N_11922);
nand U12150 (N_12150,N_10841,N_11898);
nor U12151 (N_12151,N_11872,N_11172);
xor U12152 (N_12152,N_11598,N_10915);
nand U12153 (N_12153,N_11754,N_11412);
and U12154 (N_12154,N_10824,N_11583);
and U12155 (N_12155,N_11586,N_11960);
xnor U12156 (N_12156,N_11958,N_11824);
nand U12157 (N_12157,N_11466,N_11094);
nand U12158 (N_12158,N_10888,N_10808);
xor U12159 (N_12159,N_11322,N_11110);
nand U12160 (N_12160,N_11667,N_10994);
nor U12161 (N_12161,N_11112,N_11669);
nand U12162 (N_12162,N_11827,N_11472);
nand U12163 (N_12163,N_11274,N_10972);
xor U12164 (N_12164,N_11602,N_11848);
xnor U12165 (N_12165,N_11256,N_11692);
nor U12166 (N_12166,N_11282,N_11105);
nor U12167 (N_12167,N_11346,N_11856);
or U12168 (N_12168,N_11199,N_11400);
nor U12169 (N_12169,N_11933,N_10880);
or U12170 (N_12170,N_10844,N_11957);
nor U12171 (N_12171,N_10930,N_11713);
nor U12172 (N_12172,N_11897,N_11711);
nand U12173 (N_12173,N_10946,N_11565);
or U12174 (N_12174,N_11760,N_11516);
nor U12175 (N_12175,N_11257,N_10992);
nor U12176 (N_12176,N_11859,N_11971);
xnor U12177 (N_12177,N_11611,N_11581);
nand U12178 (N_12178,N_11117,N_11661);
nand U12179 (N_12179,N_11005,N_11888);
nor U12180 (N_12180,N_11935,N_11972);
nor U12181 (N_12181,N_11788,N_11995);
xnor U12182 (N_12182,N_10904,N_11832);
nor U12183 (N_12183,N_11352,N_11884);
or U12184 (N_12184,N_11207,N_10948);
nand U12185 (N_12185,N_11852,N_11358);
nor U12186 (N_12186,N_11395,N_11141);
or U12187 (N_12187,N_11327,N_11177);
xor U12188 (N_12188,N_11396,N_11234);
nand U12189 (N_12189,N_11476,N_11276);
nor U12190 (N_12190,N_11846,N_11685);
xnor U12191 (N_12191,N_11139,N_10882);
nand U12192 (N_12192,N_11994,N_11764);
or U12193 (N_12193,N_11086,N_11751);
nand U12194 (N_12194,N_11336,N_11663);
xnor U12195 (N_12195,N_11335,N_11390);
nand U12196 (N_12196,N_10890,N_11135);
nand U12197 (N_12197,N_11200,N_11036);
nand U12198 (N_12198,N_11297,N_11134);
nand U12199 (N_12199,N_11555,N_11046);
or U12200 (N_12200,N_11183,N_10997);
nor U12201 (N_12201,N_11011,N_11526);
nand U12202 (N_12202,N_10978,N_11497);
nand U12203 (N_12203,N_11090,N_10945);
and U12204 (N_12204,N_10960,N_11265);
or U12205 (N_12205,N_11240,N_11642);
and U12206 (N_12206,N_11552,N_11580);
and U12207 (N_12207,N_11664,N_11999);
and U12208 (N_12208,N_11899,N_11331);
nor U12209 (N_12209,N_11053,N_11275);
nor U12210 (N_12210,N_10947,N_11369);
xnor U12211 (N_12211,N_11918,N_11930);
and U12212 (N_12212,N_11406,N_11576);
xnor U12213 (N_12213,N_11959,N_11837);
and U12214 (N_12214,N_10881,N_11292);
nand U12215 (N_12215,N_11178,N_11371);
or U12216 (N_12216,N_11263,N_11486);
xor U12217 (N_12217,N_11684,N_11283);
xnor U12218 (N_12218,N_11495,N_10943);
and U12219 (N_12219,N_11014,N_11686);
nand U12220 (N_12220,N_11499,N_11532);
xnor U12221 (N_12221,N_10951,N_11072);
nand U12222 (N_12222,N_10912,N_11801);
and U12223 (N_12223,N_11906,N_11704);
and U12224 (N_12224,N_11022,N_11970);
xor U12225 (N_12225,N_11301,N_11488);
nor U12226 (N_12226,N_11353,N_11991);
and U12227 (N_12227,N_11198,N_11145);
and U12228 (N_12228,N_10884,N_11035);
and U12229 (N_12229,N_11120,N_11490);
nor U12230 (N_12230,N_11190,N_11344);
nand U12231 (N_12231,N_11024,N_11755);
xor U12232 (N_12232,N_11879,N_11523);
or U12233 (N_12233,N_11128,N_11547);
and U12234 (N_12234,N_11710,N_10814);
xnor U12235 (N_12235,N_11334,N_11019);
nand U12236 (N_12236,N_11473,N_11766);
or U12237 (N_12237,N_11118,N_11505);
or U12238 (N_12238,N_11706,N_11680);
or U12239 (N_12239,N_11984,N_11615);
nor U12240 (N_12240,N_10968,N_10834);
xnor U12241 (N_12241,N_11378,N_10897);
and U12242 (N_12242,N_10896,N_11567);
xnor U12243 (N_12243,N_11730,N_11594);
or U12244 (N_12244,N_10848,N_10939);
xnor U12245 (N_12245,N_11763,N_11170);
or U12246 (N_12246,N_11870,N_11858);
nand U12247 (N_12247,N_11087,N_11592);
nor U12248 (N_12248,N_11232,N_11052);
or U12249 (N_12249,N_11538,N_11149);
and U12250 (N_12250,N_11073,N_11937);
xor U12251 (N_12251,N_10829,N_11127);
and U12252 (N_12252,N_11489,N_10934);
or U12253 (N_12253,N_10802,N_11307);
nand U12254 (N_12254,N_11437,N_10811);
xnor U12255 (N_12255,N_11812,N_11260);
nor U12256 (N_12256,N_11273,N_10923);
nor U12257 (N_12257,N_11709,N_11044);
or U12258 (N_12258,N_11708,N_11056);
nand U12259 (N_12259,N_11248,N_11182);
or U12260 (N_12260,N_10985,N_11551);
nand U12261 (N_12261,N_10998,N_11359);
xnor U12262 (N_12262,N_11681,N_11624);
xnor U12263 (N_12263,N_10843,N_10932);
or U12264 (N_12264,N_11102,N_11975);
xor U12265 (N_12265,N_11320,N_11811);
nor U12266 (N_12266,N_11144,N_11197);
and U12267 (N_12267,N_11569,N_11455);
xor U12268 (N_12268,N_11741,N_11451);
and U12269 (N_12269,N_11540,N_11590);
and U12270 (N_12270,N_11745,N_11833);
or U12271 (N_12271,N_11316,N_11861);
and U12272 (N_12272,N_11163,N_11088);
xor U12273 (N_12273,N_11857,N_11458);
or U12274 (N_12274,N_11943,N_11806);
nor U12275 (N_12275,N_11690,N_11249);
or U12276 (N_12276,N_11750,N_11165);
nor U12277 (N_12277,N_11566,N_11637);
xor U12278 (N_12278,N_11457,N_11208);
nor U12279 (N_12279,N_10955,N_11420);
or U12280 (N_12280,N_10868,N_11278);
xnor U12281 (N_12281,N_11272,N_11491);
nor U12282 (N_12282,N_11589,N_11725);
and U12283 (N_12283,N_11152,N_11875);
or U12284 (N_12284,N_11503,N_11956);
xnor U12285 (N_12285,N_11030,N_11267);
xnor U12286 (N_12286,N_11606,N_10906);
nand U12287 (N_12287,N_11456,N_11251);
xor U12288 (N_12288,N_11054,N_11723);
and U12289 (N_12289,N_10920,N_11058);
nor U12290 (N_12290,N_11368,N_11360);
xnor U12291 (N_12291,N_11379,N_11574);
nand U12292 (N_12292,N_11559,N_11610);
and U12293 (N_12293,N_11210,N_10901);
xor U12294 (N_12294,N_10990,N_10878);
or U12295 (N_12295,N_11980,N_11405);
or U12296 (N_12296,N_11939,N_11817);
or U12297 (N_12297,N_11381,N_11921);
nor U12298 (N_12298,N_11890,N_11974);
xor U12299 (N_12299,N_11338,N_11231);
or U12300 (N_12300,N_11825,N_11634);
xnor U12301 (N_12301,N_11108,N_11093);
or U12302 (N_12302,N_11732,N_11734);
or U12303 (N_12303,N_11912,N_11601);
nand U12304 (N_12304,N_10863,N_11619);
xnor U12305 (N_12305,N_11214,N_11533);
nor U12306 (N_12306,N_10870,N_10874);
xnor U12307 (N_12307,N_11293,N_11614);
xor U12308 (N_12308,N_11560,N_11607);
or U12309 (N_12309,N_11161,N_11777);
and U12310 (N_12310,N_11077,N_11259);
nand U12311 (N_12311,N_11082,N_11736);
xor U12312 (N_12312,N_11021,N_11057);
nor U12313 (N_12313,N_11880,N_11481);
xor U12314 (N_12314,N_11524,N_11843);
or U12315 (N_12315,N_10858,N_10895);
xnor U12316 (N_12316,N_11802,N_11185);
nand U12317 (N_12317,N_11013,N_10871);
xor U12318 (N_12318,N_11508,N_10898);
and U12319 (N_12319,N_11114,N_11917);
or U12320 (N_12320,N_11783,N_11596);
and U12321 (N_12321,N_11840,N_11448);
or U12322 (N_12322,N_11919,N_11786);
nor U12323 (N_12323,N_11784,N_11630);
and U12324 (N_12324,N_11398,N_11790);
or U12325 (N_12325,N_11480,N_11909);
or U12326 (N_12326,N_10818,N_11071);
nand U12327 (N_12327,N_11099,N_10864);
nand U12328 (N_12328,N_11936,N_11815);
or U12329 (N_12329,N_11217,N_11164);
nand U12330 (N_12330,N_10931,N_10928);
nor U12331 (N_12331,N_11673,N_11444);
xor U12332 (N_12332,N_11724,N_11435);
nand U12333 (N_12333,N_10823,N_11631);
nand U12334 (N_12334,N_11618,N_10975);
xnor U12335 (N_12335,N_11376,N_11031);
nand U12336 (N_12336,N_11041,N_11410);
xnor U12337 (N_12337,N_11427,N_11285);
or U12338 (N_12338,N_11967,N_11720);
or U12339 (N_12339,N_11062,N_10861);
and U12340 (N_12340,N_11781,N_11886);
or U12341 (N_12341,N_10812,N_11761);
nor U12342 (N_12342,N_11417,N_11123);
xnor U12343 (N_12343,N_10857,N_11512);
and U12344 (N_12344,N_11391,N_11885);
and U12345 (N_12345,N_10845,N_11988);
nor U12346 (N_12346,N_11985,N_11561);
nor U12347 (N_12347,N_11799,N_11151);
nor U12348 (N_12348,N_11079,N_11900);
or U12349 (N_12349,N_11699,N_11446);
nor U12350 (N_12350,N_10850,N_11542);
xnor U12351 (N_12351,N_10853,N_11209);
nand U12352 (N_12352,N_11838,N_11477);
or U12353 (N_12353,N_11961,N_11545);
nand U12354 (N_12354,N_11776,N_11775);
nor U12355 (N_12355,N_11075,N_10966);
and U12356 (N_12356,N_11115,N_11672);
nor U12357 (N_12357,N_11780,N_11515);
nor U12358 (N_12358,N_11218,N_11213);
nor U12359 (N_12359,N_11600,N_10892);
xnor U12360 (N_12360,N_11534,N_11955);
nand U12361 (N_12361,N_11716,N_11539);
nand U12362 (N_12362,N_11992,N_11803);
xor U12363 (N_12363,N_10938,N_11302);
or U12364 (N_12364,N_11098,N_11668);
or U12365 (N_12365,N_10828,N_10913);
or U12366 (N_12366,N_11212,N_11025);
nor U12367 (N_12367,N_11496,N_11903);
xnor U12368 (N_12368,N_11050,N_10807);
and U12369 (N_12369,N_11337,N_11393);
nand U12370 (N_12370,N_11430,N_11625);
and U12371 (N_12371,N_11277,N_11756);
nand U12372 (N_12372,N_11562,N_11683);
xor U12373 (N_12373,N_11350,N_11445);
nor U12374 (N_12374,N_11397,N_11950);
and U12375 (N_12375,N_11698,N_10837);
and U12376 (N_12376,N_11931,N_11284);
nor U12377 (N_12377,N_10805,N_11325);
or U12378 (N_12378,N_11148,N_11881);
nand U12379 (N_12379,N_10859,N_11928);
or U12380 (N_12380,N_11343,N_11319);
and U12381 (N_12381,N_11845,N_11658);
and U12382 (N_12382,N_11809,N_11701);
or U12383 (N_12383,N_11271,N_11416);
or U12384 (N_12384,N_11662,N_11864);
and U12385 (N_12385,N_11411,N_10921);
nor U12386 (N_12386,N_11564,N_10971);
or U12387 (N_12387,N_11882,N_11342);
nor U12388 (N_12388,N_11387,N_11184);
xor U12389 (N_12389,N_11219,N_11892);
nor U12390 (N_12390,N_11345,N_11454);
or U12391 (N_12391,N_11648,N_11947);
and U12392 (N_12392,N_11296,N_11554);
nand U12393 (N_12393,N_11652,N_11844);
nand U12394 (N_12394,N_11834,N_10852);
nor U12395 (N_12395,N_11537,N_10935);
nand U12396 (N_12396,N_11655,N_10941);
nand U12397 (N_12397,N_11541,N_11399);
xnor U12398 (N_12398,N_11223,N_11493);
and U12399 (N_12399,N_11007,N_11436);
nand U12400 (N_12400,N_11317,N_11083);
nand U12401 (N_12401,N_10902,N_11103);
nand U12402 (N_12402,N_11419,N_11129);
nand U12403 (N_12403,N_10965,N_11374);
nor U12404 (N_12404,N_11461,N_11154);
and U12405 (N_12405,N_11175,N_11987);
nand U12406 (N_12406,N_11831,N_11674);
nor U12407 (N_12407,N_11753,N_11979);
xnor U12408 (N_12408,N_11431,N_10925);
xor U12409 (N_12409,N_10873,N_11813);
and U12410 (N_12410,N_11008,N_10952);
nor U12411 (N_12411,N_11934,N_11605);
or U12412 (N_12412,N_11965,N_11328);
or U12413 (N_12413,N_11804,N_11040);
nand U12414 (N_12414,N_11865,N_10830);
and U12415 (N_12415,N_11794,N_11176);
or U12416 (N_12416,N_11235,N_11587);
xnor U12417 (N_12417,N_11111,N_11438);
nand U12418 (N_12418,N_11929,N_11722);
nor U12419 (N_12419,N_11641,N_11823);
and U12420 (N_12420,N_11498,N_11408);
or U12421 (N_12421,N_11752,N_11133);
or U12422 (N_12422,N_11385,N_10810);
and U12423 (N_12423,N_11998,N_11429);
nand U12424 (N_12424,N_11042,N_11194);
nor U12425 (N_12425,N_11380,N_11993);
nand U12426 (N_12426,N_10869,N_10886);
or U12427 (N_12427,N_10984,N_11187);
nand U12428 (N_12428,N_11206,N_11733);
xor U12429 (N_12429,N_11159,N_11027);
nor U12430 (N_12430,N_11841,N_11174);
nor U12431 (N_12431,N_11543,N_11137);
and U12432 (N_12432,N_11038,N_11573);
xor U12433 (N_12433,N_11308,N_10860);
or U12434 (N_12434,N_11948,N_10851);
and U12435 (N_12435,N_11414,N_11571);
nor U12436 (N_12436,N_11023,N_11015);
or U12437 (N_12437,N_11323,N_11778);
xnor U12438 (N_12438,N_11952,N_11908);
xor U12439 (N_12439,N_11245,N_11951);
xor U12440 (N_12440,N_11808,N_10954);
xnor U12441 (N_12441,N_11332,N_11976);
xnor U12442 (N_12442,N_11665,N_11246);
and U12443 (N_12443,N_11109,N_11850);
or U12444 (N_12444,N_11363,N_10937);
or U12445 (N_12445,N_11224,N_11717);
or U12446 (N_12446,N_11233,N_11047);
xnor U12447 (N_12447,N_11266,N_10959);
or U12448 (N_12448,N_11453,N_11983);
nor U12449 (N_12449,N_11440,N_11687);
and U12450 (N_12450,N_11584,N_11718);
or U12451 (N_12451,N_10905,N_11070);
xor U12452 (N_12452,N_11582,N_11394);
xnor U12453 (N_12453,N_11572,N_11773);
and U12454 (N_12454,N_11442,N_10926);
nand U12455 (N_12455,N_10813,N_11116);
nor U12456 (N_12456,N_11883,N_11051);
and U12457 (N_12457,N_11407,N_11742);
nand U12458 (N_12458,N_11171,N_11009);
nand U12459 (N_12459,N_11800,N_11871);
xnor U12460 (N_12460,N_11628,N_11204);
or U12461 (N_12461,N_11357,N_11604);
nand U12462 (N_12462,N_11227,N_11588);
and U12463 (N_12463,N_10991,N_11143);
nand U12464 (N_12464,N_11707,N_11449);
nor U12465 (N_12465,N_11876,N_11748);
nor U12466 (N_12466,N_10862,N_11126);
nand U12467 (N_12467,N_11001,N_11869);
xor U12468 (N_12468,N_11091,N_11441);
nand U12469 (N_12469,N_11767,N_11949);
xnor U12470 (N_12470,N_11063,N_11434);
and U12471 (N_12471,N_11160,N_11125);
nand U12472 (N_12472,N_10924,N_10821);
nor U12473 (N_12473,N_11712,N_11383);
xnor U12474 (N_12474,N_10820,N_10865);
nand U12475 (N_12475,N_11715,N_11193);
xnor U12476 (N_12476,N_11029,N_10849);
xor U12477 (N_12477,N_11520,N_11236);
nor U12478 (N_12478,N_10838,N_11492);
or U12479 (N_12479,N_11428,N_11819);
xnor U12480 (N_12480,N_11124,N_11749);
or U12481 (N_12481,N_10842,N_10989);
nand U12482 (N_12482,N_11644,N_10970);
nand U12483 (N_12483,N_11191,N_11654);
nand U12484 (N_12484,N_11096,N_11597);
nor U12485 (N_12485,N_11517,N_11938);
and U12486 (N_12486,N_11941,N_11003);
or U12487 (N_12487,N_11924,N_11037);
or U12488 (N_12488,N_11666,N_11033);
nand U12489 (N_12489,N_11968,N_11132);
or U12490 (N_12490,N_11361,N_11693);
nand U12491 (N_12491,N_11318,N_11237);
nor U12492 (N_12492,N_11645,N_11016);
nand U12493 (N_12493,N_11229,N_11017);
nor U12494 (N_12494,N_11158,N_11510);
and U12495 (N_12495,N_10940,N_11866);
or U12496 (N_12496,N_10836,N_11066);
or U12497 (N_12497,N_11484,N_11796);
nand U12498 (N_12498,N_11366,N_11617);
nand U12499 (N_12499,N_11443,N_11651);
xnor U12500 (N_12500,N_11996,N_11568);
or U12501 (N_12501,N_10833,N_11901);
or U12502 (N_12502,N_10933,N_11621);
nor U12503 (N_12503,N_11829,N_11789);
xnor U12504 (N_12504,N_11536,N_10993);
nand U12505 (N_12505,N_11261,N_11904);
xnor U12506 (N_12506,N_11312,N_11367);
nand U12507 (N_12507,N_11080,N_11746);
xnor U12508 (N_12508,N_11459,N_11306);
or U12509 (N_12509,N_11377,N_11639);
nor U12510 (N_12510,N_10967,N_10804);
or U12511 (N_12511,N_11426,N_11004);
nand U12512 (N_12512,N_11026,N_11084);
or U12513 (N_12513,N_10917,N_11660);
nand U12514 (N_12514,N_10976,N_11244);
and U12515 (N_12515,N_11836,N_11364);
nor U12516 (N_12516,N_11162,N_11304);
nor U12517 (N_12517,N_11460,N_10831);
and U12518 (N_12518,N_10883,N_11136);
or U12519 (N_12519,N_11333,N_11504);
nand U12520 (N_12520,N_11989,N_10929);
nor U12521 (N_12521,N_11622,N_11585);
nor U12522 (N_12522,N_11409,N_11913);
or U12523 (N_12523,N_11638,N_10806);
nand U12524 (N_12524,N_11326,N_11527);
or U12525 (N_12525,N_11696,N_11973);
nor U12526 (N_12526,N_11138,N_11694);
and U12527 (N_12527,N_11563,N_11375);
nand U12528 (N_12528,N_11627,N_11726);
or U12529 (N_12529,N_11782,N_11355);
nor U12530 (N_12530,N_10903,N_11675);
nand U12531 (N_12531,N_11737,N_11119);
nand U12532 (N_12532,N_11365,N_11314);
or U12533 (N_12533,N_11169,N_11531);
xnor U12534 (N_12534,N_11220,N_11415);
nand U12535 (N_12535,N_11500,N_11147);
and U12536 (N_12536,N_11069,N_11513);
nand U12537 (N_12537,N_11347,N_10809);
nand U12538 (N_12538,N_10800,N_11028);
or U12539 (N_12539,N_10907,N_11370);
nor U12540 (N_12540,N_11221,N_11215);
nor U12541 (N_12541,N_11905,N_11467);
nor U12542 (N_12542,N_10910,N_11757);
and U12543 (N_12543,N_11997,N_11146);
and U12544 (N_12544,N_11966,N_11828);
nor U12545 (N_12545,N_11779,N_10856);
nand U12546 (N_12546,N_11514,N_11577);
and U12547 (N_12547,N_10980,N_10840);
and U12548 (N_12548,N_11868,N_10826);
xnor U12549 (N_12549,N_10927,N_10977);
xor U12550 (N_12550,N_11425,N_10900);
xor U12551 (N_12551,N_11150,N_11768);
xor U12552 (N_12552,N_11068,N_11043);
and U12553 (N_12553,N_11657,N_10815);
and U12554 (N_12554,N_11386,N_11771);
or U12555 (N_12555,N_11889,N_11270);
or U12556 (N_12556,N_11682,N_11727);
and U12557 (N_12557,N_11867,N_11599);
xnor U12558 (N_12558,N_11544,N_11247);
nor U12559 (N_12559,N_11916,N_11649);
nor U12560 (N_12560,N_11575,N_11556);
xor U12561 (N_12561,N_11243,N_11603);
xnor U12562 (N_12562,N_11697,N_11373);
or U12563 (N_12563,N_10914,N_10953);
nor U12564 (N_12564,N_11432,N_11469);
and U12565 (N_12565,N_11787,N_11546);
and U12566 (N_12566,N_11620,N_11511);
xnor U12567 (N_12567,N_11269,N_11558);
nand U12568 (N_12568,N_11679,N_10891);
nand U12569 (N_12569,N_11483,N_11189);
nand U12570 (N_12570,N_11770,N_11166);
and U12571 (N_12571,N_11300,N_10942);
nand U12572 (N_12572,N_11006,N_11896);
xor U12573 (N_12573,N_11923,N_11059);
nor U12574 (N_12574,N_11303,N_11113);
nor U12575 (N_12575,N_11877,N_11167);
or U12576 (N_12576,N_11324,N_11940);
nand U12577 (N_12577,N_11688,N_11039);
nand U12578 (N_12578,N_11595,N_11348);
and U12579 (N_12579,N_11299,N_11608);
xor U12580 (N_12580,N_10922,N_10958);
nor U12581 (N_12581,N_11294,N_10875);
nor U12582 (N_12582,N_11821,N_11384);
xnor U12583 (N_12583,N_11853,N_11519);
or U12584 (N_12584,N_11820,N_11676);
or U12585 (N_12585,N_11242,N_10908);
nor U12586 (N_12586,N_11646,N_11470);
or U12587 (N_12587,N_11356,N_11895);
or U12588 (N_12588,N_10995,N_11255);
and U12589 (N_12589,N_11647,N_10822);
or U12590 (N_12590,N_11034,N_10974);
xnor U12591 (N_12591,N_11969,N_11402);
or U12592 (N_12592,N_10983,N_11810);
nor U12593 (N_12593,N_11418,N_10879);
or U12594 (N_12594,N_11305,N_11785);
xnor U12595 (N_12595,N_11677,N_11591);
and U12596 (N_12596,N_11953,N_11553);
and U12597 (N_12597,N_11452,N_10916);
and U12598 (N_12598,N_11382,N_11747);
nand U12599 (N_12599,N_11977,N_11423);
and U12600 (N_12600,N_11718,N_11149);
or U12601 (N_12601,N_11905,N_11836);
and U12602 (N_12602,N_11684,N_11515);
nand U12603 (N_12603,N_10994,N_11109);
and U12604 (N_12604,N_11846,N_11702);
xor U12605 (N_12605,N_11141,N_11242);
nand U12606 (N_12606,N_11745,N_11666);
nand U12607 (N_12607,N_11875,N_11289);
nor U12608 (N_12608,N_10860,N_11511);
or U12609 (N_12609,N_11611,N_11188);
and U12610 (N_12610,N_11146,N_11827);
or U12611 (N_12611,N_11490,N_11212);
or U12612 (N_12612,N_11895,N_10911);
and U12613 (N_12613,N_11567,N_11083);
and U12614 (N_12614,N_11866,N_11630);
xnor U12615 (N_12615,N_11230,N_11462);
xor U12616 (N_12616,N_11649,N_11085);
xnor U12617 (N_12617,N_11115,N_11989);
nor U12618 (N_12618,N_11292,N_11328);
xor U12619 (N_12619,N_11086,N_10979);
and U12620 (N_12620,N_11695,N_10903);
and U12621 (N_12621,N_11922,N_11359);
xnor U12622 (N_12622,N_11328,N_10917);
nand U12623 (N_12623,N_11410,N_11874);
or U12624 (N_12624,N_11485,N_11926);
and U12625 (N_12625,N_11364,N_11861);
or U12626 (N_12626,N_11988,N_11608);
and U12627 (N_12627,N_10989,N_11951);
and U12628 (N_12628,N_11877,N_11487);
and U12629 (N_12629,N_10849,N_11640);
nor U12630 (N_12630,N_11138,N_11364);
nand U12631 (N_12631,N_11232,N_11494);
nor U12632 (N_12632,N_11424,N_11813);
nor U12633 (N_12633,N_11478,N_11955);
xor U12634 (N_12634,N_11678,N_11135);
or U12635 (N_12635,N_11412,N_10875);
or U12636 (N_12636,N_11220,N_11977);
xor U12637 (N_12637,N_10891,N_11021);
nor U12638 (N_12638,N_11694,N_10998);
and U12639 (N_12639,N_11926,N_10867);
nor U12640 (N_12640,N_10969,N_11483);
nand U12641 (N_12641,N_10913,N_11266);
nor U12642 (N_12642,N_11235,N_10812);
xor U12643 (N_12643,N_11368,N_11382);
and U12644 (N_12644,N_11099,N_11590);
nor U12645 (N_12645,N_11470,N_11396);
nand U12646 (N_12646,N_11311,N_11589);
nand U12647 (N_12647,N_11656,N_11365);
or U12648 (N_12648,N_11353,N_11386);
nand U12649 (N_12649,N_11527,N_10931);
nand U12650 (N_12650,N_11558,N_11813);
and U12651 (N_12651,N_10999,N_11074);
nor U12652 (N_12652,N_11614,N_10966);
or U12653 (N_12653,N_11608,N_11252);
and U12654 (N_12654,N_11360,N_10961);
nand U12655 (N_12655,N_11409,N_11931);
or U12656 (N_12656,N_11945,N_10936);
or U12657 (N_12657,N_11231,N_11239);
nand U12658 (N_12658,N_11621,N_11275);
or U12659 (N_12659,N_11608,N_11954);
nand U12660 (N_12660,N_10868,N_11012);
nand U12661 (N_12661,N_11047,N_10878);
and U12662 (N_12662,N_11900,N_11151);
or U12663 (N_12663,N_11131,N_11467);
and U12664 (N_12664,N_10868,N_11524);
nand U12665 (N_12665,N_11463,N_11407);
xnor U12666 (N_12666,N_11814,N_11574);
nor U12667 (N_12667,N_11408,N_11187);
and U12668 (N_12668,N_10912,N_10953);
or U12669 (N_12669,N_10913,N_10939);
nand U12670 (N_12670,N_11724,N_10843);
nand U12671 (N_12671,N_11575,N_11705);
or U12672 (N_12672,N_11679,N_11086);
nor U12673 (N_12673,N_10945,N_11411);
xnor U12674 (N_12674,N_11756,N_11655);
nor U12675 (N_12675,N_11203,N_10846);
nor U12676 (N_12676,N_11649,N_11801);
and U12677 (N_12677,N_11390,N_11639);
or U12678 (N_12678,N_11184,N_11615);
xor U12679 (N_12679,N_11630,N_11206);
and U12680 (N_12680,N_11350,N_10817);
xor U12681 (N_12681,N_11557,N_11127);
nor U12682 (N_12682,N_11567,N_11547);
nand U12683 (N_12683,N_11120,N_11925);
nor U12684 (N_12684,N_10885,N_11379);
and U12685 (N_12685,N_10827,N_11799);
and U12686 (N_12686,N_11321,N_11989);
nor U12687 (N_12687,N_11053,N_11581);
nor U12688 (N_12688,N_10988,N_11192);
or U12689 (N_12689,N_11894,N_10983);
or U12690 (N_12690,N_10943,N_10972);
or U12691 (N_12691,N_11066,N_11341);
or U12692 (N_12692,N_11541,N_11606);
nor U12693 (N_12693,N_11877,N_10888);
and U12694 (N_12694,N_11500,N_11269);
nand U12695 (N_12695,N_11976,N_10851);
xnor U12696 (N_12696,N_11075,N_11501);
or U12697 (N_12697,N_11093,N_11942);
or U12698 (N_12698,N_11457,N_11356);
and U12699 (N_12699,N_11937,N_11479);
and U12700 (N_12700,N_11300,N_10960);
nand U12701 (N_12701,N_11749,N_11968);
or U12702 (N_12702,N_11264,N_11714);
or U12703 (N_12703,N_11376,N_11608);
xor U12704 (N_12704,N_10898,N_11613);
nand U12705 (N_12705,N_11331,N_11475);
or U12706 (N_12706,N_11504,N_11695);
and U12707 (N_12707,N_11848,N_11932);
xor U12708 (N_12708,N_11447,N_11639);
xnor U12709 (N_12709,N_11713,N_11064);
and U12710 (N_12710,N_11124,N_11106);
nand U12711 (N_12711,N_11632,N_11467);
nand U12712 (N_12712,N_11666,N_11822);
nand U12713 (N_12713,N_10844,N_11257);
xnor U12714 (N_12714,N_11529,N_11984);
and U12715 (N_12715,N_11238,N_11072);
xnor U12716 (N_12716,N_11691,N_11172);
or U12717 (N_12717,N_11696,N_11052);
nand U12718 (N_12718,N_11133,N_11565);
xnor U12719 (N_12719,N_10816,N_11165);
or U12720 (N_12720,N_11394,N_10972);
and U12721 (N_12721,N_11609,N_10869);
nor U12722 (N_12722,N_11612,N_11776);
or U12723 (N_12723,N_11832,N_11228);
nor U12724 (N_12724,N_10832,N_11434);
nor U12725 (N_12725,N_11103,N_11264);
and U12726 (N_12726,N_11715,N_11477);
and U12727 (N_12727,N_11477,N_11121);
nor U12728 (N_12728,N_11423,N_11131);
nor U12729 (N_12729,N_11922,N_11097);
nor U12730 (N_12730,N_11600,N_11632);
nor U12731 (N_12731,N_11278,N_11083);
nand U12732 (N_12732,N_10900,N_11080);
or U12733 (N_12733,N_11331,N_11885);
nand U12734 (N_12734,N_11772,N_11043);
or U12735 (N_12735,N_11905,N_11884);
xnor U12736 (N_12736,N_11200,N_11203);
or U12737 (N_12737,N_11505,N_11903);
nor U12738 (N_12738,N_11420,N_11016);
or U12739 (N_12739,N_11717,N_11450);
or U12740 (N_12740,N_11340,N_11333);
and U12741 (N_12741,N_11649,N_11686);
or U12742 (N_12742,N_11330,N_11155);
and U12743 (N_12743,N_11777,N_11369);
nand U12744 (N_12744,N_11530,N_11436);
nand U12745 (N_12745,N_11146,N_11806);
or U12746 (N_12746,N_11017,N_11469);
nor U12747 (N_12747,N_11816,N_10887);
nand U12748 (N_12748,N_11761,N_11586);
or U12749 (N_12749,N_11861,N_11920);
nor U12750 (N_12750,N_11847,N_11606);
xnor U12751 (N_12751,N_11710,N_11523);
nor U12752 (N_12752,N_11740,N_11319);
nand U12753 (N_12753,N_10930,N_10838);
nand U12754 (N_12754,N_11338,N_11426);
nor U12755 (N_12755,N_11342,N_11008);
xor U12756 (N_12756,N_11904,N_11631);
nand U12757 (N_12757,N_10995,N_11899);
and U12758 (N_12758,N_11642,N_11469);
nand U12759 (N_12759,N_11115,N_11742);
or U12760 (N_12760,N_11529,N_11942);
or U12761 (N_12761,N_11301,N_11642);
xor U12762 (N_12762,N_10826,N_10876);
or U12763 (N_12763,N_11281,N_11151);
nand U12764 (N_12764,N_11600,N_10947);
or U12765 (N_12765,N_11873,N_11380);
or U12766 (N_12766,N_11824,N_10813);
xnor U12767 (N_12767,N_11973,N_11998);
and U12768 (N_12768,N_11136,N_11194);
xor U12769 (N_12769,N_11471,N_10875);
and U12770 (N_12770,N_11338,N_11214);
nor U12771 (N_12771,N_10890,N_11087);
nand U12772 (N_12772,N_11197,N_11534);
nand U12773 (N_12773,N_11962,N_10990);
nand U12774 (N_12774,N_11018,N_11585);
xor U12775 (N_12775,N_10813,N_11412);
nand U12776 (N_12776,N_11405,N_11700);
nor U12777 (N_12777,N_11460,N_11391);
xnor U12778 (N_12778,N_11850,N_11173);
xnor U12779 (N_12779,N_11548,N_11797);
or U12780 (N_12780,N_10812,N_11526);
and U12781 (N_12781,N_11012,N_11281);
and U12782 (N_12782,N_10879,N_11780);
xor U12783 (N_12783,N_11005,N_11385);
and U12784 (N_12784,N_11405,N_11494);
or U12785 (N_12785,N_10824,N_11505);
or U12786 (N_12786,N_11142,N_11195);
or U12787 (N_12787,N_10984,N_11242);
or U12788 (N_12788,N_11026,N_10910);
xnor U12789 (N_12789,N_11736,N_11196);
and U12790 (N_12790,N_11670,N_11674);
nand U12791 (N_12791,N_11718,N_11444);
xnor U12792 (N_12792,N_11083,N_11149);
and U12793 (N_12793,N_11521,N_11913);
or U12794 (N_12794,N_11637,N_10816);
or U12795 (N_12795,N_11772,N_11826);
nor U12796 (N_12796,N_11764,N_11925);
or U12797 (N_12797,N_11601,N_11147);
nand U12798 (N_12798,N_11008,N_11041);
nor U12799 (N_12799,N_11415,N_11572);
nand U12800 (N_12800,N_11702,N_11620);
or U12801 (N_12801,N_11702,N_10978);
nand U12802 (N_12802,N_11881,N_11692);
and U12803 (N_12803,N_11370,N_11841);
or U12804 (N_12804,N_10801,N_11707);
nor U12805 (N_12805,N_11610,N_11505);
or U12806 (N_12806,N_10939,N_10823);
nor U12807 (N_12807,N_11939,N_11859);
xnor U12808 (N_12808,N_11121,N_11794);
and U12809 (N_12809,N_11491,N_11734);
nand U12810 (N_12810,N_11723,N_11027);
nor U12811 (N_12811,N_10802,N_11729);
xor U12812 (N_12812,N_11163,N_11390);
and U12813 (N_12813,N_11021,N_11431);
nand U12814 (N_12814,N_10834,N_11679);
nand U12815 (N_12815,N_11253,N_10977);
and U12816 (N_12816,N_11482,N_11739);
xnor U12817 (N_12817,N_11252,N_11978);
or U12818 (N_12818,N_11769,N_11096);
nor U12819 (N_12819,N_11046,N_11226);
nor U12820 (N_12820,N_11222,N_10816);
nand U12821 (N_12821,N_10995,N_10800);
xnor U12822 (N_12822,N_11402,N_11302);
or U12823 (N_12823,N_11292,N_10808);
or U12824 (N_12824,N_11073,N_10940);
nor U12825 (N_12825,N_11661,N_11785);
nor U12826 (N_12826,N_10960,N_11530);
nand U12827 (N_12827,N_10832,N_11637);
nor U12828 (N_12828,N_11512,N_11483);
nand U12829 (N_12829,N_11811,N_11514);
and U12830 (N_12830,N_11026,N_10892);
nand U12831 (N_12831,N_11538,N_11494);
xnor U12832 (N_12832,N_11842,N_11902);
nand U12833 (N_12833,N_11313,N_11527);
or U12834 (N_12834,N_11923,N_10930);
and U12835 (N_12835,N_11291,N_11590);
and U12836 (N_12836,N_11276,N_11847);
nor U12837 (N_12837,N_11447,N_11934);
xor U12838 (N_12838,N_11149,N_11868);
and U12839 (N_12839,N_11833,N_11912);
or U12840 (N_12840,N_11399,N_11533);
or U12841 (N_12841,N_11772,N_10979);
and U12842 (N_12842,N_10942,N_10911);
and U12843 (N_12843,N_10922,N_11023);
or U12844 (N_12844,N_11199,N_11146);
nand U12845 (N_12845,N_11807,N_11202);
and U12846 (N_12846,N_11881,N_11601);
xor U12847 (N_12847,N_10995,N_11902);
or U12848 (N_12848,N_11932,N_11624);
xnor U12849 (N_12849,N_11612,N_11230);
xor U12850 (N_12850,N_11011,N_11269);
nand U12851 (N_12851,N_11226,N_11009);
or U12852 (N_12852,N_10878,N_10946);
nand U12853 (N_12853,N_11481,N_10987);
or U12854 (N_12854,N_10962,N_11751);
and U12855 (N_12855,N_11628,N_11512);
nor U12856 (N_12856,N_10803,N_10901);
nand U12857 (N_12857,N_11527,N_11977);
and U12858 (N_12858,N_10857,N_11567);
xnor U12859 (N_12859,N_11060,N_11026);
xnor U12860 (N_12860,N_11619,N_11055);
or U12861 (N_12861,N_11542,N_11982);
and U12862 (N_12862,N_11110,N_11745);
and U12863 (N_12863,N_10896,N_11242);
nand U12864 (N_12864,N_11871,N_11244);
and U12865 (N_12865,N_11989,N_11776);
xor U12866 (N_12866,N_11190,N_11459);
or U12867 (N_12867,N_11098,N_11538);
and U12868 (N_12868,N_10893,N_11834);
and U12869 (N_12869,N_11303,N_11999);
xor U12870 (N_12870,N_10843,N_11972);
and U12871 (N_12871,N_11145,N_11927);
xnor U12872 (N_12872,N_11419,N_11580);
or U12873 (N_12873,N_11903,N_11283);
and U12874 (N_12874,N_11114,N_11095);
or U12875 (N_12875,N_10937,N_11354);
and U12876 (N_12876,N_11025,N_11573);
or U12877 (N_12877,N_11414,N_11143);
nor U12878 (N_12878,N_11535,N_11480);
xor U12879 (N_12879,N_11038,N_11133);
and U12880 (N_12880,N_11275,N_11473);
xor U12881 (N_12881,N_11228,N_11627);
nand U12882 (N_12882,N_10940,N_11681);
and U12883 (N_12883,N_11864,N_10885);
nor U12884 (N_12884,N_11284,N_11258);
and U12885 (N_12885,N_11888,N_11085);
xor U12886 (N_12886,N_11756,N_11880);
nor U12887 (N_12887,N_11870,N_10819);
nand U12888 (N_12888,N_11369,N_11568);
nand U12889 (N_12889,N_11436,N_11227);
xnor U12890 (N_12890,N_10967,N_11900);
nand U12891 (N_12891,N_11955,N_11589);
xor U12892 (N_12892,N_11620,N_11250);
and U12893 (N_12893,N_10959,N_11643);
nand U12894 (N_12894,N_11617,N_10962);
and U12895 (N_12895,N_11822,N_11466);
or U12896 (N_12896,N_10899,N_11875);
nand U12897 (N_12897,N_11475,N_10894);
or U12898 (N_12898,N_11682,N_11246);
and U12899 (N_12899,N_11332,N_11306);
and U12900 (N_12900,N_11851,N_11590);
nor U12901 (N_12901,N_11184,N_11365);
xor U12902 (N_12902,N_11182,N_11299);
xor U12903 (N_12903,N_10838,N_10885);
xnor U12904 (N_12904,N_11996,N_11691);
and U12905 (N_12905,N_11032,N_11724);
nand U12906 (N_12906,N_11103,N_11313);
nor U12907 (N_12907,N_11610,N_11658);
nand U12908 (N_12908,N_11249,N_11119);
and U12909 (N_12909,N_11267,N_11430);
and U12910 (N_12910,N_11259,N_11164);
xor U12911 (N_12911,N_10980,N_11507);
or U12912 (N_12912,N_11899,N_10978);
and U12913 (N_12913,N_11918,N_10930);
nor U12914 (N_12914,N_11659,N_11211);
and U12915 (N_12915,N_11754,N_11954);
nor U12916 (N_12916,N_10903,N_11129);
and U12917 (N_12917,N_11764,N_11274);
and U12918 (N_12918,N_11130,N_11886);
xor U12919 (N_12919,N_10844,N_11225);
or U12920 (N_12920,N_10875,N_11215);
and U12921 (N_12921,N_11905,N_11952);
xor U12922 (N_12922,N_11068,N_10858);
xor U12923 (N_12923,N_11616,N_11754);
xnor U12924 (N_12924,N_11398,N_10821);
xor U12925 (N_12925,N_11914,N_11091);
or U12926 (N_12926,N_10889,N_11742);
nand U12927 (N_12927,N_11152,N_10979);
or U12928 (N_12928,N_10805,N_11621);
xnor U12929 (N_12929,N_11984,N_11975);
or U12930 (N_12930,N_11459,N_11668);
nand U12931 (N_12931,N_11126,N_11810);
and U12932 (N_12932,N_11494,N_11425);
or U12933 (N_12933,N_11355,N_11429);
xor U12934 (N_12934,N_11062,N_10801);
nand U12935 (N_12935,N_11664,N_10843);
or U12936 (N_12936,N_11982,N_11320);
nand U12937 (N_12937,N_11505,N_11466);
or U12938 (N_12938,N_11591,N_11486);
and U12939 (N_12939,N_11908,N_11427);
or U12940 (N_12940,N_11228,N_11040);
xnor U12941 (N_12941,N_10934,N_11074);
nand U12942 (N_12942,N_11205,N_11307);
xnor U12943 (N_12943,N_11153,N_11469);
xor U12944 (N_12944,N_11977,N_11729);
nand U12945 (N_12945,N_11210,N_11232);
nand U12946 (N_12946,N_11809,N_11686);
xor U12947 (N_12947,N_10881,N_11205);
and U12948 (N_12948,N_11494,N_11074);
nand U12949 (N_12949,N_11031,N_11127);
or U12950 (N_12950,N_11843,N_11342);
nor U12951 (N_12951,N_11215,N_11073);
or U12952 (N_12952,N_11379,N_11154);
xor U12953 (N_12953,N_10827,N_11088);
and U12954 (N_12954,N_11276,N_11230);
nand U12955 (N_12955,N_11587,N_11260);
xnor U12956 (N_12956,N_11119,N_11760);
xor U12957 (N_12957,N_10889,N_11965);
nor U12958 (N_12958,N_11142,N_10850);
or U12959 (N_12959,N_11300,N_11570);
xor U12960 (N_12960,N_10980,N_11135);
or U12961 (N_12961,N_11949,N_11742);
xor U12962 (N_12962,N_11947,N_11346);
or U12963 (N_12963,N_11953,N_11794);
or U12964 (N_12964,N_11647,N_11939);
xnor U12965 (N_12965,N_11484,N_11916);
nor U12966 (N_12966,N_11030,N_11586);
or U12967 (N_12967,N_11594,N_11381);
nand U12968 (N_12968,N_11218,N_11394);
and U12969 (N_12969,N_11171,N_10938);
nand U12970 (N_12970,N_10859,N_11944);
nand U12971 (N_12971,N_10804,N_11132);
nor U12972 (N_12972,N_11500,N_10805);
xor U12973 (N_12973,N_11760,N_11434);
xor U12974 (N_12974,N_11382,N_11398);
or U12975 (N_12975,N_11057,N_11996);
xnor U12976 (N_12976,N_11324,N_10910);
xnor U12977 (N_12977,N_11447,N_11939);
or U12978 (N_12978,N_11453,N_11857);
nand U12979 (N_12979,N_11083,N_10802);
nor U12980 (N_12980,N_10894,N_11126);
and U12981 (N_12981,N_11078,N_10963);
and U12982 (N_12982,N_11689,N_10823);
or U12983 (N_12983,N_11283,N_11094);
nor U12984 (N_12984,N_10856,N_10899);
nand U12985 (N_12985,N_10908,N_11007);
nor U12986 (N_12986,N_11644,N_11180);
and U12987 (N_12987,N_11685,N_11101);
or U12988 (N_12988,N_11518,N_11754);
or U12989 (N_12989,N_11980,N_11829);
xor U12990 (N_12990,N_11362,N_11280);
xnor U12991 (N_12991,N_11830,N_11937);
nand U12992 (N_12992,N_11612,N_11622);
xnor U12993 (N_12993,N_10946,N_11664);
and U12994 (N_12994,N_10885,N_11372);
nand U12995 (N_12995,N_11361,N_10959);
or U12996 (N_12996,N_11296,N_11630);
xor U12997 (N_12997,N_11226,N_11070);
and U12998 (N_12998,N_11562,N_11161);
or U12999 (N_12999,N_10936,N_11266);
nor U13000 (N_13000,N_11034,N_11869);
nand U13001 (N_13001,N_11539,N_11801);
nor U13002 (N_13002,N_11778,N_11185);
xor U13003 (N_13003,N_11464,N_11053);
and U13004 (N_13004,N_11959,N_11554);
or U13005 (N_13005,N_11717,N_11968);
nor U13006 (N_13006,N_11593,N_11076);
or U13007 (N_13007,N_11644,N_11940);
and U13008 (N_13008,N_11402,N_11298);
xnor U13009 (N_13009,N_11233,N_11654);
nand U13010 (N_13010,N_11710,N_11744);
nand U13011 (N_13011,N_11040,N_11503);
nor U13012 (N_13012,N_11276,N_11551);
or U13013 (N_13013,N_11619,N_11277);
xnor U13014 (N_13014,N_11454,N_11412);
and U13015 (N_13015,N_10947,N_11507);
or U13016 (N_13016,N_11091,N_11891);
or U13017 (N_13017,N_11111,N_11675);
nand U13018 (N_13018,N_11485,N_11031);
or U13019 (N_13019,N_11451,N_11593);
nor U13020 (N_13020,N_11306,N_10850);
or U13021 (N_13021,N_11858,N_11682);
nor U13022 (N_13022,N_10809,N_10929);
or U13023 (N_13023,N_11443,N_10982);
nand U13024 (N_13024,N_11504,N_11572);
or U13025 (N_13025,N_11768,N_11166);
nand U13026 (N_13026,N_11671,N_11763);
xnor U13027 (N_13027,N_11430,N_11531);
nand U13028 (N_13028,N_11423,N_11560);
nand U13029 (N_13029,N_10915,N_11520);
xor U13030 (N_13030,N_11354,N_10811);
nand U13031 (N_13031,N_11851,N_11287);
xnor U13032 (N_13032,N_11377,N_11827);
or U13033 (N_13033,N_11298,N_11581);
nand U13034 (N_13034,N_11215,N_11682);
xnor U13035 (N_13035,N_11054,N_11035);
nand U13036 (N_13036,N_11468,N_11733);
and U13037 (N_13037,N_11380,N_11416);
and U13038 (N_13038,N_11992,N_11205);
nor U13039 (N_13039,N_10847,N_11138);
nor U13040 (N_13040,N_11585,N_11260);
and U13041 (N_13041,N_11971,N_11728);
or U13042 (N_13042,N_11534,N_11466);
and U13043 (N_13043,N_11106,N_11759);
nor U13044 (N_13044,N_11249,N_11856);
or U13045 (N_13045,N_11302,N_11370);
nor U13046 (N_13046,N_10992,N_11235);
nor U13047 (N_13047,N_11733,N_11724);
and U13048 (N_13048,N_11209,N_11414);
or U13049 (N_13049,N_11208,N_10856);
nor U13050 (N_13050,N_11422,N_11950);
nor U13051 (N_13051,N_11228,N_11098);
nor U13052 (N_13052,N_11061,N_11411);
and U13053 (N_13053,N_11048,N_11786);
nand U13054 (N_13054,N_10855,N_11347);
xnor U13055 (N_13055,N_11443,N_11623);
nor U13056 (N_13056,N_11793,N_11114);
and U13057 (N_13057,N_11729,N_11662);
nor U13058 (N_13058,N_10899,N_11072);
xnor U13059 (N_13059,N_10909,N_11853);
and U13060 (N_13060,N_11481,N_11472);
nor U13061 (N_13061,N_11916,N_11823);
xor U13062 (N_13062,N_11750,N_11265);
nor U13063 (N_13063,N_11291,N_11034);
and U13064 (N_13064,N_11280,N_10906);
or U13065 (N_13065,N_11635,N_11758);
and U13066 (N_13066,N_11412,N_11595);
or U13067 (N_13067,N_10860,N_11041);
and U13068 (N_13068,N_11239,N_10941);
nand U13069 (N_13069,N_11968,N_11487);
nand U13070 (N_13070,N_11609,N_10963);
xor U13071 (N_13071,N_11245,N_11784);
nand U13072 (N_13072,N_11582,N_11401);
nor U13073 (N_13073,N_11425,N_11364);
nand U13074 (N_13074,N_11591,N_11694);
and U13075 (N_13075,N_10889,N_10908);
xor U13076 (N_13076,N_11510,N_11484);
nand U13077 (N_13077,N_11013,N_11572);
nand U13078 (N_13078,N_10925,N_11837);
nor U13079 (N_13079,N_11801,N_11807);
nor U13080 (N_13080,N_11300,N_11574);
or U13081 (N_13081,N_11486,N_11158);
and U13082 (N_13082,N_11736,N_11257);
and U13083 (N_13083,N_11435,N_11396);
and U13084 (N_13084,N_11537,N_11667);
nand U13085 (N_13085,N_11475,N_11271);
or U13086 (N_13086,N_10904,N_11704);
or U13087 (N_13087,N_11396,N_11099);
nor U13088 (N_13088,N_10949,N_10849);
nor U13089 (N_13089,N_10947,N_11908);
or U13090 (N_13090,N_10963,N_11036);
or U13091 (N_13091,N_11271,N_11317);
and U13092 (N_13092,N_11269,N_11887);
and U13093 (N_13093,N_11420,N_11084);
nand U13094 (N_13094,N_11421,N_11561);
nor U13095 (N_13095,N_11690,N_11146);
nor U13096 (N_13096,N_11771,N_11659);
or U13097 (N_13097,N_11107,N_11659);
xnor U13098 (N_13098,N_11803,N_11198);
or U13099 (N_13099,N_10929,N_11386);
and U13100 (N_13100,N_11068,N_11203);
nand U13101 (N_13101,N_11074,N_11562);
nor U13102 (N_13102,N_11730,N_11436);
and U13103 (N_13103,N_11402,N_11633);
nand U13104 (N_13104,N_11499,N_11141);
and U13105 (N_13105,N_11343,N_11747);
and U13106 (N_13106,N_10928,N_11239);
nor U13107 (N_13107,N_11521,N_10836);
and U13108 (N_13108,N_11443,N_11306);
xnor U13109 (N_13109,N_11771,N_11855);
xnor U13110 (N_13110,N_11358,N_11083);
or U13111 (N_13111,N_10895,N_11606);
xnor U13112 (N_13112,N_10985,N_11983);
nand U13113 (N_13113,N_11258,N_11895);
nor U13114 (N_13114,N_11445,N_11148);
and U13115 (N_13115,N_11085,N_11468);
nand U13116 (N_13116,N_11915,N_10934);
nor U13117 (N_13117,N_10946,N_11838);
nand U13118 (N_13118,N_11006,N_10863);
nand U13119 (N_13119,N_11906,N_11337);
and U13120 (N_13120,N_11883,N_11953);
or U13121 (N_13121,N_11858,N_11894);
xor U13122 (N_13122,N_11827,N_11985);
or U13123 (N_13123,N_11470,N_11267);
xor U13124 (N_13124,N_11673,N_11331);
and U13125 (N_13125,N_10998,N_11027);
nand U13126 (N_13126,N_11413,N_11215);
xnor U13127 (N_13127,N_11217,N_11846);
or U13128 (N_13128,N_10950,N_11290);
and U13129 (N_13129,N_11610,N_11143);
and U13130 (N_13130,N_11510,N_11397);
and U13131 (N_13131,N_11507,N_11692);
nand U13132 (N_13132,N_11223,N_11451);
or U13133 (N_13133,N_11675,N_10954);
nor U13134 (N_13134,N_11883,N_11349);
and U13135 (N_13135,N_11492,N_11070);
or U13136 (N_13136,N_11379,N_11548);
nand U13137 (N_13137,N_10819,N_11740);
xor U13138 (N_13138,N_11706,N_10864);
and U13139 (N_13139,N_11609,N_11669);
nor U13140 (N_13140,N_11627,N_11286);
xor U13141 (N_13141,N_11857,N_11119);
nand U13142 (N_13142,N_11942,N_10962);
xor U13143 (N_13143,N_11750,N_11904);
and U13144 (N_13144,N_11265,N_11365);
and U13145 (N_13145,N_11396,N_11707);
or U13146 (N_13146,N_10955,N_11748);
nor U13147 (N_13147,N_11373,N_11324);
nor U13148 (N_13148,N_11812,N_11317);
and U13149 (N_13149,N_11308,N_11801);
xnor U13150 (N_13150,N_11809,N_11559);
xor U13151 (N_13151,N_10980,N_11396);
nand U13152 (N_13152,N_11013,N_11605);
nor U13153 (N_13153,N_11355,N_11319);
xor U13154 (N_13154,N_11372,N_11159);
xor U13155 (N_13155,N_11595,N_10873);
nor U13156 (N_13156,N_11390,N_11414);
nand U13157 (N_13157,N_11533,N_10824);
nand U13158 (N_13158,N_11033,N_11372);
nand U13159 (N_13159,N_11062,N_11642);
xor U13160 (N_13160,N_10894,N_11021);
and U13161 (N_13161,N_11080,N_11943);
or U13162 (N_13162,N_11105,N_11169);
or U13163 (N_13163,N_11251,N_11295);
nor U13164 (N_13164,N_11036,N_11066);
and U13165 (N_13165,N_10951,N_10934);
nor U13166 (N_13166,N_11646,N_11330);
nor U13167 (N_13167,N_11697,N_11560);
nor U13168 (N_13168,N_11058,N_11083);
and U13169 (N_13169,N_11551,N_11864);
or U13170 (N_13170,N_11586,N_11834);
nor U13171 (N_13171,N_10909,N_11544);
or U13172 (N_13172,N_11992,N_11900);
xnor U13173 (N_13173,N_11172,N_11366);
nor U13174 (N_13174,N_11726,N_11587);
xor U13175 (N_13175,N_11081,N_11925);
and U13176 (N_13176,N_10951,N_10994);
and U13177 (N_13177,N_11994,N_11124);
xor U13178 (N_13178,N_11223,N_11446);
xor U13179 (N_13179,N_10819,N_10999);
or U13180 (N_13180,N_11598,N_11130);
nor U13181 (N_13181,N_11382,N_11816);
xor U13182 (N_13182,N_11146,N_11453);
nor U13183 (N_13183,N_11842,N_11210);
nand U13184 (N_13184,N_11984,N_11212);
nand U13185 (N_13185,N_10816,N_11944);
or U13186 (N_13186,N_10939,N_11223);
nor U13187 (N_13187,N_10807,N_11714);
or U13188 (N_13188,N_10854,N_11099);
nor U13189 (N_13189,N_11312,N_11416);
or U13190 (N_13190,N_11319,N_11203);
or U13191 (N_13191,N_11753,N_11458);
and U13192 (N_13192,N_11328,N_11504);
or U13193 (N_13193,N_11295,N_10840);
nor U13194 (N_13194,N_11066,N_11845);
nor U13195 (N_13195,N_11353,N_11630);
and U13196 (N_13196,N_11192,N_10941);
nand U13197 (N_13197,N_10890,N_11065);
nor U13198 (N_13198,N_11707,N_11905);
xnor U13199 (N_13199,N_11880,N_11427);
nor U13200 (N_13200,N_12572,N_12746);
nand U13201 (N_13201,N_12742,N_12435);
or U13202 (N_13202,N_12040,N_12265);
nor U13203 (N_13203,N_12312,N_12370);
nor U13204 (N_13204,N_12847,N_12466);
xor U13205 (N_13205,N_12509,N_12108);
and U13206 (N_13206,N_12839,N_12257);
and U13207 (N_13207,N_12779,N_12415);
xnor U13208 (N_13208,N_12635,N_12800);
xor U13209 (N_13209,N_12131,N_12998);
nand U13210 (N_13210,N_12246,N_12187);
and U13211 (N_13211,N_12799,N_13174);
nor U13212 (N_13212,N_12678,N_12668);
nor U13213 (N_13213,N_12341,N_13193);
or U13214 (N_13214,N_12879,N_12983);
xor U13215 (N_13215,N_12297,N_12660);
and U13216 (N_13216,N_12756,N_12676);
and U13217 (N_13217,N_13054,N_12959);
nor U13218 (N_13218,N_13027,N_13119);
and U13219 (N_13219,N_12717,N_12145);
nand U13220 (N_13220,N_12400,N_13164);
nand U13221 (N_13221,N_12709,N_12431);
and U13222 (N_13222,N_13026,N_12147);
nand U13223 (N_13223,N_12051,N_12373);
and U13224 (N_13224,N_12149,N_13115);
nor U13225 (N_13225,N_12065,N_13044);
xor U13226 (N_13226,N_12180,N_12865);
xnor U13227 (N_13227,N_12890,N_12785);
nor U13228 (N_13228,N_12278,N_12335);
or U13229 (N_13229,N_12609,N_12809);
nor U13230 (N_13230,N_12037,N_12971);
nand U13231 (N_13231,N_13099,N_12422);
nor U13232 (N_13232,N_12176,N_12646);
or U13233 (N_13233,N_12812,N_12437);
or U13234 (N_13234,N_12551,N_12558);
xor U13235 (N_13235,N_12641,N_12100);
xor U13236 (N_13236,N_12980,N_12221);
nor U13237 (N_13237,N_12266,N_12114);
nand U13238 (N_13238,N_12392,N_12083);
nor U13239 (N_13239,N_12141,N_12394);
nor U13240 (N_13240,N_12116,N_12078);
nand U13241 (N_13241,N_12489,N_12156);
xnor U13242 (N_13242,N_12136,N_12308);
xnor U13243 (N_13243,N_12757,N_12857);
nand U13244 (N_13244,N_12640,N_12880);
nand U13245 (N_13245,N_13101,N_12218);
and U13246 (N_13246,N_13151,N_12854);
and U13247 (N_13247,N_12738,N_12500);
nand U13248 (N_13248,N_12690,N_12896);
or U13249 (N_13249,N_12902,N_12367);
and U13250 (N_13250,N_12719,N_12817);
nor U13251 (N_13251,N_12984,N_13097);
or U13252 (N_13252,N_12580,N_13182);
and U13253 (N_13253,N_12560,N_12087);
xor U13254 (N_13254,N_13178,N_12397);
nand U13255 (N_13255,N_12371,N_12516);
or U13256 (N_13256,N_13091,N_13198);
nand U13257 (N_13257,N_12689,N_13137);
xnor U13258 (N_13258,N_13006,N_12905);
xor U13259 (N_13259,N_12698,N_13087);
xnor U13260 (N_13260,N_12291,N_12128);
xnor U13261 (N_13261,N_12028,N_12589);
nor U13262 (N_13262,N_12199,N_12900);
or U13263 (N_13263,N_12164,N_12916);
nand U13264 (N_13264,N_12462,N_12425);
nand U13265 (N_13265,N_12189,N_12579);
and U13266 (N_13266,N_12869,N_12304);
nor U13267 (N_13267,N_12254,N_12039);
nor U13268 (N_13268,N_13180,N_12811);
nand U13269 (N_13269,N_12731,N_12192);
nor U13270 (N_13270,N_12781,N_12084);
nand U13271 (N_13271,N_12021,N_12845);
nand U13272 (N_13272,N_12741,N_12810);
nor U13273 (N_13273,N_12674,N_13047);
nor U13274 (N_13274,N_12612,N_13060);
xor U13275 (N_13275,N_12115,N_13138);
and U13276 (N_13276,N_12521,N_12333);
xnor U13277 (N_13277,N_12904,N_12915);
nand U13278 (N_13278,N_12836,N_12636);
xor U13279 (N_13279,N_12884,N_12958);
nand U13280 (N_13280,N_12262,N_12823);
and U13281 (N_13281,N_13077,N_12244);
nor U13282 (N_13282,N_12448,N_12961);
nor U13283 (N_13283,N_12020,N_12225);
or U13284 (N_13284,N_12602,N_12043);
or U13285 (N_13285,N_12673,N_12577);
xnor U13286 (N_13286,N_12606,N_13104);
and U13287 (N_13287,N_12728,N_12939);
or U13288 (N_13288,N_12542,N_13168);
and U13289 (N_13289,N_13022,N_12960);
nand U13290 (N_13290,N_12929,N_12699);
or U13291 (N_13291,N_13059,N_13035);
xnor U13292 (N_13292,N_12788,N_12228);
and U13293 (N_13293,N_12859,N_12918);
xnor U13294 (N_13294,N_12449,N_12909);
nor U13295 (N_13295,N_12541,N_12351);
and U13296 (N_13296,N_12970,N_12684);
nand U13297 (N_13297,N_12707,N_12376);
or U13298 (N_13298,N_12289,N_12471);
xnor U13299 (N_13299,N_12356,N_12185);
and U13300 (N_13300,N_12016,N_12398);
or U13301 (N_13301,N_12352,N_12484);
nand U13302 (N_13302,N_13149,N_13126);
or U13303 (N_13303,N_12193,N_12544);
nand U13304 (N_13304,N_13124,N_13105);
xor U13305 (N_13305,N_12241,N_12585);
xnor U13306 (N_13306,N_12327,N_13071);
xor U13307 (N_13307,N_12005,N_13025);
or U13308 (N_13308,N_12822,N_12801);
nand U13309 (N_13309,N_13037,N_12184);
and U13310 (N_13310,N_12331,N_12480);
nor U13311 (N_13311,N_12769,N_12790);
and U13312 (N_13312,N_13122,N_12569);
nand U13313 (N_13313,N_12436,N_13024);
nor U13314 (N_13314,N_12364,N_12336);
and U13315 (N_13315,N_12679,N_12619);
nor U13316 (N_13316,N_12599,N_12760);
or U13317 (N_13317,N_12063,N_12414);
nor U13318 (N_13318,N_12628,N_12104);
nand U13319 (N_13319,N_12532,N_12566);
nand U13320 (N_13320,N_12837,N_13075);
xnor U13321 (N_13321,N_12486,N_12103);
nor U13322 (N_13322,N_12598,N_12253);
or U13323 (N_13323,N_12345,N_12791);
or U13324 (N_13324,N_12066,N_12841);
and U13325 (N_13325,N_12794,N_12217);
nand U13326 (N_13326,N_13147,N_12643);
and U13327 (N_13327,N_12299,N_12664);
and U13328 (N_13328,N_12657,N_12263);
nand U13329 (N_13329,N_12219,N_12157);
or U13330 (N_13330,N_12440,N_12206);
or U13331 (N_13331,N_12752,N_13053);
and U13332 (N_13332,N_12624,N_12320);
nor U13333 (N_13333,N_12615,N_13034);
and U13334 (N_13334,N_12031,N_12284);
nand U13335 (N_13335,N_13146,N_13056);
nor U13336 (N_13336,N_12999,N_12277);
nand U13337 (N_13337,N_12737,N_12595);
nor U13338 (N_13338,N_12740,N_12618);
nor U13339 (N_13339,N_12829,N_12910);
or U13340 (N_13340,N_12766,N_12018);
nand U13341 (N_13341,N_12026,N_12549);
xor U13342 (N_13342,N_12554,N_12369);
or U13343 (N_13343,N_13181,N_12604);
xor U13344 (N_13344,N_12872,N_12947);
nand U13345 (N_13345,N_12754,N_12034);
and U13346 (N_13346,N_12213,N_12451);
xnor U13347 (N_13347,N_12974,N_13021);
xnor U13348 (N_13348,N_12639,N_13068);
nand U13349 (N_13349,N_12306,N_13094);
xor U13350 (N_13350,N_12571,N_12109);
xnor U13351 (N_13351,N_12107,N_12346);
nand U13352 (N_13352,N_12528,N_13008);
nand U13353 (N_13353,N_12223,N_12008);
or U13354 (N_13354,N_13028,N_12911);
nor U13355 (N_13355,N_13065,N_12458);
and U13356 (N_13356,N_12923,N_12121);
and U13357 (N_13357,N_12982,N_12093);
nor U13358 (N_13358,N_12565,N_13199);
nor U13359 (N_13359,N_12876,N_12897);
and U13360 (N_13360,N_12750,N_12655);
xor U13361 (N_13361,N_12832,N_12826);
nand U13362 (N_13362,N_12525,N_12416);
nand U13363 (N_13363,N_12274,N_12582);
and U13364 (N_13364,N_12503,N_13161);
nand U13365 (N_13365,N_12954,N_12322);
nor U13366 (N_13366,N_12474,N_12049);
or U13367 (N_13367,N_12077,N_12454);
xor U13368 (N_13368,N_12831,N_12975);
nor U13369 (N_13369,N_13143,N_13194);
nand U13370 (N_13370,N_13113,N_13165);
nand U13371 (N_13371,N_12751,N_12670);
xor U13372 (N_13372,N_12393,N_13114);
and U13373 (N_13373,N_12276,N_12523);
xor U13374 (N_13374,N_12361,N_12725);
nor U13375 (N_13375,N_12165,N_13196);
xnor U13376 (N_13376,N_13160,N_12723);
nand U13377 (N_13377,N_13078,N_12726);
or U13378 (N_13378,N_12634,N_12372);
nor U13379 (N_13379,N_12951,N_12137);
nand U13380 (N_13380,N_12434,N_13132);
xnor U13381 (N_13381,N_12706,N_12428);
and U13382 (N_13382,N_12380,N_12873);
and U13383 (N_13383,N_12313,N_12772);
nand U13384 (N_13384,N_12172,N_12429);
xor U13385 (N_13385,N_12889,N_12268);
or U13386 (N_13386,N_12802,N_12749);
or U13387 (N_13387,N_12041,N_12249);
nor U13388 (N_13388,N_12139,N_12882);
or U13389 (N_13389,N_12348,N_12433);
and U13390 (N_13390,N_12235,N_13179);
nor U13391 (N_13391,N_12102,N_12499);
or U13392 (N_13392,N_12941,N_13176);
or U13393 (N_13393,N_12997,N_12061);
nand U13394 (N_13394,N_12692,N_12390);
or U13395 (N_13395,N_12360,N_12405);
nand U13396 (N_13396,N_13029,N_12922);
xnor U13397 (N_13397,N_12597,N_12906);
nor U13398 (N_13398,N_12101,N_12903);
nor U13399 (N_13399,N_12968,N_12814);
nor U13400 (N_13400,N_12382,N_13145);
or U13401 (N_13401,N_12762,N_13141);
nand U13402 (N_13402,N_12470,N_12793);
nor U13403 (N_13403,N_12718,N_12122);
or U13404 (N_13404,N_12969,N_12293);
and U13405 (N_13405,N_12874,N_12009);
xnor U13406 (N_13406,N_12315,N_12753);
nor U13407 (N_13407,N_13197,N_12317);
or U13408 (N_13408,N_13066,N_12046);
xor U13409 (N_13409,N_12688,N_12144);
nor U13410 (N_13410,N_12326,N_13144);
nor U13411 (N_13411,N_12285,N_12886);
nor U13412 (N_13412,N_12167,N_12162);
xnor U13413 (N_13413,N_12849,N_12340);
nand U13414 (N_13414,N_13000,N_12893);
and U13415 (N_13415,N_12146,N_12607);
xor U13416 (N_13416,N_12888,N_12403);
nand U13417 (N_13417,N_13167,N_12052);
nor U13418 (N_13418,N_12578,N_12159);
or U13419 (N_13419,N_13023,N_12385);
and U13420 (N_13420,N_12610,N_12736);
nand U13421 (N_13421,N_12680,N_13018);
nand U13422 (N_13422,N_12778,N_12074);
nand U13423 (N_13423,N_12208,N_12868);
nand U13424 (N_13424,N_12216,N_12815);
xor U13425 (N_13425,N_12366,N_12252);
and U13426 (N_13426,N_12671,N_12409);
nor U13427 (N_13427,N_12806,N_12143);
or U13428 (N_13428,N_12224,N_12700);
nand U13429 (N_13429,N_12507,N_12447);
nand U13430 (N_13430,N_12632,N_12508);
and U13431 (N_13431,N_12432,N_12242);
xnor U13432 (N_13432,N_12659,N_13085);
nand U13433 (N_13433,N_13133,N_12803);
and U13434 (N_13434,N_12183,N_12743);
xor U13435 (N_13435,N_12482,N_12201);
nand U13436 (N_13436,N_12883,N_12197);
and U13437 (N_13437,N_12190,N_13004);
nand U13438 (N_13438,N_12761,N_12407);
and U13439 (N_13439,N_12962,N_12713);
nand U13440 (N_13440,N_12758,N_12967);
or U13441 (N_13441,N_12653,N_12933);
nand U13442 (N_13442,N_12818,N_12858);
xor U13443 (N_13443,N_12129,N_12325);
nand U13444 (N_13444,N_12605,N_12584);
nand U13445 (N_13445,N_12853,N_13019);
or U13446 (N_13446,N_12163,N_12030);
or U13447 (N_13447,N_12002,N_12358);
nand U13448 (N_13448,N_13067,N_12148);
nor U13449 (N_13449,N_12047,N_12978);
nand U13450 (N_13450,N_12734,N_12493);
nand U13451 (N_13451,N_12842,N_12044);
xnor U13452 (N_13452,N_12090,N_12838);
nand U13453 (N_13453,N_12828,N_12780);
xnor U13454 (N_13454,N_12260,N_12017);
or U13455 (N_13455,N_12126,N_12343);
xor U13456 (N_13456,N_12966,N_12965);
xor U13457 (N_13457,N_13153,N_12685);
and U13458 (N_13458,N_13128,N_12531);
nand U13459 (N_13459,N_12258,N_12981);
nand U13460 (N_13460,N_12747,N_12648);
nand U13461 (N_13461,N_12894,N_12057);
and U13462 (N_13462,N_12234,N_12901);
xor U13463 (N_13463,N_12421,N_12353);
nor U13464 (N_13464,N_12050,N_12658);
nor U13465 (N_13465,N_12158,N_12596);
and U13466 (N_13466,N_12973,N_12952);
or U13467 (N_13467,N_12730,N_12866);
nor U13468 (N_13468,N_12419,N_12567);
or U13469 (N_13469,N_12786,N_12177);
nand U13470 (N_13470,N_12070,N_12675);
and U13471 (N_13471,N_12479,N_12444);
xor U13472 (N_13472,N_12830,N_12220);
and U13473 (N_13473,N_12637,N_12209);
xor U13474 (N_13474,N_12245,N_13155);
or U13475 (N_13475,N_12179,N_13106);
xor U13476 (N_13476,N_12944,N_12387);
nor U13477 (N_13477,N_12305,N_12150);
nand U13478 (N_13478,N_12708,N_12205);
xnor U13479 (N_13479,N_12783,N_12937);
and U13480 (N_13480,N_12927,N_13057);
and U13481 (N_13481,N_12247,N_12494);
and U13482 (N_13482,N_12032,N_13039);
nor U13483 (N_13483,N_13015,N_13031);
xnor U13484 (N_13484,N_12501,N_12645);
nand U13485 (N_13485,N_12059,N_12191);
nand U13486 (N_13486,N_12468,N_12384);
xnor U13487 (N_13487,N_13142,N_12067);
nor U13488 (N_13488,N_12770,N_12357);
nor U13489 (N_13489,N_12697,N_12477);
xnor U13490 (N_13490,N_12765,N_12194);
or U13491 (N_13491,N_12776,N_12759);
nand U13492 (N_13492,N_13107,N_12112);
nor U13493 (N_13493,N_12825,N_12000);
nand U13494 (N_13494,N_12232,N_12441);
nor U13495 (N_13495,N_12467,N_12703);
and U13496 (N_13496,N_12231,N_12110);
and U13497 (N_13497,N_12427,N_13169);
nand U13498 (N_13498,N_12298,N_12069);
or U13499 (N_13499,N_13139,N_12649);
and U13500 (N_13500,N_12796,N_12138);
and U13501 (N_13501,N_13125,N_12677);
nand U13502 (N_13502,N_12006,N_12733);
or U13503 (N_13503,N_12033,N_12288);
and U13504 (N_13504,N_12086,N_12133);
xor U13505 (N_13505,N_12054,N_12096);
nand U13506 (N_13506,N_13159,N_12445);
xor U13507 (N_13507,N_12273,N_12111);
xor U13508 (N_13508,N_12993,N_12323);
or U13509 (N_13509,N_12092,N_13080);
xnor U13510 (N_13510,N_12238,N_12711);
and U13511 (N_13511,N_13157,N_12992);
nor U13512 (N_13512,N_12843,N_12586);
and U13513 (N_13513,N_13045,N_13083);
and U13514 (N_13514,N_12614,N_12472);
nand U13515 (N_13515,N_12460,N_12964);
nand U13516 (N_13516,N_12236,N_12912);
nand U13517 (N_13517,N_12774,N_13190);
and U13518 (N_13518,N_12140,N_12412);
nor U13519 (N_13519,N_13121,N_12379);
or U13520 (N_13520,N_12316,N_13017);
xor U13521 (N_13521,N_12792,N_12038);
nand U13522 (N_13522,N_12988,N_12990);
nand U13523 (N_13523,N_12946,N_12355);
nor U13524 (N_13524,N_12976,N_13082);
nand U13525 (N_13525,N_12650,N_12106);
xnor U13526 (N_13526,N_12024,N_12885);
xnor U13527 (N_13527,N_12629,N_12295);
nor U13528 (N_13528,N_12919,N_12048);
xor U13529 (N_13529,N_12099,N_12797);
nor U13530 (N_13530,N_13116,N_12058);
or U13531 (N_13531,N_12587,N_12727);
nor U13532 (N_13532,N_12204,N_12784);
nand U13533 (N_13533,N_13117,N_13014);
nand U13534 (N_13534,N_12391,N_12085);
xnor U13535 (N_13535,N_12496,N_13171);
and U13536 (N_13536,N_13062,N_13073);
nand U13537 (N_13537,N_13135,N_12617);
xor U13538 (N_13538,N_12378,N_12816);
xor U13539 (N_13539,N_12704,N_12053);
or U13540 (N_13540,N_12928,N_12514);
or U13541 (N_13541,N_12594,N_12899);
xor U13542 (N_13542,N_12592,N_12767);
nor U13543 (N_13543,N_12518,N_12022);
and U13544 (N_13544,N_12729,N_12603);
nand U13545 (N_13545,N_12491,N_12178);
nor U13546 (N_13546,N_13192,N_12691);
xor U13547 (N_13547,N_12446,N_13088);
or U13548 (N_13548,N_12036,N_12924);
nand U13549 (N_13549,N_12576,N_12365);
nor U13550 (N_13550,N_12275,N_12134);
or U13551 (N_13551,N_12004,N_12188);
or U13552 (N_13552,N_12170,N_13049);
or U13553 (N_13553,N_13150,N_12877);
xnor U13554 (N_13554,N_12120,N_12214);
nor U13555 (N_13555,N_13131,N_12226);
and U13556 (N_13556,N_12820,N_13184);
nand U13557 (N_13557,N_12042,N_12375);
and U13558 (N_13558,N_12517,N_12267);
and U13559 (N_13559,N_12536,N_13081);
nor U13560 (N_13560,N_12255,N_12846);
or U13561 (N_13561,N_13055,N_12130);
nor U13562 (N_13562,N_12504,N_12064);
and U13563 (N_13563,N_12695,N_12715);
and U13564 (N_13564,N_13038,N_12324);
or U13565 (N_13565,N_12892,N_12495);
nand U13566 (N_13566,N_12773,N_12151);
and U13567 (N_13567,N_12464,N_12280);
nor U13568 (N_13568,N_12081,N_13046);
and U13569 (N_13569,N_12283,N_12203);
nor U13570 (N_13570,N_12662,N_12694);
or U13571 (N_13571,N_12745,N_12485);
xnor U13572 (N_13572,N_12955,N_12473);
nor U13573 (N_13573,N_13009,N_12502);
and U13574 (N_13574,N_12505,N_12626);
or U13575 (N_13575,N_13092,N_12850);
and U13576 (N_13576,N_12782,N_12710);
xor U13577 (N_13577,N_12210,N_12256);
or U13578 (N_13578,N_12979,N_12511);
and U13579 (N_13579,N_12015,N_12272);
or U13580 (N_13580,N_12469,N_12557);
and U13581 (N_13581,N_12940,N_13188);
nor U13582 (N_13582,N_12233,N_12821);
and U13583 (N_13583,N_12012,N_12613);
xor U13584 (N_13584,N_12907,N_12851);
or U13585 (N_13585,N_12945,N_12406);
nor U13586 (N_13586,N_12334,N_13186);
and U13587 (N_13587,N_12702,N_13089);
or U13588 (N_13588,N_12622,N_12938);
or U13589 (N_13589,N_13013,N_13048);
xnor U13590 (N_13590,N_12001,N_12705);
nand U13591 (N_13591,N_12181,N_12195);
nor U13592 (N_13592,N_12953,N_12795);
xnor U13593 (N_13593,N_12027,N_12593);
nand U13594 (N_13594,N_12683,N_13043);
or U13595 (N_13595,N_12330,N_13050);
nand U13596 (N_13596,N_12174,N_12798);
nand U13597 (N_13597,N_12098,N_12302);
nor U13598 (N_13598,N_12153,N_12570);
xnor U13599 (N_13599,N_12534,N_12229);
xor U13600 (N_13600,N_12644,N_12867);
or U13601 (N_13601,N_12215,N_12359);
nand U13602 (N_13602,N_12332,N_12011);
nor U13603 (N_13603,N_12948,N_12995);
or U13604 (N_13604,N_12080,N_13061);
nor U13605 (N_13605,N_13109,N_12665);
xnor U13606 (N_13606,N_12463,N_12055);
nor U13607 (N_13607,N_13172,N_12986);
xor U13608 (N_13608,N_12342,N_12588);
nand U13609 (N_13609,N_13084,N_12926);
nor U13610 (N_13610,N_12014,N_12212);
nand U13611 (N_13611,N_12533,N_13064);
nor U13612 (N_13612,N_12573,N_13111);
xnor U13613 (N_13613,N_13010,N_13096);
nor U13614 (N_13614,N_12914,N_12537);
nor U13615 (N_13615,N_12744,N_12389);
nor U13616 (N_13616,N_12127,N_12339);
xor U13617 (N_13617,N_12457,N_12693);
or U13618 (N_13618,N_12555,N_12399);
nand U13619 (N_13619,N_12985,N_12424);
xor U13620 (N_13620,N_12513,N_12510);
nor U13621 (N_13621,N_12775,N_13007);
or U13622 (N_13622,N_12091,N_13070);
and U13623 (N_13623,N_12264,N_12310);
xor U13624 (N_13624,N_12386,N_12029);
nand U13625 (N_13625,N_12300,N_12721);
and U13626 (N_13626,N_12777,N_12476);
and U13627 (N_13627,N_12337,N_12413);
nor U13628 (N_13628,N_12871,N_12991);
xnor U13629 (N_13629,N_12546,N_12630);
xnor U13630 (N_13630,N_12701,N_12996);
nor U13631 (N_13631,N_12987,N_12539);
nand U13632 (N_13632,N_12519,N_12171);
nand U13633 (N_13633,N_12949,N_12418);
and U13634 (N_13634,N_12396,N_12977);
and U13635 (N_13635,N_13002,N_12529);
or U13636 (N_13636,N_12368,N_12887);
xnor U13637 (N_13637,N_12625,N_12575);
nand U13638 (N_13638,N_12520,N_12647);
xor U13639 (N_13639,N_12279,N_12600);
nor U13640 (N_13640,N_12807,N_13136);
or U13641 (N_13641,N_12819,N_12568);
and U13642 (N_13642,N_13140,N_12269);
or U13643 (N_13643,N_13162,N_12735);
nand U13644 (N_13644,N_12222,N_12908);
nor U13645 (N_13645,N_12075,N_12515);
xnor U13646 (N_13646,N_12344,N_12155);
or U13647 (N_13647,N_12724,N_13129);
or U13648 (N_13648,N_13173,N_12455);
and U13649 (N_13649,N_12667,N_12552);
xor U13650 (N_13650,N_12720,N_12089);
and U13651 (N_13651,N_12282,N_12931);
and U13652 (N_13652,N_12010,N_12363);
or U13653 (N_13653,N_12374,N_12564);
nor U13654 (N_13654,N_12714,N_12423);
or U13655 (N_13655,N_13076,N_12410);
nor U13656 (N_13656,N_12497,N_12250);
xor U13657 (N_13657,N_13086,N_12169);
xnor U13658 (N_13658,N_12656,N_12739);
xnor U13659 (N_13659,N_12082,N_12301);
nor U13660 (N_13660,N_12755,N_12286);
xor U13661 (N_13661,N_12025,N_12543);
or U13662 (N_13662,N_12712,N_13093);
nand U13663 (N_13663,N_13183,N_12994);
nor U13664 (N_13664,N_12349,N_12860);
xnor U13665 (N_13665,N_12186,N_12088);
nand U13666 (N_13666,N_12623,N_12642);
nor U13667 (N_13667,N_12608,N_12813);
nand U13668 (N_13668,N_12611,N_12898);
xor U13669 (N_13669,N_13032,N_12490);
nand U13670 (N_13670,N_13001,N_12633);
and U13671 (N_13671,N_12230,N_12475);
nor U13672 (N_13672,N_12362,N_12251);
nor U13673 (N_13673,N_12294,N_12696);
or U13674 (N_13674,N_13063,N_13177);
xnor U13675 (N_13675,N_12240,N_13079);
or U13676 (N_13676,N_12328,N_12388);
xnor U13677 (N_13677,N_12553,N_12855);
nor U13678 (N_13678,N_12942,N_12123);
and U13679 (N_13679,N_13108,N_13069);
and U13680 (N_13680,N_12459,N_12583);
or U13681 (N_13681,N_12581,N_12936);
or U13682 (N_13682,N_12338,N_12771);
nand U13683 (N_13683,N_13112,N_13040);
or U13684 (N_13684,N_12350,N_12438);
or U13685 (N_13685,N_12408,N_12045);
or U13686 (N_13686,N_12013,N_13166);
nor U13687 (N_13687,N_12654,N_12663);
nor U13688 (N_13688,N_12556,N_12307);
nor U13689 (N_13689,N_12522,N_13072);
xnor U13690 (N_13690,N_12227,N_12443);
and U13691 (N_13691,N_13130,N_12347);
nand U13692 (N_13692,N_12426,N_12060);
nand U13693 (N_13693,N_12119,N_12287);
nor U13694 (N_13694,N_12620,N_12196);
or U13695 (N_13695,N_12243,N_12561);
nor U13696 (N_13696,N_12512,N_12527);
or U13697 (N_13697,N_12453,N_12271);
nor U13698 (N_13698,N_13030,N_12125);
nand U13699 (N_13699,N_12550,N_12402);
xor U13700 (N_13700,N_12321,N_12198);
or U13701 (N_13701,N_12844,N_12878);
and U13702 (N_13702,N_12863,N_12763);
xor U13703 (N_13703,N_12161,N_13074);
and U13704 (N_13704,N_12456,N_12105);
nor U13705 (N_13705,N_12142,N_12616);
and U13706 (N_13706,N_12563,N_12804);
nand U13707 (N_13707,N_12548,N_12094);
xor U13708 (N_13708,N_12950,N_12430);
and U13709 (N_13709,N_12506,N_12805);
nand U13710 (N_13710,N_12354,N_13095);
or U13711 (N_13711,N_12019,N_12259);
xnor U13712 (N_13712,N_12113,N_12848);
xnor U13713 (N_13713,N_12411,N_12498);
nor U13714 (N_13714,N_12627,N_12652);
or U13715 (N_13715,N_13154,N_13041);
xnor U13716 (N_13716,N_12681,N_12538);
or U13717 (N_13717,N_12461,N_12535);
nor U13718 (N_13718,N_12917,N_12601);
nand U13719 (N_13719,N_12182,N_12862);
nand U13720 (N_13720,N_12827,N_12483);
and U13721 (N_13721,N_12311,N_12290);
xor U13722 (N_13722,N_12672,N_13158);
or U13723 (N_13723,N_12891,N_12824);
nor U13724 (N_13724,N_13191,N_12913);
xor U13725 (N_13725,N_12834,N_13042);
nand U13726 (N_13726,N_12682,N_12465);
nor U13727 (N_13727,N_12526,N_12478);
nand U13728 (N_13728,N_12732,N_12035);
or U13729 (N_13729,N_12442,N_12808);
and U13730 (N_13730,N_13016,N_12377);
nor U13731 (N_13731,N_12930,N_12211);
nor U13732 (N_13732,N_12547,N_13148);
xor U13733 (N_13733,N_12768,N_12202);
nor U13734 (N_13734,N_13036,N_12524);
nor U13735 (N_13735,N_13187,N_13127);
nor U13736 (N_13736,N_12237,N_12562);
or U13737 (N_13737,N_13012,N_12073);
and U13738 (N_13738,N_12117,N_12787);
xnor U13739 (N_13739,N_12023,N_12870);
nand U13740 (N_13740,N_12481,N_12932);
xor U13741 (N_13741,N_13185,N_13033);
nand U13742 (N_13742,N_12666,N_12076);
or U13743 (N_13743,N_12651,N_12166);
nand U13744 (N_13744,N_12329,N_12248);
xor U13745 (N_13745,N_13052,N_12840);
or U13746 (N_13746,N_12687,N_12861);
and U13747 (N_13747,N_13195,N_12381);
nand U13748 (N_13748,N_13156,N_12875);
xnor U13749 (N_13749,N_12920,N_12833);
xor U13750 (N_13750,N_12281,N_12835);
xnor U13751 (N_13751,N_12395,N_12881);
nor U13752 (N_13752,N_13011,N_12686);
xnor U13753 (N_13753,N_12132,N_12309);
xor U13754 (N_13754,N_12303,N_12173);
or U13755 (N_13755,N_12956,N_12439);
nand U13756 (N_13756,N_12452,N_12200);
nand U13757 (N_13757,N_12559,N_13051);
xor U13758 (N_13758,N_12852,N_13175);
nor U13759 (N_13759,N_12296,N_13058);
xor U13760 (N_13760,N_12270,N_12545);
and U13761 (N_13761,N_12487,N_13152);
or U13762 (N_13762,N_12530,N_12095);
or U13763 (N_13763,N_12160,N_13170);
or U13764 (N_13764,N_12420,N_12124);
nand U13765 (N_13765,N_12062,N_12261);
nand U13766 (N_13766,N_12097,N_13189);
xnor U13767 (N_13767,N_12056,N_12401);
nand U13768 (N_13768,N_12319,N_12488);
and U13769 (N_13769,N_12621,N_12925);
nand U13770 (N_13770,N_12631,N_12068);
xnor U13771 (N_13771,N_12921,N_12292);
nor U13772 (N_13772,N_13005,N_12935);
nand U13773 (N_13773,N_13123,N_12864);
and U13774 (N_13774,N_12540,N_12417);
or U13775 (N_13775,N_13003,N_13102);
xnor U13776 (N_13776,N_12963,N_12934);
xor U13777 (N_13777,N_12152,N_12318);
nor U13778 (N_13778,N_12314,N_13098);
and U13779 (N_13779,N_12404,N_13020);
nor U13780 (N_13780,N_12789,N_12492);
nor U13781 (N_13781,N_12895,N_12972);
and U13782 (N_13782,N_13090,N_13103);
nor U13783 (N_13783,N_12716,N_12003);
or U13784 (N_13784,N_12661,N_12135);
nand U13785 (N_13785,N_12072,N_12154);
nand U13786 (N_13786,N_12591,N_12574);
nor U13787 (N_13787,N_13163,N_12175);
and U13788 (N_13788,N_12118,N_13118);
or U13789 (N_13789,N_12748,N_12590);
nor U13790 (N_13790,N_12450,N_12943);
and U13791 (N_13791,N_12239,N_12722);
nor U13792 (N_13792,N_12764,N_12638);
nand U13793 (N_13793,N_12168,N_12669);
or U13794 (N_13794,N_12007,N_12071);
nor U13795 (N_13795,N_12856,N_12957);
xnor U13796 (N_13796,N_13120,N_12207);
nand U13797 (N_13797,N_13110,N_12383);
xnor U13798 (N_13798,N_12079,N_12989);
or U13799 (N_13799,N_13100,N_13134);
nor U13800 (N_13800,N_12422,N_12704);
nand U13801 (N_13801,N_12037,N_12591);
xor U13802 (N_13802,N_12602,N_12731);
nor U13803 (N_13803,N_13089,N_12111);
and U13804 (N_13804,N_12629,N_12133);
nor U13805 (N_13805,N_12737,N_12972);
nand U13806 (N_13806,N_12462,N_12203);
nand U13807 (N_13807,N_12468,N_12899);
nor U13808 (N_13808,N_12421,N_12791);
nor U13809 (N_13809,N_12326,N_12463);
nor U13810 (N_13810,N_13100,N_12891);
xor U13811 (N_13811,N_12659,N_12364);
xnor U13812 (N_13812,N_12057,N_13159);
nor U13813 (N_13813,N_13082,N_12502);
or U13814 (N_13814,N_12857,N_12044);
nand U13815 (N_13815,N_12058,N_13181);
xnor U13816 (N_13816,N_12001,N_12567);
nor U13817 (N_13817,N_12662,N_12159);
nor U13818 (N_13818,N_12314,N_12666);
nand U13819 (N_13819,N_13156,N_12352);
and U13820 (N_13820,N_12408,N_12390);
and U13821 (N_13821,N_12534,N_12467);
or U13822 (N_13822,N_12991,N_13033);
xnor U13823 (N_13823,N_12472,N_12920);
or U13824 (N_13824,N_12099,N_13018);
xnor U13825 (N_13825,N_12401,N_12625);
nor U13826 (N_13826,N_12888,N_12885);
and U13827 (N_13827,N_12568,N_12069);
and U13828 (N_13828,N_12690,N_12298);
nor U13829 (N_13829,N_12558,N_13117);
nand U13830 (N_13830,N_12623,N_12409);
xor U13831 (N_13831,N_12008,N_12044);
and U13832 (N_13832,N_12869,N_12916);
nand U13833 (N_13833,N_12252,N_12647);
and U13834 (N_13834,N_12880,N_12604);
or U13835 (N_13835,N_12449,N_12197);
nand U13836 (N_13836,N_12810,N_12317);
nor U13837 (N_13837,N_12281,N_12138);
and U13838 (N_13838,N_12739,N_12486);
nand U13839 (N_13839,N_12058,N_13081);
or U13840 (N_13840,N_12694,N_12692);
nand U13841 (N_13841,N_12321,N_12762);
or U13842 (N_13842,N_12276,N_13186);
or U13843 (N_13843,N_12084,N_12333);
or U13844 (N_13844,N_12533,N_12520);
or U13845 (N_13845,N_12364,N_12832);
or U13846 (N_13846,N_12470,N_12181);
and U13847 (N_13847,N_12303,N_12790);
xor U13848 (N_13848,N_12438,N_12595);
nand U13849 (N_13849,N_12787,N_12604);
nor U13850 (N_13850,N_13179,N_12288);
nand U13851 (N_13851,N_12099,N_13066);
and U13852 (N_13852,N_12620,N_12409);
and U13853 (N_13853,N_12040,N_12446);
and U13854 (N_13854,N_12790,N_12837);
nand U13855 (N_13855,N_12642,N_12131);
nor U13856 (N_13856,N_12940,N_12251);
nand U13857 (N_13857,N_12902,N_13074);
nand U13858 (N_13858,N_12575,N_12721);
or U13859 (N_13859,N_12845,N_13193);
nor U13860 (N_13860,N_12629,N_12582);
or U13861 (N_13861,N_12366,N_13039);
and U13862 (N_13862,N_12615,N_12600);
and U13863 (N_13863,N_12043,N_12434);
nor U13864 (N_13864,N_12838,N_12588);
and U13865 (N_13865,N_12718,N_12089);
and U13866 (N_13866,N_12483,N_12118);
or U13867 (N_13867,N_13135,N_12204);
or U13868 (N_13868,N_12263,N_13140);
xor U13869 (N_13869,N_12061,N_12509);
xnor U13870 (N_13870,N_12619,N_13033);
xor U13871 (N_13871,N_12959,N_13040);
or U13872 (N_13872,N_13003,N_12453);
xor U13873 (N_13873,N_12297,N_12108);
nor U13874 (N_13874,N_13001,N_13162);
nor U13875 (N_13875,N_12042,N_12378);
nand U13876 (N_13876,N_12888,N_12364);
nor U13877 (N_13877,N_12839,N_12875);
or U13878 (N_13878,N_12844,N_12776);
or U13879 (N_13879,N_12223,N_12579);
nor U13880 (N_13880,N_12891,N_12388);
and U13881 (N_13881,N_12172,N_12627);
or U13882 (N_13882,N_12690,N_12265);
nand U13883 (N_13883,N_12193,N_12245);
nor U13884 (N_13884,N_12561,N_12964);
and U13885 (N_13885,N_12075,N_12514);
nor U13886 (N_13886,N_12484,N_12083);
or U13887 (N_13887,N_12382,N_12384);
xnor U13888 (N_13888,N_12778,N_12160);
or U13889 (N_13889,N_12123,N_12163);
nor U13890 (N_13890,N_12330,N_12398);
and U13891 (N_13891,N_12311,N_13085);
or U13892 (N_13892,N_12017,N_12002);
and U13893 (N_13893,N_12742,N_12363);
and U13894 (N_13894,N_12016,N_12835);
or U13895 (N_13895,N_12423,N_12849);
nand U13896 (N_13896,N_13136,N_13089);
nor U13897 (N_13897,N_12494,N_12641);
and U13898 (N_13898,N_13054,N_12330);
and U13899 (N_13899,N_12348,N_12186);
xor U13900 (N_13900,N_12760,N_12955);
nor U13901 (N_13901,N_13109,N_12534);
nand U13902 (N_13902,N_13040,N_12673);
xor U13903 (N_13903,N_12159,N_12870);
nor U13904 (N_13904,N_12972,N_12134);
or U13905 (N_13905,N_12977,N_12242);
and U13906 (N_13906,N_12930,N_12214);
or U13907 (N_13907,N_12058,N_13146);
and U13908 (N_13908,N_12615,N_12466);
or U13909 (N_13909,N_13181,N_12359);
xor U13910 (N_13910,N_13116,N_13136);
nor U13911 (N_13911,N_12643,N_12728);
xnor U13912 (N_13912,N_12967,N_12773);
nand U13913 (N_13913,N_13003,N_12999);
or U13914 (N_13914,N_12524,N_13131);
xor U13915 (N_13915,N_12877,N_12575);
xor U13916 (N_13916,N_12658,N_12796);
nand U13917 (N_13917,N_12777,N_13019);
xor U13918 (N_13918,N_13126,N_12268);
nand U13919 (N_13919,N_12411,N_13052);
and U13920 (N_13920,N_12914,N_12627);
xnor U13921 (N_13921,N_12403,N_12763);
xor U13922 (N_13922,N_13113,N_12543);
and U13923 (N_13923,N_12711,N_12133);
xor U13924 (N_13924,N_12606,N_13022);
xor U13925 (N_13925,N_12308,N_12972);
or U13926 (N_13926,N_12119,N_12833);
nor U13927 (N_13927,N_13021,N_12445);
xnor U13928 (N_13928,N_12332,N_12699);
xor U13929 (N_13929,N_12665,N_12672);
and U13930 (N_13930,N_12679,N_12048);
nand U13931 (N_13931,N_12617,N_12449);
nand U13932 (N_13932,N_12741,N_12527);
nand U13933 (N_13933,N_12869,N_12276);
xnor U13934 (N_13934,N_12308,N_12941);
and U13935 (N_13935,N_12909,N_12231);
xor U13936 (N_13936,N_12290,N_13118);
and U13937 (N_13937,N_12144,N_12207);
and U13938 (N_13938,N_12360,N_12732);
xor U13939 (N_13939,N_12460,N_12618);
nor U13940 (N_13940,N_12029,N_12597);
nor U13941 (N_13941,N_12296,N_12435);
and U13942 (N_13942,N_12901,N_12722);
and U13943 (N_13943,N_12162,N_12105);
and U13944 (N_13944,N_12619,N_12205);
nand U13945 (N_13945,N_13096,N_12159);
nand U13946 (N_13946,N_12867,N_12522);
nor U13947 (N_13947,N_13184,N_12023);
nor U13948 (N_13948,N_12920,N_12619);
xor U13949 (N_13949,N_12135,N_12330);
nor U13950 (N_13950,N_12749,N_12441);
or U13951 (N_13951,N_12385,N_12446);
or U13952 (N_13952,N_12913,N_13029);
or U13953 (N_13953,N_13129,N_12985);
and U13954 (N_13954,N_13053,N_12077);
or U13955 (N_13955,N_12847,N_12247);
xor U13956 (N_13956,N_12434,N_12491);
nand U13957 (N_13957,N_13140,N_12404);
nand U13958 (N_13958,N_12749,N_12492);
or U13959 (N_13959,N_12849,N_12164);
or U13960 (N_13960,N_12923,N_12656);
or U13961 (N_13961,N_12930,N_12468);
xor U13962 (N_13962,N_12490,N_12366);
nand U13963 (N_13963,N_12039,N_12530);
or U13964 (N_13964,N_12092,N_12190);
nand U13965 (N_13965,N_12071,N_12682);
xnor U13966 (N_13966,N_12928,N_12094);
xnor U13967 (N_13967,N_12235,N_12703);
nor U13968 (N_13968,N_13162,N_12188);
nand U13969 (N_13969,N_12931,N_12091);
xnor U13970 (N_13970,N_12460,N_12328);
xor U13971 (N_13971,N_13078,N_12692);
nor U13972 (N_13972,N_12185,N_12002);
nor U13973 (N_13973,N_12784,N_12802);
xor U13974 (N_13974,N_12887,N_13104);
nand U13975 (N_13975,N_12554,N_12640);
xnor U13976 (N_13976,N_12503,N_13109);
xor U13977 (N_13977,N_13155,N_12881);
nor U13978 (N_13978,N_13130,N_12373);
and U13979 (N_13979,N_12946,N_12955);
nor U13980 (N_13980,N_12364,N_13102);
nand U13981 (N_13981,N_12178,N_12510);
xor U13982 (N_13982,N_13194,N_12112);
nor U13983 (N_13983,N_12789,N_12143);
or U13984 (N_13984,N_12614,N_12255);
nor U13985 (N_13985,N_12449,N_12641);
and U13986 (N_13986,N_12270,N_12184);
or U13987 (N_13987,N_12916,N_12159);
xor U13988 (N_13988,N_12481,N_12877);
and U13989 (N_13989,N_12377,N_12164);
nor U13990 (N_13990,N_12872,N_12011);
nand U13991 (N_13991,N_12618,N_12030);
nand U13992 (N_13992,N_12815,N_12683);
nor U13993 (N_13993,N_12734,N_12834);
and U13994 (N_13994,N_12104,N_12113);
nor U13995 (N_13995,N_12717,N_12552);
nor U13996 (N_13996,N_12630,N_13199);
nand U13997 (N_13997,N_12911,N_12947);
xnor U13998 (N_13998,N_12105,N_12917);
and U13999 (N_13999,N_12480,N_13116);
and U14000 (N_14000,N_12964,N_12408);
xnor U14001 (N_14001,N_12155,N_12334);
nor U14002 (N_14002,N_12382,N_12306);
and U14003 (N_14003,N_12037,N_12903);
or U14004 (N_14004,N_12784,N_12533);
nor U14005 (N_14005,N_13084,N_12079);
nand U14006 (N_14006,N_12259,N_13011);
and U14007 (N_14007,N_12285,N_12316);
nand U14008 (N_14008,N_12474,N_12835);
nor U14009 (N_14009,N_12942,N_12744);
nor U14010 (N_14010,N_12380,N_12109);
or U14011 (N_14011,N_12719,N_12316);
xor U14012 (N_14012,N_13117,N_12017);
nand U14013 (N_14013,N_12022,N_12371);
nor U14014 (N_14014,N_12662,N_12145);
and U14015 (N_14015,N_12668,N_13140);
or U14016 (N_14016,N_12414,N_12270);
or U14017 (N_14017,N_12046,N_12186);
nor U14018 (N_14018,N_12959,N_12845);
or U14019 (N_14019,N_12450,N_12961);
nand U14020 (N_14020,N_12288,N_12287);
nor U14021 (N_14021,N_13022,N_12560);
nor U14022 (N_14022,N_12827,N_12160);
nand U14023 (N_14023,N_12828,N_12614);
and U14024 (N_14024,N_12542,N_12303);
and U14025 (N_14025,N_13137,N_12072);
or U14026 (N_14026,N_12203,N_12349);
and U14027 (N_14027,N_12959,N_12601);
or U14028 (N_14028,N_13074,N_12081);
xor U14029 (N_14029,N_12924,N_13042);
or U14030 (N_14030,N_12200,N_12139);
nor U14031 (N_14031,N_12599,N_12499);
and U14032 (N_14032,N_12500,N_12732);
and U14033 (N_14033,N_12831,N_12543);
xnor U14034 (N_14034,N_12597,N_12033);
nor U14035 (N_14035,N_12577,N_12774);
or U14036 (N_14036,N_12127,N_12934);
nor U14037 (N_14037,N_12686,N_12702);
or U14038 (N_14038,N_13184,N_12487);
nand U14039 (N_14039,N_12754,N_12352);
and U14040 (N_14040,N_13127,N_12304);
nand U14041 (N_14041,N_12221,N_12287);
and U14042 (N_14042,N_12082,N_12552);
xor U14043 (N_14043,N_12972,N_12119);
nand U14044 (N_14044,N_12458,N_12004);
xor U14045 (N_14045,N_12491,N_12655);
and U14046 (N_14046,N_12907,N_13196);
xor U14047 (N_14047,N_13060,N_12470);
or U14048 (N_14048,N_13009,N_13161);
and U14049 (N_14049,N_13019,N_12801);
xor U14050 (N_14050,N_12975,N_12762);
nand U14051 (N_14051,N_12530,N_12007);
or U14052 (N_14052,N_13180,N_13134);
xnor U14053 (N_14053,N_12586,N_12350);
nor U14054 (N_14054,N_13122,N_12277);
nand U14055 (N_14055,N_12901,N_12284);
nor U14056 (N_14056,N_13186,N_12037);
xor U14057 (N_14057,N_12466,N_12343);
nor U14058 (N_14058,N_13013,N_12928);
nor U14059 (N_14059,N_12057,N_12284);
and U14060 (N_14060,N_12440,N_13029);
and U14061 (N_14061,N_12651,N_12747);
and U14062 (N_14062,N_12370,N_12636);
nand U14063 (N_14063,N_12689,N_12045);
or U14064 (N_14064,N_13027,N_13196);
xnor U14065 (N_14065,N_13002,N_12332);
nor U14066 (N_14066,N_12857,N_12870);
or U14067 (N_14067,N_12168,N_13056);
nor U14068 (N_14068,N_12687,N_12910);
nand U14069 (N_14069,N_12064,N_13005);
or U14070 (N_14070,N_13189,N_12270);
nor U14071 (N_14071,N_12977,N_12305);
or U14072 (N_14072,N_12468,N_13083);
and U14073 (N_14073,N_12975,N_12938);
nor U14074 (N_14074,N_12376,N_12052);
and U14075 (N_14075,N_12291,N_12958);
nand U14076 (N_14076,N_12375,N_12062);
nor U14077 (N_14077,N_12030,N_12365);
or U14078 (N_14078,N_12873,N_12105);
and U14079 (N_14079,N_12860,N_12680);
xnor U14080 (N_14080,N_12694,N_12503);
and U14081 (N_14081,N_12094,N_12362);
nand U14082 (N_14082,N_12654,N_12968);
nand U14083 (N_14083,N_12912,N_12874);
nor U14084 (N_14084,N_12075,N_13008);
or U14085 (N_14085,N_12962,N_12388);
xor U14086 (N_14086,N_12646,N_12333);
nor U14087 (N_14087,N_13110,N_12691);
nand U14088 (N_14088,N_12399,N_12932);
and U14089 (N_14089,N_12619,N_12707);
xor U14090 (N_14090,N_12020,N_12740);
nand U14091 (N_14091,N_12037,N_12308);
nor U14092 (N_14092,N_12607,N_12534);
nor U14093 (N_14093,N_12698,N_13105);
nand U14094 (N_14094,N_12766,N_13063);
nand U14095 (N_14095,N_12968,N_12873);
and U14096 (N_14096,N_12501,N_12181);
xor U14097 (N_14097,N_13190,N_12416);
xor U14098 (N_14098,N_12264,N_13074);
nor U14099 (N_14099,N_12774,N_12920);
nand U14100 (N_14100,N_12203,N_12807);
or U14101 (N_14101,N_12786,N_13070);
xor U14102 (N_14102,N_12921,N_12066);
or U14103 (N_14103,N_12225,N_13125);
nor U14104 (N_14104,N_13165,N_13035);
nand U14105 (N_14105,N_12432,N_12440);
xnor U14106 (N_14106,N_12697,N_12109);
xnor U14107 (N_14107,N_12549,N_12866);
or U14108 (N_14108,N_12921,N_12155);
and U14109 (N_14109,N_12141,N_12496);
nor U14110 (N_14110,N_13129,N_12803);
xor U14111 (N_14111,N_12394,N_12486);
xor U14112 (N_14112,N_12515,N_12004);
and U14113 (N_14113,N_12265,N_12196);
xnor U14114 (N_14114,N_12820,N_12169);
xor U14115 (N_14115,N_13166,N_12862);
and U14116 (N_14116,N_12888,N_12170);
nor U14117 (N_14117,N_12977,N_13064);
nand U14118 (N_14118,N_12857,N_12419);
nand U14119 (N_14119,N_13169,N_12751);
nor U14120 (N_14120,N_12629,N_12904);
nand U14121 (N_14121,N_12851,N_12402);
or U14122 (N_14122,N_12772,N_12378);
or U14123 (N_14123,N_12621,N_13015);
xor U14124 (N_14124,N_12343,N_13102);
nor U14125 (N_14125,N_13028,N_12560);
xor U14126 (N_14126,N_13169,N_12875);
and U14127 (N_14127,N_12814,N_12976);
nor U14128 (N_14128,N_12006,N_12284);
xnor U14129 (N_14129,N_13096,N_12462);
nor U14130 (N_14130,N_13031,N_13025);
nor U14131 (N_14131,N_13004,N_12184);
nand U14132 (N_14132,N_12913,N_12381);
xor U14133 (N_14133,N_13184,N_13056);
nand U14134 (N_14134,N_13059,N_12994);
nand U14135 (N_14135,N_12014,N_12307);
and U14136 (N_14136,N_12692,N_13119);
nand U14137 (N_14137,N_12960,N_12331);
xnor U14138 (N_14138,N_12385,N_12915);
nor U14139 (N_14139,N_12453,N_13119);
and U14140 (N_14140,N_12487,N_12024);
xnor U14141 (N_14141,N_13154,N_12461);
and U14142 (N_14142,N_12646,N_12503);
xnor U14143 (N_14143,N_12707,N_12003);
xor U14144 (N_14144,N_12220,N_12893);
xnor U14145 (N_14145,N_12021,N_13043);
nor U14146 (N_14146,N_12952,N_12962);
nor U14147 (N_14147,N_13182,N_12707);
or U14148 (N_14148,N_12680,N_12621);
xor U14149 (N_14149,N_12075,N_13130);
nor U14150 (N_14150,N_12723,N_12244);
or U14151 (N_14151,N_12256,N_12399);
nor U14152 (N_14152,N_12986,N_12273);
nand U14153 (N_14153,N_12505,N_12068);
nor U14154 (N_14154,N_12364,N_12776);
xnor U14155 (N_14155,N_12348,N_12582);
xor U14156 (N_14156,N_12662,N_12346);
xnor U14157 (N_14157,N_12469,N_12263);
or U14158 (N_14158,N_12852,N_13109);
and U14159 (N_14159,N_12609,N_13005);
nand U14160 (N_14160,N_12406,N_12671);
and U14161 (N_14161,N_12630,N_12645);
and U14162 (N_14162,N_12368,N_12543);
or U14163 (N_14163,N_12484,N_13195);
nand U14164 (N_14164,N_12944,N_12895);
and U14165 (N_14165,N_12714,N_12351);
and U14166 (N_14166,N_12283,N_12744);
nor U14167 (N_14167,N_13000,N_12043);
xor U14168 (N_14168,N_12882,N_12835);
or U14169 (N_14169,N_12325,N_12439);
or U14170 (N_14170,N_12488,N_12447);
and U14171 (N_14171,N_12929,N_12183);
and U14172 (N_14172,N_12570,N_12706);
nand U14173 (N_14173,N_12122,N_13171);
nor U14174 (N_14174,N_12506,N_12642);
and U14175 (N_14175,N_13000,N_12713);
nand U14176 (N_14176,N_12112,N_12889);
nor U14177 (N_14177,N_12975,N_12148);
nor U14178 (N_14178,N_12908,N_13149);
nand U14179 (N_14179,N_12759,N_12378);
or U14180 (N_14180,N_12379,N_12544);
or U14181 (N_14181,N_12079,N_12236);
nand U14182 (N_14182,N_12173,N_12483);
and U14183 (N_14183,N_12506,N_13063);
nand U14184 (N_14184,N_12557,N_13050);
nor U14185 (N_14185,N_12990,N_12315);
nor U14186 (N_14186,N_12900,N_12704);
nor U14187 (N_14187,N_12225,N_12054);
and U14188 (N_14188,N_12672,N_12406);
xor U14189 (N_14189,N_12347,N_12186);
xor U14190 (N_14190,N_12870,N_12988);
nand U14191 (N_14191,N_13144,N_12131);
or U14192 (N_14192,N_12597,N_12627);
nor U14193 (N_14193,N_12490,N_12400);
or U14194 (N_14194,N_12944,N_12907);
nor U14195 (N_14195,N_12362,N_12813);
nor U14196 (N_14196,N_12694,N_12668);
and U14197 (N_14197,N_12962,N_13061);
xor U14198 (N_14198,N_12160,N_12292);
and U14199 (N_14199,N_12390,N_13037);
xnor U14200 (N_14200,N_13130,N_13020);
xnor U14201 (N_14201,N_12403,N_12196);
nand U14202 (N_14202,N_12975,N_12237);
nand U14203 (N_14203,N_12441,N_12065);
nor U14204 (N_14204,N_13063,N_12224);
xnor U14205 (N_14205,N_13025,N_13040);
xnor U14206 (N_14206,N_12374,N_13182);
nand U14207 (N_14207,N_12935,N_13104);
nor U14208 (N_14208,N_12007,N_12447);
or U14209 (N_14209,N_12004,N_12683);
nor U14210 (N_14210,N_12276,N_12853);
xor U14211 (N_14211,N_12889,N_12013);
nor U14212 (N_14212,N_12597,N_13126);
or U14213 (N_14213,N_12925,N_13114);
xnor U14214 (N_14214,N_12492,N_12783);
nand U14215 (N_14215,N_12895,N_12828);
and U14216 (N_14216,N_12007,N_12922);
or U14217 (N_14217,N_12465,N_12403);
nor U14218 (N_14218,N_13154,N_12352);
nor U14219 (N_14219,N_12339,N_12152);
xnor U14220 (N_14220,N_12683,N_12863);
or U14221 (N_14221,N_12126,N_12853);
xor U14222 (N_14222,N_12034,N_12680);
xor U14223 (N_14223,N_12586,N_12266);
or U14224 (N_14224,N_12665,N_12106);
and U14225 (N_14225,N_12323,N_12244);
nor U14226 (N_14226,N_12560,N_12512);
and U14227 (N_14227,N_12862,N_12710);
nand U14228 (N_14228,N_12114,N_12661);
nor U14229 (N_14229,N_12876,N_12004);
xnor U14230 (N_14230,N_12650,N_12809);
nand U14231 (N_14231,N_13179,N_13178);
and U14232 (N_14232,N_13089,N_12597);
and U14233 (N_14233,N_13040,N_12471);
nor U14234 (N_14234,N_12177,N_12474);
and U14235 (N_14235,N_13065,N_12721);
nand U14236 (N_14236,N_12887,N_12457);
nand U14237 (N_14237,N_12612,N_12087);
or U14238 (N_14238,N_12245,N_12507);
nor U14239 (N_14239,N_12262,N_12868);
or U14240 (N_14240,N_13079,N_12016);
and U14241 (N_14241,N_12072,N_12231);
nand U14242 (N_14242,N_12761,N_12338);
xnor U14243 (N_14243,N_12587,N_12428);
or U14244 (N_14244,N_12420,N_12728);
or U14245 (N_14245,N_12354,N_12026);
or U14246 (N_14246,N_13165,N_12511);
and U14247 (N_14247,N_12381,N_13110);
nand U14248 (N_14248,N_12501,N_12638);
or U14249 (N_14249,N_12639,N_13180);
and U14250 (N_14250,N_12435,N_12583);
nand U14251 (N_14251,N_12954,N_13046);
and U14252 (N_14252,N_12269,N_12259);
xnor U14253 (N_14253,N_12879,N_12675);
and U14254 (N_14254,N_12649,N_12246);
nand U14255 (N_14255,N_12456,N_12981);
or U14256 (N_14256,N_12787,N_13060);
xor U14257 (N_14257,N_12380,N_12761);
and U14258 (N_14258,N_12353,N_12448);
xor U14259 (N_14259,N_12953,N_13173);
nor U14260 (N_14260,N_13173,N_12902);
xor U14261 (N_14261,N_12707,N_12625);
xnor U14262 (N_14262,N_12950,N_13103);
nand U14263 (N_14263,N_13007,N_12441);
or U14264 (N_14264,N_12983,N_12968);
nand U14265 (N_14265,N_12773,N_12531);
xor U14266 (N_14266,N_12695,N_12531);
and U14267 (N_14267,N_13126,N_12421);
or U14268 (N_14268,N_12562,N_12863);
nand U14269 (N_14269,N_12627,N_13063);
or U14270 (N_14270,N_12926,N_12303);
and U14271 (N_14271,N_12030,N_12211);
or U14272 (N_14272,N_12719,N_13029);
xor U14273 (N_14273,N_13180,N_12999);
nor U14274 (N_14274,N_12017,N_12185);
and U14275 (N_14275,N_12030,N_13086);
or U14276 (N_14276,N_12679,N_12622);
nand U14277 (N_14277,N_12344,N_12816);
or U14278 (N_14278,N_12520,N_12302);
nor U14279 (N_14279,N_12448,N_12911);
xnor U14280 (N_14280,N_13028,N_13142);
nand U14281 (N_14281,N_12597,N_13162);
nor U14282 (N_14282,N_12206,N_12696);
xnor U14283 (N_14283,N_12250,N_12555);
xor U14284 (N_14284,N_13040,N_12435);
and U14285 (N_14285,N_12592,N_13073);
or U14286 (N_14286,N_12655,N_12038);
xnor U14287 (N_14287,N_12145,N_12195);
nor U14288 (N_14288,N_12319,N_12002);
nand U14289 (N_14289,N_12880,N_12035);
xnor U14290 (N_14290,N_12247,N_12300);
nand U14291 (N_14291,N_12856,N_12110);
nand U14292 (N_14292,N_12179,N_13051);
nand U14293 (N_14293,N_12005,N_12022);
nor U14294 (N_14294,N_12991,N_12584);
nor U14295 (N_14295,N_12544,N_12982);
nor U14296 (N_14296,N_12669,N_13138);
nor U14297 (N_14297,N_12427,N_12689);
nand U14298 (N_14298,N_12841,N_13152);
and U14299 (N_14299,N_12923,N_12418);
nand U14300 (N_14300,N_12487,N_12993);
nand U14301 (N_14301,N_12457,N_12448);
nand U14302 (N_14302,N_12687,N_12429);
nand U14303 (N_14303,N_12701,N_12803);
nor U14304 (N_14304,N_12283,N_12791);
or U14305 (N_14305,N_12772,N_12458);
and U14306 (N_14306,N_12175,N_12108);
or U14307 (N_14307,N_12910,N_12725);
nand U14308 (N_14308,N_13044,N_13172);
or U14309 (N_14309,N_12286,N_13117);
and U14310 (N_14310,N_12271,N_12285);
or U14311 (N_14311,N_12716,N_12459);
or U14312 (N_14312,N_12252,N_12594);
or U14313 (N_14313,N_12508,N_12718);
or U14314 (N_14314,N_12258,N_12327);
xnor U14315 (N_14315,N_12294,N_12402);
nand U14316 (N_14316,N_12079,N_12634);
xor U14317 (N_14317,N_12001,N_12011);
or U14318 (N_14318,N_12468,N_13000);
nand U14319 (N_14319,N_12879,N_12002);
or U14320 (N_14320,N_12477,N_12521);
or U14321 (N_14321,N_13008,N_12254);
nor U14322 (N_14322,N_12543,N_12324);
or U14323 (N_14323,N_12178,N_12385);
nor U14324 (N_14324,N_12250,N_12372);
nand U14325 (N_14325,N_12114,N_12382);
nor U14326 (N_14326,N_12979,N_12843);
xor U14327 (N_14327,N_12154,N_12630);
nor U14328 (N_14328,N_13183,N_12554);
xnor U14329 (N_14329,N_12860,N_12489);
xor U14330 (N_14330,N_12558,N_12072);
and U14331 (N_14331,N_12308,N_12181);
or U14332 (N_14332,N_12297,N_12477);
nand U14333 (N_14333,N_12216,N_12342);
and U14334 (N_14334,N_12024,N_12601);
nor U14335 (N_14335,N_12849,N_13054);
and U14336 (N_14336,N_13092,N_12616);
nand U14337 (N_14337,N_12244,N_12692);
xor U14338 (N_14338,N_13118,N_13081);
nor U14339 (N_14339,N_12666,N_12210);
xnor U14340 (N_14340,N_12514,N_12849);
nand U14341 (N_14341,N_12949,N_12156);
and U14342 (N_14342,N_12474,N_12446);
nand U14343 (N_14343,N_12590,N_12964);
xnor U14344 (N_14344,N_12706,N_12332);
xor U14345 (N_14345,N_13079,N_12073);
nor U14346 (N_14346,N_12792,N_12327);
nor U14347 (N_14347,N_12169,N_12351);
and U14348 (N_14348,N_12971,N_12772);
or U14349 (N_14349,N_12241,N_12832);
xor U14350 (N_14350,N_12177,N_12234);
or U14351 (N_14351,N_12274,N_13182);
xor U14352 (N_14352,N_12998,N_12102);
xnor U14353 (N_14353,N_12104,N_13143);
xnor U14354 (N_14354,N_12338,N_12584);
nand U14355 (N_14355,N_13076,N_12361);
or U14356 (N_14356,N_12182,N_12052);
and U14357 (N_14357,N_12609,N_12032);
xnor U14358 (N_14358,N_12075,N_12001);
nor U14359 (N_14359,N_13130,N_12550);
nand U14360 (N_14360,N_12405,N_12244);
or U14361 (N_14361,N_12901,N_12402);
or U14362 (N_14362,N_12381,N_12343);
xnor U14363 (N_14363,N_12186,N_12065);
or U14364 (N_14364,N_12834,N_12799);
nor U14365 (N_14365,N_12249,N_12698);
and U14366 (N_14366,N_12649,N_12016);
nor U14367 (N_14367,N_12456,N_12226);
nor U14368 (N_14368,N_12212,N_12613);
and U14369 (N_14369,N_12917,N_12464);
xnor U14370 (N_14370,N_12747,N_12056);
xnor U14371 (N_14371,N_12108,N_13013);
nand U14372 (N_14372,N_12830,N_12945);
or U14373 (N_14373,N_12663,N_12759);
or U14374 (N_14374,N_12291,N_13150);
and U14375 (N_14375,N_12557,N_12591);
xor U14376 (N_14376,N_12556,N_12693);
xor U14377 (N_14377,N_12762,N_12108);
nor U14378 (N_14378,N_12986,N_12865);
and U14379 (N_14379,N_12161,N_12368);
nor U14380 (N_14380,N_12941,N_12145);
and U14381 (N_14381,N_12259,N_12794);
and U14382 (N_14382,N_12288,N_12983);
xnor U14383 (N_14383,N_13012,N_12036);
and U14384 (N_14384,N_12211,N_12760);
and U14385 (N_14385,N_13142,N_12828);
or U14386 (N_14386,N_12696,N_12263);
xnor U14387 (N_14387,N_12042,N_12221);
nand U14388 (N_14388,N_13193,N_12363);
nor U14389 (N_14389,N_12712,N_12978);
nor U14390 (N_14390,N_12861,N_12534);
nand U14391 (N_14391,N_12467,N_12743);
and U14392 (N_14392,N_12075,N_12119);
and U14393 (N_14393,N_12994,N_12242);
nor U14394 (N_14394,N_12981,N_12722);
or U14395 (N_14395,N_12383,N_12920);
and U14396 (N_14396,N_13085,N_12738);
nor U14397 (N_14397,N_12650,N_12695);
xnor U14398 (N_14398,N_12488,N_13126);
nor U14399 (N_14399,N_12521,N_12872);
nand U14400 (N_14400,N_14363,N_13379);
nor U14401 (N_14401,N_13786,N_14147);
or U14402 (N_14402,N_14187,N_13833);
nand U14403 (N_14403,N_13599,N_14301);
or U14404 (N_14404,N_13522,N_14331);
nand U14405 (N_14405,N_14376,N_13257);
nor U14406 (N_14406,N_14359,N_14234);
nand U14407 (N_14407,N_14083,N_14032);
xor U14408 (N_14408,N_13751,N_13406);
and U14409 (N_14409,N_14045,N_13843);
xor U14410 (N_14410,N_13651,N_13377);
or U14411 (N_14411,N_13469,N_13866);
and U14412 (N_14412,N_13810,N_14153);
and U14413 (N_14413,N_14106,N_13357);
and U14414 (N_14414,N_13796,N_13606);
xor U14415 (N_14415,N_13999,N_14097);
nand U14416 (N_14416,N_13740,N_14102);
or U14417 (N_14417,N_13712,N_13551);
nor U14418 (N_14418,N_13316,N_14167);
nor U14419 (N_14419,N_13781,N_13491);
nor U14420 (N_14420,N_13263,N_14230);
nor U14421 (N_14421,N_13371,N_13545);
xor U14422 (N_14422,N_13749,N_13592);
or U14423 (N_14423,N_13729,N_13664);
or U14424 (N_14424,N_14249,N_13397);
nand U14425 (N_14425,N_13911,N_14180);
nand U14426 (N_14426,N_14202,N_13872);
nand U14427 (N_14427,N_13791,N_13957);
nor U14428 (N_14428,N_14367,N_13875);
nand U14429 (N_14429,N_13641,N_13658);
and U14430 (N_14430,N_13531,N_14362);
and U14431 (N_14431,N_14217,N_14341);
and U14432 (N_14432,N_13314,N_14148);
xor U14433 (N_14433,N_13992,N_13832);
and U14434 (N_14434,N_13201,N_13655);
xor U14435 (N_14435,N_13958,N_13619);
nor U14436 (N_14436,N_14282,N_13925);
or U14437 (N_14437,N_14195,N_13363);
nand U14438 (N_14438,N_13825,N_13777);
or U14439 (N_14439,N_13234,N_13460);
nand U14440 (N_14440,N_13952,N_13896);
nor U14441 (N_14441,N_13799,N_13972);
xnor U14442 (N_14442,N_13643,N_13628);
nor U14443 (N_14443,N_13723,N_13552);
and U14444 (N_14444,N_13950,N_13734);
xor U14445 (N_14445,N_13550,N_13744);
and U14446 (N_14446,N_13250,N_13984);
xor U14447 (N_14447,N_13722,N_13203);
nand U14448 (N_14448,N_13515,N_13648);
and U14449 (N_14449,N_13270,N_13555);
xor U14450 (N_14450,N_14251,N_13672);
and U14451 (N_14451,N_13738,N_13918);
nand U14452 (N_14452,N_13753,N_13627);
or U14453 (N_14453,N_13822,N_13939);
or U14454 (N_14454,N_14085,N_13216);
or U14455 (N_14455,N_14063,N_14242);
and U14456 (N_14456,N_13649,N_13811);
and U14457 (N_14457,N_14084,N_13407);
and U14458 (N_14458,N_13477,N_14399);
nand U14459 (N_14459,N_14350,N_13354);
xor U14460 (N_14460,N_13541,N_14009);
xnor U14461 (N_14461,N_13674,N_14235);
and U14462 (N_14462,N_14019,N_13755);
and U14463 (N_14463,N_13965,N_14328);
xnor U14464 (N_14464,N_14040,N_14314);
and U14465 (N_14465,N_13455,N_14015);
xor U14466 (N_14466,N_13494,N_14387);
nand U14467 (N_14467,N_14238,N_14243);
nand U14468 (N_14468,N_13528,N_13580);
nand U14469 (N_14469,N_13910,N_13352);
nor U14470 (N_14470,N_14017,N_13700);
or U14471 (N_14471,N_13675,N_14397);
xor U14472 (N_14472,N_14349,N_13300);
nor U14473 (N_14473,N_13986,N_13699);
nor U14474 (N_14474,N_13548,N_13891);
xor U14475 (N_14475,N_13881,N_13233);
and U14476 (N_14476,N_13978,N_13766);
and U14477 (N_14477,N_14056,N_13959);
nor U14478 (N_14478,N_13403,N_13835);
or U14479 (N_14479,N_13677,N_14246);
nand U14480 (N_14480,N_13828,N_13594);
and U14481 (N_14481,N_14355,N_13304);
nand U14482 (N_14482,N_14393,N_14309);
or U14483 (N_14483,N_14211,N_13899);
or U14484 (N_14484,N_14285,N_13947);
and U14485 (N_14485,N_14356,N_14154);
nand U14486 (N_14486,N_13364,N_13758);
nand U14487 (N_14487,N_14104,N_14183);
nor U14488 (N_14488,N_14351,N_13754);
and U14489 (N_14489,N_13794,N_13517);
nor U14490 (N_14490,N_14173,N_13435);
or U14491 (N_14491,N_14182,N_13598);
xor U14492 (N_14492,N_13297,N_13861);
nand U14493 (N_14493,N_14171,N_14123);
nand U14494 (N_14494,N_13680,N_13622);
or U14495 (N_14495,N_13577,N_13562);
or U14496 (N_14496,N_14291,N_13306);
xnor U14497 (N_14497,N_13490,N_14346);
or U14498 (N_14498,N_14231,N_13706);
nor U14499 (N_14499,N_13211,N_14277);
xor U14500 (N_14500,N_13808,N_14087);
nand U14501 (N_14501,N_13801,N_14368);
nand U14502 (N_14502,N_14093,N_14257);
and U14503 (N_14503,N_14004,N_14262);
nand U14504 (N_14504,N_13390,N_13426);
xnor U14505 (N_14505,N_13227,N_14361);
and U14506 (N_14506,N_13804,N_13298);
xor U14507 (N_14507,N_13995,N_13800);
xnor U14508 (N_14508,N_13520,N_14013);
or U14509 (N_14509,N_14227,N_13805);
nor U14510 (N_14510,N_14021,N_13879);
or U14511 (N_14511,N_14320,N_13450);
and U14512 (N_14512,N_13242,N_13559);
xor U14513 (N_14513,N_13208,N_13750);
and U14514 (N_14514,N_13525,N_13567);
or U14515 (N_14515,N_13478,N_13793);
or U14516 (N_14516,N_13660,N_13955);
and U14517 (N_14517,N_14033,N_13220);
nand U14518 (N_14518,N_13798,N_13235);
xor U14519 (N_14519,N_13831,N_13855);
nand U14520 (N_14520,N_14364,N_13812);
nor U14521 (N_14521,N_14108,N_14354);
xor U14522 (N_14522,N_13707,N_13232);
and U14523 (N_14523,N_14221,N_14181);
nand U14524 (N_14524,N_14245,N_14207);
and U14525 (N_14525,N_13569,N_13282);
nand U14526 (N_14526,N_13412,N_14103);
or U14527 (N_14527,N_14233,N_13295);
xor U14528 (N_14528,N_13617,N_14116);
nand U14529 (N_14529,N_13761,N_13637);
nor U14530 (N_14530,N_13888,N_13358);
or U14531 (N_14531,N_14290,N_14155);
xnor U14532 (N_14532,N_13558,N_13310);
nand U14533 (N_14533,N_13671,N_14261);
nand U14534 (N_14534,N_13634,N_14258);
and U14535 (N_14535,N_13446,N_13966);
nand U14536 (N_14536,N_13587,N_13591);
nand U14537 (N_14537,N_13605,N_13432);
or U14538 (N_14538,N_14105,N_13482);
xor U14539 (N_14539,N_14090,N_13311);
xnor U14540 (N_14540,N_14111,N_13968);
nor U14541 (N_14541,N_13876,N_14037);
xor U14542 (N_14542,N_13313,N_14191);
xnor U14543 (N_14543,N_13654,N_13682);
xor U14544 (N_14544,N_13329,N_14272);
xnor U14545 (N_14545,N_13852,N_13933);
nor U14546 (N_14546,N_13401,N_14115);
nor U14547 (N_14547,N_13378,N_13676);
xnor U14548 (N_14548,N_14053,N_13607);
xnor U14549 (N_14549,N_13542,N_13644);
nor U14550 (N_14550,N_13868,N_13907);
nor U14551 (N_14551,N_13759,N_13409);
xor U14552 (N_14552,N_13302,N_14292);
or U14553 (N_14553,N_14172,N_14337);
nor U14554 (N_14554,N_14018,N_14135);
and U14555 (N_14555,N_14190,N_14216);
and U14556 (N_14556,N_13206,N_13414);
nand U14557 (N_14557,N_13813,N_14080);
or U14558 (N_14558,N_13327,N_13915);
nor U14559 (N_14559,N_14160,N_13365);
xnor U14560 (N_14560,N_14288,N_13716);
nor U14561 (N_14561,N_13554,N_13987);
nor U14562 (N_14562,N_14132,N_13486);
xor U14563 (N_14563,N_13578,N_13384);
and U14564 (N_14564,N_14138,N_13244);
and U14565 (N_14565,N_13683,N_14162);
and U14566 (N_14566,N_14247,N_13402);
nand U14567 (N_14567,N_14066,N_13274);
nand U14568 (N_14568,N_13315,N_14120);
nand U14569 (N_14569,N_14332,N_13499);
nand U14570 (N_14570,N_13974,N_13889);
nor U14571 (N_14571,N_13685,N_13293);
and U14572 (N_14572,N_14122,N_14305);
xnor U14573 (N_14573,N_13924,N_13823);
nor U14574 (N_14574,N_14077,N_13860);
or U14575 (N_14575,N_14145,N_14031);
and U14576 (N_14576,N_13757,N_14220);
and U14577 (N_14577,N_14330,N_13226);
or U14578 (N_14578,N_14300,N_14163);
or U14579 (N_14579,N_14025,N_14078);
or U14580 (N_14580,N_14137,N_13770);
and U14581 (N_14581,N_13348,N_13814);
and U14582 (N_14582,N_14392,N_13882);
nand U14583 (N_14583,N_13816,N_13321);
or U14584 (N_14584,N_14223,N_14131);
nand U14585 (N_14585,N_14192,N_13589);
or U14586 (N_14586,N_13684,N_14002);
and U14587 (N_14587,N_14201,N_13366);
nor U14588 (N_14588,N_14127,N_13593);
xnor U14589 (N_14589,N_14199,N_13439);
or U14590 (N_14590,N_13838,N_13726);
and U14591 (N_14591,N_13498,N_13693);
and U14592 (N_14592,N_14304,N_14067);
xor U14593 (N_14593,N_13615,N_13527);
xor U14594 (N_14594,N_13779,N_13850);
and U14595 (N_14595,N_14189,N_14005);
nor U14596 (N_14596,N_13919,N_13696);
nor U14597 (N_14597,N_14307,N_13420);
and U14598 (N_14598,N_13787,N_13495);
or U14599 (N_14599,N_14073,N_13846);
and U14600 (N_14600,N_14194,N_13989);
or U14601 (N_14601,N_13458,N_13291);
nand U14602 (N_14602,N_13454,N_13936);
nor U14603 (N_14603,N_13294,N_13837);
or U14604 (N_14604,N_13285,N_13510);
nor U14605 (N_14605,N_13916,N_14094);
or U14606 (N_14606,N_13570,N_13466);
or U14607 (N_14607,N_13626,N_13353);
nand U14608 (N_14608,N_13465,N_14310);
nor U14609 (N_14609,N_13610,N_13624);
and U14610 (N_14610,N_13438,N_13507);
or U14611 (N_14611,N_13476,N_13265);
xnor U14612 (N_14612,N_13202,N_14365);
or U14613 (N_14613,N_13386,N_13488);
nor U14614 (N_14614,N_14353,N_13909);
xnor U14615 (N_14615,N_14286,N_13241);
or U14616 (N_14616,N_13803,N_13767);
xnor U14617 (N_14617,N_13737,N_13739);
and U14618 (N_14618,N_13385,N_14164);
or U14619 (N_14619,N_14283,N_13728);
xor U14620 (N_14620,N_13940,N_14074);
and U14621 (N_14621,N_13322,N_13708);
nor U14622 (N_14622,N_14264,N_13782);
nor U14623 (N_14623,N_13920,N_13368);
and U14624 (N_14624,N_14139,N_14333);
nand U14625 (N_14625,N_14370,N_13701);
nor U14626 (N_14626,N_14001,N_13271);
or U14627 (N_14627,N_13411,N_13632);
and U14628 (N_14628,N_14335,N_14060);
and U14629 (N_14629,N_13393,N_14188);
or U14630 (N_14630,N_14280,N_13376);
nand U14631 (N_14631,N_14284,N_13848);
and U14632 (N_14632,N_14026,N_13746);
or U14633 (N_14633,N_13457,N_13513);
and U14634 (N_14634,N_14043,N_13917);
and U14635 (N_14635,N_14270,N_13451);
nor U14636 (N_14636,N_13893,N_14089);
and U14637 (N_14637,N_13720,N_13425);
nor U14638 (N_14638,N_14237,N_14208);
nor U14639 (N_14639,N_13663,N_13337);
and U14640 (N_14640,N_13429,N_13511);
nor U14641 (N_14641,N_14050,N_13679);
nand U14642 (N_14642,N_14383,N_13388);
and U14643 (N_14643,N_14347,N_14395);
and U14644 (N_14644,N_13897,N_14222);
xor U14645 (N_14645,N_13288,N_13949);
xnor U14646 (N_14646,N_13871,N_13341);
nor U14647 (N_14647,N_13922,N_13576);
nand U14648 (N_14648,N_13927,N_13504);
xnor U14649 (N_14649,N_13557,N_13921);
nor U14650 (N_14650,N_13309,N_13844);
nand U14651 (N_14651,N_13666,N_13264);
and U14652 (N_14652,N_13903,N_13873);
or U14653 (N_14653,N_14197,N_13284);
and U14654 (N_14654,N_13988,N_13566);
or U14655 (N_14655,N_13883,N_14338);
or U14656 (N_14656,N_13229,N_13497);
or U14657 (N_14657,N_13400,N_14006);
or U14658 (N_14658,N_13745,N_13383);
and U14659 (N_14659,N_14256,N_14129);
or U14660 (N_14660,N_13923,N_13396);
xnor U14661 (N_14661,N_14276,N_14027);
xnor U14662 (N_14662,N_13941,N_13748);
nor U14663 (N_14663,N_13392,N_14130);
nor U14664 (N_14664,N_13931,N_14390);
or U14665 (N_14665,N_13862,N_14144);
xnor U14666 (N_14666,N_14156,N_14193);
xor U14667 (N_14667,N_13456,N_13629);
and U14668 (N_14668,N_13526,N_13713);
and U14669 (N_14669,N_13360,N_13642);
nand U14670 (N_14670,N_13845,N_13289);
xor U14671 (N_14671,N_13980,N_13690);
xor U14672 (N_14672,N_14254,N_14098);
xnor U14673 (N_14673,N_14380,N_13904);
nand U14674 (N_14674,N_13913,N_14339);
nand U14675 (N_14675,N_13572,N_13342);
and U14676 (N_14676,N_13638,N_13665);
nor U14677 (N_14677,N_13568,N_13752);
nand U14678 (N_14678,N_13418,N_14125);
nand U14679 (N_14679,N_14295,N_13858);
and U14680 (N_14680,N_13765,N_14329);
nor U14681 (N_14681,N_14252,N_14287);
or U14682 (N_14682,N_13280,N_13584);
nor U14683 (N_14683,N_14134,N_13431);
xor U14684 (N_14684,N_14378,N_13333);
or U14685 (N_14685,N_13514,N_14228);
or U14686 (N_14686,N_14323,N_13829);
nand U14687 (N_14687,N_14279,N_13727);
or U14688 (N_14688,N_14313,N_13374);
or U14689 (N_14689,N_13243,N_13709);
and U14690 (N_14690,N_14034,N_13278);
nand U14691 (N_14691,N_14054,N_13417);
xnor U14692 (N_14692,N_13474,N_14340);
nand U14693 (N_14693,N_13900,N_14205);
or U14694 (N_14694,N_13603,N_13317);
nand U14695 (N_14695,N_13251,N_14336);
or U14696 (N_14696,N_13290,N_14113);
xnor U14697 (N_14697,N_13287,N_13970);
or U14698 (N_14698,N_13973,N_13349);
nand U14699 (N_14699,N_13356,N_14269);
xor U14700 (N_14700,N_13259,N_13967);
xor U14701 (N_14701,N_14236,N_13339);
and U14702 (N_14702,N_14079,N_14316);
or U14703 (N_14703,N_13611,N_13681);
xor U14704 (N_14704,N_13733,N_14263);
xor U14705 (N_14705,N_14255,N_14379);
and U14706 (N_14706,N_13224,N_14174);
nor U14707 (N_14707,N_14371,N_13631);
and U14708 (N_14708,N_14259,N_14149);
nand U14709 (N_14709,N_13275,N_14142);
nor U14710 (N_14710,N_13362,N_13864);
nor U14711 (N_14711,N_13273,N_13998);
nand U14712 (N_14712,N_14109,N_14170);
or U14713 (N_14713,N_13616,N_14049);
nand U14714 (N_14714,N_13387,N_13332);
and U14715 (N_14715,N_14317,N_13442);
and U14716 (N_14716,N_13826,N_13225);
nor U14717 (N_14717,N_13743,N_13908);
or U14718 (N_14718,N_13532,N_13207);
or U14719 (N_14719,N_13492,N_13635);
and U14720 (N_14720,N_13934,N_14360);
or U14721 (N_14721,N_13990,N_13540);
nand U14722 (N_14722,N_13874,N_14274);
and U14723 (N_14723,N_14297,N_13625);
and U14724 (N_14724,N_14126,N_14096);
xnor U14725 (N_14725,N_14152,N_13785);
xnor U14726 (N_14726,N_13715,N_13239);
nand U14727 (N_14727,N_14051,N_14334);
and U14728 (N_14728,N_14303,N_14326);
or U14729 (N_14729,N_14267,N_13350);
and U14730 (N_14730,N_13869,N_13428);
and U14731 (N_14731,N_13653,N_14151);
nor U14732 (N_14732,N_13512,N_13954);
xor U14733 (N_14733,N_13338,N_14299);
nor U14734 (N_14734,N_14281,N_13659);
xnor U14735 (N_14735,N_13276,N_13730);
or U14736 (N_14736,N_14091,N_14022);
xnor U14737 (N_14737,N_13444,N_13943);
xor U14738 (N_14738,N_13763,N_13717);
xor U14739 (N_14739,N_14374,N_13324);
nor U14740 (N_14740,N_14011,N_13612);
nor U14741 (N_14741,N_13501,N_13355);
or U14742 (N_14742,N_13292,N_13867);
xor U14743 (N_14743,N_13481,N_13347);
nand U14744 (N_14744,N_13565,N_14064);
or U14745 (N_14745,N_13668,N_14225);
xnor U14746 (N_14746,N_13771,N_13391);
or U14747 (N_14747,N_13820,N_14384);
or U14748 (N_14748,N_13212,N_14119);
nand U14749 (N_14749,N_13521,N_14061);
xnor U14750 (N_14750,N_14213,N_13691);
or U14751 (N_14751,N_14082,N_13415);
or U14752 (N_14752,N_13650,N_13518);
nand U14753 (N_14753,N_14253,N_14020);
xnor U14754 (N_14754,N_14377,N_14101);
or U14755 (N_14755,N_13381,N_13807);
or U14756 (N_14756,N_14124,N_14322);
nor U14757 (N_14757,N_13404,N_13573);
nand U14758 (N_14758,N_14128,N_14358);
and U14759 (N_14759,N_14095,N_13213);
xor U14760 (N_14760,N_13533,N_13878);
and U14761 (N_14761,N_14318,N_13496);
and U14762 (N_14762,N_13307,N_13236);
xor U14763 (N_14763,N_14143,N_14327);
and U14764 (N_14764,N_13788,N_13249);
xnor U14765 (N_14765,N_13574,N_13600);
and U14766 (N_14766,N_13932,N_13299);
xnor U14767 (N_14767,N_13710,N_13319);
nand U14768 (N_14768,N_14168,N_13703);
or U14769 (N_14769,N_13623,N_13993);
xnor U14770 (N_14770,N_13898,N_13686);
or U14771 (N_14771,N_13859,N_13543);
nor U14772 (N_14772,N_14052,N_13702);
or U14773 (N_14773,N_13238,N_14212);
and U14774 (N_14774,N_14150,N_13945);
xnor U14775 (N_14775,N_13842,N_13372);
and U14776 (N_14776,N_13468,N_13246);
nor U14777 (N_14777,N_13480,N_14315);
and U14778 (N_14778,N_13847,N_14041);
nor U14779 (N_14779,N_13613,N_13789);
or U14780 (N_14780,N_13325,N_14012);
and U14781 (N_14781,N_14271,N_14112);
or U14782 (N_14782,N_13991,N_14298);
nor U14783 (N_14783,N_14176,N_14344);
nand U14784 (N_14784,N_13942,N_13473);
nor U14785 (N_14785,N_14239,N_13818);
or U14786 (N_14786,N_13410,N_13389);
and U14787 (N_14787,N_13221,N_13215);
nor U14788 (N_14788,N_13547,N_14008);
and U14789 (N_14789,N_13445,N_13588);
and U14790 (N_14790,N_13538,N_13575);
nand U14791 (N_14791,N_13776,N_14306);
nor U14792 (N_14792,N_13985,N_13463);
xor U14793 (N_14793,N_14366,N_14047);
nand U14794 (N_14794,N_14058,N_14215);
and U14795 (N_14795,N_13618,N_13975);
nor U14796 (N_14796,N_13851,N_13506);
nor U14797 (N_14797,N_13802,N_14324);
nor U14798 (N_14798,N_14141,N_13840);
xor U14799 (N_14799,N_14072,N_14042);
nand U14800 (N_14800,N_13887,N_13930);
and U14801 (N_14801,N_13824,N_14169);
or U14802 (N_14802,N_13539,N_13886);
or U14803 (N_14803,N_13783,N_14014);
or U14804 (N_14804,N_14140,N_13398);
and U14805 (N_14805,N_13351,N_14117);
and U14806 (N_14806,N_14248,N_14110);
xor U14807 (N_14807,N_13537,N_13760);
xor U14808 (N_14808,N_14293,N_13424);
nand U14809 (N_14809,N_13633,N_14224);
and U14810 (N_14810,N_13849,N_13231);
or U14811 (N_14811,N_13583,N_14203);
or U14812 (N_14812,N_13951,N_14055);
and U14813 (N_14813,N_13335,N_13260);
xor U14814 (N_14814,N_13453,N_14178);
nor U14815 (N_14815,N_13268,N_14396);
and U14816 (N_14816,N_13948,N_13399);
and U14817 (N_14817,N_13792,N_13560);
xnor U14818 (N_14818,N_13301,N_13373);
xnor U14819 (N_14819,N_14068,N_14226);
nand U14820 (N_14820,N_14294,N_14059);
xor U14821 (N_14821,N_13914,N_13596);
nand U14822 (N_14822,N_14044,N_13895);
xnor U14823 (N_14823,N_13636,N_13331);
nor U14824 (N_14824,N_13217,N_14038);
nand U14825 (N_14825,N_13544,N_13773);
nand U14826 (N_14826,N_13762,N_14302);
and U14827 (N_14827,N_13697,N_13926);
or U14828 (N_14828,N_13894,N_13556);
and U14829 (N_14829,N_13604,N_13440);
or U14830 (N_14830,N_13956,N_13326);
xor U14831 (N_14831,N_13963,N_13819);
and U14832 (N_14832,N_13340,N_13549);
or U14833 (N_14833,N_14311,N_13841);
nor U14834 (N_14834,N_14348,N_13345);
xor U14835 (N_14835,N_13582,N_14107);
and U14836 (N_14836,N_13509,N_13983);
or U14837 (N_14837,N_13487,N_14289);
xnor U14838 (N_14838,N_14388,N_13994);
nand U14839 (N_14839,N_13443,N_13369);
and U14840 (N_14840,N_14136,N_13901);
nand U14841 (N_14841,N_13405,N_14200);
nand U14842 (N_14842,N_13736,N_14030);
or U14843 (N_14843,N_13662,N_14065);
or U14844 (N_14844,N_14133,N_13772);
xor U14845 (N_14845,N_13483,N_13964);
or U14846 (N_14846,N_13380,N_14081);
or U14847 (N_14847,N_14069,N_13254);
xnor U14848 (N_14848,N_13747,N_13422);
xnor U14849 (N_14849,N_13470,N_13602);
nor U14850 (N_14850,N_13778,N_13553);
nor U14851 (N_14851,N_14177,N_13269);
xnor U14852 (N_14852,N_13283,N_13437);
nor U14853 (N_14853,N_13630,N_14057);
nand U14854 (N_14854,N_13485,N_13503);
nor U14855 (N_14855,N_14159,N_13563);
or U14856 (N_14856,N_14024,N_13652);
xnor U14857 (N_14857,N_13856,N_14389);
or U14858 (N_14858,N_13361,N_13732);
or U14859 (N_14859,N_13689,N_13795);
or U14860 (N_14860,N_13323,N_13529);
and U14861 (N_14861,N_13769,N_13305);
and U14862 (N_14862,N_14232,N_13645);
or U14863 (N_14863,N_13976,N_13997);
nand U14864 (N_14864,N_14121,N_14325);
or U14865 (N_14865,N_13971,N_14088);
nand U14866 (N_14866,N_13996,N_13524);
xnor U14867 (N_14867,N_14244,N_14265);
xnor U14868 (N_14868,N_13977,N_13590);
xnor U14869 (N_14869,N_13597,N_13657);
nand U14870 (N_14870,N_13741,N_14118);
and U14871 (N_14871,N_13870,N_14369);
nor U14872 (N_14872,N_13230,N_13240);
nand U14873 (N_14873,N_13523,N_14273);
xnor U14874 (N_14874,N_14092,N_13834);
nand U14875 (N_14875,N_13982,N_13367);
nor U14876 (N_14876,N_14373,N_13564);
nand U14877 (N_14877,N_14023,N_13464);
nor U14878 (N_14878,N_13906,N_14296);
xor U14879 (N_14879,N_13436,N_13218);
xor U14880 (N_14880,N_14029,N_13489);
xor U14881 (N_14881,N_13375,N_14075);
nor U14882 (N_14882,N_14039,N_13938);
nor U14883 (N_14883,N_13678,N_14275);
nor U14884 (N_14884,N_14186,N_13764);
xnor U14885 (N_14885,N_13768,N_13209);
nand U14886 (N_14886,N_13423,N_13286);
or U14887 (N_14887,N_14099,N_13912);
nor U14888 (N_14888,N_13695,N_13817);
xor U14889 (N_14889,N_14210,N_13960);
nor U14890 (N_14890,N_13979,N_13711);
nand U14891 (N_14891,N_14385,N_14357);
and U14892 (N_14892,N_13595,N_13687);
or U14893 (N_14893,N_13459,N_14398);
or U14894 (N_14894,N_13719,N_14278);
or U14895 (N_14895,N_13530,N_13416);
or U14896 (N_14896,N_13266,N_14260);
and U14897 (N_14897,N_13614,N_13827);
xor U14898 (N_14898,N_13705,N_13929);
or U14899 (N_14899,N_13585,N_13780);
nor U14900 (N_14900,N_14007,N_13214);
or U14901 (N_14901,N_13673,N_13318);
nor U14902 (N_14902,N_14372,N_14241);
nor U14903 (N_14903,N_14382,N_13784);
or U14904 (N_14904,N_14048,N_13320);
nor U14905 (N_14905,N_13237,N_13735);
xnor U14906 (N_14906,N_13219,N_13502);
xor U14907 (N_14907,N_13359,N_13704);
xnor U14908 (N_14908,N_14198,N_13640);
xnor U14909 (N_14909,N_14219,N_14100);
xnor U14910 (N_14910,N_13601,N_13467);
nor U14911 (N_14911,N_13493,N_13981);
and U14912 (N_14912,N_13935,N_13336);
nand U14913 (N_14913,N_13255,N_14268);
nand U14914 (N_14914,N_13370,N_13534);
nor U14915 (N_14915,N_13519,N_13484);
or U14916 (N_14916,N_13944,N_13639);
and U14917 (N_14917,N_14161,N_13775);
nor U14918 (N_14918,N_14204,N_13721);
nand U14919 (N_14919,N_13449,N_14266);
and U14920 (N_14920,N_13247,N_13296);
nand U14921 (N_14921,N_14342,N_13688);
nand U14922 (N_14922,N_13756,N_13500);
and U14923 (N_14923,N_13885,N_13228);
and U14924 (N_14924,N_13774,N_13821);
nand U14925 (N_14925,N_13839,N_13854);
or U14926 (N_14926,N_13253,N_13252);
or U14927 (N_14927,N_14196,N_13334);
nand U14928 (N_14928,N_14000,N_13742);
nand U14929 (N_14929,N_13646,N_13508);
nor U14930 (N_14930,N_13905,N_14076);
xor U14931 (N_14931,N_13877,N_14386);
and U14932 (N_14932,N_13937,N_14214);
and U14933 (N_14933,N_13647,N_13395);
and U14934 (N_14934,N_13961,N_13441);
nand U14935 (N_14935,N_13863,N_14343);
or U14936 (N_14936,N_13731,N_13694);
xnor U14937 (N_14937,N_13797,N_13448);
and U14938 (N_14938,N_13890,N_13670);
and U14939 (N_14939,N_13516,N_13656);
or U14940 (N_14940,N_13581,N_13427);
nor U14941 (N_14941,N_13725,N_13258);
or U14942 (N_14942,N_14184,N_13222);
xnor U14943 (N_14943,N_14158,N_13579);
xnor U14944 (N_14944,N_13256,N_13267);
nor U14945 (N_14945,N_13586,N_13281);
nand U14946 (N_14946,N_14028,N_14352);
nor U14947 (N_14947,N_13308,N_13471);
nand U14948 (N_14948,N_13262,N_13880);
nor U14949 (N_14949,N_13892,N_14010);
and U14950 (N_14950,N_14179,N_14229);
nand U14951 (N_14951,N_13853,N_13447);
nand U14952 (N_14952,N_13561,N_13479);
xnor U14953 (N_14953,N_13698,N_13245);
xor U14954 (N_14954,N_13223,N_14157);
and U14955 (N_14955,N_13692,N_13928);
or U14956 (N_14956,N_13248,N_13535);
xnor U14957 (N_14957,N_13620,N_13472);
or U14958 (N_14958,N_14175,N_13204);
xor U14959 (N_14959,N_14206,N_13382);
and U14960 (N_14960,N_14070,N_13836);
nor U14961 (N_14961,N_13434,N_13884);
nand U14962 (N_14962,N_13461,N_14381);
nor U14963 (N_14963,N_13303,N_13546);
xnor U14964 (N_14964,N_13857,N_13865);
nor U14965 (N_14965,N_13343,N_13346);
nor U14966 (N_14966,N_13790,N_13205);
xnor U14967 (N_14967,N_13609,N_13969);
nand U14968 (N_14968,N_14308,N_13953);
xor U14969 (N_14969,N_14035,N_13505);
or U14970 (N_14970,N_13608,N_13419);
and U14971 (N_14971,N_14071,N_13830);
nand U14972 (N_14972,N_13430,N_13330);
or U14973 (N_14973,N_13806,N_14209);
or U14974 (N_14974,N_14319,N_13536);
and U14975 (N_14975,N_14185,N_14166);
or U14976 (N_14976,N_13815,N_13452);
nor U14977 (N_14977,N_13344,N_13661);
xor U14978 (N_14978,N_14375,N_14114);
xnor U14979 (N_14979,N_14394,N_14321);
nand U14980 (N_14980,N_13279,N_14016);
or U14981 (N_14981,N_13394,N_13669);
xor U14982 (N_14982,N_13200,N_13261);
and U14983 (N_14983,N_13714,N_14312);
nor U14984 (N_14984,N_14036,N_13312);
or U14985 (N_14985,N_13433,N_14240);
nand U14986 (N_14986,N_14345,N_14086);
nand U14987 (N_14987,N_14165,N_13962);
nor U14988 (N_14988,N_14062,N_13462);
or U14989 (N_14989,N_13621,N_13421);
nand U14990 (N_14990,N_13667,N_14391);
and U14991 (N_14991,N_13724,N_13571);
nand U14992 (N_14992,N_14003,N_14146);
or U14993 (N_14993,N_13902,N_13408);
or U14994 (N_14994,N_13413,N_14218);
nand U14995 (N_14995,N_13210,N_13475);
and U14996 (N_14996,N_14250,N_13328);
and U14997 (N_14997,N_13272,N_13718);
nand U14998 (N_14998,N_14046,N_13277);
nor U14999 (N_14999,N_13809,N_13946);
and U15000 (N_15000,N_14290,N_14007);
nand U15001 (N_15001,N_13271,N_14234);
nand U15002 (N_15002,N_14072,N_13556);
or U15003 (N_15003,N_13895,N_13592);
xor U15004 (N_15004,N_14030,N_14278);
nand U15005 (N_15005,N_14307,N_13659);
and U15006 (N_15006,N_13805,N_13317);
or U15007 (N_15007,N_13960,N_13520);
and U15008 (N_15008,N_13398,N_13822);
nand U15009 (N_15009,N_14239,N_14105);
nor U15010 (N_15010,N_13740,N_13922);
nor U15011 (N_15011,N_14171,N_14117);
and U15012 (N_15012,N_13545,N_14201);
and U15013 (N_15013,N_13722,N_14129);
xnor U15014 (N_15014,N_13954,N_14172);
nor U15015 (N_15015,N_13486,N_14399);
and U15016 (N_15016,N_14118,N_13972);
and U15017 (N_15017,N_13882,N_14131);
nand U15018 (N_15018,N_14246,N_13572);
nand U15019 (N_15019,N_14222,N_14321);
xnor U15020 (N_15020,N_14302,N_13824);
and U15021 (N_15021,N_13869,N_13947);
or U15022 (N_15022,N_13316,N_14020);
and U15023 (N_15023,N_13493,N_14077);
nor U15024 (N_15024,N_13434,N_14057);
or U15025 (N_15025,N_14251,N_13493);
or U15026 (N_15026,N_14383,N_13268);
nand U15027 (N_15027,N_14297,N_14278);
and U15028 (N_15028,N_14219,N_14344);
or U15029 (N_15029,N_13727,N_14293);
or U15030 (N_15030,N_13840,N_13876);
xor U15031 (N_15031,N_14096,N_14081);
nand U15032 (N_15032,N_13768,N_14018);
or U15033 (N_15033,N_13588,N_13209);
xnor U15034 (N_15034,N_13863,N_14035);
nand U15035 (N_15035,N_13826,N_14009);
and U15036 (N_15036,N_14176,N_14098);
or U15037 (N_15037,N_13855,N_13430);
or U15038 (N_15038,N_14308,N_13792);
or U15039 (N_15039,N_13960,N_13659);
and U15040 (N_15040,N_13215,N_13256);
xnor U15041 (N_15041,N_13515,N_13998);
nand U15042 (N_15042,N_14325,N_13660);
or U15043 (N_15043,N_13962,N_13547);
nand U15044 (N_15044,N_13971,N_14099);
or U15045 (N_15045,N_13295,N_13282);
and U15046 (N_15046,N_13606,N_13437);
or U15047 (N_15047,N_13212,N_13572);
or U15048 (N_15048,N_13863,N_14366);
xor U15049 (N_15049,N_13717,N_14198);
and U15050 (N_15050,N_13817,N_14109);
or U15051 (N_15051,N_13888,N_13740);
nand U15052 (N_15052,N_13869,N_13835);
nor U15053 (N_15053,N_14315,N_13787);
and U15054 (N_15054,N_13577,N_13404);
nand U15055 (N_15055,N_13390,N_13634);
nand U15056 (N_15056,N_13682,N_14256);
nor U15057 (N_15057,N_13686,N_13226);
and U15058 (N_15058,N_13750,N_14374);
or U15059 (N_15059,N_13564,N_14136);
or U15060 (N_15060,N_14024,N_13598);
nand U15061 (N_15061,N_13927,N_13585);
nand U15062 (N_15062,N_13547,N_13599);
nor U15063 (N_15063,N_13953,N_13414);
nand U15064 (N_15064,N_13899,N_14086);
and U15065 (N_15065,N_13926,N_13258);
xnor U15066 (N_15066,N_13892,N_13780);
nor U15067 (N_15067,N_13864,N_14300);
and U15068 (N_15068,N_13421,N_13740);
xnor U15069 (N_15069,N_13663,N_13908);
or U15070 (N_15070,N_14245,N_13546);
nor U15071 (N_15071,N_14102,N_14030);
and U15072 (N_15072,N_14111,N_13372);
nor U15073 (N_15073,N_14203,N_14316);
xor U15074 (N_15074,N_14238,N_13319);
nand U15075 (N_15075,N_13200,N_13606);
nor U15076 (N_15076,N_13871,N_13667);
nor U15077 (N_15077,N_14106,N_13637);
or U15078 (N_15078,N_13232,N_13317);
nand U15079 (N_15079,N_13437,N_13465);
and U15080 (N_15080,N_14312,N_14087);
and U15081 (N_15081,N_13542,N_14298);
xor U15082 (N_15082,N_13562,N_14230);
nor U15083 (N_15083,N_13648,N_13756);
nor U15084 (N_15084,N_13201,N_13200);
or U15085 (N_15085,N_14091,N_13254);
and U15086 (N_15086,N_13558,N_14361);
or U15087 (N_15087,N_13348,N_14291);
nand U15088 (N_15088,N_14380,N_14056);
and U15089 (N_15089,N_13319,N_13749);
and U15090 (N_15090,N_13559,N_14287);
and U15091 (N_15091,N_13492,N_13453);
and U15092 (N_15092,N_13835,N_13206);
and U15093 (N_15093,N_14111,N_13318);
nor U15094 (N_15094,N_13472,N_13939);
xor U15095 (N_15095,N_13442,N_14086);
and U15096 (N_15096,N_13829,N_14183);
nor U15097 (N_15097,N_14047,N_13264);
and U15098 (N_15098,N_13578,N_14007);
and U15099 (N_15099,N_13306,N_13236);
nand U15100 (N_15100,N_13940,N_13298);
and U15101 (N_15101,N_14228,N_14274);
or U15102 (N_15102,N_14282,N_13715);
xnor U15103 (N_15103,N_14308,N_13622);
or U15104 (N_15104,N_13459,N_13991);
nand U15105 (N_15105,N_14002,N_14104);
or U15106 (N_15106,N_13308,N_13916);
or U15107 (N_15107,N_14130,N_14371);
or U15108 (N_15108,N_14269,N_13362);
and U15109 (N_15109,N_14199,N_13831);
and U15110 (N_15110,N_13879,N_13973);
xor U15111 (N_15111,N_13665,N_14374);
xor U15112 (N_15112,N_13839,N_13315);
nor U15113 (N_15113,N_13735,N_13338);
xnor U15114 (N_15114,N_14185,N_13998);
and U15115 (N_15115,N_14023,N_14084);
xnor U15116 (N_15116,N_14093,N_13808);
nor U15117 (N_15117,N_13846,N_13660);
nor U15118 (N_15118,N_13371,N_13621);
nor U15119 (N_15119,N_14057,N_13530);
nand U15120 (N_15120,N_14155,N_13995);
xor U15121 (N_15121,N_14293,N_13776);
nor U15122 (N_15122,N_13989,N_13659);
nor U15123 (N_15123,N_13954,N_13565);
and U15124 (N_15124,N_13985,N_13311);
nor U15125 (N_15125,N_14225,N_14304);
and U15126 (N_15126,N_14140,N_13232);
nand U15127 (N_15127,N_14020,N_14117);
nor U15128 (N_15128,N_13549,N_13461);
or U15129 (N_15129,N_14358,N_14046);
and U15130 (N_15130,N_13392,N_14120);
nor U15131 (N_15131,N_14056,N_14058);
or U15132 (N_15132,N_14021,N_14284);
nor U15133 (N_15133,N_13565,N_14045);
nand U15134 (N_15134,N_14053,N_14200);
or U15135 (N_15135,N_13283,N_13712);
and U15136 (N_15136,N_14133,N_13841);
nor U15137 (N_15137,N_14363,N_13455);
nand U15138 (N_15138,N_13638,N_13434);
or U15139 (N_15139,N_14177,N_13267);
nand U15140 (N_15140,N_13266,N_14120);
or U15141 (N_15141,N_13927,N_13853);
nor U15142 (N_15142,N_13367,N_13223);
nand U15143 (N_15143,N_14074,N_13300);
xnor U15144 (N_15144,N_13362,N_13295);
nor U15145 (N_15145,N_13529,N_13559);
nand U15146 (N_15146,N_13265,N_13642);
nor U15147 (N_15147,N_13491,N_13496);
and U15148 (N_15148,N_14203,N_13817);
nor U15149 (N_15149,N_13733,N_13997);
xnor U15150 (N_15150,N_14391,N_14065);
xor U15151 (N_15151,N_13865,N_13596);
and U15152 (N_15152,N_14134,N_13762);
and U15153 (N_15153,N_14167,N_13947);
nor U15154 (N_15154,N_14202,N_13876);
or U15155 (N_15155,N_14399,N_13857);
nor U15156 (N_15156,N_13467,N_13771);
xor U15157 (N_15157,N_13512,N_13523);
or U15158 (N_15158,N_13712,N_13845);
xor U15159 (N_15159,N_14234,N_13479);
and U15160 (N_15160,N_13979,N_13826);
nand U15161 (N_15161,N_13798,N_13876);
or U15162 (N_15162,N_13591,N_13974);
nand U15163 (N_15163,N_13238,N_13757);
nand U15164 (N_15164,N_13496,N_13462);
and U15165 (N_15165,N_13755,N_13695);
nand U15166 (N_15166,N_13600,N_14238);
and U15167 (N_15167,N_13995,N_14078);
nand U15168 (N_15168,N_14093,N_14296);
and U15169 (N_15169,N_13685,N_13354);
xor U15170 (N_15170,N_13362,N_13834);
nor U15171 (N_15171,N_13886,N_13550);
and U15172 (N_15172,N_13954,N_14382);
nand U15173 (N_15173,N_13394,N_13650);
nand U15174 (N_15174,N_14314,N_13816);
xor U15175 (N_15175,N_13435,N_13769);
nand U15176 (N_15176,N_13380,N_14112);
nand U15177 (N_15177,N_13640,N_14010);
xnor U15178 (N_15178,N_13426,N_14108);
xor U15179 (N_15179,N_14211,N_14181);
xnor U15180 (N_15180,N_14316,N_14328);
nand U15181 (N_15181,N_13437,N_14209);
xnor U15182 (N_15182,N_13932,N_13315);
nand U15183 (N_15183,N_14189,N_13856);
xnor U15184 (N_15184,N_13333,N_13245);
or U15185 (N_15185,N_14270,N_14251);
or U15186 (N_15186,N_13472,N_13430);
xnor U15187 (N_15187,N_13438,N_14034);
or U15188 (N_15188,N_13380,N_13865);
nor U15189 (N_15189,N_13910,N_13888);
or U15190 (N_15190,N_13928,N_13790);
nand U15191 (N_15191,N_13606,N_13831);
xnor U15192 (N_15192,N_13590,N_13371);
or U15193 (N_15193,N_13942,N_14320);
nand U15194 (N_15194,N_14217,N_13916);
or U15195 (N_15195,N_13249,N_13419);
nor U15196 (N_15196,N_13477,N_13803);
xor U15197 (N_15197,N_14123,N_13684);
nand U15198 (N_15198,N_13799,N_13977);
nand U15199 (N_15199,N_13454,N_13222);
and U15200 (N_15200,N_13237,N_14263);
xor U15201 (N_15201,N_13380,N_14270);
nor U15202 (N_15202,N_13565,N_14235);
nor U15203 (N_15203,N_13776,N_13673);
or U15204 (N_15204,N_13780,N_14229);
and U15205 (N_15205,N_13320,N_13639);
or U15206 (N_15206,N_13631,N_14223);
and U15207 (N_15207,N_14203,N_13435);
xnor U15208 (N_15208,N_14151,N_13990);
or U15209 (N_15209,N_13592,N_14105);
and U15210 (N_15210,N_13362,N_13649);
nand U15211 (N_15211,N_13831,N_13891);
xor U15212 (N_15212,N_13980,N_13307);
xnor U15213 (N_15213,N_14094,N_14267);
nand U15214 (N_15214,N_14047,N_13463);
and U15215 (N_15215,N_14364,N_13592);
nand U15216 (N_15216,N_13996,N_13750);
or U15217 (N_15217,N_13747,N_13904);
or U15218 (N_15218,N_13743,N_14370);
or U15219 (N_15219,N_13959,N_13396);
nand U15220 (N_15220,N_14311,N_14385);
or U15221 (N_15221,N_13456,N_13788);
nor U15222 (N_15222,N_13837,N_13453);
or U15223 (N_15223,N_13541,N_13247);
nor U15224 (N_15224,N_13318,N_13943);
nor U15225 (N_15225,N_13327,N_13801);
nand U15226 (N_15226,N_13671,N_13687);
nor U15227 (N_15227,N_13564,N_13582);
nand U15228 (N_15228,N_14323,N_13654);
xnor U15229 (N_15229,N_13529,N_13966);
xor U15230 (N_15230,N_13296,N_14241);
or U15231 (N_15231,N_13746,N_13209);
nor U15232 (N_15232,N_13879,N_13707);
xnor U15233 (N_15233,N_14306,N_13792);
xnor U15234 (N_15234,N_13975,N_14159);
or U15235 (N_15235,N_14168,N_13711);
and U15236 (N_15236,N_13879,N_13305);
and U15237 (N_15237,N_14108,N_13424);
or U15238 (N_15238,N_13781,N_13554);
nor U15239 (N_15239,N_13832,N_13656);
or U15240 (N_15240,N_13341,N_13987);
or U15241 (N_15241,N_13683,N_13429);
xnor U15242 (N_15242,N_13249,N_13972);
or U15243 (N_15243,N_13264,N_14061);
or U15244 (N_15244,N_14083,N_13459);
nand U15245 (N_15245,N_14384,N_13761);
nand U15246 (N_15246,N_14005,N_13473);
nor U15247 (N_15247,N_13916,N_13694);
or U15248 (N_15248,N_14154,N_14001);
nand U15249 (N_15249,N_13455,N_14150);
xor U15250 (N_15250,N_13350,N_13893);
or U15251 (N_15251,N_14217,N_14125);
and U15252 (N_15252,N_13972,N_14012);
nor U15253 (N_15253,N_14008,N_13488);
nor U15254 (N_15254,N_14260,N_13325);
nor U15255 (N_15255,N_13923,N_13932);
nor U15256 (N_15256,N_14164,N_14377);
nand U15257 (N_15257,N_14196,N_13666);
nand U15258 (N_15258,N_14140,N_13415);
or U15259 (N_15259,N_13274,N_13598);
or U15260 (N_15260,N_13274,N_13806);
nor U15261 (N_15261,N_13746,N_13334);
or U15262 (N_15262,N_13781,N_13669);
nor U15263 (N_15263,N_13444,N_13540);
or U15264 (N_15264,N_13530,N_13641);
nand U15265 (N_15265,N_14347,N_14203);
nand U15266 (N_15266,N_13458,N_14395);
or U15267 (N_15267,N_13623,N_14354);
nand U15268 (N_15268,N_14073,N_13227);
nor U15269 (N_15269,N_13909,N_13478);
xor U15270 (N_15270,N_13576,N_13261);
or U15271 (N_15271,N_13610,N_13873);
or U15272 (N_15272,N_14251,N_14263);
and U15273 (N_15273,N_13698,N_14312);
or U15274 (N_15274,N_14004,N_14363);
nor U15275 (N_15275,N_13510,N_13580);
nor U15276 (N_15276,N_14146,N_13932);
nand U15277 (N_15277,N_13816,N_14283);
nand U15278 (N_15278,N_14068,N_13509);
xor U15279 (N_15279,N_14297,N_13439);
or U15280 (N_15280,N_14288,N_13543);
or U15281 (N_15281,N_13587,N_13246);
nand U15282 (N_15282,N_14306,N_13961);
xnor U15283 (N_15283,N_13584,N_13485);
xor U15284 (N_15284,N_14083,N_14282);
xor U15285 (N_15285,N_14124,N_13958);
xor U15286 (N_15286,N_13443,N_14064);
and U15287 (N_15287,N_13457,N_14305);
and U15288 (N_15288,N_13477,N_13348);
nand U15289 (N_15289,N_13904,N_13200);
nor U15290 (N_15290,N_13287,N_14379);
xnor U15291 (N_15291,N_14188,N_13303);
xnor U15292 (N_15292,N_14355,N_13254);
or U15293 (N_15293,N_13258,N_13240);
nand U15294 (N_15294,N_14104,N_14139);
or U15295 (N_15295,N_13291,N_13330);
and U15296 (N_15296,N_13279,N_13979);
xnor U15297 (N_15297,N_14170,N_14138);
xor U15298 (N_15298,N_13404,N_13248);
or U15299 (N_15299,N_13241,N_14176);
nor U15300 (N_15300,N_13685,N_13484);
and U15301 (N_15301,N_13668,N_13401);
and U15302 (N_15302,N_13681,N_13326);
xnor U15303 (N_15303,N_13660,N_13922);
xnor U15304 (N_15304,N_13995,N_14285);
or U15305 (N_15305,N_13781,N_14380);
nor U15306 (N_15306,N_14234,N_13330);
nor U15307 (N_15307,N_13982,N_13555);
nand U15308 (N_15308,N_13426,N_13231);
nor U15309 (N_15309,N_13927,N_14244);
and U15310 (N_15310,N_13621,N_13215);
xor U15311 (N_15311,N_14238,N_13515);
and U15312 (N_15312,N_14069,N_14198);
nor U15313 (N_15313,N_14393,N_14011);
xnor U15314 (N_15314,N_14140,N_14316);
nand U15315 (N_15315,N_14022,N_13915);
and U15316 (N_15316,N_13891,N_14268);
xnor U15317 (N_15317,N_14288,N_13954);
or U15318 (N_15318,N_14317,N_13295);
xnor U15319 (N_15319,N_13435,N_13500);
and U15320 (N_15320,N_14007,N_14231);
nand U15321 (N_15321,N_14342,N_13765);
or U15322 (N_15322,N_13942,N_13943);
or U15323 (N_15323,N_13816,N_13635);
or U15324 (N_15324,N_14043,N_13795);
and U15325 (N_15325,N_13594,N_14283);
nand U15326 (N_15326,N_14128,N_13614);
and U15327 (N_15327,N_13987,N_13464);
xor U15328 (N_15328,N_13215,N_14254);
and U15329 (N_15329,N_13880,N_13689);
xor U15330 (N_15330,N_14285,N_13411);
and U15331 (N_15331,N_13700,N_14331);
nor U15332 (N_15332,N_13934,N_13654);
xor U15333 (N_15333,N_13486,N_13974);
xnor U15334 (N_15334,N_13713,N_14354);
and U15335 (N_15335,N_14154,N_14275);
xnor U15336 (N_15336,N_13595,N_13923);
xor U15337 (N_15337,N_14080,N_13415);
nand U15338 (N_15338,N_13608,N_13432);
xor U15339 (N_15339,N_13603,N_13290);
nor U15340 (N_15340,N_13204,N_13607);
and U15341 (N_15341,N_14112,N_14227);
and U15342 (N_15342,N_13584,N_14066);
or U15343 (N_15343,N_13572,N_14028);
and U15344 (N_15344,N_13264,N_13904);
xor U15345 (N_15345,N_13312,N_13221);
xor U15346 (N_15346,N_13210,N_14372);
xnor U15347 (N_15347,N_14064,N_13923);
nand U15348 (N_15348,N_13776,N_13431);
and U15349 (N_15349,N_14020,N_14276);
or U15350 (N_15350,N_13999,N_13975);
xor U15351 (N_15351,N_13659,N_13253);
xor U15352 (N_15352,N_14160,N_14356);
and U15353 (N_15353,N_13454,N_14266);
xnor U15354 (N_15354,N_13293,N_13792);
nand U15355 (N_15355,N_13497,N_13674);
or U15356 (N_15356,N_13601,N_14049);
nor U15357 (N_15357,N_14288,N_13860);
nor U15358 (N_15358,N_13581,N_13790);
xor U15359 (N_15359,N_13827,N_13453);
or U15360 (N_15360,N_13444,N_13819);
nand U15361 (N_15361,N_14209,N_13564);
or U15362 (N_15362,N_14229,N_13499);
xor U15363 (N_15363,N_13301,N_13587);
and U15364 (N_15364,N_14246,N_13207);
xnor U15365 (N_15365,N_13561,N_13621);
or U15366 (N_15366,N_14203,N_13334);
nand U15367 (N_15367,N_13411,N_13647);
or U15368 (N_15368,N_14149,N_13803);
nand U15369 (N_15369,N_13359,N_14267);
and U15370 (N_15370,N_14360,N_14370);
xor U15371 (N_15371,N_13496,N_13619);
nor U15372 (N_15372,N_13536,N_13772);
nand U15373 (N_15373,N_14238,N_13478);
nand U15374 (N_15374,N_14272,N_13581);
xor U15375 (N_15375,N_13918,N_14024);
nor U15376 (N_15376,N_13275,N_13328);
nand U15377 (N_15377,N_13407,N_13442);
nor U15378 (N_15378,N_14336,N_14317);
xor U15379 (N_15379,N_13430,N_14215);
or U15380 (N_15380,N_13917,N_13962);
and U15381 (N_15381,N_14398,N_13790);
or U15382 (N_15382,N_14224,N_13328);
or U15383 (N_15383,N_14289,N_14081);
and U15384 (N_15384,N_14212,N_13307);
xor U15385 (N_15385,N_13474,N_13881);
and U15386 (N_15386,N_13347,N_13640);
xnor U15387 (N_15387,N_13769,N_13487);
or U15388 (N_15388,N_13630,N_14023);
nand U15389 (N_15389,N_13461,N_14342);
nor U15390 (N_15390,N_14027,N_13205);
and U15391 (N_15391,N_13975,N_13576);
or U15392 (N_15392,N_14001,N_13341);
xor U15393 (N_15393,N_13872,N_13500);
xor U15394 (N_15394,N_14372,N_13445);
nor U15395 (N_15395,N_13234,N_14260);
xor U15396 (N_15396,N_13241,N_14248);
or U15397 (N_15397,N_13856,N_14104);
and U15398 (N_15398,N_14078,N_13454);
or U15399 (N_15399,N_13435,N_13423);
nand U15400 (N_15400,N_14302,N_13634);
or U15401 (N_15401,N_14203,N_13221);
and U15402 (N_15402,N_13365,N_13219);
or U15403 (N_15403,N_14126,N_13669);
nor U15404 (N_15404,N_13563,N_13245);
or U15405 (N_15405,N_13489,N_13493);
nand U15406 (N_15406,N_14392,N_14134);
nor U15407 (N_15407,N_14105,N_13693);
nor U15408 (N_15408,N_13603,N_13533);
or U15409 (N_15409,N_13832,N_13368);
nor U15410 (N_15410,N_13754,N_14354);
and U15411 (N_15411,N_14315,N_13403);
nor U15412 (N_15412,N_13702,N_13322);
nor U15413 (N_15413,N_13924,N_14083);
or U15414 (N_15414,N_14209,N_14050);
nor U15415 (N_15415,N_13239,N_14365);
and U15416 (N_15416,N_13292,N_13447);
or U15417 (N_15417,N_13676,N_14258);
nor U15418 (N_15418,N_13798,N_14355);
or U15419 (N_15419,N_13868,N_13914);
nor U15420 (N_15420,N_13365,N_13883);
xor U15421 (N_15421,N_13660,N_14213);
and U15422 (N_15422,N_13292,N_13787);
or U15423 (N_15423,N_13438,N_14025);
xnor U15424 (N_15424,N_14258,N_13508);
xnor U15425 (N_15425,N_13385,N_13844);
nor U15426 (N_15426,N_14258,N_13569);
nand U15427 (N_15427,N_13842,N_13317);
nor U15428 (N_15428,N_14234,N_13280);
and U15429 (N_15429,N_14042,N_14133);
or U15430 (N_15430,N_14358,N_14333);
or U15431 (N_15431,N_14334,N_14105);
nor U15432 (N_15432,N_13286,N_14256);
or U15433 (N_15433,N_13868,N_13252);
or U15434 (N_15434,N_13913,N_14184);
nand U15435 (N_15435,N_13333,N_13460);
nand U15436 (N_15436,N_13442,N_13676);
xnor U15437 (N_15437,N_14209,N_14008);
or U15438 (N_15438,N_13255,N_13774);
and U15439 (N_15439,N_13312,N_14382);
nand U15440 (N_15440,N_13223,N_14296);
or U15441 (N_15441,N_14316,N_13453);
xor U15442 (N_15442,N_13859,N_13460);
or U15443 (N_15443,N_14110,N_13254);
or U15444 (N_15444,N_14119,N_14185);
xnor U15445 (N_15445,N_13573,N_13392);
nor U15446 (N_15446,N_14327,N_14128);
or U15447 (N_15447,N_13328,N_13409);
nor U15448 (N_15448,N_13874,N_14094);
nand U15449 (N_15449,N_14175,N_13654);
nand U15450 (N_15450,N_14175,N_13367);
or U15451 (N_15451,N_13342,N_14031);
nor U15452 (N_15452,N_14185,N_13927);
xnor U15453 (N_15453,N_13683,N_14169);
nor U15454 (N_15454,N_14166,N_14275);
nand U15455 (N_15455,N_14025,N_13730);
nand U15456 (N_15456,N_14346,N_13527);
nor U15457 (N_15457,N_13987,N_13531);
nand U15458 (N_15458,N_13354,N_13845);
nand U15459 (N_15459,N_13815,N_13923);
and U15460 (N_15460,N_13562,N_13504);
nor U15461 (N_15461,N_13517,N_13430);
nor U15462 (N_15462,N_14266,N_14140);
nor U15463 (N_15463,N_13889,N_13335);
xor U15464 (N_15464,N_13721,N_14045);
or U15465 (N_15465,N_13644,N_13940);
or U15466 (N_15466,N_14183,N_13568);
xor U15467 (N_15467,N_13869,N_13330);
xor U15468 (N_15468,N_14355,N_13387);
and U15469 (N_15469,N_14048,N_13789);
xnor U15470 (N_15470,N_14170,N_14031);
nand U15471 (N_15471,N_14235,N_14143);
xnor U15472 (N_15472,N_13825,N_14058);
or U15473 (N_15473,N_13255,N_13921);
xor U15474 (N_15474,N_13396,N_14153);
nor U15475 (N_15475,N_13878,N_13406);
xor U15476 (N_15476,N_13388,N_13531);
nor U15477 (N_15477,N_14099,N_13423);
or U15478 (N_15478,N_14296,N_14355);
and U15479 (N_15479,N_14390,N_13263);
nor U15480 (N_15480,N_13551,N_13980);
nor U15481 (N_15481,N_13412,N_13428);
nand U15482 (N_15482,N_14045,N_13282);
xor U15483 (N_15483,N_13400,N_14025);
or U15484 (N_15484,N_14280,N_13911);
xnor U15485 (N_15485,N_14228,N_13568);
nand U15486 (N_15486,N_13344,N_14132);
xnor U15487 (N_15487,N_13722,N_14335);
xor U15488 (N_15488,N_14326,N_13354);
or U15489 (N_15489,N_13770,N_14243);
and U15490 (N_15490,N_13290,N_14032);
nor U15491 (N_15491,N_13891,N_14316);
and U15492 (N_15492,N_13866,N_13636);
or U15493 (N_15493,N_13503,N_13856);
xor U15494 (N_15494,N_14061,N_14065);
and U15495 (N_15495,N_14060,N_14018);
nor U15496 (N_15496,N_13469,N_13877);
and U15497 (N_15497,N_13944,N_14370);
nor U15498 (N_15498,N_13575,N_14062);
or U15499 (N_15499,N_14352,N_13913);
xor U15500 (N_15500,N_13879,N_14026);
xor U15501 (N_15501,N_14286,N_13947);
and U15502 (N_15502,N_13733,N_13418);
xnor U15503 (N_15503,N_14038,N_13564);
xnor U15504 (N_15504,N_13268,N_13827);
nand U15505 (N_15505,N_13672,N_14320);
xnor U15506 (N_15506,N_13480,N_14165);
nand U15507 (N_15507,N_13247,N_13501);
or U15508 (N_15508,N_13762,N_14316);
nor U15509 (N_15509,N_13232,N_13596);
nand U15510 (N_15510,N_14226,N_13381);
xor U15511 (N_15511,N_13513,N_13369);
and U15512 (N_15512,N_14325,N_13348);
and U15513 (N_15513,N_14048,N_13697);
or U15514 (N_15514,N_13235,N_13559);
or U15515 (N_15515,N_14272,N_13966);
nand U15516 (N_15516,N_14172,N_13755);
xor U15517 (N_15517,N_14117,N_14274);
nor U15518 (N_15518,N_13225,N_13483);
or U15519 (N_15519,N_13906,N_13276);
or U15520 (N_15520,N_13967,N_14225);
nand U15521 (N_15521,N_14396,N_13526);
xnor U15522 (N_15522,N_13803,N_14335);
and U15523 (N_15523,N_13323,N_14026);
and U15524 (N_15524,N_14230,N_13415);
nand U15525 (N_15525,N_13465,N_13537);
or U15526 (N_15526,N_13327,N_13283);
xor U15527 (N_15527,N_13967,N_13868);
xnor U15528 (N_15528,N_13284,N_14139);
nor U15529 (N_15529,N_14043,N_14197);
and U15530 (N_15530,N_14291,N_14252);
nand U15531 (N_15531,N_13309,N_13437);
and U15532 (N_15532,N_13417,N_13975);
or U15533 (N_15533,N_13262,N_14345);
nor U15534 (N_15534,N_13265,N_13270);
nor U15535 (N_15535,N_13971,N_13736);
and U15536 (N_15536,N_13419,N_14126);
or U15537 (N_15537,N_14261,N_13761);
nand U15538 (N_15538,N_14101,N_13349);
xor U15539 (N_15539,N_13555,N_13671);
or U15540 (N_15540,N_13369,N_13340);
or U15541 (N_15541,N_13843,N_13779);
or U15542 (N_15542,N_13690,N_13619);
xnor U15543 (N_15543,N_14077,N_14288);
xor U15544 (N_15544,N_13470,N_13895);
xor U15545 (N_15545,N_13719,N_13866);
or U15546 (N_15546,N_13817,N_14153);
nor U15547 (N_15547,N_13856,N_13305);
nor U15548 (N_15548,N_13817,N_13262);
nor U15549 (N_15549,N_14265,N_14305);
or U15550 (N_15550,N_13804,N_13304);
nand U15551 (N_15551,N_13285,N_13779);
and U15552 (N_15552,N_13667,N_13872);
and U15553 (N_15553,N_13608,N_14133);
nand U15554 (N_15554,N_14309,N_13582);
nand U15555 (N_15555,N_14180,N_14010);
or U15556 (N_15556,N_14296,N_14335);
nor U15557 (N_15557,N_13599,N_14197);
or U15558 (N_15558,N_14019,N_13581);
nor U15559 (N_15559,N_13798,N_13837);
nand U15560 (N_15560,N_13530,N_14385);
and U15561 (N_15561,N_13254,N_14019);
and U15562 (N_15562,N_13418,N_13668);
nor U15563 (N_15563,N_13855,N_13724);
and U15564 (N_15564,N_13641,N_14154);
nor U15565 (N_15565,N_13644,N_13285);
nand U15566 (N_15566,N_13423,N_14260);
or U15567 (N_15567,N_13968,N_13639);
xor U15568 (N_15568,N_13551,N_13459);
xor U15569 (N_15569,N_13548,N_14110);
nor U15570 (N_15570,N_13624,N_14092);
and U15571 (N_15571,N_13578,N_13682);
nor U15572 (N_15572,N_14388,N_14312);
nand U15573 (N_15573,N_14070,N_13816);
nand U15574 (N_15574,N_14137,N_13981);
nor U15575 (N_15575,N_13678,N_13764);
xnor U15576 (N_15576,N_13752,N_13983);
or U15577 (N_15577,N_14143,N_14260);
and U15578 (N_15578,N_14169,N_13845);
nand U15579 (N_15579,N_13762,N_13567);
xnor U15580 (N_15580,N_13632,N_14149);
xor U15581 (N_15581,N_13331,N_13645);
or U15582 (N_15582,N_14068,N_13980);
xor U15583 (N_15583,N_14181,N_13939);
nor U15584 (N_15584,N_14213,N_13298);
nand U15585 (N_15585,N_13956,N_13980);
xor U15586 (N_15586,N_13852,N_13763);
and U15587 (N_15587,N_13652,N_14246);
xor U15588 (N_15588,N_13228,N_14360);
nor U15589 (N_15589,N_13797,N_13315);
nand U15590 (N_15590,N_13663,N_13884);
xnor U15591 (N_15591,N_13640,N_13202);
xnor U15592 (N_15592,N_14240,N_13681);
nand U15593 (N_15593,N_13479,N_14323);
nor U15594 (N_15594,N_13468,N_13703);
nand U15595 (N_15595,N_14008,N_13360);
and U15596 (N_15596,N_13431,N_13381);
nand U15597 (N_15597,N_14336,N_14204);
nand U15598 (N_15598,N_13637,N_13670);
or U15599 (N_15599,N_13306,N_13624);
nand U15600 (N_15600,N_15001,N_14979);
xor U15601 (N_15601,N_14969,N_14540);
or U15602 (N_15602,N_15166,N_15497);
or U15603 (N_15603,N_14818,N_14603);
xnor U15604 (N_15604,N_15230,N_14937);
nor U15605 (N_15605,N_14710,N_14422);
and U15606 (N_15606,N_15360,N_14994);
nor U15607 (N_15607,N_15154,N_15110);
nand U15608 (N_15608,N_15498,N_15096);
and U15609 (N_15609,N_15133,N_14441);
and U15610 (N_15610,N_15580,N_14981);
and U15611 (N_15611,N_15376,N_14401);
and U15612 (N_15612,N_14986,N_15218);
nand U15613 (N_15613,N_15045,N_14700);
xnor U15614 (N_15614,N_14703,N_15344);
xor U15615 (N_15615,N_14760,N_15517);
and U15616 (N_15616,N_15155,N_15552);
and U15617 (N_15617,N_15228,N_14565);
nand U15618 (N_15618,N_14910,N_14506);
or U15619 (N_15619,N_14694,N_15406);
nand U15620 (N_15620,N_15056,N_14460);
nor U15621 (N_15621,N_14742,N_15407);
nand U15622 (N_15622,N_15310,N_15329);
or U15623 (N_15623,N_15305,N_14610);
or U15624 (N_15624,N_14531,N_15184);
or U15625 (N_15625,N_15384,N_14504);
and U15626 (N_15626,N_15378,N_15152);
nand U15627 (N_15627,N_14799,N_15239);
and U15628 (N_15628,N_15539,N_15504);
xnor U15629 (N_15629,N_14502,N_14826);
nor U15630 (N_15630,N_15291,N_14747);
or U15631 (N_15631,N_14496,N_15182);
and U15632 (N_15632,N_15177,N_14882);
nand U15633 (N_15633,N_14663,N_15104);
nor U15634 (N_15634,N_14941,N_14998);
or U15635 (N_15635,N_15348,N_14854);
nor U15636 (N_15636,N_14491,N_14844);
and U15637 (N_15637,N_15282,N_14575);
nor U15638 (N_15638,N_14995,N_15509);
nor U15639 (N_15639,N_15060,N_14970);
and U15640 (N_15640,N_15250,N_14641);
nor U15641 (N_15641,N_14696,N_15191);
and U15642 (N_15642,N_15401,N_15074);
nand U15643 (N_15643,N_15468,N_14697);
xor U15644 (N_15644,N_15064,N_15272);
and U15645 (N_15645,N_14681,N_14613);
or U15646 (N_15646,N_14482,N_15400);
and U15647 (N_15647,N_15138,N_15506);
xnor U15648 (N_15648,N_14616,N_15253);
xor U15649 (N_15649,N_14493,N_14691);
and U15650 (N_15650,N_15345,N_15578);
xnor U15651 (N_15651,N_15148,N_15485);
and U15652 (N_15652,N_14840,N_15025);
or U15653 (N_15653,N_14608,N_15508);
nor U15654 (N_15654,N_15264,N_14604);
nor U15655 (N_15655,N_14664,N_15017);
and U15656 (N_15656,N_15099,N_15334);
and U15657 (N_15657,N_15303,N_15494);
and U15658 (N_15658,N_15240,N_14577);
nor U15659 (N_15659,N_15582,N_15313);
nor U15660 (N_15660,N_15559,N_14458);
nand U15661 (N_15661,N_14602,N_15161);
xor U15662 (N_15662,N_14545,N_15170);
nor U15663 (N_15663,N_14730,N_14606);
or U15664 (N_15664,N_15553,N_14961);
and U15665 (N_15665,N_14943,N_14815);
xor U15666 (N_15666,N_14601,N_14906);
or U15667 (N_15667,N_14476,N_14472);
nor U15668 (N_15668,N_14911,N_15091);
nor U15669 (N_15669,N_15077,N_14816);
nor U15670 (N_15670,N_15530,N_15260);
nor U15671 (N_15671,N_14657,N_14925);
and U15672 (N_15672,N_14962,N_15267);
nand U15673 (N_15673,N_15458,N_14440);
nand U15674 (N_15674,N_14558,N_15192);
xnor U15675 (N_15675,N_14876,N_14791);
nand U15676 (N_15676,N_15489,N_14438);
xor U15677 (N_15677,N_14617,N_14521);
and U15678 (N_15678,N_15076,N_15404);
xnor U15679 (N_15679,N_15548,N_14611);
and U15680 (N_15680,N_14678,N_15034);
and U15681 (N_15681,N_15123,N_14780);
and U15682 (N_15682,N_14808,N_14933);
xnor U15683 (N_15683,N_14772,N_14503);
and U15684 (N_15684,N_14661,N_14989);
or U15685 (N_15685,N_14427,N_15487);
and U15686 (N_15686,N_15531,N_14529);
and U15687 (N_15687,N_14570,N_15373);
nor U15688 (N_15688,N_15231,N_15036);
and U15689 (N_15689,N_15052,N_14542);
nand U15690 (N_15690,N_14865,N_15270);
and U15691 (N_15691,N_14701,N_15377);
xnor U15692 (N_15692,N_15335,N_14964);
nor U15693 (N_15693,N_14938,N_14966);
xor U15694 (N_15694,N_14515,N_14878);
or U15695 (N_15695,N_15281,N_15010);
or U15696 (N_15696,N_14402,N_15511);
and U15697 (N_15697,N_14477,N_15273);
and U15698 (N_15698,N_15311,N_15385);
or U15699 (N_15699,N_15143,N_14927);
and U15700 (N_15700,N_15419,N_14907);
or U15701 (N_15701,N_14492,N_15343);
or U15702 (N_15702,N_15245,N_15187);
and U15703 (N_15703,N_15368,N_14487);
and U15704 (N_15704,N_14481,N_15190);
or U15705 (N_15705,N_15212,N_14899);
or U15706 (N_15706,N_14810,N_15551);
xor U15707 (N_15707,N_15083,N_14639);
or U15708 (N_15708,N_14413,N_14766);
nand U15709 (N_15709,N_14673,N_14405);
xnor U15710 (N_15710,N_15442,N_15564);
xor U15711 (N_15711,N_14952,N_15470);
xor U15712 (N_15712,N_15082,N_15295);
and U15713 (N_15713,N_15003,N_15249);
nand U15714 (N_15714,N_14773,N_14547);
xnor U15715 (N_15715,N_15501,N_15037);
nand U15716 (N_15716,N_14588,N_15416);
and U15717 (N_15717,N_15337,N_14709);
nor U15718 (N_15718,N_14972,N_14444);
or U15719 (N_15719,N_15464,N_14853);
nand U15720 (N_15720,N_14524,N_15535);
xnor U15721 (N_15721,N_14765,N_14729);
and U15722 (N_15722,N_15292,N_15226);
nand U15723 (N_15723,N_14984,N_14722);
or U15724 (N_15724,N_15225,N_15463);
xor U15725 (N_15725,N_15537,N_15180);
or U15726 (N_15726,N_15032,N_14516);
nor U15727 (N_15727,N_14647,N_15274);
nor U15728 (N_15728,N_15132,N_15567);
or U15729 (N_15729,N_15573,N_15179);
and U15730 (N_15730,N_15069,N_15579);
and U15731 (N_15731,N_14946,N_14787);
nand U15732 (N_15732,N_14900,N_14828);
nand U15733 (N_15733,N_15205,N_14676);
and U15734 (N_15734,N_14825,N_14555);
nor U15735 (N_15735,N_15374,N_14877);
nand U15736 (N_15736,N_14692,N_14450);
and U15737 (N_15737,N_14636,N_15331);
nand U15738 (N_15738,N_15061,N_14432);
or U15739 (N_15739,N_14645,N_14586);
and U15740 (N_15740,N_15493,N_15103);
and U15741 (N_15741,N_14625,N_14716);
xnor U15742 (N_15742,N_14967,N_15043);
nand U15743 (N_15743,N_15362,N_15048);
and U15744 (N_15744,N_15302,N_15340);
or U15745 (N_15745,N_15444,N_14842);
nand U15746 (N_15746,N_14839,N_15097);
nand U15747 (N_15747,N_15262,N_14754);
or U15748 (N_15748,N_15095,N_15481);
nor U15749 (N_15749,N_15484,N_14607);
xor U15750 (N_15750,N_14426,N_14687);
nand U15751 (N_15751,N_15290,N_14939);
or U15752 (N_15752,N_15333,N_14408);
nor U15753 (N_15753,N_15561,N_15008);
or U15754 (N_15754,N_15536,N_14934);
xor U15755 (N_15755,N_14403,N_15206);
and U15756 (N_15756,N_15092,N_14598);
or U15757 (N_15757,N_14746,N_15421);
nor U15758 (N_15758,N_14424,N_15546);
and U15759 (N_15759,N_15323,N_15156);
xor U15760 (N_15760,N_15426,N_14576);
nand U15761 (N_15761,N_14761,N_14582);
nor U15762 (N_15762,N_14740,N_14439);
and U15763 (N_15763,N_14649,N_14499);
nand U15764 (N_15764,N_15558,N_15046);
nor U15765 (N_15765,N_15448,N_15107);
or U15766 (N_15766,N_14571,N_14705);
and U15767 (N_15767,N_15248,N_14612);
nor U15768 (N_15768,N_14505,N_15058);
or U15769 (N_15769,N_15146,N_14718);
nor U15770 (N_15770,N_14976,N_15460);
or U15771 (N_15771,N_15178,N_15255);
xnor U15772 (N_15772,N_15028,N_15112);
or U15773 (N_15773,N_14860,N_15284);
xor U15774 (N_15774,N_14843,N_15140);
nand U15775 (N_15775,N_14638,N_15457);
or U15776 (N_15776,N_15369,N_14759);
xor U15777 (N_15777,N_14414,N_14656);
nand U15778 (N_15778,N_14669,N_15533);
xor U15779 (N_15779,N_15306,N_14559);
nor U15780 (N_15780,N_14778,N_14707);
nand U15781 (N_15781,N_15322,N_14881);
nand U15782 (N_15782,N_15592,N_14490);
and U15783 (N_15783,N_14530,N_14659);
nand U15784 (N_15784,N_14695,N_15298);
or U15785 (N_15785,N_15007,N_14903);
or U15786 (N_15786,N_15475,N_15137);
or U15787 (N_15787,N_15529,N_14532);
xnor U15788 (N_15788,N_15173,N_15275);
or U15789 (N_15789,N_14406,N_14820);
nor U15790 (N_15790,N_14795,N_14551);
nand U15791 (N_15791,N_15365,N_15440);
xor U15792 (N_15792,N_15574,N_14862);
and U15793 (N_15793,N_14419,N_14561);
or U15794 (N_15794,N_15391,N_15486);
or U15795 (N_15795,N_15087,N_14596);
nand U15796 (N_15796,N_14640,N_15051);
nand U15797 (N_15797,N_14968,N_15382);
nor U15798 (N_15798,N_14400,N_15174);
nand U15799 (N_15799,N_14523,N_15540);
xor U15800 (N_15800,N_15241,N_14956);
nand U15801 (N_15801,N_15113,N_15328);
nor U15802 (N_15802,N_14717,N_15462);
and U15803 (N_15803,N_15522,N_14668);
or U15804 (N_15804,N_15189,N_15106);
xor U15805 (N_15805,N_14831,N_15588);
nor U15806 (N_15806,N_15167,N_15186);
and U15807 (N_15807,N_14861,N_15024);
nor U15808 (N_15808,N_15293,N_15432);
or U15809 (N_15809,N_14985,N_15049);
or U15810 (N_15810,N_14548,N_15118);
and U15811 (N_15811,N_14893,N_14800);
and U15812 (N_15812,N_15409,N_15185);
nand U15813 (N_15813,N_15346,N_15568);
nand U15814 (N_15814,N_14684,N_14553);
nor U15815 (N_15815,N_15480,N_14873);
or U15816 (N_15816,N_14999,N_15414);
nor U15817 (N_15817,N_14848,N_15317);
or U15818 (N_15818,N_15397,N_14782);
or U15819 (N_15819,N_15288,N_14660);
nor U15820 (N_15820,N_15220,N_14958);
nor U15821 (N_15821,N_14845,N_14744);
xor U15822 (N_15822,N_14855,N_15342);
xnor U15823 (N_15823,N_15236,N_14822);
nor U15824 (N_15824,N_15521,N_14654);
and U15825 (N_15825,N_15338,N_15439);
and U15826 (N_15826,N_14735,N_14887);
xor U15827 (N_15827,N_14512,N_15098);
or U15828 (N_15828,N_14856,N_14960);
xor U15829 (N_15829,N_14753,N_14779);
nor U15830 (N_15830,N_15300,N_14836);
nand U15831 (N_15831,N_15398,N_14615);
nand U15832 (N_15832,N_15483,N_15129);
and U15833 (N_15833,N_15066,N_14417);
xnor U15834 (N_15834,N_14751,N_15589);
and U15835 (N_15835,N_15027,N_15512);
or U15836 (N_15836,N_15075,N_15354);
nor U15837 (N_15837,N_15394,N_14886);
nand U15838 (N_15838,N_15315,N_14777);
xnor U15839 (N_15839,N_15015,N_14630);
and U15840 (N_15840,N_15251,N_15518);
nand U15841 (N_15841,N_15433,N_14682);
or U15842 (N_15842,N_15128,N_15570);
or U15843 (N_15843,N_14431,N_14723);
nand U15844 (N_15844,N_14788,N_14739);
or U15845 (N_15845,N_14771,N_14846);
xor U15846 (N_15846,N_15572,N_14411);
and U15847 (N_15847,N_15030,N_14734);
or U15848 (N_15848,N_14868,N_15320);
nor U15849 (N_15849,N_15516,N_15085);
or U15850 (N_15850,N_15210,N_14637);
nand U15851 (N_15851,N_15142,N_15478);
xor U15852 (N_15852,N_14724,N_15035);
and U15853 (N_15853,N_15316,N_14469);
or U15854 (N_15854,N_14445,N_15183);
nand U15855 (N_15855,N_15525,N_15209);
xnor U15856 (N_15856,N_14783,N_15285);
and U15857 (N_15857,N_14642,N_15364);
or U15858 (N_15858,N_14549,N_14809);
and U15859 (N_15859,N_14404,N_14993);
xnor U15860 (N_15860,N_15527,N_15523);
nor U15861 (N_15861,N_15078,N_15258);
and U15862 (N_15862,N_14635,N_15452);
nor U15863 (N_15863,N_14686,N_14685);
nand U15864 (N_15864,N_15247,N_14591);
and U15865 (N_15865,N_14942,N_14920);
xor U15866 (N_15866,N_15127,N_15022);
and U15867 (N_15867,N_14463,N_15353);
nor U15868 (N_15868,N_14599,N_15261);
nor U15869 (N_15869,N_14415,N_14905);
xor U15870 (N_15870,N_15555,N_15488);
xor U15871 (N_15871,N_15381,N_15164);
nor U15872 (N_15872,N_15532,N_14945);
nand U15873 (N_15873,N_15390,N_14564);
and U15874 (N_15874,N_14443,N_15150);
xnor U15875 (N_15875,N_15466,N_15188);
or U15876 (N_15876,N_15299,N_14421);
xor U15877 (N_15877,N_14631,N_14541);
nand U15878 (N_15878,N_14436,N_14892);
nor U15879 (N_15879,N_15449,N_15438);
or U15880 (N_15880,N_14947,N_14776);
nor U15881 (N_15881,N_15557,N_14447);
xor U15882 (N_15882,N_14812,N_14829);
nand U15883 (N_15883,N_14713,N_14453);
nand U15884 (N_15884,N_14715,N_15500);
xor U15885 (N_15885,N_14749,N_14748);
nor U15886 (N_15886,N_14552,N_14806);
xnor U15887 (N_15887,N_15157,N_14581);
xor U15888 (N_15888,N_14627,N_15116);
or U15889 (N_15889,N_14704,N_14841);
and U15890 (N_15890,N_14850,N_15428);
xor U15891 (N_15891,N_14519,N_14832);
xnor U15892 (N_15892,N_15542,N_14935);
or U15893 (N_15893,N_15054,N_15105);
nor U15894 (N_15894,N_14801,N_14728);
or U15895 (N_15895,N_14833,N_14955);
xor U15896 (N_15896,N_14650,N_14533);
xnor U15897 (N_15897,N_15356,N_14667);
and U15898 (N_15898,N_14917,N_15223);
and U15899 (N_15899,N_14546,N_15277);
or U15900 (N_15900,N_14464,N_15595);
xor U15901 (N_15901,N_15059,N_15294);
nor U15902 (N_15902,N_15234,N_14513);
and U15903 (N_15903,N_15203,N_15006);
xor U15904 (N_15904,N_15473,N_15510);
and U15905 (N_15905,N_14775,N_14926);
nor U15906 (N_15906,N_14467,N_14634);
nor U15907 (N_15907,N_14698,N_14852);
xor U15908 (N_15908,N_15441,N_14786);
or U15909 (N_15909,N_15243,N_14675);
nor U15910 (N_15910,N_15307,N_14908);
xor U15911 (N_15911,N_14622,N_15079);
xor U15912 (N_15912,N_15534,N_14624);
or U15913 (N_15913,N_14554,N_14921);
xnor U15914 (N_15914,N_14975,N_15431);
nand U15915 (N_15915,N_15425,N_15181);
nand U15916 (N_15916,N_14430,N_14869);
nor U15917 (N_15917,N_14407,N_15465);
nand U15918 (N_15918,N_14600,N_14435);
or U15919 (N_15919,N_14556,N_14867);
nand U15920 (N_15920,N_14517,N_14648);
or U15921 (N_15921,N_15389,N_15357);
or U15922 (N_15922,N_15594,N_15370);
nand U15923 (N_15923,N_15266,N_14671);
xor U15924 (N_15924,N_14579,N_15149);
xnor U15925 (N_15925,N_15038,N_14784);
or U15926 (N_15926,N_14567,N_14909);
and U15927 (N_15927,N_15403,N_14480);
nor U15928 (N_15928,N_15396,N_15513);
or U15929 (N_15929,N_14896,N_14619);
nor U15930 (N_15930,N_14537,N_14988);
nor U15931 (N_15931,N_15505,N_15279);
xor U15932 (N_15932,N_14583,N_15372);
nor U15933 (N_15933,N_14466,N_14456);
nand U15934 (N_15934,N_14712,N_14821);
nand U15935 (N_15935,N_15575,N_15201);
nand U15936 (N_15936,N_15101,N_14593);
xor U15937 (N_15937,N_15386,N_15366);
and U15938 (N_15938,N_14418,N_15395);
and U15939 (N_15939,N_15593,N_15122);
xnor U15940 (N_15940,N_14475,N_14699);
nor U15941 (N_15941,N_14847,N_14597);
nand U15942 (N_15942,N_15162,N_14474);
xnor U15943 (N_15943,N_14462,N_14573);
xor U15944 (N_15944,N_15053,N_15352);
nand U15945 (N_15945,N_15067,N_14498);
nand U15946 (N_15946,N_15216,N_15124);
and U15947 (N_15947,N_14535,N_14510);
or U15948 (N_15948,N_15437,N_14457);
nand U15949 (N_15949,N_14494,N_14992);
nor U15950 (N_15950,N_14623,N_15332);
nor U15951 (N_15951,N_14618,N_14539);
nor U15952 (N_15952,N_14915,N_15213);
xor U15953 (N_15953,N_14940,N_15399);
nand U15954 (N_15954,N_14769,N_15268);
and U15955 (N_15955,N_14762,N_14763);
nand U15956 (N_15956,N_15047,N_15215);
and U15957 (N_15957,N_15063,N_15565);
nand U15958 (N_15958,N_15196,N_14870);
nand U15959 (N_15959,N_14936,N_15040);
nor U15960 (N_15960,N_15005,N_14755);
nand U15961 (N_15961,N_14628,N_15229);
xor U15962 (N_15962,N_15109,N_15130);
nand U15963 (N_15963,N_15459,N_15197);
nand U15964 (N_15964,N_15090,N_14997);
nor U15965 (N_15965,N_14835,N_14904);
nand U15966 (N_15966,N_14620,N_15221);
or U15967 (N_15967,N_15126,N_14866);
nand U15968 (N_15968,N_15144,N_15584);
xnor U15969 (N_15969,N_15271,N_15217);
or U15970 (N_15970,N_15169,N_15554);
and U15971 (N_15971,N_15363,N_14774);
and U15972 (N_15972,N_15467,N_15355);
nand U15973 (N_15973,N_15193,N_15039);
nand U15974 (N_15974,N_14670,N_14589);
and U15975 (N_15975,N_14572,N_14764);
or U15976 (N_15976,N_15301,N_15469);
and U15977 (N_15977,N_15585,N_15233);
or U15978 (N_15978,N_14796,N_15312);
or U15979 (N_15979,N_14965,N_14662);
nand U15980 (N_15980,N_15265,N_15094);
and U15981 (N_15981,N_15330,N_14543);
nand U15982 (N_15982,N_14894,N_15571);
xor U15983 (N_15983,N_15490,N_15246);
or U15984 (N_15984,N_14743,N_14931);
nand U15985 (N_15985,N_15115,N_15388);
or U15986 (N_15986,N_15461,N_14720);
or U15987 (N_15987,N_15411,N_15599);
xnor U15988 (N_15988,N_14953,N_15014);
nor U15989 (N_15989,N_14811,N_14674);
xor U15990 (N_15990,N_14679,N_15450);
nand U15991 (N_15991,N_15011,N_14605);
nand U15992 (N_15992,N_14849,N_15071);
and U15993 (N_15993,N_15168,N_15111);
nand U15994 (N_15994,N_15136,N_14890);
nor U15995 (N_15995,N_14983,N_14891);
and U15996 (N_15996,N_15380,N_14461);
nor U15997 (N_15997,N_14726,N_15347);
xor U15998 (N_15998,N_14609,N_15413);
or U15999 (N_15999,N_15019,N_14789);
nor U16000 (N_16000,N_14508,N_14924);
and U16001 (N_16001,N_14485,N_15514);
and U16002 (N_16002,N_14689,N_14895);
and U16003 (N_16003,N_14804,N_15238);
or U16004 (N_16004,N_14980,N_15447);
nor U16005 (N_16005,N_14489,N_15151);
nor U16006 (N_16006,N_15072,N_14633);
xnor U16007 (N_16007,N_15254,N_15526);
xor U16008 (N_16008,N_15507,N_14817);
nor U16009 (N_16009,N_15207,N_15073);
or U16010 (N_16010,N_14859,N_15171);
nor U16011 (N_16011,N_15158,N_14758);
nand U16012 (N_16012,N_15545,N_15581);
nand U16013 (N_16013,N_15393,N_14756);
or U16014 (N_16014,N_15237,N_15445);
and U16015 (N_16015,N_15139,N_15244);
or U16016 (N_16016,N_15423,N_14442);
nor U16017 (N_16017,N_15520,N_15065);
or U16018 (N_16018,N_14932,N_14888);
or U16019 (N_16019,N_15088,N_15117);
nor U16020 (N_16020,N_14672,N_14874);
or U16021 (N_16021,N_14823,N_15576);
and U16022 (N_16022,N_15081,N_15379);
nor U16023 (N_16023,N_14518,N_14838);
nand U16024 (N_16024,N_14614,N_14963);
or U16025 (N_16025,N_15041,N_15089);
and U16026 (N_16026,N_14858,N_15418);
or U16027 (N_16027,N_15044,N_15405);
xnor U16028 (N_16028,N_15125,N_14557);
nand U16029 (N_16029,N_14478,N_14465);
or U16030 (N_16030,N_14629,N_15198);
and U16031 (N_16031,N_14626,N_14459);
nor U16032 (N_16032,N_14412,N_15222);
xor U16033 (N_16033,N_15598,N_14741);
or U16034 (N_16034,N_15278,N_14902);
nand U16035 (N_16035,N_15057,N_14454);
and U16036 (N_16036,N_15009,N_14584);
or U16037 (N_16037,N_14470,N_15451);
nand U16038 (N_16038,N_15528,N_15424);
or U16039 (N_16039,N_15204,N_14793);
nand U16040 (N_16040,N_14566,N_15590);
xor U16041 (N_16041,N_15297,N_15121);
nor U16042 (N_16042,N_15456,N_14646);
nor U16043 (N_16043,N_15029,N_15392);
xor U16044 (N_16044,N_14727,N_15358);
xnor U16045 (N_16045,N_14949,N_14562);
nand U16046 (N_16046,N_15361,N_14884);
or U16047 (N_16047,N_15435,N_14643);
nor U16048 (N_16048,N_15430,N_15482);
or U16049 (N_16049,N_15208,N_15446);
and U16050 (N_16050,N_14954,N_14733);
or U16051 (N_16051,N_15556,N_15031);
or U16052 (N_16052,N_14578,N_14658);
or U16053 (N_16053,N_14428,N_15597);
or U16054 (N_16054,N_14644,N_15420);
xnor U16055 (N_16055,N_14632,N_14864);
xor U16056 (N_16056,N_15550,N_15367);
and U16057 (N_16057,N_15199,N_14785);
xor U16058 (N_16058,N_14912,N_15235);
nand U16059 (N_16059,N_14948,N_15415);
or U16060 (N_16060,N_15214,N_14520);
or U16061 (N_16061,N_15020,N_14738);
xnor U16062 (N_16062,N_14797,N_15427);
nand U16063 (N_16063,N_15084,N_14665);
nor U16064 (N_16064,N_14452,N_14409);
nand U16065 (N_16065,N_14587,N_15256);
and U16066 (N_16066,N_14959,N_15587);
or U16067 (N_16067,N_14880,N_14794);
and U16068 (N_16068,N_15502,N_14996);
nor U16069 (N_16069,N_15195,N_14416);
and U16070 (N_16070,N_14737,N_14827);
nand U16071 (N_16071,N_14767,N_14680);
nand U16072 (N_16072,N_14770,N_14568);
or U16073 (N_16073,N_14706,N_15519);
xor U16074 (N_16074,N_15479,N_15351);
and U16075 (N_16075,N_15417,N_15375);
and U16076 (N_16076,N_14929,N_14420);
nor U16077 (N_16077,N_15309,N_14990);
xor U16078 (N_16078,N_14757,N_15153);
and U16079 (N_16079,N_14585,N_14580);
xor U16080 (N_16080,N_14928,N_15068);
and U16081 (N_16081,N_14550,N_14683);
nor U16082 (N_16082,N_14423,N_14528);
or U16083 (N_16083,N_14889,N_15326);
nor U16084 (N_16084,N_15387,N_15263);
or U16085 (N_16085,N_14792,N_15476);
nor U16086 (N_16086,N_15232,N_14819);
xor U16087 (N_16087,N_15050,N_15422);
or U16088 (N_16088,N_15100,N_15560);
nor U16089 (N_16089,N_14592,N_15120);
nand U16090 (N_16090,N_14930,N_15453);
nor U16091 (N_16091,N_15033,N_14594);
and U16092 (N_16092,N_14944,N_14527);
nor U16093 (N_16093,N_15131,N_15026);
nand U16094 (N_16094,N_14731,N_15259);
or U16095 (N_16095,N_14719,N_15495);
nand U16096 (N_16096,N_15304,N_15359);
or U16097 (N_16097,N_14536,N_14501);
nor U16098 (N_16098,N_15242,N_14863);
nand U16099 (N_16099,N_15102,N_14781);
nor U16100 (N_16100,N_14437,N_14951);
nand U16101 (N_16101,N_14805,N_15080);
or U16102 (N_16102,N_14913,N_15145);
or U16103 (N_16103,N_15165,N_14750);
or U16104 (N_16104,N_15402,N_14814);
nand U16105 (N_16105,N_15325,N_15252);
nor U16106 (N_16106,N_14725,N_14950);
and U16107 (N_16107,N_15147,N_14677);
xor U16108 (N_16108,N_14526,N_15563);
xnor U16109 (N_16109,N_15289,N_14595);
nand U16110 (N_16110,N_14433,N_15287);
and U16111 (N_16111,N_15515,N_15002);
nand U16112 (N_16112,N_15004,N_15436);
xor U16113 (N_16113,N_14977,N_15454);
and U16114 (N_16114,N_15549,N_14807);
or U16115 (N_16115,N_14834,N_14991);
nor U16116 (N_16116,N_14525,N_14473);
nor U16117 (N_16117,N_14666,N_14652);
or U16118 (N_16118,N_15499,N_15114);
and U16119 (N_16119,N_14544,N_15314);
xnor U16120 (N_16120,N_14982,N_14410);
and U16121 (N_16121,N_14973,N_15319);
nand U16122 (N_16122,N_15175,N_15224);
nand U16123 (N_16123,N_14736,N_15383);
and U16124 (N_16124,N_14569,N_15547);
or U16125 (N_16125,N_14690,N_14897);
or U16126 (N_16126,N_15159,N_15412);
nand U16127 (N_16127,N_14857,N_15491);
nor U16128 (N_16128,N_15474,N_15434);
nor U16129 (N_16129,N_15321,N_15341);
nor U16130 (N_16130,N_15566,N_14448);
and U16131 (N_16131,N_15477,N_15013);
or U16132 (N_16132,N_14497,N_14872);
nand U16133 (N_16133,N_15172,N_15296);
nor U16134 (N_16134,N_15324,N_14987);
and U16135 (N_16135,N_15562,N_15429);
xnor U16136 (N_16136,N_14449,N_14824);
nand U16137 (N_16137,N_15286,N_15443);
xnor U16138 (N_16138,N_15135,N_14813);
nor U16139 (N_16139,N_15211,N_14721);
nand U16140 (N_16140,N_15408,N_14837);
nor U16141 (N_16141,N_14790,N_15591);
or U16142 (N_16142,N_14455,N_14752);
nand U16143 (N_16143,N_14653,N_14708);
or U16144 (N_16144,N_14702,N_14509);
nand U16145 (N_16145,N_14693,N_14688);
nor U16146 (N_16146,N_14425,N_14875);
nor U16147 (N_16147,N_14471,N_15503);
and U16148 (N_16148,N_14851,N_14434);
and U16149 (N_16149,N_14957,N_15583);
and U16150 (N_16150,N_14468,N_15371);
and U16151 (N_16151,N_15062,N_15496);
and U16152 (N_16152,N_14590,N_15093);
or U16153 (N_16153,N_15163,N_15021);
and U16154 (N_16154,N_14446,N_14574);
nor U16155 (N_16155,N_15327,N_15543);
and U16156 (N_16156,N_14507,N_14522);
nand U16157 (N_16157,N_14916,N_15318);
or U16158 (N_16158,N_15524,N_15276);
xnor U16159 (N_16159,N_15269,N_14563);
nand U16160 (N_16160,N_14883,N_14768);
nor U16161 (N_16161,N_15280,N_15070);
and U16162 (N_16162,N_15176,N_15018);
and U16163 (N_16163,N_15569,N_14538);
nor U16164 (N_16164,N_15202,N_15455);
nor U16165 (N_16165,N_15596,N_14711);
nor U16166 (N_16166,N_14500,N_15108);
and U16167 (N_16167,N_15000,N_14732);
xor U16168 (N_16168,N_14745,N_15308);
nor U16169 (N_16169,N_14511,N_14655);
and U16170 (N_16170,N_15538,N_15160);
nand U16171 (N_16171,N_14971,N_14714);
xor U16172 (N_16172,N_15492,N_14488);
xor U16173 (N_16173,N_15544,N_15200);
nand U16174 (N_16174,N_14798,N_14479);
nand U16175 (N_16175,N_14919,N_15055);
and U16176 (N_16176,N_14830,N_14918);
and U16177 (N_16177,N_15016,N_14803);
xnor U16178 (N_16178,N_14978,N_14495);
xor U16179 (N_16179,N_15350,N_14560);
or U16180 (N_16180,N_15541,N_15141);
xor U16181 (N_16181,N_15086,N_14901);
nor U16182 (N_16182,N_15134,N_14885);
nand U16183 (N_16183,N_14879,N_15339);
nand U16184 (N_16184,N_14514,N_15012);
and U16185 (N_16185,N_14534,N_14451);
and U16186 (N_16186,N_15410,N_14802);
nand U16187 (N_16187,N_15023,N_14914);
xnor U16188 (N_16188,N_15349,N_14429);
xor U16189 (N_16189,N_14871,N_14898);
nand U16190 (N_16190,N_15227,N_15336);
nand U16191 (N_16191,N_15042,N_15471);
nor U16192 (N_16192,N_15194,N_15119);
nand U16193 (N_16193,N_15586,N_14923);
xnor U16194 (N_16194,N_14651,N_14483);
nor U16195 (N_16195,N_15257,N_15472);
and U16196 (N_16196,N_14486,N_15219);
nand U16197 (N_16197,N_14922,N_14621);
xor U16198 (N_16198,N_15577,N_14484);
nand U16199 (N_16199,N_14974,N_15283);
nand U16200 (N_16200,N_14602,N_15528);
and U16201 (N_16201,N_15295,N_15529);
nand U16202 (N_16202,N_15413,N_14647);
or U16203 (N_16203,N_15495,N_15065);
nand U16204 (N_16204,N_14830,N_14890);
and U16205 (N_16205,N_15103,N_15331);
xor U16206 (N_16206,N_15514,N_15411);
nand U16207 (N_16207,N_15490,N_14565);
and U16208 (N_16208,N_14898,N_14655);
nor U16209 (N_16209,N_14667,N_15420);
nand U16210 (N_16210,N_15339,N_14400);
nand U16211 (N_16211,N_14873,N_15118);
nand U16212 (N_16212,N_15359,N_14439);
nand U16213 (N_16213,N_14812,N_15381);
nand U16214 (N_16214,N_14785,N_14653);
nand U16215 (N_16215,N_14968,N_14415);
nor U16216 (N_16216,N_14830,N_14585);
or U16217 (N_16217,N_15337,N_15392);
and U16218 (N_16218,N_15039,N_14914);
or U16219 (N_16219,N_15082,N_14513);
nand U16220 (N_16220,N_14575,N_15554);
xnor U16221 (N_16221,N_15494,N_14401);
and U16222 (N_16222,N_14739,N_14555);
and U16223 (N_16223,N_15219,N_14771);
nor U16224 (N_16224,N_14950,N_14930);
nor U16225 (N_16225,N_14454,N_14601);
nand U16226 (N_16226,N_14473,N_14953);
or U16227 (N_16227,N_15250,N_15546);
or U16228 (N_16228,N_15312,N_15126);
nor U16229 (N_16229,N_15556,N_15152);
and U16230 (N_16230,N_15519,N_15033);
nand U16231 (N_16231,N_14456,N_14501);
and U16232 (N_16232,N_14778,N_15018);
nand U16233 (N_16233,N_15394,N_15597);
xnor U16234 (N_16234,N_15595,N_14659);
or U16235 (N_16235,N_14989,N_15400);
and U16236 (N_16236,N_15013,N_15531);
or U16237 (N_16237,N_15587,N_14896);
or U16238 (N_16238,N_14848,N_14676);
nand U16239 (N_16239,N_15014,N_14724);
and U16240 (N_16240,N_15268,N_14440);
or U16241 (N_16241,N_14492,N_14503);
nor U16242 (N_16242,N_15361,N_15226);
xnor U16243 (N_16243,N_14400,N_15081);
nand U16244 (N_16244,N_15436,N_14582);
nand U16245 (N_16245,N_14850,N_15370);
or U16246 (N_16246,N_15034,N_14881);
nor U16247 (N_16247,N_14695,N_15051);
xor U16248 (N_16248,N_15324,N_15556);
nor U16249 (N_16249,N_15050,N_15073);
or U16250 (N_16250,N_15522,N_15439);
nand U16251 (N_16251,N_15320,N_15419);
or U16252 (N_16252,N_15557,N_15244);
nor U16253 (N_16253,N_14922,N_15019);
or U16254 (N_16254,N_15238,N_14486);
and U16255 (N_16255,N_14944,N_15177);
xor U16256 (N_16256,N_15465,N_15474);
nand U16257 (N_16257,N_15212,N_15248);
nor U16258 (N_16258,N_15282,N_14840);
and U16259 (N_16259,N_14614,N_15308);
or U16260 (N_16260,N_15560,N_15186);
and U16261 (N_16261,N_14511,N_14460);
and U16262 (N_16262,N_14460,N_15296);
and U16263 (N_16263,N_14999,N_15169);
nand U16264 (N_16264,N_15557,N_14979);
nor U16265 (N_16265,N_14503,N_15319);
and U16266 (N_16266,N_14968,N_14433);
or U16267 (N_16267,N_15577,N_14817);
or U16268 (N_16268,N_14944,N_14882);
xor U16269 (N_16269,N_14958,N_14409);
nor U16270 (N_16270,N_15277,N_14592);
xor U16271 (N_16271,N_14626,N_15297);
xnor U16272 (N_16272,N_15439,N_15228);
or U16273 (N_16273,N_14607,N_15251);
nand U16274 (N_16274,N_14850,N_14722);
nand U16275 (N_16275,N_14403,N_15150);
xor U16276 (N_16276,N_14979,N_15287);
nor U16277 (N_16277,N_15491,N_15373);
and U16278 (N_16278,N_14882,N_15370);
or U16279 (N_16279,N_15016,N_15061);
and U16280 (N_16280,N_14612,N_14794);
or U16281 (N_16281,N_14845,N_14792);
and U16282 (N_16282,N_15596,N_15099);
nand U16283 (N_16283,N_14529,N_15165);
nand U16284 (N_16284,N_15092,N_14420);
nand U16285 (N_16285,N_15388,N_14857);
nand U16286 (N_16286,N_14859,N_14935);
or U16287 (N_16287,N_15388,N_14545);
or U16288 (N_16288,N_14630,N_14836);
or U16289 (N_16289,N_15051,N_15527);
or U16290 (N_16290,N_14591,N_14755);
or U16291 (N_16291,N_15548,N_14746);
xor U16292 (N_16292,N_15354,N_15256);
nand U16293 (N_16293,N_14533,N_14500);
or U16294 (N_16294,N_14774,N_14542);
or U16295 (N_16295,N_14464,N_14898);
nor U16296 (N_16296,N_15348,N_15090);
nand U16297 (N_16297,N_14757,N_14905);
nand U16298 (N_16298,N_15293,N_15138);
nand U16299 (N_16299,N_15336,N_15303);
or U16300 (N_16300,N_15278,N_15161);
nand U16301 (N_16301,N_15027,N_14632);
xnor U16302 (N_16302,N_14664,N_15377);
xnor U16303 (N_16303,N_15187,N_15102);
xor U16304 (N_16304,N_14481,N_14677);
nand U16305 (N_16305,N_15124,N_15347);
and U16306 (N_16306,N_14939,N_15389);
nor U16307 (N_16307,N_15147,N_14454);
or U16308 (N_16308,N_14928,N_14894);
xnor U16309 (N_16309,N_15183,N_15180);
nand U16310 (N_16310,N_14442,N_14738);
and U16311 (N_16311,N_15008,N_15406);
nor U16312 (N_16312,N_15201,N_14980);
xnor U16313 (N_16313,N_14935,N_15399);
nand U16314 (N_16314,N_15282,N_15524);
nand U16315 (N_16315,N_14983,N_15232);
xor U16316 (N_16316,N_14845,N_14814);
xnor U16317 (N_16317,N_14414,N_15270);
and U16318 (N_16318,N_15098,N_15048);
or U16319 (N_16319,N_14873,N_15412);
xor U16320 (N_16320,N_15269,N_14670);
xnor U16321 (N_16321,N_14646,N_15246);
nor U16322 (N_16322,N_15456,N_15225);
nor U16323 (N_16323,N_15102,N_14516);
and U16324 (N_16324,N_14600,N_15423);
xnor U16325 (N_16325,N_14504,N_14965);
nand U16326 (N_16326,N_14669,N_14466);
nand U16327 (N_16327,N_15127,N_15425);
and U16328 (N_16328,N_15146,N_15186);
or U16329 (N_16329,N_14450,N_14751);
xor U16330 (N_16330,N_15220,N_15416);
and U16331 (N_16331,N_15184,N_15509);
nand U16332 (N_16332,N_14700,N_14493);
and U16333 (N_16333,N_14964,N_15507);
or U16334 (N_16334,N_14738,N_14638);
nor U16335 (N_16335,N_15010,N_14923);
xor U16336 (N_16336,N_14500,N_14972);
nand U16337 (N_16337,N_15462,N_15381);
xnor U16338 (N_16338,N_15573,N_15399);
and U16339 (N_16339,N_14681,N_15559);
nand U16340 (N_16340,N_15064,N_15390);
nand U16341 (N_16341,N_14807,N_15018);
and U16342 (N_16342,N_15189,N_14417);
nor U16343 (N_16343,N_15587,N_15484);
and U16344 (N_16344,N_14489,N_15090);
xnor U16345 (N_16345,N_15443,N_14534);
and U16346 (N_16346,N_15146,N_14644);
nor U16347 (N_16347,N_14657,N_15145);
or U16348 (N_16348,N_15448,N_14717);
nand U16349 (N_16349,N_14949,N_14778);
nand U16350 (N_16350,N_15132,N_14716);
or U16351 (N_16351,N_14592,N_14928);
nor U16352 (N_16352,N_14845,N_15140);
nand U16353 (N_16353,N_14457,N_15116);
nor U16354 (N_16354,N_15068,N_15066);
or U16355 (N_16355,N_15176,N_15189);
nor U16356 (N_16356,N_14996,N_14836);
nor U16357 (N_16357,N_14444,N_14963);
or U16358 (N_16358,N_14676,N_15395);
nor U16359 (N_16359,N_15313,N_14809);
nand U16360 (N_16360,N_14646,N_14574);
or U16361 (N_16361,N_15585,N_15490);
and U16362 (N_16362,N_15350,N_15066);
nor U16363 (N_16363,N_14937,N_14429);
and U16364 (N_16364,N_15162,N_14867);
xor U16365 (N_16365,N_15326,N_15192);
nand U16366 (N_16366,N_15203,N_15478);
nor U16367 (N_16367,N_14815,N_14640);
or U16368 (N_16368,N_14480,N_14573);
xnor U16369 (N_16369,N_15566,N_14626);
or U16370 (N_16370,N_15113,N_15307);
nand U16371 (N_16371,N_14997,N_14428);
nand U16372 (N_16372,N_15520,N_14675);
nand U16373 (N_16373,N_14870,N_14569);
or U16374 (N_16374,N_15360,N_15415);
nor U16375 (N_16375,N_14774,N_14752);
or U16376 (N_16376,N_14938,N_15017);
nor U16377 (N_16377,N_14582,N_15239);
or U16378 (N_16378,N_14408,N_14849);
and U16379 (N_16379,N_15066,N_15061);
or U16380 (N_16380,N_15157,N_15050);
nor U16381 (N_16381,N_14489,N_14712);
and U16382 (N_16382,N_14906,N_15184);
nor U16383 (N_16383,N_15126,N_15415);
nand U16384 (N_16384,N_14558,N_15006);
and U16385 (N_16385,N_14562,N_14420);
nand U16386 (N_16386,N_15019,N_14710);
nor U16387 (N_16387,N_14688,N_14813);
nand U16388 (N_16388,N_15405,N_14456);
nor U16389 (N_16389,N_14695,N_15421);
or U16390 (N_16390,N_14411,N_14908);
xnor U16391 (N_16391,N_14724,N_14602);
nor U16392 (N_16392,N_14999,N_14660);
and U16393 (N_16393,N_14647,N_14429);
xor U16394 (N_16394,N_14637,N_14486);
or U16395 (N_16395,N_14783,N_14776);
and U16396 (N_16396,N_15561,N_15178);
and U16397 (N_16397,N_15105,N_14602);
and U16398 (N_16398,N_15313,N_14822);
nor U16399 (N_16399,N_14588,N_14433);
xnor U16400 (N_16400,N_14883,N_14690);
nand U16401 (N_16401,N_15512,N_15156);
nand U16402 (N_16402,N_15249,N_15096);
and U16403 (N_16403,N_14880,N_14949);
nand U16404 (N_16404,N_14589,N_14970);
nand U16405 (N_16405,N_15428,N_15287);
xnor U16406 (N_16406,N_15546,N_14915);
nand U16407 (N_16407,N_14746,N_15408);
xnor U16408 (N_16408,N_15396,N_15479);
and U16409 (N_16409,N_15134,N_15452);
xor U16410 (N_16410,N_15005,N_14617);
nor U16411 (N_16411,N_14874,N_15247);
and U16412 (N_16412,N_15391,N_15054);
nor U16413 (N_16413,N_15284,N_15582);
or U16414 (N_16414,N_14403,N_15585);
or U16415 (N_16415,N_14919,N_15554);
xor U16416 (N_16416,N_15594,N_14885);
nand U16417 (N_16417,N_15122,N_14518);
nor U16418 (N_16418,N_14592,N_15115);
or U16419 (N_16419,N_15207,N_15149);
nand U16420 (N_16420,N_14811,N_14559);
and U16421 (N_16421,N_14807,N_15216);
xor U16422 (N_16422,N_14483,N_14997);
xnor U16423 (N_16423,N_15222,N_15082);
xnor U16424 (N_16424,N_14697,N_15272);
nor U16425 (N_16425,N_15506,N_14747);
or U16426 (N_16426,N_14948,N_14642);
or U16427 (N_16427,N_14791,N_15129);
nor U16428 (N_16428,N_15289,N_14995);
nor U16429 (N_16429,N_15009,N_14667);
and U16430 (N_16430,N_14823,N_14618);
nand U16431 (N_16431,N_14988,N_14540);
nor U16432 (N_16432,N_15370,N_14870);
xnor U16433 (N_16433,N_14558,N_15514);
nor U16434 (N_16434,N_14448,N_14914);
and U16435 (N_16435,N_15591,N_15192);
or U16436 (N_16436,N_14475,N_14756);
and U16437 (N_16437,N_15167,N_14580);
and U16438 (N_16438,N_15544,N_15527);
nor U16439 (N_16439,N_14606,N_14967);
xnor U16440 (N_16440,N_14880,N_15381);
nor U16441 (N_16441,N_15171,N_14990);
xnor U16442 (N_16442,N_15015,N_15037);
and U16443 (N_16443,N_14701,N_14876);
nand U16444 (N_16444,N_14856,N_15339);
xnor U16445 (N_16445,N_15101,N_15015);
xor U16446 (N_16446,N_15166,N_15058);
or U16447 (N_16447,N_15203,N_15556);
xor U16448 (N_16448,N_14588,N_15243);
xnor U16449 (N_16449,N_15391,N_14507);
and U16450 (N_16450,N_14491,N_14967);
and U16451 (N_16451,N_15176,N_15041);
nand U16452 (N_16452,N_15120,N_15385);
and U16453 (N_16453,N_14509,N_15146);
xor U16454 (N_16454,N_14905,N_15593);
nor U16455 (N_16455,N_14827,N_14847);
xor U16456 (N_16456,N_15511,N_15587);
nor U16457 (N_16457,N_14735,N_14723);
or U16458 (N_16458,N_14530,N_15441);
nand U16459 (N_16459,N_15182,N_15585);
nor U16460 (N_16460,N_14764,N_14760);
or U16461 (N_16461,N_15560,N_15273);
nor U16462 (N_16462,N_15091,N_14675);
nand U16463 (N_16463,N_15490,N_15429);
nor U16464 (N_16464,N_15280,N_15091);
xnor U16465 (N_16465,N_14491,N_14785);
nor U16466 (N_16466,N_14525,N_14432);
xor U16467 (N_16467,N_14637,N_14830);
and U16468 (N_16468,N_15252,N_14837);
and U16469 (N_16469,N_14656,N_14676);
nor U16470 (N_16470,N_15228,N_15096);
and U16471 (N_16471,N_15239,N_15476);
nand U16472 (N_16472,N_14773,N_14530);
nand U16473 (N_16473,N_14407,N_14470);
or U16474 (N_16474,N_14551,N_15263);
and U16475 (N_16475,N_14765,N_15026);
nand U16476 (N_16476,N_14637,N_15275);
nor U16477 (N_16477,N_14635,N_14407);
xnor U16478 (N_16478,N_15581,N_14542);
and U16479 (N_16479,N_15531,N_14441);
nand U16480 (N_16480,N_15046,N_14826);
and U16481 (N_16481,N_14939,N_14433);
nand U16482 (N_16482,N_14921,N_15448);
nand U16483 (N_16483,N_15363,N_15103);
xor U16484 (N_16484,N_14846,N_15222);
or U16485 (N_16485,N_14859,N_15544);
or U16486 (N_16486,N_15032,N_14850);
or U16487 (N_16487,N_14510,N_15420);
or U16488 (N_16488,N_15132,N_15000);
and U16489 (N_16489,N_15195,N_15465);
and U16490 (N_16490,N_15344,N_15137);
and U16491 (N_16491,N_15010,N_15595);
or U16492 (N_16492,N_15040,N_15093);
and U16493 (N_16493,N_14558,N_14633);
or U16494 (N_16494,N_15029,N_15490);
or U16495 (N_16495,N_15344,N_15143);
nor U16496 (N_16496,N_15247,N_14937);
or U16497 (N_16497,N_14954,N_15449);
xnor U16498 (N_16498,N_15325,N_14519);
and U16499 (N_16499,N_15446,N_15309);
nand U16500 (N_16500,N_15371,N_15245);
or U16501 (N_16501,N_14517,N_14785);
and U16502 (N_16502,N_14608,N_15228);
nor U16503 (N_16503,N_14576,N_14824);
and U16504 (N_16504,N_15509,N_15268);
or U16505 (N_16505,N_15407,N_14599);
and U16506 (N_16506,N_14564,N_14524);
or U16507 (N_16507,N_15027,N_14980);
nand U16508 (N_16508,N_15426,N_14736);
nand U16509 (N_16509,N_15523,N_14902);
and U16510 (N_16510,N_14897,N_14460);
nor U16511 (N_16511,N_14913,N_14543);
xnor U16512 (N_16512,N_14575,N_14573);
xor U16513 (N_16513,N_14424,N_14683);
nor U16514 (N_16514,N_14519,N_14898);
or U16515 (N_16515,N_15502,N_15395);
nand U16516 (N_16516,N_14613,N_15367);
nor U16517 (N_16517,N_15295,N_14745);
xor U16518 (N_16518,N_15406,N_14992);
xnor U16519 (N_16519,N_15390,N_15038);
nand U16520 (N_16520,N_14540,N_14984);
or U16521 (N_16521,N_14612,N_15566);
nor U16522 (N_16522,N_15356,N_14476);
or U16523 (N_16523,N_15475,N_15590);
nor U16524 (N_16524,N_15454,N_14555);
nor U16525 (N_16525,N_15069,N_14922);
or U16526 (N_16526,N_15257,N_15246);
xor U16527 (N_16527,N_15171,N_14965);
or U16528 (N_16528,N_14569,N_15402);
xnor U16529 (N_16529,N_15304,N_14651);
xnor U16530 (N_16530,N_14971,N_15425);
nand U16531 (N_16531,N_14821,N_15260);
or U16532 (N_16532,N_15077,N_15215);
and U16533 (N_16533,N_15170,N_14488);
nand U16534 (N_16534,N_15224,N_15440);
xor U16535 (N_16535,N_14757,N_14823);
nor U16536 (N_16536,N_15186,N_15283);
nand U16537 (N_16537,N_15308,N_15508);
and U16538 (N_16538,N_14453,N_14972);
xor U16539 (N_16539,N_14411,N_15157);
nor U16540 (N_16540,N_15592,N_14998);
xnor U16541 (N_16541,N_15027,N_14818);
nor U16542 (N_16542,N_14627,N_14664);
xnor U16543 (N_16543,N_15544,N_15573);
nor U16544 (N_16544,N_15109,N_14930);
nand U16545 (N_16545,N_14847,N_14510);
and U16546 (N_16546,N_15025,N_14961);
nor U16547 (N_16547,N_15403,N_14934);
or U16548 (N_16548,N_15423,N_14687);
nand U16549 (N_16549,N_14614,N_15343);
and U16550 (N_16550,N_15027,N_14410);
nand U16551 (N_16551,N_14784,N_15123);
and U16552 (N_16552,N_14906,N_15588);
xnor U16553 (N_16553,N_14737,N_15478);
and U16554 (N_16554,N_14522,N_15375);
xnor U16555 (N_16555,N_15187,N_14495);
nand U16556 (N_16556,N_14578,N_14442);
nor U16557 (N_16557,N_15057,N_15020);
and U16558 (N_16558,N_15354,N_15195);
and U16559 (N_16559,N_15323,N_15043);
xnor U16560 (N_16560,N_15319,N_15479);
nor U16561 (N_16561,N_14858,N_15169);
nor U16562 (N_16562,N_14897,N_14515);
or U16563 (N_16563,N_14758,N_15554);
nor U16564 (N_16564,N_15178,N_15045);
nand U16565 (N_16565,N_15272,N_14707);
nand U16566 (N_16566,N_15460,N_15119);
xor U16567 (N_16567,N_15123,N_14437);
or U16568 (N_16568,N_15326,N_14490);
xor U16569 (N_16569,N_14888,N_14815);
or U16570 (N_16570,N_15336,N_15447);
nand U16571 (N_16571,N_15300,N_15193);
nor U16572 (N_16572,N_15540,N_14637);
nand U16573 (N_16573,N_14615,N_15095);
or U16574 (N_16574,N_15063,N_14926);
xor U16575 (N_16575,N_14567,N_15506);
or U16576 (N_16576,N_15041,N_14556);
nor U16577 (N_16577,N_14710,N_15282);
nor U16578 (N_16578,N_14938,N_15590);
xnor U16579 (N_16579,N_15386,N_14521);
nand U16580 (N_16580,N_14618,N_14734);
xor U16581 (N_16581,N_14592,N_14690);
or U16582 (N_16582,N_15028,N_15380);
nor U16583 (N_16583,N_14820,N_15168);
nor U16584 (N_16584,N_14889,N_15290);
or U16585 (N_16585,N_15458,N_15203);
or U16586 (N_16586,N_14556,N_14887);
and U16587 (N_16587,N_15597,N_14767);
and U16588 (N_16588,N_14470,N_15244);
nor U16589 (N_16589,N_14456,N_15537);
nor U16590 (N_16590,N_14824,N_15204);
xor U16591 (N_16591,N_15541,N_14981);
xor U16592 (N_16592,N_15421,N_14933);
and U16593 (N_16593,N_15131,N_14816);
and U16594 (N_16594,N_15579,N_14991);
xor U16595 (N_16595,N_15295,N_14746);
or U16596 (N_16596,N_15424,N_15270);
xor U16597 (N_16597,N_14748,N_15181);
nand U16598 (N_16598,N_14688,N_15355);
nand U16599 (N_16599,N_14401,N_15344);
nand U16600 (N_16600,N_14655,N_15319);
xnor U16601 (N_16601,N_14615,N_14814);
xor U16602 (N_16602,N_14620,N_14600);
nor U16603 (N_16603,N_14808,N_14940);
nor U16604 (N_16604,N_15402,N_15082);
or U16605 (N_16605,N_14654,N_15282);
or U16606 (N_16606,N_14723,N_14958);
and U16607 (N_16607,N_15027,N_14415);
xnor U16608 (N_16608,N_14972,N_14471);
xor U16609 (N_16609,N_15212,N_15041);
nand U16610 (N_16610,N_15514,N_14835);
xnor U16611 (N_16611,N_15445,N_14785);
nor U16612 (N_16612,N_15576,N_14939);
or U16613 (N_16613,N_14587,N_14900);
nor U16614 (N_16614,N_14906,N_15445);
or U16615 (N_16615,N_14701,N_14592);
or U16616 (N_16616,N_14872,N_15245);
nor U16617 (N_16617,N_15479,N_15362);
or U16618 (N_16618,N_15340,N_14767);
xor U16619 (N_16619,N_14736,N_14556);
and U16620 (N_16620,N_15318,N_14660);
nor U16621 (N_16621,N_14461,N_14893);
and U16622 (N_16622,N_14494,N_15546);
nor U16623 (N_16623,N_14448,N_15383);
or U16624 (N_16624,N_15356,N_15338);
and U16625 (N_16625,N_15142,N_14907);
or U16626 (N_16626,N_14805,N_14657);
or U16627 (N_16627,N_14874,N_15598);
or U16628 (N_16628,N_15030,N_14691);
or U16629 (N_16629,N_14781,N_15217);
nor U16630 (N_16630,N_15157,N_15237);
xnor U16631 (N_16631,N_14716,N_15033);
or U16632 (N_16632,N_14700,N_14943);
and U16633 (N_16633,N_14970,N_14866);
and U16634 (N_16634,N_14689,N_14433);
and U16635 (N_16635,N_14681,N_15075);
xor U16636 (N_16636,N_14884,N_14960);
nor U16637 (N_16637,N_15218,N_14723);
xnor U16638 (N_16638,N_15511,N_14916);
and U16639 (N_16639,N_14619,N_14522);
or U16640 (N_16640,N_14979,N_14672);
and U16641 (N_16641,N_15566,N_15131);
xnor U16642 (N_16642,N_15176,N_14787);
nand U16643 (N_16643,N_14608,N_14878);
or U16644 (N_16644,N_15352,N_15149);
or U16645 (N_16645,N_15519,N_15339);
nand U16646 (N_16646,N_15393,N_15223);
and U16647 (N_16647,N_14666,N_15002);
and U16648 (N_16648,N_15387,N_15316);
nand U16649 (N_16649,N_14616,N_14641);
and U16650 (N_16650,N_15043,N_15574);
or U16651 (N_16651,N_15088,N_14985);
and U16652 (N_16652,N_14489,N_14456);
and U16653 (N_16653,N_14771,N_14639);
xnor U16654 (N_16654,N_14576,N_15471);
xnor U16655 (N_16655,N_14939,N_15217);
or U16656 (N_16656,N_14677,N_15514);
nor U16657 (N_16657,N_14459,N_14737);
nand U16658 (N_16658,N_14791,N_14930);
or U16659 (N_16659,N_15386,N_14873);
xor U16660 (N_16660,N_14831,N_14627);
nor U16661 (N_16661,N_14881,N_15109);
and U16662 (N_16662,N_15499,N_14717);
or U16663 (N_16663,N_14814,N_15063);
or U16664 (N_16664,N_14861,N_15246);
nand U16665 (N_16665,N_15174,N_15402);
xnor U16666 (N_16666,N_15403,N_15227);
xnor U16667 (N_16667,N_14863,N_14834);
nor U16668 (N_16668,N_14956,N_15416);
nor U16669 (N_16669,N_15107,N_14885);
xnor U16670 (N_16670,N_15382,N_15565);
and U16671 (N_16671,N_15388,N_15298);
nor U16672 (N_16672,N_14970,N_15193);
and U16673 (N_16673,N_15165,N_14966);
or U16674 (N_16674,N_15594,N_15035);
and U16675 (N_16675,N_15301,N_14601);
and U16676 (N_16676,N_14407,N_14488);
xnor U16677 (N_16677,N_14971,N_14405);
xor U16678 (N_16678,N_15467,N_15212);
nand U16679 (N_16679,N_14455,N_14579);
xnor U16680 (N_16680,N_14798,N_14413);
and U16681 (N_16681,N_15267,N_15433);
nor U16682 (N_16682,N_15521,N_15028);
nor U16683 (N_16683,N_15061,N_14775);
nand U16684 (N_16684,N_15203,N_15360);
and U16685 (N_16685,N_14540,N_14512);
and U16686 (N_16686,N_14796,N_14504);
and U16687 (N_16687,N_14708,N_14468);
nand U16688 (N_16688,N_14701,N_14603);
xor U16689 (N_16689,N_14835,N_15313);
nor U16690 (N_16690,N_15455,N_15512);
nor U16691 (N_16691,N_15427,N_14694);
or U16692 (N_16692,N_15237,N_15330);
nor U16693 (N_16693,N_14491,N_15139);
xor U16694 (N_16694,N_14525,N_15065);
or U16695 (N_16695,N_15328,N_15065);
nand U16696 (N_16696,N_15120,N_15051);
nor U16697 (N_16697,N_14691,N_14835);
nand U16698 (N_16698,N_14851,N_15085);
or U16699 (N_16699,N_14854,N_14838);
or U16700 (N_16700,N_14542,N_14714);
nor U16701 (N_16701,N_15030,N_14824);
or U16702 (N_16702,N_14505,N_14616);
and U16703 (N_16703,N_14915,N_15457);
or U16704 (N_16704,N_15533,N_15567);
and U16705 (N_16705,N_14997,N_15505);
and U16706 (N_16706,N_14472,N_14682);
or U16707 (N_16707,N_14437,N_15141);
xor U16708 (N_16708,N_14447,N_14746);
nand U16709 (N_16709,N_14697,N_15164);
nand U16710 (N_16710,N_15525,N_15219);
xnor U16711 (N_16711,N_15340,N_14979);
nand U16712 (N_16712,N_14822,N_14508);
or U16713 (N_16713,N_14809,N_14997);
nor U16714 (N_16714,N_15463,N_14436);
nand U16715 (N_16715,N_15526,N_15432);
nand U16716 (N_16716,N_15545,N_15293);
and U16717 (N_16717,N_15276,N_15235);
or U16718 (N_16718,N_15347,N_15033);
nor U16719 (N_16719,N_14767,N_14973);
xor U16720 (N_16720,N_15480,N_15308);
xnor U16721 (N_16721,N_15128,N_15586);
or U16722 (N_16722,N_14565,N_15516);
and U16723 (N_16723,N_15329,N_15225);
nand U16724 (N_16724,N_15159,N_15076);
and U16725 (N_16725,N_15452,N_15508);
xnor U16726 (N_16726,N_15205,N_14963);
or U16727 (N_16727,N_14876,N_15436);
xor U16728 (N_16728,N_15506,N_15423);
and U16729 (N_16729,N_14541,N_14860);
nand U16730 (N_16730,N_15514,N_14658);
or U16731 (N_16731,N_15494,N_15358);
and U16732 (N_16732,N_15019,N_15450);
xnor U16733 (N_16733,N_15197,N_14747);
xor U16734 (N_16734,N_14966,N_15535);
and U16735 (N_16735,N_15019,N_14909);
or U16736 (N_16736,N_14497,N_14960);
or U16737 (N_16737,N_14509,N_15578);
or U16738 (N_16738,N_14521,N_14717);
and U16739 (N_16739,N_14430,N_14665);
nor U16740 (N_16740,N_15587,N_14895);
nor U16741 (N_16741,N_14586,N_15331);
xor U16742 (N_16742,N_14530,N_15210);
xnor U16743 (N_16743,N_14749,N_14619);
nand U16744 (N_16744,N_15436,N_15560);
or U16745 (N_16745,N_15004,N_14695);
and U16746 (N_16746,N_15493,N_15535);
xor U16747 (N_16747,N_14891,N_15450);
and U16748 (N_16748,N_15011,N_14967);
nand U16749 (N_16749,N_14623,N_14402);
nor U16750 (N_16750,N_14916,N_15018);
nand U16751 (N_16751,N_14815,N_15562);
xor U16752 (N_16752,N_14969,N_14700);
or U16753 (N_16753,N_14554,N_15549);
xor U16754 (N_16754,N_15545,N_14951);
nor U16755 (N_16755,N_15544,N_15354);
xnor U16756 (N_16756,N_14671,N_15582);
nor U16757 (N_16757,N_14548,N_14605);
xor U16758 (N_16758,N_15128,N_14921);
or U16759 (N_16759,N_14803,N_14564);
xor U16760 (N_16760,N_15321,N_14670);
or U16761 (N_16761,N_14404,N_14850);
and U16762 (N_16762,N_15128,N_15113);
and U16763 (N_16763,N_14781,N_15377);
or U16764 (N_16764,N_15374,N_14947);
nand U16765 (N_16765,N_15223,N_15020);
and U16766 (N_16766,N_14686,N_14665);
and U16767 (N_16767,N_14722,N_15321);
or U16768 (N_16768,N_14620,N_14454);
nor U16769 (N_16769,N_14673,N_15406);
xor U16770 (N_16770,N_15500,N_14550);
and U16771 (N_16771,N_15172,N_15322);
and U16772 (N_16772,N_15340,N_15146);
or U16773 (N_16773,N_15572,N_14410);
nor U16774 (N_16774,N_15510,N_14843);
xnor U16775 (N_16775,N_15400,N_14871);
nand U16776 (N_16776,N_14822,N_15425);
nor U16777 (N_16777,N_14988,N_14499);
nor U16778 (N_16778,N_14445,N_15330);
or U16779 (N_16779,N_15023,N_14966);
and U16780 (N_16780,N_14659,N_14893);
xnor U16781 (N_16781,N_14967,N_14814);
xnor U16782 (N_16782,N_14793,N_14556);
or U16783 (N_16783,N_15100,N_15447);
and U16784 (N_16784,N_15570,N_14546);
or U16785 (N_16785,N_15444,N_14524);
nand U16786 (N_16786,N_15396,N_15578);
or U16787 (N_16787,N_15262,N_14661);
nand U16788 (N_16788,N_15135,N_14655);
nand U16789 (N_16789,N_15039,N_14928);
and U16790 (N_16790,N_14411,N_15319);
nor U16791 (N_16791,N_15044,N_14998);
and U16792 (N_16792,N_14801,N_15186);
or U16793 (N_16793,N_14584,N_15337);
or U16794 (N_16794,N_14926,N_14626);
and U16795 (N_16795,N_14637,N_15048);
xor U16796 (N_16796,N_15440,N_15199);
and U16797 (N_16797,N_15431,N_15089);
nand U16798 (N_16798,N_15360,N_14557);
or U16799 (N_16799,N_15533,N_15544);
and U16800 (N_16800,N_16445,N_15768);
xnor U16801 (N_16801,N_15608,N_16170);
and U16802 (N_16802,N_16252,N_16706);
and U16803 (N_16803,N_16021,N_16485);
nor U16804 (N_16804,N_15615,N_16773);
and U16805 (N_16805,N_16640,N_16369);
and U16806 (N_16806,N_15761,N_15917);
nor U16807 (N_16807,N_16226,N_15728);
and U16808 (N_16808,N_15907,N_16276);
nand U16809 (N_16809,N_16266,N_15685);
nand U16810 (N_16810,N_16623,N_16158);
and U16811 (N_16811,N_15625,N_15734);
or U16812 (N_16812,N_15683,N_16253);
nor U16813 (N_16813,N_16559,N_16557);
or U16814 (N_16814,N_16499,N_15966);
or U16815 (N_16815,N_16663,N_16272);
nand U16816 (N_16816,N_16182,N_16138);
xnor U16817 (N_16817,N_16674,N_15813);
and U16818 (N_16818,N_16354,N_15969);
or U16819 (N_16819,N_15717,N_15808);
nor U16820 (N_16820,N_16651,N_16704);
xor U16821 (N_16821,N_15864,N_15601);
or U16822 (N_16822,N_15949,N_15933);
and U16823 (N_16823,N_16524,N_16289);
nand U16824 (N_16824,N_16782,N_15991);
or U16825 (N_16825,N_16144,N_16028);
xnor U16826 (N_16826,N_15779,N_16145);
and U16827 (N_16827,N_16468,N_15684);
nand U16828 (N_16828,N_15651,N_15707);
or U16829 (N_16829,N_15981,N_16480);
and U16830 (N_16830,N_15918,N_16127);
nand U16831 (N_16831,N_16373,N_15692);
nand U16832 (N_16832,N_15843,N_16408);
nor U16833 (N_16833,N_16049,N_15983);
or U16834 (N_16834,N_15993,N_15944);
and U16835 (N_16835,N_16300,N_16361);
xor U16836 (N_16836,N_16549,N_16647);
or U16837 (N_16837,N_16722,N_15925);
or U16838 (N_16838,N_16515,N_15657);
and U16839 (N_16839,N_16626,N_16173);
or U16840 (N_16840,N_16481,N_16619);
xnor U16841 (N_16841,N_16379,N_15787);
nand U16842 (N_16842,N_15622,N_15614);
and U16843 (N_16843,N_16677,N_16032);
or U16844 (N_16844,N_16727,N_15992);
xnor U16845 (N_16845,N_16255,N_15904);
or U16846 (N_16846,N_15617,N_16737);
nor U16847 (N_16847,N_15816,N_16080);
and U16848 (N_16848,N_15915,N_15901);
nor U16849 (N_16849,N_15961,N_15940);
xor U16850 (N_16850,N_16458,N_16486);
xnor U16851 (N_16851,N_15696,N_16537);
xnor U16852 (N_16852,N_16746,N_16405);
or U16853 (N_16853,N_16420,N_16086);
and U16854 (N_16854,N_15935,N_15871);
or U16855 (N_16855,N_16579,N_16281);
or U16856 (N_16856,N_15912,N_16271);
or U16857 (N_16857,N_15656,N_16261);
xor U16858 (N_16858,N_16510,N_16417);
or U16859 (N_16859,N_16701,N_15667);
and U16860 (N_16860,N_15703,N_16358);
nand U16861 (N_16861,N_16694,N_16375);
and U16862 (N_16862,N_16406,N_16464);
xnor U16863 (N_16863,N_16079,N_15633);
and U16864 (N_16864,N_16196,N_16284);
nand U16865 (N_16865,N_16713,N_16344);
or U16866 (N_16866,N_15611,N_16539);
or U16867 (N_16867,N_15788,N_16584);
or U16868 (N_16868,N_16120,N_16421);
nand U16869 (N_16869,N_16591,N_15932);
or U16870 (N_16870,N_16229,N_16195);
xnor U16871 (N_16871,N_15950,N_16243);
and U16872 (N_16872,N_15835,N_16102);
and U16873 (N_16873,N_15664,N_15756);
xnor U16874 (N_16874,N_16787,N_16556);
and U16875 (N_16875,N_16317,N_16491);
nor U16876 (N_16876,N_15892,N_16301);
and U16877 (N_16877,N_16180,N_16561);
xnor U16878 (N_16878,N_16767,N_16149);
and U16879 (N_16879,N_15934,N_16048);
and U16880 (N_16880,N_15709,N_16413);
nor U16881 (N_16881,N_16328,N_15609);
nand U16882 (N_16882,N_15905,N_16497);
nand U16883 (N_16883,N_16137,N_16741);
or U16884 (N_16884,N_16297,N_16026);
xor U16885 (N_16885,N_16702,N_16568);
xor U16886 (N_16886,N_15706,N_16207);
xnor U16887 (N_16887,N_16681,N_15930);
xnor U16888 (N_16888,N_16334,N_16431);
xnor U16889 (N_16889,N_16618,N_15699);
nand U16890 (N_16890,N_15986,N_16685);
nor U16891 (N_16891,N_16365,N_16296);
or U16892 (N_16892,N_16501,N_16397);
or U16893 (N_16893,N_16633,N_16477);
nand U16894 (N_16894,N_16454,N_15749);
and U16895 (N_16895,N_16130,N_16277);
nor U16896 (N_16896,N_16081,N_16331);
xnor U16897 (N_16897,N_15919,N_16747);
nor U16898 (N_16898,N_16402,N_16333);
nand U16899 (N_16899,N_15739,N_16189);
or U16900 (N_16900,N_15795,N_16059);
nand U16901 (N_16901,N_16472,N_15896);
nand U16902 (N_16902,N_16245,N_16583);
nor U16903 (N_16903,N_15790,N_16469);
nor U16904 (N_16904,N_16363,N_16439);
nand U16905 (N_16905,N_16309,N_16199);
and U16906 (N_16906,N_16325,N_15635);
or U16907 (N_16907,N_16033,N_16001);
xnor U16908 (N_16908,N_16605,N_15658);
or U16909 (N_16909,N_16471,N_16490);
nand U16910 (N_16910,N_16603,N_16257);
or U16911 (N_16911,N_16070,N_16311);
or U16912 (N_16912,N_16762,N_16686);
nor U16913 (N_16913,N_15946,N_16526);
nor U16914 (N_16914,N_16629,N_16225);
nor U16915 (N_16915,N_15829,N_16565);
nor U16916 (N_16916,N_16576,N_16153);
or U16917 (N_16917,N_16476,N_16724);
and U16918 (N_16918,N_16030,N_16745);
and U16919 (N_16919,N_15920,N_15888);
nand U16920 (N_16920,N_16505,N_16409);
nand U16921 (N_16921,N_16139,N_15856);
and U16922 (N_16922,N_16768,N_16577);
nor U16923 (N_16923,N_16793,N_16422);
and U16924 (N_16924,N_15724,N_15807);
nand U16925 (N_16925,N_16212,N_16097);
xnor U16926 (N_16926,N_16438,N_16661);
nand U16927 (N_16927,N_15840,N_16588);
nand U16928 (N_16928,N_16269,N_16073);
nor U16929 (N_16929,N_16209,N_16185);
or U16930 (N_16930,N_16792,N_16174);
xnor U16931 (N_16931,N_15889,N_16446);
nand U16932 (N_16932,N_16135,N_15841);
or U16933 (N_16933,N_16660,N_16087);
and U16934 (N_16934,N_16104,N_15883);
nor U16935 (N_16935,N_16377,N_15603);
or U16936 (N_16936,N_15942,N_16432);
xor U16937 (N_16937,N_16419,N_16456);
xnor U16938 (N_16938,N_16532,N_16460);
nand U16939 (N_16939,N_16649,N_16543);
nand U16940 (N_16940,N_16718,N_16278);
nand U16941 (N_16941,N_16042,N_15887);
and U16942 (N_16942,N_16453,N_15859);
nand U16943 (N_16943,N_16436,N_16098);
and U16944 (N_16944,N_16125,N_16089);
nor U16945 (N_16945,N_16769,N_15763);
nor U16946 (N_16946,N_16115,N_16766);
xnor U16947 (N_16947,N_16750,N_15774);
nor U16948 (N_16948,N_15792,N_16239);
nor U16949 (N_16949,N_16017,N_16298);
or U16950 (N_16950,N_16063,N_16217);
nand U16951 (N_16951,N_15827,N_16085);
nor U16952 (N_16952,N_15860,N_15936);
or U16953 (N_16953,N_16128,N_16250);
nand U16954 (N_16954,N_15722,N_16614);
and U16955 (N_16955,N_16423,N_15893);
xor U16956 (N_16956,N_15955,N_16323);
nor U16957 (N_16957,N_16178,N_16279);
nor U16958 (N_16958,N_15804,N_16611);
xnor U16959 (N_16959,N_16644,N_16562);
xor U16960 (N_16960,N_16554,N_16440);
nor U16961 (N_16961,N_15967,N_16601);
and U16962 (N_16962,N_16659,N_16000);
nand U16963 (N_16963,N_16112,N_15778);
nor U16964 (N_16964,N_16005,N_16610);
or U16965 (N_16965,N_16014,N_16292);
nor U16966 (N_16966,N_15680,N_15838);
and U16967 (N_16967,N_16634,N_15604);
or U16968 (N_16968,N_16581,N_15988);
xor U16969 (N_16969,N_15819,N_16188);
nand U16970 (N_16970,N_16072,N_16461);
xnor U16971 (N_16971,N_16675,N_15874);
nor U16972 (N_16972,N_16056,N_15947);
or U16973 (N_16973,N_16078,N_16721);
and U16974 (N_16974,N_16639,N_15861);
and U16975 (N_16975,N_15708,N_16381);
nand U16976 (N_16976,N_15714,N_16183);
nor U16977 (N_16977,N_16224,N_16343);
xnor U16978 (N_16978,N_16606,N_16484);
or U16979 (N_16979,N_16513,N_15785);
nand U16980 (N_16980,N_16564,N_16667);
and U16981 (N_16981,N_16683,N_15948);
xor U16982 (N_16982,N_16003,N_15953);
nand U16983 (N_16983,N_16506,N_16441);
xnor U16984 (N_16984,N_15814,N_16372);
or U16985 (N_16985,N_16617,N_16038);
nand U16986 (N_16986,N_16470,N_15784);
nand U16987 (N_16987,N_16206,N_16449);
nor U16988 (N_16988,N_16107,N_16155);
and U16989 (N_16989,N_15849,N_16430);
nand U16990 (N_16990,N_16246,N_15994);
nand U16991 (N_16991,N_15830,N_15735);
nor U16992 (N_16992,N_15914,N_16540);
or U16993 (N_16993,N_15738,N_15980);
nor U16994 (N_16994,N_15674,N_16714);
xor U16995 (N_16995,N_15605,N_16777);
and U16996 (N_16996,N_16530,N_16013);
xnor U16997 (N_16997,N_15764,N_16315);
xor U16998 (N_16998,N_15971,N_15854);
and U16999 (N_16999,N_15984,N_16223);
or U17000 (N_17000,N_16172,N_15832);
or U17001 (N_17001,N_15652,N_16558);
nor U17002 (N_17002,N_16553,N_15660);
nand U17003 (N_17003,N_16216,N_15850);
and U17004 (N_17004,N_16758,N_16717);
or U17005 (N_17005,N_16244,N_15770);
or U17006 (N_17006,N_16126,N_16351);
nor U17007 (N_17007,N_15853,N_15817);
nand U17008 (N_17008,N_15700,N_16798);
nor U17009 (N_17009,N_16036,N_15688);
and U17010 (N_17010,N_16455,N_15720);
nor U17011 (N_17011,N_15767,N_16040);
nor U17012 (N_17012,N_16176,N_15847);
nor U17013 (N_17013,N_15643,N_15675);
nor U17014 (N_17014,N_16242,N_16636);
nand U17015 (N_17015,N_16010,N_16574);
nand U17016 (N_17016,N_15741,N_16504);
nand U17017 (N_17017,N_16218,N_16482);
and U17018 (N_17018,N_15711,N_16437);
nand U17019 (N_17019,N_15818,N_15836);
nand U17020 (N_17020,N_16164,N_16113);
and U17021 (N_17021,N_16177,N_16641);
xnor U17022 (N_17022,N_16052,N_16376);
or U17023 (N_17023,N_16140,N_15793);
xnor U17024 (N_17024,N_16096,N_16488);
nor U17025 (N_17025,N_16592,N_16313);
xor U17026 (N_17026,N_15673,N_15783);
nand U17027 (N_17027,N_16692,N_15978);
and U17028 (N_17028,N_16141,N_16114);
or U17029 (N_17029,N_15958,N_16214);
nor U17030 (N_17030,N_16290,N_16754);
or U17031 (N_17031,N_16693,N_16100);
and U17032 (N_17032,N_16106,N_15968);
nand U17033 (N_17033,N_16654,N_16400);
nor U17034 (N_17034,N_15801,N_16682);
nor U17035 (N_17035,N_16573,N_16303);
or U17036 (N_17036,N_16690,N_15822);
nand U17037 (N_17037,N_15713,N_16123);
nand U17038 (N_17038,N_16774,N_16625);
nor U17039 (N_17039,N_16710,N_15977);
and U17040 (N_17040,N_15771,N_16738);
nand U17041 (N_17041,N_16563,N_16353);
or U17042 (N_17042,N_15661,N_16370);
or U17043 (N_17043,N_16221,N_15931);
or U17044 (N_17044,N_16382,N_15899);
nand U17045 (N_17045,N_15910,N_16088);
xnor U17046 (N_17046,N_15655,N_15881);
and U17047 (N_17047,N_16496,N_16753);
xor U17048 (N_17048,N_15780,N_15782);
nand U17049 (N_17049,N_15624,N_16548);
nand U17050 (N_17050,N_16638,N_16656);
xnor U17051 (N_17051,N_16023,N_16414);
nand U17052 (N_17052,N_16035,N_15911);
and U17053 (N_17053,N_16270,N_16055);
nor U17054 (N_17054,N_15921,N_16121);
xor U17055 (N_17055,N_16555,N_16703);
nand U17056 (N_17056,N_15799,N_15639);
nor U17057 (N_17057,N_16509,N_16143);
or U17058 (N_17058,N_15902,N_15974);
xnor U17059 (N_17059,N_15922,N_15939);
xor U17060 (N_17060,N_15619,N_16230);
nand U17061 (N_17061,N_15662,N_16529);
and U17062 (N_17062,N_15710,N_16047);
nand U17063 (N_17063,N_16719,N_16186);
xor U17064 (N_17064,N_16580,N_15694);
xor U17065 (N_17065,N_16181,N_16355);
or U17066 (N_17066,N_16022,N_16346);
xnor U17067 (N_17067,N_15898,N_16428);
nor U17068 (N_17068,N_16628,N_16776);
and U17069 (N_17069,N_16103,N_16027);
and U17070 (N_17070,N_16029,N_16763);
or U17071 (N_17071,N_16528,N_16533);
nand U17072 (N_17072,N_15646,N_15929);
nor U17073 (N_17073,N_16755,N_16462);
nor U17074 (N_17074,N_16142,N_16286);
xnor U17075 (N_17075,N_16489,N_15721);
nor U17076 (N_17076,N_15951,N_16388);
nor U17077 (N_17077,N_15890,N_16359);
and U17078 (N_17078,N_16064,N_16546);
xor U17079 (N_17079,N_16262,N_15626);
nand U17080 (N_17080,N_16374,N_15679);
and U17081 (N_17081,N_15867,N_16607);
or U17082 (N_17082,N_15669,N_16390);
and U17083 (N_17083,N_15800,N_15612);
xor U17084 (N_17084,N_16119,N_16552);
and U17085 (N_17085,N_16740,N_16691);
or U17086 (N_17086,N_16234,N_16341);
nor U17087 (N_17087,N_15677,N_15803);
and U17088 (N_17088,N_16507,N_16569);
nor U17089 (N_17089,N_16254,N_16407);
or U17090 (N_17090,N_16646,N_16697);
nand U17091 (N_17091,N_16612,N_16247);
and U17092 (N_17092,N_15797,N_16648);
or U17093 (N_17093,N_16129,N_16688);
nor U17094 (N_17094,N_15610,N_16796);
and U17095 (N_17095,N_16412,N_16175);
xnor U17096 (N_17096,N_15642,N_15653);
or U17097 (N_17097,N_16770,N_16163);
or U17098 (N_17098,N_16179,N_16789);
or U17099 (N_17099,N_16215,N_16248);
nand U17100 (N_17100,N_15820,N_15682);
nand U17101 (N_17101,N_15909,N_16002);
or U17102 (N_17102,N_15760,N_16208);
nor U17103 (N_17103,N_16091,N_15810);
xor U17104 (N_17104,N_16589,N_16122);
nand U17105 (N_17105,N_16016,N_15952);
nand U17106 (N_17106,N_16124,N_16475);
or U17107 (N_17107,N_15897,N_16671);
or U17108 (N_17108,N_16752,N_15607);
nor U17109 (N_17109,N_16168,N_15863);
xor U17110 (N_17110,N_15727,N_16594);
or U17111 (N_17111,N_15839,N_16264);
xnor U17112 (N_17112,N_16053,N_16586);
nor U17113 (N_17113,N_15776,N_16167);
and U17114 (N_17114,N_15731,N_15875);
or U17115 (N_17115,N_16117,N_16424);
xnor U17116 (N_17116,N_16771,N_16136);
nand U17117 (N_17117,N_15647,N_16024);
nand U17118 (N_17118,N_16165,N_16500);
xor U17119 (N_17119,N_16044,N_16735);
nor U17120 (N_17120,N_16517,N_16492);
nand U17121 (N_17121,N_15891,N_16335);
nand U17122 (N_17122,N_16338,N_16133);
or U17123 (N_17123,N_16783,N_16156);
and U17124 (N_17124,N_16161,N_16725);
or U17125 (N_17125,N_15945,N_16067);
or U17126 (N_17126,N_16670,N_15719);
nand U17127 (N_17127,N_16146,N_16518);
and U17128 (N_17128,N_16307,N_16527);
nor U17129 (N_17129,N_15999,N_16268);
or U17130 (N_17130,N_16095,N_16729);
nor U17131 (N_17131,N_16742,N_16452);
nand U17132 (N_17132,N_15926,N_16319);
nand U17133 (N_17133,N_15798,N_16060);
xor U17134 (N_17134,N_16194,N_16635);
xor U17135 (N_17135,N_15924,N_16200);
and U17136 (N_17136,N_15730,N_16795);
and U17137 (N_17137,N_16760,N_16698);
nand U17138 (N_17138,N_16578,N_16544);
nand U17139 (N_17139,N_16273,N_16520);
xor U17140 (N_17140,N_15781,N_15777);
xnor U17141 (N_17141,N_16267,N_16609);
xor U17142 (N_17142,N_16571,N_16700);
nor U17143 (N_17143,N_15962,N_15668);
nor U17144 (N_17144,N_16160,N_16534);
and U17145 (N_17145,N_15878,N_16711);
xor U17146 (N_17146,N_16061,N_16237);
and U17147 (N_17147,N_16368,N_16726);
nand U17148 (N_17148,N_16318,N_16616);
xor U17149 (N_17149,N_16068,N_16728);
nand U17150 (N_17150,N_16545,N_16339);
nand U17151 (N_17151,N_16316,N_16386);
xnor U17152 (N_17152,N_16627,N_16321);
nand U17153 (N_17153,N_16778,N_15895);
and U17154 (N_17154,N_15670,N_16094);
and U17155 (N_17155,N_16797,N_15636);
or U17156 (N_17156,N_15715,N_16380);
and U17157 (N_17157,N_15631,N_16330);
and U17158 (N_17158,N_15866,N_16288);
nand U17159 (N_17159,N_16680,N_15690);
xor U17160 (N_17160,N_16415,N_16756);
xnor U17161 (N_17161,N_16707,N_15630);
nand U17162 (N_17162,N_15732,N_15737);
nor U17163 (N_17163,N_16672,N_15759);
or U17164 (N_17164,N_16759,N_15654);
nand U17165 (N_17165,N_15848,N_16066);
nor U17166 (N_17166,N_15824,N_16716);
or U17167 (N_17167,N_16418,N_15620);
nor U17168 (N_17168,N_16111,N_15663);
and U17169 (N_17169,N_16345,N_15857);
nor U17170 (N_17170,N_15937,N_16522);
nand U17171 (N_17171,N_15766,N_16652);
or U17172 (N_17172,N_16399,N_16630);
xnor U17173 (N_17173,N_16525,N_16642);
and U17174 (N_17174,N_15873,N_16493);
or U17175 (N_17175,N_15855,N_16512);
nand U17176 (N_17176,N_16433,N_16590);
or U17177 (N_17177,N_15632,N_16450);
and U17178 (N_17178,N_16587,N_16169);
xor U17179 (N_17179,N_15870,N_16478);
nor U17180 (N_17180,N_16679,N_16008);
and U17181 (N_17181,N_15970,N_16779);
nor U17182 (N_17182,N_16781,N_16790);
or U17183 (N_17183,N_16508,N_16668);
nand U17184 (N_17184,N_16235,N_15954);
or U17185 (N_17185,N_15851,N_15960);
nand U17186 (N_17186,N_16371,N_15746);
nand U17187 (N_17187,N_16132,N_15882);
nor U17188 (N_17188,N_16238,N_16147);
or U17189 (N_17189,N_16219,N_16205);
xnor U17190 (N_17190,N_15621,N_16190);
nand U17191 (N_17191,N_16302,N_16547);
and U17192 (N_17192,N_16503,N_15877);
nand U17193 (N_17193,N_16511,N_15627);
nand U17194 (N_17194,N_15600,N_16602);
nor U17195 (N_17195,N_16093,N_15865);
or U17196 (N_17196,N_16232,N_16249);
nor U17197 (N_17197,N_15762,N_16551);
and U17198 (N_17198,N_16632,N_16360);
nand U17199 (N_17199,N_16187,N_15858);
xor U17200 (N_17200,N_15938,N_16083);
nor U17201 (N_17201,N_16084,N_16069);
and U17202 (N_17202,N_16733,N_15640);
or U17203 (N_17203,N_16712,N_15606);
nor U17204 (N_17204,N_15957,N_15894);
or U17205 (N_17205,N_15743,N_16523);
or U17206 (N_17206,N_15973,N_16231);
nand U17207 (N_17207,N_16669,N_15740);
nor U17208 (N_17208,N_16152,N_16657);
or U17209 (N_17209,N_16171,N_16608);
nor U17210 (N_17210,N_16166,N_16516);
nand U17211 (N_17211,N_16090,N_16401);
and U17212 (N_17212,N_16715,N_15775);
xnor U17213 (N_17213,N_15963,N_16356);
or U17214 (N_17214,N_16236,N_15691);
or U17215 (N_17215,N_16101,N_16696);
nand U17216 (N_17216,N_15965,N_15876);
or U17217 (N_17217,N_16521,N_16039);
or U17218 (N_17218,N_16336,N_16324);
and U17219 (N_17219,N_15834,N_16025);
xor U17220 (N_17220,N_16184,N_16465);
or U17221 (N_17221,N_15976,N_16799);
or U17222 (N_17222,N_15659,N_15754);
nand U17223 (N_17223,N_15687,N_16435);
or U17224 (N_17224,N_16201,N_16673);
xnor U17225 (N_17225,N_16191,N_15791);
nor U17226 (N_17226,N_16282,N_15701);
or U17227 (N_17227,N_16567,N_16151);
and U17228 (N_17228,N_16535,N_16411);
and U17229 (N_17229,N_15880,N_16031);
xor U17230 (N_17230,N_16599,N_16463);
nand U17231 (N_17231,N_15979,N_16265);
nor U17232 (N_17232,N_16637,N_15733);
or U17233 (N_17233,N_16082,N_16731);
nor U17234 (N_17234,N_16220,N_15618);
xor U17235 (N_17235,N_15811,N_16004);
nor U17236 (N_17236,N_15886,N_16597);
or U17237 (N_17237,N_15686,N_15725);
nand U17238 (N_17238,N_15900,N_16352);
xnor U17239 (N_17239,N_16110,N_16695);
and U17240 (N_17240,N_15786,N_15765);
nand U17241 (N_17241,N_15671,N_15695);
xor U17242 (N_17242,N_15828,N_16020);
nor U17243 (N_17243,N_16314,N_16426);
and U17244 (N_17244,N_15906,N_16786);
or U17245 (N_17245,N_16054,N_16784);
or U17246 (N_17246,N_16404,N_15805);
nand U17247 (N_17247,N_16598,N_16560);
xnor U17248 (N_17248,N_16037,N_16474);
nor U17249 (N_17249,N_16310,N_16071);
and U17250 (N_17250,N_16012,N_16210);
nor U17251 (N_17251,N_15681,N_15943);
nor U17252 (N_17252,N_15985,N_15744);
nand U17253 (N_17253,N_15602,N_15815);
and U17254 (N_17254,N_16322,N_16451);
or U17255 (N_17255,N_16764,N_16312);
or U17256 (N_17256,N_16631,N_15745);
and U17257 (N_17257,N_16263,N_16748);
nor U17258 (N_17258,N_16393,N_16429);
nand U17259 (N_17259,N_15821,N_15672);
nor U17260 (N_17260,N_15613,N_16791);
nor U17261 (N_17261,N_16709,N_16285);
nand U17262 (N_17262,N_15794,N_16678);
xnor U17263 (N_17263,N_16378,N_15809);
or U17264 (N_17264,N_16109,N_16699);
and U17265 (N_17265,N_16076,N_16739);
nor U17266 (N_17266,N_16519,N_15996);
and U17267 (N_17267,N_16157,N_16751);
and U17268 (N_17268,N_16118,N_16251);
nor U17269 (N_17269,N_15846,N_16665);
or U17270 (N_17270,N_15616,N_16327);
nand U17271 (N_17271,N_15644,N_15903);
or U17272 (N_17272,N_16459,N_16720);
and U17273 (N_17273,N_15634,N_16708);
and U17274 (N_17274,N_16442,N_15693);
nor U17275 (N_17275,N_16466,N_16193);
nor U17276 (N_17276,N_16655,N_16582);
and U17277 (N_17277,N_16357,N_16241);
and U17278 (N_17278,N_16730,N_16495);
and U17279 (N_17279,N_15702,N_16585);
and U17280 (N_17280,N_16050,N_15812);
xnor U17281 (N_17281,N_16457,N_16542);
nand U17282 (N_17282,N_15806,N_16099);
xnor U17283 (N_17283,N_16502,N_15997);
nor U17284 (N_17284,N_16662,N_15650);
nand U17285 (N_17285,N_15758,N_16350);
and U17286 (N_17286,N_16222,N_16596);
and U17287 (N_17287,N_15869,N_16615);
xnor U17288 (N_17288,N_16593,N_15729);
nand U17289 (N_17289,N_16233,N_16444);
nand U17290 (N_17290,N_16689,N_16074);
xor U17291 (N_17291,N_15712,N_16306);
or U17292 (N_17292,N_16366,N_16600);
nand U17293 (N_17293,N_16150,N_15789);
xnor U17294 (N_17294,N_16391,N_16498);
nor U17295 (N_17295,N_16041,N_16613);
or U17296 (N_17296,N_15975,N_16595);
or U17297 (N_17297,N_16337,N_16622);
or U17298 (N_17298,N_15748,N_15972);
nand U17299 (N_17299,N_15990,N_16794);
nor U17300 (N_17300,N_16051,N_16620);
xor U17301 (N_17301,N_15927,N_15665);
nand U17302 (N_17302,N_16448,N_15773);
nand U17303 (N_17303,N_16364,N_16019);
or U17304 (N_17304,N_16566,N_16275);
or U17305 (N_17305,N_16294,N_15862);
nand U17306 (N_17306,N_16342,N_16131);
and U17307 (N_17307,N_15989,N_15796);
nand U17308 (N_17308,N_16398,N_15879);
nand U17309 (N_17309,N_16162,N_16514);
and U17310 (N_17310,N_16676,N_15941);
or U17311 (N_17311,N_16394,N_16467);
or U17312 (N_17312,N_15751,N_16204);
or U17313 (N_17313,N_15908,N_15747);
and U17314 (N_17314,N_15666,N_16780);
xnor U17315 (N_17315,N_16228,N_15802);
nand U17316 (N_17316,N_16447,N_15697);
xor U17317 (N_17317,N_16202,N_15649);
xnor U17318 (N_17318,N_16541,N_16732);
nor U17319 (N_17319,N_16329,N_16105);
nor U17320 (N_17320,N_16075,N_15956);
xor U17321 (N_17321,N_16295,N_16396);
nand U17322 (N_17322,N_15648,N_16159);
and U17323 (N_17323,N_16604,N_16736);
nor U17324 (N_17324,N_16256,N_15629);
nand U17325 (N_17325,N_16326,N_16154);
or U17326 (N_17326,N_16108,N_16291);
nand U17327 (N_17327,N_16258,N_15837);
nor U17328 (N_17328,N_15844,N_16650);
nor U17329 (N_17329,N_15959,N_15913);
nand U17330 (N_17330,N_16487,N_16362);
or U17331 (N_17331,N_15826,N_15753);
nor U17332 (N_17332,N_15678,N_16009);
xnor U17333 (N_17333,N_15750,N_16757);
and U17334 (N_17334,N_16621,N_16643);
nor U17335 (N_17335,N_15995,N_16664);
xnor U17336 (N_17336,N_16658,N_16211);
nor U17337 (N_17337,N_15645,N_16425);
and U17338 (N_17338,N_15755,N_16575);
and U17339 (N_17339,N_16416,N_16772);
or U17340 (N_17340,N_16198,N_16058);
and U17341 (N_17341,N_16744,N_15769);
or U17342 (N_17342,N_16293,N_16483);
or U17343 (N_17343,N_16570,N_16213);
nor U17344 (N_17344,N_15987,N_15833);
xnor U17345 (N_17345,N_15823,N_16645);
nor U17346 (N_17346,N_15772,N_16494);
xor U17347 (N_17347,N_16092,N_15868);
and U17348 (N_17348,N_15872,N_15964);
xor U17349 (N_17349,N_16305,N_16384);
or U17350 (N_17350,N_15736,N_16043);
or U17351 (N_17351,N_16705,N_16287);
nor U17352 (N_17352,N_15752,N_16259);
or U17353 (N_17353,N_16134,N_16410);
and U17354 (N_17354,N_16260,N_16192);
xor U17355 (N_17355,N_16348,N_16045);
nor U17356 (N_17356,N_16687,N_16240);
xnor U17357 (N_17357,N_15742,N_16057);
and U17358 (N_17358,N_16389,N_16734);
and U17359 (N_17359,N_16203,N_15923);
or U17360 (N_17360,N_16197,N_16340);
and U17361 (N_17361,N_16749,N_15885);
or U17362 (N_17362,N_15842,N_15637);
and U17363 (N_17363,N_16443,N_15845);
nor U17364 (N_17364,N_16387,N_16320);
xnor U17365 (N_17365,N_15638,N_16385);
xor U17366 (N_17366,N_16684,N_15757);
xor U17367 (N_17367,N_15831,N_16299);
xor U17368 (N_17368,N_16034,N_15628);
nand U17369 (N_17369,N_16046,N_16367);
nor U17370 (N_17370,N_16274,N_16653);
or U17371 (N_17371,N_15825,N_16536);
nand U17372 (N_17372,N_15704,N_16392);
or U17373 (N_17373,N_15698,N_16788);
nor U17374 (N_17374,N_16765,N_16403);
xnor U17375 (N_17375,N_16280,N_16434);
or U17376 (N_17376,N_15718,N_16006);
nor U17377 (N_17377,N_16148,N_15641);
or U17378 (N_17378,N_16538,N_16116);
nor U17379 (N_17379,N_16743,N_16304);
and U17380 (N_17380,N_15884,N_16227);
or U17381 (N_17381,N_16283,N_16018);
or U17382 (N_17382,N_16349,N_16347);
or U17383 (N_17383,N_15928,N_16011);
or U17384 (N_17384,N_16531,N_15623);
or U17385 (N_17385,N_16550,N_16427);
xnor U17386 (N_17386,N_15726,N_16395);
nor U17387 (N_17387,N_16332,N_15998);
nand U17388 (N_17388,N_15982,N_16572);
nor U17389 (N_17389,N_15916,N_16723);
xor U17390 (N_17390,N_16775,N_16785);
nor U17391 (N_17391,N_16065,N_16007);
or U17392 (N_17392,N_16383,N_16015);
nor U17393 (N_17393,N_16624,N_15689);
or U17394 (N_17394,N_16479,N_15716);
or U17395 (N_17395,N_15676,N_16473);
nor U17396 (N_17396,N_16308,N_16761);
and U17397 (N_17397,N_15705,N_16062);
nor U17398 (N_17398,N_16666,N_15723);
or U17399 (N_17399,N_16077,N_15852);
nor U17400 (N_17400,N_15627,N_15981);
xor U17401 (N_17401,N_16005,N_16368);
nand U17402 (N_17402,N_16390,N_15861);
and U17403 (N_17403,N_16323,N_15838);
or U17404 (N_17404,N_15748,N_16160);
nand U17405 (N_17405,N_15776,N_16587);
nand U17406 (N_17406,N_15860,N_16171);
xor U17407 (N_17407,N_15672,N_16095);
nor U17408 (N_17408,N_15626,N_15619);
xnor U17409 (N_17409,N_16461,N_15786);
nor U17410 (N_17410,N_16129,N_16717);
nor U17411 (N_17411,N_16269,N_15979);
nand U17412 (N_17412,N_15873,N_16506);
xor U17413 (N_17413,N_16090,N_16322);
xor U17414 (N_17414,N_16057,N_16657);
or U17415 (N_17415,N_16406,N_16444);
nor U17416 (N_17416,N_16161,N_16497);
and U17417 (N_17417,N_16672,N_16292);
xor U17418 (N_17418,N_15926,N_16252);
nand U17419 (N_17419,N_16641,N_16425);
xnor U17420 (N_17420,N_15846,N_16056);
xor U17421 (N_17421,N_16702,N_16116);
nor U17422 (N_17422,N_16100,N_16666);
nand U17423 (N_17423,N_16386,N_16655);
nand U17424 (N_17424,N_16095,N_16464);
or U17425 (N_17425,N_16050,N_15732);
nand U17426 (N_17426,N_16440,N_16450);
nor U17427 (N_17427,N_16370,N_15754);
and U17428 (N_17428,N_15702,N_16592);
or U17429 (N_17429,N_16168,N_16322);
and U17430 (N_17430,N_15856,N_16500);
xnor U17431 (N_17431,N_15627,N_15831);
and U17432 (N_17432,N_16755,N_16098);
nor U17433 (N_17433,N_16253,N_16744);
xnor U17434 (N_17434,N_16336,N_15825);
nor U17435 (N_17435,N_16283,N_15697);
xnor U17436 (N_17436,N_15924,N_16309);
nand U17437 (N_17437,N_16274,N_15837);
or U17438 (N_17438,N_16540,N_16640);
nand U17439 (N_17439,N_16694,N_16257);
and U17440 (N_17440,N_15799,N_15850);
and U17441 (N_17441,N_16713,N_16185);
nand U17442 (N_17442,N_15917,N_16317);
and U17443 (N_17443,N_16519,N_16224);
and U17444 (N_17444,N_16620,N_16518);
nor U17445 (N_17445,N_16785,N_16132);
and U17446 (N_17446,N_16489,N_16190);
or U17447 (N_17447,N_16213,N_16656);
and U17448 (N_17448,N_16074,N_16302);
nand U17449 (N_17449,N_16392,N_16010);
nor U17450 (N_17450,N_16065,N_16346);
xor U17451 (N_17451,N_16693,N_16189);
nand U17452 (N_17452,N_16787,N_15823);
or U17453 (N_17453,N_15687,N_16065);
xor U17454 (N_17454,N_16201,N_16769);
or U17455 (N_17455,N_16253,N_15713);
or U17456 (N_17456,N_16049,N_16538);
or U17457 (N_17457,N_16083,N_16679);
xnor U17458 (N_17458,N_16469,N_16348);
nor U17459 (N_17459,N_16389,N_16260);
and U17460 (N_17460,N_16348,N_15726);
or U17461 (N_17461,N_15932,N_16644);
or U17462 (N_17462,N_15889,N_16164);
nand U17463 (N_17463,N_16519,N_16210);
or U17464 (N_17464,N_16510,N_15867);
or U17465 (N_17465,N_16041,N_15931);
nand U17466 (N_17466,N_15829,N_16474);
and U17467 (N_17467,N_16158,N_15840);
or U17468 (N_17468,N_16710,N_16731);
or U17469 (N_17469,N_16415,N_15769);
nor U17470 (N_17470,N_16468,N_16408);
and U17471 (N_17471,N_16757,N_16303);
or U17472 (N_17472,N_15913,N_16302);
and U17473 (N_17473,N_16240,N_15920);
nand U17474 (N_17474,N_16384,N_16349);
or U17475 (N_17475,N_16753,N_15838);
or U17476 (N_17476,N_15776,N_16007);
and U17477 (N_17477,N_16260,N_16583);
or U17478 (N_17478,N_16353,N_15666);
xor U17479 (N_17479,N_15994,N_16455);
nand U17480 (N_17480,N_16378,N_16744);
nand U17481 (N_17481,N_16448,N_16705);
nor U17482 (N_17482,N_16245,N_16703);
nor U17483 (N_17483,N_15734,N_16044);
and U17484 (N_17484,N_15814,N_16081);
xnor U17485 (N_17485,N_16665,N_15640);
nand U17486 (N_17486,N_16734,N_15895);
or U17487 (N_17487,N_15901,N_16795);
nor U17488 (N_17488,N_16117,N_16637);
or U17489 (N_17489,N_15742,N_16343);
and U17490 (N_17490,N_16215,N_16323);
nor U17491 (N_17491,N_16634,N_15845);
xnor U17492 (N_17492,N_16722,N_16341);
and U17493 (N_17493,N_16186,N_16053);
or U17494 (N_17494,N_16025,N_15927);
or U17495 (N_17495,N_16672,N_16474);
and U17496 (N_17496,N_15723,N_16769);
nor U17497 (N_17497,N_16678,N_15612);
and U17498 (N_17498,N_16685,N_16533);
nand U17499 (N_17499,N_15773,N_16150);
nand U17500 (N_17500,N_15648,N_15980);
nand U17501 (N_17501,N_16578,N_16668);
or U17502 (N_17502,N_16378,N_16629);
or U17503 (N_17503,N_16458,N_16016);
or U17504 (N_17504,N_16312,N_16089);
and U17505 (N_17505,N_15672,N_16414);
nand U17506 (N_17506,N_16623,N_16442);
and U17507 (N_17507,N_16578,N_16120);
and U17508 (N_17508,N_16355,N_15647);
and U17509 (N_17509,N_15627,N_15641);
and U17510 (N_17510,N_15905,N_16755);
or U17511 (N_17511,N_16072,N_16744);
nand U17512 (N_17512,N_15618,N_15941);
nand U17513 (N_17513,N_16391,N_16264);
xor U17514 (N_17514,N_16744,N_15920);
or U17515 (N_17515,N_16609,N_16123);
xor U17516 (N_17516,N_16673,N_16444);
xnor U17517 (N_17517,N_16053,N_16593);
xor U17518 (N_17518,N_15765,N_15912);
nand U17519 (N_17519,N_16184,N_16634);
nor U17520 (N_17520,N_16045,N_15764);
and U17521 (N_17521,N_15859,N_16563);
and U17522 (N_17522,N_16091,N_16711);
nor U17523 (N_17523,N_16780,N_16411);
and U17524 (N_17524,N_15765,N_16536);
nor U17525 (N_17525,N_16289,N_16459);
xor U17526 (N_17526,N_15912,N_16775);
and U17527 (N_17527,N_16422,N_16072);
nor U17528 (N_17528,N_16642,N_15879);
and U17529 (N_17529,N_16276,N_16481);
and U17530 (N_17530,N_16177,N_16381);
and U17531 (N_17531,N_16689,N_16208);
nand U17532 (N_17532,N_16727,N_15999);
nand U17533 (N_17533,N_16643,N_16045);
nand U17534 (N_17534,N_16603,N_16400);
and U17535 (N_17535,N_16781,N_16476);
xnor U17536 (N_17536,N_15998,N_16407);
nand U17537 (N_17537,N_16191,N_16640);
xor U17538 (N_17538,N_15917,N_16565);
nand U17539 (N_17539,N_16789,N_16112);
nor U17540 (N_17540,N_16031,N_16049);
and U17541 (N_17541,N_16748,N_16593);
or U17542 (N_17542,N_16097,N_16290);
or U17543 (N_17543,N_16335,N_16655);
xor U17544 (N_17544,N_16279,N_16347);
nand U17545 (N_17545,N_16178,N_16385);
xor U17546 (N_17546,N_15841,N_16735);
nor U17547 (N_17547,N_16111,N_16458);
nor U17548 (N_17548,N_16326,N_16065);
nor U17549 (N_17549,N_15660,N_16515);
and U17550 (N_17550,N_16175,N_16178);
or U17551 (N_17551,N_15802,N_16787);
and U17552 (N_17552,N_15693,N_16160);
and U17553 (N_17553,N_16154,N_15931);
or U17554 (N_17554,N_15991,N_15746);
or U17555 (N_17555,N_15932,N_15873);
nor U17556 (N_17556,N_15902,N_16757);
nor U17557 (N_17557,N_15969,N_15985);
nor U17558 (N_17558,N_16434,N_16697);
and U17559 (N_17559,N_15849,N_16266);
and U17560 (N_17560,N_15861,N_16541);
nor U17561 (N_17561,N_15704,N_15613);
or U17562 (N_17562,N_16493,N_16441);
or U17563 (N_17563,N_15747,N_16398);
nor U17564 (N_17564,N_16211,N_15896);
or U17565 (N_17565,N_15835,N_16129);
nand U17566 (N_17566,N_15714,N_16486);
nor U17567 (N_17567,N_16401,N_15951);
or U17568 (N_17568,N_16346,N_16550);
or U17569 (N_17569,N_15947,N_16019);
nand U17570 (N_17570,N_16392,N_15869);
xor U17571 (N_17571,N_15996,N_16015);
xnor U17572 (N_17572,N_16272,N_15620);
and U17573 (N_17573,N_15629,N_16595);
nand U17574 (N_17574,N_16254,N_16621);
nand U17575 (N_17575,N_16763,N_16709);
xor U17576 (N_17576,N_16100,N_15929);
nor U17577 (N_17577,N_16337,N_15908);
nand U17578 (N_17578,N_16432,N_16131);
nor U17579 (N_17579,N_16726,N_16543);
or U17580 (N_17580,N_16556,N_16201);
and U17581 (N_17581,N_15944,N_16168);
and U17582 (N_17582,N_16689,N_16583);
and U17583 (N_17583,N_16325,N_15754);
and U17584 (N_17584,N_16214,N_16191);
nor U17585 (N_17585,N_16153,N_16787);
nand U17586 (N_17586,N_16439,N_16210);
or U17587 (N_17587,N_16148,N_15642);
and U17588 (N_17588,N_15625,N_16053);
nand U17589 (N_17589,N_16076,N_16165);
xor U17590 (N_17590,N_16036,N_16570);
nand U17591 (N_17591,N_15906,N_16092);
and U17592 (N_17592,N_15722,N_16353);
nand U17593 (N_17593,N_15928,N_16291);
and U17594 (N_17594,N_16064,N_16396);
nor U17595 (N_17595,N_15608,N_16394);
and U17596 (N_17596,N_15897,N_16430);
nand U17597 (N_17597,N_15845,N_15826);
nand U17598 (N_17598,N_16492,N_16426);
nand U17599 (N_17599,N_15835,N_16398);
nand U17600 (N_17600,N_16333,N_16080);
nor U17601 (N_17601,N_16737,N_16289);
nor U17602 (N_17602,N_15757,N_16314);
xnor U17603 (N_17603,N_16373,N_16220);
or U17604 (N_17604,N_16558,N_16380);
nand U17605 (N_17605,N_15776,N_15915);
nor U17606 (N_17606,N_15681,N_15768);
nor U17607 (N_17607,N_15801,N_16151);
and U17608 (N_17608,N_16590,N_15904);
xnor U17609 (N_17609,N_16613,N_16259);
nand U17610 (N_17610,N_15635,N_16079);
and U17611 (N_17611,N_16295,N_16040);
and U17612 (N_17612,N_16129,N_16661);
nor U17613 (N_17613,N_15610,N_15998);
or U17614 (N_17614,N_15972,N_16760);
or U17615 (N_17615,N_15602,N_15681);
xnor U17616 (N_17616,N_16726,N_15768);
xnor U17617 (N_17617,N_16650,N_16627);
or U17618 (N_17618,N_15925,N_16400);
nand U17619 (N_17619,N_16538,N_15961);
nand U17620 (N_17620,N_15914,N_16570);
and U17621 (N_17621,N_16065,N_16410);
or U17622 (N_17622,N_16423,N_16782);
nand U17623 (N_17623,N_16100,N_16670);
or U17624 (N_17624,N_16331,N_16614);
and U17625 (N_17625,N_16112,N_15632);
or U17626 (N_17626,N_16278,N_15636);
nand U17627 (N_17627,N_16771,N_15749);
and U17628 (N_17628,N_16063,N_16074);
xnor U17629 (N_17629,N_15867,N_15836);
xor U17630 (N_17630,N_16115,N_16782);
or U17631 (N_17631,N_15849,N_16184);
xor U17632 (N_17632,N_15907,N_16592);
or U17633 (N_17633,N_16527,N_16101);
nor U17634 (N_17634,N_16596,N_16685);
nand U17635 (N_17635,N_15725,N_15774);
or U17636 (N_17636,N_16419,N_15662);
or U17637 (N_17637,N_16301,N_16172);
and U17638 (N_17638,N_15711,N_16516);
nand U17639 (N_17639,N_16475,N_16467);
nand U17640 (N_17640,N_16200,N_16487);
nand U17641 (N_17641,N_16080,N_16607);
or U17642 (N_17642,N_15990,N_16348);
and U17643 (N_17643,N_15930,N_16355);
and U17644 (N_17644,N_15654,N_15793);
xor U17645 (N_17645,N_15609,N_16551);
xnor U17646 (N_17646,N_15913,N_16065);
or U17647 (N_17647,N_16250,N_15806);
or U17648 (N_17648,N_16154,N_16764);
nand U17649 (N_17649,N_16017,N_16570);
nand U17650 (N_17650,N_16286,N_16484);
nand U17651 (N_17651,N_16786,N_16197);
nand U17652 (N_17652,N_16700,N_16437);
or U17653 (N_17653,N_16427,N_16224);
and U17654 (N_17654,N_16101,N_16492);
or U17655 (N_17655,N_16379,N_15600);
nand U17656 (N_17656,N_16731,N_15690);
and U17657 (N_17657,N_16199,N_16340);
and U17658 (N_17658,N_16200,N_16135);
or U17659 (N_17659,N_16529,N_16675);
and U17660 (N_17660,N_15807,N_16266);
and U17661 (N_17661,N_15930,N_16656);
nand U17662 (N_17662,N_16190,N_16614);
and U17663 (N_17663,N_16690,N_15999);
or U17664 (N_17664,N_16157,N_16546);
or U17665 (N_17665,N_16354,N_15877);
xnor U17666 (N_17666,N_15929,N_16309);
and U17667 (N_17667,N_16396,N_16403);
or U17668 (N_17668,N_16714,N_16176);
xnor U17669 (N_17669,N_16072,N_15712);
or U17670 (N_17670,N_15983,N_16625);
xnor U17671 (N_17671,N_16579,N_16441);
nand U17672 (N_17672,N_15608,N_16417);
or U17673 (N_17673,N_16782,N_16066);
xnor U17674 (N_17674,N_15919,N_15652);
nor U17675 (N_17675,N_16612,N_16765);
and U17676 (N_17676,N_16502,N_16244);
nor U17677 (N_17677,N_15924,N_15812);
nand U17678 (N_17678,N_16550,N_15872);
nor U17679 (N_17679,N_16535,N_15603);
nor U17680 (N_17680,N_15973,N_16343);
xnor U17681 (N_17681,N_16541,N_15673);
nand U17682 (N_17682,N_16010,N_16609);
or U17683 (N_17683,N_16293,N_16352);
and U17684 (N_17684,N_15854,N_15728);
or U17685 (N_17685,N_15636,N_16175);
and U17686 (N_17686,N_16113,N_16363);
nor U17687 (N_17687,N_16385,N_16136);
xor U17688 (N_17688,N_15949,N_15763);
and U17689 (N_17689,N_16144,N_15696);
and U17690 (N_17690,N_15711,N_16512);
or U17691 (N_17691,N_16210,N_15951);
nand U17692 (N_17692,N_15832,N_16757);
xor U17693 (N_17693,N_16695,N_15717);
nand U17694 (N_17694,N_16650,N_16285);
nand U17695 (N_17695,N_15676,N_16001);
nand U17696 (N_17696,N_15635,N_16765);
xnor U17697 (N_17697,N_16021,N_16698);
xnor U17698 (N_17698,N_16015,N_15829);
nor U17699 (N_17699,N_15925,N_15726);
xor U17700 (N_17700,N_16456,N_16470);
nor U17701 (N_17701,N_16264,N_16586);
and U17702 (N_17702,N_15873,N_16368);
nand U17703 (N_17703,N_16784,N_15686);
xor U17704 (N_17704,N_16394,N_16148);
xor U17705 (N_17705,N_16619,N_16588);
and U17706 (N_17706,N_16721,N_16788);
and U17707 (N_17707,N_16524,N_15745);
or U17708 (N_17708,N_15727,N_15814);
nor U17709 (N_17709,N_16016,N_15913);
and U17710 (N_17710,N_16564,N_16379);
xor U17711 (N_17711,N_16579,N_16453);
nor U17712 (N_17712,N_16379,N_16586);
nor U17713 (N_17713,N_15832,N_15636);
or U17714 (N_17714,N_16495,N_15676);
or U17715 (N_17715,N_15653,N_16650);
or U17716 (N_17716,N_16322,N_16088);
nor U17717 (N_17717,N_16371,N_16255);
and U17718 (N_17718,N_15929,N_16063);
and U17719 (N_17719,N_16263,N_15892);
nand U17720 (N_17720,N_16731,N_15727);
nand U17721 (N_17721,N_16197,N_16120);
or U17722 (N_17722,N_16269,N_16382);
xnor U17723 (N_17723,N_16086,N_16074);
nor U17724 (N_17724,N_16361,N_16075);
nand U17725 (N_17725,N_16569,N_16543);
nand U17726 (N_17726,N_16760,N_15612);
nand U17727 (N_17727,N_15993,N_15620);
nor U17728 (N_17728,N_15960,N_16172);
or U17729 (N_17729,N_16747,N_15861);
xor U17730 (N_17730,N_16656,N_16537);
nor U17731 (N_17731,N_16345,N_16368);
nor U17732 (N_17732,N_16490,N_15916);
xor U17733 (N_17733,N_16411,N_16235);
and U17734 (N_17734,N_15611,N_16768);
xor U17735 (N_17735,N_16144,N_16564);
or U17736 (N_17736,N_15905,N_16407);
and U17737 (N_17737,N_16759,N_16303);
nand U17738 (N_17738,N_16202,N_15882);
xor U17739 (N_17739,N_16110,N_16468);
nor U17740 (N_17740,N_16276,N_15811);
and U17741 (N_17741,N_16439,N_16493);
nor U17742 (N_17742,N_16293,N_16599);
xnor U17743 (N_17743,N_16004,N_15704);
xor U17744 (N_17744,N_16290,N_16570);
or U17745 (N_17745,N_16302,N_15980);
and U17746 (N_17746,N_15646,N_16756);
and U17747 (N_17747,N_16766,N_16347);
nand U17748 (N_17748,N_16539,N_15656);
nand U17749 (N_17749,N_15796,N_16705);
nor U17750 (N_17750,N_16500,N_16464);
or U17751 (N_17751,N_15850,N_16418);
or U17752 (N_17752,N_15602,N_15924);
nand U17753 (N_17753,N_15630,N_16460);
and U17754 (N_17754,N_16411,N_16295);
nor U17755 (N_17755,N_15958,N_16159);
and U17756 (N_17756,N_15810,N_16504);
and U17757 (N_17757,N_16357,N_16326);
and U17758 (N_17758,N_16669,N_15714);
nand U17759 (N_17759,N_16547,N_15627);
nor U17760 (N_17760,N_15891,N_15602);
nor U17761 (N_17761,N_16590,N_16034);
nor U17762 (N_17762,N_16326,N_16147);
xor U17763 (N_17763,N_16143,N_16692);
or U17764 (N_17764,N_16656,N_16136);
or U17765 (N_17765,N_16251,N_15758);
or U17766 (N_17766,N_16507,N_16755);
nand U17767 (N_17767,N_15659,N_15614);
nor U17768 (N_17768,N_15678,N_16546);
xnor U17769 (N_17769,N_16264,N_16685);
nor U17770 (N_17770,N_15645,N_16111);
or U17771 (N_17771,N_16286,N_15791);
nor U17772 (N_17772,N_15843,N_16771);
or U17773 (N_17773,N_16461,N_15851);
xor U17774 (N_17774,N_15864,N_16705);
nand U17775 (N_17775,N_16535,N_15815);
nand U17776 (N_17776,N_15701,N_16122);
xnor U17777 (N_17777,N_16620,N_15779);
nor U17778 (N_17778,N_16139,N_16246);
or U17779 (N_17779,N_16080,N_15825);
nand U17780 (N_17780,N_15603,N_16317);
nor U17781 (N_17781,N_16583,N_16784);
nand U17782 (N_17782,N_16230,N_15906);
nor U17783 (N_17783,N_16343,N_16393);
nor U17784 (N_17784,N_16266,N_16278);
or U17785 (N_17785,N_16534,N_16317);
and U17786 (N_17786,N_16402,N_16661);
xnor U17787 (N_17787,N_15784,N_16336);
nand U17788 (N_17788,N_16481,N_15984);
nand U17789 (N_17789,N_15808,N_16301);
nand U17790 (N_17790,N_15927,N_16313);
xor U17791 (N_17791,N_15794,N_16278);
nor U17792 (N_17792,N_15964,N_15737);
and U17793 (N_17793,N_15858,N_15930);
and U17794 (N_17794,N_16528,N_16590);
or U17795 (N_17795,N_16344,N_16515);
or U17796 (N_17796,N_16145,N_16094);
or U17797 (N_17797,N_16604,N_16003);
or U17798 (N_17798,N_16233,N_16188);
xnor U17799 (N_17799,N_15981,N_15796);
nand U17800 (N_17800,N_16709,N_16120);
nand U17801 (N_17801,N_16555,N_16210);
xnor U17802 (N_17802,N_16642,N_15947);
or U17803 (N_17803,N_15787,N_15771);
xor U17804 (N_17804,N_15823,N_16793);
or U17805 (N_17805,N_15617,N_15658);
or U17806 (N_17806,N_16578,N_15850);
xnor U17807 (N_17807,N_15952,N_15808);
nand U17808 (N_17808,N_15649,N_16638);
xnor U17809 (N_17809,N_16071,N_16088);
nor U17810 (N_17810,N_16694,N_15748);
xor U17811 (N_17811,N_16300,N_15722);
or U17812 (N_17812,N_16574,N_15752);
and U17813 (N_17813,N_16734,N_15906);
and U17814 (N_17814,N_15775,N_16265);
xor U17815 (N_17815,N_15906,N_16252);
and U17816 (N_17816,N_16120,N_16208);
and U17817 (N_17817,N_15973,N_15784);
or U17818 (N_17818,N_15655,N_15604);
and U17819 (N_17819,N_16719,N_15720);
nand U17820 (N_17820,N_16324,N_16309);
or U17821 (N_17821,N_16179,N_16191);
and U17822 (N_17822,N_16676,N_15827);
nor U17823 (N_17823,N_16192,N_16345);
nand U17824 (N_17824,N_16636,N_15981);
or U17825 (N_17825,N_15624,N_16131);
xor U17826 (N_17826,N_15787,N_15850);
and U17827 (N_17827,N_16311,N_16795);
nand U17828 (N_17828,N_16757,N_16064);
xor U17829 (N_17829,N_15607,N_16165);
xnor U17830 (N_17830,N_15745,N_16456);
nand U17831 (N_17831,N_16232,N_16409);
or U17832 (N_17832,N_15888,N_15765);
xnor U17833 (N_17833,N_16787,N_15687);
xnor U17834 (N_17834,N_15932,N_15984);
or U17835 (N_17835,N_16795,N_16286);
xor U17836 (N_17836,N_15774,N_15700);
xnor U17837 (N_17837,N_16392,N_16319);
nor U17838 (N_17838,N_16560,N_15717);
or U17839 (N_17839,N_15891,N_16088);
xnor U17840 (N_17840,N_15828,N_16588);
nand U17841 (N_17841,N_16065,N_16248);
and U17842 (N_17842,N_15746,N_16696);
nand U17843 (N_17843,N_16624,N_16424);
or U17844 (N_17844,N_16126,N_16671);
nand U17845 (N_17845,N_15872,N_16696);
nand U17846 (N_17846,N_16094,N_15646);
nand U17847 (N_17847,N_15916,N_15998);
and U17848 (N_17848,N_15954,N_16292);
nor U17849 (N_17849,N_16147,N_16384);
xor U17850 (N_17850,N_15978,N_16731);
nor U17851 (N_17851,N_15650,N_16145);
xnor U17852 (N_17852,N_16633,N_16272);
xor U17853 (N_17853,N_16302,N_15775);
nor U17854 (N_17854,N_15853,N_16418);
or U17855 (N_17855,N_16537,N_16412);
and U17856 (N_17856,N_16702,N_16575);
nor U17857 (N_17857,N_16665,N_15758);
or U17858 (N_17858,N_16622,N_16663);
nor U17859 (N_17859,N_16747,N_16386);
nor U17860 (N_17860,N_16380,N_15670);
nand U17861 (N_17861,N_15892,N_16086);
nor U17862 (N_17862,N_16185,N_16739);
and U17863 (N_17863,N_16470,N_15810);
nor U17864 (N_17864,N_16532,N_16638);
nand U17865 (N_17865,N_15995,N_16662);
nor U17866 (N_17866,N_16366,N_16156);
xnor U17867 (N_17867,N_15639,N_16118);
and U17868 (N_17868,N_16045,N_16599);
and U17869 (N_17869,N_16498,N_16180);
nor U17870 (N_17870,N_16544,N_16269);
or U17871 (N_17871,N_16504,N_16731);
or U17872 (N_17872,N_16044,N_16657);
xor U17873 (N_17873,N_16481,N_16650);
nand U17874 (N_17874,N_16284,N_16627);
nor U17875 (N_17875,N_16614,N_16011);
and U17876 (N_17876,N_15822,N_16744);
and U17877 (N_17877,N_15876,N_16627);
nor U17878 (N_17878,N_16421,N_16208);
and U17879 (N_17879,N_16028,N_16520);
nor U17880 (N_17880,N_16646,N_15886);
nor U17881 (N_17881,N_16287,N_16342);
xor U17882 (N_17882,N_15941,N_15721);
nand U17883 (N_17883,N_16254,N_16680);
nand U17884 (N_17884,N_15676,N_16268);
nor U17885 (N_17885,N_16493,N_16380);
xnor U17886 (N_17886,N_16628,N_16655);
nor U17887 (N_17887,N_16296,N_16598);
xor U17888 (N_17888,N_16483,N_15847);
xnor U17889 (N_17889,N_15964,N_16345);
nor U17890 (N_17890,N_16693,N_16481);
and U17891 (N_17891,N_16216,N_16524);
nor U17892 (N_17892,N_15937,N_15602);
nand U17893 (N_17893,N_15775,N_16107);
nor U17894 (N_17894,N_16226,N_15791);
nor U17895 (N_17895,N_15957,N_16334);
xnor U17896 (N_17896,N_15908,N_16169);
and U17897 (N_17897,N_16402,N_16787);
nor U17898 (N_17898,N_15850,N_16509);
nand U17899 (N_17899,N_15988,N_16445);
and U17900 (N_17900,N_15880,N_15988);
nor U17901 (N_17901,N_16103,N_16630);
and U17902 (N_17902,N_15634,N_16705);
or U17903 (N_17903,N_16789,N_16735);
or U17904 (N_17904,N_16586,N_16698);
nor U17905 (N_17905,N_16027,N_16322);
xnor U17906 (N_17906,N_16348,N_15603);
and U17907 (N_17907,N_15714,N_16391);
and U17908 (N_17908,N_16410,N_15837);
xor U17909 (N_17909,N_15728,N_16516);
xnor U17910 (N_17910,N_16783,N_15860);
xnor U17911 (N_17911,N_15955,N_15720);
and U17912 (N_17912,N_15617,N_16093);
nor U17913 (N_17913,N_15827,N_15953);
or U17914 (N_17914,N_16639,N_15958);
or U17915 (N_17915,N_16290,N_15786);
and U17916 (N_17916,N_15969,N_15958);
nor U17917 (N_17917,N_15888,N_15786);
nor U17918 (N_17918,N_15988,N_16665);
nand U17919 (N_17919,N_15928,N_16445);
xor U17920 (N_17920,N_15924,N_16409);
and U17921 (N_17921,N_16552,N_15791);
nand U17922 (N_17922,N_16328,N_15809);
nand U17923 (N_17923,N_15789,N_15675);
or U17924 (N_17924,N_16196,N_16267);
and U17925 (N_17925,N_16591,N_16560);
nor U17926 (N_17926,N_15691,N_16141);
nand U17927 (N_17927,N_15772,N_15958);
nand U17928 (N_17928,N_16271,N_16339);
xor U17929 (N_17929,N_16553,N_16222);
nor U17930 (N_17930,N_16430,N_16744);
or U17931 (N_17931,N_15747,N_15660);
nand U17932 (N_17932,N_16752,N_16742);
and U17933 (N_17933,N_16262,N_15830);
and U17934 (N_17934,N_15926,N_16249);
or U17935 (N_17935,N_16663,N_16132);
and U17936 (N_17936,N_16410,N_16465);
nand U17937 (N_17937,N_15879,N_16448);
xor U17938 (N_17938,N_15772,N_16611);
xor U17939 (N_17939,N_16466,N_15980);
or U17940 (N_17940,N_16484,N_15839);
nor U17941 (N_17941,N_16634,N_16254);
nand U17942 (N_17942,N_16215,N_16770);
nand U17943 (N_17943,N_16631,N_15655);
nand U17944 (N_17944,N_16658,N_16111);
nand U17945 (N_17945,N_15914,N_15981);
nand U17946 (N_17946,N_15971,N_15960);
nor U17947 (N_17947,N_16467,N_16095);
xnor U17948 (N_17948,N_16673,N_15774);
and U17949 (N_17949,N_16438,N_16057);
or U17950 (N_17950,N_15635,N_15729);
or U17951 (N_17951,N_16125,N_15964);
and U17952 (N_17952,N_16041,N_15696);
nor U17953 (N_17953,N_16645,N_15640);
nand U17954 (N_17954,N_16792,N_16162);
nand U17955 (N_17955,N_16717,N_15833);
nor U17956 (N_17956,N_16019,N_16705);
nand U17957 (N_17957,N_16172,N_15848);
nor U17958 (N_17958,N_16340,N_16661);
xnor U17959 (N_17959,N_15939,N_16641);
nor U17960 (N_17960,N_15796,N_16458);
or U17961 (N_17961,N_16589,N_15615);
and U17962 (N_17962,N_16085,N_16009);
nor U17963 (N_17963,N_16135,N_15981);
xor U17964 (N_17964,N_16726,N_16775);
xor U17965 (N_17965,N_16126,N_16641);
xnor U17966 (N_17966,N_15855,N_16027);
nand U17967 (N_17967,N_16127,N_16345);
nand U17968 (N_17968,N_16584,N_15964);
and U17969 (N_17969,N_15870,N_16691);
and U17970 (N_17970,N_15764,N_16546);
nand U17971 (N_17971,N_16430,N_15807);
xnor U17972 (N_17972,N_15636,N_16419);
or U17973 (N_17973,N_16587,N_16138);
and U17974 (N_17974,N_16556,N_16796);
xor U17975 (N_17975,N_15748,N_16479);
and U17976 (N_17976,N_16347,N_16407);
xnor U17977 (N_17977,N_16347,N_16697);
nand U17978 (N_17978,N_16288,N_16263);
and U17979 (N_17979,N_15999,N_15760);
or U17980 (N_17980,N_16324,N_16788);
xnor U17981 (N_17981,N_16132,N_15940);
xor U17982 (N_17982,N_16242,N_16503);
nor U17983 (N_17983,N_15961,N_15827);
nand U17984 (N_17984,N_15994,N_16609);
nor U17985 (N_17985,N_16607,N_16528);
nor U17986 (N_17986,N_15915,N_16396);
nand U17987 (N_17987,N_15707,N_16579);
or U17988 (N_17988,N_16795,N_15916);
nand U17989 (N_17989,N_15820,N_15782);
xnor U17990 (N_17990,N_16485,N_15910);
and U17991 (N_17991,N_16167,N_16103);
and U17992 (N_17992,N_16121,N_16506);
nor U17993 (N_17993,N_15862,N_15744);
nor U17994 (N_17994,N_15840,N_16136);
xor U17995 (N_17995,N_16075,N_16427);
nor U17996 (N_17996,N_16684,N_15695);
and U17997 (N_17997,N_16736,N_16524);
and U17998 (N_17998,N_16412,N_15816);
nor U17999 (N_17999,N_16113,N_15719);
nor U18000 (N_18000,N_16873,N_17907);
nor U18001 (N_18001,N_17580,N_17596);
nand U18002 (N_18002,N_17105,N_17024);
nand U18003 (N_18003,N_16939,N_17204);
xnor U18004 (N_18004,N_16947,N_17566);
and U18005 (N_18005,N_17794,N_17952);
xor U18006 (N_18006,N_17149,N_17466);
xnor U18007 (N_18007,N_16833,N_16837);
and U18008 (N_18008,N_17749,N_16842);
nand U18009 (N_18009,N_17012,N_17525);
nor U18010 (N_18010,N_17348,N_17927);
and U18011 (N_18011,N_17064,N_17916);
and U18012 (N_18012,N_17038,N_17751);
nand U18013 (N_18013,N_17013,N_17532);
xor U18014 (N_18014,N_16806,N_17948);
xor U18015 (N_18015,N_17023,N_17594);
xnor U18016 (N_18016,N_17787,N_17186);
and U18017 (N_18017,N_17263,N_17944);
and U18018 (N_18018,N_16908,N_17392);
nor U18019 (N_18019,N_16984,N_17576);
nand U18020 (N_18020,N_17494,N_17543);
xor U18021 (N_18021,N_17557,N_17837);
and U18022 (N_18022,N_17774,N_17314);
nor U18023 (N_18023,N_17715,N_17334);
nand U18024 (N_18024,N_17175,N_17694);
and U18025 (N_18025,N_17299,N_17629);
or U18026 (N_18026,N_17193,N_17757);
nand U18027 (N_18027,N_17841,N_16962);
or U18028 (N_18028,N_17981,N_17853);
or U18029 (N_18029,N_17535,N_16825);
or U18030 (N_18030,N_17579,N_17796);
nor U18031 (N_18031,N_17605,N_17914);
and U18032 (N_18032,N_17360,N_17830);
nor U18033 (N_18033,N_16860,N_17262);
nor U18034 (N_18034,N_17848,N_17681);
nand U18035 (N_18035,N_17985,N_17875);
nor U18036 (N_18036,N_16988,N_16986);
and U18037 (N_18037,N_17975,N_17775);
nor U18038 (N_18038,N_17992,N_16994);
nor U18039 (N_18039,N_17808,N_17635);
and U18040 (N_18040,N_17705,N_17316);
and U18041 (N_18041,N_17849,N_17281);
nor U18042 (N_18042,N_17219,N_16802);
xor U18043 (N_18043,N_17955,N_17147);
nand U18044 (N_18044,N_17998,N_17061);
nand U18045 (N_18045,N_16999,N_17212);
and U18046 (N_18046,N_17523,N_16901);
xor U18047 (N_18047,N_17722,N_17154);
nand U18048 (N_18048,N_17156,N_16876);
xnor U18049 (N_18049,N_17151,N_17721);
or U18050 (N_18050,N_17781,N_17202);
and U18051 (N_18051,N_17055,N_16905);
xor U18052 (N_18052,N_17936,N_17469);
xor U18053 (N_18053,N_17168,N_17832);
or U18054 (N_18054,N_17960,N_17661);
and U18055 (N_18055,N_17941,N_16808);
nand U18056 (N_18056,N_17477,N_17111);
nand U18057 (N_18057,N_17329,N_17620);
nand U18058 (N_18058,N_17686,N_16963);
or U18059 (N_18059,N_16928,N_17044);
nor U18060 (N_18060,N_17632,N_17009);
nand U18061 (N_18061,N_17707,N_17275);
and U18062 (N_18062,N_17199,N_17207);
xor U18063 (N_18063,N_17593,N_16869);
or U18064 (N_18064,N_17685,N_17339);
and U18065 (N_18065,N_17083,N_17714);
or U18066 (N_18066,N_17654,N_17835);
or U18067 (N_18067,N_17609,N_17133);
nand U18068 (N_18068,N_17652,N_17903);
nor U18069 (N_18069,N_17514,N_17834);
and U18070 (N_18070,N_17935,N_17324);
xnor U18071 (N_18071,N_17607,N_17759);
and U18072 (N_18072,N_17585,N_17229);
and U18073 (N_18073,N_17291,N_17860);
and U18074 (N_18074,N_17045,N_17847);
nand U18075 (N_18075,N_17724,N_16971);
nor U18076 (N_18076,N_17448,N_17277);
or U18077 (N_18077,N_17239,N_17542);
xnor U18078 (N_18078,N_16820,N_17531);
and U18079 (N_18079,N_16840,N_17288);
xnor U18080 (N_18080,N_17185,N_17420);
nor U18081 (N_18081,N_17919,N_17565);
and U18082 (N_18082,N_17822,N_17490);
nand U18083 (N_18083,N_17273,N_16867);
nor U18084 (N_18084,N_17245,N_17079);
nor U18085 (N_18085,N_17192,N_17680);
xor U18086 (N_18086,N_17592,N_17457);
or U18087 (N_18087,N_17340,N_16883);
xor U18088 (N_18088,N_17588,N_17416);
or U18089 (N_18089,N_17280,N_16979);
nand U18090 (N_18090,N_17399,N_17268);
nor U18091 (N_18091,N_17062,N_17125);
xnor U18092 (N_18092,N_17816,N_17638);
nor U18093 (N_18093,N_17740,N_17495);
or U18094 (N_18094,N_16903,N_17300);
nor U18095 (N_18095,N_17896,N_17571);
or U18096 (N_18096,N_17616,N_17028);
nand U18097 (N_18097,N_17351,N_17518);
nor U18098 (N_18098,N_17224,N_17918);
nand U18099 (N_18099,N_17226,N_17929);
nor U18100 (N_18100,N_17379,N_17556);
or U18101 (N_18101,N_17797,N_17536);
xnor U18102 (N_18102,N_16991,N_17122);
or U18103 (N_18103,N_16951,N_17790);
and U18104 (N_18104,N_17406,N_17421);
or U18105 (N_18105,N_17545,N_17615);
nor U18106 (N_18106,N_17396,N_17027);
and U18107 (N_18107,N_17695,N_17109);
and U18108 (N_18108,N_17793,N_17780);
nand U18109 (N_18109,N_17075,N_16940);
and U18110 (N_18110,N_17754,N_17387);
and U18111 (N_18111,N_17890,N_17252);
or U18112 (N_18112,N_17343,N_16900);
and U18113 (N_18113,N_17684,N_17672);
or U18114 (N_18114,N_17561,N_17323);
nand U18115 (N_18115,N_16865,N_17679);
nand U18116 (N_18116,N_17934,N_17957);
xor U18117 (N_18117,N_17050,N_17641);
nor U18118 (N_18118,N_16987,N_17519);
and U18119 (N_18119,N_16923,N_17368);
nor U18120 (N_18120,N_17104,N_17866);
xor U18121 (N_18121,N_17507,N_17008);
nor U18122 (N_18122,N_17237,N_17559);
nand U18123 (N_18123,N_17713,N_17209);
and U18124 (N_18124,N_17655,N_17215);
or U18125 (N_18125,N_17491,N_17692);
or U18126 (N_18126,N_17459,N_17879);
xnor U18127 (N_18127,N_17259,N_17824);
nand U18128 (N_18128,N_16972,N_17270);
nor U18129 (N_18129,N_16936,N_17395);
nor U18130 (N_18130,N_17385,N_17389);
and U18131 (N_18131,N_17931,N_17337);
and U18132 (N_18132,N_17123,N_17538);
nand U18133 (N_18133,N_17070,N_16879);
and U18134 (N_18134,N_17984,N_16980);
nand U18135 (N_18135,N_17446,N_17746);
xor U18136 (N_18136,N_17434,N_17547);
nor U18137 (N_18137,N_16834,N_16841);
or U18138 (N_18138,N_17068,N_17319);
xor U18139 (N_18139,N_17905,N_17372);
and U18140 (N_18140,N_17789,N_17294);
xor U18141 (N_18141,N_17014,N_17806);
nor U18142 (N_18142,N_17241,N_17658);
or U18143 (N_18143,N_17540,N_17529);
xnor U18144 (N_18144,N_17731,N_16891);
xnor U18145 (N_18145,N_17912,N_17814);
nand U18146 (N_18146,N_17190,N_17520);
xnor U18147 (N_18147,N_16998,N_17206);
nor U18148 (N_18148,N_17110,N_16819);
and U18149 (N_18149,N_17465,N_17819);
nand U18150 (N_18150,N_17115,N_16911);
nor U18151 (N_18151,N_17058,N_17622);
nand U18152 (N_18152,N_16904,N_16843);
or U18153 (N_18153,N_17167,N_16890);
nand U18154 (N_18154,N_17312,N_17455);
and U18155 (N_18155,N_17287,N_16956);
and U18156 (N_18156,N_17902,N_17646);
or U18157 (N_18157,N_17327,N_17753);
and U18158 (N_18158,N_17969,N_17765);
or U18159 (N_18159,N_17102,N_16858);
xnor U18160 (N_18160,N_17415,N_17234);
xnor U18161 (N_18161,N_17388,N_17255);
xor U18162 (N_18162,N_16801,N_16823);
xnor U18163 (N_18163,N_17002,N_17898);
nand U18164 (N_18164,N_17437,N_17997);
xnor U18165 (N_18165,N_17733,N_17682);
nor U18166 (N_18166,N_16992,N_17251);
xnor U18167 (N_18167,N_17698,N_17893);
xor U18168 (N_18168,N_17369,N_17601);
nor U18169 (N_18169,N_17137,N_17712);
nor U18170 (N_18170,N_17030,N_17864);
and U18171 (N_18171,N_17475,N_17748);
nor U18172 (N_18172,N_16946,N_17553);
or U18173 (N_18173,N_17752,N_17894);
and U18174 (N_18174,N_16927,N_17656);
nor U18175 (N_18175,N_17815,N_17026);
nor U18176 (N_18176,N_17021,N_17092);
nand U18177 (N_18177,N_17569,N_17498);
and U18178 (N_18178,N_17552,N_17135);
and U18179 (N_18179,N_17600,N_17584);
and U18180 (N_18180,N_17513,N_17054);
xor U18181 (N_18181,N_17230,N_17106);
nor U18182 (N_18182,N_17734,N_17924);
and U18183 (N_18183,N_17842,N_17155);
nand U18184 (N_18184,N_17820,N_17803);
nand U18185 (N_18185,N_17625,N_17745);
or U18186 (N_18186,N_17729,N_17143);
and U18187 (N_18187,N_17423,N_17769);
and U18188 (N_18188,N_16916,N_17057);
nand U18189 (N_18189,N_17160,N_17505);
nor U18190 (N_18190,N_17967,N_17333);
xor U18191 (N_18191,N_17511,N_17589);
and U18192 (N_18192,N_17180,N_17930);
and U18193 (N_18193,N_17474,N_17227);
and U18194 (N_18194,N_17476,N_17425);
xnor U18195 (N_18195,N_16982,N_16978);
nor U18196 (N_18196,N_17693,N_17791);
nand U18197 (N_18197,N_17611,N_17077);
xnor U18198 (N_18198,N_17770,N_17739);
xnor U18199 (N_18199,N_17763,N_17108);
and U18200 (N_18200,N_16934,N_17639);
xor U18201 (N_18201,N_17619,N_17315);
nand U18202 (N_18202,N_17517,N_16824);
nand U18203 (N_18203,N_16925,N_17440);
and U18204 (N_18204,N_17481,N_17855);
xnor U18205 (N_18205,N_17242,N_17604);
or U18206 (N_18206,N_17318,N_17341);
nor U18207 (N_18207,N_17376,N_17492);
or U18208 (N_18208,N_17696,N_16969);
xnor U18209 (N_18209,N_17979,N_17673);
xor U18210 (N_18210,N_17216,N_17628);
nor U18211 (N_18211,N_16881,N_17405);
and U18212 (N_18212,N_17362,N_17117);
nor U18213 (N_18213,N_17331,N_17441);
or U18214 (N_18214,N_17524,N_17456);
nor U18215 (N_18215,N_17301,N_17867);
or U18216 (N_18216,N_16870,N_17537);
or U18217 (N_18217,N_17886,N_17954);
xor U18218 (N_18218,N_17210,N_17412);
or U18219 (N_18219,N_17962,N_17188);
and U18220 (N_18220,N_17617,N_17355);
and U18221 (N_18221,N_17195,N_17141);
nand U18222 (N_18222,N_17786,N_17627);
nor U18223 (N_18223,N_17504,N_17506);
and U18224 (N_18224,N_17873,N_17272);
or U18225 (N_18225,N_17031,N_17131);
xnor U18226 (N_18226,N_17874,N_17484);
or U18227 (N_18227,N_17640,N_17451);
or U18228 (N_18228,N_17303,N_17119);
nor U18229 (N_18229,N_17982,N_17183);
or U18230 (N_18230,N_17309,N_17403);
xnor U18231 (N_18231,N_17450,N_17478);
xor U18232 (N_18232,N_17367,N_16892);
xor U18233 (N_18233,N_17238,N_17839);
xor U18234 (N_18234,N_17101,N_17633);
and U18235 (N_18235,N_17427,N_17727);
and U18236 (N_18236,N_17688,N_17699);
nand U18237 (N_18237,N_17845,N_16924);
nand U18238 (N_18238,N_17097,N_17560);
nand U18239 (N_18239,N_17868,N_17583);
xor U18240 (N_18240,N_17697,N_17900);
and U18241 (N_18241,N_16844,N_17533);
nor U18242 (N_18242,N_17244,N_17282);
nand U18243 (N_18243,N_17232,N_17431);
or U18244 (N_18244,N_17438,N_17939);
nand U18245 (N_18245,N_17426,N_16929);
and U18246 (N_18246,N_17349,N_17574);
or U18247 (N_18247,N_17701,N_17043);
or U18248 (N_18248,N_17813,N_17452);
and U18249 (N_18249,N_17503,N_17771);
xnor U18250 (N_18250,N_16800,N_17366);
nor U18251 (N_18251,N_17920,N_16831);
or U18252 (N_18252,N_17821,N_17591);
xor U18253 (N_18253,N_17338,N_17500);
xor U18254 (N_18254,N_17735,N_16915);
xor U18255 (N_18255,N_17443,N_17643);
and U18256 (N_18256,N_16889,N_17926);
and U18257 (N_18257,N_16897,N_17410);
xnor U18258 (N_18258,N_17080,N_17090);
xnor U18259 (N_18259,N_17674,N_17218);
and U18260 (N_18260,N_17597,N_17269);
and U18261 (N_18261,N_17100,N_17140);
nor U18262 (N_18262,N_17463,N_17851);
or U18263 (N_18263,N_17169,N_17827);
and U18264 (N_18264,N_16931,N_17074);
xnor U18265 (N_18265,N_17187,N_17884);
or U18266 (N_18266,N_17785,N_16866);
or U18267 (N_18267,N_17419,N_17980);
xor U18268 (N_18268,N_16826,N_17240);
or U18269 (N_18269,N_17728,N_17171);
xor U18270 (N_18270,N_17810,N_17302);
or U18271 (N_18271,N_17346,N_17034);
nand U18272 (N_18272,N_17800,N_17677);
or U18273 (N_18273,N_17634,N_17081);
xor U18274 (N_18274,N_17344,N_16909);
or U18275 (N_18275,N_17648,N_17678);
xor U18276 (N_18276,N_17788,N_17250);
nand U18277 (N_18277,N_17046,N_16964);
nand U18278 (N_18278,N_17805,N_17342);
and U18279 (N_18279,N_17949,N_17052);
or U18280 (N_18280,N_17345,N_17235);
or U18281 (N_18281,N_17888,N_17606);
and U18282 (N_18282,N_16933,N_17430);
nor U18283 (N_18283,N_17161,N_17243);
and U18284 (N_18284,N_16974,N_17139);
and U18285 (N_18285,N_17144,N_17248);
nor U18286 (N_18286,N_16938,N_17809);
nor U18287 (N_18287,N_17741,N_17153);
and U18288 (N_18288,N_17764,N_17700);
or U18289 (N_18289,N_17462,N_17332);
and U18290 (N_18290,N_17354,N_17295);
nor U18291 (N_18291,N_17082,N_16863);
and U18292 (N_18292,N_17947,N_16828);
nand U18293 (N_18293,N_16850,N_17099);
nand U18294 (N_18294,N_17817,N_17717);
xnor U18295 (N_18295,N_17899,N_17464);
or U18296 (N_18296,N_17356,N_17471);
and U18297 (N_18297,N_17065,N_17653);
and U18298 (N_18298,N_16912,N_16937);
and U18299 (N_18299,N_16849,N_17132);
xor U18300 (N_18300,N_17577,N_16935);
or U18301 (N_18301,N_17482,N_16910);
nand U18302 (N_18302,N_17130,N_17095);
nand U18303 (N_18303,N_17363,N_17546);
and U18304 (N_18304,N_17278,N_17084);
and U18305 (N_18305,N_17792,N_17378);
nand U18306 (N_18306,N_17675,N_16948);
nand U18307 (N_18307,N_17965,N_17370);
nor U18308 (N_18308,N_16875,N_16817);
or U18309 (N_18309,N_17779,N_17623);
xor U18310 (N_18310,N_17689,N_16906);
and U18311 (N_18311,N_17078,N_16965);
nor U18312 (N_18312,N_17222,N_16932);
nand U18313 (N_18313,N_17863,N_17937);
or U18314 (N_18314,N_17447,N_17196);
nor U18315 (N_18315,N_17650,N_17308);
nand U18316 (N_18316,N_17129,N_17995);
or U18317 (N_18317,N_17178,N_17214);
nand U18318 (N_18318,N_17386,N_16966);
xor U18319 (N_18319,N_17066,N_17758);
xor U18320 (N_18320,N_17157,N_17003);
xnor U18321 (N_18321,N_17258,N_17005);
and U18322 (N_18322,N_17645,N_16917);
nand U18323 (N_18323,N_16861,N_17124);
xor U18324 (N_18324,N_17439,N_17261);
nand U18325 (N_18325,N_17946,N_16815);
nand U18326 (N_18326,N_17019,N_17534);
and U18327 (N_18327,N_17823,N_16914);
and U18328 (N_18328,N_17691,N_17993);
and U18329 (N_18329,N_17750,N_17549);
and U18330 (N_18330,N_16955,N_17148);
nand U18331 (N_18331,N_17307,N_16821);
nand U18332 (N_18332,N_16885,N_16894);
or U18333 (N_18333,N_17198,N_17709);
xor U18334 (N_18334,N_16997,N_17858);
and U18335 (N_18335,N_17554,N_17558);
and U18336 (N_18336,N_17444,N_16822);
and U18337 (N_18337,N_17970,N_17225);
xnor U18338 (N_18338,N_17550,N_17357);
xor U18339 (N_18339,N_17040,N_17578);
nand U18340 (N_18340,N_17564,N_17649);
and U18341 (N_18341,N_16827,N_16830);
and U18342 (N_18342,N_17467,N_17671);
nor U18343 (N_18343,N_17901,N_16967);
or U18344 (N_18344,N_17121,N_17906);
or U18345 (N_18345,N_17398,N_16942);
xnor U18346 (N_18346,N_16816,N_16989);
and U18347 (N_18347,N_17966,N_17710);
or U18348 (N_18348,N_17666,N_17271);
or U18349 (N_18349,N_17502,N_16859);
and U18350 (N_18350,N_16958,N_16913);
and U18351 (N_18351,N_17613,N_17742);
and U18352 (N_18352,N_17913,N_17795);
nand U18353 (N_18353,N_16871,N_16968);
nor U18354 (N_18354,N_17850,N_17350);
nand U18355 (N_18355,N_17726,N_17220);
nor U18356 (N_18356,N_17973,N_16945);
nor U18357 (N_18357,N_17644,N_17397);
nor U18358 (N_18358,N_17048,N_17544);
nand U18359 (N_18359,N_17166,N_17266);
nand U18360 (N_18360,N_17497,N_17371);
nor U18361 (N_18361,N_16898,N_17018);
nand U18362 (N_18362,N_17449,N_17411);
xor U18363 (N_18363,N_17223,N_16954);
nand U18364 (N_18364,N_17811,N_17630);
or U18365 (N_18365,N_17732,N_17516);
and U18366 (N_18366,N_16853,N_16976);
nor U18367 (N_18367,N_16977,N_17022);
or U18368 (N_18368,N_17381,N_17798);
nand U18369 (N_18369,N_17784,N_17310);
or U18370 (N_18370,N_17059,N_17383);
or U18371 (N_18371,N_17076,N_17265);
nand U18372 (N_18372,N_17833,N_16839);
or U18373 (N_18373,N_16835,N_17352);
xor U18374 (N_18374,N_17487,N_17828);
or U18375 (N_18375,N_16926,N_17932);
nor U18376 (N_18376,N_16810,N_17642);
and U18377 (N_18377,N_17994,N_17723);
and U18378 (N_18378,N_17407,N_17000);
and U18379 (N_18379,N_17624,N_17923);
or U18380 (N_18380,N_17767,N_17877);
or U18381 (N_18381,N_17353,N_17088);
xnor U18382 (N_18382,N_17568,N_16922);
nor U18383 (N_18383,N_17881,N_17460);
nand U18384 (N_18384,N_17861,N_17203);
or U18385 (N_18385,N_17826,N_17736);
nand U18386 (N_18386,N_16868,N_17401);
and U18387 (N_18387,N_17473,N_16949);
or U18388 (N_18388,N_17610,N_16872);
and U18389 (N_18389,N_16895,N_17608);
nand U18390 (N_18390,N_17683,N_17246);
nor U18391 (N_18391,N_17174,N_17961);
nand U18392 (N_18392,N_17114,N_16851);
nand U18393 (N_18393,N_17404,N_17486);
nor U18394 (N_18394,N_16996,N_17762);
nor U18395 (N_18395,N_17085,N_17172);
nand U18396 (N_18396,N_17660,N_17442);
or U18397 (N_18397,N_17221,N_17335);
or U18398 (N_18398,N_17205,N_17871);
xnor U18399 (N_18399,N_17690,N_17637);
and U18400 (N_18400,N_17951,N_17096);
xor U18401 (N_18401,N_17041,N_17181);
nor U18402 (N_18402,N_17807,N_17772);
nand U18403 (N_18403,N_16959,N_16957);
nor U18404 (N_18404,N_17020,N_17093);
nor U18405 (N_18405,N_16930,N_17522);
nor U18406 (N_18406,N_17159,N_17321);
nand U18407 (N_18407,N_16856,N_17971);
nand U18408 (N_18408,N_17164,N_17029);
and U18409 (N_18409,N_17976,N_17508);
xnor U18410 (N_18410,N_17445,N_17428);
nor U18411 (N_18411,N_16941,N_17283);
nand U18412 (N_18412,N_17483,N_17977);
nand U18413 (N_18413,N_17778,N_17777);
nand U18414 (N_18414,N_17528,N_17687);
nand U18415 (N_18415,N_17978,N_17359);
xnor U18416 (N_18416,N_17162,N_17933);
nand U18417 (N_18417,N_17738,N_17662);
xnor U18418 (N_18418,N_17182,N_17602);
or U18419 (N_18419,N_17213,N_17004);
xor U18420 (N_18420,N_17422,N_17704);
nor U18421 (N_18421,N_17264,N_17136);
and U18422 (N_18422,N_17328,N_17865);
xnor U18423 (N_18423,N_17959,N_17663);
nor U18424 (N_18424,N_17211,N_17454);
nor U18425 (N_18425,N_17152,N_17988);
xnor U18426 (N_18426,N_17720,N_17501);
xnor U18427 (N_18427,N_17711,N_17260);
or U18428 (N_18428,N_17856,N_17228);
or U18429 (N_18429,N_16896,N_17468);
or U18430 (N_18430,N_17703,N_17032);
xor U18431 (N_18431,N_17072,N_17107);
nand U18432 (N_18432,N_17067,N_17541);
or U18433 (N_18433,N_16848,N_17113);
nand U18434 (N_18434,N_17825,N_17526);
nor U18435 (N_18435,N_17317,N_17485);
nor U18436 (N_18436,N_17876,N_16952);
xor U18437 (N_18437,N_17049,N_17581);
nor U18438 (N_18438,N_17963,N_16953);
and U18439 (N_18439,N_16864,N_17279);
and U18440 (N_18440,N_17293,N_17840);
nand U18441 (N_18441,N_17968,N_17891);
and U18442 (N_18442,N_17163,N_17567);
or U18443 (N_18443,N_16852,N_17480);
xnor U18444 (N_18444,N_17458,N_17882);
nor U18445 (N_18445,N_17033,N_17725);
nor U18446 (N_18446,N_17200,N_17016);
and U18447 (N_18447,N_17737,N_17852);
or U18448 (N_18448,N_17393,N_17669);
or U18449 (N_18449,N_16803,N_17313);
nand U18450 (N_18450,N_17173,N_17320);
nand U18451 (N_18451,N_17037,N_17925);
and U18452 (N_18452,N_17897,N_17380);
nor U18453 (N_18453,N_17184,N_17756);
or U18454 (N_18454,N_17880,N_17285);
xnor U18455 (N_18455,N_17194,N_17702);
or U18456 (N_18456,N_17290,N_17358);
xor U18457 (N_18457,N_17414,N_17436);
and U18458 (N_18458,N_17659,N_16981);
nand U18459 (N_18459,N_17094,N_17289);
or U18460 (N_18460,N_17986,N_17667);
or U18461 (N_18461,N_17292,N_17253);
or U18462 (N_18462,N_17394,N_17869);
nand U18463 (N_18463,N_17938,N_17296);
or U18464 (N_18464,N_17257,N_17035);
or U18465 (N_18465,N_17744,N_17073);
xor U18466 (N_18466,N_17562,N_17208);
nor U18467 (N_18467,N_17010,N_17413);
and U18468 (N_18468,N_17563,N_17249);
nor U18469 (N_18469,N_16944,N_16862);
nor U18470 (N_18470,N_17036,N_17719);
nand U18471 (N_18471,N_17461,N_16995);
nor U18472 (N_18472,N_17138,N_16857);
nor U18473 (N_18473,N_17964,N_16813);
or U18474 (N_18474,N_17862,N_16893);
nor U18475 (N_18475,N_17972,N_17595);
xnor U18476 (N_18476,N_17887,N_17325);
xor U18477 (N_18477,N_17015,N_17176);
xor U18478 (N_18478,N_17857,N_16921);
and U18479 (N_18479,N_17470,N_17274);
or U18480 (N_18480,N_16907,N_16832);
nand U18481 (N_18481,N_17958,N_17112);
nor U18482 (N_18482,N_17063,N_17071);
nand U18483 (N_18483,N_17829,N_17527);
nor U18484 (N_18484,N_17373,N_17170);
nor U18485 (N_18485,N_16811,N_17311);
or U18486 (N_18486,N_17618,N_17911);
nor U18487 (N_18487,N_17165,N_17942);
or U18488 (N_18488,N_16818,N_17472);
or U18489 (N_18489,N_16918,N_17991);
and U18490 (N_18490,N_17217,N_17391);
or U18491 (N_18491,N_17120,N_16836);
nand U18492 (N_18492,N_17515,N_17665);
nand U18493 (N_18493,N_17989,N_17651);
nand U18494 (N_18494,N_17818,N_17676);
or U18495 (N_18495,N_17718,N_17051);
or U18496 (N_18496,N_17776,N_16960);
or U18497 (N_18497,N_17429,N_17706);
nand U18498 (N_18498,N_17956,N_16814);
nand U18499 (N_18499,N_17773,N_17400);
or U18500 (N_18500,N_17424,N_16970);
and U18501 (N_18501,N_17990,N_17364);
nand U18502 (N_18502,N_17843,N_17582);
and U18503 (N_18503,N_17365,N_17326);
nand U18504 (N_18504,N_17298,N_17859);
xor U18505 (N_18505,N_17996,N_17747);
and U18506 (N_18506,N_17755,N_16847);
nor U18507 (N_18507,N_17304,N_17103);
nand U18508 (N_18508,N_17512,N_17432);
or U18509 (N_18509,N_17118,N_17134);
nor U18510 (N_18510,N_17587,N_17011);
xor U18511 (N_18511,N_17042,N_17158);
nand U18512 (N_18512,N_17276,N_17760);
xor U18513 (N_18513,N_17347,N_17382);
or U18514 (N_18514,N_17586,N_17191);
nand U18515 (N_18515,N_16812,N_17039);
or U18516 (N_18516,N_17453,N_17889);
xnor U18517 (N_18517,N_17590,N_17878);
or U18518 (N_18518,N_17128,N_17730);
nor U18519 (N_18519,N_17069,N_17086);
nor U18520 (N_18520,N_17716,N_17708);
and U18521 (N_18521,N_16950,N_17390);
xnor U18522 (N_18522,N_17603,N_17831);
nor U18523 (N_18523,N_17496,N_16829);
xor U18524 (N_18524,N_17091,N_16973);
xor U18525 (N_18525,N_17007,N_17917);
xor U18526 (N_18526,N_17247,N_17499);
nand U18527 (N_18527,N_17087,N_17521);
xor U18528 (N_18528,N_17614,N_16805);
xnor U18529 (N_18529,N_16943,N_17284);
nand U18530 (N_18530,N_17885,N_17836);
nor U18531 (N_18531,N_17621,N_17987);
nor U18532 (N_18532,N_17402,N_16888);
nand U18533 (N_18533,N_17940,N_17001);
or U18534 (N_18534,N_17375,N_16809);
xnor U18535 (N_18535,N_17539,N_17626);
nand U18536 (N_18536,N_16884,N_16975);
and U18537 (N_18537,N_17922,N_17838);
xor U18538 (N_18538,N_17322,N_17053);
and U18539 (N_18539,N_17417,N_17126);
nand U18540 (N_18540,N_17572,N_17297);
nand U18541 (N_18541,N_16899,N_16919);
xnor U18542 (N_18542,N_16990,N_17197);
or U18543 (N_18543,N_17573,N_17384);
xnor U18544 (N_18544,N_17599,N_17256);
and U18545 (N_18545,N_17999,N_17636);
xor U18546 (N_18546,N_17768,N_17928);
nor U18547 (N_18547,N_17142,N_17017);
and U18548 (N_18548,N_17953,N_16993);
nor U18549 (N_18549,N_17060,N_17025);
nand U18550 (N_18550,N_16874,N_17361);
nor U18551 (N_18551,N_17409,N_17943);
or U18552 (N_18552,N_17179,N_17330);
and U18553 (N_18553,N_17915,N_17804);
nor U18554 (N_18554,N_17983,N_17575);
and U18555 (N_18555,N_17670,N_17548);
or U18556 (N_18556,N_17146,N_17904);
xnor U18557 (N_18557,N_17846,N_17267);
or U18558 (N_18558,N_17530,N_16807);
nand U18559 (N_18559,N_17761,N_17056);
or U18560 (N_18560,N_17089,N_17555);
nand U18561 (N_18561,N_16804,N_17374);
or U18562 (N_18562,N_16878,N_17201);
or U18563 (N_18563,N_17950,N_17974);
or U18564 (N_18564,N_17177,N_17892);
nor U18565 (N_18565,N_16882,N_16887);
nor U18566 (N_18566,N_17306,N_17945);
and U18567 (N_18567,N_17657,N_17612);
and U18568 (N_18568,N_17664,N_17479);
xnor U18569 (N_18569,N_17233,N_16920);
and U18570 (N_18570,N_17254,N_17435);
and U18571 (N_18571,N_17872,N_16880);
nor U18572 (N_18572,N_17551,N_17408);
xnor U18573 (N_18573,N_16985,N_17489);
or U18574 (N_18574,N_17799,N_16854);
nor U18575 (N_18575,N_17418,N_17509);
and U18576 (N_18576,N_17116,N_17286);
or U18577 (N_18577,N_17766,N_17631);
and U18578 (N_18578,N_17844,N_16838);
and U18579 (N_18579,N_17570,N_17870);
nand U18580 (N_18580,N_17908,N_17909);
nor U18581 (N_18581,N_17743,N_17801);
or U18582 (N_18582,N_17145,N_17802);
nand U18583 (N_18583,N_17493,N_17883);
nor U18584 (N_18584,N_17236,N_17510);
xor U18585 (N_18585,N_17006,N_17488);
nand U18586 (N_18586,N_16886,N_17668);
and U18587 (N_18587,N_17782,N_17231);
and U18588 (N_18588,N_17336,N_16845);
xnor U18589 (N_18589,N_17098,N_17921);
or U18590 (N_18590,N_17433,N_17189);
and U18591 (N_18591,N_17047,N_17895);
nor U18592 (N_18592,N_16902,N_16983);
xnor U18593 (N_18593,N_17910,N_16846);
and U18594 (N_18594,N_16855,N_17812);
and U18595 (N_18595,N_17598,N_16877);
nor U18596 (N_18596,N_17783,N_17854);
xnor U18597 (N_18597,N_16961,N_17305);
and U18598 (N_18598,N_17647,N_17127);
xor U18599 (N_18599,N_17377,N_17150);
or U18600 (N_18600,N_17790,N_17914);
xnor U18601 (N_18601,N_17095,N_17546);
xnor U18602 (N_18602,N_17916,N_17686);
nor U18603 (N_18603,N_17554,N_17290);
and U18604 (N_18604,N_17516,N_17595);
and U18605 (N_18605,N_16995,N_17756);
nand U18606 (N_18606,N_17774,N_17557);
and U18607 (N_18607,N_17534,N_16876);
or U18608 (N_18608,N_16896,N_16958);
and U18609 (N_18609,N_17704,N_17329);
or U18610 (N_18610,N_17863,N_17162);
or U18611 (N_18611,N_17491,N_17251);
xor U18612 (N_18612,N_17836,N_17877);
nand U18613 (N_18613,N_17079,N_17870);
and U18614 (N_18614,N_17783,N_17241);
xnor U18615 (N_18615,N_17466,N_17503);
or U18616 (N_18616,N_17685,N_17364);
nand U18617 (N_18617,N_17812,N_17136);
nand U18618 (N_18618,N_16849,N_17724);
and U18619 (N_18619,N_17934,N_17405);
or U18620 (N_18620,N_17893,N_16867);
nor U18621 (N_18621,N_17457,N_17453);
xnor U18622 (N_18622,N_17793,N_17130);
and U18623 (N_18623,N_17006,N_17824);
nor U18624 (N_18624,N_17667,N_17503);
or U18625 (N_18625,N_17738,N_17657);
xor U18626 (N_18626,N_17342,N_16818);
or U18627 (N_18627,N_17989,N_17798);
or U18628 (N_18628,N_16887,N_17135);
and U18629 (N_18629,N_17602,N_17354);
nor U18630 (N_18630,N_17103,N_17795);
xnor U18631 (N_18631,N_17094,N_17651);
xor U18632 (N_18632,N_17827,N_17065);
and U18633 (N_18633,N_17167,N_17716);
nor U18634 (N_18634,N_17974,N_17826);
xor U18635 (N_18635,N_17697,N_17039);
or U18636 (N_18636,N_16920,N_17915);
and U18637 (N_18637,N_17075,N_17727);
xnor U18638 (N_18638,N_17224,N_17638);
nand U18639 (N_18639,N_16986,N_16814);
nor U18640 (N_18640,N_17455,N_17832);
nor U18641 (N_18641,N_16940,N_17000);
or U18642 (N_18642,N_17314,N_17191);
xor U18643 (N_18643,N_17940,N_17154);
nor U18644 (N_18644,N_17123,N_17877);
or U18645 (N_18645,N_16956,N_17911);
nor U18646 (N_18646,N_16833,N_17145);
nor U18647 (N_18647,N_16840,N_17081);
nand U18648 (N_18648,N_17017,N_17337);
or U18649 (N_18649,N_17880,N_17152);
xnor U18650 (N_18650,N_17642,N_17002);
nor U18651 (N_18651,N_17704,N_17550);
xor U18652 (N_18652,N_16956,N_17816);
or U18653 (N_18653,N_17965,N_17719);
xnor U18654 (N_18654,N_17206,N_17610);
nand U18655 (N_18655,N_17604,N_17857);
nand U18656 (N_18656,N_17176,N_17721);
or U18657 (N_18657,N_17529,N_17708);
xor U18658 (N_18658,N_17397,N_17728);
nand U18659 (N_18659,N_17540,N_17816);
or U18660 (N_18660,N_17648,N_17619);
and U18661 (N_18661,N_17806,N_17921);
and U18662 (N_18662,N_17467,N_17979);
and U18663 (N_18663,N_17261,N_17340);
nor U18664 (N_18664,N_17898,N_16805);
nand U18665 (N_18665,N_16916,N_16835);
and U18666 (N_18666,N_17138,N_17814);
or U18667 (N_18667,N_17872,N_17262);
nand U18668 (N_18668,N_17666,N_17922);
xnor U18669 (N_18669,N_17820,N_17328);
or U18670 (N_18670,N_17309,N_17478);
nand U18671 (N_18671,N_17610,N_17023);
or U18672 (N_18672,N_17696,N_17756);
nand U18673 (N_18673,N_17421,N_17051);
xnor U18674 (N_18674,N_16897,N_17034);
nand U18675 (N_18675,N_17532,N_17956);
nor U18676 (N_18676,N_17667,N_17923);
xnor U18677 (N_18677,N_17547,N_17679);
nand U18678 (N_18678,N_16899,N_17647);
xor U18679 (N_18679,N_17043,N_17659);
xor U18680 (N_18680,N_17371,N_16800);
nor U18681 (N_18681,N_17128,N_17622);
nor U18682 (N_18682,N_16985,N_17403);
or U18683 (N_18683,N_17311,N_17630);
and U18684 (N_18684,N_16804,N_17361);
and U18685 (N_18685,N_17581,N_17717);
xor U18686 (N_18686,N_17003,N_17908);
xor U18687 (N_18687,N_17984,N_16921);
xnor U18688 (N_18688,N_17316,N_17036);
and U18689 (N_18689,N_16843,N_16921);
xnor U18690 (N_18690,N_17820,N_16954);
and U18691 (N_18691,N_17132,N_17681);
and U18692 (N_18692,N_17896,N_17072);
nor U18693 (N_18693,N_17590,N_17680);
or U18694 (N_18694,N_17268,N_17331);
nand U18695 (N_18695,N_17765,N_17915);
nand U18696 (N_18696,N_17922,N_17950);
or U18697 (N_18697,N_17127,N_17945);
nor U18698 (N_18698,N_17650,N_16921);
nand U18699 (N_18699,N_17706,N_17000);
xor U18700 (N_18700,N_17855,N_17222);
or U18701 (N_18701,N_17203,N_17385);
nand U18702 (N_18702,N_17226,N_17526);
or U18703 (N_18703,N_17209,N_17440);
or U18704 (N_18704,N_17836,N_17307);
nand U18705 (N_18705,N_17864,N_17533);
xnor U18706 (N_18706,N_17620,N_17445);
xor U18707 (N_18707,N_16807,N_17886);
nand U18708 (N_18708,N_17617,N_17439);
and U18709 (N_18709,N_17889,N_17010);
and U18710 (N_18710,N_17197,N_16930);
and U18711 (N_18711,N_17918,N_17568);
xnor U18712 (N_18712,N_17788,N_17231);
and U18713 (N_18713,N_17564,N_17881);
nand U18714 (N_18714,N_17759,N_17071);
or U18715 (N_18715,N_16921,N_17064);
or U18716 (N_18716,N_16891,N_17586);
nor U18717 (N_18717,N_16873,N_17479);
or U18718 (N_18718,N_17206,N_17378);
nor U18719 (N_18719,N_17783,N_17677);
xnor U18720 (N_18720,N_17954,N_17498);
nand U18721 (N_18721,N_17749,N_16870);
nor U18722 (N_18722,N_17456,N_17087);
xor U18723 (N_18723,N_17294,N_17785);
nor U18724 (N_18724,N_16800,N_16949);
xnor U18725 (N_18725,N_17387,N_17504);
and U18726 (N_18726,N_17011,N_17447);
nand U18727 (N_18727,N_17295,N_17580);
or U18728 (N_18728,N_17334,N_17686);
nor U18729 (N_18729,N_17633,N_17484);
and U18730 (N_18730,N_16951,N_17210);
nor U18731 (N_18731,N_17502,N_17750);
xnor U18732 (N_18732,N_17025,N_17379);
or U18733 (N_18733,N_17019,N_17415);
nor U18734 (N_18734,N_16943,N_17430);
nand U18735 (N_18735,N_17798,N_17251);
nand U18736 (N_18736,N_17530,N_17529);
xnor U18737 (N_18737,N_17435,N_17946);
nor U18738 (N_18738,N_17788,N_17492);
nor U18739 (N_18739,N_17024,N_17658);
nor U18740 (N_18740,N_17427,N_17589);
or U18741 (N_18741,N_17855,N_17184);
and U18742 (N_18742,N_16834,N_17453);
nor U18743 (N_18743,N_17856,N_17891);
nand U18744 (N_18744,N_17480,N_17029);
nand U18745 (N_18745,N_17538,N_17673);
or U18746 (N_18746,N_16805,N_17006);
xor U18747 (N_18747,N_17165,N_17642);
xnor U18748 (N_18748,N_17147,N_17788);
and U18749 (N_18749,N_16872,N_16852);
nand U18750 (N_18750,N_17069,N_17823);
xnor U18751 (N_18751,N_16876,N_17019);
xnor U18752 (N_18752,N_17747,N_17292);
nor U18753 (N_18753,N_17252,N_17670);
xor U18754 (N_18754,N_17563,N_17418);
nor U18755 (N_18755,N_17269,N_17409);
nand U18756 (N_18756,N_16976,N_17962);
and U18757 (N_18757,N_17289,N_17461);
nor U18758 (N_18758,N_17037,N_16910);
nor U18759 (N_18759,N_16824,N_17755);
and U18760 (N_18760,N_17935,N_17030);
and U18761 (N_18761,N_17955,N_16992);
nor U18762 (N_18762,N_16819,N_17619);
or U18763 (N_18763,N_17877,N_17184);
or U18764 (N_18764,N_16986,N_17162);
xor U18765 (N_18765,N_17731,N_17098);
or U18766 (N_18766,N_17047,N_17473);
nand U18767 (N_18767,N_17546,N_17952);
nand U18768 (N_18768,N_17362,N_17540);
or U18769 (N_18769,N_17231,N_17484);
xor U18770 (N_18770,N_17965,N_17861);
nor U18771 (N_18771,N_17220,N_17542);
nand U18772 (N_18772,N_17730,N_17337);
and U18773 (N_18773,N_17424,N_17802);
xnor U18774 (N_18774,N_17680,N_17352);
or U18775 (N_18775,N_17555,N_17562);
xor U18776 (N_18776,N_17538,N_17564);
xor U18777 (N_18777,N_17389,N_17582);
nor U18778 (N_18778,N_17212,N_17382);
nand U18779 (N_18779,N_17350,N_17847);
nand U18780 (N_18780,N_17235,N_17211);
nand U18781 (N_18781,N_17660,N_16803);
nand U18782 (N_18782,N_16844,N_17996);
nor U18783 (N_18783,N_16853,N_17669);
nor U18784 (N_18784,N_17687,N_17677);
nand U18785 (N_18785,N_17052,N_17942);
or U18786 (N_18786,N_17981,N_17458);
nand U18787 (N_18787,N_17374,N_17597);
nand U18788 (N_18788,N_17016,N_17306);
or U18789 (N_18789,N_17087,N_17988);
xor U18790 (N_18790,N_16868,N_17668);
nand U18791 (N_18791,N_17235,N_16967);
xnor U18792 (N_18792,N_17318,N_17292);
xor U18793 (N_18793,N_17749,N_17609);
nor U18794 (N_18794,N_17599,N_17867);
and U18795 (N_18795,N_17214,N_17199);
and U18796 (N_18796,N_17497,N_16959);
xor U18797 (N_18797,N_17486,N_17994);
xor U18798 (N_18798,N_17791,N_16988);
and U18799 (N_18799,N_16992,N_17503);
or U18800 (N_18800,N_16916,N_17808);
or U18801 (N_18801,N_17133,N_17200);
or U18802 (N_18802,N_17242,N_16911);
xnor U18803 (N_18803,N_17375,N_17273);
nor U18804 (N_18804,N_17626,N_17571);
nand U18805 (N_18805,N_16978,N_17676);
or U18806 (N_18806,N_17184,N_17288);
or U18807 (N_18807,N_17778,N_17282);
xnor U18808 (N_18808,N_16883,N_17191);
or U18809 (N_18809,N_17538,N_17748);
and U18810 (N_18810,N_17558,N_16809);
or U18811 (N_18811,N_17905,N_16886);
nor U18812 (N_18812,N_16875,N_17373);
nand U18813 (N_18813,N_17494,N_17422);
and U18814 (N_18814,N_17607,N_16843);
or U18815 (N_18815,N_17493,N_17898);
nand U18816 (N_18816,N_17320,N_17108);
xor U18817 (N_18817,N_16985,N_17422);
xor U18818 (N_18818,N_17967,N_17852);
and U18819 (N_18819,N_17231,N_17994);
nand U18820 (N_18820,N_17644,N_17842);
xnor U18821 (N_18821,N_17708,N_17719);
and U18822 (N_18822,N_17812,N_17251);
nand U18823 (N_18823,N_17354,N_17682);
nand U18824 (N_18824,N_17631,N_17990);
nor U18825 (N_18825,N_17682,N_17323);
nand U18826 (N_18826,N_17762,N_17854);
nand U18827 (N_18827,N_17673,N_17678);
and U18828 (N_18828,N_17452,N_16976);
and U18829 (N_18829,N_17321,N_17432);
and U18830 (N_18830,N_17622,N_17812);
or U18831 (N_18831,N_17510,N_17322);
or U18832 (N_18832,N_17567,N_17597);
xnor U18833 (N_18833,N_17366,N_16958);
xor U18834 (N_18834,N_17303,N_17208);
xor U18835 (N_18835,N_17689,N_17678);
xnor U18836 (N_18836,N_17496,N_16839);
and U18837 (N_18837,N_17645,N_17986);
and U18838 (N_18838,N_16802,N_17184);
nor U18839 (N_18839,N_17553,N_17856);
nand U18840 (N_18840,N_17778,N_17272);
xor U18841 (N_18841,N_16812,N_17774);
xor U18842 (N_18842,N_17221,N_17736);
or U18843 (N_18843,N_17944,N_17772);
xor U18844 (N_18844,N_16907,N_16822);
nor U18845 (N_18845,N_17979,N_17207);
xnor U18846 (N_18846,N_17491,N_16969);
nand U18847 (N_18847,N_17418,N_17736);
nor U18848 (N_18848,N_17086,N_16977);
nand U18849 (N_18849,N_17831,N_17645);
or U18850 (N_18850,N_17887,N_17300);
or U18851 (N_18851,N_17748,N_16819);
nand U18852 (N_18852,N_17421,N_16943);
nor U18853 (N_18853,N_17267,N_17576);
and U18854 (N_18854,N_17036,N_17413);
nor U18855 (N_18855,N_17445,N_17458);
and U18856 (N_18856,N_16942,N_16814);
and U18857 (N_18857,N_17750,N_17920);
or U18858 (N_18858,N_17170,N_17707);
and U18859 (N_18859,N_17264,N_16921);
xor U18860 (N_18860,N_17471,N_17848);
xnor U18861 (N_18861,N_17887,N_17705);
nor U18862 (N_18862,N_17574,N_17640);
xor U18863 (N_18863,N_17662,N_17438);
or U18864 (N_18864,N_16877,N_17860);
nor U18865 (N_18865,N_17774,N_17354);
nand U18866 (N_18866,N_17746,N_16817);
or U18867 (N_18867,N_17315,N_17982);
or U18868 (N_18868,N_17911,N_17876);
or U18869 (N_18869,N_17373,N_17624);
and U18870 (N_18870,N_17772,N_17983);
or U18871 (N_18871,N_17893,N_17697);
or U18872 (N_18872,N_16845,N_17504);
and U18873 (N_18873,N_17094,N_17920);
nand U18874 (N_18874,N_16959,N_17327);
or U18875 (N_18875,N_17990,N_17034);
nor U18876 (N_18876,N_17638,N_17655);
nand U18877 (N_18877,N_17225,N_17438);
nor U18878 (N_18878,N_17145,N_17760);
nor U18879 (N_18879,N_16897,N_16924);
xor U18880 (N_18880,N_17762,N_17298);
or U18881 (N_18881,N_17734,N_17482);
or U18882 (N_18882,N_17338,N_17386);
xor U18883 (N_18883,N_17476,N_17766);
or U18884 (N_18884,N_17289,N_16992);
or U18885 (N_18885,N_17677,N_17932);
xnor U18886 (N_18886,N_17604,N_17163);
or U18887 (N_18887,N_16971,N_17943);
and U18888 (N_18888,N_17749,N_17034);
nor U18889 (N_18889,N_17882,N_16924);
and U18890 (N_18890,N_17042,N_17292);
nor U18891 (N_18891,N_17394,N_17266);
nand U18892 (N_18892,N_17424,N_17259);
xor U18893 (N_18893,N_17676,N_17885);
xnor U18894 (N_18894,N_17241,N_17488);
and U18895 (N_18895,N_17456,N_17284);
nor U18896 (N_18896,N_17573,N_17953);
and U18897 (N_18897,N_17984,N_17647);
nor U18898 (N_18898,N_17987,N_17691);
nand U18899 (N_18899,N_17416,N_17328);
nor U18900 (N_18900,N_16945,N_17786);
and U18901 (N_18901,N_17650,N_17790);
nand U18902 (N_18902,N_17241,N_17189);
nand U18903 (N_18903,N_17847,N_17470);
or U18904 (N_18904,N_17741,N_17900);
nand U18905 (N_18905,N_17630,N_16875);
nand U18906 (N_18906,N_17653,N_17939);
nand U18907 (N_18907,N_17527,N_17980);
nor U18908 (N_18908,N_17740,N_17406);
nand U18909 (N_18909,N_17406,N_17951);
or U18910 (N_18910,N_17236,N_17969);
and U18911 (N_18911,N_17791,N_17630);
xnor U18912 (N_18912,N_17986,N_17638);
xor U18913 (N_18913,N_17918,N_17221);
and U18914 (N_18914,N_16827,N_17028);
and U18915 (N_18915,N_17783,N_17488);
and U18916 (N_18916,N_16927,N_17187);
xnor U18917 (N_18917,N_16995,N_17605);
nor U18918 (N_18918,N_17184,N_16827);
or U18919 (N_18919,N_17519,N_17372);
nor U18920 (N_18920,N_17192,N_17329);
or U18921 (N_18921,N_17687,N_17044);
nor U18922 (N_18922,N_16927,N_17757);
nor U18923 (N_18923,N_17060,N_17621);
nor U18924 (N_18924,N_17717,N_16955);
xnor U18925 (N_18925,N_17600,N_16931);
xnor U18926 (N_18926,N_17217,N_17680);
xnor U18927 (N_18927,N_17627,N_17626);
xnor U18928 (N_18928,N_17648,N_17952);
nand U18929 (N_18929,N_17475,N_16808);
nor U18930 (N_18930,N_17470,N_17559);
or U18931 (N_18931,N_17677,N_17619);
and U18932 (N_18932,N_17166,N_17242);
and U18933 (N_18933,N_17199,N_17539);
xor U18934 (N_18934,N_17122,N_17688);
xnor U18935 (N_18935,N_17868,N_17947);
nor U18936 (N_18936,N_16814,N_17397);
or U18937 (N_18937,N_16972,N_17592);
nand U18938 (N_18938,N_17760,N_17477);
or U18939 (N_18939,N_17987,N_16966);
or U18940 (N_18940,N_16999,N_17019);
nand U18941 (N_18941,N_17633,N_17692);
xnor U18942 (N_18942,N_17569,N_17419);
nor U18943 (N_18943,N_17778,N_16828);
nand U18944 (N_18944,N_17752,N_17847);
xor U18945 (N_18945,N_16887,N_16857);
nand U18946 (N_18946,N_17952,N_17488);
nor U18947 (N_18947,N_17481,N_17984);
or U18948 (N_18948,N_17733,N_16874);
nand U18949 (N_18949,N_17102,N_17738);
xor U18950 (N_18950,N_16974,N_17132);
or U18951 (N_18951,N_17053,N_17542);
nor U18952 (N_18952,N_17984,N_17360);
nor U18953 (N_18953,N_17365,N_17789);
and U18954 (N_18954,N_17984,N_17635);
and U18955 (N_18955,N_17522,N_17574);
or U18956 (N_18956,N_17801,N_17218);
nand U18957 (N_18957,N_16942,N_16838);
and U18958 (N_18958,N_17826,N_17376);
nand U18959 (N_18959,N_16881,N_16937);
nand U18960 (N_18960,N_17966,N_17206);
or U18961 (N_18961,N_16814,N_17619);
or U18962 (N_18962,N_17714,N_17858);
or U18963 (N_18963,N_17460,N_17706);
nor U18964 (N_18964,N_17934,N_17467);
or U18965 (N_18965,N_17703,N_17992);
xnor U18966 (N_18966,N_17727,N_17602);
and U18967 (N_18967,N_17735,N_17837);
xnor U18968 (N_18968,N_16883,N_17461);
nor U18969 (N_18969,N_17536,N_17468);
or U18970 (N_18970,N_17416,N_17126);
nor U18971 (N_18971,N_16811,N_16843);
xnor U18972 (N_18972,N_17094,N_17565);
nand U18973 (N_18973,N_17021,N_17253);
xnor U18974 (N_18974,N_16870,N_17002);
nand U18975 (N_18975,N_16942,N_16891);
and U18976 (N_18976,N_17368,N_17140);
nand U18977 (N_18977,N_16909,N_17682);
xnor U18978 (N_18978,N_17387,N_17958);
xnor U18979 (N_18979,N_17333,N_17889);
and U18980 (N_18980,N_16821,N_17962);
xor U18981 (N_18981,N_17278,N_17790);
and U18982 (N_18982,N_17384,N_16826);
nand U18983 (N_18983,N_17418,N_17103);
and U18984 (N_18984,N_17600,N_17820);
or U18985 (N_18985,N_17034,N_16843);
and U18986 (N_18986,N_17054,N_17966);
or U18987 (N_18987,N_17374,N_16815);
nor U18988 (N_18988,N_17126,N_17946);
xor U18989 (N_18989,N_17586,N_16836);
xor U18990 (N_18990,N_17449,N_17112);
or U18991 (N_18991,N_17228,N_17379);
and U18992 (N_18992,N_17431,N_17132);
and U18993 (N_18993,N_17403,N_17778);
xnor U18994 (N_18994,N_16943,N_16979);
nor U18995 (N_18995,N_16846,N_17162);
or U18996 (N_18996,N_17601,N_17638);
or U18997 (N_18997,N_17629,N_17333);
or U18998 (N_18998,N_17498,N_17105);
xnor U18999 (N_18999,N_17025,N_17843);
nand U19000 (N_19000,N_17379,N_17351);
and U19001 (N_19001,N_17104,N_17357);
nand U19002 (N_19002,N_16891,N_17071);
nor U19003 (N_19003,N_17534,N_17135);
nor U19004 (N_19004,N_17879,N_17283);
xnor U19005 (N_19005,N_17210,N_17765);
or U19006 (N_19006,N_16923,N_17214);
xor U19007 (N_19007,N_17864,N_17919);
nand U19008 (N_19008,N_17039,N_17276);
nor U19009 (N_19009,N_17752,N_16839);
and U19010 (N_19010,N_17543,N_17243);
xnor U19011 (N_19011,N_17529,N_17868);
xnor U19012 (N_19012,N_16800,N_16802);
and U19013 (N_19013,N_17364,N_17506);
xor U19014 (N_19014,N_17771,N_17501);
nor U19015 (N_19015,N_17140,N_17985);
nor U19016 (N_19016,N_17145,N_16998);
or U19017 (N_19017,N_17216,N_17150);
and U19018 (N_19018,N_17000,N_16910);
xnor U19019 (N_19019,N_17120,N_16938);
and U19020 (N_19020,N_17316,N_17399);
nor U19021 (N_19021,N_17682,N_16906);
nor U19022 (N_19022,N_17958,N_16921);
and U19023 (N_19023,N_17598,N_17029);
nor U19024 (N_19024,N_17969,N_17731);
nor U19025 (N_19025,N_17747,N_16812);
nand U19026 (N_19026,N_16851,N_17232);
xnor U19027 (N_19027,N_17308,N_17728);
xor U19028 (N_19028,N_17318,N_17238);
nor U19029 (N_19029,N_17700,N_17137);
xor U19030 (N_19030,N_17722,N_17044);
nand U19031 (N_19031,N_17886,N_16886);
nand U19032 (N_19032,N_17500,N_17709);
nor U19033 (N_19033,N_17487,N_17717);
or U19034 (N_19034,N_17533,N_17449);
nand U19035 (N_19035,N_17914,N_16836);
nand U19036 (N_19036,N_16998,N_16882);
and U19037 (N_19037,N_17080,N_17165);
nor U19038 (N_19038,N_17084,N_16964);
nor U19039 (N_19039,N_17800,N_16880);
or U19040 (N_19040,N_17790,N_17855);
xor U19041 (N_19041,N_17381,N_17032);
nor U19042 (N_19042,N_17065,N_17911);
nand U19043 (N_19043,N_17500,N_17970);
nor U19044 (N_19044,N_17239,N_17256);
and U19045 (N_19045,N_16817,N_17510);
nor U19046 (N_19046,N_17829,N_17360);
or U19047 (N_19047,N_17197,N_17703);
or U19048 (N_19048,N_17184,N_17591);
nand U19049 (N_19049,N_17185,N_16873);
or U19050 (N_19050,N_16959,N_17942);
nand U19051 (N_19051,N_17364,N_17017);
and U19052 (N_19052,N_17800,N_16906);
xnor U19053 (N_19053,N_17995,N_17730);
and U19054 (N_19054,N_17796,N_17026);
nor U19055 (N_19055,N_17166,N_17169);
and U19056 (N_19056,N_17308,N_17406);
and U19057 (N_19057,N_17135,N_17986);
xor U19058 (N_19058,N_17736,N_17491);
nor U19059 (N_19059,N_16816,N_17750);
or U19060 (N_19060,N_17969,N_17549);
nand U19061 (N_19061,N_17006,N_17129);
or U19062 (N_19062,N_17851,N_17464);
or U19063 (N_19063,N_17088,N_17097);
xor U19064 (N_19064,N_17792,N_17912);
nand U19065 (N_19065,N_17482,N_16919);
nand U19066 (N_19066,N_17898,N_17660);
and U19067 (N_19067,N_16887,N_17061);
and U19068 (N_19068,N_17331,N_16942);
and U19069 (N_19069,N_17485,N_16986);
nand U19070 (N_19070,N_17167,N_17704);
xor U19071 (N_19071,N_17828,N_17814);
nor U19072 (N_19072,N_17861,N_16903);
nand U19073 (N_19073,N_17566,N_17899);
nand U19074 (N_19074,N_17292,N_17235);
xnor U19075 (N_19075,N_16860,N_17348);
xor U19076 (N_19076,N_17504,N_16917);
xnor U19077 (N_19077,N_17427,N_17285);
nor U19078 (N_19078,N_17559,N_17806);
nor U19079 (N_19079,N_17463,N_16840);
or U19080 (N_19080,N_17899,N_17569);
xnor U19081 (N_19081,N_17571,N_17660);
nor U19082 (N_19082,N_17034,N_17524);
xor U19083 (N_19083,N_17587,N_16851);
or U19084 (N_19084,N_17340,N_17916);
xor U19085 (N_19085,N_16839,N_17075);
xor U19086 (N_19086,N_17480,N_17843);
nand U19087 (N_19087,N_16937,N_17378);
and U19088 (N_19088,N_17387,N_17182);
or U19089 (N_19089,N_17915,N_17424);
and U19090 (N_19090,N_17920,N_17913);
nand U19091 (N_19091,N_17332,N_17257);
or U19092 (N_19092,N_16863,N_17409);
xor U19093 (N_19093,N_17429,N_17679);
nor U19094 (N_19094,N_17192,N_16906);
and U19095 (N_19095,N_16993,N_17167);
and U19096 (N_19096,N_17889,N_17743);
nand U19097 (N_19097,N_16810,N_17820);
or U19098 (N_19098,N_17934,N_17593);
xnor U19099 (N_19099,N_16972,N_17859);
xnor U19100 (N_19100,N_17388,N_16964);
xnor U19101 (N_19101,N_16894,N_17687);
nand U19102 (N_19102,N_17725,N_17254);
or U19103 (N_19103,N_17957,N_17169);
nand U19104 (N_19104,N_17630,N_17291);
or U19105 (N_19105,N_17313,N_17674);
or U19106 (N_19106,N_17198,N_17068);
nor U19107 (N_19107,N_16936,N_16887);
nor U19108 (N_19108,N_16847,N_17442);
nor U19109 (N_19109,N_16904,N_17341);
and U19110 (N_19110,N_17399,N_17838);
nand U19111 (N_19111,N_17311,N_17038);
and U19112 (N_19112,N_17120,N_16961);
xnor U19113 (N_19113,N_16922,N_17791);
and U19114 (N_19114,N_17759,N_17929);
and U19115 (N_19115,N_17666,N_16820);
or U19116 (N_19116,N_17975,N_17948);
xnor U19117 (N_19117,N_17508,N_17194);
nor U19118 (N_19118,N_17994,N_17700);
xor U19119 (N_19119,N_17761,N_17568);
nor U19120 (N_19120,N_16930,N_17006);
and U19121 (N_19121,N_17482,N_17154);
or U19122 (N_19122,N_17303,N_17774);
nor U19123 (N_19123,N_17558,N_17975);
or U19124 (N_19124,N_17272,N_17681);
nand U19125 (N_19125,N_17378,N_17702);
and U19126 (N_19126,N_16822,N_17676);
or U19127 (N_19127,N_17294,N_17228);
nand U19128 (N_19128,N_17829,N_16800);
or U19129 (N_19129,N_17266,N_17991);
and U19130 (N_19130,N_17318,N_17277);
and U19131 (N_19131,N_17672,N_17316);
xnor U19132 (N_19132,N_16931,N_17972);
xnor U19133 (N_19133,N_17551,N_17237);
nand U19134 (N_19134,N_16829,N_17377);
nand U19135 (N_19135,N_17086,N_17976);
nor U19136 (N_19136,N_17266,N_16947);
xnor U19137 (N_19137,N_17604,N_17288);
xor U19138 (N_19138,N_17184,N_16879);
xnor U19139 (N_19139,N_17032,N_17339);
or U19140 (N_19140,N_17039,N_17512);
nand U19141 (N_19141,N_17921,N_17387);
xnor U19142 (N_19142,N_16863,N_17891);
or U19143 (N_19143,N_17375,N_17499);
nand U19144 (N_19144,N_17772,N_16972);
and U19145 (N_19145,N_17153,N_17772);
nand U19146 (N_19146,N_17732,N_17950);
xor U19147 (N_19147,N_17818,N_17205);
nand U19148 (N_19148,N_17460,N_17462);
and U19149 (N_19149,N_16976,N_17665);
and U19150 (N_19150,N_17636,N_17548);
or U19151 (N_19151,N_17152,N_17062);
or U19152 (N_19152,N_17975,N_17092);
nor U19153 (N_19153,N_17424,N_17169);
or U19154 (N_19154,N_17421,N_17162);
or U19155 (N_19155,N_17405,N_17685);
xor U19156 (N_19156,N_17598,N_17527);
nand U19157 (N_19157,N_17395,N_17129);
and U19158 (N_19158,N_17080,N_17910);
xor U19159 (N_19159,N_17294,N_16915);
nor U19160 (N_19160,N_17902,N_16890);
nand U19161 (N_19161,N_17172,N_17618);
and U19162 (N_19162,N_17135,N_17310);
and U19163 (N_19163,N_17583,N_17262);
or U19164 (N_19164,N_16981,N_17972);
nand U19165 (N_19165,N_17452,N_17777);
nor U19166 (N_19166,N_17654,N_16802);
nand U19167 (N_19167,N_17210,N_17860);
nand U19168 (N_19168,N_17427,N_17701);
and U19169 (N_19169,N_17818,N_17105);
nand U19170 (N_19170,N_17702,N_17751);
nor U19171 (N_19171,N_16901,N_17853);
and U19172 (N_19172,N_16882,N_17379);
or U19173 (N_19173,N_17408,N_17635);
nor U19174 (N_19174,N_16971,N_17664);
or U19175 (N_19175,N_17145,N_17898);
nand U19176 (N_19176,N_17644,N_17951);
nor U19177 (N_19177,N_17639,N_17185);
xnor U19178 (N_19178,N_17652,N_17536);
and U19179 (N_19179,N_17479,N_17102);
xnor U19180 (N_19180,N_17873,N_17213);
nand U19181 (N_19181,N_17110,N_17175);
nand U19182 (N_19182,N_17868,N_17767);
xnor U19183 (N_19183,N_17634,N_17200);
nand U19184 (N_19184,N_17836,N_17949);
nand U19185 (N_19185,N_16801,N_17844);
nor U19186 (N_19186,N_17769,N_17540);
or U19187 (N_19187,N_17198,N_17264);
nand U19188 (N_19188,N_17242,N_16850);
nand U19189 (N_19189,N_16824,N_17167);
nor U19190 (N_19190,N_17437,N_17692);
xnor U19191 (N_19191,N_17816,N_16884);
xor U19192 (N_19192,N_17491,N_17195);
or U19193 (N_19193,N_17951,N_17250);
xor U19194 (N_19194,N_17265,N_17622);
nand U19195 (N_19195,N_17626,N_17317);
xor U19196 (N_19196,N_17926,N_17402);
and U19197 (N_19197,N_17940,N_17296);
nor U19198 (N_19198,N_17436,N_17755);
and U19199 (N_19199,N_16993,N_16847);
nand U19200 (N_19200,N_18680,N_19046);
xnor U19201 (N_19201,N_18788,N_18704);
xor U19202 (N_19202,N_19035,N_18777);
nor U19203 (N_19203,N_18911,N_18370);
and U19204 (N_19204,N_18290,N_18278);
and U19205 (N_19205,N_19168,N_18147);
xnor U19206 (N_19206,N_18252,N_18211);
xor U19207 (N_19207,N_18347,N_18664);
nand U19208 (N_19208,N_18677,N_18433);
and U19209 (N_19209,N_18652,N_18140);
nand U19210 (N_19210,N_18700,N_18453);
nor U19211 (N_19211,N_18507,N_19186);
xor U19212 (N_19212,N_19111,N_19073);
xnor U19213 (N_19213,N_18263,N_18932);
nor U19214 (N_19214,N_18653,N_18670);
nor U19215 (N_19215,N_18172,N_18513);
xor U19216 (N_19216,N_18241,N_19127);
nand U19217 (N_19217,N_18512,N_18387);
nand U19218 (N_19218,N_19055,N_18767);
or U19219 (N_19219,N_18371,N_18941);
and U19220 (N_19220,N_18951,N_18958);
or U19221 (N_19221,N_18599,N_18683);
nor U19222 (N_19222,N_19032,N_18609);
or U19223 (N_19223,N_18378,N_18000);
or U19224 (N_19224,N_19157,N_18296);
or U19225 (N_19225,N_18090,N_19140);
or U19226 (N_19226,N_18117,N_18836);
or U19227 (N_19227,N_18108,N_18353);
or U19228 (N_19228,N_18082,N_18058);
xnor U19229 (N_19229,N_18176,N_18658);
nand U19230 (N_19230,N_18448,N_18632);
and U19231 (N_19231,N_18874,N_18754);
nand U19232 (N_19232,N_18391,N_18327);
xor U19233 (N_19233,N_18721,N_18746);
nor U19234 (N_19234,N_18210,N_18188);
nor U19235 (N_19235,N_18690,N_18167);
or U19236 (N_19236,N_19091,N_18847);
xnor U19237 (N_19237,N_18399,N_18019);
and U19238 (N_19238,N_18569,N_18612);
and U19239 (N_19239,N_18666,N_18150);
and U19240 (N_19240,N_19120,N_18462);
nand U19241 (N_19241,N_18947,N_18741);
xor U19242 (N_19242,N_18618,N_18503);
nand U19243 (N_19243,N_18185,N_18711);
nor U19244 (N_19244,N_18029,N_18887);
xor U19245 (N_19245,N_19106,N_18458);
or U19246 (N_19246,N_18998,N_18732);
xnor U19247 (N_19247,N_18723,N_18872);
nand U19248 (N_19248,N_18647,N_19143);
xor U19249 (N_19249,N_18002,N_19003);
xnor U19250 (N_19250,N_19151,N_18339);
or U19251 (N_19251,N_18235,N_18648);
nand U19252 (N_19252,N_18913,N_19085);
nor U19253 (N_19253,N_18303,N_18970);
nand U19254 (N_19254,N_18109,N_18497);
nor U19255 (N_19255,N_18114,N_18194);
or U19256 (N_19256,N_18145,N_18756);
nor U19257 (N_19257,N_18480,N_18705);
nand U19258 (N_19258,N_18243,N_18769);
nor U19259 (N_19259,N_19137,N_19083);
nand U19260 (N_19260,N_18505,N_18372);
xor U19261 (N_19261,N_18094,N_18801);
xor U19262 (N_19262,N_19029,N_19113);
nand U19263 (N_19263,N_18013,N_18990);
or U19264 (N_19264,N_18304,N_18203);
nor U19265 (N_19265,N_18464,N_19198);
nor U19266 (N_19266,N_19133,N_18280);
nand U19267 (N_19267,N_18447,N_19049);
nand U19268 (N_19268,N_18824,N_18600);
nand U19269 (N_19269,N_18725,N_18139);
xor U19270 (N_19270,N_19084,N_18411);
nor U19271 (N_19271,N_19199,N_18567);
nand U19272 (N_19272,N_18922,N_18467);
nor U19273 (N_19273,N_18423,N_18548);
and U19274 (N_19274,N_18486,N_18316);
nor U19275 (N_19275,N_18456,N_18675);
and U19276 (N_19276,N_18535,N_18573);
and U19277 (N_19277,N_18071,N_19043);
xnor U19278 (N_19278,N_19172,N_19053);
nand U19279 (N_19279,N_18460,N_18551);
and U19280 (N_19280,N_18668,N_19128);
nand U19281 (N_19281,N_18182,N_18662);
nand U19282 (N_19282,N_18734,N_19148);
nor U19283 (N_19283,N_18770,N_19004);
nor U19284 (N_19284,N_18492,N_18413);
xnor U19285 (N_19285,N_18006,N_18076);
nor U19286 (N_19286,N_18988,N_18527);
xnor U19287 (N_19287,N_19044,N_18868);
nor U19288 (N_19288,N_19033,N_18978);
and U19289 (N_19289,N_19045,N_18603);
and U19290 (N_19290,N_18628,N_19058);
nand U19291 (N_19291,N_18793,N_18157);
or U19292 (N_19292,N_19016,N_18475);
nor U19293 (N_19293,N_18436,N_18125);
xor U19294 (N_19294,N_18825,N_18067);
nand U19295 (N_19295,N_18576,N_18400);
and U19296 (N_19296,N_18786,N_18574);
nor U19297 (N_19297,N_18397,N_18291);
nand U19298 (N_19298,N_18279,N_18834);
xor U19299 (N_19299,N_18803,N_18636);
and U19300 (N_19300,N_18816,N_19006);
and U19301 (N_19301,N_18995,N_18223);
xor U19302 (N_19302,N_18098,N_18258);
nand U19303 (N_19303,N_18866,N_19162);
or U19304 (N_19304,N_18719,N_18650);
and U19305 (N_19305,N_18953,N_18017);
nand U19306 (N_19306,N_19015,N_18848);
and U19307 (N_19307,N_18283,N_18539);
or U19308 (N_19308,N_19070,N_19017);
and U19309 (N_19309,N_18643,N_18078);
and U19310 (N_19310,N_19138,N_18495);
or U19311 (N_19311,N_18102,N_18530);
xnor U19312 (N_19312,N_19178,N_18766);
xor U19313 (N_19313,N_18457,N_18350);
or U19314 (N_19314,N_18357,N_18035);
xor U19315 (N_19315,N_18107,N_18274);
nor U19316 (N_19316,N_18251,N_18165);
xnor U19317 (N_19317,N_18169,N_18917);
xor U19318 (N_19318,N_18536,N_19009);
and U19319 (N_19319,N_19052,N_18760);
nand U19320 (N_19320,N_18807,N_18861);
and U19321 (N_19321,N_18601,N_18620);
nor U19322 (N_19322,N_18038,N_18763);
xor U19323 (N_19323,N_19107,N_18928);
and U19324 (N_19324,N_18369,N_18684);
nor U19325 (N_19325,N_18465,N_18199);
or U19326 (N_19326,N_18575,N_18987);
xnor U19327 (N_19327,N_18743,N_19077);
nand U19328 (N_19328,N_19144,N_18320);
xor U19329 (N_19329,N_19161,N_18722);
or U19330 (N_19330,N_19062,N_19153);
nor U19331 (N_19331,N_18174,N_18384);
xor U19332 (N_19332,N_18914,N_19010);
nor U19333 (N_19333,N_18656,N_18819);
nor U19334 (N_19334,N_19089,N_18120);
nor U19335 (N_19335,N_18924,N_18552);
and U19336 (N_19336,N_18500,N_19019);
and U19337 (N_19337,N_19163,N_18715);
or U19338 (N_19338,N_18118,N_18748);
or U19339 (N_19339,N_19002,N_19166);
nand U19340 (N_19340,N_19050,N_18133);
or U19341 (N_19341,N_18129,N_18485);
nand U19342 (N_19342,N_18882,N_18810);
nor U19343 (N_19343,N_18192,N_18744);
xor U19344 (N_19344,N_18328,N_19109);
xor U19345 (N_19345,N_18001,N_19170);
and U19346 (N_19346,N_19125,N_18967);
nand U19347 (N_19347,N_18916,N_18317);
nor U19348 (N_19348,N_18402,N_18592);
xor U19349 (N_19349,N_18173,N_18965);
and U19350 (N_19350,N_18420,N_18589);
or U19351 (N_19351,N_18162,N_18918);
and U19352 (N_19352,N_18128,N_18968);
or U19353 (N_19353,N_19005,N_18583);
nand U19354 (N_19354,N_18640,N_19150);
nor U19355 (N_19355,N_18113,N_18307);
nor U19356 (N_19356,N_18534,N_19056);
and U19357 (N_19357,N_18005,N_18343);
xor U19358 (N_19358,N_18231,N_18940);
xnor U19359 (N_19359,N_19087,N_18451);
xor U19360 (N_19360,N_18952,N_18850);
and U19361 (N_19361,N_18047,N_18031);
and U19362 (N_19362,N_18946,N_18022);
xnor U19363 (N_19363,N_18494,N_18352);
nand U19364 (N_19364,N_18896,N_18706);
xnor U19365 (N_19365,N_18131,N_18935);
or U19366 (N_19366,N_18020,N_18586);
nor U19367 (N_19367,N_19123,N_18196);
nor U19368 (N_19368,N_18622,N_18613);
nand U19369 (N_19369,N_18178,N_18212);
or U19370 (N_19370,N_18832,N_18220);
and U19371 (N_19371,N_19187,N_18753);
nor U19372 (N_19372,N_19040,N_18966);
or U19373 (N_19373,N_19078,N_18452);
or U19374 (N_19374,N_18151,N_18837);
xor U19375 (N_19375,N_18103,N_19102);
or U19376 (N_19376,N_18830,N_18531);
nand U19377 (N_19377,N_18481,N_18389);
or U19378 (N_19378,N_18828,N_18380);
or U19379 (N_19379,N_18667,N_18214);
and U19380 (N_19380,N_18230,N_18374);
and U19381 (N_19381,N_18835,N_19051);
xnor U19382 (N_19382,N_18973,N_18406);
or U19383 (N_19383,N_18046,N_18685);
xor U19384 (N_19384,N_18607,N_18137);
xnor U19385 (N_19385,N_18703,N_18687);
nand U19386 (N_19386,N_18269,N_18617);
xnor U19387 (N_19387,N_18862,N_18471);
and U19388 (N_19388,N_18469,N_18542);
xnor U19389 (N_19389,N_18564,N_18289);
and U19390 (N_19390,N_18818,N_18854);
nor U19391 (N_19391,N_18004,N_18015);
nand U19392 (N_19392,N_18493,N_18135);
or U19393 (N_19393,N_18245,N_18487);
and U19394 (N_19394,N_18392,N_18859);
or U19395 (N_19395,N_18900,N_18356);
xor U19396 (N_19396,N_19088,N_18334);
xor U19397 (N_19397,N_18915,N_18362);
nor U19398 (N_19398,N_18877,N_18483);
and U19399 (N_19399,N_18180,N_18663);
and U19400 (N_19400,N_18043,N_18961);
and U19401 (N_19401,N_18419,N_18511);
nor U19402 (N_19402,N_18611,N_19020);
or U19403 (N_19403,N_18669,N_18478);
xor U19404 (N_19404,N_18578,N_18979);
and U19405 (N_19405,N_18297,N_19098);
xor U19406 (N_19406,N_18085,N_19007);
nand U19407 (N_19407,N_18799,N_19175);
nor U19408 (N_19408,N_18555,N_19159);
nor U19409 (N_19409,N_18365,N_18383);
or U19410 (N_19410,N_18518,N_18106);
nor U19411 (N_19411,N_18443,N_18812);
and U19412 (N_19412,N_18123,N_18954);
xnor U19413 (N_19413,N_18745,N_18591);
and U19414 (N_19414,N_18697,N_18116);
nand U19415 (N_19415,N_18974,N_18184);
and U19416 (N_19416,N_18509,N_18727);
nand U19417 (N_19417,N_19066,N_18735);
nand U19418 (N_19418,N_18689,N_18152);
or U19419 (N_19419,N_18295,N_18064);
or U19420 (N_19420,N_18260,N_18999);
and U19421 (N_19421,N_18065,N_18168);
xnor U19422 (N_19422,N_18285,N_18257);
nand U19423 (N_19423,N_18858,N_18124);
or U19424 (N_19424,N_18733,N_18962);
or U19425 (N_19425,N_18774,N_18712);
nor U19426 (N_19426,N_18694,N_18610);
nor U19427 (N_19427,N_19105,N_18189);
nand U19428 (N_19428,N_18336,N_18948);
xnor U19429 (N_19429,N_19195,N_18281);
or U19430 (N_19430,N_18883,N_18351);
nand U19431 (N_19431,N_18193,N_18331);
nor U19432 (N_19432,N_18813,N_18287);
nand U19433 (N_19433,N_19026,N_18556);
xor U19434 (N_19434,N_18254,N_18201);
xnor U19435 (N_19435,N_18190,N_19146);
xnor U19436 (N_19436,N_18313,N_19037);
nor U19437 (N_19437,N_19174,N_18377);
nor U19438 (N_19438,N_18375,N_18814);
nand U19439 (N_19439,N_18797,N_18726);
or U19440 (N_19440,N_18606,N_18981);
and U19441 (N_19441,N_19108,N_18657);
and U19442 (N_19442,N_18440,N_18943);
xor U19443 (N_19443,N_18691,N_18826);
or U19444 (N_19444,N_18454,N_18096);
nor U19445 (N_19445,N_19156,N_18839);
or U19446 (N_19446,N_18104,N_18122);
xnor U19447 (N_19447,N_19031,N_18790);
or U19448 (N_19448,N_18893,N_18891);
xor U19449 (N_19449,N_18517,N_18747);
or U19450 (N_19450,N_19099,N_18795);
and U19451 (N_19451,N_18288,N_18246);
and U19452 (N_19452,N_19145,N_18787);
or U19453 (N_19453,N_19132,N_18142);
and U19454 (N_19454,N_18267,N_19071);
xor U19455 (N_19455,N_19193,N_18649);
or U19456 (N_19456,N_18616,N_18851);
and U19457 (N_19457,N_18298,N_18055);
or U19458 (N_19458,N_18582,N_19072);
and U19459 (N_19459,N_18265,N_18838);
or U19460 (N_19460,N_18815,N_18218);
xnor U19461 (N_19461,N_18547,N_18554);
or U19462 (N_19462,N_18292,N_18804);
nand U19463 (N_19463,N_18525,N_18580);
and U19464 (N_19464,N_18084,N_18991);
nand U19465 (N_19465,N_18286,N_18401);
and U19466 (N_19466,N_19180,N_18003);
or U19467 (N_19467,N_18233,N_18864);
nor U19468 (N_19468,N_18863,N_18642);
and U19469 (N_19469,N_18061,N_18529);
and U19470 (N_19470,N_18366,N_18639);
and U19471 (N_19471,N_18829,N_18476);
xnor U19472 (N_19472,N_18659,N_18852);
xor U19473 (N_19473,N_18489,N_18321);
and U19474 (N_19474,N_18431,N_18775);
nor U19475 (N_19475,N_19131,N_18468);
and U19476 (N_19476,N_18040,N_18802);
and U19477 (N_19477,N_18594,N_18771);
and U19478 (N_19478,N_18092,N_18225);
and U19479 (N_19479,N_18596,N_18593);
nand U19480 (N_19480,N_18115,N_18718);
nand U19481 (N_19481,N_18635,N_19154);
or U19482 (N_19482,N_19068,N_18361);
or U19483 (N_19483,N_18543,N_19039);
nor U19484 (N_19484,N_18256,N_18134);
nand U19485 (N_19485,N_18992,N_18242);
or U19486 (N_19486,N_19014,N_19185);
nor U19487 (N_19487,N_18409,N_18976);
and U19488 (N_19488,N_18164,N_18259);
or U19489 (N_19489,N_18014,N_18563);
nand U19490 (N_19490,N_18198,N_18678);
nand U19491 (N_19491,N_19025,N_18363);
nand U19492 (N_19492,N_18466,N_18410);
nor U19493 (N_19493,N_18111,N_18206);
nand U19494 (N_19494,N_18950,N_18936);
or U19495 (N_19495,N_18024,N_18630);
and U19496 (N_19496,N_18121,N_19101);
and U19497 (N_19497,N_18300,N_18341);
or U19498 (N_19498,N_18626,N_18780);
and U19499 (N_19499,N_18472,N_19116);
nand U19500 (N_19500,N_19122,N_18105);
or U19501 (N_19501,N_18544,N_18876);
xnor U19502 (N_19502,N_18840,N_18739);
nand U19503 (N_19503,N_18429,N_19104);
or U19504 (N_19504,N_19184,N_18444);
and U19505 (N_19505,N_18960,N_18405);
and U19506 (N_19506,N_18025,N_18731);
xor U19507 (N_19507,N_18785,N_18737);
and U19508 (N_19508,N_18983,N_18446);
nor U19509 (N_19509,N_18337,N_18095);
nor U19510 (N_19510,N_18833,N_19008);
nor U19511 (N_19511,N_19169,N_18081);
nand U19512 (N_19512,N_19047,N_18089);
or U19513 (N_19513,N_19189,N_18742);
xor U19514 (N_19514,N_18759,N_18421);
or U19515 (N_19515,N_19096,N_18811);
xnor U19516 (N_19516,N_18101,N_18821);
xnor U19517 (N_19517,N_18736,N_19112);
and U19518 (N_19518,N_18672,N_18926);
nor U19519 (N_19519,N_18424,N_18126);
nor U19520 (N_19520,N_18349,N_18415);
nand U19521 (N_19521,N_19069,N_18056);
xnor U19522 (N_19522,N_19110,N_18942);
or U19523 (N_19523,N_18264,N_18156);
nand U19524 (N_19524,N_18282,N_19065);
nand U19525 (N_19525,N_19158,N_18927);
xor U19526 (N_19526,N_18197,N_19011);
nand U19527 (N_19527,N_18088,N_18418);
xor U19528 (N_19528,N_18323,N_18087);
xnor U19529 (N_19529,N_18515,N_18007);
or U19530 (N_19530,N_19130,N_18239);
xor U19531 (N_19531,N_18959,N_18100);
nand U19532 (N_19532,N_18021,N_18955);
nor U19533 (N_19533,N_18909,N_18855);
xnor U19534 (N_19534,N_18030,N_19124);
nor U19535 (N_19535,N_19061,N_19028);
nand U19536 (N_19536,N_18018,N_18546);
or U19537 (N_19537,N_18699,N_18902);
or U19538 (N_19538,N_19177,N_18127);
nor U19539 (N_19539,N_18545,N_18183);
and U19540 (N_19540,N_19181,N_18041);
xnor U19541 (N_19541,N_18524,N_18276);
or U19542 (N_19542,N_18571,N_18997);
and U19543 (N_19543,N_18262,N_19013);
nand U19544 (N_19544,N_18474,N_18880);
or U19545 (N_19545,N_18890,N_18161);
nand U19546 (N_19546,N_18499,N_18665);
or U19547 (N_19547,N_18310,N_18332);
or U19548 (N_19548,N_19034,N_18034);
and U19549 (N_19549,N_19194,N_18937);
or U19550 (N_19550,N_18390,N_18625);
nor U19551 (N_19551,N_18207,N_18314);
nor U19552 (N_19552,N_18093,N_18590);
or U19553 (N_19553,N_18160,N_18273);
nand U19554 (N_19554,N_18329,N_18645);
and U19555 (N_19555,N_19060,N_18956);
nor U19556 (N_19556,N_18870,N_18261);
or U19557 (N_19557,N_18050,N_18794);
or U19558 (N_19558,N_18213,N_18195);
nor U19559 (N_19559,N_18473,N_18395);
nor U19560 (N_19560,N_18408,N_18520);
nor U19561 (N_19561,N_18376,N_18271);
nand U19562 (N_19562,N_18187,N_18538);
xor U19563 (N_19563,N_18541,N_18920);
or U19564 (N_19564,N_18853,N_18439);
xor U19565 (N_19565,N_18655,N_19059);
or U19566 (N_19566,N_18779,N_18631);
and U19567 (N_19567,N_19192,N_18026);
and U19568 (N_19568,N_18910,N_18903);
and U19569 (N_19569,N_18738,N_18386);
xnor U19570 (N_19570,N_18333,N_19152);
and U19571 (N_19571,N_18191,N_18340);
or U19572 (N_19572,N_18709,N_18430);
and U19573 (N_19573,N_18776,N_18412);
and U19574 (N_19574,N_18367,N_19190);
nor U19575 (N_19575,N_18805,N_18063);
or U19576 (N_19576,N_19082,N_19095);
xor U19577 (N_19577,N_18634,N_18994);
nor U19578 (N_19578,N_18681,N_18895);
xor U19579 (N_19579,N_18843,N_18660);
or U19580 (N_19580,N_18526,N_19048);
or U19581 (N_19581,N_18345,N_18240);
nand U19582 (N_19582,N_18354,N_18484);
or U19583 (N_19583,N_18588,N_18049);
nand U19584 (N_19584,N_18938,N_18856);
nand U19585 (N_19585,N_19173,N_19054);
xor U19586 (N_19586,N_18984,N_18986);
nand U19587 (N_19587,N_18570,N_18335);
and U19588 (N_19588,N_18388,N_19147);
or U19589 (N_19589,N_18729,N_18865);
and U19590 (N_19590,N_18130,N_18579);
xnor U19591 (N_19591,N_18309,N_18584);
nor U19592 (N_19592,N_18867,N_18751);
and U19593 (N_19593,N_18514,N_18757);
nand U19594 (N_19594,N_18908,N_18166);
nand U19595 (N_19595,N_18459,N_18934);
or U19596 (N_19596,N_18077,N_18688);
and U19597 (N_19597,N_18654,N_18360);
or U19598 (N_19598,N_18572,N_18266);
nand U19599 (N_19599,N_18428,N_18977);
and U19600 (N_19600,N_18153,N_18414);
nand U19601 (N_19601,N_18841,N_18426);
xor U19602 (N_19602,N_18605,N_18091);
nand U19603 (N_19603,N_18702,N_18708);
nor U19604 (N_19604,N_18238,N_19135);
or U19605 (N_19605,N_18247,N_18502);
and U19606 (N_19606,N_18009,N_18671);
xor U19607 (N_19607,N_18846,N_18996);
or U19608 (N_19608,N_18215,N_18425);
or U19609 (N_19609,N_18396,N_19119);
and U19610 (N_19610,N_18097,N_19183);
nand U19611 (N_19611,N_18604,N_18901);
nand U19612 (N_19612,N_18698,N_19076);
nor U19613 (N_19613,N_18629,N_19182);
nand U19614 (N_19614,N_18422,N_18559);
nor U19615 (N_19615,N_18205,N_19118);
nand U19616 (N_19616,N_19036,N_18749);
and U19617 (N_19617,N_18159,N_18033);
xnor U19618 (N_19618,N_18523,N_18772);
or U19619 (N_19619,N_18522,N_18796);
and U19620 (N_19620,N_18208,N_18326);
or U19621 (N_19621,N_18470,N_19001);
or U19622 (N_19622,N_18886,N_18519);
xor U19623 (N_19623,N_18268,N_18540);
nand U19624 (N_19624,N_18608,N_18822);
and U19625 (N_19625,N_19023,N_18404);
nand U19626 (N_19626,N_18250,N_19149);
and U19627 (N_19627,N_19075,N_18714);
nor U19628 (N_19628,N_18562,N_18558);
nand U19629 (N_19629,N_18849,N_18060);
nand U19630 (N_19630,N_18442,N_18831);
or U19631 (N_19631,N_19081,N_18975);
xor U19632 (N_19632,N_18148,N_18342);
or U19633 (N_19633,N_19018,N_18227);
nand U19634 (N_19634,N_19041,N_18221);
and U19635 (N_19635,N_18045,N_19134);
or U19636 (N_19636,N_18270,N_18037);
nor U19637 (N_19637,N_18504,N_19171);
nand U19638 (N_19638,N_19165,N_18324);
or U19639 (N_19639,N_18869,N_18477);
nor U19640 (N_19640,N_18302,N_18028);
nor U19641 (N_19641,N_18209,N_18528);
xnor U19642 (N_19642,N_18305,N_18565);
xnor U19643 (N_19643,N_18012,N_18598);
nor U19644 (N_19644,N_18696,N_18817);
xor U19645 (N_19645,N_18784,N_18075);
xnor U19646 (N_19646,N_18237,N_18646);
or U19647 (N_19647,N_19139,N_18549);
or U19648 (N_19648,N_19191,N_18294);
xor U19649 (N_19649,N_18724,N_18624);
and U19650 (N_19650,N_18016,N_18044);
or U19651 (N_19651,N_18186,N_18764);
or U19652 (N_19652,N_19155,N_18144);
or U19653 (N_19653,N_18441,N_18945);
xor U19654 (N_19654,N_18881,N_18933);
and U19655 (N_19655,N_18894,N_18510);
nand U19656 (N_19656,N_18445,N_18778);
xnor U19657 (N_19657,N_18730,N_19063);
or U19658 (N_19658,N_18750,N_18236);
or U19659 (N_19659,N_18312,N_18944);
and U19660 (N_19660,N_18823,N_18762);
nand U19661 (N_19661,N_18765,N_19074);
xnor U19662 (N_19662,N_18053,N_18434);
or U19663 (N_19663,N_18720,N_18679);
xnor U19664 (N_19664,N_18330,N_18929);
xnor U19665 (N_19665,N_18619,N_18068);
nor U19666 (N_19666,N_18897,N_18532);
or U19667 (N_19667,N_18781,N_18232);
nor U19668 (N_19668,N_18407,N_18381);
and U19669 (N_19669,N_18898,N_18394);
or U19670 (N_19670,N_18170,N_18516);
and U19671 (N_19671,N_18073,N_18385);
or U19672 (N_19672,N_18806,N_19115);
or U19673 (N_19673,N_18463,N_19103);
nand U19674 (N_19674,N_18713,N_18949);
nand U19675 (N_19675,N_18686,N_18226);
nand U19676 (N_19676,N_18553,N_18857);
nand U19677 (N_19677,N_18931,N_18054);
or U19678 (N_19678,N_18338,N_18435);
and U19679 (N_19679,N_18740,N_18980);
xnor U19680 (N_19680,N_18368,N_18925);
or U19681 (N_19681,N_19022,N_19114);
and U19682 (N_19682,N_18752,N_18498);
xnor U19683 (N_19683,N_18216,N_18318);
and U19684 (N_19684,N_18234,N_18717);
nor U19685 (N_19685,N_19097,N_18845);
nor U19686 (N_19686,N_18820,N_18202);
and U19687 (N_19687,N_18889,N_18373);
nor U19688 (N_19688,N_18461,N_18141);
and U19689 (N_19689,N_18827,N_18964);
and U19690 (N_19690,N_18673,N_18971);
nand U19691 (N_19691,N_18921,N_18661);
nor U19692 (N_19692,N_18930,N_18792);
nand U19693 (N_19693,N_18358,N_18982);
and U19694 (N_19694,N_18651,N_18299);
or U19695 (N_19695,N_19021,N_18627);
and U19696 (N_19696,N_18557,N_18782);
xor U19697 (N_19697,N_18229,N_19027);
xnor U19698 (N_19698,N_18072,N_18884);
nor U19699 (N_19699,N_19079,N_18132);
nand U19700 (N_19700,N_18348,N_19086);
and U19701 (N_19701,N_19117,N_18032);
and U19702 (N_19702,N_18885,N_18253);
nor U19703 (N_19703,N_18615,N_18939);
nand U19704 (N_19704,N_18809,N_18011);
nor U19705 (N_19705,N_18993,N_18306);
or U19706 (N_19706,N_19141,N_18427);
and U19707 (N_19707,N_18985,N_18879);
and U19708 (N_19708,N_18842,N_18755);
nor U19709 (N_19709,N_19042,N_18905);
xor U19710 (N_19710,N_19090,N_18682);
xor U19711 (N_19711,N_18293,N_18692);
xor U19712 (N_19712,N_18888,N_19057);
xnor U19713 (N_19713,N_18989,N_19100);
xnor U19714 (N_19714,N_18906,N_18346);
and U19715 (N_19715,N_18158,N_18701);
or U19716 (N_19716,N_18496,N_18912);
xor U19717 (N_19717,N_18871,N_18641);
nor U19718 (N_19718,N_18875,N_18716);
nand U19719 (N_19719,N_18693,N_18069);
and U19720 (N_19720,N_18566,N_18783);
nor U19721 (N_19721,N_18907,N_18344);
nor U19722 (N_19722,N_18179,N_18163);
nor U19723 (N_19723,N_19179,N_18146);
and U19724 (N_19724,N_18758,N_18136);
nand U19725 (N_19725,N_18217,N_19196);
or U19726 (N_19726,N_18311,N_18919);
xnor U19727 (N_19727,N_18490,N_19197);
and U19728 (N_19728,N_19129,N_19000);
nor U19729 (N_19729,N_18581,N_18143);
nor U19730 (N_19730,N_18550,N_19038);
and U19731 (N_19731,N_18437,N_18432);
xor U19732 (N_19732,N_18359,N_18171);
or U19733 (N_19733,N_18074,N_18355);
or U19734 (N_19734,N_18284,N_18438);
and U19735 (N_19735,N_18789,N_18450);
nor U19736 (N_19736,N_19160,N_18325);
or U19737 (N_19737,N_18508,N_18768);
xor U19738 (N_19738,N_18248,N_18079);
nor U19739 (N_19739,N_18963,N_18644);
xor U19740 (N_19740,N_18393,N_18561);
or U19741 (N_19741,N_18479,N_18059);
nand U19742 (N_19742,N_18577,N_18923);
and U19743 (N_19743,N_18506,N_18277);
nand U19744 (N_19744,N_18791,N_18449);
nor U19745 (N_19745,N_18904,N_18695);
and U19746 (N_19746,N_18382,N_18637);
and U19747 (N_19747,N_19024,N_18023);
and U19748 (N_19748,N_18379,N_18860);
nand U19749 (N_19749,N_18597,N_18301);
or U19750 (N_19750,N_19136,N_18244);
or U19751 (N_19751,N_18800,N_18112);
nor U19752 (N_19752,N_19164,N_18537);
and U19753 (N_19753,N_19030,N_18455);
nor U19754 (N_19754,N_18482,N_18315);
xnor U19755 (N_19755,N_18204,N_18623);
and U19756 (N_19756,N_18272,N_18501);
and U19757 (N_19757,N_18728,N_18521);
nand U19758 (N_19758,N_18080,N_18674);
nand U19759 (N_19759,N_18892,N_18957);
nor U19760 (N_19760,N_18761,N_18398);
nor U19761 (N_19761,N_19093,N_18039);
nand U19762 (N_19762,N_18052,N_18222);
nand U19763 (N_19763,N_18086,N_18491);
nand U19764 (N_19764,N_18417,N_19121);
xnor U19765 (N_19765,N_18322,N_18181);
or U19766 (N_19766,N_19064,N_18585);
xnor U19767 (N_19767,N_18416,N_18036);
or U19768 (N_19768,N_19094,N_19092);
xor U19769 (N_19769,N_18488,N_19067);
xor U19770 (N_19770,N_18844,N_18051);
or U19771 (N_19771,N_18533,N_19167);
nor U19772 (N_19772,N_18676,N_18707);
xor U19773 (N_19773,N_19188,N_18621);
xor U19774 (N_19774,N_19126,N_19142);
nor U19775 (N_19775,N_18010,N_18099);
nand U19776 (N_19776,N_19012,N_18899);
nor U19777 (N_19777,N_18119,N_18008);
or U19778 (N_19778,N_18138,N_18560);
nor U19779 (N_19779,N_18249,N_18175);
nor U19780 (N_19780,N_18048,N_18972);
nand U19781 (N_19781,N_18638,N_18154);
and U19782 (N_19782,N_18319,N_18155);
or U19783 (N_19783,N_18595,N_18403);
nor U19784 (N_19784,N_18587,N_18224);
xnor U19785 (N_19785,N_19176,N_18602);
xor U19786 (N_19786,N_18878,N_18969);
xnor U19787 (N_19787,N_18070,N_18228);
xor U19788 (N_19788,N_18614,N_18568);
and U19789 (N_19789,N_18200,N_18042);
xor U19790 (N_19790,N_18710,N_18219);
or U19791 (N_19791,N_18633,N_18066);
and U19792 (N_19792,N_18057,N_18083);
nand U19793 (N_19793,N_18808,N_19080);
xnor U19794 (N_19794,N_18027,N_18177);
nor U19795 (N_19795,N_18364,N_18308);
nand U19796 (N_19796,N_18149,N_18062);
nor U19797 (N_19797,N_18275,N_18873);
or U19798 (N_19798,N_18255,N_18110);
xnor U19799 (N_19799,N_18798,N_18773);
or U19800 (N_19800,N_18672,N_18671);
and U19801 (N_19801,N_18417,N_19134);
nor U19802 (N_19802,N_18736,N_18307);
xor U19803 (N_19803,N_18978,N_18043);
nand U19804 (N_19804,N_18440,N_18699);
or U19805 (N_19805,N_18213,N_18383);
xor U19806 (N_19806,N_18099,N_19158);
nor U19807 (N_19807,N_18880,N_18428);
nand U19808 (N_19808,N_18169,N_18643);
nand U19809 (N_19809,N_18342,N_18934);
nand U19810 (N_19810,N_18303,N_18766);
nand U19811 (N_19811,N_18420,N_18113);
or U19812 (N_19812,N_18028,N_18918);
xnor U19813 (N_19813,N_18227,N_18628);
or U19814 (N_19814,N_18269,N_18636);
and U19815 (N_19815,N_18578,N_18076);
xor U19816 (N_19816,N_18924,N_18939);
or U19817 (N_19817,N_18012,N_18437);
or U19818 (N_19818,N_18374,N_18318);
or U19819 (N_19819,N_19080,N_18867);
and U19820 (N_19820,N_18615,N_19106);
xor U19821 (N_19821,N_18006,N_18658);
or U19822 (N_19822,N_18120,N_18124);
or U19823 (N_19823,N_18779,N_18394);
xnor U19824 (N_19824,N_18944,N_18562);
nand U19825 (N_19825,N_18083,N_18045);
or U19826 (N_19826,N_18434,N_19054);
nand U19827 (N_19827,N_18043,N_18183);
nand U19828 (N_19828,N_18547,N_18332);
and U19829 (N_19829,N_19005,N_19066);
or U19830 (N_19830,N_18999,N_18332);
nor U19831 (N_19831,N_18702,N_18710);
nand U19832 (N_19832,N_18896,N_18069);
nand U19833 (N_19833,N_18878,N_18100);
nand U19834 (N_19834,N_19079,N_18644);
nor U19835 (N_19835,N_18411,N_18870);
nor U19836 (N_19836,N_18410,N_18343);
nand U19837 (N_19837,N_18141,N_19022);
nand U19838 (N_19838,N_18928,N_18772);
nand U19839 (N_19839,N_18819,N_18234);
xnor U19840 (N_19840,N_18555,N_18576);
and U19841 (N_19841,N_18206,N_18456);
xnor U19842 (N_19842,N_18625,N_18600);
nand U19843 (N_19843,N_18735,N_18357);
nor U19844 (N_19844,N_18605,N_19076);
nand U19845 (N_19845,N_18161,N_18703);
xnor U19846 (N_19846,N_18301,N_18445);
xnor U19847 (N_19847,N_19114,N_19093);
nor U19848 (N_19848,N_18568,N_19187);
nand U19849 (N_19849,N_18949,N_18139);
nor U19850 (N_19850,N_18341,N_18015);
or U19851 (N_19851,N_18008,N_18865);
nor U19852 (N_19852,N_18709,N_18901);
and U19853 (N_19853,N_18352,N_18603);
nand U19854 (N_19854,N_18821,N_19175);
nor U19855 (N_19855,N_18441,N_18433);
nand U19856 (N_19856,N_18092,N_18404);
nor U19857 (N_19857,N_18332,N_18601);
nand U19858 (N_19858,N_18904,N_18323);
nand U19859 (N_19859,N_19154,N_18761);
nand U19860 (N_19860,N_19121,N_19026);
or U19861 (N_19861,N_19147,N_18672);
xor U19862 (N_19862,N_18468,N_18952);
nand U19863 (N_19863,N_18352,N_18703);
nand U19864 (N_19864,N_18664,N_18450);
xnor U19865 (N_19865,N_18327,N_19193);
nor U19866 (N_19866,N_18256,N_18348);
nor U19867 (N_19867,N_18111,N_18261);
and U19868 (N_19868,N_18841,N_18863);
nand U19869 (N_19869,N_18077,N_18170);
nor U19870 (N_19870,N_18006,N_18926);
nor U19871 (N_19871,N_18737,N_18651);
nor U19872 (N_19872,N_18854,N_18162);
nor U19873 (N_19873,N_18952,N_18168);
or U19874 (N_19874,N_18183,N_18864);
nor U19875 (N_19875,N_18044,N_18462);
nand U19876 (N_19876,N_18163,N_18666);
and U19877 (N_19877,N_19188,N_18835);
xnor U19878 (N_19878,N_18337,N_19145);
and U19879 (N_19879,N_18813,N_18367);
nand U19880 (N_19880,N_18271,N_18819);
nor U19881 (N_19881,N_18066,N_18459);
nor U19882 (N_19882,N_18577,N_18910);
xor U19883 (N_19883,N_18733,N_18885);
nand U19884 (N_19884,N_18019,N_18966);
nor U19885 (N_19885,N_18036,N_18738);
or U19886 (N_19886,N_18920,N_18336);
and U19887 (N_19887,N_18124,N_18956);
or U19888 (N_19888,N_18976,N_18347);
nor U19889 (N_19889,N_18204,N_18978);
nand U19890 (N_19890,N_18990,N_18075);
nor U19891 (N_19891,N_18797,N_18651);
nor U19892 (N_19892,N_18512,N_18426);
nand U19893 (N_19893,N_18216,N_18495);
and U19894 (N_19894,N_18278,N_18866);
or U19895 (N_19895,N_18226,N_18546);
nand U19896 (N_19896,N_18469,N_18071);
xnor U19897 (N_19897,N_18304,N_18666);
xnor U19898 (N_19898,N_18852,N_18898);
and U19899 (N_19899,N_18115,N_18608);
or U19900 (N_19900,N_18433,N_18710);
or U19901 (N_19901,N_18671,N_18347);
or U19902 (N_19902,N_18855,N_18535);
or U19903 (N_19903,N_18172,N_18921);
xor U19904 (N_19904,N_18612,N_18496);
nor U19905 (N_19905,N_18539,N_18846);
xor U19906 (N_19906,N_18111,N_18805);
nand U19907 (N_19907,N_18048,N_19013);
nand U19908 (N_19908,N_18991,N_18364);
and U19909 (N_19909,N_18345,N_18720);
xnor U19910 (N_19910,N_18713,N_18519);
and U19911 (N_19911,N_18182,N_18375);
and U19912 (N_19912,N_18343,N_19195);
xnor U19913 (N_19913,N_18056,N_18044);
or U19914 (N_19914,N_18570,N_18128);
nor U19915 (N_19915,N_18338,N_18450);
and U19916 (N_19916,N_18634,N_18023);
and U19917 (N_19917,N_18602,N_19084);
xnor U19918 (N_19918,N_18636,N_18799);
and U19919 (N_19919,N_18043,N_18794);
nor U19920 (N_19920,N_19164,N_18620);
or U19921 (N_19921,N_19143,N_18315);
nor U19922 (N_19922,N_19100,N_18315);
or U19923 (N_19923,N_18959,N_18127);
nor U19924 (N_19924,N_18791,N_18235);
nor U19925 (N_19925,N_18886,N_18305);
xnor U19926 (N_19926,N_18156,N_19072);
and U19927 (N_19927,N_19046,N_18031);
or U19928 (N_19928,N_18074,N_19179);
nor U19929 (N_19929,N_18565,N_18498);
xor U19930 (N_19930,N_19126,N_19149);
nand U19931 (N_19931,N_19057,N_18321);
nand U19932 (N_19932,N_18981,N_18526);
nand U19933 (N_19933,N_18766,N_18809);
nand U19934 (N_19934,N_18480,N_18476);
xnor U19935 (N_19935,N_19154,N_18047);
nor U19936 (N_19936,N_19056,N_18469);
nor U19937 (N_19937,N_18431,N_18457);
or U19938 (N_19938,N_18743,N_18347);
or U19939 (N_19939,N_18749,N_18454);
xor U19940 (N_19940,N_18254,N_18478);
nand U19941 (N_19941,N_18659,N_18813);
or U19942 (N_19942,N_18514,N_18120);
and U19943 (N_19943,N_18236,N_18088);
xor U19944 (N_19944,N_18720,N_18009);
nand U19945 (N_19945,N_18228,N_18063);
and U19946 (N_19946,N_18218,N_18948);
nor U19947 (N_19947,N_18447,N_19013);
and U19948 (N_19948,N_18640,N_19178);
nand U19949 (N_19949,N_18320,N_18896);
and U19950 (N_19950,N_18509,N_18743);
xnor U19951 (N_19951,N_19108,N_18940);
nand U19952 (N_19952,N_18000,N_18489);
or U19953 (N_19953,N_18851,N_18221);
nor U19954 (N_19954,N_19107,N_18435);
nor U19955 (N_19955,N_18712,N_18661);
nand U19956 (N_19956,N_18733,N_18246);
or U19957 (N_19957,N_18226,N_18244);
and U19958 (N_19958,N_18625,N_18837);
or U19959 (N_19959,N_18864,N_18846);
and U19960 (N_19960,N_18754,N_18517);
or U19961 (N_19961,N_19059,N_18455);
or U19962 (N_19962,N_18912,N_18526);
nand U19963 (N_19963,N_18782,N_18602);
and U19964 (N_19964,N_18786,N_18228);
and U19965 (N_19965,N_18510,N_19198);
and U19966 (N_19966,N_19173,N_19063);
xor U19967 (N_19967,N_18021,N_18532);
and U19968 (N_19968,N_18364,N_18460);
nand U19969 (N_19969,N_18654,N_19044);
or U19970 (N_19970,N_18080,N_18227);
or U19971 (N_19971,N_18323,N_19080);
and U19972 (N_19972,N_18890,N_18932);
nand U19973 (N_19973,N_19117,N_18452);
nand U19974 (N_19974,N_19045,N_18403);
or U19975 (N_19975,N_18504,N_18765);
or U19976 (N_19976,N_18982,N_18795);
nand U19977 (N_19977,N_18173,N_18078);
and U19978 (N_19978,N_19014,N_19181);
nor U19979 (N_19979,N_18644,N_18975);
and U19980 (N_19980,N_18819,N_18706);
nand U19981 (N_19981,N_18991,N_18715);
nand U19982 (N_19982,N_18499,N_18414);
xor U19983 (N_19983,N_18389,N_18121);
or U19984 (N_19984,N_18203,N_18699);
and U19985 (N_19985,N_18820,N_19077);
nor U19986 (N_19986,N_18864,N_18925);
nor U19987 (N_19987,N_18406,N_19169);
nand U19988 (N_19988,N_18797,N_18996);
or U19989 (N_19989,N_19190,N_18920);
and U19990 (N_19990,N_18370,N_19027);
or U19991 (N_19991,N_18954,N_18164);
nor U19992 (N_19992,N_18088,N_18573);
and U19993 (N_19993,N_18831,N_18542);
nand U19994 (N_19994,N_18680,N_18155);
or U19995 (N_19995,N_18924,N_18475);
or U19996 (N_19996,N_18662,N_18941);
xor U19997 (N_19997,N_18944,N_18619);
nor U19998 (N_19998,N_18055,N_19159);
nand U19999 (N_19999,N_18258,N_18145);
or U20000 (N_20000,N_18314,N_19077);
nor U20001 (N_20001,N_19054,N_18250);
nor U20002 (N_20002,N_19183,N_18322);
and U20003 (N_20003,N_18009,N_19192);
nor U20004 (N_20004,N_18076,N_19043);
or U20005 (N_20005,N_18175,N_18453);
or U20006 (N_20006,N_18077,N_18194);
xor U20007 (N_20007,N_18550,N_18636);
or U20008 (N_20008,N_18288,N_18194);
nand U20009 (N_20009,N_18411,N_18127);
xnor U20010 (N_20010,N_18958,N_18727);
nor U20011 (N_20011,N_18224,N_18647);
or U20012 (N_20012,N_19157,N_18348);
nand U20013 (N_20013,N_18151,N_18924);
nor U20014 (N_20014,N_18346,N_18410);
nor U20015 (N_20015,N_19013,N_18660);
and U20016 (N_20016,N_18425,N_18832);
or U20017 (N_20017,N_19166,N_19072);
and U20018 (N_20018,N_18078,N_18147);
nor U20019 (N_20019,N_18736,N_18538);
nand U20020 (N_20020,N_18352,N_18885);
and U20021 (N_20021,N_19103,N_18919);
nand U20022 (N_20022,N_18301,N_18217);
and U20023 (N_20023,N_18070,N_18317);
and U20024 (N_20024,N_18669,N_18427);
nand U20025 (N_20025,N_18984,N_18415);
nor U20026 (N_20026,N_19080,N_18604);
nand U20027 (N_20027,N_18171,N_18585);
nor U20028 (N_20028,N_18497,N_19194);
nand U20029 (N_20029,N_18703,N_18615);
xnor U20030 (N_20030,N_18114,N_18751);
and U20031 (N_20031,N_18912,N_18557);
or U20032 (N_20032,N_18912,N_18295);
nor U20033 (N_20033,N_18877,N_18459);
xnor U20034 (N_20034,N_18756,N_18063);
or U20035 (N_20035,N_19040,N_18339);
nand U20036 (N_20036,N_19173,N_18433);
or U20037 (N_20037,N_18515,N_18237);
and U20038 (N_20038,N_18522,N_18590);
or U20039 (N_20039,N_18590,N_18509);
nor U20040 (N_20040,N_18675,N_18966);
or U20041 (N_20041,N_18472,N_18890);
or U20042 (N_20042,N_18010,N_18446);
or U20043 (N_20043,N_18043,N_18370);
and U20044 (N_20044,N_18389,N_18302);
nand U20045 (N_20045,N_19129,N_18892);
and U20046 (N_20046,N_18677,N_19105);
nand U20047 (N_20047,N_18286,N_18671);
or U20048 (N_20048,N_19192,N_18662);
or U20049 (N_20049,N_18750,N_18310);
and U20050 (N_20050,N_18907,N_18878);
nand U20051 (N_20051,N_19079,N_19086);
nand U20052 (N_20052,N_18449,N_18956);
nand U20053 (N_20053,N_18015,N_18545);
xor U20054 (N_20054,N_18635,N_18874);
nor U20055 (N_20055,N_19126,N_18760);
and U20056 (N_20056,N_18230,N_18470);
or U20057 (N_20057,N_18609,N_18121);
and U20058 (N_20058,N_18955,N_18484);
nor U20059 (N_20059,N_18132,N_18159);
xor U20060 (N_20060,N_18867,N_18499);
xor U20061 (N_20061,N_18485,N_18775);
nor U20062 (N_20062,N_19118,N_19039);
nor U20063 (N_20063,N_18887,N_19054);
and U20064 (N_20064,N_18171,N_18200);
and U20065 (N_20065,N_18642,N_18831);
nand U20066 (N_20066,N_18603,N_18828);
nand U20067 (N_20067,N_18558,N_18214);
nor U20068 (N_20068,N_18184,N_18333);
nand U20069 (N_20069,N_19118,N_18767);
and U20070 (N_20070,N_18989,N_18563);
or U20071 (N_20071,N_18423,N_18220);
xor U20072 (N_20072,N_18034,N_18202);
or U20073 (N_20073,N_18793,N_19043);
nand U20074 (N_20074,N_18175,N_19183);
xnor U20075 (N_20075,N_18447,N_18546);
nor U20076 (N_20076,N_18916,N_19167);
nor U20077 (N_20077,N_18213,N_18580);
or U20078 (N_20078,N_18104,N_18271);
and U20079 (N_20079,N_18016,N_18606);
or U20080 (N_20080,N_19089,N_19109);
and U20081 (N_20081,N_18963,N_18533);
xnor U20082 (N_20082,N_19012,N_19050);
xor U20083 (N_20083,N_18064,N_19188);
and U20084 (N_20084,N_18971,N_18739);
and U20085 (N_20085,N_18986,N_18514);
or U20086 (N_20086,N_18940,N_18475);
or U20087 (N_20087,N_19100,N_18131);
nor U20088 (N_20088,N_18943,N_18584);
nor U20089 (N_20089,N_18433,N_18956);
xnor U20090 (N_20090,N_18715,N_18888);
or U20091 (N_20091,N_18813,N_18555);
nor U20092 (N_20092,N_18130,N_18307);
xor U20093 (N_20093,N_18563,N_19007);
nor U20094 (N_20094,N_18860,N_18063);
xor U20095 (N_20095,N_18818,N_18612);
nor U20096 (N_20096,N_18551,N_18319);
nor U20097 (N_20097,N_18695,N_18053);
nand U20098 (N_20098,N_18708,N_18536);
or U20099 (N_20099,N_18882,N_18073);
xnor U20100 (N_20100,N_19120,N_18099);
nor U20101 (N_20101,N_18561,N_18493);
xor U20102 (N_20102,N_19032,N_18465);
nor U20103 (N_20103,N_18162,N_18668);
nor U20104 (N_20104,N_18469,N_18595);
or U20105 (N_20105,N_18191,N_18980);
nand U20106 (N_20106,N_18570,N_18351);
xnor U20107 (N_20107,N_18348,N_18405);
xor U20108 (N_20108,N_18196,N_18580);
nor U20109 (N_20109,N_19146,N_18403);
or U20110 (N_20110,N_19023,N_18187);
and U20111 (N_20111,N_18394,N_18964);
xnor U20112 (N_20112,N_18483,N_18722);
nand U20113 (N_20113,N_18995,N_18954);
nor U20114 (N_20114,N_18515,N_18620);
nand U20115 (N_20115,N_18160,N_18535);
xnor U20116 (N_20116,N_18068,N_18418);
nor U20117 (N_20117,N_18730,N_18458);
and U20118 (N_20118,N_18739,N_18287);
nor U20119 (N_20119,N_18732,N_18996);
or U20120 (N_20120,N_19002,N_18771);
nand U20121 (N_20121,N_19081,N_18869);
nand U20122 (N_20122,N_18516,N_18045);
nor U20123 (N_20123,N_18987,N_18195);
nand U20124 (N_20124,N_19047,N_18342);
and U20125 (N_20125,N_18153,N_18304);
and U20126 (N_20126,N_18632,N_18909);
nor U20127 (N_20127,N_18498,N_19121);
nand U20128 (N_20128,N_18645,N_18790);
and U20129 (N_20129,N_18940,N_18830);
nor U20130 (N_20130,N_18020,N_18738);
nand U20131 (N_20131,N_18410,N_18629);
and U20132 (N_20132,N_18648,N_18018);
and U20133 (N_20133,N_18691,N_18093);
nand U20134 (N_20134,N_18300,N_18611);
nand U20135 (N_20135,N_18771,N_18724);
nor U20136 (N_20136,N_18756,N_18559);
and U20137 (N_20137,N_18949,N_18975);
nand U20138 (N_20138,N_19199,N_18122);
nand U20139 (N_20139,N_18578,N_18855);
nand U20140 (N_20140,N_19133,N_18345);
and U20141 (N_20141,N_18011,N_18479);
xnor U20142 (N_20142,N_18125,N_18855);
xor U20143 (N_20143,N_18730,N_18878);
and U20144 (N_20144,N_18606,N_18494);
xnor U20145 (N_20145,N_18300,N_18409);
and U20146 (N_20146,N_18038,N_19121);
or U20147 (N_20147,N_18667,N_18891);
nor U20148 (N_20148,N_18237,N_18828);
xnor U20149 (N_20149,N_18017,N_18685);
xnor U20150 (N_20150,N_18182,N_18458);
or U20151 (N_20151,N_18122,N_18011);
and U20152 (N_20152,N_18153,N_18188);
nor U20153 (N_20153,N_18782,N_18544);
and U20154 (N_20154,N_18935,N_18446);
nand U20155 (N_20155,N_18469,N_18847);
nor U20156 (N_20156,N_19113,N_18295);
and U20157 (N_20157,N_18220,N_18148);
and U20158 (N_20158,N_18412,N_18818);
or U20159 (N_20159,N_18922,N_18195);
or U20160 (N_20160,N_19070,N_18775);
or U20161 (N_20161,N_18384,N_18371);
nor U20162 (N_20162,N_19138,N_18572);
nor U20163 (N_20163,N_18465,N_18445);
nand U20164 (N_20164,N_18789,N_18173);
and U20165 (N_20165,N_18673,N_18427);
xnor U20166 (N_20166,N_19005,N_18277);
nand U20167 (N_20167,N_18565,N_18362);
nor U20168 (N_20168,N_19095,N_18186);
nand U20169 (N_20169,N_18143,N_18914);
nand U20170 (N_20170,N_18784,N_18114);
or U20171 (N_20171,N_18392,N_18571);
or U20172 (N_20172,N_19060,N_19079);
nand U20173 (N_20173,N_18308,N_18413);
nand U20174 (N_20174,N_18892,N_18148);
xnor U20175 (N_20175,N_18993,N_18547);
nand U20176 (N_20176,N_18274,N_18949);
and U20177 (N_20177,N_18126,N_18210);
nand U20178 (N_20178,N_19197,N_18237);
nand U20179 (N_20179,N_18025,N_19027);
and U20180 (N_20180,N_18130,N_18630);
or U20181 (N_20181,N_18837,N_19062);
xnor U20182 (N_20182,N_18905,N_19024);
and U20183 (N_20183,N_18788,N_18580);
and U20184 (N_20184,N_18562,N_18612);
and U20185 (N_20185,N_18815,N_18262);
and U20186 (N_20186,N_18885,N_18947);
nand U20187 (N_20187,N_19063,N_18618);
or U20188 (N_20188,N_18132,N_18365);
or U20189 (N_20189,N_18268,N_18880);
or U20190 (N_20190,N_19041,N_18274);
or U20191 (N_20191,N_18699,N_18139);
nand U20192 (N_20192,N_19010,N_18525);
nor U20193 (N_20193,N_18276,N_19179);
xnor U20194 (N_20194,N_18566,N_19008);
and U20195 (N_20195,N_18659,N_18049);
nand U20196 (N_20196,N_18020,N_18449);
xor U20197 (N_20197,N_18500,N_18819);
nand U20198 (N_20198,N_18238,N_18331);
nor U20199 (N_20199,N_18926,N_18159);
and U20200 (N_20200,N_18935,N_18327);
xor U20201 (N_20201,N_18648,N_18033);
and U20202 (N_20202,N_18638,N_19179);
or U20203 (N_20203,N_18003,N_18968);
and U20204 (N_20204,N_18401,N_18843);
xnor U20205 (N_20205,N_18224,N_18982);
xnor U20206 (N_20206,N_18284,N_18809);
and U20207 (N_20207,N_18960,N_19123);
nand U20208 (N_20208,N_18857,N_18995);
nor U20209 (N_20209,N_18601,N_18530);
nor U20210 (N_20210,N_18957,N_18970);
or U20211 (N_20211,N_19090,N_18831);
xnor U20212 (N_20212,N_18131,N_18196);
xnor U20213 (N_20213,N_18816,N_18112);
or U20214 (N_20214,N_18554,N_18943);
or U20215 (N_20215,N_19045,N_19173);
or U20216 (N_20216,N_18586,N_18814);
nor U20217 (N_20217,N_18784,N_18504);
nor U20218 (N_20218,N_18919,N_18300);
nor U20219 (N_20219,N_18815,N_18799);
xor U20220 (N_20220,N_18166,N_18981);
xnor U20221 (N_20221,N_19199,N_18712);
nand U20222 (N_20222,N_18388,N_19048);
and U20223 (N_20223,N_19098,N_18148);
nor U20224 (N_20224,N_18998,N_18703);
nor U20225 (N_20225,N_18922,N_18030);
and U20226 (N_20226,N_18291,N_18507);
nand U20227 (N_20227,N_18392,N_18835);
nor U20228 (N_20228,N_18400,N_18667);
or U20229 (N_20229,N_18758,N_18009);
or U20230 (N_20230,N_18964,N_18085);
xnor U20231 (N_20231,N_18659,N_18416);
or U20232 (N_20232,N_19007,N_18365);
nor U20233 (N_20233,N_18618,N_18062);
nor U20234 (N_20234,N_18610,N_18128);
nand U20235 (N_20235,N_19050,N_18966);
nor U20236 (N_20236,N_18360,N_18587);
nor U20237 (N_20237,N_18069,N_18940);
and U20238 (N_20238,N_19045,N_18437);
xnor U20239 (N_20239,N_18709,N_18036);
or U20240 (N_20240,N_18352,N_18697);
nand U20241 (N_20241,N_19058,N_18233);
or U20242 (N_20242,N_18715,N_18712);
nand U20243 (N_20243,N_18706,N_18561);
or U20244 (N_20244,N_18263,N_18348);
and U20245 (N_20245,N_18563,N_18833);
or U20246 (N_20246,N_18348,N_18479);
nand U20247 (N_20247,N_18230,N_18024);
or U20248 (N_20248,N_18960,N_18764);
and U20249 (N_20249,N_19052,N_18223);
xnor U20250 (N_20250,N_18143,N_18150);
nor U20251 (N_20251,N_18581,N_18975);
nand U20252 (N_20252,N_18414,N_18481);
nor U20253 (N_20253,N_18157,N_18251);
xnor U20254 (N_20254,N_18701,N_19033);
xnor U20255 (N_20255,N_18801,N_18783);
nand U20256 (N_20256,N_19020,N_18020);
nand U20257 (N_20257,N_18575,N_18287);
nor U20258 (N_20258,N_18652,N_19069);
and U20259 (N_20259,N_18262,N_18909);
or U20260 (N_20260,N_19083,N_18130);
nor U20261 (N_20261,N_18998,N_18027);
and U20262 (N_20262,N_18118,N_18756);
xnor U20263 (N_20263,N_18810,N_18878);
or U20264 (N_20264,N_18324,N_19183);
or U20265 (N_20265,N_18132,N_18012);
nor U20266 (N_20266,N_18651,N_18378);
nand U20267 (N_20267,N_18514,N_18546);
or U20268 (N_20268,N_19101,N_18030);
or U20269 (N_20269,N_18420,N_18934);
xor U20270 (N_20270,N_18432,N_18656);
xor U20271 (N_20271,N_19017,N_19192);
nor U20272 (N_20272,N_19159,N_18116);
nand U20273 (N_20273,N_18492,N_18054);
xor U20274 (N_20274,N_19172,N_18847);
nor U20275 (N_20275,N_19199,N_18285);
nand U20276 (N_20276,N_18814,N_18427);
xnor U20277 (N_20277,N_19050,N_18521);
nor U20278 (N_20278,N_18109,N_19165);
nor U20279 (N_20279,N_18763,N_18064);
xnor U20280 (N_20280,N_18069,N_18417);
nand U20281 (N_20281,N_18495,N_18575);
and U20282 (N_20282,N_18853,N_18307);
or U20283 (N_20283,N_18668,N_18313);
or U20284 (N_20284,N_18019,N_18598);
nand U20285 (N_20285,N_18928,N_18669);
xnor U20286 (N_20286,N_18880,N_18832);
xor U20287 (N_20287,N_18086,N_19134);
nand U20288 (N_20288,N_19142,N_18253);
nor U20289 (N_20289,N_18041,N_18378);
and U20290 (N_20290,N_18452,N_18629);
and U20291 (N_20291,N_18234,N_18405);
nand U20292 (N_20292,N_18060,N_18272);
or U20293 (N_20293,N_18621,N_18704);
nor U20294 (N_20294,N_18296,N_18078);
and U20295 (N_20295,N_18410,N_19198);
and U20296 (N_20296,N_18859,N_18095);
nor U20297 (N_20297,N_18988,N_18472);
nor U20298 (N_20298,N_18666,N_19184);
nand U20299 (N_20299,N_18682,N_19185);
xor U20300 (N_20300,N_18008,N_18881);
nor U20301 (N_20301,N_18531,N_18220);
or U20302 (N_20302,N_18144,N_18848);
nand U20303 (N_20303,N_18898,N_18331);
nand U20304 (N_20304,N_18917,N_18096);
and U20305 (N_20305,N_18900,N_18552);
and U20306 (N_20306,N_19030,N_18790);
xnor U20307 (N_20307,N_19133,N_19037);
and U20308 (N_20308,N_18236,N_18425);
nor U20309 (N_20309,N_18794,N_19123);
xnor U20310 (N_20310,N_18181,N_18875);
xnor U20311 (N_20311,N_19067,N_18699);
xnor U20312 (N_20312,N_18647,N_18163);
xor U20313 (N_20313,N_18549,N_18381);
nor U20314 (N_20314,N_18246,N_18046);
xor U20315 (N_20315,N_18565,N_18031);
nor U20316 (N_20316,N_18980,N_19079);
nand U20317 (N_20317,N_18291,N_18846);
and U20318 (N_20318,N_18771,N_18782);
nor U20319 (N_20319,N_18451,N_18775);
nand U20320 (N_20320,N_18138,N_18531);
and U20321 (N_20321,N_18418,N_18023);
nand U20322 (N_20322,N_18149,N_18309);
nor U20323 (N_20323,N_18510,N_18423);
or U20324 (N_20324,N_18863,N_19174);
nand U20325 (N_20325,N_18515,N_18375);
nand U20326 (N_20326,N_18977,N_19179);
nand U20327 (N_20327,N_18573,N_18004);
nand U20328 (N_20328,N_18327,N_18376);
and U20329 (N_20329,N_18848,N_18333);
nand U20330 (N_20330,N_18903,N_18024);
xnor U20331 (N_20331,N_18161,N_18414);
or U20332 (N_20332,N_18246,N_18426);
xor U20333 (N_20333,N_18248,N_18351);
nor U20334 (N_20334,N_18003,N_18177);
xnor U20335 (N_20335,N_18255,N_18964);
nor U20336 (N_20336,N_18173,N_18418);
nand U20337 (N_20337,N_18801,N_18960);
and U20338 (N_20338,N_19037,N_18782);
and U20339 (N_20339,N_18969,N_18205);
and U20340 (N_20340,N_18534,N_18868);
or U20341 (N_20341,N_18858,N_18806);
and U20342 (N_20342,N_18134,N_18211);
nor U20343 (N_20343,N_18939,N_18060);
or U20344 (N_20344,N_18458,N_18040);
or U20345 (N_20345,N_18978,N_18414);
xor U20346 (N_20346,N_19144,N_19190);
xor U20347 (N_20347,N_18268,N_18710);
nor U20348 (N_20348,N_18645,N_19165);
or U20349 (N_20349,N_19176,N_18039);
nor U20350 (N_20350,N_18042,N_18898);
nand U20351 (N_20351,N_18317,N_18398);
and U20352 (N_20352,N_18818,N_18083);
xnor U20353 (N_20353,N_19143,N_18463);
nand U20354 (N_20354,N_18035,N_18257);
and U20355 (N_20355,N_18169,N_18130);
xnor U20356 (N_20356,N_18827,N_18663);
xor U20357 (N_20357,N_18289,N_18949);
xor U20358 (N_20358,N_18886,N_18217);
nand U20359 (N_20359,N_18086,N_18027);
nand U20360 (N_20360,N_19085,N_18575);
nor U20361 (N_20361,N_18557,N_19177);
or U20362 (N_20362,N_18827,N_18244);
or U20363 (N_20363,N_18954,N_18111);
or U20364 (N_20364,N_18254,N_18119);
xor U20365 (N_20365,N_18463,N_18897);
nand U20366 (N_20366,N_18325,N_18271);
or U20367 (N_20367,N_18519,N_19078);
xnor U20368 (N_20368,N_18052,N_18929);
or U20369 (N_20369,N_18130,N_18375);
nor U20370 (N_20370,N_18588,N_18799);
nor U20371 (N_20371,N_18252,N_19185);
and U20372 (N_20372,N_18782,N_18829);
nand U20373 (N_20373,N_19132,N_18583);
nand U20374 (N_20374,N_18540,N_18104);
and U20375 (N_20375,N_18569,N_18443);
and U20376 (N_20376,N_18752,N_18901);
nor U20377 (N_20377,N_18741,N_18813);
or U20378 (N_20378,N_19169,N_18924);
or U20379 (N_20379,N_18733,N_18799);
nor U20380 (N_20380,N_19092,N_19057);
or U20381 (N_20381,N_18763,N_18879);
nor U20382 (N_20382,N_18348,N_18636);
nor U20383 (N_20383,N_18991,N_18010);
or U20384 (N_20384,N_18532,N_19066);
xnor U20385 (N_20385,N_18481,N_18141);
or U20386 (N_20386,N_19088,N_18810);
or U20387 (N_20387,N_18464,N_18841);
nor U20388 (N_20388,N_19139,N_18419);
or U20389 (N_20389,N_18456,N_18919);
or U20390 (N_20390,N_18411,N_19055);
nor U20391 (N_20391,N_18968,N_18786);
or U20392 (N_20392,N_18418,N_19067);
nand U20393 (N_20393,N_18041,N_19148);
xor U20394 (N_20394,N_18878,N_19175);
nor U20395 (N_20395,N_18975,N_18917);
and U20396 (N_20396,N_18522,N_18808);
and U20397 (N_20397,N_18530,N_18638);
and U20398 (N_20398,N_18452,N_18943);
or U20399 (N_20399,N_18339,N_19152);
xor U20400 (N_20400,N_19991,N_19333);
nor U20401 (N_20401,N_20006,N_19579);
and U20402 (N_20402,N_19852,N_20280);
nand U20403 (N_20403,N_19557,N_19335);
nor U20404 (N_20404,N_19986,N_19535);
or U20405 (N_20405,N_19483,N_19355);
or U20406 (N_20406,N_19366,N_20003);
nor U20407 (N_20407,N_19570,N_19866);
nor U20408 (N_20408,N_19624,N_19241);
or U20409 (N_20409,N_19423,N_19350);
or U20410 (N_20410,N_19467,N_19916);
and U20411 (N_20411,N_20007,N_19735);
nand U20412 (N_20412,N_19386,N_20374);
nand U20413 (N_20413,N_19950,N_19396);
and U20414 (N_20414,N_19864,N_20246);
or U20415 (N_20415,N_20061,N_19356);
nand U20416 (N_20416,N_19717,N_19723);
and U20417 (N_20417,N_20148,N_19446);
nor U20418 (N_20418,N_20213,N_20321);
and U20419 (N_20419,N_19304,N_20153);
and U20420 (N_20420,N_20342,N_19381);
nand U20421 (N_20421,N_19913,N_20134);
nor U20422 (N_20422,N_20305,N_19251);
nor U20423 (N_20423,N_19865,N_19987);
or U20424 (N_20424,N_19258,N_19501);
and U20425 (N_20425,N_20326,N_19341);
xor U20426 (N_20426,N_19897,N_19325);
xnor U20427 (N_20427,N_19281,N_19202);
xor U20428 (N_20428,N_19395,N_20051);
or U20429 (N_20429,N_19364,N_20230);
nand U20430 (N_20430,N_19972,N_20236);
or U20431 (N_20431,N_19232,N_19351);
and U20432 (N_20432,N_19317,N_20347);
xnor U20433 (N_20433,N_19431,N_19323);
xor U20434 (N_20434,N_19985,N_19294);
or U20435 (N_20435,N_20244,N_19316);
nor U20436 (N_20436,N_19550,N_19222);
or U20437 (N_20437,N_20385,N_19538);
and U20438 (N_20438,N_20351,N_19681);
xor U20439 (N_20439,N_20093,N_20319);
or U20440 (N_20440,N_19766,N_19715);
nand U20441 (N_20441,N_19754,N_19418);
nor U20442 (N_20442,N_20025,N_19272);
nor U20443 (N_20443,N_19552,N_19684);
or U20444 (N_20444,N_19266,N_19697);
xnor U20445 (N_20445,N_19937,N_20005);
nor U20446 (N_20446,N_20376,N_19758);
nand U20447 (N_20447,N_20212,N_19569);
nor U20448 (N_20448,N_19466,N_19971);
xor U20449 (N_20449,N_19597,N_19828);
xor U20450 (N_20450,N_19360,N_19435);
and U20451 (N_20451,N_19876,N_20111);
nor U20452 (N_20452,N_19737,N_20096);
or U20453 (N_20453,N_19405,N_19474);
and U20454 (N_20454,N_19330,N_19773);
nand U20455 (N_20455,N_19906,N_19776);
nand U20456 (N_20456,N_19635,N_19973);
and U20457 (N_20457,N_19449,N_19771);
nor U20458 (N_20458,N_20090,N_20106);
nand U20459 (N_20459,N_20195,N_19795);
and U20460 (N_20460,N_20306,N_19512);
or U20461 (N_20461,N_20085,N_19677);
and U20462 (N_20462,N_19461,N_19701);
nand U20463 (N_20463,N_19373,N_20249);
and U20464 (N_20464,N_20227,N_19228);
xor U20465 (N_20465,N_19755,N_19902);
xor U20466 (N_20466,N_19277,N_19205);
xor U20467 (N_20467,N_20270,N_20181);
or U20468 (N_20468,N_20395,N_19947);
and U20469 (N_20469,N_20063,N_20026);
nand U20470 (N_20470,N_19582,N_19941);
xnor U20471 (N_20471,N_19200,N_20384);
nand U20472 (N_20472,N_19939,N_19777);
or U20473 (N_20473,N_19887,N_19514);
or U20474 (N_20474,N_19695,N_20002);
or U20475 (N_20475,N_19548,N_20140);
or U20476 (N_20476,N_19475,N_19756);
nor U20477 (N_20477,N_19860,N_19470);
xor U20478 (N_20478,N_20170,N_20372);
and U20479 (N_20479,N_20393,N_19940);
and U20480 (N_20480,N_19440,N_20233);
nor U20481 (N_20481,N_19920,N_19314);
nand U20482 (N_20482,N_19797,N_20194);
and U20483 (N_20483,N_20108,N_19734);
or U20484 (N_20484,N_19690,N_20293);
xnor U20485 (N_20485,N_19741,N_19370);
nand U20486 (N_20486,N_19551,N_19286);
or U20487 (N_20487,N_20127,N_19278);
nand U20488 (N_20488,N_19555,N_19320);
or U20489 (N_20489,N_19539,N_19398);
or U20490 (N_20490,N_19517,N_19713);
xnor U20491 (N_20491,N_19375,N_19781);
and U20492 (N_20492,N_20067,N_19763);
or U20493 (N_20493,N_19420,N_19826);
nor U20494 (N_20494,N_19660,N_19993);
xor U20495 (N_20495,N_19340,N_20359);
xor U20496 (N_20496,N_19667,N_19457);
and U20497 (N_20497,N_20253,N_19237);
or U20498 (N_20498,N_20069,N_20091);
nor U20499 (N_20499,N_20028,N_20240);
and U20500 (N_20500,N_19979,N_19785);
nor U20501 (N_20501,N_20114,N_20373);
xnor U20502 (N_20502,N_19290,N_19665);
nand U20503 (N_20503,N_20183,N_20049);
nor U20504 (N_20504,N_19306,N_19401);
nor U20505 (N_20505,N_19556,N_19641);
nand U20506 (N_20506,N_19430,N_19425);
and U20507 (N_20507,N_19962,N_19309);
and U20508 (N_20508,N_19465,N_19632);
or U20509 (N_20509,N_19458,N_20116);
or U20510 (N_20510,N_19663,N_19308);
and U20511 (N_20511,N_19793,N_20320);
or U20512 (N_20512,N_20179,N_19943);
nand U20513 (N_20513,N_19583,N_19289);
xor U20514 (N_20514,N_19918,N_19217);
nor U20515 (N_20515,N_20316,N_19898);
nand U20516 (N_20516,N_20142,N_20291);
xnor U20517 (N_20517,N_19293,N_20295);
and U20518 (N_20518,N_19447,N_19969);
nor U20519 (N_20519,N_20394,N_19409);
nand U20520 (N_20520,N_19592,N_20272);
nand U20521 (N_20521,N_19923,N_19774);
nand U20522 (N_20522,N_19662,N_19786);
xnor U20523 (N_20523,N_19203,N_19807);
xnor U20524 (N_20524,N_20038,N_19218);
or U20525 (N_20525,N_19675,N_19576);
xnor U20526 (N_20526,N_19213,N_19863);
nand U20527 (N_20527,N_20135,N_20109);
nand U20528 (N_20528,N_20363,N_19903);
xnor U20529 (N_20529,N_19368,N_20024);
and U20530 (N_20530,N_20251,N_19329);
nand U20531 (N_20531,N_20260,N_19254);
and U20532 (N_20532,N_20149,N_19464);
xnor U20533 (N_20533,N_19647,N_19818);
or U20534 (N_20534,N_19910,N_20035);
nand U20535 (N_20535,N_19589,N_19646);
xnor U20536 (N_20536,N_19770,N_19305);
nand U20537 (N_20537,N_19451,N_20014);
nand U20538 (N_20538,N_19869,N_20123);
nand U20539 (N_20539,N_20274,N_19421);
nor U20540 (N_20540,N_19578,N_19437);
or U20541 (N_20541,N_20083,N_19426);
and U20542 (N_20542,N_19242,N_19714);
xnor U20543 (N_20543,N_19740,N_19788);
or U20544 (N_20544,N_19498,N_19678);
or U20545 (N_20545,N_19264,N_19959);
or U20546 (N_20546,N_19958,N_19400);
xnor U20547 (N_20547,N_20268,N_20141);
nand U20548 (N_20548,N_19670,N_19843);
nand U20549 (N_20549,N_19736,N_19315);
or U20550 (N_20550,N_19605,N_20339);
or U20551 (N_20551,N_19768,N_19416);
nor U20552 (N_20552,N_19683,N_19616);
and U20553 (N_20553,N_20180,N_19702);
and U20554 (N_20554,N_19919,N_19566);
nand U20555 (N_20555,N_19933,N_19964);
xnor U20556 (N_20556,N_20278,N_20378);
or U20557 (N_20557,N_19673,N_19637);
nor U20558 (N_20558,N_19821,N_19659);
or U20559 (N_20559,N_20380,N_19925);
and U20560 (N_20560,N_20329,N_19493);
nand U20561 (N_20561,N_19927,N_19250);
and U20562 (N_20562,N_19263,N_19230);
xnor U20563 (N_20563,N_19995,N_20330);
and U20564 (N_20564,N_19604,N_19994);
nand U20565 (N_20565,N_19444,N_20344);
nand U20566 (N_20566,N_19561,N_20082);
nor U20567 (N_20567,N_19298,N_20059);
and U20568 (N_20568,N_19879,N_20033);
nor U20569 (N_20569,N_19705,N_19388);
or U20570 (N_20570,N_19233,N_19626);
nand U20571 (N_20571,N_19509,N_20232);
and U20572 (N_20572,N_20346,N_19982);
nor U20573 (N_20573,N_19328,N_20084);
nand U20574 (N_20574,N_19438,N_19562);
nor U20575 (N_20575,N_19434,N_20036);
xnor U20576 (N_20576,N_19645,N_19724);
or U20577 (N_20577,N_19759,N_19584);
nand U20578 (N_20578,N_19393,N_19600);
and U20579 (N_20579,N_20095,N_20275);
and U20580 (N_20580,N_19299,N_20110);
or U20581 (N_20581,N_19274,N_19489);
nand U20582 (N_20582,N_19238,N_20099);
and U20583 (N_20583,N_19862,N_20340);
and U20584 (N_20584,N_19729,N_19427);
xnor U20585 (N_20585,N_19255,N_19883);
or U20586 (N_20586,N_19669,N_19997);
and U20587 (N_20587,N_19471,N_19956);
nand U20588 (N_20588,N_19836,N_19837);
and U20589 (N_20589,N_20118,N_20216);
or U20590 (N_20590,N_20048,N_19819);
or U20591 (N_20591,N_19376,N_19392);
nor U20592 (N_20592,N_19804,N_19436);
or U20593 (N_20593,N_19407,N_19347);
nand U20594 (N_20594,N_19270,N_19841);
or U20595 (N_20595,N_19224,N_19379);
nor U20596 (N_20596,N_20365,N_19303);
nand U20597 (N_20597,N_19780,N_20105);
nand U20598 (N_20598,N_19634,N_19811);
and U20599 (N_20599,N_19901,N_19382);
and U20600 (N_20600,N_19215,N_20369);
nor U20601 (N_20601,N_19404,N_19282);
nand U20602 (N_20602,N_19743,N_19301);
and U20603 (N_20603,N_19784,N_19412);
and U20604 (N_20604,N_20196,N_20054);
and U20605 (N_20605,N_20277,N_20345);
xnor U20606 (N_20606,N_19428,N_20327);
and U20607 (N_20607,N_19322,N_19899);
or U20608 (N_20608,N_20081,N_19686);
nand U20609 (N_20609,N_19861,N_19545);
nand U20610 (N_20610,N_20097,N_20064);
and U20611 (N_20611,N_20331,N_19806);
nand U20612 (N_20612,N_19511,N_20279);
and U20613 (N_20613,N_19761,N_20021);
or U20614 (N_20614,N_20050,N_19651);
or U20615 (N_20615,N_19935,N_20386);
xor U20616 (N_20616,N_19846,N_20042);
nor U20617 (N_20617,N_20087,N_20168);
or U20618 (N_20618,N_19374,N_19480);
and U20619 (N_20619,N_20205,N_19324);
nand U20620 (N_20620,N_19508,N_19515);
and U20621 (N_20621,N_19952,N_19267);
nand U20622 (N_20622,N_19287,N_20158);
and U20623 (N_20623,N_19623,N_19990);
xor U20624 (N_20624,N_19648,N_20052);
and U20625 (N_20625,N_19629,N_19853);
nor U20626 (N_20626,N_19738,N_20368);
and U20627 (N_20627,N_19731,N_19767);
xnor U20628 (N_20628,N_19297,N_19621);
nor U20629 (N_20629,N_19881,N_19989);
nand U20630 (N_20630,N_20258,N_20334);
or U20631 (N_20631,N_20350,N_20112);
nor U20632 (N_20632,N_19833,N_19674);
nor U20633 (N_20633,N_20335,N_19915);
nand U20634 (N_20634,N_19248,N_20103);
nand U20635 (N_20635,N_20217,N_19394);
xnor U20636 (N_20636,N_19571,N_20147);
and U20637 (N_20637,N_19479,N_19572);
nand U20638 (N_20638,N_19809,N_20030);
xor U20639 (N_20639,N_20391,N_19808);
or U20640 (N_20640,N_20190,N_19478);
or U20641 (N_20641,N_20264,N_20381);
and U20642 (N_20642,N_19856,N_20294);
or U20643 (N_20643,N_19868,N_20269);
or U20644 (N_20644,N_20377,N_20337);
xor U20645 (N_20645,N_19300,N_19219);
nand U20646 (N_20646,N_19454,N_19500);
xnor U20647 (N_20647,N_19588,N_20176);
nand U20648 (N_20648,N_20143,N_20150);
nor U20649 (N_20649,N_19851,N_19574);
or U20650 (N_20650,N_20125,N_20089);
nor U20651 (N_20651,N_19829,N_19399);
nor U20652 (N_20652,N_20178,N_19975);
xor U20653 (N_20653,N_19456,N_20129);
nand U20654 (N_20654,N_19492,N_19234);
and U20655 (N_20655,N_19658,N_20145);
xor U20656 (N_20656,N_20088,N_19854);
and U20657 (N_20657,N_19358,N_20322);
xnor U20658 (N_20658,N_19611,N_20262);
nor U20659 (N_20659,N_19365,N_20100);
or U20660 (N_20660,N_19628,N_19513);
nand U20661 (N_20661,N_19614,N_19619);
xor U20662 (N_20662,N_19960,N_20016);
or U20663 (N_20663,N_19452,N_20201);
xor U20664 (N_20664,N_19602,N_19594);
xnor U20665 (N_20665,N_19657,N_19321);
and U20666 (N_20666,N_19253,N_19271);
or U20667 (N_20667,N_19585,N_19847);
and U20668 (N_20668,N_19649,N_19859);
xor U20669 (N_20669,N_19671,N_19835);
xor U20670 (N_20670,N_20017,N_19565);
or U20671 (N_20671,N_19380,N_19812);
xnor U20672 (N_20672,N_19803,N_19344);
xnor U20673 (N_20673,N_19802,N_19815);
nand U20674 (N_20674,N_19432,N_19936);
xnor U20675 (N_20675,N_20189,N_20164);
xnor U20676 (N_20676,N_19229,N_20389);
nand U20677 (N_20677,N_19769,N_20323);
xnor U20678 (N_20678,N_19867,N_20120);
or U20679 (N_20679,N_20199,N_19482);
nand U20680 (N_20680,N_19591,N_19728);
or U20681 (N_20681,N_19424,N_20130);
xor U20682 (N_20682,N_19595,N_19313);
xnor U20683 (N_20683,N_20161,N_20229);
and U20684 (N_20684,N_20068,N_19599);
nand U20685 (N_20685,N_20259,N_20200);
nor U20686 (N_20686,N_19790,N_20318);
and U20687 (N_20687,N_19699,N_19696);
nor U20688 (N_20688,N_19210,N_19996);
or U20689 (N_20689,N_20098,N_19485);
xor U20690 (N_20690,N_19832,N_19617);
and U20691 (N_20691,N_20072,N_19433);
or U20692 (N_20692,N_19656,N_19844);
xnor U20693 (N_20693,N_20008,N_20165);
xnor U20694 (N_20694,N_19966,N_20160);
or U20695 (N_20695,N_19268,N_20273);
xnor U20696 (N_20696,N_19885,N_20167);
xor U20697 (N_20697,N_19782,N_20202);
and U20698 (N_20698,N_19486,N_19760);
nor U20699 (N_20699,N_20324,N_19503);
nand U20700 (N_20700,N_19718,N_19842);
nand U20701 (N_20701,N_20392,N_19801);
or U20702 (N_20702,N_20012,N_19544);
nand U20703 (N_20703,N_20211,N_19295);
xor U20704 (N_20704,N_19291,N_19462);
xor U20705 (N_20705,N_19654,N_19820);
nor U20706 (N_20706,N_20267,N_19612);
and U20707 (N_20707,N_19516,N_19810);
xnor U20708 (N_20708,N_19922,N_19911);
nand U20709 (N_20709,N_20358,N_19463);
nand U20710 (N_20710,N_20029,N_19402);
nand U20711 (N_20711,N_20107,N_19792);
nand U20712 (N_20712,N_19223,N_19257);
nand U20713 (N_20713,N_19273,N_19694);
nor U20714 (N_20714,N_19746,N_20155);
xor U20715 (N_20715,N_19698,N_20283);
nand U20716 (N_20716,N_20124,N_19757);
or U20717 (N_20717,N_19615,N_20182);
and U20718 (N_20718,N_19904,N_19926);
xnor U20719 (N_20719,N_19775,N_19858);
or U20720 (N_20720,N_20299,N_19676);
nand U20721 (N_20721,N_19722,N_20309);
nand U20722 (N_20722,N_20056,N_20075);
nand U20723 (N_20723,N_20060,N_20173);
nor U20724 (N_20724,N_19794,N_19469);
or U20725 (N_20725,N_19288,N_19563);
and U20726 (N_20726,N_19442,N_20250);
nor U20727 (N_20727,N_19888,N_19598);
or U20728 (N_20728,N_19530,N_20325);
xnor U20729 (N_20729,N_19840,N_20362);
nor U20730 (N_20730,N_19607,N_19417);
xnor U20731 (N_20731,N_19895,N_19639);
nand U20732 (N_20732,N_19453,N_20276);
or U20733 (N_20733,N_20198,N_19216);
and U20734 (N_20734,N_19824,N_19664);
or U20735 (N_20735,N_20288,N_19929);
xor U20736 (N_20736,N_20137,N_20242);
xor U20737 (N_20737,N_19725,N_20210);
nor U20738 (N_20738,N_20315,N_20333);
xor U20739 (N_20739,N_19256,N_19526);
nand U20740 (N_20740,N_19988,N_19871);
or U20741 (N_20741,N_19744,N_20353);
xnor U20742 (N_20742,N_20261,N_20296);
xor U20743 (N_20743,N_19640,N_19601);
nand U20744 (N_20744,N_19227,N_19596);
and U20745 (N_20745,N_20071,N_19630);
and U20746 (N_20746,N_20151,N_19719);
xnor U20747 (N_20747,N_19798,N_19965);
nor U20748 (N_20748,N_19870,N_20045);
nand U20749 (N_20749,N_19525,N_19727);
xnor U20750 (N_20750,N_20207,N_19226);
nor U20751 (N_20751,N_19873,N_20304);
or U20752 (N_20752,N_20080,N_20128);
nor U20753 (N_20753,N_19528,N_19560);
xnor U20754 (N_20754,N_19814,N_19712);
xnor U20755 (N_20755,N_19799,N_20214);
or U20756 (N_20756,N_19613,N_20265);
nor U20757 (N_20757,N_20254,N_20101);
or U20758 (N_20758,N_20222,N_19261);
nand U20759 (N_20759,N_19312,N_19575);
xor U20760 (N_20760,N_19473,N_19796);
and U20761 (N_20761,N_20215,N_19685);
nor U20762 (N_20762,N_19504,N_19917);
or U20763 (N_20763,N_19331,N_19208);
nand U20764 (N_20764,N_19772,N_19706);
nor U20765 (N_20765,N_19779,N_19558);
xnor U20766 (N_20766,N_19886,N_20022);
or U20767 (N_20767,N_19448,N_19337);
xnor U20768 (N_20768,N_20018,N_20188);
xnor U20769 (N_20769,N_19580,N_19800);
nand U20770 (N_20770,N_20184,N_19816);
nand U20771 (N_20771,N_20397,N_19638);
xnor U20772 (N_20772,N_20197,N_20286);
xnor U20773 (N_20773,N_19502,N_20307);
and U20774 (N_20774,N_20037,N_19679);
nand U20775 (N_20775,N_19534,N_19764);
or U20776 (N_20776,N_19371,N_19912);
or U20777 (N_20777,N_19524,N_19472);
nor U20778 (N_20778,N_19240,N_19276);
or U20779 (N_20779,N_19932,N_20354);
nor U20780 (N_20780,N_19220,N_19532);
xnor U20781 (N_20781,N_20154,N_19978);
nand U20782 (N_20782,N_19951,N_19488);
xor U20783 (N_20783,N_19443,N_20078);
and U20784 (N_20784,N_19823,N_19327);
nand U20785 (N_20785,N_19924,N_19239);
xnor U20786 (N_20786,N_19593,N_20065);
nand U20787 (N_20787,N_20144,N_19541);
nor U20788 (N_20788,N_19839,N_19419);
and U20789 (N_20789,N_19791,N_20185);
nand U20790 (N_20790,N_20079,N_20241);
and U20791 (N_20791,N_20379,N_19296);
nor U20792 (N_20792,N_20218,N_20203);
nand U20793 (N_20793,N_19813,N_19201);
xor U20794 (N_20794,N_19415,N_20302);
and U20795 (N_20795,N_19577,N_20290);
and U20796 (N_20796,N_19682,N_20138);
xor U20797 (N_20797,N_20177,N_19930);
or U20798 (N_20798,N_20073,N_20255);
nand U20799 (N_20799,N_20383,N_20220);
and U20800 (N_20800,N_20292,N_19477);
nor U20801 (N_20801,N_20131,N_20387);
xor U20802 (N_20802,N_19450,N_19225);
and U20803 (N_20803,N_19362,N_20297);
and U20804 (N_20804,N_19211,N_19494);
nor U20805 (N_20805,N_20226,N_19609);
xnor U20806 (N_20806,N_19908,N_19302);
and U20807 (N_20807,N_19311,N_20219);
and U20808 (N_20808,N_20187,N_19636);
or U20809 (N_20809,N_19716,N_19822);
nor U20810 (N_20810,N_20360,N_20338);
and U20811 (N_20811,N_20169,N_19389);
xnor U20812 (N_20812,N_20370,N_19586);
or U20813 (N_20813,N_20062,N_20015);
and U20814 (N_20814,N_20361,N_20238);
nor U20815 (N_20815,N_19893,N_19455);
or U20816 (N_20816,N_20192,N_19652);
nor U20817 (N_20817,N_20044,N_19610);
xor U20818 (N_20818,N_19490,N_19590);
nor U20819 (N_20819,N_19949,N_20396);
or U20820 (N_20820,N_20136,N_19247);
xnor U20821 (N_20821,N_19285,N_19506);
xor U20822 (N_20822,N_19880,N_20077);
nor U20823 (N_20823,N_19280,N_19339);
nand U20824 (N_20824,N_20284,N_20133);
nand U20825 (N_20825,N_19606,N_19397);
and U20826 (N_20826,N_19954,N_20332);
xor U20827 (N_20827,N_20235,N_20175);
or U20828 (N_20828,N_19390,N_20032);
and U20829 (N_20829,N_19338,N_19359);
nand U20830 (N_20830,N_19945,N_19882);
nor U20831 (N_20831,N_20171,N_20303);
nand U20832 (N_20832,N_19762,N_19896);
nand U20833 (N_20833,N_20245,N_19739);
or U20834 (N_20834,N_20122,N_20209);
or U20835 (N_20835,N_19789,N_20282);
or U20836 (N_20836,N_19907,N_20191);
nor U20837 (N_20837,N_19948,N_19387);
or U20838 (N_20838,N_20019,N_19672);
and U20839 (N_20839,N_20011,N_19441);
or U20840 (N_20840,N_19934,N_19711);
xnor U20841 (N_20841,N_19353,N_19522);
nand U20842 (N_20842,N_20057,N_19292);
or U20843 (N_20843,N_20186,N_20031);
xor U20844 (N_20844,N_19567,N_19332);
nor U20845 (N_20845,N_20020,N_19495);
nand U20846 (N_20846,N_19805,N_20058);
xor U20847 (N_20847,N_19889,N_19547);
and U20848 (N_20848,N_20266,N_20094);
nand U20849 (N_20849,N_19825,N_19529);
or U20850 (N_20850,N_20314,N_19284);
and U20851 (N_20851,N_20162,N_19413);
nand U20852 (N_20852,N_19827,N_19977);
xor U20853 (N_20853,N_19349,N_19783);
and U20854 (N_20854,N_19909,N_19279);
and U20855 (N_20855,N_19720,N_19408);
or U20856 (N_20856,N_20356,N_19850);
xnor U20857 (N_20857,N_19765,N_20070);
nand U20858 (N_20858,N_19981,N_19403);
or U20859 (N_20859,N_19236,N_20121);
xnor U20860 (N_20860,N_19752,N_20119);
and U20861 (N_20861,N_19944,N_19894);
xor U20862 (N_20862,N_19406,N_19377);
nor U20863 (N_20863,N_19384,N_20364);
xor U20864 (N_20864,N_19687,N_19980);
and U20865 (N_20865,N_19603,N_19206);
nor U20866 (N_20866,N_19688,N_20300);
nor U20867 (N_20867,N_19265,N_19905);
nor U20868 (N_20868,N_20074,N_19207);
xor U20869 (N_20869,N_19942,N_19703);
nor U20870 (N_20870,N_20113,N_19875);
or U20871 (N_20871,N_19733,N_20352);
and U20872 (N_20872,N_20086,N_20009);
nor U20873 (N_20873,N_20013,N_19491);
nor U20874 (N_20874,N_19378,N_20102);
xor U20875 (N_20875,N_20263,N_20301);
and U20876 (N_20876,N_20204,N_19747);
nand U20877 (N_20877,N_19385,N_19559);
xnor U20878 (N_20878,N_20132,N_19573);
nand U20879 (N_20879,N_20231,N_19543);
or U20880 (N_20880,N_20001,N_20023);
nand U20881 (N_20881,N_19643,N_19410);
xor U20882 (N_20882,N_19546,N_19505);
nor U20883 (N_20883,N_19343,N_19983);
xnor U20884 (N_20884,N_19348,N_19357);
nor U20885 (N_20885,N_20041,N_20066);
and U20886 (N_20886,N_20206,N_19642);
nand U20887 (N_20887,N_20055,N_19721);
nand U20888 (N_20888,N_19751,N_20043);
and U20889 (N_20889,N_20243,N_19468);
nor U20890 (N_20890,N_19890,N_19817);
xor U20891 (N_20891,N_19914,N_19487);
nor U20892 (N_20892,N_20355,N_19831);
and U20893 (N_20893,N_19521,N_20298);
nor U20894 (N_20894,N_19633,N_20341);
nor U20895 (N_20895,N_20234,N_20285);
and U20896 (N_20896,N_19587,N_19476);
nand U20897 (N_20897,N_19892,N_20256);
xor U20898 (N_20898,N_20046,N_19984);
xor U20899 (N_20899,N_19748,N_20371);
nand U20900 (N_20900,N_20163,N_19655);
nand U20901 (N_20901,N_19554,N_19957);
nor U20902 (N_20902,N_19622,N_19872);
nor U20903 (N_20903,N_20117,N_19260);
or U20904 (N_20904,N_19310,N_20399);
or U20905 (N_20905,N_19921,N_19520);
nor U20906 (N_20906,N_19531,N_19422);
and U20907 (N_20907,N_20126,N_19245);
or U20908 (N_20908,N_20349,N_19283);
xor U20909 (N_20909,N_19787,N_19383);
xnor U20910 (N_20910,N_19668,N_20348);
or U20911 (N_20911,N_20115,N_19484);
or U20912 (N_20912,N_20193,N_19745);
and U20913 (N_20913,N_19523,N_20310);
nor U20914 (N_20914,N_19710,N_19691);
and U20915 (N_20915,N_19369,N_20040);
and U20916 (N_20916,N_19644,N_19708);
nor U20917 (N_20917,N_19212,N_20004);
nor U20918 (N_20918,N_19753,N_19650);
nor U20919 (N_20919,N_20336,N_20271);
and U20920 (N_20920,N_19429,N_20159);
nand U20921 (N_20921,N_19661,N_19334);
xor U20922 (N_20922,N_19537,N_19931);
xnor U20923 (N_20923,N_19269,N_20252);
or U20924 (N_20924,N_19346,N_19411);
and U20925 (N_20925,N_20146,N_19834);
or U20926 (N_20926,N_19845,N_20237);
xor U20927 (N_20927,N_19518,N_20313);
and U20928 (N_20928,N_19946,N_19700);
or U20929 (N_20929,N_19726,N_19608);
or U20930 (N_20930,N_19848,N_19354);
nand U20931 (N_20931,N_19884,N_19414);
nor U20932 (N_20932,N_19221,N_19459);
nor U20933 (N_20933,N_19900,N_20156);
nand U20934 (N_20934,N_19857,N_19627);
nand U20935 (N_20935,N_19542,N_19707);
or U20936 (N_20936,N_19246,N_19838);
nor U20937 (N_20937,N_19625,N_20000);
nor U20938 (N_20938,N_19999,N_19704);
nor U20939 (N_20939,N_19439,N_19938);
nand U20940 (N_20940,N_20257,N_19961);
nor U20941 (N_20941,N_19666,N_19874);
or U20942 (N_20942,N_19970,N_20104);
xnor U20943 (N_20943,N_20367,N_19549);
xor U20944 (N_20944,N_19877,N_19568);
nand U20945 (N_20945,N_20308,N_19214);
nand U20946 (N_20946,N_20228,N_19732);
or U20947 (N_20947,N_19445,N_19345);
and U20948 (N_20948,N_20390,N_19262);
xnor U20949 (N_20949,N_19361,N_19778);
nor U20950 (N_20950,N_19564,N_19849);
or U20951 (N_20951,N_20223,N_19878);
nand U20952 (N_20952,N_19618,N_20092);
nor U20953 (N_20953,N_19510,N_19527);
xnor U20954 (N_20954,N_20311,N_19620);
nand U20955 (N_20955,N_20027,N_19249);
nand U20956 (N_20956,N_19497,N_20166);
nor U20957 (N_20957,N_19204,N_19967);
and U20958 (N_20958,N_19460,N_20289);
nand U20959 (N_20959,N_19750,N_19749);
nor U20960 (N_20960,N_20312,N_20076);
or U20961 (N_20961,N_19507,N_20248);
nor U20962 (N_20962,N_20034,N_20398);
and U20963 (N_20963,N_19209,N_19689);
nand U20964 (N_20964,N_20328,N_19692);
xor U20965 (N_20965,N_19243,N_19275);
or U20966 (N_20966,N_19992,N_19553);
or U20967 (N_20967,N_19955,N_20172);
and U20968 (N_20968,N_20366,N_20053);
nand U20969 (N_20969,N_19391,N_19631);
nand U20970 (N_20970,N_19367,N_20208);
and U20971 (N_20971,N_20157,N_19519);
nor U20972 (N_20972,N_20247,N_19693);
and U20973 (N_20973,N_20039,N_20225);
nor U20974 (N_20974,N_19342,N_20343);
and U20975 (N_20975,N_19953,N_19974);
xor U20976 (N_20976,N_19653,N_19742);
xor U20977 (N_20977,N_19231,N_19326);
xor U20978 (N_20978,N_19318,N_20357);
and U20979 (N_20979,N_19976,N_19891);
xnor U20980 (N_20980,N_19963,N_19307);
nand U20981 (N_20981,N_19968,N_19533);
and U20982 (N_20982,N_19252,N_19830);
or U20983 (N_20983,N_20224,N_20174);
nor U20984 (N_20984,N_19481,N_19499);
nand U20985 (N_20985,N_19855,N_19352);
nand U20986 (N_20986,N_19998,N_19536);
nor U20987 (N_20987,N_20010,N_19680);
xnor U20988 (N_20988,N_20388,N_19540);
and U20989 (N_20989,N_20047,N_19581);
and U20990 (N_20990,N_19319,N_19730);
and U20991 (N_20991,N_20221,N_20281);
and U20992 (N_20992,N_20382,N_19709);
xnor U20993 (N_20993,N_19244,N_20152);
nand U20994 (N_20994,N_20375,N_20287);
nor U20995 (N_20995,N_19235,N_20239);
nor U20996 (N_20996,N_20139,N_19363);
nor U20997 (N_20997,N_19928,N_19372);
xor U20998 (N_20998,N_20317,N_19259);
nor U20999 (N_20999,N_19496,N_19336);
nand U21000 (N_21000,N_19705,N_19843);
nor U21001 (N_21001,N_19450,N_19803);
xnor U21002 (N_21002,N_19224,N_20127);
or U21003 (N_21003,N_20068,N_20326);
and U21004 (N_21004,N_19507,N_19413);
or U21005 (N_21005,N_20386,N_19300);
xor U21006 (N_21006,N_20173,N_19950);
xor U21007 (N_21007,N_20178,N_20117);
or U21008 (N_21008,N_19493,N_19312);
nor U21009 (N_21009,N_19735,N_20322);
nor U21010 (N_21010,N_19420,N_19288);
nand U21011 (N_21011,N_19284,N_19645);
xor U21012 (N_21012,N_20163,N_19996);
xor U21013 (N_21013,N_19900,N_19559);
or U21014 (N_21014,N_19423,N_19470);
nand U21015 (N_21015,N_19758,N_20083);
nand U21016 (N_21016,N_20027,N_20170);
nand U21017 (N_21017,N_19912,N_19546);
xnor U21018 (N_21018,N_19607,N_20071);
nand U21019 (N_21019,N_20139,N_20368);
nand U21020 (N_21020,N_20382,N_19660);
and U21021 (N_21021,N_19796,N_19870);
and U21022 (N_21022,N_20047,N_20131);
and U21023 (N_21023,N_19277,N_19523);
or U21024 (N_21024,N_19409,N_19578);
nor U21025 (N_21025,N_19603,N_20383);
and U21026 (N_21026,N_19683,N_19527);
xor U21027 (N_21027,N_19458,N_19460);
nand U21028 (N_21028,N_19319,N_19348);
xor U21029 (N_21029,N_19980,N_19930);
xnor U21030 (N_21030,N_19679,N_20231);
nor U21031 (N_21031,N_19770,N_20088);
or U21032 (N_21032,N_20118,N_19486);
or U21033 (N_21033,N_20309,N_19545);
nand U21034 (N_21034,N_20090,N_19975);
nor U21035 (N_21035,N_19286,N_20040);
xnor U21036 (N_21036,N_19808,N_19478);
or U21037 (N_21037,N_19942,N_20349);
nand U21038 (N_21038,N_19995,N_19486);
nor U21039 (N_21039,N_20375,N_19269);
and U21040 (N_21040,N_20136,N_19632);
nand U21041 (N_21041,N_19938,N_19763);
or U21042 (N_21042,N_19762,N_19600);
nor U21043 (N_21043,N_19498,N_19922);
and U21044 (N_21044,N_19634,N_19337);
xor U21045 (N_21045,N_20255,N_20246);
nand U21046 (N_21046,N_19758,N_20112);
xnor U21047 (N_21047,N_19641,N_19308);
or U21048 (N_21048,N_20093,N_19863);
nor U21049 (N_21049,N_19703,N_19430);
xnor U21050 (N_21050,N_20227,N_19456);
and U21051 (N_21051,N_19229,N_19390);
or U21052 (N_21052,N_19475,N_20136);
or U21053 (N_21053,N_19351,N_20054);
nand U21054 (N_21054,N_19510,N_19565);
nor U21055 (N_21055,N_20112,N_19641);
nor U21056 (N_21056,N_20220,N_20362);
and U21057 (N_21057,N_19833,N_20245);
nand U21058 (N_21058,N_19941,N_19314);
nor U21059 (N_21059,N_19987,N_19835);
nand U21060 (N_21060,N_19598,N_20269);
xnor U21061 (N_21061,N_19744,N_20184);
and U21062 (N_21062,N_19923,N_20291);
and U21063 (N_21063,N_20172,N_19252);
and U21064 (N_21064,N_20033,N_19615);
or U21065 (N_21065,N_19746,N_19852);
nand U21066 (N_21066,N_20244,N_20231);
nor U21067 (N_21067,N_19293,N_20002);
and U21068 (N_21068,N_19819,N_20265);
nand U21069 (N_21069,N_20009,N_19793);
or U21070 (N_21070,N_19557,N_19594);
or U21071 (N_21071,N_19775,N_20379);
xnor U21072 (N_21072,N_19750,N_20047);
and U21073 (N_21073,N_19787,N_19410);
or U21074 (N_21074,N_20193,N_19229);
nor U21075 (N_21075,N_19528,N_19421);
nor U21076 (N_21076,N_19347,N_20196);
nand U21077 (N_21077,N_19875,N_19586);
xnor U21078 (N_21078,N_19361,N_19293);
nor U21079 (N_21079,N_19478,N_20181);
and U21080 (N_21080,N_20113,N_19261);
and U21081 (N_21081,N_19340,N_19641);
nor U21082 (N_21082,N_19536,N_19767);
nand U21083 (N_21083,N_19674,N_19755);
nor U21084 (N_21084,N_19503,N_20195);
nor U21085 (N_21085,N_19402,N_20207);
nor U21086 (N_21086,N_19982,N_19749);
and U21087 (N_21087,N_20264,N_19242);
nand U21088 (N_21088,N_19617,N_20129);
nor U21089 (N_21089,N_19419,N_19917);
nand U21090 (N_21090,N_19282,N_20193);
nor U21091 (N_21091,N_20013,N_19912);
or U21092 (N_21092,N_20003,N_20237);
or U21093 (N_21093,N_19908,N_20151);
or U21094 (N_21094,N_19208,N_20071);
xor U21095 (N_21095,N_19649,N_19904);
and U21096 (N_21096,N_19891,N_19672);
nor U21097 (N_21097,N_20243,N_19515);
nor U21098 (N_21098,N_19876,N_19540);
xnor U21099 (N_21099,N_20185,N_20295);
xor U21100 (N_21100,N_19666,N_20158);
nand U21101 (N_21101,N_19380,N_19212);
and U21102 (N_21102,N_19214,N_20091);
nor U21103 (N_21103,N_19809,N_19383);
and U21104 (N_21104,N_20306,N_19856);
nor U21105 (N_21105,N_19625,N_19256);
nor U21106 (N_21106,N_19985,N_20234);
xnor U21107 (N_21107,N_20017,N_19449);
nor U21108 (N_21108,N_19550,N_19682);
and U21109 (N_21109,N_19965,N_19780);
and U21110 (N_21110,N_20274,N_20310);
and U21111 (N_21111,N_19536,N_20056);
or U21112 (N_21112,N_20145,N_19523);
or U21113 (N_21113,N_19555,N_19818);
nand U21114 (N_21114,N_20034,N_19296);
or U21115 (N_21115,N_19625,N_20259);
xor U21116 (N_21116,N_19980,N_20022);
and U21117 (N_21117,N_20136,N_19457);
and U21118 (N_21118,N_20296,N_19230);
xor U21119 (N_21119,N_20248,N_20251);
nor U21120 (N_21120,N_20357,N_20050);
and U21121 (N_21121,N_19425,N_19346);
xnor U21122 (N_21122,N_19673,N_19221);
xor U21123 (N_21123,N_19921,N_19735);
nand U21124 (N_21124,N_20347,N_20228);
nand U21125 (N_21125,N_19895,N_19969);
nor U21126 (N_21126,N_19227,N_19613);
nor U21127 (N_21127,N_19228,N_19740);
xnor U21128 (N_21128,N_20236,N_20267);
and U21129 (N_21129,N_19520,N_19554);
or U21130 (N_21130,N_19268,N_20014);
xnor U21131 (N_21131,N_19502,N_20163);
and U21132 (N_21132,N_19571,N_19281);
nor U21133 (N_21133,N_19278,N_19628);
xnor U21134 (N_21134,N_19295,N_19291);
xnor U21135 (N_21135,N_20211,N_20208);
and U21136 (N_21136,N_20206,N_19585);
nor U21137 (N_21137,N_19744,N_20340);
and U21138 (N_21138,N_19701,N_19948);
and U21139 (N_21139,N_20177,N_19424);
nand U21140 (N_21140,N_19422,N_20080);
nand U21141 (N_21141,N_20357,N_19923);
xnor U21142 (N_21142,N_19418,N_20015);
xor U21143 (N_21143,N_20165,N_19214);
or U21144 (N_21144,N_20118,N_19332);
nand U21145 (N_21145,N_19987,N_19854);
or U21146 (N_21146,N_19871,N_19729);
or U21147 (N_21147,N_19756,N_20313);
nand U21148 (N_21148,N_19480,N_20038);
or U21149 (N_21149,N_19369,N_19366);
nand U21150 (N_21150,N_19843,N_19674);
nand U21151 (N_21151,N_20329,N_20158);
nand U21152 (N_21152,N_19941,N_19864);
xnor U21153 (N_21153,N_19668,N_19380);
nand U21154 (N_21154,N_19885,N_20125);
xor U21155 (N_21155,N_19898,N_19925);
nand U21156 (N_21156,N_19389,N_19374);
nor U21157 (N_21157,N_19358,N_19325);
and U21158 (N_21158,N_19737,N_19674);
xor U21159 (N_21159,N_19492,N_19604);
and U21160 (N_21160,N_19861,N_19505);
or U21161 (N_21161,N_20213,N_19413);
nand U21162 (N_21162,N_19250,N_19735);
nand U21163 (N_21163,N_19574,N_19654);
or U21164 (N_21164,N_19492,N_19819);
and U21165 (N_21165,N_20256,N_19402);
nor U21166 (N_21166,N_20083,N_19755);
xnor U21167 (N_21167,N_19976,N_19718);
or U21168 (N_21168,N_20113,N_20221);
nand U21169 (N_21169,N_20280,N_20234);
or U21170 (N_21170,N_20169,N_19896);
nand U21171 (N_21171,N_19518,N_20172);
or U21172 (N_21172,N_19986,N_19229);
nor U21173 (N_21173,N_19906,N_19984);
and U21174 (N_21174,N_19420,N_19481);
nor U21175 (N_21175,N_19374,N_20003);
nor U21176 (N_21176,N_20183,N_20163);
xor U21177 (N_21177,N_19286,N_19438);
nor U21178 (N_21178,N_20272,N_19455);
or U21179 (N_21179,N_20297,N_20098);
nand U21180 (N_21180,N_19232,N_19353);
or U21181 (N_21181,N_19428,N_19864);
and U21182 (N_21182,N_19768,N_19458);
nand U21183 (N_21183,N_19915,N_19835);
nor U21184 (N_21184,N_20205,N_19781);
xor U21185 (N_21185,N_19530,N_20368);
and U21186 (N_21186,N_19355,N_20245);
and U21187 (N_21187,N_19307,N_20177);
nand U21188 (N_21188,N_20319,N_19730);
or U21189 (N_21189,N_19748,N_20018);
nand U21190 (N_21190,N_19564,N_19442);
nand U21191 (N_21191,N_19832,N_19633);
and U21192 (N_21192,N_19829,N_19416);
or U21193 (N_21193,N_20143,N_20084);
or U21194 (N_21194,N_19539,N_19270);
nand U21195 (N_21195,N_19423,N_19444);
or U21196 (N_21196,N_19720,N_19571);
and U21197 (N_21197,N_19202,N_19911);
nor U21198 (N_21198,N_20145,N_19599);
xnor U21199 (N_21199,N_19730,N_19822);
nor U21200 (N_21200,N_20294,N_19294);
nor U21201 (N_21201,N_19542,N_20333);
nor U21202 (N_21202,N_20273,N_20275);
nor U21203 (N_21203,N_20350,N_19291);
nor U21204 (N_21204,N_19262,N_19811);
and U21205 (N_21205,N_19347,N_20169);
and U21206 (N_21206,N_20099,N_19837);
or U21207 (N_21207,N_19445,N_19430);
and U21208 (N_21208,N_19699,N_20050);
nor U21209 (N_21209,N_20338,N_20286);
nand U21210 (N_21210,N_19300,N_19357);
or U21211 (N_21211,N_19544,N_19771);
nand U21212 (N_21212,N_19984,N_19345);
and U21213 (N_21213,N_19951,N_20035);
or U21214 (N_21214,N_19450,N_19264);
nand U21215 (N_21215,N_19609,N_20001);
nor U21216 (N_21216,N_19984,N_19234);
nand U21217 (N_21217,N_19785,N_19564);
xor U21218 (N_21218,N_20202,N_19421);
nand U21219 (N_21219,N_19509,N_19379);
nand U21220 (N_21220,N_19967,N_19732);
nor U21221 (N_21221,N_19985,N_19660);
xnor U21222 (N_21222,N_19876,N_20203);
xnor U21223 (N_21223,N_19788,N_19801);
and U21224 (N_21224,N_19249,N_19775);
nand U21225 (N_21225,N_19372,N_19902);
and U21226 (N_21226,N_19581,N_19459);
nor U21227 (N_21227,N_20162,N_19743);
or U21228 (N_21228,N_20032,N_19833);
nor U21229 (N_21229,N_20194,N_19439);
nor U21230 (N_21230,N_20026,N_19269);
xnor U21231 (N_21231,N_20272,N_20377);
nor U21232 (N_21232,N_19919,N_19861);
xor U21233 (N_21233,N_19362,N_19713);
or U21234 (N_21234,N_20053,N_19740);
or U21235 (N_21235,N_20214,N_19638);
nor U21236 (N_21236,N_19302,N_19792);
nand U21237 (N_21237,N_19475,N_20144);
and U21238 (N_21238,N_20324,N_20157);
or U21239 (N_21239,N_19356,N_19400);
xnor U21240 (N_21240,N_19542,N_20138);
and U21241 (N_21241,N_19602,N_19386);
xor U21242 (N_21242,N_19468,N_20154);
nand U21243 (N_21243,N_20266,N_20314);
or U21244 (N_21244,N_20335,N_19351);
nor U21245 (N_21245,N_19237,N_19328);
nor U21246 (N_21246,N_19256,N_20053);
and U21247 (N_21247,N_19987,N_19766);
or U21248 (N_21248,N_19420,N_19672);
nand U21249 (N_21249,N_19800,N_19332);
nor U21250 (N_21250,N_19201,N_19766);
nor U21251 (N_21251,N_20038,N_19289);
and U21252 (N_21252,N_20260,N_19847);
xnor U21253 (N_21253,N_19978,N_20263);
xor U21254 (N_21254,N_19781,N_20169);
nand U21255 (N_21255,N_19872,N_19412);
or U21256 (N_21256,N_19416,N_19524);
nor U21257 (N_21257,N_19884,N_20297);
or U21258 (N_21258,N_20356,N_20144);
nor U21259 (N_21259,N_20148,N_19442);
xnor U21260 (N_21260,N_19658,N_19719);
nor U21261 (N_21261,N_20328,N_19876);
nor U21262 (N_21262,N_20371,N_19826);
and U21263 (N_21263,N_19733,N_20110);
or U21264 (N_21264,N_19254,N_19532);
or U21265 (N_21265,N_19852,N_19417);
nor U21266 (N_21266,N_19873,N_19870);
xnor U21267 (N_21267,N_20304,N_19825);
and U21268 (N_21268,N_19721,N_19610);
or U21269 (N_21269,N_19449,N_20321);
nor U21270 (N_21270,N_19574,N_19378);
or U21271 (N_21271,N_20003,N_19570);
xnor U21272 (N_21272,N_20011,N_19773);
and U21273 (N_21273,N_20083,N_20324);
xor U21274 (N_21274,N_19621,N_19559);
and U21275 (N_21275,N_19853,N_20205);
xnor U21276 (N_21276,N_19953,N_19554);
or U21277 (N_21277,N_20104,N_19821);
nand U21278 (N_21278,N_19309,N_20176);
nor U21279 (N_21279,N_19943,N_19485);
nand U21280 (N_21280,N_19944,N_20241);
nand U21281 (N_21281,N_20111,N_19946);
nand U21282 (N_21282,N_20353,N_20289);
and U21283 (N_21283,N_19561,N_19315);
xor U21284 (N_21284,N_19442,N_19664);
and U21285 (N_21285,N_20331,N_20038);
nand U21286 (N_21286,N_19764,N_20161);
and U21287 (N_21287,N_20097,N_19625);
nand U21288 (N_21288,N_20371,N_19611);
xnor U21289 (N_21289,N_19612,N_19335);
nand U21290 (N_21290,N_20353,N_19427);
or U21291 (N_21291,N_19261,N_19662);
and U21292 (N_21292,N_19220,N_19440);
and U21293 (N_21293,N_19727,N_19521);
xnor U21294 (N_21294,N_19440,N_20123);
and U21295 (N_21295,N_19785,N_19911);
or U21296 (N_21296,N_19376,N_19221);
or U21297 (N_21297,N_19531,N_19411);
nand U21298 (N_21298,N_20102,N_20316);
and U21299 (N_21299,N_20095,N_20341);
nand U21300 (N_21300,N_19237,N_20258);
or U21301 (N_21301,N_19608,N_19378);
nand U21302 (N_21302,N_20274,N_19280);
or U21303 (N_21303,N_20384,N_20253);
xnor U21304 (N_21304,N_20260,N_19695);
or U21305 (N_21305,N_19610,N_19293);
and U21306 (N_21306,N_19499,N_20339);
and U21307 (N_21307,N_19313,N_20174);
and U21308 (N_21308,N_19603,N_19586);
and U21309 (N_21309,N_19764,N_19306);
and U21310 (N_21310,N_20127,N_19334);
and U21311 (N_21311,N_19419,N_20220);
and U21312 (N_21312,N_19600,N_20183);
xnor U21313 (N_21313,N_19949,N_19833);
nor U21314 (N_21314,N_19743,N_19527);
or U21315 (N_21315,N_19333,N_20272);
and U21316 (N_21316,N_19224,N_19490);
nand U21317 (N_21317,N_19509,N_19610);
and U21318 (N_21318,N_20265,N_19909);
xor U21319 (N_21319,N_20215,N_20155);
nor U21320 (N_21320,N_19555,N_19838);
xnor U21321 (N_21321,N_19519,N_19459);
nor U21322 (N_21322,N_19273,N_20230);
or U21323 (N_21323,N_19988,N_20314);
nand U21324 (N_21324,N_19219,N_20311);
nor U21325 (N_21325,N_20006,N_19274);
nand U21326 (N_21326,N_20310,N_19494);
nor U21327 (N_21327,N_19305,N_19950);
and U21328 (N_21328,N_19886,N_19847);
nor U21329 (N_21329,N_20083,N_19681);
and U21330 (N_21330,N_19925,N_20302);
or U21331 (N_21331,N_19736,N_19342);
xor U21332 (N_21332,N_19614,N_19347);
nor U21333 (N_21333,N_19733,N_19339);
xor U21334 (N_21334,N_19771,N_19303);
xor U21335 (N_21335,N_20246,N_20299);
nand U21336 (N_21336,N_20154,N_19415);
nand U21337 (N_21337,N_19989,N_19529);
nand U21338 (N_21338,N_19704,N_19633);
nand U21339 (N_21339,N_20154,N_19525);
nor U21340 (N_21340,N_19946,N_19342);
or U21341 (N_21341,N_19293,N_20390);
nor U21342 (N_21342,N_19756,N_19803);
nor U21343 (N_21343,N_19213,N_19356);
and U21344 (N_21344,N_19273,N_20341);
or U21345 (N_21345,N_19753,N_19602);
nand U21346 (N_21346,N_19466,N_20103);
nor U21347 (N_21347,N_19950,N_19749);
nand U21348 (N_21348,N_19751,N_19780);
and U21349 (N_21349,N_20064,N_19263);
nand U21350 (N_21350,N_19759,N_19899);
xor U21351 (N_21351,N_19276,N_19644);
nand U21352 (N_21352,N_19300,N_19883);
or U21353 (N_21353,N_20096,N_20185);
and U21354 (N_21354,N_20028,N_19953);
nand U21355 (N_21355,N_19343,N_19248);
or U21356 (N_21356,N_20222,N_19896);
xnor U21357 (N_21357,N_19382,N_19984);
nor U21358 (N_21358,N_19226,N_20344);
nor U21359 (N_21359,N_20204,N_19214);
xnor U21360 (N_21360,N_20228,N_19379);
or U21361 (N_21361,N_19889,N_19914);
and U21362 (N_21362,N_19232,N_19893);
nor U21363 (N_21363,N_19897,N_19542);
nor U21364 (N_21364,N_19771,N_19250);
nand U21365 (N_21365,N_19933,N_19759);
nor U21366 (N_21366,N_20333,N_19516);
xor U21367 (N_21367,N_19247,N_19358);
and U21368 (N_21368,N_19275,N_20301);
and U21369 (N_21369,N_19352,N_20206);
nand U21370 (N_21370,N_19332,N_19848);
nand U21371 (N_21371,N_19859,N_19598);
nor U21372 (N_21372,N_20393,N_19931);
nor U21373 (N_21373,N_19443,N_20115);
nand U21374 (N_21374,N_19777,N_19753);
and U21375 (N_21375,N_19506,N_19267);
nand U21376 (N_21376,N_20146,N_19562);
or U21377 (N_21377,N_19746,N_19799);
and U21378 (N_21378,N_20050,N_20332);
nor U21379 (N_21379,N_19941,N_19916);
nand U21380 (N_21380,N_19822,N_19727);
xnor U21381 (N_21381,N_19542,N_19638);
nor U21382 (N_21382,N_20181,N_20263);
nand U21383 (N_21383,N_19594,N_19457);
nor U21384 (N_21384,N_20108,N_20020);
nor U21385 (N_21385,N_20032,N_19813);
or U21386 (N_21386,N_19829,N_20393);
nor U21387 (N_21387,N_19253,N_20075);
xor U21388 (N_21388,N_19312,N_19349);
and U21389 (N_21389,N_19998,N_20195);
nand U21390 (N_21390,N_20147,N_20152);
xnor U21391 (N_21391,N_19535,N_20084);
and U21392 (N_21392,N_19897,N_19431);
and U21393 (N_21393,N_20181,N_20100);
and U21394 (N_21394,N_19267,N_19804);
and U21395 (N_21395,N_20032,N_19220);
xnor U21396 (N_21396,N_20265,N_19935);
or U21397 (N_21397,N_20209,N_20274);
nor U21398 (N_21398,N_20232,N_19832);
or U21399 (N_21399,N_20357,N_20047);
nand U21400 (N_21400,N_19306,N_19696);
xnor U21401 (N_21401,N_20176,N_20167);
and U21402 (N_21402,N_19844,N_20369);
xnor U21403 (N_21403,N_20150,N_19328);
xor U21404 (N_21404,N_19827,N_19575);
and U21405 (N_21405,N_19563,N_19721);
or U21406 (N_21406,N_19421,N_19843);
and U21407 (N_21407,N_20234,N_20213);
xor U21408 (N_21408,N_19442,N_19624);
nor U21409 (N_21409,N_19505,N_19706);
or U21410 (N_21410,N_19452,N_20026);
nor U21411 (N_21411,N_19451,N_19836);
or U21412 (N_21412,N_19286,N_20223);
nor U21413 (N_21413,N_20329,N_20236);
and U21414 (N_21414,N_20211,N_20248);
nor U21415 (N_21415,N_20287,N_19910);
xor U21416 (N_21416,N_20098,N_19564);
or U21417 (N_21417,N_19531,N_19659);
nand U21418 (N_21418,N_19547,N_19899);
xnor U21419 (N_21419,N_19418,N_19675);
xor U21420 (N_21420,N_19504,N_20360);
xor U21421 (N_21421,N_19522,N_20186);
or U21422 (N_21422,N_19352,N_19751);
or U21423 (N_21423,N_19950,N_19354);
and U21424 (N_21424,N_19613,N_19660);
xor U21425 (N_21425,N_19571,N_19371);
nor U21426 (N_21426,N_19462,N_20159);
and U21427 (N_21427,N_20028,N_19512);
nor U21428 (N_21428,N_19333,N_20226);
nor U21429 (N_21429,N_19214,N_19830);
and U21430 (N_21430,N_19900,N_19206);
nand U21431 (N_21431,N_19798,N_20113);
nor U21432 (N_21432,N_19591,N_20100);
nand U21433 (N_21433,N_19995,N_19423);
nor U21434 (N_21434,N_19741,N_19775);
nor U21435 (N_21435,N_19357,N_20275);
or U21436 (N_21436,N_19573,N_19824);
xor U21437 (N_21437,N_20060,N_19839);
nor U21438 (N_21438,N_19692,N_19552);
or U21439 (N_21439,N_19475,N_20340);
nor U21440 (N_21440,N_19673,N_19787);
xor U21441 (N_21441,N_19874,N_19633);
or U21442 (N_21442,N_20204,N_19745);
xor U21443 (N_21443,N_20185,N_20393);
or U21444 (N_21444,N_19551,N_19573);
nor U21445 (N_21445,N_19257,N_19721);
or U21446 (N_21446,N_20031,N_20037);
or U21447 (N_21447,N_20171,N_20187);
and U21448 (N_21448,N_19682,N_20269);
nor U21449 (N_21449,N_20302,N_19660);
or U21450 (N_21450,N_19437,N_20160);
nor U21451 (N_21451,N_20146,N_19255);
nand U21452 (N_21452,N_19511,N_20222);
and U21453 (N_21453,N_19679,N_19680);
nor U21454 (N_21454,N_20125,N_19792);
nand U21455 (N_21455,N_19776,N_19921);
and U21456 (N_21456,N_19239,N_19894);
or U21457 (N_21457,N_20139,N_19579);
xor U21458 (N_21458,N_19667,N_20303);
nand U21459 (N_21459,N_20042,N_19881);
nand U21460 (N_21460,N_20195,N_19823);
nor U21461 (N_21461,N_19491,N_19851);
nand U21462 (N_21462,N_19565,N_19848);
and U21463 (N_21463,N_19439,N_20018);
xor U21464 (N_21464,N_19853,N_20039);
nor U21465 (N_21465,N_19338,N_20348);
and U21466 (N_21466,N_20340,N_19530);
xor U21467 (N_21467,N_19319,N_19362);
and U21468 (N_21468,N_19642,N_19595);
or U21469 (N_21469,N_19777,N_19910);
xnor U21470 (N_21470,N_19432,N_19445);
xnor U21471 (N_21471,N_20125,N_19508);
and U21472 (N_21472,N_19988,N_19347);
nor U21473 (N_21473,N_20397,N_19559);
nand U21474 (N_21474,N_19228,N_19476);
nor U21475 (N_21475,N_19208,N_19962);
and U21476 (N_21476,N_19596,N_19231);
nand U21477 (N_21477,N_19523,N_19662);
and U21478 (N_21478,N_19215,N_19974);
and U21479 (N_21479,N_19708,N_19505);
nor U21480 (N_21480,N_20047,N_20024);
nor U21481 (N_21481,N_19852,N_19506);
or U21482 (N_21482,N_19941,N_20252);
xor U21483 (N_21483,N_19400,N_19287);
nor U21484 (N_21484,N_20006,N_19830);
and U21485 (N_21485,N_20055,N_19509);
or U21486 (N_21486,N_20318,N_19858);
and U21487 (N_21487,N_19751,N_20279);
nor U21488 (N_21488,N_20309,N_20310);
nor U21489 (N_21489,N_20369,N_19243);
nand U21490 (N_21490,N_19266,N_19868);
nor U21491 (N_21491,N_19635,N_19750);
or U21492 (N_21492,N_20345,N_19242);
and U21493 (N_21493,N_20180,N_19926);
xnor U21494 (N_21494,N_19983,N_19623);
nand U21495 (N_21495,N_19542,N_19793);
or U21496 (N_21496,N_20077,N_20066);
and U21497 (N_21497,N_19536,N_19738);
or U21498 (N_21498,N_20046,N_19353);
nor U21499 (N_21499,N_19845,N_20171);
xor U21500 (N_21500,N_19544,N_19422);
xor U21501 (N_21501,N_19708,N_19918);
xnor U21502 (N_21502,N_20315,N_19281);
nand U21503 (N_21503,N_19799,N_20372);
and U21504 (N_21504,N_19576,N_19832);
nor U21505 (N_21505,N_20168,N_19886);
nand U21506 (N_21506,N_19832,N_19744);
nor U21507 (N_21507,N_19986,N_19527);
nor U21508 (N_21508,N_19214,N_19556);
nand U21509 (N_21509,N_19579,N_20145);
nor U21510 (N_21510,N_19985,N_19359);
xor U21511 (N_21511,N_20097,N_19600);
and U21512 (N_21512,N_19740,N_19871);
xor U21513 (N_21513,N_19230,N_19207);
nand U21514 (N_21514,N_20358,N_19480);
nand U21515 (N_21515,N_19861,N_19984);
nor U21516 (N_21516,N_19755,N_19696);
or U21517 (N_21517,N_19296,N_19915);
nand U21518 (N_21518,N_19504,N_20199);
nand U21519 (N_21519,N_20202,N_19608);
or U21520 (N_21520,N_19489,N_19964);
xor U21521 (N_21521,N_19323,N_20164);
and U21522 (N_21522,N_19877,N_19201);
nor U21523 (N_21523,N_19433,N_20397);
or U21524 (N_21524,N_19695,N_19518);
nand U21525 (N_21525,N_19463,N_19285);
and U21526 (N_21526,N_19778,N_19713);
and U21527 (N_21527,N_20085,N_19369);
nor U21528 (N_21528,N_19697,N_19968);
or U21529 (N_21529,N_19615,N_19812);
xnor U21530 (N_21530,N_19767,N_19284);
xnor U21531 (N_21531,N_20149,N_20317);
xor U21532 (N_21532,N_19949,N_20200);
and U21533 (N_21533,N_19457,N_19370);
nor U21534 (N_21534,N_20354,N_20198);
nor U21535 (N_21535,N_20079,N_20009);
nand U21536 (N_21536,N_19910,N_20239);
and U21537 (N_21537,N_19853,N_20251);
xnor U21538 (N_21538,N_19244,N_19253);
xor U21539 (N_21539,N_19948,N_19271);
nor U21540 (N_21540,N_19336,N_19550);
nand U21541 (N_21541,N_19575,N_19948);
nor U21542 (N_21542,N_20230,N_19370);
or U21543 (N_21543,N_19229,N_19387);
and U21544 (N_21544,N_19611,N_19972);
and U21545 (N_21545,N_19762,N_19612);
or U21546 (N_21546,N_19399,N_19759);
or U21547 (N_21547,N_19221,N_20317);
and U21548 (N_21548,N_20263,N_19795);
or U21549 (N_21549,N_19320,N_20114);
xnor U21550 (N_21550,N_20059,N_19771);
xnor U21551 (N_21551,N_19651,N_19799);
or U21552 (N_21552,N_19846,N_19852);
xor U21553 (N_21553,N_19849,N_19655);
nor U21554 (N_21554,N_19757,N_19372);
or U21555 (N_21555,N_19564,N_19942);
nand U21556 (N_21556,N_20369,N_19857);
or U21557 (N_21557,N_20370,N_19705);
nor U21558 (N_21558,N_20309,N_19820);
nor U21559 (N_21559,N_20203,N_20122);
and U21560 (N_21560,N_20271,N_20329);
or U21561 (N_21561,N_20116,N_19505);
and U21562 (N_21562,N_19814,N_19256);
or U21563 (N_21563,N_20127,N_20317);
and U21564 (N_21564,N_19638,N_19753);
and U21565 (N_21565,N_19903,N_20263);
xnor U21566 (N_21566,N_19690,N_19625);
or U21567 (N_21567,N_19913,N_19206);
and U21568 (N_21568,N_19572,N_20020);
nand U21569 (N_21569,N_19647,N_19626);
nor U21570 (N_21570,N_19279,N_19974);
xor U21571 (N_21571,N_19736,N_19684);
nor U21572 (N_21572,N_19782,N_19275);
or U21573 (N_21573,N_19458,N_19922);
and U21574 (N_21574,N_19352,N_19542);
nand U21575 (N_21575,N_19836,N_20310);
and U21576 (N_21576,N_20004,N_20361);
and U21577 (N_21577,N_20021,N_19873);
nand U21578 (N_21578,N_20151,N_19288);
nand U21579 (N_21579,N_19632,N_19849);
and U21580 (N_21580,N_20191,N_20119);
nor U21581 (N_21581,N_19901,N_20299);
or U21582 (N_21582,N_20329,N_20007);
and U21583 (N_21583,N_19321,N_19214);
and U21584 (N_21584,N_20162,N_19448);
or U21585 (N_21585,N_20108,N_20136);
and U21586 (N_21586,N_19918,N_20244);
or U21587 (N_21587,N_19362,N_19509);
and U21588 (N_21588,N_19712,N_19799);
nor U21589 (N_21589,N_19292,N_19476);
nand U21590 (N_21590,N_19618,N_19764);
nor U21591 (N_21591,N_19930,N_19766);
nor U21592 (N_21592,N_19707,N_19357);
nand U21593 (N_21593,N_19335,N_19601);
or U21594 (N_21594,N_20365,N_19373);
nor U21595 (N_21595,N_19605,N_19742);
or U21596 (N_21596,N_20206,N_19300);
or U21597 (N_21597,N_19364,N_19394);
or U21598 (N_21598,N_19450,N_20388);
nand U21599 (N_21599,N_19942,N_20194);
nor U21600 (N_21600,N_21012,N_21033);
nand U21601 (N_21601,N_21567,N_21558);
and U21602 (N_21602,N_20996,N_20455);
xor U21603 (N_21603,N_21083,N_20418);
and U21604 (N_21604,N_20952,N_20497);
or U21605 (N_21605,N_21159,N_20929);
xor U21606 (N_21606,N_20905,N_21163);
or U21607 (N_21607,N_20627,N_21552);
nor U21608 (N_21608,N_21421,N_21042);
nor U21609 (N_21609,N_21341,N_20687);
xor U21610 (N_21610,N_21238,N_21144);
nor U21611 (N_21611,N_21371,N_21284);
nand U21612 (N_21612,N_20628,N_21126);
nor U21613 (N_21613,N_21069,N_21576);
and U21614 (N_21614,N_21178,N_20931);
xor U21615 (N_21615,N_21079,N_21363);
or U21616 (N_21616,N_21258,N_20988);
nor U21617 (N_21617,N_20583,N_20566);
or U21618 (N_21618,N_21278,N_21344);
xor U21619 (N_21619,N_21564,N_20726);
nand U21620 (N_21620,N_20942,N_21256);
nor U21621 (N_21621,N_20724,N_21044);
xor U21622 (N_21622,N_21264,N_21195);
or U21623 (N_21623,N_20846,N_21243);
and U21624 (N_21624,N_21285,N_20619);
and U21625 (N_21625,N_20748,N_20880);
nand U21626 (N_21626,N_20705,N_21336);
nand U21627 (N_21627,N_20556,N_21403);
nand U21628 (N_21628,N_20822,N_21112);
nor U21629 (N_21629,N_21132,N_20993);
xor U21630 (N_21630,N_21067,N_21034);
nand U21631 (N_21631,N_20449,N_21321);
and U21632 (N_21632,N_21490,N_20768);
and U21633 (N_21633,N_20648,N_21199);
nand U21634 (N_21634,N_21375,N_21223);
xor U21635 (N_21635,N_20960,N_20432);
or U21636 (N_21636,N_21398,N_20824);
nand U21637 (N_21637,N_20843,N_20511);
or U21638 (N_21638,N_20832,N_20646);
or U21639 (N_21639,N_21347,N_21152);
nand U21640 (N_21640,N_21242,N_21145);
nand U21641 (N_21641,N_20489,N_20634);
and U21642 (N_21642,N_21353,N_21110);
or U21643 (N_21643,N_20459,N_20538);
xor U21644 (N_21644,N_21364,N_20710);
nand U21645 (N_21645,N_21376,N_21198);
nor U21646 (N_21646,N_21357,N_20468);
and U21647 (N_21647,N_20563,N_21451);
or U21648 (N_21648,N_20947,N_21460);
xor U21649 (N_21649,N_20678,N_20503);
nand U21650 (N_21650,N_21372,N_20829);
nor U21651 (N_21651,N_21032,N_20665);
and U21652 (N_21652,N_21596,N_21471);
xnor U21653 (N_21653,N_20883,N_20464);
nor U21654 (N_21654,N_20903,N_20407);
xnor U21655 (N_21655,N_21327,N_20535);
or U21656 (N_21656,N_21399,N_21547);
nor U21657 (N_21657,N_20744,N_21131);
or U21658 (N_21658,N_21158,N_21501);
xor U21659 (N_21659,N_21052,N_20991);
or U21660 (N_21660,N_20777,N_21526);
or U21661 (N_21661,N_21397,N_21387);
xnor U21662 (N_21662,N_20488,N_21553);
nand U21663 (N_21663,N_21239,N_20995);
nand U21664 (N_21664,N_21443,N_21568);
and U21665 (N_21665,N_20764,N_20486);
xnor U21666 (N_21666,N_21200,N_20805);
nor U21667 (N_21667,N_20827,N_21165);
or U21668 (N_21668,N_20708,N_21204);
or U21669 (N_21669,N_20601,N_21454);
nand U21670 (N_21670,N_20636,N_21280);
and U21671 (N_21671,N_20493,N_21154);
or U21672 (N_21672,N_21486,N_20474);
xnor U21673 (N_21673,N_21205,N_21367);
and U21674 (N_21674,N_21080,N_21217);
and U21675 (N_21675,N_21170,N_21149);
nor U21676 (N_21676,N_20850,N_21493);
nand U21677 (N_21677,N_21188,N_21477);
nand U21678 (N_21678,N_21293,N_21054);
nand U21679 (N_21679,N_21255,N_21107);
nand U21680 (N_21680,N_21301,N_21449);
nor U21681 (N_21681,N_20879,N_20997);
xor U21682 (N_21682,N_20500,N_20689);
nor U21683 (N_21683,N_20626,N_20783);
nand U21684 (N_21684,N_20616,N_21410);
nor U21685 (N_21685,N_21361,N_21459);
or U21686 (N_21686,N_21378,N_21402);
xnor U21687 (N_21687,N_21318,N_21478);
or U21688 (N_21688,N_20809,N_21431);
xnor U21689 (N_21689,N_21434,N_20732);
or U21690 (N_21690,N_20717,N_21332);
or U21691 (N_21691,N_21342,N_20467);
or U21692 (N_21692,N_20696,N_20450);
xor U21693 (N_21693,N_20693,N_20526);
nand U21694 (N_21694,N_21190,N_21382);
xnor U21695 (N_21695,N_20871,N_20965);
nand U21696 (N_21696,N_21545,N_21295);
and U21697 (N_21697,N_21540,N_20508);
and U21698 (N_21698,N_21550,N_20772);
xnor U21699 (N_21699,N_21005,N_21302);
nand U21700 (N_21700,N_20800,N_20999);
and U21701 (N_21701,N_21051,N_21157);
or U21702 (N_21702,N_20845,N_21294);
and U21703 (N_21703,N_20848,N_20752);
nand U21704 (N_21704,N_21554,N_20913);
xor U21705 (N_21705,N_21487,N_20823);
nand U21706 (N_21706,N_21053,N_20596);
or U21707 (N_21707,N_21134,N_20509);
nand U21708 (N_21708,N_21578,N_20498);
xnor U21709 (N_21709,N_20760,N_21214);
and U21710 (N_21710,N_21368,N_21580);
nand U21711 (N_21711,N_20941,N_21024);
nor U21712 (N_21712,N_21062,N_20821);
or U21713 (N_21713,N_21193,N_20719);
and U21714 (N_21714,N_21068,N_20590);
nand U21715 (N_21715,N_21065,N_21337);
or U21716 (N_21716,N_20715,N_21511);
nor U21717 (N_21717,N_20423,N_20766);
xnor U21718 (N_21718,N_20876,N_21524);
or U21719 (N_21719,N_20698,N_20501);
and U21720 (N_21720,N_21521,N_21581);
xor U21721 (N_21721,N_21356,N_21251);
or U21722 (N_21722,N_20473,N_20944);
or U21723 (N_21723,N_21424,N_20651);
nand U21724 (N_21724,N_21074,N_20557);
nor U21725 (N_21725,N_21426,N_20525);
nand U21726 (N_21726,N_20638,N_20551);
nor U21727 (N_21727,N_20516,N_20674);
nand U21728 (N_21728,N_21324,N_20666);
nand U21729 (N_21729,N_20737,N_21279);
or U21730 (N_21730,N_20412,N_21537);
or U21731 (N_21731,N_21202,N_20523);
nand U21732 (N_21732,N_21452,N_21435);
nand U21733 (N_21733,N_21287,N_20973);
nor U21734 (N_21734,N_20611,N_20537);
and U21735 (N_21735,N_20544,N_21589);
nand U21736 (N_21736,N_20998,N_20411);
nand U21737 (N_21737,N_21555,N_21076);
and U21738 (N_21738,N_21089,N_21234);
or U21739 (N_21739,N_21441,N_20452);
nand U21740 (N_21740,N_20545,N_20830);
and U21741 (N_21741,N_21465,N_21470);
nor U21742 (N_21742,N_20495,N_20750);
nor U21743 (N_21743,N_21182,N_20925);
or U21744 (N_21744,N_20703,N_21007);
xor U21745 (N_21745,N_21308,N_20499);
nor U21746 (N_21746,N_20527,N_21040);
nand U21747 (N_21747,N_20533,N_20416);
nand U21748 (N_21748,N_20856,N_20943);
or U21749 (N_21749,N_20740,N_21420);
nor U21750 (N_21750,N_21483,N_20854);
nand U21751 (N_21751,N_21320,N_21267);
nand U21752 (N_21752,N_21469,N_21139);
and U21753 (N_21753,N_20958,N_21050);
and U21754 (N_21754,N_20536,N_21366);
xnor U21755 (N_21755,N_20797,N_21395);
nor U21756 (N_21756,N_20977,N_20658);
or U21757 (N_21757,N_20804,N_21014);
or U21758 (N_21758,N_21522,N_21533);
nand U21759 (N_21759,N_20409,N_20463);
and U21760 (N_21760,N_21077,N_20655);
nor U21761 (N_21761,N_21586,N_20915);
xor U21762 (N_21762,N_21212,N_21473);
nor U21763 (N_21763,N_20962,N_21060);
nand U21764 (N_21764,N_21096,N_20639);
or U21765 (N_21765,N_21240,N_20801);
nand U21766 (N_21766,N_20948,N_20788);
xnor U21767 (N_21767,N_20600,N_21381);
or U21768 (N_21768,N_20755,N_21230);
nand U21769 (N_21769,N_21528,N_21281);
or U21770 (N_21770,N_21343,N_21128);
xnor U21771 (N_21771,N_21447,N_21373);
nor U21772 (N_21772,N_20951,N_21146);
nor U21773 (N_21773,N_21500,N_21006);
nand U21774 (N_21774,N_21036,N_21136);
nor U21775 (N_21775,N_20402,N_21057);
and U21776 (N_21776,N_21481,N_21135);
or U21777 (N_21777,N_21197,N_20881);
or U21778 (N_21778,N_21098,N_20555);
nor U21779 (N_21779,N_21291,N_20751);
and U21780 (N_21780,N_20625,N_20866);
xor U21781 (N_21781,N_21229,N_20673);
nor U21782 (N_21782,N_20796,N_20442);
nor U21783 (N_21783,N_20733,N_20632);
and U21784 (N_21784,N_20849,N_20613);
nor U21785 (N_21785,N_21133,N_21520);
xor U21786 (N_21786,N_21549,N_20546);
nor U21787 (N_21787,N_20579,N_21075);
or U21788 (N_21788,N_21322,N_21506);
nand U21789 (N_21789,N_21249,N_20835);
nand U21790 (N_21790,N_20707,N_20818);
or U21791 (N_21791,N_21020,N_20863);
nor U21792 (N_21792,N_20685,N_20400);
and U21793 (N_21793,N_20867,N_20743);
nor U21794 (N_21794,N_20424,N_20940);
and U21795 (N_21795,N_20790,N_20812);
xnor U21796 (N_21796,N_21400,N_21315);
nor U21797 (N_21797,N_20736,N_20885);
nand U21798 (N_21798,N_20815,N_21411);
nand U21799 (N_21799,N_20587,N_20695);
and U21800 (N_21800,N_20574,N_20819);
or U21801 (N_21801,N_20785,N_21233);
nor U21802 (N_21802,N_20820,N_20584);
and U21803 (N_21803,N_21358,N_21235);
and U21804 (N_21804,N_20969,N_21335);
xnor U21805 (N_21805,N_20979,N_20485);
nor U21806 (N_21806,N_21252,N_20923);
nor U21807 (N_21807,N_20445,N_21408);
or U21808 (N_21808,N_20742,N_20477);
and U21809 (N_21809,N_21140,N_20427);
nor U21810 (N_21810,N_21307,N_20599);
xor U21811 (N_21811,N_21265,N_21203);
nor U21812 (N_21812,N_20478,N_21531);
xor U21813 (N_21813,N_20562,N_20496);
xnor U21814 (N_21814,N_21365,N_21438);
nand U21815 (N_21815,N_20571,N_21428);
and U21816 (N_21816,N_20623,N_20505);
nor U21817 (N_21817,N_21104,N_21328);
and U21818 (N_21818,N_21565,N_21406);
or U21819 (N_21819,N_20921,N_20592);
xor U21820 (N_21820,N_20482,N_20875);
nand U21821 (N_21821,N_20422,N_21466);
or U21822 (N_21822,N_20614,N_20549);
and U21823 (N_21823,N_21515,N_21563);
nand U21824 (N_21824,N_21458,N_20591);
xnor U21825 (N_21825,N_21008,N_21560);
and U21826 (N_21826,N_20607,N_21495);
and U21827 (N_21827,N_20519,N_20847);
xor U21828 (N_21828,N_20435,N_20798);
and U21829 (N_21829,N_21121,N_20458);
nor U21830 (N_21830,N_20730,N_20679);
or U21831 (N_21831,N_20887,N_20837);
nor U21832 (N_21832,N_20975,N_20582);
xnor U21833 (N_21833,N_21569,N_20520);
and U21834 (N_21834,N_21031,N_21268);
xnor U21835 (N_21835,N_20775,N_21215);
or U21836 (N_21836,N_21102,N_21009);
nand U21837 (N_21837,N_20677,N_21226);
and U21838 (N_21838,N_20441,N_21177);
nor U21839 (N_21839,N_20690,N_21507);
and U21840 (N_21840,N_20568,N_21496);
nand U21841 (N_21841,N_21021,N_21038);
nand U21842 (N_21842,N_21409,N_21385);
or U21843 (N_21843,N_21220,N_20675);
nand U21844 (N_21844,N_21290,N_21105);
nor U21845 (N_21845,N_20753,N_21173);
or U21846 (N_21846,N_21196,N_20859);
nand U21847 (N_21847,N_21108,N_20428);
nor U21848 (N_21848,N_20460,N_21359);
and U21849 (N_21849,N_21035,N_20565);
nor U21850 (N_21850,N_21303,N_21599);
xnor U21851 (N_21851,N_21103,N_21260);
and U21852 (N_21852,N_20963,N_20990);
and U21853 (N_21853,N_20652,N_21266);
xor U21854 (N_21854,N_20763,N_20588);
xnor U21855 (N_21855,N_21194,N_21039);
or U21856 (N_21856,N_20774,N_21116);
and U21857 (N_21857,N_21244,N_21000);
and U21858 (N_21858,N_20589,N_21001);
and U21859 (N_21859,N_20810,N_21527);
nor U21860 (N_21860,N_20624,N_21575);
and U21861 (N_21861,N_20932,N_20984);
nor U21862 (N_21862,N_21429,N_21374);
nand U21863 (N_21863,N_20831,N_20598);
nand U21864 (N_21864,N_20955,N_20443);
nand U21865 (N_21865,N_21319,N_20781);
nand U21866 (N_21866,N_21254,N_21418);
xnor U21867 (N_21867,N_21587,N_20640);
and U21868 (N_21868,N_21043,N_20976);
or U21869 (N_21869,N_21172,N_20686);
nor U21870 (N_21870,N_20912,N_21440);
nand U21871 (N_21871,N_20425,N_20731);
xnor U21872 (N_21872,N_21088,N_20811);
or U21873 (N_21873,N_21415,N_21407);
or U21874 (N_21874,N_20992,N_21384);
and U21875 (N_21875,N_21480,N_21432);
nand U21876 (N_21876,N_21461,N_21349);
or U21877 (N_21877,N_21138,N_21595);
nand U21878 (N_21878,N_20644,N_21472);
and U21879 (N_21879,N_20886,N_21227);
or U21880 (N_21880,N_20681,N_21147);
nand U21881 (N_21881,N_20844,N_20670);
or U21882 (N_21882,N_20808,N_20608);
and U21883 (N_21883,N_21379,N_20580);
and U21884 (N_21884,N_20662,N_20807);
nand U21885 (N_21885,N_20668,N_21518);
nand U21886 (N_21886,N_20454,N_20889);
xor U21887 (N_21887,N_21277,N_21130);
or U21888 (N_21888,N_20471,N_20688);
xor U21889 (N_21889,N_20938,N_20891);
and U21890 (N_21890,N_20758,N_21106);
nor U21891 (N_21891,N_20865,N_21354);
nor U21892 (N_21892,N_21548,N_21175);
or U21893 (N_21893,N_21257,N_20487);
and U21894 (N_21894,N_20517,N_21456);
xor U21895 (N_21895,N_21161,N_21115);
nand U21896 (N_21896,N_20694,N_20862);
xor U21897 (N_21897,N_21142,N_20709);
xnor U21898 (N_21898,N_21232,N_21562);
xnor U21899 (N_21899,N_20720,N_21445);
xnor U21900 (N_21900,N_20475,N_20833);
xor U21901 (N_21901,N_20540,N_21283);
nor U21902 (N_21902,N_20405,N_21093);
and U21903 (N_21903,N_20633,N_20767);
xnor U21904 (N_21904,N_20415,N_20577);
xnor U21905 (N_21905,N_21355,N_20602);
and U21906 (N_21906,N_21352,N_20586);
xor U21907 (N_21907,N_20739,N_20661);
xnor U21908 (N_21908,N_21391,N_20855);
nor U21909 (N_21909,N_20410,N_21591);
and U21910 (N_21910,N_20466,N_20784);
nor U21911 (N_21911,N_21476,N_20672);
and U21912 (N_21912,N_20786,N_20641);
and U21913 (N_21913,N_20572,N_21179);
xnor U21914 (N_21914,N_20869,N_21164);
nand U21915 (N_21915,N_21312,N_20792);
xnor U21916 (N_21916,N_20570,N_20595);
nor U21917 (N_21917,N_21572,N_20447);
or U21918 (N_21918,N_20649,N_20558);
or U21919 (N_21919,N_21148,N_21597);
and U21920 (N_21920,N_21166,N_20836);
xnor U21921 (N_21921,N_21081,N_21412);
nor U21922 (N_21922,N_20789,N_20895);
and U21923 (N_21923,N_21530,N_21228);
xor U21924 (N_21924,N_20567,N_21346);
nor U21925 (N_21925,N_21503,N_21248);
xnor U21926 (N_21926,N_21467,N_21143);
or U21927 (N_21927,N_21025,N_20453);
nor U21928 (N_21928,N_20906,N_21383);
nand U21929 (N_21929,N_20594,N_20515);
nor U21930 (N_21930,N_20841,N_21213);
or U21931 (N_21931,N_20461,N_20787);
and U21932 (N_21932,N_20877,N_20946);
or U21933 (N_21933,N_21123,N_20816);
and U21934 (N_21934,N_20882,N_20456);
nand U21935 (N_21935,N_21386,N_21221);
and U21936 (N_21936,N_20791,N_21329);
nor U21937 (N_21937,N_20437,N_20914);
and U21938 (N_21938,N_20989,N_20433);
nand U21939 (N_21939,N_20878,N_21072);
nand U21940 (N_21940,N_21274,N_20706);
and U21941 (N_21941,N_21369,N_20934);
and U21942 (N_21942,N_21593,N_20650);
and U21943 (N_21943,N_20770,N_21331);
and U21944 (N_21944,N_20484,N_20884);
and U21945 (N_21945,N_21180,N_20704);
nand U21946 (N_21946,N_20617,N_20585);
nand U21947 (N_21947,N_20403,N_21063);
and U21948 (N_21948,N_21022,N_21396);
nand U21949 (N_21949,N_21070,N_20725);
nor U21950 (N_21950,N_20431,N_20899);
xor U21951 (N_21951,N_20900,N_21594);
or U21952 (N_21952,N_21026,N_21086);
and U21953 (N_21953,N_21423,N_20518);
and U21954 (N_21954,N_20968,N_20683);
or U21955 (N_21955,N_20699,N_20953);
xor U21956 (N_21956,N_21117,N_20971);
and U21957 (N_21957,N_21574,N_20684);
or U21958 (N_21958,N_21219,N_20552);
and U21959 (N_21959,N_21097,N_20637);
xnor U21960 (N_21960,N_21111,N_21275);
nor U21961 (N_21961,N_20604,N_20994);
or U21962 (N_21962,N_20860,N_21512);
nand U21963 (N_21963,N_20697,N_20794);
and U21964 (N_21964,N_21253,N_21330);
and U21965 (N_21965,N_20762,N_21546);
xor U21966 (N_21966,N_21168,N_20864);
xor U21967 (N_21967,N_21150,N_20711);
nor U21968 (N_21968,N_21090,N_20956);
and U21969 (N_21969,N_21282,N_21084);
nor U21970 (N_21970,N_21125,N_20539);
nor U21971 (N_21971,N_20434,N_21417);
and U21972 (N_21972,N_21141,N_21541);
nand U21973 (N_21973,N_20701,N_21119);
nand U21974 (N_21974,N_20547,N_20978);
or U21975 (N_21975,N_21362,N_21059);
and U21976 (N_21976,N_20669,N_21120);
or U21977 (N_21977,N_20676,N_21183);
and U21978 (N_21978,N_21049,N_21245);
nor U21979 (N_21979,N_20605,N_21448);
nor U21980 (N_21980,N_20754,N_21311);
nand U21981 (N_21981,N_20723,N_20982);
nor U21982 (N_21982,N_20561,N_20840);
or U21983 (N_21983,N_21113,N_21210);
or U21984 (N_21984,N_21151,N_21078);
xor U21985 (N_21985,N_21351,N_20512);
xnor U21986 (N_21986,N_20890,N_20436);
nor U21987 (N_21987,N_20735,N_21534);
and U21988 (N_21988,N_20950,N_20597);
xor U21989 (N_21989,N_20448,N_20911);
and U21990 (N_21990,N_21450,N_20825);
or U21991 (N_21991,N_20747,N_21551);
or U21992 (N_21992,N_21455,N_21047);
and U21993 (N_21993,N_20813,N_20964);
nor U21994 (N_21994,N_21442,N_21394);
and U21995 (N_21995,N_20575,N_21114);
and U21996 (N_21996,N_21348,N_21488);
and U21997 (N_21997,N_21066,N_20446);
xnor U21998 (N_21998,N_21339,N_20749);
or U21999 (N_21999,N_20761,N_20653);
nor U22000 (N_22000,N_20606,N_20927);
nor U22001 (N_22001,N_20874,N_21590);
nand U22002 (N_22002,N_20635,N_21262);
nand U22003 (N_22003,N_21388,N_21457);
xnor U22004 (N_22004,N_21377,N_21504);
or U22005 (N_22005,N_21389,N_20907);
xor U22006 (N_22006,N_21211,N_21261);
and U22007 (N_22007,N_21422,N_20550);
nor U22008 (N_22008,N_21027,N_20507);
nand U22009 (N_22009,N_20799,N_21118);
and U22010 (N_22010,N_20838,N_21216);
or U22011 (N_22011,N_21246,N_20554);
or U22012 (N_22012,N_20985,N_21030);
or U22013 (N_22013,N_21316,N_20406);
and U22014 (N_22014,N_21505,N_21538);
xor U22015 (N_22015,N_21297,N_20986);
nor U22016 (N_22016,N_20439,N_20691);
nor U22017 (N_22017,N_20667,N_20759);
nand U22018 (N_22018,N_20657,N_21559);
or U22019 (N_22019,N_21498,N_21122);
nand U22020 (N_22020,N_21092,N_20444);
nand U22021 (N_22021,N_21491,N_20462);
or U22022 (N_22022,N_20842,N_21543);
and U22023 (N_22023,N_21592,N_21517);
xnor U22024 (N_22024,N_21259,N_20414);
xnor U22025 (N_22025,N_20893,N_20472);
nor U22026 (N_22026,N_21071,N_21174);
or U22027 (N_22027,N_20937,N_21087);
or U22028 (N_22028,N_20618,N_21288);
and U22029 (N_22029,N_21588,N_20802);
or U22030 (N_22030,N_20839,N_20404);
or U22031 (N_22031,N_21037,N_21162);
or U22032 (N_22032,N_20778,N_20541);
and U22033 (N_22033,N_20757,N_20528);
nand U22034 (N_22034,N_21082,N_21208);
and U22035 (N_22035,N_21045,N_21181);
xor U22036 (N_22036,N_20873,N_20479);
and U22037 (N_22037,N_21556,N_20620);
nand U22038 (N_22038,N_21317,N_21479);
nor U22039 (N_22039,N_21323,N_21276);
nor U22040 (N_22040,N_20987,N_21514);
and U22041 (N_22041,N_20957,N_20714);
nand U22042 (N_22042,N_21091,N_20569);
and U22043 (N_22043,N_21156,N_21513);
nor U22044 (N_22044,N_20920,N_21313);
nor U22045 (N_22045,N_21444,N_20700);
and U22046 (N_22046,N_20573,N_20776);
xnor U22047 (N_22047,N_21425,N_21056);
or U22048 (N_22048,N_21536,N_20560);
xor U22049 (N_22049,N_20896,N_20413);
or U22050 (N_22050,N_21094,N_20936);
nand U22051 (N_22051,N_21101,N_20902);
xnor U22052 (N_22052,N_20967,N_21304);
or U22053 (N_22053,N_20919,N_21224);
nand U22054 (N_22054,N_20659,N_21340);
nor U22055 (N_22055,N_20918,N_21502);
nor U22056 (N_22056,N_21222,N_21338);
xor U22057 (N_22057,N_20401,N_20513);
or U22058 (N_22058,N_21334,N_21430);
and U22059 (N_22059,N_20481,N_21207);
and U22060 (N_22060,N_21539,N_21137);
nand U22061 (N_22061,N_21237,N_21029);
and U22062 (N_22062,N_20780,N_20692);
or U22063 (N_22063,N_20622,N_21011);
nor U22064 (N_22064,N_20852,N_21160);
or U22065 (N_22065,N_20904,N_21585);
xor U22066 (N_22066,N_20782,N_20532);
or U22067 (N_22067,N_20745,N_20916);
xnor U22068 (N_22068,N_20609,N_20974);
nand U22069 (N_22069,N_20972,N_20712);
and U22070 (N_22070,N_21250,N_21015);
xnor U22071 (N_22071,N_21484,N_20949);
and U22072 (N_22072,N_21298,N_20945);
or U22073 (N_22073,N_20510,N_21129);
xnor U22074 (N_22074,N_20421,N_21273);
nor U22075 (N_22075,N_20793,N_20576);
and U22076 (N_22076,N_21350,N_21299);
or U22077 (N_22077,N_21176,N_21532);
and U22078 (N_22078,N_21271,N_20734);
nor U22079 (N_22079,N_21463,N_20621);
nand U22080 (N_22080,N_20491,N_20542);
and U22081 (N_22081,N_21492,N_20480);
nor U22082 (N_22082,N_21535,N_20983);
and U22083 (N_22083,N_20728,N_20476);
or U22084 (N_22084,N_21579,N_21064);
nor U22085 (N_22085,N_21292,N_20814);
nand U22086 (N_22086,N_20494,N_21414);
nor U22087 (N_22087,N_20910,N_21542);
xnor U22088 (N_22088,N_21437,N_20769);
or U22089 (N_22089,N_21345,N_21416);
nand U22090 (N_22090,N_21523,N_20664);
nor U22091 (N_22091,N_21085,N_20660);
xor U22092 (N_22092,N_21055,N_21169);
and U22093 (N_22093,N_20828,N_21494);
or U22094 (N_22094,N_21392,N_20917);
nor U22095 (N_22095,N_21048,N_20935);
nor U22096 (N_22096,N_21582,N_20765);
nor U22097 (N_22097,N_21405,N_21003);
nand U22098 (N_22098,N_20451,N_21419);
nor U22099 (N_22099,N_21571,N_20746);
nand U22100 (N_22100,N_21557,N_21510);
nand U22101 (N_22101,N_20438,N_21439);
nor U22102 (N_22102,N_21573,N_20612);
nand U22103 (N_22103,N_21413,N_21270);
xnor U22104 (N_22104,N_20771,N_21446);
xor U22105 (N_22105,N_21225,N_20506);
nor U22106 (N_22106,N_21529,N_20966);
nor U22107 (N_22107,N_21013,N_20522);
nand U22108 (N_22108,N_20631,N_20908);
or U22109 (N_22109,N_20870,N_21171);
or U22110 (N_22110,N_21186,N_20469);
xnor U22111 (N_22111,N_21241,N_21497);
nand U22112 (N_22112,N_21247,N_20564);
xnor U22113 (N_22113,N_20716,N_21236);
and U22114 (N_22114,N_20826,N_21436);
nand U22115 (N_22115,N_20857,N_20663);
nor U22116 (N_22116,N_21427,N_20718);
and U22117 (N_22117,N_20817,N_21028);
xnor U22118 (N_22118,N_21489,N_21453);
or U22119 (N_22119,N_21577,N_20898);
or U22120 (N_22120,N_20702,N_21192);
nor U22121 (N_22121,N_21390,N_21201);
xnor U22122 (N_22122,N_20642,N_20514);
nand U22123 (N_22123,N_21468,N_20529);
xor U22124 (N_22124,N_21561,N_20954);
nor U22125 (N_22125,N_20901,N_20713);
or U22126 (N_22126,N_21499,N_20970);
nand U22127 (N_22127,N_20593,N_20470);
and U22128 (N_22128,N_20680,N_20795);
and U22129 (N_22129,N_20922,N_20806);
xnor U22130 (N_22130,N_21004,N_20543);
and U22131 (N_22131,N_21041,N_20853);
xor U22132 (N_22132,N_21109,N_21095);
xor U22133 (N_22133,N_20483,N_20417);
and U22134 (N_22134,N_21509,N_20615);
and U22135 (N_22135,N_20722,N_21019);
or U22136 (N_22136,N_21016,N_20980);
and U22137 (N_22137,N_20408,N_21218);
nor U22138 (N_22138,N_20531,N_20741);
xnor U22139 (N_22139,N_20779,N_21401);
nor U22140 (N_22140,N_21464,N_21516);
or U22141 (N_22141,N_21127,N_20897);
nand U22142 (N_22142,N_20868,N_20430);
nand U22143 (N_22143,N_21380,N_21570);
and U22144 (N_22144,N_21010,N_20656);
or U22145 (N_22145,N_21309,N_20727);
or U22146 (N_22146,N_21475,N_20872);
or U22147 (N_22147,N_20524,N_21508);
nand U22148 (N_22148,N_21360,N_21404);
xor U22149 (N_22149,N_21286,N_21289);
or U22150 (N_22150,N_20803,N_21058);
xor U22151 (N_22151,N_20610,N_21314);
or U22152 (N_22152,N_20534,N_21370);
or U22153 (N_22153,N_21474,N_20420);
nand U22154 (N_22154,N_20490,N_20581);
nor U22155 (N_22155,N_20981,N_21269);
xnor U22156 (N_22156,N_21100,N_20603);
and U22157 (N_22157,N_21525,N_20933);
or U22158 (N_22158,N_20930,N_21584);
nor U22159 (N_22159,N_20721,N_21333);
and U22160 (N_22160,N_21023,N_20504);
nand U22161 (N_22161,N_20926,N_21187);
nor U22162 (N_22162,N_21300,N_20548);
nor U22163 (N_22163,N_21153,N_21306);
nand U22164 (N_22164,N_21099,N_20861);
nor U22165 (N_22165,N_20671,N_21017);
xor U22166 (N_22166,N_21184,N_20851);
xor U22167 (N_22167,N_20888,N_20457);
or U22168 (N_22168,N_21544,N_21598);
or U22169 (N_22169,N_21002,N_20939);
xnor U22170 (N_22170,N_20440,N_21073);
nor U22171 (N_22171,N_21305,N_20729);
or U22172 (N_22172,N_20924,N_21482);
nor U22173 (N_22173,N_20909,N_20834);
xnor U22174 (N_22174,N_20892,N_21191);
xnor U22175 (N_22175,N_20521,N_21185);
xnor U22176 (N_22176,N_20773,N_21263);
xor U22177 (N_22177,N_21326,N_20429);
or U22178 (N_22178,N_21018,N_21189);
xnor U22179 (N_22179,N_21046,N_21462);
xnor U22180 (N_22180,N_21566,N_20465);
or U22181 (N_22181,N_21325,N_21310);
nand U22182 (N_22182,N_21124,N_20578);
nand U22183 (N_22183,N_20426,N_21272);
or U22184 (N_22184,N_20756,N_21209);
xor U22185 (N_22185,N_20559,N_21393);
nand U22186 (N_22186,N_20654,N_20961);
or U22187 (N_22187,N_20629,N_20858);
nor U22188 (N_22188,N_20419,N_20959);
and U22189 (N_22189,N_20553,N_21519);
and U22190 (N_22190,N_21155,N_20647);
or U22191 (N_22191,N_21061,N_21167);
nor U22192 (N_22192,N_21583,N_21433);
nor U22193 (N_22193,N_20643,N_21485);
nand U22194 (N_22194,N_20928,N_20738);
or U22195 (N_22195,N_20492,N_20630);
nor U22196 (N_22196,N_20645,N_20502);
nand U22197 (N_22197,N_21231,N_21206);
and U22198 (N_22198,N_21296,N_20530);
nor U22199 (N_22199,N_20682,N_20894);
nor U22200 (N_22200,N_20474,N_21280);
nor U22201 (N_22201,N_21243,N_21298);
or U22202 (N_22202,N_20720,N_20731);
nand U22203 (N_22203,N_20887,N_21158);
and U22204 (N_22204,N_21159,N_20434);
xor U22205 (N_22205,N_20848,N_21031);
nand U22206 (N_22206,N_21008,N_20482);
or U22207 (N_22207,N_20430,N_21244);
nor U22208 (N_22208,N_20573,N_21334);
nor U22209 (N_22209,N_21190,N_20934);
xor U22210 (N_22210,N_21378,N_21019);
nand U22211 (N_22211,N_20936,N_21585);
nor U22212 (N_22212,N_21346,N_20539);
nand U22213 (N_22213,N_21566,N_20724);
nor U22214 (N_22214,N_21445,N_21009);
and U22215 (N_22215,N_20951,N_21326);
nor U22216 (N_22216,N_21513,N_21594);
nor U22217 (N_22217,N_21165,N_20512);
or U22218 (N_22218,N_21325,N_21088);
nand U22219 (N_22219,N_20418,N_21172);
xor U22220 (N_22220,N_20854,N_20407);
nand U22221 (N_22221,N_21370,N_21384);
or U22222 (N_22222,N_21098,N_20437);
or U22223 (N_22223,N_21476,N_21486);
or U22224 (N_22224,N_21145,N_21296);
nor U22225 (N_22225,N_21230,N_20527);
xor U22226 (N_22226,N_21340,N_21137);
nor U22227 (N_22227,N_20984,N_20463);
xor U22228 (N_22228,N_21127,N_20596);
nand U22229 (N_22229,N_20473,N_20722);
and U22230 (N_22230,N_20782,N_20661);
xnor U22231 (N_22231,N_21384,N_21305);
nor U22232 (N_22232,N_20977,N_21495);
nand U22233 (N_22233,N_20514,N_21380);
or U22234 (N_22234,N_20862,N_20784);
and U22235 (N_22235,N_21351,N_20703);
and U22236 (N_22236,N_20522,N_20429);
nor U22237 (N_22237,N_21048,N_20983);
and U22238 (N_22238,N_21299,N_20600);
nor U22239 (N_22239,N_21066,N_21202);
or U22240 (N_22240,N_21097,N_20765);
nand U22241 (N_22241,N_21503,N_21378);
and U22242 (N_22242,N_21449,N_21430);
xnor U22243 (N_22243,N_21292,N_21162);
and U22244 (N_22244,N_21013,N_21514);
xnor U22245 (N_22245,N_21238,N_20982);
nand U22246 (N_22246,N_20477,N_21594);
nand U22247 (N_22247,N_20460,N_21401);
xnor U22248 (N_22248,N_20446,N_20469);
nand U22249 (N_22249,N_21037,N_20882);
and U22250 (N_22250,N_20961,N_20607);
nand U22251 (N_22251,N_20459,N_21456);
nand U22252 (N_22252,N_21475,N_21355);
and U22253 (N_22253,N_20628,N_20757);
nand U22254 (N_22254,N_20711,N_21549);
nor U22255 (N_22255,N_21590,N_21077);
or U22256 (N_22256,N_21411,N_20990);
and U22257 (N_22257,N_21186,N_21538);
or U22258 (N_22258,N_21278,N_21496);
nand U22259 (N_22259,N_21339,N_20452);
nand U22260 (N_22260,N_21145,N_20927);
xnor U22261 (N_22261,N_20499,N_21068);
nor U22262 (N_22262,N_21031,N_21122);
or U22263 (N_22263,N_21172,N_20438);
and U22264 (N_22264,N_21393,N_20683);
and U22265 (N_22265,N_21151,N_20857);
and U22266 (N_22266,N_20588,N_21151);
or U22267 (N_22267,N_20547,N_20419);
or U22268 (N_22268,N_20740,N_20929);
xor U22269 (N_22269,N_20845,N_21596);
nor U22270 (N_22270,N_20574,N_20704);
nor U22271 (N_22271,N_21349,N_20443);
nand U22272 (N_22272,N_21064,N_21444);
nor U22273 (N_22273,N_21258,N_20813);
or U22274 (N_22274,N_21350,N_21595);
or U22275 (N_22275,N_20858,N_20531);
nand U22276 (N_22276,N_20699,N_20892);
xnor U22277 (N_22277,N_20827,N_21320);
xnor U22278 (N_22278,N_20733,N_21507);
nand U22279 (N_22279,N_20906,N_20688);
nor U22280 (N_22280,N_21492,N_21311);
nand U22281 (N_22281,N_21131,N_20929);
nor U22282 (N_22282,N_21309,N_21588);
and U22283 (N_22283,N_21036,N_21251);
nor U22284 (N_22284,N_21525,N_21521);
nor U22285 (N_22285,N_21086,N_21523);
nand U22286 (N_22286,N_21173,N_21576);
nor U22287 (N_22287,N_20707,N_21201);
xor U22288 (N_22288,N_21424,N_20546);
nor U22289 (N_22289,N_20882,N_21586);
nand U22290 (N_22290,N_20888,N_20688);
nand U22291 (N_22291,N_20680,N_21486);
and U22292 (N_22292,N_20982,N_20750);
nor U22293 (N_22293,N_20485,N_20831);
nor U22294 (N_22294,N_21209,N_21524);
nor U22295 (N_22295,N_20496,N_20800);
xnor U22296 (N_22296,N_20504,N_21181);
and U22297 (N_22297,N_21095,N_20416);
nor U22298 (N_22298,N_20522,N_20943);
or U22299 (N_22299,N_20928,N_21327);
nor U22300 (N_22300,N_21287,N_21495);
and U22301 (N_22301,N_21481,N_20530);
nand U22302 (N_22302,N_21206,N_20907);
nand U22303 (N_22303,N_21327,N_21107);
nand U22304 (N_22304,N_20870,N_20437);
and U22305 (N_22305,N_21365,N_20582);
or U22306 (N_22306,N_21337,N_21582);
nor U22307 (N_22307,N_21546,N_20413);
nor U22308 (N_22308,N_20782,N_20960);
nor U22309 (N_22309,N_21331,N_21426);
or U22310 (N_22310,N_20860,N_20771);
or U22311 (N_22311,N_20510,N_21415);
xor U22312 (N_22312,N_20435,N_20610);
xnor U22313 (N_22313,N_20545,N_21377);
and U22314 (N_22314,N_20505,N_21230);
nor U22315 (N_22315,N_21216,N_21273);
and U22316 (N_22316,N_21015,N_21074);
or U22317 (N_22317,N_20706,N_21108);
and U22318 (N_22318,N_21375,N_20483);
or U22319 (N_22319,N_21156,N_21050);
or U22320 (N_22320,N_20877,N_20695);
or U22321 (N_22321,N_21057,N_20910);
nor U22322 (N_22322,N_20543,N_20873);
nor U22323 (N_22323,N_20978,N_20564);
nor U22324 (N_22324,N_21489,N_21341);
nand U22325 (N_22325,N_21134,N_20416);
and U22326 (N_22326,N_20727,N_21154);
xnor U22327 (N_22327,N_21150,N_20856);
nand U22328 (N_22328,N_20601,N_21531);
xnor U22329 (N_22329,N_21326,N_21166);
and U22330 (N_22330,N_21244,N_20953);
nand U22331 (N_22331,N_20626,N_21182);
and U22332 (N_22332,N_20407,N_20981);
xor U22333 (N_22333,N_20602,N_20736);
or U22334 (N_22334,N_20766,N_21059);
nor U22335 (N_22335,N_20662,N_20576);
nand U22336 (N_22336,N_20826,N_20821);
and U22337 (N_22337,N_20498,N_20820);
xnor U22338 (N_22338,N_21073,N_20978);
nor U22339 (N_22339,N_21385,N_21534);
or U22340 (N_22340,N_21329,N_20970);
or U22341 (N_22341,N_20458,N_20632);
nor U22342 (N_22342,N_20826,N_20921);
and U22343 (N_22343,N_21373,N_20718);
nand U22344 (N_22344,N_20620,N_20609);
or U22345 (N_22345,N_21453,N_21002);
and U22346 (N_22346,N_20998,N_21531);
or U22347 (N_22347,N_20959,N_20639);
nand U22348 (N_22348,N_21506,N_20414);
nand U22349 (N_22349,N_20535,N_21347);
or U22350 (N_22350,N_20976,N_20806);
and U22351 (N_22351,N_20634,N_20547);
xor U22352 (N_22352,N_21382,N_21505);
or U22353 (N_22353,N_21312,N_21001);
nor U22354 (N_22354,N_20670,N_21525);
and U22355 (N_22355,N_20868,N_21081);
xor U22356 (N_22356,N_21567,N_20939);
nor U22357 (N_22357,N_20782,N_21160);
nor U22358 (N_22358,N_20781,N_20432);
xor U22359 (N_22359,N_20454,N_21482);
nor U22360 (N_22360,N_21089,N_20635);
xor U22361 (N_22361,N_21212,N_20510);
nand U22362 (N_22362,N_21136,N_20522);
nand U22363 (N_22363,N_20779,N_21526);
or U22364 (N_22364,N_20485,N_20816);
nand U22365 (N_22365,N_20800,N_21070);
and U22366 (N_22366,N_21346,N_20456);
or U22367 (N_22367,N_20608,N_21325);
or U22368 (N_22368,N_20948,N_20828);
nor U22369 (N_22369,N_20485,N_20923);
or U22370 (N_22370,N_20617,N_21029);
nand U22371 (N_22371,N_20481,N_21084);
nand U22372 (N_22372,N_20957,N_20563);
nor U22373 (N_22373,N_21380,N_21183);
nor U22374 (N_22374,N_21104,N_20688);
and U22375 (N_22375,N_20511,N_21395);
nor U22376 (N_22376,N_21379,N_20428);
nand U22377 (N_22377,N_20441,N_20525);
and U22378 (N_22378,N_21092,N_20877);
xor U22379 (N_22379,N_21319,N_21471);
xor U22380 (N_22380,N_21136,N_21508);
and U22381 (N_22381,N_21028,N_21446);
and U22382 (N_22382,N_20440,N_21117);
or U22383 (N_22383,N_21133,N_21148);
and U22384 (N_22384,N_21299,N_21166);
or U22385 (N_22385,N_20636,N_21376);
xor U22386 (N_22386,N_20558,N_20763);
or U22387 (N_22387,N_21516,N_21531);
nand U22388 (N_22388,N_20861,N_20701);
xnor U22389 (N_22389,N_20492,N_21480);
and U22390 (N_22390,N_20765,N_20528);
xnor U22391 (N_22391,N_20751,N_21409);
nand U22392 (N_22392,N_21294,N_21432);
nand U22393 (N_22393,N_21309,N_21519);
xor U22394 (N_22394,N_21482,N_21063);
or U22395 (N_22395,N_21325,N_21315);
nand U22396 (N_22396,N_20879,N_20454);
xnor U22397 (N_22397,N_20437,N_21266);
nor U22398 (N_22398,N_20775,N_21462);
nor U22399 (N_22399,N_21107,N_21114);
nand U22400 (N_22400,N_20645,N_20480);
nand U22401 (N_22401,N_20725,N_21133);
nor U22402 (N_22402,N_21171,N_21308);
and U22403 (N_22403,N_21521,N_21095);
nor U22404 (N_22404,N_20942,N_20472);
nand U22405 (N_22405,N_21166,N_20909);
nor U22406 (N_22406,N_20914,N_21376);
and U22407 (N_22407,N_20418,N_21552);
xnor U22408 (N_22408,N_21322,N_20624);
or U22409 (N_22409,N_21353,N_20770);
and U22410 (N_22410,N_21459,N_20767);
and U22411 (N_22411,N_21148,N_21519);
and U22412 (N_22412,N_20787,N_20719);
or U22413 (N_22413,N_21344,N_21546);
or U22414 (N_22414,N_21179,N_20850);
nor U22415 (N_22415,N_20477,N_20942);
nand U22416 (N_22416,N_20867,N_21423);
nand U22417 (N_22417,N_20856,N_21479);
nand U22418 (N_22418,N_21053,N_21000);
nor U22419 (N_22419,N_20715,N_20637);
or U22420 (N_22420,N_20739,N_21492);
xnor U22421 (N_22421,N_20644,N_21002);
and U22422 (N_22422,N_21206,N_20567);
nor U22423 (N_22423,N_21008,N_20745);
and U22424 (N_22424,N_20624,N_20401);
xor U22425 (N_22425,N_21026,N_21084);
and U22426 (N_22426,N_21592,N_20947);
and U22427 (N_22427,N_20401,N_21530);
and U22428 (N_22428,N_21267,N_21158);
xor U22429 (N_22429,N_21295,N_20566);
or U22430 (N_22430,N_21283,N_21192);
nand U22431 (N_22431,N_21591,N_21561);
xor U22432 (N_22432,N_21588,N_20943);
xor U22433 (N_22433,N_20615,N_21402);
nand U22434 (N_22434,N_20604,N_21006);
and U22435 (N_22435,N_21080,N_21308);
nand U22436 (N_22436,N_20946,N_21077);
xor U22437 (N_22437,N_20646,N_20909);
and U22438 (N_22438,N_21510,N_20829);
xor U22439 (N_22439,N_20818,N_21520);
xor U22440 (N_22440,N_21109,N_21381);
xor U22441 (N_22441,N_20842,N_20597);
nand U22442 (N_22442,N_21178,N_21578);
nand U22443 (N_22443,N_20714,N_20831);
xor U22444 (N_22444,N_21378,N_21249);
xnor U22445 (N_22445,N_20700,N_21418);
nand U22446 (N_22446,N_20829,N_21566);
or U22447 (N_22447,N_20407,N_20598);
nand U22448 (N_22448,N_21337,N_20574);
nand U22449 (N_22449,N_21409,N_21383);
xnor U22450 (N_22450,N_20970,N_21479);
or U22451 (N_22451,N_21076,N_21297);
xnor U22452 (N_22452,N_20555,N_20793);
and U22453 (N_22453,N_20985,N_20455);
xor U22454 (N_22454,N_21548,N_21123);
and U22455 (N_22455,N_21340,N_20927);
xnor U22456 (N_22456,N_21218,N_20542);
xnor U22457 (N_22457,N_20526,N_20779);
or U22458 (N_22458,N_20643,N_20613);
nor U22459 (N_22459,N_20485,N_21109);
or U22460 (N_22460,N_20799,N_21029);
nand U22461 (N_22461,N_21249,N_21482);
nand U22462 (N_22462,N_21088,N_20498);
xor U22463 (N_22463,N_21271,N_21204);
or U22464 (N_22464,N_21172,N_20896);
or U22465 (N_22465,N_20455,N_20792);
nand U22466 (N_22466,N_20826,N_20879);
nand U22467 (N_22467,N_20738,N_21101);
and U22468 (N_22468,N_21101,N_20499);
nand U22469 (N_22469,N_21401,N_21321);
xor U22470 (N_22470,N_21043,N_21284);
nand U22471 (N_22471,N_20916,N_21441);
xnor U22472 (N_22472,N_21322,N_20938);
and U22473 (N_22473,N_21557,N_20561);
or U22474 (N_22474,N_20773,N_20556);
or U22475 (N_22475,N_21155,N_21107);
or U22476 (N_22476,N_20857,N_20684);
nand U22477 (N_22477,N_20980,N_20687);
nand U22478 (N_22478,N_20418,N_20875);
or U22479 (N_22479,N_20577,N_21235);
nor U22480 (N_22480,N_21222,N_20838);
xor U22481 (N_22481,N_20864,N_20423);
and U22482 (N_22482,N_21164,N_20498);
nand U22483 (N_22483,N_20445,N_21087);
and U22484 (N_22484,N_20901,N_20424);
nand U22485 (N_22485,N_20552,N_21245);
or U22486 (N_22486,N_21178,N_21090);
and U22487 (N_22487,N_21535,N_20662);
and U22488 (N_22488,N_21164,N_20995);
and U22489 (N_22489,N_20601,N_21492);
or U22490 (N_22490,N_21171,N_20716);
nor U22491 (N_22491,N_20457,N_21264);
and U22492 (N_22492,N_21002,N_20618);
xnor U22493 (N_22493,N_21201,N_20530);
or U22494 (N_22494,N_21488,N_21361);
xnor U22495 (N_22495,N_20999,N_21536);
and U22496 (N_22496,N_20992,N_20586);
nor U22497 (N_22497,N_20806,N_21597);
xnor U22498 (N_22498,N_21004,N_20919);
or U22499 (N_22499,N_21325,N_21469);
and U22500 (N_22500,N_21448,N_21275);
or U22501 (N_22501,N_20410,N_20810);
and U22502 (N_22502,N_21084,N_20917);
nor U22503 (N_22503,N_21384,N_21141);
xor U22504 (N_22504,N_21352,N_20445);
and U22505 (N_22505,N_21480,N_20904);
xor U22506 (N_22506,N_20736,N_20797);
and U22507 (N_22507,N_20466,N_21247);
nor U22508 (N_22508,N_20810,N_20545);
and U22509 (N_22509,N_21491,N_20690);
nand U22510 (N_22510,N_21183,N_21305);
nor U22511 (N_22511,N_21532,N_20974);
or U22512 (N_22512,N_20839,N_20957);
or U22513 (N_22513,N_21151,N_20880);
xor U22514 (N_22514,N_21332,N_21483);
nand U22515 (N_22515,N_21303,N_21445);
xor U22516 (N_22516,N_21551,N_20979);
and U22517 (N_22517,N_21402,N_21025);
xor U22518 (N_22518,N_21169,N_20530);
nor U22519 (N_22519,N_20403,N_20557);
nand U22520 (N_22520,N_20873,N_21495);
xor U22521 (N_22521,N_21498,N_20548);
nor U22522 (N_22522,N_21538,N_21104);
or U22523 (N_22523,N_20407,N_21133);
xor U22524 (N_22524,N_20812,N_21498);
or U22525 (N_22525,N_20866,N_20796);
xnor U22526 (N_22526,N_20569,N_21573);
nor U22527 (N_22527,N_21350,N_20851);
or U22528 (N_22528,N_21266,N_21255);
nand U22529 (N_22529,N_20400,N_20571);
nor U22530 (N_22530,N_20409,N_21454);
nand U22531 (N_22531,N_21402,N_21299);
or U22532 (N_22532,N_21066,N_20912);
xnor U22533 (N_22533,N_20416,N_20587);
and U22534 (N_22534,N_20477,N_21212);
nand U22535 (N_22535,N_21060,N_20463);
xor U22536 (N_22536,N_20847,N_20863);
nor U22537 (N_22537,N_20400,N_20551);
or U22538 (N_22538,N_20966,N_20526);
nor U22539 (N_22539,N_20836,N_21203);
nand U22540 (N_22540,N_20688,N_20723);
nor U22541 (N_22541,N_21207,N_20826);
or U22542 (N_22542,N_20757,N_20868);
nand U22543 (N_22543,N_20555,N_21177);
nand U22544 (N_22544,N_21278,N_21233);
and U22545 (N_22545,N_20768,N_20982);
and U22546 (N_22546,N_21479,N_20556);
nor U22547 (N_22547,N_21537,N_20739);
and U22548 (N_22548,N_20944,N_20685);
xor U22549 (N_22549,N_20657,N_20833);
xnor U22550 (N_22550,N_20870,N_20898);
and U22551 (N_22551,N_20543,N_21172);
nand U22552 (N_22552,N_20524,N_20854);
and U22553 (N_22553,N_20741,N_20634);
nor U22554 (N_22554,N_20772,N_21266);
and U22555 (N_22555,N_21564,N_20592);
and U22556 (N_22556,N_20805,N_21500);
or U22557 (N_22557,N_20402,N_21015);
nand U22558 (N_22558,N_20970,N_21168);
nand U22559 (N_22559,N_21272,N_21339);
nor U22560 (N_22560,N_21498,N_20806);
or U22561 (N_22561,N_21036,N_21427);
or U22562 (N_22562,N_20757,N_20524);
xor U22563 (N_22563,N_20806,N_20613);
and U22564 (N_22564,N_21546,N_21085);
or U22565 (N_22565,N_21294,N_21227);
nor U22566 (N_22566,N_20996,N_21094);
or U22567 (N_22567,N_20575,N_21160);
and U22568 (N_22568,N_21479,N_21556);
xor U22569 (N_22569,N_21024,N_20745);
nor U22570 (N_22570,N_20639,N_21040);
or U22571 (N_22571,N_21515,N_21043);
nor U22572 (N_22572,N_21416,N_21237);
or U22573 (N_22573,N_21163,N_21292);
and U22574 (N_22574,N_21298,N_21392);
nand U22575 (N_22575,N_20480,N_21143);
nor U22576 (N_22576,N_21495,N_21321);
xor U22577 (N_22577,N_20640,N_20911);
nor U22578 (N_22578,N_21536,N_20424);
or U22579 (N_22579,N_21291,N_21506);
nor U22580 (N_22580,N_21518,N_21204);
or U22581 (N_22581,N_20796,N_20746);
nand U22582 (N_22582,N_20791,N_21233);
nand U22583 (N_22583,N_20933,N_20850);
nand U22584 (N_22584,N_20824,N_21173);
and U22585 (N_22585,N_21373,N_21240);
xor U22586 (N_22586,N_21378,N_20725);
xnor U22587 (N_22587,N_21258,N_20727);
nor U22588 (N_22588,N_21311,N_21501);
or U22589 (N_22589,N_20501,N_20900);
nand U22590 (N_22590,N_21400,N_20908);
nor U22591 (N_22591,N_20565,N_21020);
and U22592 (N_22592,N_21327,N_20665);
nor U22593 (N_22593,N_20721,N_20606);
and U22594 (N_22594,N_21305,N_21459);
or U22595 (N_22595,N_21208,N_21345);
nor U22596 (N_22596,N_20728,N_20444);
and U22597 (N_22597,N_21520,N_20685);
nor U22598 (N_22598,N_20891,N_20474);
xnor U22599 (N_22599,N_21302,N_21177);
or U22600 (N_22600,N_21382,N_21575);
nand U22601 (N_22601,N_20745,N_20766);
nor U22602 (N_22602,N_21472,N_20818);
nor U22603 (N_22603,N_20974,N_21235);
nor U22604 (N_22604,N_21573,N_20862);
nand U22605 (N_22605,N_20770,N_20862);
xor U22606 (N_22606,N_20824,N_20432);
nor U22607 (N_22607,N_21388,N_20624);
xnor U22608 (N_22608,N_21219,N_21483);
xnor U22609 (N_22609,N_20462,N_20986);
or U22610 (N_22610,N_20437,N_21026);
and U22611 (N_22611,N_21119,N_20714);
nand U22612 (N_22612,N_21519,N_21424);
and U22613 (N_22613,N_20574,N_21362);
nor U22614 (N_22614,N_20420,N_21543);
nand U22615 (N_22615,N_21180,N_21404);
and U22616 (N_22616,N_20643,N_21228);
or U22617 (N_22617,N_20885,N_20464);
nand U22618 (N_22618,N_21140,N_20408);
nand U22619 (N_22619,N_21296,N_21113);
nand U22620 (N_22620,N_20637,N_21412);
or U22621 (N_22621,N_21404,N_20455);
xor U22622 (N_22622,N_20498,N_21057);
or U22623 (N_22623,N_20776,N_20968);
and U22624 (N_22624,N_20735,N_21327);
or U22625 (N_22625,N_20656,N_20465);
nor U22626 (N_22626,N_21435,N_20531);
nor U22627 (N_22627,N_20945,N_20853);
nor U22628 (N_22628,N_21082,N_20628);
nor U22629 (N_22629,N_21349,N_20892);
nand U22630 (N_22630,N_20466,N_20727);
or U22631 (N_22631,N_20699,N_21074);
and U22632 (N_22632,N_21290,N_20997);
or U22633 (N_22633,N_21156,N_20676);
xor U22634 (N_22634,N_21474,N_21035);
nand U22635 (N_22635,N_20559,N_20413);
nand U22636 (N_22636,N_21552,N_20404);
or U22637 (N_22637,N_20679,N_21424);
xnor U22638 (N_22638,N_20875,N_20973);
and U22639 (N_22639,N_21416,N_21454);
or U22640 (N_22640,N_21256,N_20961);
or U22641 (N_22641,N_20538,N_20505);
nand U22642 (N_22642,N_20861,N_21275);
nand U22643 (N_22643,N_21154,N_20675);
or U22644 (N_22644,N_21277,N_21093);
nand U22645 (N_22645,N_20874,N_20640);
nor U22646 (N_22646,N_20402,N_21278);
nor U22647 (N_22647,N_21089,N_20464);
xnor U22648 (N_22648,N_20832,N_20682);
nor U22649 (N_22649,N_20781,N_20697);
xnor U22650 (N_22650,N_21558,N_21466);
and U22651 (N_22651,N_20614,N_20846);
and U22652 (N_22652,N_20400,N_20949);
xnor U22653 (N_22653,N_20420,N_20983);
xnor U22654 (N_22654,N_21466,N_20576);
xnor U22655 (N_22655,N_21361,N_21304);
nor U22656 (N_22656,N_21384,N_21405);
nor U22657 (N_22657,N_21429,N_20940);
nor U22658 (N_22658,N_21557,N_21488);
nand U22659 (N_22659,N_20929,N_21186);
nor U22660 (N_22660,N_21587,N_20957);
and U22661 (N_22661,N_20439,N_21093);
xor U22662 (N_22662,N_21533,N_21039);
nor U22663 (N_22663,N_21020,N_21347);
nand U22664 (N_22664,N_20904,N_20920);
or U22665 (N_22665,N_20811,N_20689);
nor U22666 (N_22666,N_21344,N_21218);
nand U22667 (N_22667,N_20967,N_20817);
or U22668 (N_22668,N_20595,N_21479);
nand U22669 (N_22669,N_20591,N_20766);
or U22670 (N_22670,N_20995,N_20781);
nor U22671 (N_22671,N_21406,N_20643);
or U22672 (N_22672,N_20646,N_20999);
and U22673 (N_22673,N_20899,N_20407);
and U22674 (N_22674,N_21541,N_20731);
nor U22675 (N_22675,N_20976,N_20967);
nor U22676 (N_22676,N_21063,N_21132);
xnor U22677 (N_22677,N_21047,N_20842);
nand U22678 (N_22678,N_20970,N_21449);
or U22679 (N_22679,N_21597,N_21234);
and U22680 (N_22680,N_20794,N_20995);
or U22681 (N_22681,N_21029,N_20645);
xor U22682 (N_22682,N_20701,N_20568);
xnor U22683 (N_22683,N_21547,N_21518);
or U22684 (N_22684,N_20560,N_20504);
nor U22685 (N_22685,N_20930,N_21131);
and U22686 (N_22686,N_20497,N_21527);
and U22687 (N_22687,N_20672,N_20784);
or U22688 (N_22688,N_21325,N_20685);
and U22689 (N_22689,N_20826,N_21088);
or U22690 (N_22690,N_21397,N_21297);
xnor U22691 (N_22691,N_20652,N_20703);
and U22692 (N_22692,N_20588,N_21111);
nor U22693 (N_22693,N_20464,N_21167);
nor U22694 (N_22694,N_21211,N_20989);
xnor U22695 (N_22695,N_20423,N_21284);
xor U22696 (N_22696,N_21382,N_21078);
nor U22697 (N_22697,N_20524,N_21128);
and U22698 (N_22698,N_20429,N_20518);
xnor U22699 (N_22699,N_21356,N_20929);
nor U22700 (N_22700,N_21413,N_20858);
nand U22701 (N_22701,N_21468,N_21083);
nor U22702 (N_22702,N_20666,N_21017);
nand U22703 (N_22703,N_21434,N_20810);
and U22704 (N_22704,N_21562,N_21042);
nand U22705 (N_22705,N_21257,N_20824);
or U22706 (N_22706,N_20942,N_21485);
or U22707 (N_22707,N_21220,N_20582);
nor U22708 (N_22708,N_20651,N_21350);
nor U22709 (N_22709,N_21540,N_21225);
or U22710 (N_22710,N_21410,N_20787);
nor U22711 (N_22711,N_21354,N_21128);
or U22712 (N_22712,N_20452,N_20824);
and U22713 (N_22713,N_21413,N_21471);
or U22714 (N_22714,N_21517,N_20955);
xor U22715 (N_22715,N_21016,N_21252);
xnor U22716 (N_22716,N_21491,N_21586);
nand U22717 (N_22717,N_21002,N_20506);
nor U22718 (N_22718,N_20627,N_20886);
or U22719 (N_22719,N_20631,N_21165);
and U22720 (N_22720,N_21127,N_21524);
and U22721 (N_22721,N_21338,N_21054);
and U22722 (N_22722,N_20658,N_20867);
nor U22723 (N_22723,N_20432,N_20430);
xor U22724 (N_22724,N_21504,N_20479);
nand U22725 (N_22725,N_21152,N_20939);
xnor U22726 (N_22726,N_20665,N_20435);
and U22727 (N_22727,N_21509,N_20479);
and U22728 (N_22728,N_21508,N_20693);
xor U22729 (N_22729,N_20984,N_20884);
or U22730 (N_22730,N_20737,N_21340);
or U22731 (N_22731,N_21251,N_21305);
or U22732 (N_22732,N_20833,N_20828);
and U22733 (N_22733,N_20549,N_21154);
nor U22734 (N_22734,N_21040,N_20537);
and U22735 (N_22735,N_21159,N_21054);
nand U22736 (N_22736,N_20609,N_20522);
nor U22737 (N_22737,N_20888,N_21552);
or U22738 (N_22738,N_21286,N_20540);
or U22739 (N_22739,N_21209,N_21029);
nand U22740 (N_22740,N_21263,N_21422);
or U22741 (N_22741,N_20565,N_21583);
xnor U22742 (N_22742,N_21463,N_21479);
nand U22743 (N_22743,N_21322,N_20744);
xor U22744 (N_22744,N_21064,N_21387);
and U22745 (N_22745,N_21043,N_21483);
or U22746 (N_22746,N_21297,N_21434);
and U22747 (N_22747,N_21549,N_21034);
and U22748 (N_22748,N_20619,N_20411);
or U22749 (N_22749,N_20458,N_20843);
nor U22750 (N_22750,N_21399,N_20938);
xnor U22751 (N_22751,N_21420,N_20658);
nor U22752 (N_22752,N_21044,N_21002);
xor U22753 (N_22753,N_21425,N_20684);
and U22754 (N_22754,N_21347,N_20529);
nor U22755 (N_22755,N_21445,N_20888);
nand U22756 (N_22756,N_21365,N_20950);
or U22757 (N_22757,N_20677,N_20466);
and U22758 (N_22758,N_20967,N_21189);
and U22759 (N_22759,N_20497,N_20503);
xor U22760 (N_22760,N_21583,N_21391);
and U22761 (N_22761,N_21407,N_21305);
xor U22762 (N_22762,N_20991,N_21059);
xor U22763 (N_22763,N_20613,N_20666);
nor U22764 (N_22764,N_20877,N_21023);
nor U22765 (N_22765,N_21505,N_21421);
and U22766 (N_22766,N_21426,N_21519);
and U22767 (N_22767,N_20632,N_21233);
nand U22768 (N_22768,N_20664,N_21467);
and U22769 (N_22769,N_20889,N_21393);
nand U22770 (N_22770,N_21391,N_20568);
or U22771 (N_22771,N_21041,N_21581);
and U22772 (N_22772,N_21241,N_21575);
nor U22773 (N_22773,N_20981,N_21077);
xnor U22774 (N_22774,N_21257,N_20927);
or U22775 (N_22775,N_21238,N_20452);
and U22776 (N_22776,N_21205,N_21438);
and U22777 (N_22777,N_21146,N_21515);
xnor U22778 (N_22778,N_21385,N_20697);
nor U22779 (N_22779,N_21113,N_21215);
or U22780 (N_22780,N_20875,N_20649);
nor U22781 (N_22781,N_20489,N_20762);
or U22782 (N_22782,N_20730,N_21590);
or U22783 (N_22783,N_20894,N_21240);
or U22784 (N_22784,N_20645,N_21013);
nor U22785 (N_22785,N_20817,N_20861);
xor U22786 (N_22786,N_21171,N_20824);
and U22787 (N_22787,N_21506,N_21062);
and U22788 (N_22788,N_21580,N_21034);
nand U22789 (N_22789,N_21341,N_21586);
nor U22790 (N_22790,N_21438,N_21496);
and U22791 (N_22791,N_21430,N_20690);
and U22792 (N_22792,N_21429,N_21495);
and U22793 (N_22793,N_20957,N_20956);
nand U22794 (N_22794,N_21194,N_20559);
or U22795 (N_22795,N_20900,N_20454);
nand U22796 (N_22796,N_21008,N_20497);
nand U22797 (N_22797,N_21211,N_20450);
and U22798 (N_22798,N_20514,N_21474);
nand U22799 (N_22799,N_21187,N_20588);
nor U22800 (N_22800,N_21698,N_21715);
and U22801 (N_22801,N_22041,N_21788);
nand U22802 (N_22802,N_22001,N_22641);
or U22803 (N_22803,N_21737,N_22584);
and U22804 (N_22804,N_22429,N_21779);
nor U22805 (N_22805,N_22455,N_22249);
and U22806 (N_22806,N_22714,N_21869);
xnor U22807 (N_22807,N_22534,N_22637);
nand U22808 (N_22808,N_21725,N_22361);
nor U22809 (N_22809,N_21927,N_21906);
xor U22810 (N_22810,N_21833,N_21603);
xnor U22811 (N_22811,N_22113,N_21935);
nor U22812 (N_22812,N_22576,N_21842);
nor U22813 (N_22813,N_22563,N_21898);
or U22814 (N_22814,N_22508,N_22524);
nand U22815 (N_22815,N_22203,N_22522);
nor U22816 (N_22816,N_22512,N_22426);
or U22817 (N_22817,N_22246,N_22515);
nand U22818 (N_22818,N_22077,N_21630);
and U22819 (N_22819,N_22171,N_21885);
xor U22820 (N_22820,N_22464,N_21621);
xor U22821 (N_22821,N_21772,N_21728);
nor U22822 (N_22822,N_21937,N_22706);
nand U22823 (N_22823,N_22782,N_22290);
nand U22824 (N_22824,N_22720,N_22540);
or U22825 (N_22825,N_22125,N_21673);
xor U22826 (N_22826,N_21993,N_22561);
xor U22827 (N_22827,N_21997,N_21735);
nand U22828 (N_22828,N_21696,N_22598);
xnor U22829 (N_22829,N_22309,N_22371);
nand U22830 (N_22830,N_22437,N_22082);
nor U22831 (N_22831,N_22240,N_22183);
xnor U22832 (N_22832,N_22003,N_22640);
nand U22833 (N_22833,N_22397,N_21734);
nand U22834 (N_22834,N_22228,N_22140);
nor U22835 (N_22835,N_22034,N_21754);
xor U22836 (N_22836,N_21675,N_22078);
and U22837 (N_22837,N_22635,N_22324);
nand U22838 (N_22838,N_22416,N_22449);
nand U22839 (N_22839,N_22732,N_22578);
or U22840 (N_22840,N_22749,N_22492);
nor U22841 (N_22841,N_22054,N_22618);
nand U22842 (N_22842,N_22157,N_21671);
xnor U22843 (N_22843,N_22353,N_22208);
nand U22844 (N_22844,N_21821,N_22334);
nor U22845 (N_22845,N_22690,N_21979);
nand U22846 (N_22846,N_21652,N_22495);
and U22847 (N_22847,N_22271,N_22647);
or U22848 (N_22848,N_21686,N_21960);
nor U22849 (N_22849,N_21990,N_22337);
xor U22850 (N_22850,N_22493,N_21877);
nor U22851 (N_22851,N_21895,N_22155);
or U22852 (N_22852,N_21773,N_21766);
xnor U22853 (N_22853,N_22322,N_22306);
and U22854 (N_22854,N_22636,N_22548);
xor U22855 (N_22855,N_22025,N_22259);
xnor U22856 (N_22856,N_22106,N_22650);
nor U22857 (N_22857,N_21792,N_21701);
xnor U22858 (N_22858,N_21981,N_22141);
or U22859 (N_22859,N_22553,N_22002);
xor U22860 (N_22860,N_21825,N_22332);
nor U22861 (N_22861,N_21782,N_22623);
nor U22862 (N_22862,N_21609,N_21670);
xnor U22863 (N_22863,N_22606,N_22651);
or U22864 (N_22864,N_21640,N_22162);
nor U22865 (N_22865,N_22533,N_22664);
xnor U22866 (N_22866,N_21819,N_22724);
nor U22867 (N_22867,N_22199,N_22787);
xnor U22868 (N_22868,N_22472,N_21957);
or U22869 (N_22869,N_21996,N_22164);
nor U22870 (N_22870,N_22719,N_22267);
nand U22871 (N_22871,N_22676,N_22317);
or U22872 (N_22872,N_22746,N_21796);
nand U22873 (N_22873,N_21864,N_22407);
or U22874 (N_22874,N_22536,N_21991);
or U22875 (N_22875,N_22212,N_21969);
nor U22876 (N_22876,N_22795,N_21827);
nor U22877 (N_22877,N_22462,N_21767);
xor U22878 (N_22878,N_22476,N_22757);
and U22879 (N_22879,N_22142,N_22594);
or U22880 (N_22880,N_21722,N_21970);
or U22881 (N_22881,N_22642,N_21843);
and U22882 (N_22882,N_22513,N_22559);
nor U22883 (N_22883,N_22277,N_22167);
xor U22884 (N_22884,N_21817,N_22575);
nor U22885 (N_22885,N_22187,N_22585);
nor U22886 (N_22886,N_22511,N_22778);
or U22887 (N_22887,N_22110,N_22065);
and U22888 (N_22888,N_22304,N_21933);
nand U22889 (N_22889,N_21758,N_22202);
and U22890 (N_22890,N_22435,N_22535);
xor U22891 (N_22891,N_21880,N_22423);
nor U22892 (N_22892,N_22530,N_22539);
and U22893 (N_22893,N_22410,N_22051);
nand U22894 (N_22894,N_22627,N_22399);
nand U22895 (N_22895,N_22252,N_22481);
and U22896 (N_22896,N_22273,N_21795);
or U22897 (N_22897,N_22008,N_22209);
nor U22898 (N_22898,N_21623,N_21915);
and U22899 (N_22899,N_21862,N_22752);
xnor U22900 (N_22900,N_21651,N_21676);
or U22901 (N_22901,N_21820,N_21672);
or U22902 (N_22902,N_22613,N_22698);
nor U22903 (N_22903,N_22204,N_21804);
nor U22904 (N_22904,N_22269,N_21811);
and U22905 (N_22905,N_22300,N_22684);
xnor U22906 (N_22906,N_22100,N_22340);
nand U22907 (N_22907,N_22088,N_21658);
or U22908 (N_22908,N_21884,N_22083);
and U22909 (N_22909,N_22031,N_21908);
and U22910 (N_22910,N_21963,N_22089);
and U22911 (N_22911,N_22079,N_22033);
and U22912 (N_22912,N_22315,N_22682);
nand U22913 (N_22913,N_21780,N_21617);
or U22914 (N_22914,N_22499,N_22130);
nor U22915 (N_22915,N_21988,N_21926);
or U22916 (N_22916,N_22438,N_22750);
xor U22917 (N_22917,N_22017,N_22289);
or U22918 (N_22918,N_21822,N_21685);
nand U22919 (N_22919,N_22781,N_22327);
or U22920 (N_22920,N_22056,N_22342);
and U22921 (N_22921,N_22663,N_21755);
nor U22922 (N_22922,N_21624,N_22629);
or U22923 (N_22923,N_22086,N_21732);
nand U22924 (N_22924,N_22726,N_22200);
and U22925 (N_22925,N_22292,N_22729);
nand U22926 (N_22926,N_22517,N_22461);
nand U22927 (N_22927,N_22264,N_22619);
nand U22928 (N_22928,N_22117,N_22700);
and U22929 (N_22929,N_22712,N_21756);
and U22930 (N_22930,N_22295,N_21622);
and U22931 (N_22931,N_22433,N_22213);
and U22932 (N_22932,N_22220,N_22677);
nor U22933 (N_22933,N_22709,N_22186);
nand U22934 (N_22934,N_22256,N_22783);
nor U22935 (N_22935,N_21687,N_22715);
nor U22936 (N_22936,N_21919,N_22689);
nor U22937 (N_22937,N_21921,N_22010);
nand U22938 (N_22938,N_21995,N_22154);
and U22939 (N_22939,N_22695,N_22731);
xnor U22940 (N_22940,N_22344,N_21816);
and U22941 (N_22941,N_22345,N_21787);
nor U22942 (N_22942,N_21809,N_22143);
and U22943 (N_22943,N_21992,N_21753);
nand U22944 (N_22944,N_22255,N_22601);
or U22945 (N_22945,N_21860,N_22582);
nand U22946 (N_22946,N_22049,N_21693);
nor U22947 (N_22947,N_21896,N_22374);
and U22948 (N_22948,N_21628,N_21920);
nand U22949 (N_22949,N_22272,N_21930);
nand U22950 (N_22950,N_22378,N_22740);
xor U22951 (N_22951,N_21646,N_22068);
or U22952 (N_22952,N_22453,N_22401);
xnor U22953 (N_22953,N_22591,N_22355);
or U22954 (N_22954,N_21914,N_22080);
nor U22955 (N_22955,N_22074,N_22149);
or U22956 (N_22956,N_22097,N_22705);
nor U22957 (N_22957,N_22391,N_22483);
xnor U22958 (N_22958,N_22330,N_22069);
nand U22959 (N_22959,N_22580,N_22674);
nor U22960 (N_22960,N_22040,N_21677);
or U22961 (N_22961,N_22620,N_21964);
or U22962 (N_22962,N_21611,N_22737);
or U22963 (N_22963,N_21974,N_22274);
and U22964 (N_22964,N_21936,N_22501);
and U22965 (N_22965,N_22741,N_22287);
and U22966 (N_22966,N_22667,N_21657);
nand U22967 (N_22967,N_21901,N_21710);
and U22968 (N_22968,N_22116,N_21961);
or U22969 (N_22969,N_22214,N_22013);
or U22970 (N_22970,N_22058,N_22331);
and U22971 (N_22971,N_22075,N_21912);
or U22972 (N_22972,N_21934,N_22136);
nor U22973 (N_22973,N_21805,N_22567);
or U22974 (N_22974,N_21859,N_22454);
and U22975 (N_22975,N_22793,N_21813);
and U22976 (N_22976,N_21695,N_22777);
xnor U22977 (N_22977,N_22526,N_22180);
nor U22978 (N_22978,N_22465,N_22450);
or U22979 (N_22979,N_22218,N_22679);
or U22980 (N_22980,N_22172,N_21784);
nor U22981 (N_22981,N_22788,N_22248);
xor U22982 (N_22982,N_22016,N_22047);
xor U22983 (N_22983,N_22656,N_22798);
or U22984 (N_22984,N_22105,N_22188);
and U22985 (N_22985,N_22538,N_22494);
nor U22986 (N_22986,N_22283,N_21789);
nor U22987 (N_22987,N_21633,N_21812);
nand U22988 (N_22988,N_22158,N_22525);
or U22989 (N_22989,N_22500,N_22456);
and U22990 (N_22990,N_21956,N_21939);
and U22991 (N_22991,N_22247,N_22092);
nor U22992 (N_22992,N_22422,N_21700);
nand U22993 (N_22993,N_22442,N_21694);
nor U22994 (N_22994,N_21600,N_21712);
nand U22995 (N_22995,N_22261,N_21691);
nand U22996 (N_22996,N_22742,N_22268);
and U22997 (N_22997,N_22792,N_22759);
and U22998 (N_22998,N_22485,N_21959);
nor U22999 (N_22999,N_22748,N_22581);
nand U23000 (N_23000,N_22614,N_22138);
xnor U23001 (N_23001,N_22329,N_21669);
or U23002 (N_23002,N_22443,N_22626);
or U23003 (N_23003,N_22021,N_22736);
xnor U23004 (N_23004,N_21840,N_22266);
nand U23005 (N_23005,N_21604,N_22560);
xor U23006 (N_23006,N_22558,N_22196);
or U23007 (N_23007,N_21650,N_22791);
nor U23008 (N_23008,N_21619,N_22572);
nand U23009 (N_23009,N_21983,N_22408);
or U23010 (N_23010,N_21713,N_22146);
nand U23011 (N_23011,N_22383,N_22160);
and U23012 (N_23012,N_21846,N_22789);
and U23013 (N_23013,N_22281,N_21994);
xnor U23014 (N_23014,N_22184,N_21891);
nor U23015 (N_23015,N_22230,N_22545);
and U23016 (N_23016,N_21972,N_21639);
and U23017 (N_23017,N_21797,N_22012);
nand U23018 (N_23018,N_22707,N_22771);
and U23019 (N_23019,N_22103,N_22451);
nor U23020 (N_23020,N_22519,N_21853);
and U23021 (N_23021,N_21897,N_22617);
nand U23022 (N_23022,N_22381,N_22367);
or U23023 (N_23023,N_22402,N_21836);
or U23024 (N_23024,N_22231,N_22071);
or U23025 (N_23025,N_21865,N_22338);
and U23026 (N_23026,N_22681,N_22648);
or U23027 (N_23027,N_21616,N_21943);
nor U23028 (N_23028,N_22109,N_21718);
or U23029 (N_23029,N_21791,N_22480);
nor U23030 (N_23030,N_22760,N_22320);
or U23031 (N_23031,N_22646,N_21966);
and U23032 (N_23032,N_22587,N_22112);
nor U23033 (N_23033,N_22615,N_21626);
and U23034 (N_23034,N_22111,N_22035);
or U23035 (N_23035,N_22593,N_21740);
xnor U23036 (N_23036,N_22504,N_21705);
or U23037 (N_23037,N_22717,N_22296);
and U23038 (N_23038,N_21602,N_22496);
xnor U23039 (N_23039,N_22745,N_21931);
nand U23040 (N_23040,N_22120,N_21913);
nand U23041 (N_23041,N_21902,N_22751);
nand U23042 (N_23042,N_21634,N_22762);
or U23043 (N_23043,N_22467,N_22301);
or U23044 (N_23044,N_22168,N_22721);
and U23045 (N_23045,N_22704,N_22521);
nor U23046 (N_23046,N_21823,N_21726);
and U23047 (N_23047,N_21803,N_21783);
nand U23048 (N_23048,N_21775,N_22032);
and U23049 (N_23049,N_22665,N_22063);
nand U23050 (N_23050,N_22232,N_22725);
nor U23051 (N_23051,N_21965,N_21882);
nor U23052 (N_23052,N_22282,N_22215);
xor U23053 (N_23053,N_22179,N_22308);
nor U23054 (N_23054,N_22257,N_22400);
xor U23055 (N_23055,N_22680,N_22101);
or U23056 (N_23056,N_22452,N_22328);
nor U23057 (N_23057,N_21973,N_21781);
or U23058 (N_23058,N_21746,N_21644);
xor U23059 (N_23059,N_21948,N_22417);
xor U23060 (N_23060,N_22191,N_22609);
nand U23061 (N_23061,N_22436,N_21759);
nand U23062 (N_23062,N_22299,N_21978);
or U23063 (N_23063,N_22389,N_22727);
or U23064 (N_23064,N_22121,N_22505);
nor U23065 (N_23065,N_21684,N_22176);
nand U23066 (N_23066,N_21774,N_21723);
and U23067 (N_23067,N_21830,N_22094);
or U23068 (N_23068,N_21757,N_21818);
and U23069 (N_23069,N_22182,N_21777);
nor U23070 (N_23070,N_22586,N_22119);
xnor U23071 (N_23071,N_21731,N_22550);
or U23072 (N_23072,N_22362,N_22592);
nor U23073 (N_23073,N_21851,N_21601);
or U23074 (N_23074,N_22258,N_22225);
xnor U23075 (N_23075,N_22786,N_22658);
or U23076 (N_23076,N_22175,N_22036);
xnor U23077 (N_23077,N_22547,N_22693);
nor U23078 (N_23078,N_22507,N_21717);
nor U23079 (N_23079,N_22661,N_22790);
or U23080 (N_23080,N_22754,N_21867);
nor U23081 (N_23081,N_21852,N_22686);
or U23082 (N_23082,N_22173,N_22672);
and U23083 (N_23083,N_22552,N_21697);
nor U23084 (N_23084,N_22118,N_21932);
nand U23085 (N_23085,N_22562,N_22769);
xor U23086 (N_23086,N_22625,N_22411);
xnor U23087 (N_23087,N_22370,N_21635);
nand U23088 (N_23088,N_21798,N_21769);
and U23089 (N_23089,N_22514,N_22703);
and U23090 (N_23090,N_22303,N_22166);
or U23091 (N_23091,N_22316,N_22102);
nand U23092 (N_23092,N_22604,N_22603);
nor U23093 (N_23093,N_21665,N_22053);
xor U23094 (N_23094,N_22350,N_22662);
or U23095 (N_23095,N_21627,N_21614);
xnor U23096 (N_23096,N_21952,N_22081);
or U23097 (N_23097,N_22730,N_21742);
and U23098 (N_23098,N_22395,N_22284);
nand U23099 (N_23099,N_22057,N_22073);
xor U23100 (N_23100,N_22628,N_21748);
and U23101 (N_23101,N_22753,N_22042);
xor U23102 (N_23102,N_22294,N_22276);
xnor U23103 (N_23103,N_21709,N_21692);
and U23104 (N_23104,N_22197,N_22000);
xnor U23105 (N_23105,N_22445,N_21968);
and U23106 (N_23106,N_22211,N_22062);
or U23107 (N_23107,N_21947,N_21987);
and U23108 (N_23108,N_22755,N_22744);
nand U23109 (N_23109,N_22201,N_22305);
xnor U23110 (N_23110,N_22134,N_22460);
or U23111 (N_23111,N_21631,N_21763);
or U23112 (N_23112,N_21660,N_22471);
and U23113 (N_23113,N_22043,N_22262);
nand U23114 (N_23114,N_22019,N_22349);
xor U23115 (N_23115,N_22368,N_22531);
xor U23116 (N_23116,N_21745,N_22660);
xnor U23117 (N_23117,N_22687,N_22696);
nor U23118 (N_23118,N_22532,N_22588);
or U23119 (N_23119,N_22775,N_22557);
nor U23120 (N_23120,N_22597,N_21719);
and U23121 (N_23121,N_21951,N_22655);
xor U23122 (N_23122,N_21662,N_22346);
xnor U23123 (N_23123,N_22336,N_22747);
or U23124 (N_23124,N_22612,N_21986);
or U23125 (N_23125,N_22392,N_22313);
nand U23126 (N_23126,N_22425,N_22242);
nor U23127 (N_23127,N_21893,N_22052);
or U23128 (N_23128,N_21708,N_22260);
nor U23129 (N_23129,N_21958,N_22288);
and U23130 (N_23130,N_21615,N_22473);
and U23131 (N_23131,N_22489,N_22607);
nor U23132 (N_23132,N_22796,N_22067);
nand U23133 (N_23133,N_22219,N_21738);
nand U23134 (N_23134,N_22321,N_22127);
nor U23135 (N_23135,N_22055,N_22520);
or U23136 (N_23136,N_22608,N_21678);
nand U23137 (N_23137,N_22333,N_22644);
xor U23138 (N_23138,N_22007,N_21873);
and U23139 (N_23139,N_22546,N_22773);
nand U23140 (N_23140,N_21883,N_22132);
or U23141 (N_23141,N_22666,N_22469);
nor U23142 (N_23142,N_22649,N_22470);
or U23143 (N_23143,N_22275,N_22030);
and U23144 (N_23144,N_22076,N_22050);
and U23145 (N_23145,N_22135,N_22236);
nand U23146 (N_23146,N_21924,N_21998);
and U23147 (N_23147,N_22551,N_22005);
xor U23148 (N_23148,N_22683,N_22066);
xnor U23149 (N_23149,N_22574,N_22434);
or U23150 (N_23150,N_22348,N_21989);
and U23151 (N_23151,N_22064,N_21858);
nand U23152 (N_23152,N_22278,N_21648);
nor U23153 (N_23153,N_22447,N_22312);
or U23154 (N_23154,N_21724,N_22799);
xor U23155 (N_23155,N_21629,N_21810);
nor U23156 (N_23156,N_21730,N_22169);
xor U23157 (N_23157,N_22446,N_22375);
xnor U23158 (N_23158,N_21929,N_22339);
or U23159 (N_23159,N_22029,N_22654);
or U23160 (N_23160,N_22060,N_22221);
nand U23161 (N_23161,N_22178,N_22291);
nand U23162 (N_23162,N_22293,N_22600);
or U23163 (N_23163,N_21977,N_21950);
nand U23164 (N_23164,N_21638,N_22390);
nand U23165 (N_23165,N_22621,N_21849);
nand U23166 (N_23166,N_21838,N_21829);
and U23167 (N_23167,N_22385,N_22554);
and U23168 (N_23168,N_21793,N_22373);
or U23169 (N_23169,N_22285,N_21702);
and U23170 (N_23170,N_22602,N_21917);
and U23171 (N_23171,N_22251,N_22205);
nor U23172 (N_23172,N_22711,N_22227);
xnor U23173 (N_23173,N_22038,N_21949);
nor U23174 (N_23174,N_22364,N_22444);
or U23175 (N_23175,N_21940,N_22095);
or U23176 (N_23176,N_22756,N_22765);
or U23177 (N_23177,N_22510,N_22688);
xor U23178 (N_23178,N_22234,N_22743);
nand U23179 (N_23179,N_22023,N_22413);
nand U23180 (N_23180,N_22718,N_22441);
xor U23181 (N_23181,N_22766,N_21982);
nor U23182 (N_23182,N_21881,N_21802);
xor U23183 (N_23183,N_22235,N_22122);
nor U23184 (N_23184,N_22194,N_22631);
or U23185 (N_23185,N_21925,N_21720);
xor U23186 (N_23186,N_22542,N_22678);
xnor U23187 (N_23187,N_22114,N_21826);
xor U23188 (N_23188,N_22670,N_22502);
nand U23189 (N_23189,N_21645,N_21688);
or U23190 (N_23190,N_22431,N_21890);
nand U23191 (N_23191,N_21668,N_22376);
or U23192 (N_23192,N_21942,N_21871);
or U23193 (N_23193,N_22384,N_22497);
nor U23194 (N_23194,N_22352,N_22009);
and U23195 (N_23195,N_22566,N_22541);
xor U23196 (N_23196,N_21834,N_21916);
xor U23197 (N_23197,N_21620,N_21945);
xor U23198 (N_23198,N_22516,N_22244);
nor U23199 (N_23199,N_21636,N_21768);
xor U23200 (N_23200,N_22466,N_22326);
nor U23201 (N_23201,N_22659,N_22430);
or U23202 (N_23202,N_22129,N_22222);
or U23203 (N_23203,N_22457,N_21607);
nand U23204 (N_23204,N_21721,N_22193);
xor U23205 (N_23205,N_22414,N_22239);
nor U23206 (N_23206,N_21855,N_21649);
xnor U23207 (N_23207,N_22366,N_21727);
nand U23208 (N_23208,N_22616,N_21806);
nand U23209 (N_23209,N_22440,N_22794);
nor U23210 (N_23210,N_22543,N_21703);
or U23211 (N_23211,N_22710,N_22137);
or U23212 (N_23212,N_21706,N_22098);
and U23213 (N_23213,N_22590,N_22772);
and U23214 (N_23214,N_22653,N_22024);
and U23215 (N_23215,N_22537,N_22128);
or U23216 (N_23216,N_21841,N_22528);
and U23217 (N_23217,N_21661,N_21610);
or U23218 (N_23218,N_22358,N_22223);
and U23219 (N_23219,N_22639,N_21962);
nor U23220 (N_23220,N_21887,N_21923);
and U23221 (N_23221,N_21976,N_22382);
and U23222 (N_23222,N_21786,N_21606);
nand U23223 (N_23223,N_22685,N_22571);
and U23224 (N_23224,N_22488,N_22174);
nand U23225 (N_23225,N_22216,N_21928);
nand U23226 (N_23226,N_22046,N_21886);
or U23227 (N_23227,N_22018,N_22280);
nor U23228 (N_23228,N_22697,N_22398);
and U23229 (N_23229,N_22377,N_22396);
nor U23230 (N_23230,N_22096,N_22409);
or U23231 (N_23231,N_21761,N_22011);
and U23232 (N_23232,N_22702,N_22104);
or U23233 (N_23233,N_22523,N_22421);
xor U23234 (N_23234,N_22151,N_22153);
nand U23235 (N_23235,N_22090,N_21953);
nand U23236 (N_23236,N_22671,N_21946);
or U23237 (N_23237,N_21866,N_22152);
xor U23238 (N_23238,N_22739,N_22486);
nand U23239 (N_23239,N_22319,N_21613);
and U23240 (N_23240,N_22403,N_22379);
nand U23241 (N_23241,N_21716,N_21655);
nand U23242 (N_23242,N_22785,N_22124);
nor U23243 (N_23243,N_21642,N_21918);
nor U23244 (N_23244,N_22701,N_21764);
xor U23245 (N_23245,N_22527,N_21922);
nor U23246 (N_23246,N_22028,N_22004);
xor U23247 (N_23247,N_22716,N_22549);
xnor U23248 (N_23248,N_22779,N_22190);
nor U23249 (N_23249,N_21828,N_22570);
or U23250 (N_23250,N_22263,N_22484);
or U23251 (N_23251,N_22091,N_22439);
nor U23252 (N_23252,N_22224,N_21659);
xor U23253 (N_23253,N_22314,N_22185);
or U23254 (N_23254,N_22694,N_21778);
and U23255 (N_23255,N_22797,N_22432);
and U23256 (N_23256,N_22226,N_21683);
nand U23257 (N_23257,N_22503,N_22238);
nor U23258 (N_23258,N_22363,N_22045);
nor U23259 (N_23259,N_21605,N_22579);
nor U23260 (N_23260,N_22144,N_21899);
or U23261 (N_23261,N_21618,N_21870);
nand U23262 (N_23262,N_22764,N_22310);
xor U23263 (N_23263,N_21868,N_22150);
xor U23264 (N_23264,N_22298,N_21888);
or U23265 (N_23265,N_22477,N_22165);
or U23266 (N_23266,N_21743,N_21625);
nor U23267 (N_23267,N_21744,N_22634);
nand U23268 (N_23268,N_21707,N_22323);
or U23269 (N_23269,N_22335,N_22487);
and U23270 (N_23270,N_22723,N_21679);
nand U23271 (N_23271,N_21835,N_22669);
nand U23272 (N_23272,N_21831,N_22633);
nor U23273 (N_23273,N_21801,N_22254);
and U23274 (N_23274,N_21656,N_22325);
or U23275 (N_23275,N_22675,N_21837);
nand U23276 (N_23276,N_22192,N_22148);
or U23277 (N_23277,N_22386,N_22630);
and U23278 (N_23278,N_22357,N_22177);
and U23279 (N_23279,N_22624,N_22084);
and U23280 (N_23280,N_22573,N_22037);
nand U23281 (N_23281,N_22768,N_22015);
or U23282 (N_23282,N_22229,N_21844);
nand U23283 (N_23283,N_21785,N_22206);
nor U23284 (N_23284,N_22428,N_21938);
or U23285 (N_23285,N_22761,N_21879);
or U23286 (N_23286,N_21876,N_21848);
nand U23287 (N_23287,N_21653,N_22595);
nor U23288 (N_23288,N_22479,N_21680);
and U23289 (N_23289,N_21663,N_22448);
nor U23290 (N_23290,N_21971,N_21892);
nor U23291 (N_23291,N_21714,N_22691);
nand U23292 (N_23292,N_21643,N_22245);
nor U23293 (N_23293,N_22115,N_22020);
xor U23294 (N_23294,N_22555,N_21790);
nand U23295 (N_23295,N_21944,N_21807);
nand U23296 (N_23296,N_22406,N_21741);
nor U23297 (N_23297,N_22093,N_21750);
xor U23298 (N_23298,N_22307,N_22354);
or U23299 (N_23299,N_22758,N_22270);
or U23300 (N_23300,N_21808,N_22347);
or U23301 (N_23301,N_22380,N_22356);
nand U23302 (N_23302,N_21681,N_21954);
xnor U23303 (N_23303,N_22404,N_22061);
xor U23304 (N_23304,N_22605,N_22145);
nor U23305 (N_23305,N_21711,N_22072);
xnor U23306 (N_23306,N_21911,N_22133);
nor U23307 (N_23307,N_21894,N_22468);
nor U23308 (N_23308,N_21900,N_22474);
xor U23309 (N_23309,N_21752,N_22123);
nand U23310 (N_23310,N_22564,N_21857);
and U23311 (N_23311,N_22770,N_21682);
xnor U23312 (N_23312,N_21907,N_22774);
and U23313 (N_23313,N_22387,N_22611);
and U23314 (N_23314,N_22596,N_21874);
nor U23315 (N_23315,N_22159,N_21861);
nand U23316 (N_23316,N_22207,N_21910);
and U23317 (N_23317,N_21751,N_21889);
xor U23318 (N_23318,N_22708,N_22728);
or U23319 (N_23319,N_21975,N_22394);
or U23320 (N_23320,N_22099,N_22343);
nor U23321 (N_23321,N_21955,N_21760);
or U23322 (N_23322,N_21839,N_21739);
nand U23323 (N_23323,N_22427,N_22735);
or U23324 (N_23324,N_21800,N_22217);
nor U23325 (N_23325,N_22643,N_21667);
nand U23326 (N_23326,N_21666,N_22070);
or U23327 (N_23327,N_22279,N_21690);
xnor U23328 (N_23328,N_22738,N_22022);
or U23329 (N_23329,N_21664,N_22302);
nor U23330 (N_23330,N_22044,N_22233);
xor U23331 (N_23331,N_22645,N_22048);
nand U23332 (N_23332,N_22565,N_22763);
xor U23333 (N_23333,N_22250,N_21674);
nand U23334 (N_23334,N_22265,N_22418);
xnor U23335 (N_23335,N_22006,N_22420);
xor U23336 (N_23336,N_22506,N_22419);
nor U23337 (N_23337,N_22297,N_21771);
and U23338 (N_23338,N_21704,N_21875);
nor U23339 (N_23339,N_22170,N_21824);
xnor U23340 (N_23340,N_21905,N_22189);
or U23341 (N_23341,N_22341,N_22589);
and U23342 (N_23342,N_22610,N_21967);
or U23343 (N_23343,N_21647,N_22014);
or U23344 (N_23344,N_22498,N_21729);
or U23345 (N_23345,N_21984,N_22622);
xnor U23346 (N_23346,N_21856,N_21854);
nand U23347 (N_23347,N_22780,N_22478);
xnor U23348 (N_23348,N_22087,N_22463);
nor U23349 (N_23349,N_22286,N_21632);
and U23350 (N_23350,N_22241,N_22556);
or U23351 (N_23351,N_22568,N_22163);
xnor U23352 (N_23352,N_22509,N_21832);
nor U23353 (N_23353,N_22156,N_21776);
nand U23354 (N_23354,N_22784,N_21749);
nor U23355 (N_23355,N_22237,N_22424);
and U23356 (N_23356,N_21999,N_21815);
nor U23357 (N_23357,N_22161,N_22482);
nor U23358 (N_23358,N_22311,N_22147);
nor U23359 (N_23359,N_22027,N_22318);
nor U23360 (N_23360,N_22393,N_22458);
or U23361 (N_23361,N_22372,N_21794);
nor U23362 (N_23362,N_22491,N_22360);
and U23363 (N_23363,N_22692,N_21814);
nand U23364 (N_23364,N_22388,N_21872);
nand U23365 (N_23365,N_22733,N_22652);
nor U23366 (N_23366,N_22351,N_22131);
and U23367 (N_23367,N_22365,N_22039);
xor U23368 (N_23368,N_22776,N_21845);
nand U23369 (N_23369,N_22668,N_22544);
nor U23370 (N_23370,N_22405,N_22734);
nor U23371 (N_23371,N_22459,N_21608);
xnor U23372 (N_23372,N_21941,N_22139);
xnor U23373 (N_23373,N_22085,N_22475);
xnor U23374 (N_23374,N_22359,N_22599);
and U23375 (N_23375,N_22673,N_22059);
nor U23376 (N_23376,N_22490,N_21641);
or U23377 (N_23377,N_22253,N_21904);
or U23378 (N_23378,N_22638,N_21799);
and U23379 (N_23379,N_21770,N_21733);
xor U23380 (N_23380,N_21612,N_21850);
or U23381 (N_23381,N_21689,N_22632);
nand U23382 (N_23382,N_22126,N_22108);
xor U23383 (N_23383,N_22699,N_22713);
xnor U23384 (N_23384,N_22412,N_22569);
nor U23385 (N_23385,N_22722,N_22583);
and U23386 (N_23386,N_21878,N_21699);
nand U23387 (N_23387,N_21637,N_22107);
and U23388 (N_23388,N_21736,N_21863);
nand U23389 (N_23389,N_22415,N_21747);
or U23390 (N_23390,N_21985,N_22243);
or U23391 (N_23391,N_21765,N_22657);
nor U23392 (N_23392,N_21654,N_21847);
or U23393 (N_23393,N_21980,N_21903);
and U23394 (N_23394,N_22577,N_21909);
nor U23395 (N_23395,N_21762,N_22518);
nor U23396 (N_23396,N_22181,N_22369);
or U23397 (N_23397,N_22026,N_22529);
nand U23398 (N_23398,N_22195,N_22767);
or U23399 (N_23399,N_22198,N_22210);
xnor U23400 (N_23400,N_21949,N_22441);
nor U23401 (N_23401,N_22518,N_22745);
or U23402 (N_23402,N_21887,N_22651);
xor U23403 (N_23403,N_22493,N_22035);
xnor U23404 (N_23404,N_22620,N_21729);
nor U23405 (N_23405,N_21893,N_22508);
nor U23406 (N_23406,N_22629,N_22171);
nand U23407 (N_23407,N_21978,N_22136);
and U23408 (N_23408,N_22400,N_22266);
and U23409 (N_23409,N_22756,N_21749);
xor U23410 (N_23410,N_21627,N_21945);
or U23411 (N_23411,N_21725,N_22114);
nand U23412 (N_23412,N_21851,N_22743);
or U23413 (N_23413,N_22769,N_21834);
or U23414 (N_23414,N_22326,N_22755);
nand U23415 (N_23415,N_22331,N_22141);
nand U23416 (N_23416,N_22015,N_21703);
and U23417 (N_23417,N_21696,N_22239);
nor U23418 (N_23418,N_22528,N_22334);
and U23419 (N_23419,N_22626,N_22671);
nand U23420 (N_23420,N_21826,N_22008);
and U23421 (N_23421,N_22674,N_22743);
nor U23422 (N_23422,N_22668,N_22657);
and U23423 (N_23423,N_22497,N_22344);
or U23424 (N_23424,N_21755,N_22745);
or U23425 (N_23425,N_21941,N_21945);
and U23426 (N_23426,N_22080,N_22020);
xor U23427 (N_23427,N_21793,N_21845);
nand U23428 (N_23428,N_21804,N_22534);
nand U23429 (N_23429,N_22348,N_22285);
and U23430 (N_23430,N_21688,N_22105);
xnor U23431 (N_23431,N_21753,N_22006);
and U23432 (N_23432,N_21714,N_21922);
xor U23433 (N_23433,N_22172,N_22205);
xor U23434 (N_23434,N_22742,N_22711);
nand U23435 (N_23435,N_21809,N_22444);
xnor U23436 (N_23436,N_22188,N_22485);
and U23437 (N_23437,N_21732,N_22709);
and U23438 (N_23438,N_22069,N_22214);
and U23439 (N_23439,N_22191,N_21851);
xor U23440 (N_23440,N_22687,N_22312);
or U23441 (N_23441,N_21607,N_22180);
nor U23442 (N_23442,N_21690,N_22223);
nand U23443 (N_23443,N_22507,N_22362);
nand U23444 (N_23444,N_22496,N_22511);
nand U23445 (N_23445,N_21734,N_21676);
or U23446 (N_23446,N_21752,N_21845);
nand U23447 (N_23447,N_21809,N_22438);
and U23448 (N_23448,N_22688,N_22549);
and U23449 (N_23449,N_21915,N_22267);
nor U23450 (N_23450,N_22713,N_22338);
and U23451 (N_23451,N_21705,N_22165);
nor U23452 (N_23452,N_21856,N_22061);
and U23453 (N_23453,N_22592,N_22498);
nand U23454 (N_23454,N_22499,N_21623);
or U23455 (N_23455,N_21686,N_21970);
nor U23456 (N_23456,N_22533,N_21733);
or U23457 (N_23457,N_21843,N_22557);
and U23458 (N_23458,N_22487,N_22292);
and U23459 (N_23459,N_22396,N_21814);
or U23460 (N_23460,N_22421,N_22578);
and U23461 (N_23461,N_21793,N_21780);
or U23462 (N_23462,N_22210,N_22378);
nand U23463 (N_23463,N_22502,N_22184);
nand U23464 (N_23464,N_22369,N_21875);
and U23465 (N_23465,N_22241,N_22363);
or U23466 (N_23466,N_21622,N_21884);
xnor U23467 (N_23467,N_22711,N_22540);
or U23468 (N_23468,N_21934,N_21728);
nand U23469 (N_23469,N_22107,N_21822);
nand U23470 (N_23470,N_22471,N_21940);
or U23471 (N_23471,N_21804,N_22121);
nand U23472 (N_23472,N_22124,N_22493);
xor U23473 (N_23473,N_22613,N_22172);
xor U23474 (N_23474,N_22536,N_22527);
and U23475 (N_23475,N_21752,N_21673);
nor U23476 (N_23476,N_22430,N_22013);
nor U23477 (N_23477,N_21718,N_22187);
and U23478 (N_23478,N_22797,N_22114);
nand U23479 (N_23479,N_22235,N_22715);
or U23480 (N_23480,N_22407,N_21721);
or U23481 (N_23481,N_21999,N_22792);
xor U23482 (N_23482,N_22663,N_21752);
or U23483 (N_23483,N_22010,N_22482);
xnor U23484 (N_23484,N_21914,N_21844);
xor U23485 (N_23485,N_22623,N_22706);
and U23486 (N_23486,N_22254,N_21737);
and U23487 (N_23487,N_21718,N_22582);
nor U23488 (N_23488,N_22539,N_22482);
nand U23489 (N_23489,N_22190,N_22198);
or U23490 (N_23490,N_22794,N_22056);
nand U23491 (N_23491,N_21667,N_21943);
and U23492 (N_23492,N_22543,N_22601);
and U23493 (N_23493,N_21820,N_22600);
xnor U23494 (N_23494,N_22158,N_22748);
nor U23495 (N_23495,N_22761,N_22053);
or U23496 (N_23496,N_22178,N_21794);
nor U23497 (N_23497,N_22093,N_22096);
nor U23498 (N_23498,N_22752,N_22109);
nor U23499 (N_23499,N_22080,N_22700);
nand U23500 (N_23500,N_22181,N_21919);
or U23501 (N_23501,N_21790,N_22583);
or U23502 (N_23502,N_21670,N_21647);
xnor U23503 (N_23503,N_22288,N_22565);
and U23504 (N_23504,N_22514,N_22323);
or U23505 (N_23505,N_22541,N_21992);
nand U23506 (N_23506,N_22239,N_21958);
or U23507 (N_23507,N_22655,N_22342);
xnor U23508 (N_23508,N_21706,N_21747);
or U23509 (N_23509,N_21889,N_22578);
nor U23510 (N_23510,N_22561,N_21668);
nor U23511 (N_23511,N_22732,N_22030);
nand U23512 (N_23512,N_22490,N_22642);
and U23513 (N_23513,N_21870,N_22570);
or U23514 (N_23514,N_22267,N_21856);
or U23515 (N_23515,N_22075,N_22099);
nand U23516 (N_23516,N_22464,N_22525);
nor U23517 (N_23517,N_21802,N_21962);
and U23518 (N_23518,N_22608,N_21645);
xnor U23519 (N_23519,N_21837,N_21631);
nand U23520 (N_23520,N_22780,N_22662);
or U23521 (N_23521,N_21910,N_22702);
or U23522 (N_23522,N_21771,N_21710);
or U23523 (N_23523,N_22577,N_22598);
nor U23524 (N_23524,N_21987,N_22268);
or U23525 (N_23525,N_22226,N_21771);
nand U23526 (N_23526,N_22454,N_22485);
nor U23527 (N_23527,N_22263,N_22382);
nor U23528 (N_23528,N_22484,N_21604);
and U23529 (N_23529,N_22757,N_21624);
nand U23530 (N_23530,N_22588,N_22331);
xnor U23531 (N_23531,N_22256,N_22071);
or U23532 (N_23532,N_22632,N_22262);
nand U23533 (N_23533,N_21713,N_22775);
xnor U23534 (N_23534,N_22675,N_22693);
and U23535 (N_23535,N_22731,N_21937);
xor U23536 (N_23536,N_21858,N_22135);
and U23537 (N_23537,N_21609,N_22092);
nor U23538 (N_23538,N_22687,N_22374);
xnor U23539 (N_23539,N_22047,N_22647);
nor U23540 (N_23540,N_21852,N_22567);
or U23541 (N_23541,N_22463,N_22508);
and U23542 (N_23542,N_22414,N_21748);
nand U23543 (N_23543,N_22187,N_22269);
nand U23544 (N_23544,N_22592,N_22573);
nor U23545 (N_23545,N_22105,N_22539);
xnor U23546 (N_23546,N_22757,N_22141);
or U23547 (N_23547,N_21936,N_22696);
nand U23548 (N_23548,N_22229,N_22204);
or U23549 (N_23549,N_22630,N_22380);
and U23550 (N_23550,N_22162,N_22799);
xor U23551 (N_23551,N_22520,N_22370);
xnor U23552 (N_23552,N_21899,N_21990);
and U23553 (N_23553,N_22193,N_22552);
nand U23554 (N_23554,N_22347,N_22239);
nor U23555 (N_23555,N_22342,N_22404);
or U23556 (N_23556,N_22769,N_22243);
xor U23557 (N_23557,N_21955,N_21697);
and U23558 (N_23558,N_22036,N_21763);
nand U23559 (N_23559,N_22039,N_22215);
or U23560 (N_23560,N_22733,N_22281);
nor U23561 (N_23561,N_22338,N_22681);
nor U23562 (N_23562,N_22573,N_22094);
xnor U23563 (N_23563,N_22350,N_22436);
or U23564 (N_23564,N_22663,N_22646);
nand U23565 (N_23565,N_21952,N_22715);
nor U23566 (N_23566,N_21696,N_22619);
and U23567 (N_23567,N_22333,N_21857);
and U23568 (N_23568,N_22764,N_21933);
nor U23569 (N_23569,N_21912,N_22687);
xnor U23570 (N_23570,N_22036,N_21812);
xor U23571 (N_23571,N_21931,N_21882);
and U23572 (N_23572,N_22095,N_21958);
nor U23573 (N_23573,N_22415,N_21898);
or U23574 (N_23574,N_22197,N_21687);
or U23575 (N_23575,N_22581,N_22306);
nor U23576 (N_23576,N_22763,N_22544);
xor U23577 (N_23577,N_22740,N_21681);
nor U23578 (N_23578,N_22717,N_22014);
nand U23579 (N_23579,N_22083,N_22536);
nand U23580 (N_23580,N_22719,N_21854);
xnor U23581 (N_23581,N_22405,N_22564);
xnor U23582 (N_23582,N_22686,N_21712);
xor U23583 (N_23583,N_21785,N_22237);
nand U23584 (N_23584,N_22570,N_22703);
nor U23585 (N_23585,N_22660,N_22103);
and U23586 (N_23586,N_22690,N_21707);
nand U23587 (N_23587,N_22556,N_21841);
nor U23588 (N_23588,N_21734,N_22340);
nor U23589 (N_23589,N_21787,N_22032);
nor U23590 (N_23590,N_22753,N_22015);
or U23591 (N_23591,N_22571,N_21758);
or U23592 (N_23592,N_21755,N_22381);
and U23593 (N_23593,N_22742,N_22282);
or U23594 (N_23594,N_22013,N_22600);
nor U23595 (N_23595,N_21962,N_21672);
nand U23596 (N_23596,N_21915,N_22069);
or U23597 (N_23597,N_22602,N_22734);
xnor U23598 (N_23598,N_22160,N_21666);
nand U23599 (N_23599,N_22047,N_22600);
nand U23600 (N_23600,N_21977,N_22658);
or U23601 (N_23601,N_22094,N_21666);
or U23602 (N_23602,N_22670,N_21982);
nand U23603 (N_23603,N_22228,N_21763);
nand U23604 (N_23604,N_22087,N_22151);
xor U23605 (N_23605,N_21942,N_21605);
xnor U23606 (N_23606,N_21726,N_22667);
nor U23607 (N_23607,N_21669,N_21991);
and U23608 (N_23608,N_22300,N_22526);
xor U23609 (N_23609,N_22315,N_21784);
nor U23610 (N_23610,N_22064,N_22602);
nor U23611 (N_23611,N_21915,N_21665);
nand U23612 (N_23612,N_22446,N_22726);
and U23613 (N_23613,N_22339,N_21825);
nor U23614 (N_23614,N_21652,N_21702);
xor U23615 (N_23615,N_22422,N_22399);
nor U23616 (N_23616,N_21676,N_21602);
and U23617 (N_23617,N_22288,N_22263);
nand U23618 (N_23618,N_21876,N_22729);
nor U23619 (N_23619,N_22683,N_22319);
nand U23620 (N_23620,N_21981,N_21930);
and U23621 (N_23621,N_22098,N_22043);
and U23622 (N_23622,N_22147,N_21609);
or U23623 (N_23623,N_21999,N_21838);
and U23624 (N_23624,N_21613,N_22452);
xor U23625 (N_23625,N_22485,N_22588);
and U23626 (N_23626,N_22064,N_21932);
nand U23627 (N_23627,N_21661,N_22792);
nand U23628 (N_23628,N_22410,N_22174);
and U23629 (N_23629,N_22042,N_22345);
xnor U23630 (N_23630,N_22128,N_22147);
or U23631 (N_23631,N_22255,N_21638);
nor U23632 (N_23632,N_22294,N_22462);
nand U23633 (N_23633,N_22748,N_22250);
xnor U23634 (N_23634,N_22377,N_22694);
nand U23635 (N_23635,N_21710,N_22536);
or U23636 (N_23636,N_21660,N_21711);
nand U23637 (N_23637,N_22298,N_22660);
or U23638 (N_23638,N_22504,N_22623);
nand U23639 (N_23639,N_22019,N_22544);
nand U23640 (N_23640,N_22315,N_21712);
nand U23641 (N_23641,N_22065,N_22686);
and U23642 (N_23642,N_22425,N_21618);
or U23643 (N_23643,N_22444,N_21921);
nor U23644 (N_23644,N_22596,N_22397);
nand U23645 (N_23645,N_21651,N_21919);
xnor U23646 (N_23646,N_22673,N_22419);
nor U23647 (N_23647,N_22702,N_22021);
nand U23648 (N_23648,N_22634,N_21871);
and U23649 (N_23649,N_22057,N_22394);
nor U23650 (N_23650,N_21916,N_22075);
or U23651 (N_23651,N_22771,N_22724);
and U23652 (N_23652,N_22500,N_22407);
or U23653 (N_23653,N_22336,N_22286);
or U23654 (N_23654,N_22313,N_21862);
and U23655 (N_23655,N_22651,N_21668);
nand U23656 (N_23656,N_22462,N_22777);
xnor U23657 (N_23657,N_22108,N_21950);
or U23658 (N_23658,N_22133,N_21935);
and U23659 (N_23659,N_22096,N_22658);
and U23660 (N_23660,N_21770,N_22073);
xnor U23661 (N_23661,N_21781,N_22040);
nor U23662 (N_23662,N_21884,N_22390);
or U23663 (N_23663,N_22377,N_21757);
and U23664 (N_23664,N_22777,N_22400);
or U23665 (N_23665,N_22661,N_22397);
and U23666 (N_23666,N_22605,N_21844);
and U23667 (N_23667,N_22333,N_22043);
and U23668 (N_23668,N_21624,N_22711);
or U23669 (N_23669,N_22263,N_21740);
or U23670 (N_23670,N_21778,N_22474);
xnor U23671 (N_23671,N_22053,N_21714);
nand U23672 (N_23672,N_22488,N_21799);
or U23673 (N_23673,N_21699,N_21970);
and U23674 (N_23674,N_22695,N_22670);
nand U23675 (N_23675,N_22411,N_22148);
nor U23676 (N_23676,N_21683,N_22618);
or U23677 (N_23677,N_21972,N_22085);
xnor U23678 (N_23678,N_21709,N_21991);
and U23679 (N_23679,N_21956,N_22572);
xor U23680 (N_23680,N_22180,N_22472);
nand U23681 (N_23681,N_22108,N_21951);
or U23682 (N_23682,N_22038,N_22104);
or U23683 (N_23683,N_21953,N_21986);
nor U23684 (N_23684,N_21671,N_22000);
nand U23685 (N_23685,N_22779,N_21772);
nand U23686 (N_23686,N_21979,N_22644);
xnor U23687 (N_23687,N_22502,N_21641);
and U23688 (N_23688,N_21921,N_22017);
or U23689 (N_23689,N_22794,N_22391);
xnor U23690 (N_23690,N_22168,N_21940);
xor U23691 (N_23691,N_22332,N_21986);
or U23692 (N_23692,N_21786,N_21728);
or U23693 (N_23693,N_22399,N_21914);
xor U23694 (N_23694,N_21933,N_21986);
xnor U23695 (N_23695,N_21869,N_22315);
nand U23696 (N_23696,N_22293,N_21999);
and U23697 (N_23697,N_22226,N_22380);
nor U23698 (N_23698,N_22623,N_21623);
nor U23699 (N_23699,N_21721,N_22314);
or U23700 (N_23700,N_22644,N_22069);
and U23701 (N_23701,N_22651,N_21647);
or U23702 (N_23702,N_22499,N_21960);
and U23703 (N_23703,N_22317,N_21951);
nor U23704 (N_23704,N_21766,N_22080);
nand U23705 (N_23705,N_22721,N_21985);
xnor U23706 (N_23706,N_21904,N_22720);
and U23707 (N_23707,N_22515,N_22379);
nor U23708 (N_23708,N_22001,N_22073);
xnor U23709 (N_23709,N_21713,N_22795);
nor U23710 (N_23710,N_21696,N_22343);
and U23711 (N_23711,N_21778,N_22111);
and U23712 (N_23712,N_22149,N_22377);
and U23713 (N_23713,N_21794,N_22037);
or U23714 (N_23714,N_21634,N_22160);
or U23715 (N_23715,N_22222,N_22368);
nand U23716 (N_23716,N_22155,N_22338);
xor U23717 (N_23717,N_22053,N_22721);
and U23718 (N_23718,N_21667,N_22325);
nand U23719 (N_23719,N_22031,N_22018);
xnor U23720 (N_23720,N_22670,N_22656);
nand U23721 (N_23721,N_22608,N_21840);
and U23722 (N_23722,N_22728,N_22333);
or U23723 (N_23723,N_22343,N_21963);
or U23724 (N_23724,N_22719,N_22430);
nor U23725 (N_23725,N_22378,N_21959);
and U23726 (N_23726,N_21816,N_22729);
xor U23727 (N_23727,N_22342,N_21849);
nor U23728 (N_23728,N_22125,N_22563);
nand U23729 (N_23729,N_22065,N_21733);
and U23730 (N_23730,N_21895,N_22515);
xor U23731 (N_23731,N_22422,N_22630);
xor U23732 (N_23732,N_22584,N_22459);
and U23733 (N_23733,N_22011,N_21794);
nor U23734 (N_23734,N_22542,N_21709);
nand U23735 (N_23735,N_22275,N_22767);
xor U23736 (N_23736,N_22787,N_21843);
or U23737 (N_23737,N_21628,N_21708);
nand U23738 (N_23738,N_21985,N_21816);
xnor U23739 (N_23739,N_22087,N_22300);
nor U23740 (N_23740,N_21883,N_22447);
or U23741 (N_23741,N_22356,N_22257);
or U23742 (N_23742,N_21696,N_22307);
nor U23743 (N_23743,N_22528,N_21820);
nor U23744 (N_23744,N_22796,N_22438);
nor U23745 (N_23745,N_22663,N_21964);
nor U23746 (N_23746,N_22527,N_22440);
or U23747 (N_23747,N_22514,N_22385);
or U23748 (N_23748,N_21860,N_22025);
and U23749 (N_23749,N_22737,N_22066);
and U23750 (N_23750,N_21655,N_22189);
xor U23751 (N_23751,N_21951,N_22756);
or U23752 (N_23752,N_21977,N_22538);
nor U23753 (N_23753,N_22315,N_22455);
nand U23754 (N_23754,N_22295,N_22072);
nor U23755 (N_23755,N_22711,N_22741);
xnor U23756 (N_23756,N_22301,N_21866);
nand U23757 (N_23757,N_21795,N_21712);
xnor U23758 (N_23758,N_21632,N_21997);
nand U23759 (N_23759,N_22516,N_22046);
nand U23760 (N_23760,N_22531,N_22060);
nor U23761 (N_23761,N_22283,N_22390);
and U23762 (N_23762,N_21875,N_21886);
or U23763 (N_23763,N_22598,N_22736);
and U23764 (N_23764,N_22103,N_22295);
or U23765 (N_23765,N_22608,N_22188);
or U23766 (N_23766,N_21991,N_22404);
xor U23767 (N_23767,N_22581,N_21942);
nor U23768 (N_23768,N_22141,N_21853);
or U23769 (N_23769,N_21740,N_22070);
and U23770 (N_23770,N_21711,N_22764);
or U23771 (N_23771,N_22432,N_22353);
xnor U23772 (N_23772,N_21862,N_22509);
nor U23773 (N_23773,N_22179,N_22485);
or U23774 (N_23774,N_21969,N_22570);
nand U23775 (N_23775,N_21701,N_22363);
or U23776 (N_23776,N_22227,N_22007);
or U23777 (N_23777,N_21800,N_22586);
nor U23778 (N_23778,N_21631,N_22256);
xnor U23779 (N_23779,N_21949,N_22159);
xor U23780 (N_23780,N_22198,N_22186);
xnor U23781 (N_23781,N_22708,N_22069);
xnor U23782 (N_23782,N_22455,N_22136);
nand U23783 (N_23783,N_22171,N_21825);
xnor U23784 (N_23784,N_21762,N_21926);
or U23785 (N_23785,N_21986,N_22772);
nand U23786 (N_23786,N_22392,N_22396);
and U23787 (N_23787,N_22518,N_21908);
xnor U23788 (N_23788,N_22762,N_22630);
xor U23789 (N_23789,N_22235,N_22129);
nand U23790 (N_23790,N_22515,N_22431);
nand U23791 (N_23791,N_22202,N_21664);
nand U23792 (N_23792,N_21698,N_22646);
xnor U23793 (N_23793,N_21904,N_21758);
nor U23794 (N_23794,N_22241,N_21802);
or U23795 (N_23795,N_21732,N_22786);
xnor U23796 (N_23796,N_22760,N_22030);
and U23797 (N_23797,N_22461,N_21604);
nand U23798 (N_23798,N_21740,N_22359);
or U23799 (N_23799,N_22258,N_22235);
nor U23800 (N_23800,N_22753,N_22166);
nor U23801 (N_23801,N_21899,N_22021);
or U23802 (N_23802,N_21731,N_21711);
and U23803 (N_23803,N_22532,N_22362);
xnor U23804 (N_23804,N_22376,N_21779);
or U23805 (N_23805,N_22595,N_22029);
xor U23806 (N_23806,N_22261,N_21802);
or U23807 (N_23807,N_22623,N_22269);
nor U23808 (N_23808,N_22343,N_22035);
nor U23809 (N_23809,N_21871,N_21818);
or U23810 (N_23810,N_21950,N_22596);
nand U23811 (N_23811,N_22326,N_21692);
xnor U23812 (N_23812,N_22433,N_21603);
xor U23813 (N_23813,N_21739,N_22694);
xnor U23814 (N_23814,N_22372,N_22497);
nand U23815 (N_23815,N_21736,N_22402);
nor U23816 (N_23816,N_22019,N_21929);
xor U23817 (N_23817,N_22157,N_21739);
xnor U23818 (N_23818,N_22680,N_21679);
nor U23819 (N_23819,N_22276,N_22386);
and U23820 (N_23820,N_22310,N_22488);
or U23821 (N_23821,N_22027,N_22227);
xnor U23822 (N_23822,N_22001,N_22311);
nand U23823 (N_23823,N_22668,N_22633);
or U23824 (N_23824,N_21828,N_22433);
and U23825 (N_23825,N_21823,N_22368);
nand U23826 (N_23826,N_22694,N_21711);
nor U23827 (N_23827,N_21635,N_22690);
nand U23828 (N_23828,N_22091,N_21687);
or U23829 (N_23829,N_22237,N_22783);
nand U23830 (N_23830,N_22080,N_22245);
xor U23831 (N_23831,N_22617,N_22544);
xor U23832 (N_23832,N_22783,N_21685);
or U23833 (N_23833,N_22792,N_22361);
nand U23834 (N_23834,N_21723,N_22530);
xor U23835 (N_23835,N_22589,N_22322);
or U23836 (N_23836,N_21707,N_22326);
nand U23837 (N_23837,N_22567,N_21759);
and U23838 (N_23838,N_21797,N_22342);
nand U23839 (N_23839,N_21860,N_21609);
nand U23840 (N_23840,N_22602,N_21790);
or U23841 (N_23841,N_22241,N_22338);
xor U23842 (N_23842,N_21889,N_22289);
xor U23843 (N_23843,N_22382,N_21716);
xnor U23844 (N_23844,N_22370,N_22245);
and U23845 (N_23845,N_21856,N_22793);
nor U23846 (N_23846,N_21730,N_22379);
and U23847 (N_23847,N_22070,N_22642);
or U23848 (N_23848,N_22122,N_21629);
xnor U23849 (N_23849,N_22216,N_21790);
nand U23850 (N_23850,N_21605,N_22355);
nor U23851 (N_23851,N_21663,N_21954);
or U23852 (N_23852,N_21716,N_22166);
xnor U23853 (N_23853,N_22617,N_21754);
nor U23854 (N_23854,N_21750,N_22733);
xnor U23855 (N_23855,N_21831,N_21890);
xor U23856 (N_23856,N_22442,N_21824);
nor U23857 (N_23857,N_21770,N_22634);
or U23858 (N_23858,N_22617,N_22005);
nor U23859 (N_23859,N_21924,N_22596);
nand U23860 (N_23860,N_21812,N_21655);
nand U23861 (N_23861,N_22336,N_21890);
or U23862 (N_23862,N_22635,N_22164);
or U23863 (N_23863,N_21929,N_22279);
xor U23864 (N_23864,N_22553,N_22241);
nand U23865 (N_23865,N_21745,N_22483);
nand U23866 (N_23866,N_22729,N_22623);
xor U23867 (N_23867,N_21754,N_22342);
or U23868 (N_23868,N_21744,N_21942);
nor U23869 (N_23869,N_22018,N_21739);
xor U23870 (N_23870,N_22405,N_21998);
nor U23871 (N_23871,N_21827,N_22192);
and U23872 (N_23872,N_21907,N_22105);
nor U23873 (N_23873,N_22096,N_22423);
nand U23874 (N_23874,N_21863,N_21985);
or U23875 (N_23875,N_22420,N_22590);
nor U23876 (N_23876,N_21778,N_22677);
xnor U23877 (N_23877,N_21985,N_22295);
xor U23878 (N_23878,N_21711,N_21812);
or U23879 (N_23879,N_22018,N_21892);
xnor U23880 (N_23880,N_21952,N_22154);
nand U23881 (N_23881,N_22286,N_22533);
xnor U23882 (N_23882,N_22394,N_22016);
nand U23883 (N_23883,N_22641,N_21951);
xnor U23884 (N_23884,N_22238,N_22792);
nor U23885 (N_23885,N_22559,N_22603);
nor U23886 (N_23886,N_22569,N_21862);
nor U23887 (N_23887,N_21802,N_22347);
xnor U23888 (N_23888,N_22564,N_22470);
and U23889 (N_23889,N_22191,N_22695);
and U23890 (N_23890,N_22752,N_22635);
and U23891 (N_23891,N_22228,N_22112);
and U23892 (N_23892,N_22530,N_21905);
nand U23893 (N_23893,N_22029,N_22658);
or U23894 (N_23894,N_22732,N_22379);
or U23895 (N_23895,N_22735,N_22330);
and U23896 (N_23896,N_22624,N_22391);
or U23897 (N_23897,N_21961,N_22790);
and U23898 (N_23898,N_21934,N_22768);
nand U23899 (N_23899,N_22146,N_21842);
xnor U23900 (N_23900,N_22633,N_22512);
nor U23901 (N_23901,N_22519,N_21992);
xor U23902 (N_23902,N_22117,N_22508);
nor U23903 (N_23903,N_22290,N_22267);
and U23904 (N_23904,N_22530,N_22282);
nor U23905 (N_23905,N_21818,N_22786);
nor U23906 (N_23906,N_21845,N_22793);
nand U23907 (N_23907,N_22611,N_22624);
nand U23908 (N_23908,N_22280,N_22504);
and U23909 (N_23909,N_21758,N_22527);
or U23910 (N_23910,N_22257,N_22797);
xnor U23911 (N_23911,N_21670,N_22732);
nand U23912 (N_23912,N_22684,N_22760);
and U23913 (N_23913,N_21622,N_21797);
or U23914 (N_23914,N_22275,N_22617);
and U23915 (N_23915,N_22171,N_22723);
or U23916 (N_23916,N_22367,N_22429);
or U23917 (N_23917,N_22391,N_22225);
nor U23918 (N_23918,N_22547,N_22359);
nand U23919 (N_23919,N_22265,N_22403);
nor U23920 (N_23920,N_22448,N_21670);
or U23921 (N_23921,N_21931,N_21947);
nand U23922 (N_23922,N_22609,N_22530);
nand U23923 (N_23923,N_22795,N_21751);
nand U23924 (N_23924,N_22528,N_22055);
and U23925 (N_23925,N_22284,N_22541);
and U23926 (N_23926,N_22200,N_22739);
or U23927 (N_23927,N_22740,N_22245);
nand U23928 (N_23928,N_21628,N_22724);
and U23929 (N_23929,N_22613,N_22227);
nand U23930 (N_23930,N_21862,N_22221);
xnor U23931 (N_23931,N_22253,N_22148);
xor U23932 (N_23932,N_22046,N_22055);
or U23933 (N_23933,N_22199,N_22051);
nor U23934 (N_23934,N_22007,N_22218);
or U23935 (N_23935,N_21888,N_22307);
or U23936 (N_23936,N_22457,N_21864);
nor U23937 (N_23937,N_21658,N_22175);
nor U23938 (N_23938,N_21891,N_21975);
or U23939 (N_23939,N_21731,N_21881);
nor U23940 (N_23940,N_22267,N_22701);
or U23941 (N_23941,N_22157,N_22359);
and U23942 (N_23942,N_21848,N_22587);
or U23943 (N_23943,N_22517,N_22235);
or U23944 (N_23944,N_22577,N_22466);
or U23945 (N_23945,N_22126,N_21959);
xnor U23946 (N_23946,N_21808,N_22251);
xnor U23947 (N_23947,N_21972,N_22319);
nor U23948 (N_23948,N_22323,N_22050);
nor U23949 (N_23949,N_22796,N_22576);
nand U23950 (N_23950,N_22299,N_22270);
or U23951 (N_23951,N_22187,N_22312);
xor U23952 (N_23952,N_21986,N_21678);
nor U23953 (N_23953,N_22617,N_22585);
and U23954 (N_23954,N_22301,N_21832);
and U23955 (N_23955,N_22155,N_22328);
xnor U23956 (N_23956,N_22109,N_22261);
or U23957 (N_23957,N_21716,N_22234);
or U23958 (N_23958,N_22436,N_22271);
xor U23959 (N_23959,N_22632,N_22737);
or U23960 (N_23960,N_22433,N_22028);
and U23961 (N_23961,N_21823,N_21677);
or U23962 (N_23962,N_22340,N_22391);
nand U23963 (N_23963,N_22357,N_22499);
or U23964 (N_23964,N_21724,N_22056);
nor U23965 (N_23965,N_22285,N_22168);
nor U23966 (N_23966,N_22439,N_22677);
nor U23967 (N_23967,N_22430,N_21927);
and U23968 (N_23968,N_22610,N_21926);
nand U23969 (N_23969,N_21854,N_22306);
nor U23970 (N_23970,N_21680,N_22743);
or U23971 (N_23971,N_22311,N_22186);
and U23972 (N_23972,N_22547,N_21680);
nand U23973 (N_23973,N_22047,N_22159);
xnor U23974 (N_23974,N_22699,N_21946);
or U23975 (N_23975,N_22552,N_22315);
nor U23976 (N_23976,N_22264,N_21613);
nor U23977 (N_23977,N_21702,N_21832);
and U23978 (N_23978,N_22494,N_22033);
nand U23979 (N_23979,N_21602,N_22552);
nor U23980 (N_23980,N_22269,N_22231);
nor U23981 (N_23981,N_21821,N_21745);
or U23982 (N_23982,N_21699,N_22285);
or U23983 (N_23983,N_22575,N_22031);
nor U23984 (N_23984,N_22328,N_22344);
nand U23985 (N_23985,N_22445,N_22088);
nand U23986 (N_23986,N_22404,N_21828);
and U23987 (N_23987,N_22718,N_21669);
nor U23988 (N_23988,N_22039,N_22247);
and U23989 (N_23989,N_22513,N_22405);
nor U23990 (N_23990,N_22685,N_21789);
or U23991 (N_23991,N_22205,N_22474);
and U23992 (N_23992,N_22514,N_21688);
or U23993 (N_23993,N_22483,N_22173);
nand U23994 (N_23994,N_22413,N_22766);
xor U23995 (N_23995,N_21857,N_22070);
xor U23996 (N_23996,N_22362,N_22633);
nor U23997 (N_23997,N_22087,N_21687);
nor U23998 (N_23998,N_22794,N_22692);
nand U23999 (N_23999,N_22113,N_21600);
and U24000 (N_24000,N_23640,N_23958);
nor U24001 (N_24001,N_23292,N_23672);
nor U24002 (N_24002,N_23616,N_23871);
xor U24003 (N_24003,N_23595,N_23645);
and U24004 (N_24004,N_22840,N_23873);
xor U24005 (N_24005,N_22977,N_23074);
xnor U24006 (N_24006,N_23164,N_23160);
nand U24007 (N_24007,N_23850,N_23932);
nand U24008 (N_24008,N_23085,N_23834);
xnor U24009 (N_24009,N_23100,N_23108);
xor U24010 (N_24010,N_23131,N_23297);
xor U24011 (N_24011,N_23156,N_23760);
nor U24012 (N_24012,N_23343,N_22836);
nor U24013 (N_24013,N_23321,N_23878);
or U24014 (N_24014,N_22981,N_23233);
nor U24015 (N_24015,N_22829,N_23408);
or U24016 (N_24016,N_23307,N_23094);
nor U24017 (N_24017,N_23203,N_23554);
nand U24018 (N_24018,N_23263,N_22884);
and U24019 (N_24019,N_23064,N_22983);
xor U24020 (N_24020,N_23116,N_23114);
or U24021 (N_24021,N_23334,N_23308);
xnor U24022 (N_24022,N_23994,N_22864);
nand U24023 (N_24023,N_23257,N_22990);
nor U24024 (N_24024,N_23588,N_23712);
xor U24025 (N_24025,N_23806,N_23232);
nand U24026 (N_24026,N_23681,N_23522);
or U24027 (N_24027,N_22926,N_23811);
nor U24028 (N_24028,N_23813,N_23080);
nor U24029 (N_24029,N_23193,N_23793);
xor U24030 (N_24030,N_23048,N_23599);
or U24031 (N_24031,N_23832,N_23743);
or U24032 (N_24032,N_23722,N_23728);
or U24033 (N_24033,N_23779,N_23853);
and U24034 (N_24034,N_22949,N_22959);
nand U24035 (N_24035,N_23208,N_23837);
nor U24036 (N_24036,N_23367,N_22814);
or U24037 (N_24037,N_23059,N_23194);
xor U24038 (N_24038,N_22890,N_22966);
nand U24039 (N_24039,N_23130,N_23610);
nand U24040 (N_24040,N_23823,N_23955);
or U24041 (N_24041,N_23357,N_22872);
xnor U24042 (N_24042,N_22995,N_23521);
nand U24043 (N_24043,N_23763,N_22916);
and U24044 (N_24044,N_23010,N_23315);
nor U24045 (N_24045,N_23364,N_23920);
nor U24046 (N_24046,N_23634,N_22954);
nor U24047 (N_24047,N_23851,N_22936);
xor U24048 (N_24048,N_23002,N_23272);
or U24049 (N_24049,N_22904,N_23846);
nor U24050 (N_24050,N_23584,N_23504);
or U24051 (N_24051,N_23035,N_23692);
nor U24052 (N_24052,N_23173,N_23426);
nor U24053 (N_24053,N_23065,N_23559);
nand U24054 (N_24054,N_23799,N_23106);
nor U24055 (N_24055,N_22964,N_23686);
xnor U24056 (N_24056,N_23467,N_22928);
or U24057 (N_24057,N_22824,N_23548);
xor U24058 (N_24058,N_23754,N_23387);
and U24059 (N_24059,N_23933,N_22871);
nand U24060 (N_24060,N_22813,N_23583);
nor U24061 (N_24061,N_23298,N_23586);
nand U24062 (N_24062,N_22897,N_22997);
nand U24063 (N_24063,N_23344,N_22933);
and U24064 (N_24064,N_23733,N_23455);
nor U24065 (N_24065,N_22886,N_23024);
nor U24066 (N_24066,N_22901,N_23135);
nor U24067 (N_24067,N_23903,N_23775);
xnor U24068 (N_24068,N_23565,N_23628);
nor U24069 (N_24069,N_23975,N_22988);
or U24070 (N_24070,N_23786,N_23183);
nor U24071 (N_24071,N_22856,N_23673);
nand U24072 (N_24072,N_23355,N_23789);
or U24073 (N_24073,N_23362,N_23037);
xnor U24074 (N_24074,N_23503,N_23757);
nand U24075 (N_24075,N_23539,N_23657);
xnor U24076 (N_24076,N_23600,N_23350);
or U24077 (N_24077,N_23711,N_22918);
nor U24078 (N_24078,N_23568,N_22908);
or U24079 (N_24079,N_23047,N_23907);
and U24080 (N_24080,N_23354,N_22939);
nand U24081 (N_24081,N_23258,N_22946);
and U24082 (N_24082,N_23166,N_23524);
and U24083 (N_24083,N_23397,N_23454);
and U24084 (N_24084,N_23378,N_23824);
nor U24085 (N_24085,N_23324,N_23801);
nand U24086 (N_24086,N_23674,N_23865);
nor U24087 (N_24087,N_23732,N_23566);
nand U24088 (N_24088,N_23778,N_23854);
xnor U24089 (N_24089,N_23874,N_23316);
and U24090 (N_24090,N_22931,N_23279);
xnor U24091 (N_24091,N_23146,N_23076);
nor U24092 (N_24092,N_23236,N_23300);
xnor U24093 (N_24093,N_22878,N_23159);
and U24094 (N_24094,N_23015,N_23511);
and U24095 (N_24095,N_23639,N_23137);
and U24096 (N_24096,N_23613,N_23946);
xor U24097 (N_24097,N_23147,N_23912);
nor U24098 (N_24098,N_23444,N_22861);
nand U24099 (N_24099,N_23162,N_22980);
nand U24100 (N_24100,N_23723,N_23480);
and U24101 (N_24101,N_22852,N_22903);
nand U24102 (N_24102,N_23424,N_22960);
nand U24103 (N_24103,N_23005,N_23758);
nand U24104 (N_24104,N_22827,N_23677);
nand U24105 (N_24105,N_23215,N_22831);
and U24106 (N_24106,N_23935,N_22888);
or U24107 (N_24107,N_23301,N_23211);
xor U24108 (N_24108,N_23451,N_23384);
nand U24109 (N_24109,N_23704,N_23143);
nand U24110 (N_24110,N_23688,N_23109);
nor U24111 (N_24111,N_23859,N_23916);
or U24112 (N_24112,N_23585,N_22867);
and U24113 (N_24113,N_23663,N_23111);
or U24114 (N_24114,N_23502,N_22837);
and U24115 (N_24115,N_23520,N_23073);
and U24116 (N_24116,N_22819,N_23881);
or U24117 (N_24117,N_23171,N_23242);
nand U24118 (N_24118,N_22889,N_22943);
or U24119 (N_24119,N_23908,N_23306);
nor U24120 (N_24120,N_23372,N_23371);
and U24121 (N_24121,N_23345,N_23581);
xor U24122 (N_24122,N_23549,N_22893);
xnor U24123 (N_24123,N_23626,N_23910);
or U24124 (N_24124,N_23656,N_23918);
or U24125 (N_24125,N_23134,N_23883);
and U24126 (N_24126,N_23369,N_23980);
xor U24127 (N_24127,N_23181,N_23996);
nand U24128 (N_24128,N_23814,N_23529);
and U24129 (N_24129,N_23478,N_23057);
nand U24130 (N_24130,N_22941,N_23133);
nand U24131 (N_24131,N_23995,N_23552);
nor U24132 (N_24132,N_22838,N_23984);
nand U24133 (N_24133,N_23738,N_23553);
or U24134 (N_24134,N_23497,N_23598);
nor U24135 (N_24135,N_23070,N_23273);
nand U24136 (N_24136,N_23465,N_23101);
and U24137 (N_24137,N_23311,N_23039);
nor U24138 (N_24138,N_23981,N_23287);
nand U24139 (N_24139,N_22935,N_23031);
xor U24140 (N_24140,N_23151,N_23400);
nor U24141 (N_24141,N_23185,N_23468);
nand U24142 (N_24142,N_23170,N_23014);
xnor U24143 (N_24143,N_23830,N_23685);
or U24144 (N_24144,N_22880,N_23937);
nand U24145 (N_24145,N_23964,N_23642);
or U24146 (N_24146,N_22951,N_23180);
nor U24147 (N_24147,N_23612,N_23796);
xor U24148 (N_24148,N_22968,N_23774);
xor U24149 (N_24149,N_23827,N_23155);
and U24150 (N_24150,N_23188,N_23620);
nand U24151 (N_24151,N_22821,N_23911);
nand U24152 (N_24152,N_22967,N_23093);
and U24153 (N_24153,N_22952,N_23800);
xnor U24154 (N_24154,N_23337,N_23127);
or U24155 (N_24155,N_23041,N_23317);
nand U24156 (N_24156,N_23228,N_23973);
or U24157 (N_24157,N_23962,N_23264);
and U24158 (N_24158,N_23421,N_23636);
nand U24159 (N_24159,N_23154,N_23060);
xor U24160 (N_24160,N_23680,N_23373);
or U24161 (N_24161,N_23082,N_23998);
nor U24162 (N_24162,N_23144,N_22934);
xnor U24163 (N_24163,N_22874,N_22921);
or U24164 (N_24164,N_22866,N_23709);
nor U24165 (N_24165,N_22991,N_23516);
nand U24166 (N_24166,N_23990,N_23420);
nor U24167 (N_24167,N_23847,N_23915);
or U24168 (N_24168,N_23449,N_23152);
and U24169 (N_24169,N_23744,N_23826);
and U24170 (N_24170,N_23785,N_23679);
and U24171 (N_24171,N_23756,N_23036);
nor U24172 (N_24172,N_23312,N_23466);
and U24173 (N_24173,N_22812,N_23508);
xnor U24174 (N_24174,N_23238,N_23992);
nand U24175 (N_24175,N_23158,N_23077);
and U24176 (N_24176,N_22854,N_23071);
nand U24177 (N_24177,N_23967,N_22932);
nor U24178 (N_24178,N_23719,N_23835);
or U24179 (N_24179,N_23459,N_23447);
nand U24180 (N_24180,N_23771,N_23296);
xor U24181 (N_24181,N_23410,N_23021);
nor U24182 (N_24182,N_23087,N_22850);
xnor U24183 (N_24183,N_23470,N_23752);
nand U24184 (N_24184,N_23107,N_23831);
xnor U24185 (N_24185,N_22863,N_23987);
nand U24186 (N_24186,N_23435,N_23249);
and U24187 (N_24187,N_23028,N_23366);
xnor U24188 (N_24188,N_23533,N_23291);
xnor U24189 (N_24189,N_23913,N_23944);
nor U24190 (N_24190,N_23286,N_23671);
nand U24191 (N_24191,N_22800,N_22809);
xor U24192 (N_24192,N_23360,N_23842);
or U24193 (N_24193,N_23545,N_22815);
or U24194 (N_24194,N_23525,N_23033);
nor U24195 (N_24195,N_23901,N_22999);
xor U24196 (N_24196,N_23690,N_23977);
nand U24197 (N_24197,N_23968,N_23319);
and U24198 (N_24198,N_23490,N_22896);
nand U24199 (N_24199,N_23187,N_23798);
nor U24200 (N_24200,N_23611,N_23948);
xor U24201 (N_24201,N_22975,N_23498);
nor U24202 (N_24202,N_23112,N_23083);
xor U24203 (N_24203,N_23304,N_23848);
or U24204 (N_24204,N_23284,N_23969);
or U24205 (N_24205,N_23575,N_23833);
or U24206 (N_24206,N_22826,N_23906);
and U24207 (N_24207,N_23807,N_22868);
and U24208 (N_24208,N_23177,N_22883);
xor U24209 (N_24209,N_23066,N_23416);
nor U24210 (N_24210,N_23501,N_22876);
xor U24211 (N_24211,N_22998,N_22974);
nor U24212 (N_24212,N_23392,N_23804);
xnor U24213 (N_24213,N_23641,N_23541);
nand U24214 (N_24214,N_23358,N_23528);
nand U24215 (N_24215,N_23245,N_23638);
and U24216 (N_24216,N_23186,N_23515);
nor U24217 (N_24217,N_23042,N_22845);
nand U24218 (N_24218,N_23463,N_23044);
and U24219 (N_24219,N_23412,N_23687);
nand U24220 (N_24220,N_23658,N_23052);
xnor U24221 (N_24221,N_23009,N_23700);
nand U24222 (N_24222,N_23067,N_23457);
xnor U24223 (N_24223,N_23894,N_23182);
and U24224 (N_24224,N_23787,N_23550);
nand U24225 (N_24225,N_23691,N_23406);
and U24226 (N_24226,N_23934,N_22963);
or U24227 (N_24227,N_23736,N_23885);
nor U24228 (N_24228,N_23381,N_22839);
or U24229 (N_24229,N_23202,N_23303);
or U24230 (N_24230,N_23051,N_23239);
and U24231 (N_24231,N_23790,N_22920);
and U24232 (N_24232,N_23900,N_23828);
or U24233 (N_24233,N_23606,N_23684);
xor U24234 (N_24234,N_23999,N_22816);
nand U24235 (N_24235,N_23570,N_23072);
nor U24236 (N_24236,N_23056,N_23621);
and U24237 (N_24237,N_23049,N_23241);
and U24238 (N_24238,N_23902,N_22873);
nand U24239 (N_24239,N_23841,N_23678);
xnor U24240 (N_24240,N_23172,N_23812);
or U24241 (N_24241,N_23212,N_23061);
nor U24242 (N_24242,N_22808,N_23485);
xor U24243 (N_24243,N_23689,N_23759);
and U24244 (N_24244,N_23414,N_23329);
nor U24245 (N_24245,N_23008,N_23267);
xnor U24246 (N_24246,N_23727,N_23513);
or U24247 (N_24247,N_23394,N_23276);
or U24248 (N_24248,N_23479,N_23805);
and U24249 (N_24249,N_23573,N_23011);
xnor U24250 (N_24250,N_23949,N_22911);
nor U24251 (N_24251,N_23305,N_23320);
and U24252 (N_24252,N_23322,N_22848);
or U24253 (N_24253,N_23555,N_23310);
nor U24254 (N_24254,N_23735,N_23278);
xor U24255 (N_24255,N_23510,N_23484);
or U24256 (N_24256,N_23708,N_23268);
nor U24257 (N_24257,N_23572,N_23880);
or U24258 (N_24258,N_22942,N_23930);
nand U24259 (N_24259,N_23262,N_23333);
nand U24260 (N_24260,N_23803,N_23139);
nor U24261 (N_24261,N_23748,N_23250);
xor U24262 (N_24262,N_23741,N_23149);
and U24263 (N_24263,N_22803,N_22818);
nor U24264 (N_24264,N_23132,N_23084);
or U24265 (N_24265,N_23492,N_23959);
or U24266 (N_24266,N_22979,N_22962);
nor U24267 (N_24267,N_23119,N_23075);
nand U24268 (N_24268,N_23536,N_22804);
nor U24269 (N_24269,N_23161,N_22913);
and U24270 (N_24270,N_23025,N_23818);
and U24271 (N_24271,N_22969,N_22844);
xnor U24272 (N_24272,N_23237,N_23974);
nor U24273 (N_24273,N_23197,N_23365);
and U24274 (N_24274,N_22860,N_23404);
xnor U24275 (N_24275,N_23473,N_22853);
or U24276 (N_24276,N_23225,N_23676);
nand U24277 (N_24277,N_23402,N_22875);
or U24278 (N_24278,N_23544,N_23019);
or U24279 (N_24279,N_23509,N_23419);
or U24280 (N_24280,N_23474,N_22955);
or U24281 (N_24281,N_23283,N_23456);
xor U24282 (N_24282,N_23899,N_23703);
nor U24283 (N_24283,N_22938,N_23890);
nand U24284 (N_24284,N_23956,N_22891);
and U24285 (N_24285,N_22817,N_23705);
or U24286 (N_24286,N_23802,N_23997);
nor U24287 (N_24287,N_22811,N_23448);
and U24288 (N_24288,N_23450,N_23399);
nand U24289 (N_24289,N_23795,N_23349);
and U24290 (N_24290,N_23363,N_23532);
xor U24291 (N_24291,N_23603,N_23755);
nand U24292 (N_24292,N_23213,N_23328);
and U24293 (N_24293,N_23167,N_23175);
nor U24294 (N_24294,N_23654,N_23593);
xor U24295 (N_24295,N_23353,N_23983);
xor U24296 (N_24296,N_23863,N_23441);
nand U24297 (N_24297,N_23209,N_23269);
nand U24298 (N_24298,N_23050,N_23817);
nor U24299 (N_24299,N_23942,N_23624);
nand U24300 (N_24300,N_23729,N_23648);
nor U24301 (N_24301,N_23221,N_22833);
xor U24302 (N_24302,N_22892,N_23618);
and U24303 (N_24303,N_23655,N_23157);
xor U24304 (N_24304,N_23274,N_23730);
or U24305 (N_24305,N_23427,N_23110);
nand U24306 (N_24306,N_23602,N_23462);
nor U24307 (N_24307,N_23564,N_23163);
nand U24308 (N_24308,N_22956,N_22994);
xnor U24309 (N_24309,N_23409,N_22828);
nor U24310 (N_24310,N_23088,N_23856);
nor U24311 (N_24311,N_23742,N_22810);
nor U24312 (N_24312,N_23380,N_23179);
nor U24313 (N_24313,N_22985,N_23433);
xor U24314 (N_24314,N_23458,N_23103);
xor U24315 (N_24315,N_23198,N_23206);
or U24316 (N_24316,N_22993,N_22825);
and U24317 (N_24317,N_23396,N_23821);
or U24318 (N_24318,N_23255,N_22881);
nand U24319 (N_24319,N_23769,N_23643);
xnor U24320 (N_24320,N_23385,N_23725);
nand U24321 (N_24321,N_23707,N_22865);
nand U24322 (N_24322,N_23556,N_23991);
nor U24323 (N_24323,N_23335,N_22971);
nor U24324 (N_24324,N_22907,N_23418);
nand U24325 (N_24325,N_23391,N_22929);
nand U24326 (N_24326,N_23816,N_23453);
or U24327 (N_24327,N_23226,N_23375);
or U24328 (N_24328,N_23794,N_23081);
or U24329 (N_24329,N_22970,N_23809);
or U24330 (N_24330,N_23557,N_23840);
nand U24331 (N_24331,N_23862,N_23222);
nand U24332 (N_24332,N_23190,N_23289);
or U24333 (N_24333,N_23766,N_22937);
and U24334 (N_24334,N_23931,N_23004);
or U24335 (N_24335,N_23428,N_23204);
nor U24336 (N_24336,N_23650,N_23034);
xnor U24337 (N_24337,N_23285,N_23675);
xor U24338 (N_24338,N_23029,N_23105);
nand U24339 (N_24339,N_23099,N_23526);
xor U24340 (N_24340,N_23280,N_22957);
nand U24341 (N_24341,N_23483,N_23045);
or U24342 (N_24342,N_22905,N_23122);
and U24343 (N_24343,N_23040,N_23235);
or U24344 (N_24344,N_23383,N_23434);
or U24345 (N_24345,N_22986,N_23003);
nand U24346 (N_24346,N_23251,N_23710);
or U24347 (N_24347,N_23253,N_22961);
and U24348 (N_24348,N_23013,N_23950);
nor U24349 (N_24349,N_23887,N_23904);
nor U24350 (N_24350,N_22855,N_23721);
nand U24351 (N_24351,N_23150,N_23342);
nand U24352 (N_24352,N_23500,N_23140);
xnor U24353 (N_24353,N_23351,N_22849);
and U24354 (N_24354,N_23749,N_23696);
or U24355 (N_24355,N_23682,N_23102);
nand U24356 (N_24356,N_22944,N_23248);
nor U24357 (N_24357,N_23220,N_23617);
or U24358 (N_24358,N_23475,N_23032);
nor U24359 (N_24359,N_23978,N_23615);
nor U24360 (N_24360,N_23368,N_23398);
and U24361 (N_24361,N_23293,N_23507);
nand U24362 (N_24362,N_22978,N_22885);
nor U24363 (N_24363,N_23561,N_23726);
and U24364 (N_24364,N_23244,N_23954);
nand U24365 (N_24365,N_23781,N_23499);
and U24366 (N_24366,N_23169,N_23866);
xor U24367 (N_24367,N_23266,N_23195);
and U24368 (N_24368,N_23924,N_23129);
nand U24369 (N_24369,N_23165,N_23772);
xor U24370 (N_24370,N_23423,N_23252);
nor U24371 (N_24371,N_23926,N_23623);
and U24372 (N_24372,N_23819,N_23745);
xor U24373 (N_24373,N_23095,N_23256);
nor U24374 (N_24374,N_23571,N_23563);
and U24375 (N_24375,N_23401,N_23895);
xor U24376 (N_24376,N_23000,N_23440);
or U24377 (N_24377,N_23928,N_23651);
nor U24378 (N_24378,N_23693,N_23096);
xnor U24379 (N_24379,N_23092,N_23331);
xnor U24380 (N_24380,N_23243,N_23713);
or U24381 (N_24381,N_23218,N_23168);
nand U24382 (N_24382,N_23845,N_23068);
nand U24383 (N_24383,N_23591,N_23761);
or U24384 (N_24384,N_23893,N_23558);
nand U24385 (N_24385,N_23486,N_23622);
or U24386 (N_24386,N_22912,N_23914);
or U24387 (N_24387,N_23174,N_23718);
nor U24388 (N_24388,N_22820,N_23952);
nor U24389 (N_24389,N_23471,N_23091);
or U24390 (N_24390,N_23788,N_23697);
nor U24391 (N_24391,N_23960,N_23302);
or U24392 (N_24392,N_22882,N_22987);
xor U24393 (N_24393,N_23875,N_23377);
xnor U24394 (N_24394,N_23927,N_23259);
or U24395 (N_24395,N_23046,N_23016);
nor U24396 (N_24396,N_23849,N_22894);
nor U24397 (N_24397,N_23210,N_23936);
nor U24398 (N_24398,N_23431,N_23724);
xnor U24399 (N_24399,N_23604,N_23281);
and U24400 (N_24400,N_23652,N_23275);
and U24401 (N_24401,N_22859,N_23348);
nand U24402 (N_24402,N_22940,N_23124);
or U24403 (N_24403,N_23988,N_22841);
or U24404 (N_24404,N_23970,N_23701);
and U24405 (N_24405,N_23825,N_23026);
nor U24406 (N_24406,N_22898,N_23627);
nand U24407 (N_24407,N_22914,N_23971);
nand U24408 (N_24408,N_23247,N_23205);
nand U24409 (N_24409,N_23393,N_23432);
xnor U24410 (N_24410,N_23415,N_23646);
nor U24411 (N_24411,N_23079,N_22976);
and U24412 (N_24412,N_23597,N_23452);
nor U24413 (N_24413,N_23868,N_22806);
nand U24414 (N_24414,N_23038,N_23097);
or U24415 (N_24415,N_23184,N_23104);
nand U24416 (N_24416,N_22910,N_23909);
and U24417 (N_24417,N_23551,N_23265);
and U24418 (N_24418,N_23231,N_23477);
or U24419 (N_24419,N_23260,N_23148);
nor U24420 (N_24420,N_23439,N_23940);
nand U24421 (N_24421,N_23808,N_23633);
nor U24422 (N_24422,N_23666,N_23596);
nor U24423 (N_24423,N_22973,N_23058);
nor U24424 (N_24424,N_23229,N_23753);
nor U24425 (N_24425,N_23659,N_22925);
xnor U24426 (N_24426,N_23720,N_23547);
nor U24427 (N_24427,N_23582,N_23495);
xor U24428 (N_24428,N_23632,N_23715);
or U24429 (N_24429,N_22862,N_23086);
nand U24430 (N_24430,N_22846,N_23411);
xor U24431 (N_24431,N_23879,N_23607);
xor U24432 (N_24432,N_22950,N_22984);
or U24433 (N_24433,N_23294,N_23142);
nand U24434 (N_24434,N_23240,N_23496);
or U24435 (N_24435,N_23487,N_23882);
and U24436 (N_24436,N_23517,N_23519);
and U24437 (N_24437,N_23531,N_23538);
xnor U24438 (N_24438,N_22917,N_23989);
xor U24439 (N_24439,N_23698,N_23339);
nand U24440 (N_24440,N_23390,N_23299);
or U24441 (N_24441,N_23867,N_22842);
nand U24442 (N_24442,N_23768,N_22919);
or U24443 (N_24443,N_23437,N_23017);
xor U24444 (N_24444,N_23601,N_23647);
nand U24445 (N_24445,N_23023,N_23965);
nand U24446 (N_24446,N_23336,N_23332);
xnor U24447 (N_24447,N_23629,N_23614);
xor U24448 (N_24448,N_22989,N_23939);
or U24449 (N_24449,N_23762,N_23491);
nand U24450 (N_24450,N_23843,N_23224);
and U24451 (N_24451,N_23138,N_22887);
and U24452 (N_24452,N_23979,N_23637);
xor U24453 (N_24453,N_23941,N_23395);
nand U24454 (N_24454,N_23443,N_23018);
nand U24455 (N_24455,N_23683,N_23660);
and U24456 (N_24456,N_22858,N_23295);
nor U24457 (N_24457,N_23667,N_23792);
nor U24458 (N_24458,N_23578,N_23562);
and U24459 (N_24459,N_23635,N_23694);
xor U24460 (N_24460,N_23630,N_23844);
and U24461 (N_24461,N_23864,N_23925);
and U24462 (N_24462,N_23417,N_22895);
xor U24463 (N_24463,N_23838,N_23461);
xor U24464 (N_24464,N_23746,N_23855);
and U24465 (N_24465,N_23505,N_22948);
nand U24466 (N_24466,N_22992,N_23196);
nor U24467 (N_24467,N_23653,N_23318);
nand U24468 (N_24468,N_23118,N_23670);
nand U24469 (N_24469,N_23922,N_23580);
nand U24470 (N_24470,N_22924,N_23888);
nand U24471 (N_24471,N_23889,N_23714);
nand U24472 (N_24472,N_22879,N_23176);
nand U24473 (N_24473,N_23886,N_23460);
xor U24474 (N_24474,N_23413,N_23063);
nand U24475 (N_24475,N_23442,N_23608);
nand U24476 (N_24476,N_22982,N_23445);
nand U24477 (N_24477,N_22947,N_23747);
nand U24478 (N_24478,N_23429,N_23523);
and U24479 (N_24479,N_23810,N_22877);
or U24480 (N_24480,N_23852,N_23527);
nand U24481 (N_24481,N_22945,N_23054);
and U24482 (N_24482,N_23780,N_23227);
xnor U24483 (N_24483,N_23199,N_23386);
nand U24484 (N_24484,N_23030,N_23783);
nand U24485 (N_24485,N_22801,N_22958);
nand U24486 (N_24486,N_23717,N_23777);
and U24487 (N_24487,N_23546,N_23271);
nand U24488 (N_24488,N_23961,N_22953);
nor U24489 (N_24489,N_23488,N_23201);
and U24490 (N_24490,N_23619,N_23731);
nor U24491 (N_24491,N_22902,N_23223);
nor U24492 (N_24492,N_23055,N_23773);
or U24493 (N_24493,N_23929,N_23716);
or U24494 (N_24494,N_23542,N_23153);
xnor U24495 (N_24495,N_22851,N_23569);
nor U24496 (N_24496,N_23876,N_23543);
or U24497 (N_24497,N_23217,N_23270);
xnor U24498 (N_24498,N_22930,N_23776);
and U24499 (N_24499,N_23346,N_23207);
or U24500 (N_24500,N_23027,N_23007);
and U24501 (N_24501,N_23494,N_23425);
and U24502 (N_24502,N_23530,N_22972);
nand U24503 (N_24503,N_23644,N_23782);
xnor U24504 (N_24504,N_23309,N_23963);
nand U24505 (N_24505,N_23089,N_22847);
xor U24506 (N_24506,N_22805,N_23966);
nor U24507 (N_24507,N_23277,N_23001);
nor U24508 (N_24508,N_23506,N_23669);
nand U24509 (N_24509,N_23976,N_23330);
xor U24510 (N_24510,N_23115,N_23382);
xnor U24511 (N_24511,N_23784,N_23189);
xor U24512 (N_24512,N_23359,N_22834);
nor U24513 (N_24513,N_23313,N_23290);
or U24514 (N_24514,N_23403,N_23739);
xnor U24515 (N_24515,N_22802,N_22830);
nor U24516 (N_24516,N_23216,N_23662);
nand U24517 (N_24517,N_23534,N_23191);
xor U24518 (N_24518,N_23869,N_23896);
nor U24519 (N_24519,N_23469,N_23797);
nand U24520 (N_24520,N_22922,N_23605);
and U24521 (N_24521,N_23518,N_23476);
nand U24522 (N_24522,N_22927,N_23514);
xnor U24523 (N_24523,N_23897,N_23388);
nand U24524 (N_24524,N_23537,N_23957);
or U24525 (N_24525,N_22869,N_23917);
and U24526 (N_24526,N_23857,N_23587);
xor U24527 (N_24527,N_23136,N_23993);
nor U24528 (N_24528,N_23664,N_23512);
nand U24529 (N_24529,N_23472,N_23438);
xnor U24530 (N_24530,N_23945,N_22906);
nand U24531 (N_24531,N_23200,N_23625);
and U24532 (N_24532,N_23861,N_23829);
or U24533 (N_24533,N_23436,N_23069);
and U24534 (N_24534,N_23261,N_23858);
nor U24535 (N_24535,N_23078,N_23567);
xnor U24536 (N_24536,N_23341,N_23986);
nand U24537 (N_24537,N_23422,N_23590);
xnor U24538 (N_24538,N_23376,N_23117);
xor U24539 (N_24539,N_23668,N_23839);
and U24540 (N_24540,N_23234,N_23836);
nand U24541 (N_24541,N_23985,N_22900);
xnor U24542 (N_24542,N_23430,N_23884);
nor U24543 (N_24543,N_23356,N_22915);
nor U24544 (N_24544,N_23246,N_23230);
xnor U24545 (N_24545,N_23090,N_22823);
xnor U24546 (N_24546,N_23405,N_23020);
nand U24547 (N_24547,N_23338,N_23815);
nand U24548 (N_24548,N_23870,N_23750);
or U24549 (N_24549,N_23631,N_23765);
and U24550 (N_24550,N_23022,N_22923);
nor U24551 (N_24551,N_23898,N_23347);
xor U24552 (N_24552,N_22909,N_23282);
nor U24553 (N_24553,N_23951,N_23120);
nor U24554 (N_24554,N_23325,N_23589);
and U24555 (N_24555,N_23737,N_23577);
and U24556 (N_24556,N_23592,N_23126);
nand U24557 (N_24557,N_23953,N_23288);
nand U24558 (N_24558,N_23481,N_23877);
and U24559 (N_24559,N_23493,N_23125);
xor U24560 (N_24560,N_23764,N_23374);
and U24561 (N_24561,N_22832,N_23113);
nor U24562 (N_24562,N_23489,N_23327);
nand U24563 (N_24563,N_23695,N_23574);
nor U24564 (N_24564,N_23921,N_23389);
nor U24565 (N_24565,N_23098,N_22807);
nand U24566 (N_24566,N_23361,N_23326);
nand U24567 (N_24567,N_22965,N_23464);
or U24568 (N_24568,N_23560,N_23919);
nor U24569 (N_24569,N_23649,N_23482);
nor U24570 (N_24570,N_23751,N_23972);
and U24571 (N_24571,N_23535,N_23872);
nand U24572 (N_24572,N_23006,N_22835);
and U24573 (N_24573,N_23314,N_23012);
xnor U24574 (N_24574,N_23770,N_23609);
nor U24575 (N_24575,N_23123,N_22843);
nand U24576 (N_24576,N_23340,N_22822);
or U24577 (N_24577,N_23576,N_23923);
nand U24578 (N_24578,N_23791,N_23214);
xor U24579 (N_24579,N_23407,N_23947);
or U24580 (N_24580,N_23891,N_23702);
nor U24581 (N_24581,N_23323,N_23352);
nand U24582 (N_24582,N_23699,N_22857);
nor U24583 (N_24583,N_23860,N_23579);
xnor U24584 (N_24584,N_23053,N_23379);
or U24585 (N_24585,N_22870,N_23062);
nand U24586 (N_24586,N_23446,N_23594);
or U24587 (N_24587,N_23661,N_23043);
or U24588 (N_24588,N_23370,N_23540);
nand U24589 (N_24589,N_23192,N_23145);
nor U24590 (N_24590,N_23892,N_23740);
nand U24591 (N_24591,N_23178,N_23767);
and U24592 (N_24592,N_23734,N_23665);
nand U24593 (N_24593,N_22899,N_23943);
nand U24594 (N_24594,N_23121,N_23219);
nor U24595 (N_24595,N_23905,N_23254);
xor U24596 (N_24596,N_23822,N_23128);
nand U24597 (N_24597,N_23141,N_22996);
nand U24598 (N_24598,N_23706,N_23938);
nand U24599 (N_24599,N_23982,N_23820);
nand U24600 (N_24600,N_23670,N_23133);
nor U24601 (N_24601,N_23404,N_23602);
and U24602 (N_24602,N_23034,N_23802);
xnor U24603 (N_24603,N_22978,N_23514);
and U24604 (N_24604,N_23079,N_23353);
nor U24605 (N_24605,N_22953,N_23997);
xor U24606 (N_24606,N_23509,N_23225);
and U24607 (N_24607,N_23681,N_23431);
or U24608 (N_24608,N_23686,N_23806);
nor U24609 (N_24609,N_23323,N_22896);
or U24610 (N_24610,N_23741,N_22808);
xor U24611 (N_24611,N_23806,N_23032);
and U24612 (N_24612,N_23751,N_23403);
and U24613 (N_24613,N_23476,N_23384);
nand U24614 (N_24614,N_23008,N_23127);
nand U24615 (N_24615,N_23287,N_22811);
nand U24616 (N_24616,N_23957,N_23413);
xnor U24617 (N_24617,N_23335,N_23781);
or U24618 (N_24618,N_23704,N_23024);
or U24619 (N_24619,N_23351,N_23253);
xor U24620 (N_24620,N_23996,N_23257);
nor U24621 (N_24621,N_23177,N_23108);
xnor U24622 (N_24622,N_22885,N_23721);
nand U24623 (N_24623,N_22816,N_22937);
or U24624 (N_24624,N_23480,N_23163);
xnor U24625 (N_24625,N_22868,N_23613);
and U24626 (N_24626,N_23677,N_23565);
nor U24627 (N_24627,N_22963,N_23918);
xnor U24628 (N_24628,N_23085,N_23209);
nor U24629 (N_24629,N_23045,N_23233);
nor U24630 (N_24630,N_23300,N_23042);
and U24631 (N_24631,N_23866,N_23053);
and U24632 (N_24632,N_23529,N_23586);
nor U24633 (N_24633,N_23701,N_23698);
or U24634 (N_24634,N_23144,N_23413);
nor U24635 (N_24635,N_23632,N_23678);
or U24636 (N_24636,N_23387,N_23567);
nand U24637 (N_24637,N_23771,N_22856);
nand U24638 (N_24638,N_23656,N_23630);
and U24639 (N_24639,N_23613,N_23118);
nor U24640 (N_24640,N_23506,N_23366);
or U24641 (N_24641,N_22967,N_23571);
nor U24642 (N_24642,N_22859,N_23307);
or U24643 (N_24643,N_23231,N_23311);
nor U24644 (N_24644,N_23462,N_23912);
nand U24645 (N_24645,N_23470,N_23721);
nor U24646 (N_24646,N_22885,N_23298);
nand U24647 (N_24647,N_23228,N_23893);
or U24648 (N_24648,N_23684,N_23205);
xnor U24649 (N_24649,N_23678,N_22846);
xor U24650 (N_24650,N_23839,N_23048);
or U24651 (N_24651,N_23002,N_23970);
and U24652 (N_24652,N_23484,N_23697);
nand U24653 (N_24653,N_23680,N_23125);
or U24654 (N_24654,N_23477,N_23481);
nor U24655 (N_24655,N_23466,N_23485);
or U24656 (N_24656,N_23686,N_23058);
nand U24657 (N_24657,N_23700,N_23997);
or U24658 (N_24658,N_22958,N_23045);
nor U24659 (N_24659,N_23985,N_23315);
nor U24660 (N_24660,N_23424,N_23253);
and U24661 (N_24661,N_23420,N_23241);
or U24662 (N_24662,N_23003,N_23251);
or U24663 (N_24663,N_23927,N_23043);
and U24664 (N_24664,N_23293,N_23157);
nand U24665 (N_24665,N_23683,N_23030);
nand U24666 (N_24666,N_23617,N_22959);
nor U24667 (N_24667,N_23260,N_23789);
nand U24668 (N_24668,N_23898,N_23836);
nand U24669 (N_24669,N_23846,N_23676);
and U24670 (N_24670,N_23316,N_23415);
xnor U24671 (N_24671,N_23938,N_23068);
or U24672 (N_24672,N_23761,N_23954);
xnor U24673 (N_24673,N_23483,N_23900);
or U24674 (N_24674,N_23933,N_23781);
xor U24675 (N_24675,N_23294,N_22928);
or U24676 (N_24676,N_23337,N_23943);
and U24677 (N_24677,N_23962,N_23236);
nand U24678 (N_24678,N_22886,N_23935);
or U24679 (N_24679,N_22817,N_23301);
and U24680 (N_24680,N_23608,N_23309);
and U24681 (N_24681,N_23174,N_23319);
and U24682 (N_24682,N_23504,N_23807);
xnor U24683 (N_24683,N_23748,N_22846);
xor U24684 (N_24684,N_23889,N_23111);
xnor U24685 (N_24685,N_22935,N_23122);
nor U24686 (N_24686,N_23546,N_23811);
nor U24687 (N_24687,N_23600,N_23471);
nand U24688 (N_24688,N_23704,N_23769);
nor U24689 (N_24689,N_23443,N_23377);
xor U24690 (N_24690,N_23824,N_22919);
nand U24691 (N_24691,N_23663,N_23532);
nor U24692 (N_24692,N_23182,N_23610);
or U24693 (N_24693,N_23910,N_23181);
nand U24694 (N_24694,N_23368,N_23685);
or U24695 (N_24695,N_23173,N_23174);
and U24696 (N_24696,N_23991,N_23982);
and U24697 (N_24697,N_23678,N_23197);
xnor U24698 (N_24698,N_22970,N_23408);
nand U24699 (N_24699,N_22930,N_23631);
or U24700 (N_24700,N_23390,N_23050);
nand U24701 (N_24701,N_23386,N_23857);
and U24702 (N_24702,N_23080,N_23386);
and U24703 (N_24703,N_23432,N_23264);
or U24704 (N_24704,N_23313,N_23126);
nor U24705 (N_24705,N_23207,N_23712);
or U24706 (N_24706,N_23462,N_23683);
or U24707 (N_24707,N_23415,N_23495);
or U24708 (N_24708,N_23556,N_23314);
nor U24709 (N_24709,N_23842,N_22958);
nand U24710 (N_24710,N_22882,N_23902);
and U24711 (N_24711,N_22830,N_23618);
xor U24712 (N_24712,N_23693,N_23422);
and U24713 (N_24713,N_22815,N_23854);
nor U24714 (N_24714,N_23421,N_22998);
and U24715 (N_24715,N_23551,N_23668);
xnor U24716 (N_24716,N_23430,N_23510);
nor U24717 (N_24717,N_22964,N_23037);
nand U24718 (N_24718,N_23537,N_23946);
and U24719 (N_24719,N_23497,N_23279);
nor U24720 (N_24720,N_23547,N_23133);
or U24721 (N_24721,N_23476,N_23870);
nor U24722 (N_24722,N_23870,N_22894);
nand U24723 (N_24723,N_22807,N_23623);
xor U24724 (N_24724,N_22932,N_23641);
or U24725 (N_24725,N_23189,N_23353);
nor U24726 (N_24726,N_23121,N_23169);
and U24727 (N_24727,N_22919,N_22889);
nor U24728 (N_24728,N_23084,N_23975);
xor U24729 (N_24729,N_23105,N_23096);
nand U24730 (N_24730,N_23807,N_23551);
nand U24731 (N_24731,N_23966,N_23103);
xor U24732 (N_24732,N_23015,N_23521);
nand U24733 (N_24733,N_23468,N_23808);
and U24734 (N_24734,N_22909,N_23602);
nor U24735 (N_24735,N_23196,N_23047);
nand U24736 (N_24736,N_23728,N_23138);
nand U24737 (N_24737,N_23884,N_23997);
xnor U24738 (N_24738,N_22924,N_23954);
nand U24739 (N_24739,N_23726,N_23633);
or U24740 (N_24740,N_23345,N_23493);
nor U24741 (N_24741,N_23156,N_23341);
xnor U24742 (N_24742,N_23681,N_23295);
xnor U24743 (N_24743,N_23432,N_22890);
and U24744 (N_24744,N_23566,N_23856);
nor U24745 (N_24745,N_22823,N_23022);
nand U24746 (N_24746,N_23506,N_23039);
xor U24747 (N_24747,N_23204,N_23601);
and U24748 (N_24748,N_23847,N_23730);
nor U24749 (N_24749,N_22989,N_23390);
or U24750 (N_24750,N_23812,N_23985);
nand U24751 (N_24751,N_23150,N_23327);
nor U24752 (N_24752,N_23098,N_23505);
xnor U24753 (N_24753,N_23680,N_22932);
and U24754 (N_24754,N_22864,N_23882);
nor U24755 (N_24755,N_23667,N_23354);
xor U24756 (N_24756,N_23964,N_23083);
and U24757 (N_24757,N_23111,N_23897);
and U24758 (N_24758,N_23138,N_23788);
xor U24759 (N_24759,N_23317,N_23042);
nand U24760 (N_24760,N_23957,N_23324);
nand U24761 (N_24761,N_23112,N_22854);
xnor U24762 (N_24762,N_23894,N_23987);
or U24763 (N_24763,N_23424,N_23613);
and U24764 (N_24764,N_23696,N_23052);
xor U24765 (N_24765,N_23356,N_23092);
and U24766 (N_24766,N_23423,N_23067);
xnor U24767 (N_24767,N_23108,N_23842);
and U24768 (N_24768,N_23535,N_23596);
and U24769 (N_24769,N_23134,N_23766);
or U24770 (N_24770,N_23793,N_23317);
nor U24771 (N_24771,N_23219,N_23020);
and U24772 (N_24772,N_23660,N_23400);
nand U24773 (N_24773,N_23509,N_23948);
xnor U24774 (N_24774,N_23539,N_23339);
nand U24775 (N_24775,N_23505,N_23936);
xor U24776 (N_24776,N_23853,N_22948);
xnor U24777 (N_24777,N_23471,N_23571);
or U24778 (N_24778,N_23055,N_23012);
nor U24779 (N_24779,N_23031,N_23516);
and U24780 (N_24780,N_23442,N_23489);
xnor U24781 (N_24781,N_23041,N_23248);
xnor U24782 (N_24782,N_23788,N_22889);
nor U24783 (N_24783,N_23442,N_23454);
xnor U24784 (N_24784,N_23001,N_22881);
xnor U24785 (N_24785,N_22962,N_23678);
nand U24786 (N_24786,N_23545,N_23983);
xnor U24787 (N_24787,N_23070,N_23169);
nor U24788 (N_24788,N_23459,N_23903);
xnor U24789 (N_24789,N_23838,N_23155);
xnor U24790 (N_24790,N_23297,N_22945);
xor U24791 (N_24791,N_23387,N_23176);
xor U24792 (N_24792,N_23322,N_23501);
nand U24793 (N_24793,N_23023,N_23117);
xnor U24794 (N_24794,N_23148,N_23704);
xnor U24795 (N_24795,N_23146,N_23441);
nand U24796 (N_24796,N_23938,N_23698);
xor U24797 (N_24797,N_23469,N_23197);
nand U24798 (N_24798,N_23815,N_23097);
and U24799 (N_24799,N_23341,N_23756);
nand U24800 (N_24800,N_23329,N_23475);
and U24801 (N_24801,N_23194,N_23619);
nand U24802 (N_24802,N_23430,N_23879);
or U24803 (N_24803,N_23781,N_22947);
and U24804 (N_24804,N_22841,N_22949);
and U24805 (N_24805,N_23187,N_22966);
nand U24806 (N_24806,N_23647,N_22864);
xnor U24807 (N_24807,N_23512,N_23830);
xor U24808 (N_24808,N_23326,N_23126);
nor U24809 (N_24809,N_23512,N_23807);
xor U24810 (N_24810,N_23400,N_23063);
xor U24811 (N_24811,N_23492,N_22800);
or U24812 (N_24812,N_23282,N_23110);
nor U24813 (N_24813,N_22876,N_23330);
or U24814 (N_24814,N_23428,N_23962);
and U24815 (N_24815,N_22864,N_23030);
nand U24816 (N_24816,N_23619,N_22839);
nand U24817 (N_24817,N_23872,N_23209);
nand U24818 (N_24818,N_23207,N_23539);
xnor U24819 (N_24819,N_23731,N_23533);
xnor U24820 (N_24820,N_23935,N_23852);
nand U24821 (N_24821,N_23823,N_23226);
or U24822 (N_24822,N_23784,N_22852);
nor U24823 (N_24823,N_23948,N_23745);
xnor U24824 (N_24824,N_23076,N_22817);
xor U24825 (N_24825,N_23303,N_23769);
or U24826 (N_24826,N_23053,N_23455);
nor U24827 (N_24827,N_23818,N_23213);
nor U24828 (N_24828,N_23188,N_23250);
xnor U24829 (N_24829,N_23793,N_23529);
xnor U24830 (N_24830,N_23483,N_23204);
and U24831 (N_24831,N_23103,N_23631);
nor U24832 (N_24832,N_23791,N_22803);
and U24833 (N_24833,N_23470,N_23962);
or U24834 (N_24834,N_23092,N_23195);
nand U24835 (N_24835,N_23485,N_23513);
xor U24836 (N_24836,N_22900,N_23283);
nand U24837 (N_24837,N_23222,N_23560);
and U24838 (N_24838,N_23195,N_23827);
xor U24839 (N_24839,N_23166,N_22955);
xnor U24840 (N_24840,N_23562,N_23418);
or U24841 (N_24841,N_23968,N_23470);
nor U24842 (N_24842,N_23993,N_23513);
nand U24843 (N_24843,N_22912,N_23654);
or U24844 (N_24844,N_23803,N_23383);
or U24845 (N_24845,N_22904,N_23308);
nand U24846 (N_24846,N_23250,N_23382);
xnor U24847 (N_24847,N_23822,N_22957);
or U24848 (N_24848,N_23288,N_23646);
nor U24849 (N_24849,N_23858,N_23568);
nand U24850 (N_24850,N_23289,N_23612);
and U24851 (N_24851,N_22893,N_22921);
nand U24852 (N_24852,N_23652,N_23612);
nand U24853 (N_24853,N_23797,N_23026);
nand U24854 (N_24854,N_23589,N_23709);
or U24855 (N_24855,N_23440,N_23294);
nor U24856 (N_24856,N_23612,N_23635);
or U24857 (N_24857,N_23905,N_23633);
nor U24858 (N_24858,N_22915,N_23390);
or U24859 (N_24859,N_23736,N_23289);
or U24860 (N_24860,N_23026,N_23986);
nor U24861 (N_24861,N_23074,N_22890);
nand U24862 (N_24862,N_22839,N_23754);
nand U24863 (N_24863,N_23114,N_23261);
or U24864 (N_24864,N_23357,N_23317);
and U24865 (N_24865,N_23137,N_23774);
nor U24866 (N_24866,N_22994,N_23936);
and U24867 (N_24867,N_23522,N_22955);
xor U24868 (N_24868,N_23230,N_23420);
and U24869 (N_24869,N_23433,N_23681);
nand U24870 (N_24870,N_23393,N_23216);
xnor U24871 (N_24871,N_23045,N_23923);
nand U24872 (N_24872,N_23395,N_23273);
nor U24873 (N_24873,N_23315,N_23156);
nand U24874 (N_24874,N_23340,N_23365);
and U24875 (N_24875,N_23481,N_23168);
or U24876 (N_24876,N_23698,N_23088);
nand U24877 (N_24877,N_23277,N_23475);
nor U24878 (N_24878,N_23276,N_22919);
and U24879 (N_24879,N_23571,N_23110);
xnor U24880 (N_24880,N_23801,N_23886);
and U24881 (N_24881,N_23196,N_23739);
nor U24882 (N_24882,N_23336,N_23441);
nand U24883 (N_24883,N_23292,N_23694);
or U24884 (N_24884,N_23854,N_23205);
and U24885 (N_24885,N_23741,N_23126);
or U24886 (N_24886,N_23120,N_23577);
nand U24887 (N_24887,N_23906,N_23850);
nand U24888 (N_24888,N_23733,N_22859);
and U24889 (N_24889,N_23575,N_23347);
or U24890 (N_24890,N_23157,N_23985);
xnor U24891 (N_24891,N_23918,N_23411);
or U24892 (N_24892,N_23265,N_23550);
nor U24893 (N_24893,N_23445,N_23539);
and U24894 (N_24894,N_23106,N_23825);
and U24895 (N_24895,N_23561,N_23730);
or U24896 (N_24896,N_23629,N_23130);
or U24897 (N_24897,N_23031,N_22980);
xor U24898 (N_24898,N_23864,N_23875);
nand U24899 (N_24899,N_23371,N_23640);
nand U24900 (N_24900,N_23103,N_23514);
nor U24901 (N_24901,N_23030,N_22989);
nor U24902 (N_24902,N_23041,N_23191);
and U24903 (N_24903,N_23726,N_23052);
xor U24904 (N_24904,N_22956,N_23069);
and U24905 (N_24905,N_23297,N_22929);
and U24906 (N_24906,N_23281,N_23778);
and U24907 (N_24907,N_23361,N_23403);
or U24908 (N_24908,N_23534,N_23572);
nor U24909 (N_24909,N_23818,N_22959);
xor U24910 (N_24910,N_23986,N_22952);
xnor U24911 (N_24911,N_23687,N_22868);
nand U24912 (N_24912,N_23052,N_23837);
or U24913 (N_24913,N_23045,N_23453);
or U24914 (N_24914,N_23726,N_23094);
and U24915 (N_24915,N_23311,N_23509);
and U24916 (N_24916,N_22945,N_23755);
nand U24917 (N_24917,N_23103,N_23406);
xor U24918 (N_24918,N_22882,N_23559);
nor U24919 (N_24919,N_23424,N_23024);
and U24920 (N_24920,N_22847,N_23661);
xor U24921 (N_24921,N_23504,N_23649);
xor U24922 (N_24922,N_23736,N_23151);
nand U24923 (N_24923,N_23619,N_23516);
and U24924 (N_24924,N_23742,N_23972);
and U24925 (N_24925,N_23625,N_23125);
xnor U24926 (N_24926,N_23036,N_23890);
nand U24927 (N_24927,N_23192,N_23305);
or U24928 (N_24928,N_23483,N_22990);
xnor U24929 (N_24929,N_22915,N_22824);
or U24930 (N_24930,N_23138,N_23962);
or U24931 (N_24931,N_23018,N_22851);
xor U24932 (N_24932,N_23164,N_23329);
nor U24933 (N_24933,N_23669,N_23941);
nand U24934 (N_24934,N_23769,N_23931);
or U24935 (N_24935,N_23588,N_23500);
nand U24936 (N_24936,N_23095,N_23223);
nand U24937 (N_24937,N_22982,N_23123);
xor U24938 (N_24938,N_23766,N_23333);
or U24939 (N_24939,N_23661,N_23013);
xor U24940 (N_24940,N_22974,N_23190);
xor U24941 (N_24941,N_23521,N_23666);
nand U24942 (N_24942,N_23533,N_23879);
nand U24943 (N_24943,N_23158,N_23929);
nor U24944 (N_24944,N_23583,N_23843);
nand U24945 (N_24945,N_23795,N_23696);
and U24946 (N_24946,N_23788,N_23242);
nand U24947 (N_24947,N_23143,N_23781);
nor U24948 (N_24948,N_23393,N_23210);
nor U24949 (N_24949,N_22948,N_23334);
or U24950 (N_24950,N_23479,N_23914);
or U24951 (N_24951,N_23707,N_22812);
nor U24952 (N_24952,N_23151,N_22964);
xor U24953 (N_24953,N_23119,N_23508);
nor U24954 (N_24954,N_23308,N_23655);
nor U24955 (N_24955,N_23537,N_23183);
and U24956 (N_24956,N_23175,N_22841);
or U24957 (N_24957,N_23674,N_22898);
xnor U24958 (N_24958,N_23913,N_23888);
nor U24959 (N_24959,N_23775,N_23362);
or U24960 (N_24960,N_23597,N_23951);
and U24961 (N_24961,N_23326,N_23810);
and U24962 (N_24962,N_23801,N_23262);
nand U24963 (N_24963,N_22988,N_23255);
or U24964 (N_24964,N_23328,N_23293);
and U24965 (N_24965,N_23479,N_22976);
and U24966 (N_24966,N_22851,N_23586);
or U24967 (N_24967,N_23617,N_22953);
nor U24968 (N_24968,N_23204,N_23077);
xnor U24969 (N_24969,N_23216,N_23643);
or U24970 (N_24970,N_23642,N_23439);
xor U24971 (N_24971,N_23023,N_22939);
xor U24972 (N_24972,N_23242,N_23305);
and U24973 (N_24973,N_23487,N_23165);
and U24974 (N_24974,N_22818,N_22957);
xnor U24975 (N_24975,N_23288,N_22899);
nor U24976 (N_24976,N_23818,N_23468);
nand U24977 (N_24977,N_23304,N_23001);
nand U24978 (N_24978,N_23692,N_22869);
or U24979 (N_24979,N_23439,N_23712);
nand U24980 (N_24980,N_23474,N_23904);
nand U24981 (N_24981,N_23186,N_23927);
xnor U24982 (N_24982,N_23744,N_23495);
and U24983 (N_24983,N_23117,N_23242);
and U24984 (N_24984,N_23294,N_23826);
or U24985 (N_24985,N_23026,N_23547);
nor U24986 (N_24986,N_23106,N_23590);
nand U24987 (N_24987,N_23370,N_22818);
nor U24988 (N_24988,N_23031,N_23289);
nor U24989 (N_24989,N_23201,N_23097);
xnor U24990 (N_24990,N_23491,N_23940);
or U24991 (N_24991,N_22818,N_23257);
nand U24992 (N_24992,N_23199,N_23986);
xor U24993 (N_24993,N_23437,N_23645);
xor U24994 (N_24994,N_23920,N_23251);
nand U24995 (N_24995,N_23457,N_23778);
xnor U24996 (N_24996,N_23047,N_22972);
xnor U24997 (N_24997,N_23261,N_23619);
nor U24998 (N_24998,N_23859,N_23953);
xor U24999 (N_24999,N_23699,N_23718);
xnor U25000 (N_25000,N_23524,N_23444);
nor U25001 (N_25001,N_23136,N_23963);
or U25002 (N_25002,N_23781,N_23749);
and U25003 (N_25003,N_23307,N_23578);
and U25004 (N_25004,N_23207,N_22819);
xor U25005 (N_25005,N_23713,N_23429);
or U25006 (N_25006,N_23536,N_23157);
or U25007 (N_25007,N_23052,N_23566);
nor U25008 (N_25008,N_23228,N_23974);
and U25009 (N_25009,N_23025,N_23310);
or U25010 (N_25010,N_23961,N_23212);
and U25011 (N_25011,N_23964,N_23158);
nand U25012 (N_25012,N_22930,N_23023);
nor U25013 (N_25013,N_23373,N_23687);
xnor U25014 (N_25014,N_23234,N_23448);
or U25015 (N_25015,N_23468,N_22846);
or U25016 (N_25016,N_23037,N_23700);
xor U25017 (N_25017,N_23747,N_23136);
and U25018 (N_25018,N_23671,N_22974);
nand U25019 (N_25019,N_23485,N_22949);
nand U25020 (N_25020,N_23912,N_23600);
xor U25021 (N_25021,N_23743,N_22878);
and U25022 (N_25022,N_23874,N_22869);
xnor U25023 (N_25023,N_23340,N_23772);
and U25024 (N_25024,N_23848,N_23513);
nor U25025 (N_25025,N_23703,N_23778);
xnor U25026 (N_25026,N_23481,N_23358);
nor U25027 (N_25027,N_23466,N_23247);
nand U25028 (N_25028,N_23454,N_22842);
or U25029 (N_25029,N_22811,N_22954);
xor U25030 (N_25030,N_23984,N_23053);
or U25031 (N_25031,N_23613,N_23926);
nor U25032 (N_25032,N_23693,N_23592);
xor U25033 (N_25033,N_23428,N_23063);
xor U25034 (N_25034,N_23486,N_23168);
and U25035 (N_25035,N_22890,N_22837);
or U25036 (N_25036,N_23351,N_23119);
nor U25037 (N_25037,N_23208,N_23716);
and U25038 (N_25038,N_23754,N_23716);
nand U25039 (N_25039,N_23781,N_23543);
xor U25040 (N_25040,N_23374,N_22816);
or U25041 (N_25041,N_23590,N_22834);
nor U25042 (N_25042,N_23357,N_23803);
xnor U25043 (N_25043,N_23925,N_22981);
nor U25044 (N_25044,N_23167,N_23285);
or U25045 (N_25045,N_23039,N_23553);
xnor U25046 (N_25046,N_22980,N_23006);
and U25047 (N_25047,N_23365,N_23462);
xnor U25048 (N_25048,N_23609,N_23815);
nand U25049 (N_25049,N_23860,N_22816);
nand U25050 (N_25050,N_23790,N_23245);
and U25051 (N_25051,N_23531,N_23163);
nand U25052 (N_25052,N_22969,N_23421);
or U25053 (N_25053,N_22856,N_23246);
and U25054 (N_25054,N_23716,N_23939);
nor U25055 (N_25055,N_23438,N_23744);
and U25056 (N_25056,N_23948,N_23468);
nor U25057 (N_25057,N_23925,N_23717);
nand U25058 (N_25058,N_23155,N_23970);
nand U25059 (N_25059,N_22816,N_23367);
nor U25060 (N_25060,N_22883,N_23270);
and U25061 (N_25061,N_23284,N_23557);
nand U25062 (N_25062,N_23613,N_23793);
or U25063 (N_25063,N_23821,N_23569);
or U25064 (N_25064,N_23625,N_23832);
nor U25065 (N_25065,N_23586,N_23808);
and U25066 (N_25066,N_23468,N_22907);
and U25067 (N_25067,N_23241,N_23955);
xor U25068 (N_25068,N_23025,N_23647);
or U25069 (N_25069,N_22857,N_23700);
or U25070 (N_25070,N_23728,N_23855);
nor U25071 (N_25071,N_23443,N_22999);
nand U25072 (N_25072,N_22925,N_23972);
xor U25073 (N_25073,N_23232,N_23178);
nor U25074 (N_25074,N_23735,N_22897);
or U25075 (N_25075,N_23445,N_23439);
and U25076 (N_25076,N_23467,N_23248);
and U25077 (N_25077,N_23592,N_23563);
xnor U25078 (N_25078,N_23848,N_23308);
or U25079 (N_25079,N_23530,N_23406);
nor U25080 (N_25080,N_22842,N_23653);
and U25081 (N_25081,N_23899,N_22847);
nor U25082 (N_25082,N_23246,N_23280);
and U25083 (N_25083,N_23151,N_23640);
or U25084 (N_25084,N_23359,N_23744);
and U25085 (N_25085,N_23445,N_23462);
nor U25086 (N_25086,N_23599,N_22953);
nor U25087 (N_25087,N_23850,N_22980);
and U25088 (N_25088,N_22900,N_23022);
xnor U25089 (N_25089,N_23964,N_23286);
and U25090 (N_25090,N_23022,N_23273);
nand U25091 (N_25091,N_23336,N_23518);
and U25092 (N_25092,N_23163,N_22834);
xnor U25093 (N_25093,N_22884,N_22930);
and U25094 (N_25094,N_23165,N_23619);
or U25095 (N_25095,N_23386,N_23631);
nor U25096 (N_25096,N_23968,N_23750);
xor U25097 (N_25097,N_23094,N_22939);
nand U25098 (N_25098,N_22837,N_23519);
nor U25099 (N_25099,N_22864,N_22946);
xnor U25100 (N_25100,N_22918,N_23236);
nor U25101 (N_25101,N_23743,N_23024);
nor U25102 (N_25102,N_23530,N_23527);
or U25103 (N_25103,N_23458,N_23109);
and U25104 (N_25104,N_22838,N_23319);
and U25105 (N_25105,N_22842,N_23830);
and U25106 (N_25106,N_23562,N_22927);
or U25107 (N_25107,N_23173,N_23171);
nor U25108 (N_25108,N_23323,N_23496);
xor U25109 (N_25109,N_23797,N_23030);
and U25110 (N_25110,N_23843,N_22952);
or U25111 (N_25111,N_23563,N_23407);
nor U25112 (N_25112,N_22984,N_23142);
xnor U25113 (N_25113,N_23789,N_23108);
nand U25114 (N_25114,N_22944,N_23482);
or U25115 (N_25115,N_23961,N_23259);
and U25116 (N_25116,N_23701,N_23204);
xor U25117 (N_25117,N_23155,N_23239);
and U25118 (N_25118,N_23585,N_23458);
xnor U25119 (N_25119,N_23092,N_23330);
and U25120 (N_25120,N_23967,N_23867);
and U25121 (N_25121,N_22947,N_23568);
nand U25122 (N_25122,N_22828,N_23207);
and U25123 (N_25123,N_22863,N_22982);
nand U25124 (N_25124,N_23182,N_23308);
and U25125 (N_25125,N_23584,N_23371);
nor U25126 (N_25126,N_23226,N_23570);
xnor U25127 (N_25127,N_23477,N_23431);
xor U25128 (N_25128,N_23296,N_23574);
nor U25129 (N_25129,N_23732,N_23482);
and U25130 (N_25130,N_23401,N_22806);
or U25131 (N_25131,N_23803,N_23872);
nand U25132 (N_25132,N_23991,N_23876);
xor U25133 (N_25133,N_23371,N_23888);
and U25134 (N_25134,N_22871,N_22807);
xnor U25135 (N_25135,N_23570,N_23816);
nor U25136 (N_25136,N_23011,N_22983);
xnor U25137 (N_25137,N_22962,N_23763);
nor U25138 (N_25138,N_23103,N_23827);
xnor U25139 (N_25139,N_23862,N_23124);
and U25140 (N_25140,N_23480,N_23926);
xor U25141 (N_25141,N_23301,N_23049);
xor U25142 (N_25142,N_23715,N_23457);
xnor U25143 (N_25143,N_23462,N_23082);
nor U25144 (N_25144,N_23154,N_23421);
xnor U25145 (N_25145,N_23933,N_23054);
xor U25146 (N_25146,N_23277,N_23754);
nor U25147 (N_25147,N_23525,N_23928);
nand U25148 (N_25148,N_23688,N_23505);
nor U25149 (N_25149,N_23256,N_22874);
nand U25150 (N_25150,N_23720,N_23965);
xnor U25151 (N_25151,N_22969,N_23757);
nor U25152 (N_25152,N_22964,N_22808);
or U25153 (N_25153,N_23711,N_23623);
or U25154 (N_25154,N_23209,N_23952);
xor U25155 (N_25155,N_23573,N_23841);
nor U25156 (N_25156,N_23377,N_23376);
nor U25157 (N_25157,N_23506,N_23621);
or U25158 (N_25158,N_23932,N_23323);
nand U25159 (N_25159,N_23464,N_22941);
nand U25160 (N_25160,N_23620,N_23098);
nand U25161 (N_25161,N_23470,N_22908);
and U25162 (N_25162,N_23101,N_23313);
or U25163 (N_25163,N_22829,N_23301);
xnor U25164 (N_25164,N_22991,N_23397);
nand U25165 (N_25165,N_23860,N_23081);
and U25166 (N_25166,N_23938,N_23161);
xnor U25167 (N_25167,N_23098,N_23550);
nor U25168 (N_25168,N_23928,N_23438);
xnor U25169 (N_25169,N_23686,N_23413);
or U25170 (N_25170,N_23520,N_23308);
xor U25171 (N_25171,N_23184,N_23140);
or U25172 (N_25172,N_23021,N_23681);
and U25173 (N_25173,N_23670,N_23578);
or U25174 (N_25174,N_23568,N_23637);
and U25175 (N_25175,N_23125,N_23148);
nor U25176 (N_25176,N_22947,N_23437);
and U25177 (N_25177,N_23331,N_23591);
or U25178 (N_25178,N_23703,N_23307);
nor U25179 (N_25179,N_23820,N_23881);
xnor U25180 (N_25180,N_23152,N_23539);
and U25181 (N_25181,N_23200,N_23604);
nand U25182 (N_25182,N_23447,N_23310);
and U25183 (N_25183,N_23494,N_23455);
nand U25184 (N_25184,N_23861,N_23898);
and U25185 (N_25185,N_23540,N_23240);
nand U25186 (N_25186,N_23289,N_22993);
nand U25187 (N_25187,N_23565,N_23668);
xor U25188 (N_25188,N_23868,N_23069);
and U25189 (N_25189,N_23468,N_23472);
nand U25190 (N_25190,N_23329,N_23059);
nand U25191 (N_25191,N_23669,N_23500);
nand U25192 (N_25192,N_23180,N_23888);
nand U25193 (N_25193,N_22881,N_23479);
nand U25194 (N_25194,N_22912,N_23628);
and U25195 (N_25195,N_23487,N_23479);
nand U25196 (N_25196,N_23883,N_23885);
nand U25197 (N_25197,N_22922,N_23385);
or U25198 (N_25198,N_22886,N_23239);
and U25199 (N_25199,N_23858,N_23284);
nand U25200 (N_25200,N_25197,N_24877);
or U25201 (N_25201,N_24575,N_24313);
and U25202 (N_25202,N_24826,N_24646);
nor U25203 (N_25203,N_24344,N_25100);
nor U25204 (N_25204,N_24043,N_24704);
xor U25205 (N_25205,N_24483,N_24198);
xor U25206 (N_25206,N_24723,N_24712);
or U25207 (N_25207,N_24276,N_24657);
xor U25208 (N_25208,N_24599,N_24267);
nand U25209 (N_25209,N_24223,N_24967);
and U25210 (N_25210,N_24938,N_24536);
nand U25211 (N_25211,N_24190,N_24025);
xor U25212 (N_25212,N_25175,N_24399);
nor U25213 (N_25213,N_24560,N_24376);
and U25214 (N_25214,N_24838,N_24858);
xor U25215 (N_25215,N_25014,N_24435);
and U25216 (N_25216,N_24624,N_24266);
nor U25217 (N_25217,N_24887,N_24587);
nor U25218 (N_25218,N_24749,N_24264);
and U25219 (N_25219,N_24208,N_24500);
nand U25220 (N_25220,N_24908,N_24841);
nor U25221 (N_25221,N_25180,N_24679);
nand U25222 (N_25222,N_24300,N_24662);
and U25223 (N_25223,N_24386,N_24547);
nand U25224 (N_25224,N_24345,N_24821);
or U25225 (N_25225,N_24041,N_24305);
xor U25226 (N_25226,N_24647,N_24224);
nand U25227 (N_25227,N_24971,N_24144);
or U25228 (N_25228,N_24335,N_25138);
nor U25229 (N_25229,N_24894,N_24576);
nor U25230 (N_25230,N_25061,N_24367);
nand U25231 (N_25231,N_24660,N_25086);
nor U25232 (N_25232,N_24930,N_24308);
and U25233 (N_25233,N_24180,N_24436);
or U25234 (N_25234,N_24869,N_25163);
nor U25235 (N_25235,N_25105,N_24847);
nand U25236 (N_25236,N_24853,N_24814);
and U25237 (N_25237,N_25004,N_24382);
nor U25238 (N_25238,N_24282,N_24607);
or U25239 (N_25239,N_24685,N_24842);
or U25240 (N_25240,N_24066,N_24178);
or U25241 (N_25241,N_25150,N_24013);
nand U25242 (N_25242,N_24102,N_24966);
or U25243 (N_25243,N_25085,N_24922);
nor U25244 (N_25244,N_24824,N_24788);
nand U25245 (N_25245,N_24298,N_24811);
nor U25246 (N_25246,N_24242,N_24863);
xnor U25247 (N_25247,N_24935,N_25081);
or U25248 (N_25248,N_25152,N_24537);
and U25249 (N_25249,N_24825,N_24548);
or U25250 (N_25250,N_24727,N_24565);
or U25251 (N_25251,N_25063,N_25065);
nand U25252 (N_25252,N_24453,N_24911);
nand U25253 (N_25253,N_25096,N_24076);
nor U25254 (N_25254,N_25189,N_25076);
xnor U25255 (N_25255,N_24918,N_24172);
nand U25256 (N_25256,N_24176,N_24441);
and U25257 (N_25257,N_24095,N_24862);
and U25258 (N_25258,N_24580,N_24529);
nor U25259 (N_25259,N_25083,N_24110);
or U25260 (N_25260,N_24125,N_25160);
or U25261 (N_25261,N_24014,N_24752);
nand U25262 (N_25262,N_24538,N_24249);
xor U25263 (N_25263,N_24810,N_24087);
or U25264 (N_25264,N_24527,N_25003);
nor U25265 (N_25265,N_24852,N_24868);
and U25266 (N_25266,N_24322,N_24316);
nand U25267 (N_25267,N_24762,N_24092);
nor U25268 (N_25268,N_24986,N_24212);
nor U25269 (N_25269,N_24141,N_24118);
and U25270 (N_25270,N_25088,N_24388);
and U25271 (N_25271,N_24238,N_24107);
nand U25272 (N_25272,N_24042,N_25069);
and U25273 (N_25273,N_24237,N_24126);
nand U25274 (N_25274,N_24627,N_24928);
nor U25275 (N_25275,N_24256,N_25046);
nand U25276 (N_25276,N_24876,N_24979);
and U25277 (N_25277,N_24162,N_24086);
and U25278 (N_25278,N_24691,N_24395);
or U25279 (N_25279,N_24579,N_24705);
nor U25280 (N_25280,N_24796,N_24807);
or U25281 (N_25281,N_24173,N_24800);
and U25282 (N_25282,N_24121,N_24596);
xor U25283 (N_25283,N_25055,N_24904);
and U25284 (N_25284,N_24301,N_24027);
nand U25285 (N_25285,N_25198,N_24571);
xor U25286 (N_25286,N_24912,N_24044);
xnor U25287 (N_25287,N_24955,N_24650);
xnor U25288 (N_25288,N_24372,N_24953);
nand U25289 (N_25289,N_24433,N_24974);
nand U25290 (N_25290,N_24693,N_25114);
xnor U25291 (N_25291,N_24247,N_24845);
and U25292 (N_25292,N_24377,N_24613);
xor U25293 (N_25293,N_24706,N_24248);
nor U25294 (N_25294,N_24612,N_24989);
nor U25295 (N_25295,N_25178,N_24010);
and U25296 (N_25296,N_25157,N_24584);
and U25297 (N_25297,N_24421,N_25002);
or U25298 (N_25298,N_24499,N_24332);
or U25299 (N_25299,N_24915,N_25130);
nand U25300 (N_25300,N_24420,N_24883);
or U25301 (N_25301,N_24397,N_24898);
xor U25302 (N_25302,N_24558,N_25171);
or U25303 (N_25303,N_24431,N_25037);
xor U25304 (N_25304,N_24713,N_24336);
or U25305 (N_25305,N_24188,N_24664);
or U25306 (N_25306,N_24504,N_24848);
xor U25307 (N_25307,N_25191,N_24396);
nand U25308 (N_25308,N_25054,N_24556);
nand U25309 (N_25309,N_25186,N_25190);
nand U25310 (N_25310,N_24018,N_24775);
nand U25311 (N_25311,N_24849,N_24972);
nor U25312 (N_25312,N_25077,N_24632);
xor U25313 (N_25313,N_25050,N_24150);
or U25314 (N_25314,N_24402,N_24220);
nor U25315 (N_25315,N_25124,N_24780);
or U25316 (N_25316,N_24988,N_25030);
or U25317 (N_25317,N_24302,N_24473);
nand U25318 (N_25318,N_24668,N_24231);
xor U25319 (N_25319,N_24429,N_24774);
and U25320 (N_25320,N_24658,N_24490);
xnor U25321 (N_25321,N_24460,N_24213);
nor U25322 (N_25322,N_24506,N_24736);
nand U25323 (N_25323,N_24003,N_24861);
nand U25324 (N_25324,N_24748,N_24046);
xor U25325 (N_25325,N_24724,N_24589);
xnor U25326 (N_25326,N_24535,N_24641);
and U25327 (N_25327,N_24370,N_24128);
or U25328 (N_25328,N_25068,N_24326);
or U25329 (N_25329,N_24378,N_24284);
or U25330 (N_25330,N_25079,N_24899);
or U25331 (N_25331,N_24151,N_24757);
nand U25332 (N_25332,N_24562,N_24457);
or U25333 (N_25333,N_24754,N_24735);
xnor U25334 (N_25334,N_24552,N_24358);
xor U25335 (N_25335,N_24525,N_24005);
or U25336 (N_25336,N_24709,N_24717);
and U25337 (N_25337,N_24227,N_25128);
xnor U25338 (N_25338,N_24278,N_24608);
nand U25339 (N_25339,N_24982,N_24343);
xor U25340 (N_25340,N_25052,N_24152);
xnor U25341 (N_25341,N_24689,N_24291);
nand U25342 (N_25342,N_24487,N_24446);
nand U25343 (N_25343,N_24255,N_24037);
nand U25344 (N_25344,N_24885,N_24716);
or U25345 (N_25345,N_24634,N_24744);
nor U25346 (N_25346,N_24207,N_24884);
nor U25347 (N_25347,N_25182,N_24969);
nand U25348 (N_25348,N_24452,N_25194);
xor U25349 (N_25349,N_24232,N_24732);
and U25350 (N_25350,N_25013,N_24430);
nor U25351 (N_25351,N_24671,N_24163);
nor U25352 (N_25352,N_24828,N_24745);
and U25353 (N_25353,N_24482,N_24342);
nand U25354 (N_25354,N_24447,N_25159);
xnor U25355 (N_25355,N_24577,N_25170);
xor U25356 (N_25356,N_24352,N_24476);
xor U25357 (N_25357,N_24604,N_24054);
xor U25358 (N_25358,N_25093,N_25035);
nor U25359 (N_25359,N_24687,N_24669);
or U25360 (N_25360,N_25108,N_24792);
and U25361 (N_25361,N_24077,N_24550);
nor U25362 (N_25362,N_24813,N_24035);
nand U25363 (N_25363,N_24667,N_24827);
xnor U25364 (N_25364,N_24361,N_24914);
or U25365 (N_25365,N_24139,N_24878);
or U25366 (N_25366,N_25045,N_25110);
or U25367 (N_25367,N_24517,N_25167);
or U25368 (N_25368,N_24177,N_24722);
nor U25369 (N_25369,N_24374,N_24357);
nand U25370 (N_25370,N_24015,N_25078);
nor U25371 (N_25371,N_25067,N_24844);
xor U25372 (N_25372,N_25192,N_24130);
nand U25373 (N_25373,N_24870,N_24082);
and U25374 (N_25374,N_24038,N_24566);
and U25375 (N_25375,N_24590,N_24407);
xnor U25376 (N_25376,N_25010,N_24683);
or U25377 (N_25377,N_24965,N_25195);
or U25378 (N_25378,N_24049,N_24696);
nor U25379 (N_25379,N_24002,N_24170);
nor U25380 (N_25380,N_24616,N_24184);
nor U25381 (N_25381,N_24896,N_24715);
or U25382 (N_25382,N_24823,N_24970);
nand U25383 (N_25383,N_24602,N_24321);
xor U25384 (N_25384,N_25144,N_24202);
nand U25385 (N_25385,N_24663,N_24428);
nor U25386 (N_25386,N_24611,N_24893);
nor U25387 (N_25387,N_25120,N_24498);
xor U25388 (N_25388,N_24697,N_24366);
or U25389 (N_25389,N_24155,N_24065);
or U25390 (N_25390,N_24931,N_24491);
and U25391 (N_25391,N_24103,N_24078);
nor U25392 (N_25392,N_24281,N_24992);
xnor U25393 (N_25393,N_24161,N_24618);
nand U25394 (N_25394,N_24750,N_24761);
nor U25395 (N_25395,N_24069,N_24888);
and U25396 (N_25396,N_24629,N_24983);
nor U25397 (N_25397,N_24633,N_25087);
xnor U25398 (N_25398,N_24711,N_24261);
nor U25399 (N_25399,N_24021,N_24872);
and U25400 (N_25400,N_24245,N_24528);
nand U25401 (N_25401,N_24623,N_24976);
or U25402 (N_25402,N_24354,N_24648);
xor U25403 (N_25403,N_25156,N_25143);
or U25404 (N_25404,N_24785,N_24910);
or U25405 (N_25405,N_24568,N_24234);
xor U25406 (N_25406,N_24230,N_25173);
and U25407 (N_25407,N_24606,N_24288);
nand U25408 (N_25408,N_24140,N_24977);
xor U25409 (N_25409,N_24494,N_25089);
xor U25410 (N_25410,N_25099,N_24119);
and U25411 (N_25411,N_24383,N_24007);
nand U25412 (N_25412,N_25176,N_24698);
xnor U25413 (N_25413,N_24085,N_24625);
and U25414 (N_25414,N_25084,N_24600);
nand U25415 (N_25415,N_24142,N_24747);
and U25416 (N_25416,N_24100,N_24090);
xor U25417 (N_25417,N_25172,N_25074);
nand U25418 (N_25418,N_24790,N_24450);
nand U25419 (N_25419,N_24751,N_24993);
nor U25420 (N_25420,N_24240,N_25095);
nand U25421 (N_25421,N_24419,N_24991);
and U25422 (N_25422,N_25132,N_24763);
or U25423 (N_25423,N_24053,N_24501);
and U25424 (N_25424,N_24665,N_24465);
nor U25425 (N_25425,N_24192,N_24471);
and U25426 (N_25426,N_24124,N_24760);
or U25427 (N_25427,N_24205,N_24975);
or U25428 (N_25428,N_25059,N_24941);
nor U25429 (N_25429,N_25036,N_24505);
nor U25430 (N_25430,N_24225,N_24017);
and U25431 (N_25431,N_24182,N_24478);
nand U25432 (N_25432,N_24289,N_24403);
xnor U25433 (N_25433,N_24112,N_24617);
or U25434 (N_25434,N_25162,N_24574);
nand U25435 (N_25435,N_24416,N_24166);
nand U25436 (N_25436,N_25001,N_24864);
and U25437 (N_25437,N_25134,N_24635);
or U25438 (N_25438,N_24319,N_24593);
or U25439 (N_25439,N_24806,N_24831);
or U25440 (N_25440,N_24001,N_24269);
xnor U25441 (N_25441,N_24742,N_24059);
and U25442 (N_25442,N_24531,N_24680);
or U25443 (N_25443,N_24939,N_24226);
and U25444 (N_25444,N_24060,N_24275);
xor U25445 (N_25445,N_24642,N_24116);
or U25446 (N_25446,N_24443,N_24432);
or U25447 (N_25447,N_24294,N_24157);
xor U25448 (N_25448,N_24486,N_24214);
nand U25449 (N_25449,N_24138,N_24109);
xor U25450 (N_25450,N_24349,N_24555);
nand U25451 (N_25451,N_25053,N_24659);
nor U25452 (N_25452,N_24767,N_25022);
and U25453 (N_25453,N_24945,N_24250);
nor U25454 (N_25454,N_24561,N_24995);
and U25455 (N_25455,N_24011,N_24306);
nor U25456 (N_25456,N_24328,N_25181);
or U25457 (N_25457,N_24253,N_24964);
and U25458 (N_25458,N_25148,N_24519);
nor U25459 (N_25459,N_24064,N_25111);
nand U25460 (N_25460,N_24364,N_24263);
and U25461 (N_25461,N_24228,N_24047);
and U25462 (N_25462,N_24962,N_24181);
xnor U25463 (N_25463,N_25109,N_24191);
nor U25464 (N_25464,N_24619,N_24802);
or U25465 (N_25465,N_24426,N_24200);
nand U25466 (N_25466,N_24739,N_25155);
nand U25467 (N_25467,N_24470,N_25048);
or U25468 (N_25468,N_24148,N_24083);
nand U25469 (N_25469,N_24690,N_24406);
nor U25470 (N_25470,N_24394,N_24472);
or U25471 (N_25471,N_24120,N_24892);
nand U25472 (N_25472,N_24401,N_25141);
nand U25473 (N_25473,N_25188,N_24028);
nor U25474 (N_25474,N_24008,N_24147);
or U25475 (N_25475,N_24673,N_24438);
or U25476 (N_25476,N_24503,N_24681);
and U25477 (N_25477,N_24515,N_24895);
nor U25478 (N_25478,N_24956,N_24424);
nand U25479 (N_25479,N_25016,N_24265);
nand U25480 (N_25480,N_24016,N_24084);
nor U25481 (N_25481,N_24886,N_25137);
xor U25482 (N_25482,N_24303,N_24521);
xor U25483 (N_25483,N_24423,N_24277);
xnor U25484 (N_25484,N_24973,N_25165);
and U25485 (N_25485,N_24094,N_25106);
and U25486 (N_25486,N_24943,N_24039);
nand U25487 (N_25487,N_24067,N_24652);
nor U25488 (N_25488,N_24929,N_24413);
and U25489 (N_25489,N_25071,N_24645);
xnor U25490 (N_25490,N_24738,N_24818);
nor U25491 (N_25491,N_24009,N_24540);
or U25492 (N_25492,N_24179,N_24360);
xnor U25493 (N_25493,N_24781,N_24135);
nand U25494 (N_25494,N_24753,N_25112);
nand U25495 (N_25495,N_24809,N_25153);
nor U25496 (N_25496,N_24497,N_24081);
and U25497 (N_25497,N_24553,N_24570);
xnor U25498 (N_25498,N_24317,N_24398);
or U25499 (N_25499,N_24740,N_24820);
nor U25500 (N_25500,N_24508,N_25184);
nor U25501 (N_25501,N_24907,N_25140);
and U25502 (N_25502,N_25019,N_24541);
nand U25503 (N_25503,N_24734,N_24857);
and U25504 (N_25504,N_24835,N_25070);
or U25505 (N_25505,N_24113,N_24631);
and U25506 (N_25506,N_24355,N_24985);
nor U25507 (N_25507,N_25161,N_24375);
nor U25508 (N_25508,N_24614,N_24451);
xor U25509 (N_25509,N_24477,N_24871);
nor U25510 (N_25510,N_25121,N_24479);
xnor U25511 (N_25511,N_24408,N_24856);
nor U25512 (N_25512,N_25135,N_24115);
and U25513 (N_25513,N_24867,N_24987);
or U25514 (N_25514,N_24731,N_24649);
xnor U25515 (N_25515,N_24379,N_24549);
xnor U25516 (N_25516,N_24158,N_24514);
nor U25517 (N_25517,N_24105,N_24485);
nor U25518 (N_25518,N_24484,N_24789);
nand U25519 (N_25519,N_24311,N_25018);
xor U25520 (N_25520,N_25107,N_25015);
or U25521 (N_25521,N_24033,N_24511);
and U25522 (N_25522,N_24159,N_25094);
nor U25523 (N_25523,N_24071,N_24244);
xor U25524 (N_25524,N_24628,N_25064);
xor U25525 (N_25525,N_24595,N_24341);
xnor U25526 (N_25526,N_24427,N_25028);
and U25527 (N_25527,N_24675,N_24239);
and U25528 (N_25528,N_24193,N_25080);
and U25529 (N_25529,N_24339,N_24546);
xnor U25530 (N_25530,N_24651,N_24850);
or U25531 (N_25531,N_25139,N_24522);
or U25532 (N_25532,N_24353,N_24145);
nor U25533 (N_25533,N_24798,N_24733);
and U25534 (N_25534,N_24165,N_24620);
nand U25535 (N_25535,N_24097,N_24846);
and U25536 (N_25536,N_24605,N_24925);
nor U25537 (N_25537,N_24154,N_24463);
or U25538 (N_25538,N_24695,N_24369);
nand U25539 (N_25539,N_25166,N_24672);
or U25540 (N_25540,N_24666,N_24307);
or U25541 (N_25541,N_25193,N_24480);
xnor U25542 (N_25542,N_24510,N_24567);
nor U25543 (N_25543,N_24146,N_24949);
nor U25544 (N_25544,N_24944,N_25098);
nor U25545 (N_25545,N_24834,N_24304);
or U25546 (N_25546,N_24725,N_24801);
nor U25547 (N_25547,N_24822,N_24578);
nand U25548 (N_25548,N_24688,N_24072);
xnor U25549 (N_25549,N_25122,N_24475);
nor U25550 (N_25550,N_24338,N_24458);
xor U25551 (N_25551,N_24833,N_24678);
or U25552 (N_25552,N_24891,N_24805);
xnor U25553 (N_25553,N_24917,N_24773);
nor U25554 (N_25554,N_25020,N_24293);
xnor U25555 (N_25555,N_25091,N_24051);
and U25556 (N_25556,N_24919,N_24902);
or U25557 (N_25557,N_24554,N_24609);
and U25558 (N_25558,N_24246,N_24900);
nand U25559 (N_25559,N_24699,N_24252);
and U25560 (N_25560,N_24088,N_24829);
nand U25561 (N_25561,N_24999,N_24004);
nand U25562 (N_25562,N_25117,N_25103);
and U25563 (N_25563,N_24099,N_24653);
or U25564 (N_25564,N_25072,N_24559);
nand U25565 (N_25565,N_24012,N_24786);
and U25566 (N_25566,N_24516,N_25168);
and U25567 (N_25567,N_24312,N_24371);
and U25568 (N_25568,N_24320,N_25012);
or U25569 (N_25569,N_24075,N_24462);
nor U25570 (N_25570,N_24981,N_24889);
xnor U25571 (N_25571,N_24409,N_24405);
nand U25572 (N_25572,N_24348,N_24643);
nor U25573 (N_25573,N_24836,N_24933);
nand U25574 (N_25574,N_24639,N_24461);
nor U25575 (N_25575,N_25123,N_24700);
and U25576 (N_25576,N_24728,N_24502);
and U25577 (N_25577,N_24185,N_24074);
and U25578 (N_25578,N_24350,N_24737);
or U25579 (N_25579,N_24318,N_24656);
or U25580 (N_25580,N_24947,N_24765);
nor U25581 (N_25581,N_24950,N_24417);
nor U25582 (N_25582,N_24030,N_24840);
nand U25583 (N_25583,N_24913,N_25142);
xnor U25584 (N_25584,N_24260,N_24539);
and U25585 (N_25585,N_25126,N_24542);
nand U25586 (N_25586,N_24272,N_24636);
xor U25587 (N_25587,N_24286,N_24123);
nor U25588 (N_25588,N_24839,N_24381);
nor U25589 (N_25589,N_24544,N_24410);
xnor U25590 (N_25590,N_24023,N_25174);
or U25591 (N_25591,N_24601,N_24880);
nand U25592 (N_25592,N_24936,N_24832);
xnor U25593 (N_25593,N_24351,N_24456);
nand U25594 (N_25594,N_24903,N_24127);
nand U25595 (N_25595,N_24564,N_24873);
and U25596 (N_25596,N_24916,N_24056);
or U25597 (N_25597,N_25177,N_25187);
and U25598 (N_25598,N_24229,N_25090);
nand U25599 (N_25599,N_24026,N_24812);
xnor U25600 (N_25600,N_24766,N_25154);
nor U25601 (N_25601,N_24325,N_24143);
nand U25602 (N_25602,N_24957,N_24093);
xor U25603 (N_25603,N_24927,N_24776);
xnor U25604 (N_25604,N_24759,N_24134);
nor U25605 (N_25605,N_24389,N_24106);
and U25606 (N_25606,N_24924,N_25102);
and U25607 (N_25607,N_24048,N_24032);
xnor U25608 (N_25608,N_25127,N_24132);
nand U25609 (N_25609,N_25136,N_24440);
nand U25610 (N_25610,N_24670,N_24183);
nand U25611 (N_25611,N_24187,N_24117);
or U25612 (N_25612,N_24445,N_24206);
xnor U25613 (N_25613,N_24512,N_24236);
nor U25614 (N_25614,N_24865,N_24794);
xnor U25615 (N_25615,N_25023,N_24783);
xnor U25616 (N_25616,N_24797,N_24464);
nand U25617 (N_25617,N_24960,N_24569);
nor U25618 (N_25618,N_24948,N_24830);
xnor U25619 (N_25619,N_24040,N_24215);
xor U25620 (N_25620,N_25196,N_24387);
xnor U25621 (N_25621,N_25158,N_24283);
xnor U25622 (N_25622,N_25104,N_24203);
nor U25623 (N_25623,N_24996,N_24233);
xnor U25624 (N_25624,N_24347,N_24391);
and U25625 (N_25625,N_25075,N_25043);
xor U25626 (N_25626,N_25118,N_25031);
and U25627 (N_25627,N_25033,N_25062);
nor U25628 (N_25628,N_24029,N_24923);
xnor U25629 (N_25629,N_24337,N_24677);
or U25630 (N_25630,N_25021,N_24474);
or U25631 (N_25631,N_24518,N_24764);
nand U25632 (N_25632,N_24052,N_24721);
xor U25633 (N_25633,N_24031,N_25006);
nor U25634 (N_25634,N_24241,N_24926);
nor U25635 (N_25635,N_24720,N_24467);
nand U25636 (N_25636,N_24909,N_24079);
nor U25637 (N_25637,N_25044,N_24285);
xnor U25638 (N_25638,N_24591,N_24920);
and U25639 (N_25639,N_24454,N_24194);
nor U25640 (N_25640,N_24210,N_24598);
nand U25641 (N_25641,N_24603,N_24661);
and U25642 (N_25642,N_24171,N_24492);
and U25643 (N_25643,N_24310,N_25058);
and U25644 (N_25644,N_25034,N_24644);
xor U25645 (N_25645,N_24582,N_24630);
xor U25646 (N_25646,N_24058,N_24133);
nand U25647 (N_25647,N_24777,N_24034);
or U25648 (N_25648,N_25060,N_24175);
xor U25649 (N_25649,N_24297,N_24509);
xnor U25650 (N_25650,N_24978,N_24637);
xor U25651 (N_25651,N_25024,N_24994);
nor U25652 (N_25652,N_24062,N_24686);
xnor U25653 (N_25653,N_24874,N_24984);
nor U25654 (N_25654,N_24533,N_24217);
or U25655 (N_25655,N_24875,N_24692);
nand U25656 (N_25656,N_24622,N_24674);
nor U25657 (N_25657,N_24280,N_24437);
or U25658 (N_25658,N_24346,N_24149);
or U25659 (N_25659,N_24329,N_24418);
nor U25660 (N_25660,N_24890,N_24520);
or U25661 (N_25661,N_24136,N_24543);
nor U25662 (N_25662,N_25026,N_24299);
xor U25663 (N_25663,N_24070,N_24530);
nor U25664 (N_25664,N_24201,N_24489);
nand U25665 (N_25665,N_24131,N_24755);
and U25666 (N_25666,N_24524,N_24455);
xnor U25667 (N_25667,N_25097,N_24586);
and U25668 (N_25668,N_24096,N_24222);
or U25669 (N_25669,N_24694,N_25009);
nand U25670 (N_25670,N_25101,N_24684);
nand U25671 (N_25671,N_24768,N_24816);
xnor U25672 (N_25672,N_24854,N_24111);
nor U25673 (N_25673,N_24024,N_24218);
or U25674 (N_25674,N_24340,N_24710);
nor U25675 (N_25675,N_24434,N_24771);
nor U25676 (N_25676,N_24583,N_24330);
xnor U25677 (N_25677,N_25131,N_24160);
nand U25678 (N_25678,N_25082,N_24209);
nand U25679 (N_25679,N_24174,N_24439);
nor U25680 (N_25680,N_24468,N_24036);
or U25681 (N_25681,N_24385,N_24414);
nor U25682 (N_25682,N_24726,N_24638);
and U25683 (N_25683,N_24496,N_24592);
xor U25684 (N_25684,N_25042,N_24980);
nand U25685 (N_25685,N_24251,N_24729);
xor U25686 (N_25686,N_24268,N_24513);
xnor U25687 (N_25687,N_24309,N_24196);
or U25688 (N_25688,N_24020,N_24881);
and U25689 (N_25689,N_24940,N_25183);
nand U25690 (N_25690,N_24958,N_24101);
and U25691 (N_25691,N_24257,N_25113);
and U25692 (N_25692,N_24221,N_24073);
nand U25693 (N_25693,N_24164,N_25185);
or U25694 (N_25694,N_24156,N_24216);
and U25695 (N_25695,N_25133,N_24815);
nand U25696 (N_25696,N_25116,N_25049);
or U25697 (N_25697,N_24235,N_24314);
or U25698 (N_25698,N_24855,N_24585);
xor U25699 (N_25699,N_24270,N_24756);
and U25700 (N_25700,N_24167,N_24315);
nand U25701 (N_25701,N_25017,N_24019);
and U25702 (N_25702,N_24779,N_25129);
xnor U25703 (N_25703,N_24334,N_24104);
nor U25704 (N_25704,N_24271,N_24851);
nand U25705 (N_25705,N_24168,N_24803);
or U25706 (N_25706,N_25149,N_25151);
or U25707 (N_25707,N_24262,N_24581);
and U25708 (N_25708,N_24997,N_24404);
and U25709 (N_25709,N_24860,N_24295);
xnor U25710 (N_25710,N_24392,N_24859);
xor U25711 (N_25711,N_24843,N_24934);
and U25712 (N_25712,N_24718,N_24791);
or U25713 (N_25713,N_24534,N_24481);
xor U25714 (N_25714,N_25092,N_24195);
and U25715 (N_25715,N_24243,N_24122);
xor U25716 (N_25716,N_24782,N_24610);
nor U25717 (N_25717,N_24746,N_24708);
xnor U25718 (N_25718,N_24954,N_24459);
nor U25719 (N_25719,N_25169,N_24719);
nor U25720 (N_25720,N_24837,N_25057);
xor U25721 (N_25721,N_24682,N_24055);
nor U25722 (N_25722,N_24959,N_24006);
or U25723 (N_25723,N_24921,N_25199);
nand U25724 (N_25724,N_24057,N_24365);
nor U25725 (N_25725,N_24563,N_24507);
xor U25726 (N_25726,N_24654,N_24784);
xnor U25727 (N_25727,N_24951,N_24961);
or U25728 (N_25728,N_24000,N_24089);
xnor U25729 (N_25729,N_24324,N_24626);
nor U25730 (N_25730,N_24068,N_24597);
or U25731 (N_25731,N_24292,N_24572);
nand U25732 (N_25732,N_24061,N_24091);
xnor U25733 (N_25733,N_24819,N_24879);
xor U25734 (N_25734,N_24703,N_24290);
or U25735 (N_25735,N_24523,N_24532);
xnor U25736 (N_25736,N_24990,N_24808);
xor U25737 (N_25737,N_25038,N_24199);
and U25738 (N_25738,N_25066,N_24741);
xnor U25739 (N_25739,N_24274,N_24045);
xnor U25740 (N_25740,N_24362,N_24787);
xnor U25741 (N_25741,N_24770,N_24137);
or U25742 (N_25742,N_24129,N_24080);
xnor U25743 (N_25743,N_24793,N_24799);
xor U25744 (N_25744,N_25040,N_24866);
and U25745 (N_25745,N_24588,N_25027);
xnor U25746 (N_25746,N_24169,N_24551);
nor U25747 (N_25747,N_24259,N_25007);
xnor U25748 (N_25748,N_24714,N_24442);
nor U25749 (N_25749,N_25025,N_24197);
nand U25750 (N_25750,N_24906,N_24393);
nor U25751 (N_25751,N_24368,N_24153);
or U25752 (N_25752,N_25041,N_25005);
or U25753 (N_25753,N_24098,N_25147);
or U25754 (N_25754,N_24937,N_24817);
nor U25755 (N_25755,N_24730,N_24707);
and U25756 (N_25756,N_25119,N_24287);
nand U25757 (N_25757,N_24411,N_24495);
or U25758 (N_25758,N_24380,N_24108);
and U25759 (N_25759,N_24331,N_24573);
nand U25760 (N_25760,N_24743,N_25047);
nor U25761 (N_25761,N_25008,N_25179);
nand U25762 (N_25762,N_25164,N_24621);
nand U25763 (N_25763,N_24882,N_24758);
and U25764 (N_25764,N_24327,N_24279);
and U25765 (N_25765,N_25145,N_24114);
and U25766 (N_25766,N_24412,N_24998);
nor U25767 (N_25767,N_25011,N_24356);
or U25768 (N_25768,N_24373,N_24219);
and U25769 (N_25769,N_24422,N_24701);
nand U25770 (N_25770,N_24384,N_24390);
xnor U25771 (N_25771,N_24425,N_24469);
and U25772 (N_25772,N_24211,N_24296);
or U25773 (N_25773,N_25146,N_24258);
nand U25774 (N_25774,N_24615,N_24905);
xor U25775 (N_25775,N_24968,N_25000);
and U25776 (N_25776,N_24640,N_25032);
and U25777 (N_25777,N_24063,N_24557);
and U25778 (N_25778,N_24778,N_24448);
or U25779 (N_25779,N_24189,N_25051);
xnor U25780 (N_25780,N_24942,N_24359);
and U25781 (N_25781,N_24526,N_24323);
nor U25782 (N_25782,N_24022,N_24676);
nand U25783 (N_25783,N_24254,N_24769);
nand U25784 (N_25784,N_24946,N_24594);
or U25785 (N_25785,N_24655,N_25115);
or U25786 (N_25786,N_24897,N_24204);
nand U25787 (N_25787,N_24952,N_24772);
nand U25788 (N_25788,N_24901,N_24932);
xor U25789 (N_25789,N_25073,N_24804);
xor U25790 (N_25790,N_24333,N_24963);
nand U25791 (N_25791,N_24415,N_24400);
and U25792 (N_25792,N_24795,N_25029);
or U25793 (N_25793,N_24449,N_25056);
and U25794 (N_25794,N_24444,N_24493);
nor U25795 (N_25795,N_25039,N_24488);
and U25796 (N_25796,N_25125,N_24273);
nand U25797 (N_25797,N_24363,N_24545);
nor U25798 (N_25798,N_24702,N_24050);
or U25799 (N_25799,N_24186,N_24466);
nand U25800 (N_25800,N_24921,N_24304);
nor U25801 (N_25801,N_24620,N_24140);
or U25802 (N_25802,N_24901,N_24004);
xor U25803 (N_25803,N_24724,N_25148);
xor U25804 (N_25804,N_25055,N_25182);
xor U25805 (N_25805,N_24718,N_24562);
xnor U25806 (N_25806,N_24897,N_24532);
xor U25807 (N_25807,N_24794,N_24042);
and U25808 (N_25808,N_24015,N_24287);
nand U25809 (N_25809,N_24830,N_24708);
and U25810 (N_25810,N_24224,N_24746);
nand U25811 (N_25811,N_24043,N_24834);
and U25812 (N_25812,N_24062,N_24375);
xor U25813 (N_25813,N_25152,N_24145);
or U25814 (N_25814,N_24249,N_24098);
or U25815 (N_25815,N_24783,N_24817);
nor U25816 (N_25816,N_24709,N_24050);
nor U25817 (N_25817,N_24695,N_24164);
nand U25818 (N_25818,N_25033,N_24406);
or U25819 (N_25819,N_24667,N_24294);
xnor U25820 (N_25820,N_24402,N_24383);
or U25821 (N_25821,N_24377,N_24035);
xor U25822 (N_25822,N_24053,N_24370);
or U25823 (N_25823,N_24911,N_24881);
nand U25824 (N_25824,N_24911,N_24826);
nor U25825 (N_25825,N_25036,N_24456);
nand U25826 (N_25826,N_24229,N_24796);
nor U25827 (N_25827,N_24704,N_24024);
xnor U25828 (N_25828,N_24079,N_24205);
nand U25829 (N_25829,N_24749,N_25138);
nand U25830 (N_25830,N_24083,N_24363);
xnor U25831 (N_25831,N_24382,N_25166);
nand U25832 (N_25832,N_24770,N_24545);
or U25833 (N_25833,N_24558,N_24472);
xnor U25834 (N_25834,N_24844,N_25063);
and U25835 (N_25835,N_25012,N_25108);
nor U25836 (N_25836,N_24217,N_24807);
and U25837 (N_25837,N_24188,N_24875);
nand U25838 (N_25838,N_24081,N_24863);
and U25839 (N_25839,N_24031,N_24585);
nand U25840 (N_25840,N_24340,N_24053);
and U25841 (N_25841,N_24533,N_24152);
and U25842 (N_25842,N_24704,N_24052);
nand U25843 (N_25843,N_25145,N_24300);
or U25844 (N_25844,N_25028,N_24768);
and U25845 (N_25845,N_25188,N_25171);
and U25846 (N_25846,N_24123,N_25195);
xnor U25847 (N_25847,N_24453,N_24234);
nand U25848 (N_25848,N_25111,N_24129);
and U25849 (N_25849,N_24014,N_24210);
xnor U25850 (N_25850,N_24728,N_24921);
nor U25851 (N_25851,N_24650,N_25149);
nor U25852 (N_25852,N_24109,N_24949);
nor U25853 (N_25853,N_25049,N_24282);
xor U25854 (N_25854,N_24718,N_24280);
nand U25855 (N_25855,N_25056,N_24868);
nor U25856 (N_25856,N_24598,N_24191);
or U25857 (N_25857,N_24449,N_24096);
nor U25858 (N_25858,N_24533,N_24466);
and U25859 (N_25859,N_25002,N_24842);
nor U25860 (N_25860,N_24332,N_24306);
or U25861 (N_25861,N_24922,N_24941);
and U25862 (N_25862,N_25076,N_24841);
and U25863 (N_25863,N_24080,N_24696);
nand U25864 (N_25864,N_24301,N_24559);
and U25865 (N_25865,N_24052,N_24281);
nor U25866 (N_25866,N_24067,N_24726);
nand U25867 (N_25867,N_24058,N_25057);
or U25868 (N_25868,N_24339,N_24472);
or U25869 (N_25869,N_24470,N_25121);
or U25870 (N_25870,N_24279,N_25007);
xnor U25871 (N_25871,N_24449,N_24776);
nor U25872 (N_25872,N_24026,N_24340);
or U25873 (N_25873,N_24700,N_24486);
xnor U25874 (N_25874,N_25115,N_24048);
nand U25875 (N_25875,N_24148,N_24372);
and U25876 (N_25876,N_24658,N_24963);
nand U25877 (N_25877,N_24745,N_24379);
nor U25878 (N_25878,N_24424,N_24669);
nor U25879 (N_25879,N_24446,N_25055);
xnor U25880 (N_25880,N_24106,N_24102);
nor U25881 (N_25881,N_24711,N_24905);
nand U25882 (N_25882,N_24885,N_24539);
nor U25883 (N_25883,N_24340,N_24571);
xnor U25884 (N_25884,N_24178,N_24602);
nand U25885 (N_25885,N_24214,N_24234);
and U25886 (N_25886,N_24682,N_24885);
or U25887 (N_25887,N_24887,N_24996);
nand U25888 (N_25888,N_24792,N_24209);
nand U25889 (N_25889,N_25180,N_25033);
and U25890 (N_25890,N_24303,N_24307);
and U25891 (N_25891,N_24830,N_25157);
xor U25892 (N_25892,N_24585,N_24547);
nor U25893 (N_25893,N_24249,N_25112);
or U25894 (N_25894,N_24586,N_24809);
nand U25895 (N_25895,N_24988,N_24249);
or U25896 (N_25896,N_24241,N_24375);
nor U25897 (N_25897,N_24720,N_25066);
and U25898 (N_25898,N_24257,N_24756);
nand U25899 (N_25899,N_24867,N_24307);
xor U25900 (N_25900,N_24855,N_24380);
and U25901 (N_25901,N_24806,N_24161);
nand U25902 (N_25902,N_25034,N_24570);
nor U25903 (N_25903,N_25096,N_24495);
nand U25904 (N_25904,N_24609,N_24093);
xnor U25905 (N_25905,N_25094,N_24344);
or U25906 (N_25906,N_24621,N_24833);
or U25907 (N_25907,N_24623,N_24594);
and U25908 (N_25908,N_24310,N_24087);
or U25909 (N_25909,N_25188,N_24054);
or U25910 (N_25910,N_25159,N_24452);
nor U25911 (N_25911,N_24524,N_24408);
or U25912 (N_25912,N_24179,N_25163);
or U25913 (N_25913,N_24338,N_25046);
or U25914 (N_25914,N_24829,N_24547);
nor U25915 (N_25915,N_24251,N_24512);
nor U25916 (N_25916,N_24653,N_24825);
and U25917 (N_25917,N_24237,N_25146);
and U25918 (N_25918,N_24209,N_24249);
and U25919 (N_25919,N_24210,N_24259);
nand U25920 (N_25920,N_24467,N_25113);
xor U25921 (N_25921,N_24395,N_25170);
nand U25922 (N_25922,N_24618,N_24013);
nor U25923 (N_25923,N_24443,N_24250);
xnor U25924 (N_25924,N_24797,N_24509);
nand U25925 (N_25925,N_24639,N_24336);
nand U25926 (N_25926,N_25056,N_24751);
or U25927 (N_25927,N_24442,N_24238);
nand U25928 (N_25928,N_24680,N_24760);
and U25929 (N_25929,N_24177,N_25188);
or U25930 (N_25930,N_24346,N_24184);
nor U25931 (N_25931,N_24820,N_24177);
nand U25932 (N_25932,N_24962,N_24060);
xnor U25933 (N_25933,N_25079,N_24886);
or U25934 (N_25934,N_24609,N_25052);
and U25935 (N_25935,N_24010,N_24630);
xor U25936 (N_25936,N_24450,N_24589);
and U25937 (N_25937,N_24110,N_24721);
nand U25938 (N_25938,N_24620,N_24610);
or U25939 (N_25939,N_24422,N_25185);
nand U25940 (N_25940,N_24601,N_25140);
or U25941 (N_25941,N_24765,N_24009);
or U25942 (N_25942,N_24125,N_24304);
and U25943 (N_25943,N_25114,N_24959);
xnor U25944 (N_25944,N_24450,N_25038);
and U25945 (N_25945,N_24884,N_24043);
and U25946 (N_25946,N_24247,N_24647);
and U25947 (N_25947,N_24550,N_24272);
or U25948 (N_25948,N_24889,N_24732);
nor U25949 (N_25949,N_24588,N_24052);
nor U25950 (N_25950,N_24050,N_25038);
nor U25951 (N_25951,N_24542,N_25041);
nand U25952 (N_25952,N_24562,N_24481);
xnor U25953 (N_25953,N_24313,N_25137);
nor U25954 (N_25954,N_24034,N_24046);
or U25955 (N_25955,N_24637,N_24933);
nand U25956 (N_25956,N_24931,N_24279);
nand U25957 (N_25957,N_24804,N_24466);
and U25958 (N_25958,N_24036,N_25166);
nand U25959 (N_25959,N_24632,N_25197);
and U25960 (N_25960,N_24206,N_24096);
nand U25961 (N_25961,N_25139,N_24584);
or U25962 (N_25962,N_24780,N_25148);
nor U25963 (N_25963,N_24721,N_24532);
nand U25964 (N_25964,N_24370,N_24979);
nand U25965 (N_25965,N_24223,N_24017);
or U25966 (N_25966,N_24603,N_24748);
xnor U25967 (N_25967,N_24758,N_24959);
xnor U25968 (N_25968,N_25172,N_24599);
xnor U25969 (N_25969,N_25180,N_24907);
or U25970 (N_25970,N_24618,N_24758);
or U25971 (N_25971,N_24087,N_25044);
or U25972 (N_25972,N_24934,N_25105);
nand U25973 (N_25973,N_24045,N_24150);
or U25974 (N_25974,N_24359,N_24573);
or U25975 (N_25975,N_24851,N_24340);
xnor U25976 (N_25976,N_24924,N_24867);
or U25977 (N_25977,N_24946,N_24817);
or U25978 (N_25978,N_24385,N_25193);
or U25979 (N_25979,N_24288,N_24202);
nor U25980 (N_25980,N_24573,N_24559);
and U25981 (N_25981,N_24467,N_24974);
xnor U25982 (N_25982,N_24625,N_24998);
nand U25983 (N_25983,N_24149,N_24053);
and U25984 (N_25984,N_24554,N_24483);
or U25985 (N_25985,N_25191,N_24260);
nor U25986 (N_25986,N_24718,N_24248);
nand U25987 (N_25987,N_24355,N_24738);
or U25988 (N_25988,N_24341,N_24910);
xnor U25989 (N_25989,N_24269,N_24118);
and U25990 (N_25990,N_24762,N_24094);
nor U25991 (N_25991,N_24028,N_24420);
or U25992 (N_25992,N_24718,N_24986);
nand U25993 (N_25993,N_24407,N_25183);
and U25994 (N_25994,N_24700,N_25163);
nor U25995 (N_25995,N_24151,N_24616);
and U25996 (N_25996,N_24507,N_24957);
xor U25997 (N_25997,N_24192,N_24016);
or U25998 (N_25998,N_25116,N_24856);
xor U25999 (N_25999,N_25106,N_24623);
nor U26000 (N_26000,N_24439,N_24927);
or U26001 (N_26001,N_25180,N_24409);
or U26002 (N_26002,N_24368,N_24911);
nor U26003 (N_26003,N_25040,N_25031);
or U26004 (N_26004,N_24841,N_24933);
and U26005 (N_26005,N_24824,N_24143);
xor U26006 (N_26006,N_24275,N_24895);
nor U26007 (N_26007,N_24694,N_25031);
xor U26008 (N_26008,N_25188,N_24753);
xor U26009 (N_26009,N_24843,N_24951);
xor U26010 (N_26010,N_24665,N_24798);
and U26011 (N_26011,N_25079,N_24847);
xor U26012 (N_26012,N_25084,N_24449);
nor U26013 (N_26013,N_24489,N_24915);
xnor U26014 (N_26014,N_25002,N_24963);
xnor U26015 (N_26015,N_24760,N_25109);
xor U26016 (N_26016,N_25041,N_24061);
nand U26017 (N_26017,N_24266,N_24943);
xnor U26018 (N_26018,N_24863,N_24424);
xnor U26019 (N_26019,N_24178,N_24475);
or U26020 (N_26020,N_24860,N_24959);
and U26021 (N_26021,N_25182,N_24623);
and U26022 (N_26022,N_24485,N_24534);
or U26023 (N_26023,N_24014,N_24943);
and U26024 (N_26024,N_24294,N_24710);
nand U26025 (N_26025,N_24728,N_24977);
and U26026 (N_26026,N_24886,N_24286);
and U26027 (N_26027,N_24584,N_24960);
nor U26028 (N_26028,N_24679,N_24462);
xnor U26029 (N_26029,N_24487,N_24358);
and U26030 (N_26030,N_24618,N_24933);
nand U26031 (N_26031,N_24289,N_24543);
and U26032 (N_26032,N_25096,N_24164);
nand U26033 (N_26033,N_24968,N_25002);
xnor U26034 (N_26034,N_24613,N_24692);
or U26035 (N_26035,N_24959,N_24545);
or U26036 (N_26036,N_24672,N_25017);
or U26037 (N_26037,N_24945,N_24986);
xnor U26038 (N_26038,N_24045,N_24795);
nor U26039 (N_26039,N_24354,N_24227);
xor U26040 (N_26040,N_24871,N_24176);
nand U26041 (N_26041,N_24924,N_24435);
nor U26042 (N_26042,N_24865,N_24524);
nand U26043 (N_26043,N_24267,N_24344);
or U26044 (N_26044,N_24885,N_25077);
xor U26045 (N_26045,N_24038,N_24133);
or U26046 (N_26046,N_24862,N_24662);
xnor U26047 (N_26047,N_24403,N_24276);
and U26048 (N_26048,N_24573,N_25046);
and U26049 (N_26049,N_24318,N_24892);
and U26050 (N_26050,N_24899,N_24322);
nand U26051 (N_26051,N_24575,N_24301);
nand U26052 (N_26052,N_24944,N_24325);
xor U26053 (N_26053,N_24741,N_24751);
and U26054 (N_26054,N_24188,N_25156);
nand U26055 (N_26055,N_24509,N_25054);
xnor U26056 (N_26056,N_24705,N_24998);
and U26057 (N_26057,N_24420,N_24401);
nand U26058 (N_26058,N_24977,N_24724);
and U26059 (N_26059,N_24432,N_24299);
nor U26060 (N_26060,N_24975,N_24996);
or U26061 (N_26061,N_24448,N_24796);
or U26062 (N_26062,N_24327,N_24526);
or U26063 (N_26063,N_24254,N_24365);
or U26064 (N_26064,N_24177,N_24331);
or U26065 (N_26065,N_24211,N_25067);
and U26066 (N_26066,N_25190,N_24774);
or U26067 (N_26067,N_24459,N_24392);
nor U26068 (N_26068,N_24897,N_25158);
xor U26069 (N_26069,N_24486,N_25146);
nor U26070 (N_26070,N_25112,N_24507);
nand U26071 (N_26071,N_25060,N_25012);
and U26072 (N_26072,N_24958,N_24282);
nand U26073 (N_26073,N_24797,N_24144);
and U26074 (N_26074,N_24951,N_25056);
and U26075 (N_26075,N_24624,N_24211);
nor U26076 (N_26076,N_24936,N_24194);
nand U26077 (N_26077,N_24048,N_24160);
and U26078 (N_26078,N_24154,N_24719);
nand U26079 (N_26079,N_24554,N_24678);
xnor U26080 (N_26080,N_24316,N_25068);
nor U26081 (N_26081,N_24820,N_24660);
xor U26082 (N_26082,N_24511,N_24142);
nor U26083 (N_26083,N_24416,N_24468);
nor U26084 (N_26084,N_24755,N_24673);
xnor U26085 (N_26085,N_25068,N_24235);
or U26086 (N_26086,N_24181,N_25110);
nand U26087 (N_26087,N_24694,N_24639);
nand U26088 (N_26088,N_24358,N_24850);
nor U26089 (N_26089,N_24960,N_24810);
nor U26090 (N_26090,N_24705,N_24727);
and U26091 (N_26091,N_24883,N_24647);
nor U26092 (N_26092,N_24634,N_24840);
and U26093 (N_26093,N_24385,N_24152);
nor U26094 (N_26094,N_25143,N_24103);
xnor U26095 (N_26095,N_24876,N_24566);
nand U26096 (N_26096,N_24668,N_24843);
xnor U26097 (N_26097,N_24410,N_24826);
nand U26098 (N_26098,N_24210,N_24825);
nor U26099 (N_26099,N_24439,N_24724);
nor U26100 (N_26100,N_24931,N_24683);
nor U26101 (N_26101,N_24283,N_24770);
or U26102 (N_26102,N_25190,N_24464);
nand U26103 (N_26103,N_24040,N_24098);
nor U26104 (N_26104,N_24625,N_24587);
nor U26105 (N_26105,N_24507,N_24722);
or U26106 (N_26106,N_24424,N_24484);
nor U26107 (N_26107,N_24822,N_24466);
or U26108 (N_26108,N_25064,N_24395);
or U26109 (N_26109,N_25198,N_24872);
xor U26110 (N_26110,N_25166,N_25156);
and U26111 (N_26111,N_24540,N_24763);
or U26112 (N_26112,N_24944,N_25075);
and U26113 (N_26113,N_24813,N_24877);
nand U26114 (N_26114,N_25054,N_24921);
nand U26115 (N_26115,N_24131,N_24337);
nor U26116 (N_26116,N_24566,N_24111);
xor U26117 (N_26117,N_24349,N_24584);
nor U26118 (N_26118,N_24680,N_25116);
nand U26119 (N_26119,N_25135,N_24806);
and U26120 (N_26120,N_24168,N_24595);
nor U26121 (N_26121,N_25130,N_25034);
xnor U26122 (N_26122,N_24683,N_24315);
xor U26123 (N_26123,N_24561,N_24042);
and U26124 (N_26124,N_24089,N_24852);
xor U26125 (N_26125,N_24293,N_24634);
nor U26126 (N_26126,N_24734,N_25144);
nand U26127 (N_26127,N_24282,N_25180);
nor U26128 (N_26128,N_24063,N_25139);
and U26129 (N_26129,N_24657,N_24998);
and U26130 (N_26130,N_24934,N_24079);
and U26131 (N_26131,N_24134,N_24651);
nor U26132 (N_26132,N_24843,N_24764);
nor U26133 (N_26133,N_24802,N_24638);
and U26134 (N_26134,N_24173,N_24256);
nand U26135 (N_26135,N_24130,N_24929);
and U26136 (N_26136,N_24399,N_24207);
and U26137 (N_26137,N_24834,N_24704);
or U26138 (N_26138,N_24600,N_24792);
and U26139 (N_26139,N_24868,N_25156);
nand U26140 (N_26140,N_24756,N_24721);
or U26141 (N_26141,N_24509,N_24914);
and U26142 (N_26142,N_24486,N_24196);
and U26143 (N_26143,N_24388,N_24735);
or U26144 (N_26144,N_24514,N_24898);
nor U26145 (N_26145,N_24415,N_24096);
or U26146 (N_26146,N_24461,N_24646);
nor U26147 (N_26147,N_24483,N_24398);
and U26148 (N_26148,N_25049,N_24873);
nand U26149 (N_26149,N_25087,N_25152);
nor U26150 (N_26150,N_24961,N_24089);
nand U26151 (N_26151,N_24193,N_24593);
or U26152 (N_26152,N_25100,N_24865);
and U26153 (N_26153,N_24290,N_25183);
and U26154 (N_26154,N_24525,N_24126);
or U26155 (N_26155,N_25047,N_24474);
nand U26156 (N_26156,N_24550,N_25107);
nand U26157 (N_26157,N_25065,N_24379);
or U26158 (N_26158,N_24198,N_24813);
nor U26159 (N_26159,N_25121,N_25123);
nor U26160 (N_26160,N_24174,N_24797);
xnor U26161 (N_26161,N_24626,N_24371);
or U26162 (N_26162,N_25180,N_24941);
and U26163 (N_26163,N_24043,N_24560);
nor U26164 (N_26164,N_24701,N_24839);
nand U26165 (N_26165,N_24455,N_25053);
and U26166 (N_26166,N_24803,N_24479);
nand U26167 (N_26167,N_24496,N_24642);
and U26168 (N_26168,N_24197,N_25192);
and U26169 (N_26169,N_25020,N_24101);
xor U26170 (N_26170,N_24198,N_24493);
nand U26171 (N_26171,N_24983,N_24582);
nand U26172 (N_26172,N_25070,N_24798);
xnor U26173 (N_26173,N_24446,N_24439);
nor U26174 (N_26174,N_24800,N_24821);
xnor U26175 (N_26175,N_24938,N_24867);
xnor U26176 (N_26176,N_24113,N_24635);
and U26177 (N_26177,N_24719,N_24692);
nand U26178 (N_26178,N_24845,N_24215);
nand U26179 (N_26179,N_24980,N_25136);
and U26180 (N_26180,N_24988,N_24759);
nor U26181 (N_26181,N_24491,N_24223);
nand U26182 (N_26182,N_24202,N_24807);
or U26183 (N_26183,N_24547,N_24652);
or U26184 (N_26184,N_24359,N_24781);
and U26185 (N_26185,N_25015,N_24896);
xnor U26186 (N_26186,N_25141,N_24265);
nor U26187 (N_26187,N_24754,N_24147);
xnor U26188 (N_26188,N_25094,N_24351);
xnor U26189 (N_26189,N_24196,N_24745);
nor U26190 (N_26190,N_24513,N_24711);
nor U26191 (N_26191,N_24384,N_24696);
and U26192 (N_26192,N_24379,N_24313);
or U26193 (N_26193,N_24260,N_24062);
nand U26194 (N_26194,N_24072,N_24110);
nand U26195 (N_26195,N_24415,N_24566);
or U26196 (N_26196,N_24097,N_24054);
xnor U26197 (N_26197,N_24480,N_25117);
xor U26198 (N_26198,N_25076,N_25088);
and U26199 (N_26199,N_24222,N_24627);
nor U26200 (N_26200,N_24821,N_24090);
nor U26201 (N_26201,N_25001,N_24956);
nor U26202 (N_26202,N_24023,N_24254);
nor U26203 (N_26203,N_24411,N_24285);
xnor U26204 (N_26204,N_24507,N_24573);
or U26205 (N_26205,N_24291,N_24823);
nand U26206 (N_26206,N_24471,N_24564);
and U26207 (N_26207,N_24235,N_25158);
nand U26208 (N_26208,N_24862,N_24114);
xor U26209 (N_26209,N_25039,N_24583);
or U26210 (N_26210,N_24183,N_24492);
nor U26211 (N_26211,N_24370,N_24501);
nor U26212 (N_26212,N_24975,N_24030);
or U26213 (N_26213,N_24954,N_24487);
or U26214 (N_26214,N_24820,N_24651);
or U26215 (N_26215,N_24476,N_24148);
or U26216 (N_26216,N_25081,N_24724);
nor U26217 (N_26217,N_24256,N_24376);
or U26218 (N_26218,N_25110,N_24316);
and U26219 (N_26219,N_24382,N_25057);
xor U26220 (N_26220,N_24673,N_24682);
nand U26221 (N_26221,N_24545,N_24397);
or U26222 (N_26222,N_24837,N_24004);
nand U26223 (N_26223,N_24839,N_24657);
xnor U26224 (N_26224,N_24328,N_24804);
or U26225 (N_26225,N_24245,N_24559);
nor U26226 (N_26226,N_24936,N_24038);
nand U26227 (N_26227,N_24324,N_24873);
nand U26228 (N_26228,N_24371,N_24955);
nor U26229 (N_26229,N_24906,N_24670);
xor U26230 (N_26230,N_24322,N_24513);
nor U26231 (N_26231,N_24625,N_24704);
xor U26232 (N_26232,N_24898,N_24409);
and U26233 (N_26233,N_24896,N_24906);
nand U26234 (N_26234,N_24980,N_24604);
nand U26235 (N_26235,N_24886,N_24712);
nor U26236 (N_26236,N_24621,N_24765);
or U26237 (N_26237,N_24330,N_24728);
or U26238 (N_26238,N_25053,N_24165);
nor U26239 (N_26239,N_24862,N_24808);
nor U26240 (N_26240,N_25194,N_25079);
and U26241 (N_26241,N_24589,N_24634);
nand U26242 (N_26242,N_24042,N_24823);
or U26243 (N_26243,N_24760,N_24004);
nand U26244 (N_26244,N_24806,N_24559);
or U26245 (N_26245,N_24753,N_24365);
nand U26246 (N_26246,N_24135,N_24050);
nand U26247 (N_26247,N_24364,N_24701);
or U26248 (N_26248,N_24858,N_24647);
xnor U26249 (N_26249,N_24279,N_25070);
or U26250 (N_26250,N_24884,N_25173);
xnor U26251 (N_26251,N_24685,N_25056);
or U26252 (N_26252,N_24033,N_24426);
or U26253 (N_26253,N_24822,N_24656);
and U26254 (N_26254,N_25180,N_24089);
and U26255 (N_26255,N_24034,N_24397);
nor U26256 (N_26256,N_25167,N_24399);
nand U26257 (N_26257,N_24783,N_24035);
nand U26258 (N_26258,N_24755,N_24813);
or U26259 (N_26259,N_24572,N_24408);
nor U26260 (N_26260,N_24105,N_24827);
nand U26261 (N_26261,N_24282,N_24091);
nand U26262 (N_26262,N_24443,N_24337);
xor U26263 (N_26263,N_25064,N_24865);
or U26264 (N_26264,N_24199,N_24331);
nand U26265 (N_26265,N_24013,N_25186);
nand U26266 (N_26266,N_24080,N_24754);
and U26267 (N_26267,N_24894,N_25171);
nor U26268 (N_26268,N_24414,N_24837);
or U26269 (N_26269,N_24850,N_24166);
nor U26270 (N_26270,N_24975,N_24286);
nand U26271 (N_26271,N_24689,N_24598);
nand U26272 (N_26272,N_25032,N_24567);
or U26273 (N_26273,N_24903,N_25119);
and U26274 (N_26274,N_25162,N_24644);
or U26275 (N_26275,N_25143,N_24942);
xor U26276 (N_26276,N_24768,N_25034);
nor U26277 (N_26277,N_24867,N_25128);
and U26278 (N_26278,N_24941,N_24450);
and U26279 (N_26279,N_25106,N_24714);
nor U26280 (N_26280,N_24580,N_25067);
and U26281 (N_26281,N_24395,N_24383);
or U26282 (N_26282,N_24584,N_24660);
xor U26283 (N_26283,N_24787,N_24828);
xor U26284 (N_26284,N_24531,N_25193);
xor U26285 (N_26285,N_24439,N_25030);
xnor U26286 (N_26286,N_24999,N_24909);
and U26287 (N_26287,N_25098,N_24789);
xnor U26288 (N_26288,N_24964,N_24943);
xnor U26289 (N_26289,N_24343,N_24909);
xnor U26290 (N_26290,N_25042,N_24016);
and U26291 (N_26291,N_24186,N_25167);
and U26292 (N_26292,N_24137,N_24369);
or U26293 (N_26293,N_24181,N_24246);
or U26294 (N_26294,N_25122,N_24309);
nor U26295 (N_26295,N_24245,N_24843);
nand U26296 (N_26296,N_24367,N_24180);
or U26297 (N_26297,N_24290,N_24464);
nor U26298 (N_26298,N_25184,N_24642);
xor U26299 (N_26299,N_24339,N_24808);
nand U26300 (N_26300,N_24008,N_25036);
or U26301 (N_26301,N_24987,N_24657);
nand U26302 (N_26302,N_24285,N_24088);
xnor U26303 (N_26303,N_24793,N_25132);
nand U26304 (N_26304,N_24932,N_24005);
and U26305 (N_26305,N_24040,N_24123);
and U26306 (N_26306,N_24531,N_25066);
or U26307 (N_26307,N_24865,N_25172);
and U26308 (N_26308,N_24917,N_24211);
and U26309 (N_26309,N_24940,N_24925);
and U26310 (N_26310,N_24394,N_24888);
or U26311 (N_26311,N_24872,N_24122);
and U26312 (N_26312,N_24535,N_24883);
nand U26313 (N_26313,N_24728,N_24363);
or U26314 (N_26314,N_24415,N_24832);
and U26315 (N_26315,N_24091,N_24729);
nand U26316 (N_26316,N_24621,N_24131);
xnor U26317 (N_26317,N_24395,N_24431);
nand U26318 (N_26318,N_24563,N_24379);
nand U26319 (N_26319,N_24238,N_24588);
and U26320 (N_26320,N_24189,N_24535);
nand U26321 (N_26321,N_25054,N_24267);
xor U26322 (N_26322,N_24995,N_24213);
xor U26323 (N_26323,N_24031,N_24373);
nor U26324 (N_26324,N_24638,N_25034);
and U26325 (N_26325,N_24516,N_24466);
xor U26326 (N_26326,N_24083,N_24799);
nor U26327 (N_26327,N_24142,N_24390);
and U26328 (N_26328,N_24165,N_24852);
nor U26329 (N_26329,N_24846,N_24339);
or U26330 (N_26330,N_24320,N_24319);
and U26331 (N_26331,N_24469,N_24352);
xor U26332 (N_26332,N_24409,N_24142);
nor U26333 (N_26333,N_24675,N_24432);
xor U26334 (N_26334,N_24413,N_24659);
nand U26335 (N_26335,N_24694,N_24552);
and U26336 (N_26336,N_24295,N_24182);
nor U26337 (N_26337,N_24388,N_24045);
nand U26338 (N_26338,N_24054,N_24926);
and U26339 (N_26339,N_24256,N_25186);
xnor U26340 (N_26340,N_24083,N_25196);
nand U26341 (N_26341,N_25030,N_24242);
and U26342 (N_26342,N_24158,N_24489);
and U26343 (N_26343,N_24435,N_25150);
nand U26344 (N_26344,N_25011,N_24351);
nand U26345 (N_26345,N_25155,N_24524);
and U26346 (N_26346,N_25010,N_24506);
xor U26347 (N_26347,N_24393,N_24061);
nand U26348 (N_26348,N_24690,N_24147);
and U26349 (N_26349,N_24470,N_25056);
nand U26350 (N_26350,N_24426,N_24474);
nand U26351 (N_26351,N_24401,N_24160);
nor U26352 (N_26352,N_24594,N_25192);
xor U26353 (N_26353,N_24269,N_24957);
or U26354 (N_26354,N_25194,N_24424);
nand U26355 (N_26355,N_24743,N_24828);
and U26356 (N_26356,N_24797,N_24664);
and U26357 (N_26357,N_24710,N_24086);
and U26358 (N_26358,N_24256,N_24877);
nor U26359 (N_26359,N_24943,N_25101);
nor U26360 (N_26360,N_24910,N_24398);
or U26361 (N_26361,N_24013,N_24280);
or U26362 (N_26362,N_24413,N_24431);
or U26363 (N_26363,N_24085,N_24323);
nor U26364 (N_26364,N_24727,N_25192);
or U26365 (N_26365,N_25139,N_24622);
xnor U26366 (N_26366,N_24973,N_25196);
nand U26367 (N_26367,N_24784,N_24079);
or U26368 (N_26368,N_24957,N_24152);
or U26369 (N_26369,N_24863,N_24302);
nor U26370 (N_26370,N_25005,N_24641);
nor U26371 (N_26371,N_25061,N_24106);
xnor U26372 (N_26372,N_25002,N_24444);
xnor U26373 (N_26373,N_24176,N_24241);
or U26374 (N_26374,N_24398,N_25048);
and U26375 (N_26375,N_25162,N_24155);
nand U26376 (N_26376,N_24603,N_24639);
and U26377 (N_26377,N_24508,N_25065);
nor U26378 (N_26378,N_25072,N_24220);
and U26379 (N_26379,N_25014,N_24515);
nor U26380 (N_26380,N_24190,N_25091);
or U26381 (N_26381,N_24179,N_24792);
nor U26382 (N_26382,N_24942,N_24130);
nor U26383 (N_26383,N_24631,N_24603);
and U26384 (N_26384,N_24668,N_25153);
and U26385 (N_26385,N_24992,N_24891);
nor U26386 (N_26386,N_25048,N_24409);
nor U26387 (N_26387,N_24743,N_24779);
nor U26388 (N_26388,N_24969,N_24948);
xnor U26389 (N_26389,N_24972,N_24453);
and U26390 (N_26390,N_24959,N_24676);
and U26391 (N_26391,N_24615,N_24323);
xor U26392 (N_26392,N_25030,N_24780);
or U26393 (N_26393,N_24441,N_24397);
nand U26394 (N_26394,N_24492,N_24765);
or U26395 (N_26395,N_24201,N_24059);
xor U26396 (N_26396,N_24546,N_25112);
or U26397 (N_26397,N_25100,N_24799);
and U26398 (N_26398,N_24417,N_24401);
nor U26399 (N_26399,N_24634,N_24733);
xor U26400 (N_26400,N_25877,N_25999);
xnor U26401 (N_26401,N_26017,N_25384);
xor U26402 (N_26402,N_26334,N_25235);
and U26403 (N_26403,N_25699,N_26300);
xnor U26404 (N_26404,N_26071,N_26099);
or U26405 (N_26405,N_25731,N_26100);
and U26406 (N_26406,N_26356,N_26085);
and U26407 (N_26407,N_25272,N_25471);
or U26408 (N_26408,N_25629,N_26053);
nand U26409 (N_26409,N_25211,N_26113);
nand U26410 (N_26410,N_25212,N_25214);
nand U26411 (N_26411,N_25422,N_25917);
nor U26412 (N_26412,N_25291,N_25777);
xor U26413 (N_26413,N_25279,N_25789);
nor U26414 (N_26414,N_25889,N_25926);
or U26415 (N_26415,N_26149,N_26117);
xnor U26416 (N_26416,N_25319,N_25876);
nor U26417 (N_26417,N_25571,N_25636);
nand U26418 (N_26418,N_26339,N_26175);
nor U26419 (N_26419,N_26010,N_25643);
or U26420 (N_26420,N_26033,N_25770);
nor U26421 (N_26421,N_25537,N_25750);
or U26422 (N_26422,N_25252,N_25732);
nand U26423 (N_26423,N_25897,N_25846);
or U26424 (N_26424,N_26314,N_26170);
xor U26425 (N_26425,N_25254,N_25695);
and U26426 (N_26426,N_25968,N_25485);
or U26427 (N_26427,N_26058,N_25891);
nand U26428 (N_26428,N_25628,N_25826);
xor U26429 (N_26429,N_26063,N_25786);
nand U26430 (N_26430,N_25307,N_26227);
and U26431 (N_26431,N_25317,N_26250);
nand U26432 (N_26432,N_26044,N_26275);
or U26433 (N_26433,N_26026,N_25765);
and U26434 (N_26434,N_25405,N_26056);
nand U26435 (N_26435,N_26179,N_25792);
nor U26436 (N_26436,N_25784,N_25654);
xnor U26437 (N_26437,N_26370,N_26315);
nand U26438 (N_26438,N_25675,N_25218);
or U26439 (N_26439,N_25697,N_26320);
nor U26440 (N_26440,N_25231,N_26125);
nor U26441 (N_26441,N_26341,N_26062);
nand U26442 (N_26442,N_25271,N_26078);
nand U26443 (N_26443,N_25873,N_26245);
or U26444 (N_26444,N_26073,N_26121);
and U26445 (N_26445,N_26309,N_25508);
xor U26446 (N_26446,N_25599,N_25756);
nor U26447 (N_26447,N_25552,N_25812);
nor U26448 (N_26448,N_25386,N_25658);
xnor U26449 (N_26449,N_26131,N_25364);
nand U26450 (N_26450,N_25259,N_25866);
xor U26451 (N_26451,N_25350,N_25443);
nor U26452 (N_26452,N_26292,N_26031);
or U26453 (N_26453,N_26198,N_26304);
nand U26454 (N_26454,N_25389,N_25738);
and U26455 (N_26455,N_25742,N_26182);
xor U26456 (N_26456,N_26301,N_25296);
and U26457 (N_26457,N_26365,N_25703);
and U26458 (N_26458,N_25779,N_26360);
nand U26459 (N_26459,N_26248,N_26258);
and U26460 (N_26460,N_26388,N_25404);
or U26461 (N_26461,N_26393,N_26381);
and U26462 (N_26462,N_26311,N_25817);
or U26463 (N_26463,N_25318,N_26352);
nand U26464 (N_26464,N_25572,N_25514);
xnor U26465 (N_26465,N_26359,N_25990);
or U26466 (N_26466,N_25694,N_25379);
or U26467 (N_26467,N_26016,N_25493);
or U26468 (N_26468,N_25338,N_25544);
and U26469 (N_26469,N_25382,N_26180);
or U26470 (N_26470,N_26181,N_26118);
or U26471 (N_26471,N_26389,N_26174);
or U26472 (N_26472,N_25295,N_25505);
nor U26473 (N_26473,N_25881,N_25400);
and U26474 (N_26474,N_25360,N_25958);
and U26475 (N_26475,N_25700,N_25362);
or U26476 (N_26476,N_26143,N_25258);
or U26477 (N_26477,N_25547,N_25988);
and U26478 (N_26478,N_25676,N_26255);
nor U26479 (N_26479,N_25240,N_26080);
nand U26480 (N_26480,N_25649,N_26355);
nor U26481 (N_26481,N_25455,N_26236);
or U26482 (N_26482,N_25530,N_26338);
and U26483 (N_26483,N_25806,N_25504);
or U26484 (N_26484,N_25913,N_25666);
xnor U26485 (N_26485,N_25322,N_25932);
and U26486 (N_26486,N_26027,N_25783);
xnor U26487 (N_26487,N_26169,N_25767);
or U26488 (N_26488,N_26200,N_25205);
nor U26489 (N_26489,N_25439,N_26270);
and U26490 (N_26490,N_26242,N_26086);
xor U26491 (N_26491,N_25298,N_26251);
nand U26492 (N_26492,N_25527,N_25744);
or U26493 (N_26493,N_25314,N_26142);
xor U26494 (N_26494,N_25287,N_26029);
nand U26495 (N_26495,N_25663,N_25621);
or U26496 (N_26496,N_25626,N_26145);
nand U26497 (N_26497,N_26120,N_25385);
or U26498 (N_26498,N_26244,N_25224);
and U26499 (N_26499,N_25822,N_25936);
xor U26500 (N_26500,N_25850,N_25907);
nand U26501 (N_26501,N_25660,N_25785);
nand U26502 (N_26502,N_25887,N_25466);
nand U26503 (N_26503,N_25664,N_25243);
and U26504 (N_26504,N_25920,N_25661);
or U26505 (N_26505,N_25288,N_26280);
nor U26506 (N_26506,N_26246,N_26018);
or U26507 (N_26507,N_26337,N_26096);
and U26508 (N_26508,N_25332,N_25885);
nor U26509 (N_26509,N_25946,N_26264);
nand U26510 (N_26510,N_25373,N_25994);
or U26511 (N_26511,N_25472,N_26231);
xor U26512 (N_26512,N_25325,N_25462);
xor U26513 (N_26513,N_26165,N_26230);
or U26514 (N_26514,N_25824,N_26290);
and U26515 (N_26515,N_25232,N_25698);
or U26516 (N_26516,N_25359,N_25247);
or U26517 (N_26517,N_25449,N_25239);
and U26518 (N_26518,N_26291,N_25622);
xnor U26519 (N_26519,N_25509,N_25925);
xor U26520 (N_26520,N_26005,N_26187);
xor U26521 (N_26521,N_25497,N_26384);
or U26522 (N_26522,N_25667,N_25865);
or U26523 (N_26523,N_26302,N_25375);
nand U26524 (N_26524,N_26235,N_26043);
and U26525 (N_26525,N_25945,N_26303);
or U26526 (N_26526,N_25760,N_25363);
xnor U26527 (N_26527,N_25965,N_26048);
nor U26528 (N_26528,N_26249,N_25982);
and U26529 (N_26529,N_26276,N_25816);
nand U26530 (N_26530,N_26067,N_25450);
nor U26531 (N_26531,N_25486,N_25969);
xnor U26532 (N_26532,N_26011,N_25774);
or U26533 (N_26533,N_25949,N_25975);
or U26534 (N_26534,N_25955,N_25627);
nor U26535 (N_26535,N_25202,N_25559);
or U26536 (N_26536,N_25430,N_25499);
nor U26537 (N_26537,N_25226,N_26069);
nor U26538 (N_26538,N_25294,N_25457);
nor U26539 (N_26539,N_25733,N_26003);
xor U26540 (N_26540,N_26344,N_26247);
or U26541 (N_26541,N_25707,N_25903);
and U26542 (N_26542,N_25345,N_26329);
nand U26543 (N_26543,N_25267,N_25227);
nand U26544 (N_26544,N_25365,N_25281);
and U26545 (N_26545,N_25619,N_25483);
or U26546 (N_26546,N_25591,N_26277);
nand U26547 (N_26547,N_25854,N_25396);
nand U26548 (N_26548,N_25321,N_25584);
or U26549 (N_26549,N_26177,N_25432);
or U26550 (N_26550,N_25401,N_26188);
nor U26551 (N_26551,N_25723,N_26195);
xor U26552 (N_26552,N_25574,N_25358);
nor U26553 (N_26553,N_25724,N_26133);
and U26554 (N_26554,N_25280,N_25650);
and U26555 (N_26555,N_25573,N_25800);
or U26556 (N_26556,N_25640,N_25519);
and U26557 (N_26557,N_26036,N_25894);
nand U26558 (N_26558,N_25589,N_25753);
nor U26559 (N_26559,N_25392,N_25919);
nor U26560 (N_26560,N_26295,N_26317);
nor U26561 (N_26561,N_26353,N_25613);
nor U26562 (N_26562,N_25554,N_26183);
or U26563 (N_26563,N_25778,N_25859);
xnor U26564 (N_26564,N_25209,N_25904);
or U26565 (N_26565,N_26094,N_26112);
or U26566 (N_26566,N_26054,N_26111);
nor U26567 (N_26567,N_26345,N_25905);
nor U26568 (N_26568,N_25938,N_26367);
and U26569 (N_26569,N_25306,N_26268);
xor U26570 (N_26570,N_26101,N_25704);
and U26571 (N_26571,N_26382,N_25830);
and U26572 (N_26572,N_25569,N_26077);
nor U26573 (N_26573,N_25266,N_25371);
nand U26574 (N_26574,N_25293,N_25701);
and U26575 (N_26575,N_25470,N_25997);
or U26576 (N_26576,N_26226,N_25839);
nand U26577 (N_26577,N_25270,N_25869);
and U26578 (N_26578,N_25313,N_25334);
nand U26579 (N_26579,N_25229,N_26399);
xor U26580 (N_26580,N_26283,N_26252);
xnor U26581 (N_26581,N_25217,N_26202);
nor U26582 (N_26582,N_25335,N_25407);
nor U26583 (N_26583,N_25683,N_25542);
and U26584 (N_26584,N_25568,N_26066);
nor U26585 (N_26585,N_25290,N_25617);
nand U26586 (N_26586,N_26013,N_25503);
xnor U26587 (N_26587,N_25600,N_26284);
nand U26588 (N_26588,N_25529,N_25441);
nand U26589 (N_26589,N_26278,N_25987);
nor U26590 (N_26590,N_26137,N_26162);
nand U26591 (N_26591,N_25951,N_25838);
and U26592 (N_26592,N_26271,N_25981);
or U26593 (N_26593,N_25608,N_25299);
xor U26594 (N_26594,N_26070,N_26164);
nand U26595 (N_26595,N_25459,N_26241);
xnor U26596 (N_26596,N_26342,N_26158);
or U26597 (N_26597,N_25448,N_26260);
and U26598 (N_26598,N_25525,N_25856);
xor U26599 (N_26599,N_25870,N_26316);
and U26600 (N_26600,N_25603,N_25347);
nor U26601 (N_26601,N_25934,N_25840);
nor U26602 (N_26602,N_25394,N_25312);
nand U26603 (N_26603,N_25357,N_25984);
nand U26604 (N_26604,N_26343,N_26037);
nor U26605 (N_26605,N_25346,N_25727);
nand U26606 (N_26606,N_25581,N_26377);
and U26607 (N_26607,N_25369,N_26034);
nor U26608 (N_26608,N_26197,N_25353);
nand U26609 (N_26609,N_25549,N_26108);
or U26610 (N_26610,N_25688,N_25341);
or U26611 (N_26611,N_25630,N_25620);
or U26612 (N_26612,N_25759,N_25370);
and U26613 (N_26613,N_25853,N_26153);
or U26614 (N_26614,N_25673,N_25921);
or U26615 (N_26615,N_25849,N_25625);
nor U26616 (N_26616,N_25219,N_25234);
or U26617 (N_26617,N_26322,N_26259);
nand U26618 (N_26618,N_25745,N_25842);
or U26619 (N_26619,N_25883,N_25241);
and U26620 (N_26620,N_25397,N_26239);
xnor U26621 (N_26621,N_26361,N_25526);
xnor U26622 (N_26622,N_25912,N_26354);
nor U26623 (N_26623,N_25828,N_26084);
nor U26624 (N_26624,N_25693,N_26104);
nand U26625 (N_26625,N_26055,N_25749);
and U26626 (N_26626,N_26233,N_26256);
nand U26627 (N_26627,N_25606,N_25751);
nand U26628 (N_26628,N_26079,N_25893);
or U26629 (N_26629,N_26293,N_25875);
and U26630 (N_26630,N_25425,N_26038);
xnor U26631 (N_26631,N_25300,N_25825);
or U26632 (N_26632,N_25539,N_26159);
nand U26633 (N_26633,N_26046,N_25413);
nand U26634 (N_26634,N_25278,N_25222);
nand U26635 (N_26635,N_26385,N_26193);
or U26636 (N_26636,N_25930,N_25916);
or U26637 (N_26637,N_26088,N_26160);
xnor U26638 (N_26638,N_25680,N_26000);
and U26639 (N_26639,N_26220,N_25478);
nand U26640 (N_26640,N_25808,N_25395);
and U26641 (N_26641,N_26081,N_25705);
xnor U26642 (N_26642,N_25948,N_25467);
and U26643 (N_26643,N_25769,N_26152);
or U26644 (N_26644,N_25431,N_25316);
nor U26645 (N_26645,N_25845,N_25378);
or U26646 (N_26646,N_25655,N_25924);
nand U26647 (N_26647,N_25538,N_25811);
nor U26648 (N_26648,N_26391,N_25766);
nor U26649 (N_26649,N_25343,N_25858);
xor U26650 (N_26650,N_26171,N_25900);
nor U26651 (N_26651,N_26068,N_26082);
nor U26652 (N_26652,N_25922,N_25669);
nor U26653 (N_26653,N_26306,N_25420);
nor U26654 (N_26654,N_25297,N_25273);
and U26655 (N_26655,N_25755,N_25963);
xor U26656 (N_26656,N_25253,N_26379);
nor U26657 (N_26657,N_25292,N_26190);
xor U26658 (N_26658,N_25793,N_26281);
xor U26659 (N_26659,N_26098,N_25479);
and U26660 (N_26660,N_26138,N_26051);
or U26661 (N_26661,N_25444,N_25960);
nor U26662 (N_26662,N_25412,N_25996);
and U26663 (N_26663,N_25943,N_25595);
nand U26664 (N_26664,N_26115,N_25713);
or U26665 (N_26665,N_26285,N_26299);
xor U26666 (N_26666,N_26228,N_25635);
xnor U26667 (N_26667,N_25532,N_25377);
xnor U26668 (N_26668,N_26206,N_25477);
nor U26669 (N_26669,N_26330,N_26185);
nor U26670 (N_26670,N_25860,N_25427);
xor U26671 (N_26671,N_26254,N_26340);
or U26672 (N_26672,N_25484,N_25237);
nand U26673 (N_26673,N_26363,N_25668);
and U26674 (N_26674,N_25788,N_25607);
nor U26675 (N_26675,N_25631,N_25686);
nand U26676 (N_26676,N_26097,N_26229);
nand U26677 (N_26677,N_25764,N_25367);
nand U26678 (N_26678,N_25515,N_25458);
nand U26679 (N_26679,N_26168,N_25349);
xor U26680 (N_26680,N_26176,N_25594);
and U26681 (N_26681,N_25843,N_25415);
and U26682 (N_26682,N_25524,N_25787);
and U26683 (N_26683,N_26023,N_25414);
xnor U26684 (N_26684,N_25593,N_25993);
or U26685 (N_26685,N_25953,N_25895);
nor U26686 (N_26686,N_25940,N_25440);
and U26687 (N_26687,N_25548,N_25762);
xor U26688 (N_26688,N_25339,N_26074);
nor U26689 (N_26689,N_26321,N_25588);
xor U26690 (N_26690,N_26147,N_25671);
or U26691 (N_26691,N_26007,N_25248);
or U26692 (N_26692,N_25952,N_26394);
and U26693 (N_26693,N_25225,N_25761);
nand U26694 (N_26694,N_26167,N_26201);
nand U26695 (N_26695,N_25864,N_25565);
nand U26696 (N_26696,N_26144,N_25327);
nand U26697 (N_26697,N_25399,N_25383);
nand U26698 (N_26698,N_25429,N_25475);
and U26699 (N_26699,N_25374,N_25637);
nand U26700 (N_26700,N_25329,N_25402);
nand U26701 (N_26701,N_25714,N_25657);
xnor U26702 (N_26702,N_26154,N_25550);
and U26703 (N_26703,N_26217,N_26375);
nand U26704 (N_26704,N_26265,N_25433);
or U26705 (N_26705,N_25391,N_25735);
and U26706 (N_26706,N_25268,N_26150);
or U26707 (N_26707,N_25465,N_25496);
or U26708 (N_26708,N_25301,N_26061);
and U26709 (N_26709,N_26312,N_25692);
and U26710 (N_26710,N_25545,N_26351);
xnor U26711 (N_26711,N_26323,N_25791);
or U26712 (N_26712,N_25957,N_25721);
xnor U26713 (N_26713,N_25715,N_25973);
nand U26714 (N_26714,N_25336,N_25330);
xor U26715 (N_26715,N_25265,N_25555);
or U26716 (N_26716,N_26273,N_25685);
nand U26717 (N_26717,N_25743,N_25421);
nor U26718 (N_26718,N_25909,N_25315);
xnor U26719 (N_26719,N_25653,N_25390);
and U26720 (N_26720,N_26136,N_26274);
nor U26721 (N_26721,N_25618,N_26040);
nor U26722 (N_26722,N_25827,N_25469);
or U26723 (N_26723,N_25736,N_25602);
or U26724 (N_26724,N_25690,N_25203);
nand U26725 (N_26725,N_25795,N_25340);
and U26726 (N_26726,N_25255,N_26199);
nor U26727 (N_26727,N_25481,N_25566);
and U26728 (N_26728,N_26373,N_26376);
or U26729 (N_26729,N_25983,N_26173);
nor U26730 (N_26730,N_25651,N_25771);
nor U26731 (N_26731,N_25490,N_26269);
and U26732 (N_26732,N_25644,N_25416);
or U26733 (N_26733,N_25236,N_26024);
and U26734 (N_26734,N_26395,N_26127);
or U26735 (N_26735,N_25614,N_25763);
nor U26736 (N_26736,N_25546,N_25473);
or U26737 (N_26737,N_26272,N_25906);
and U26738 (N_26738,N_25815,N_25516);
and U26739 (N_26739,N_25342,N_26155);
xnor U26740 (N_26740,N_26090,N_25977);
and U26741 (N_26741,N_25564,N_26189);
or U26742 (N_26742,N_26124,N_25276);
xnor U26743 (N_26743,N_25747,N_26119);
xor U26744 (N_26744,N_25634,N_25813);
or U26745 (N_26745,N_25797,N_25890);
nand U26746 (N_26746,N_25985,N_26042);
nor U26747 (N_26747,N_26093,N_25451);
xnor U26748 (N_26748,N_26207,N_25201);
nor U26749 (N_26749,N_25674,N_26369);
and U26750 (N_26750,N_25752,N_25494);
or U26751 (N_26751,N_25352,N_25204);
nor U26752 (N_26752,N_25935,N_26390);
or U26753 (N_26753,N_26348,N_26065);
and U26754 (N_26754,N_25491,N_25579);
xnor U26755 (N_26755,N_26214,N_25261);
and U26756 (N_26756,N_25944,N_25652);
and U26757 (N_26757,N_26279,N_25615);
nor U26758 (N_26758,N_25523,N_26267);
nand U26759 (N_26759,N_25659,N_25482);
nor U26760 (N_26760,N_25580,N_25512);
and U26761 (N_26761,N_25230,N_25646);
and U26762 (N_26762,N_25739,N_25645);
nor U26763 (N_26763,N_25463,N_25772);
nor U26764 (N_26764,N_25454,N_25452);
and U26765 (N_26765,N_25972,N_25820);
nand U26766 (N_26766,N_25851,N_25711);
xor U26767 (N_26767,N_25289,N_25708);
nand U26768 (N_26768,N_25453,N_25333);
xor U26769 (N_26769,N_26057,N_25689);
or U26770 (N_26770,N_25223,N_25959);
xor U26771 (N_26771,N_25388,N_25956);
or U26772 (N_26772,N_26366,N_25246);
xor U26773 (N_26773,N_25758,N_25709);
xor U26774 (N_26774,N_25801,N_26371);
nand U26775 (N_26775,N_25264,N_25961);
or U26776 (N_26776,N_26151,N_25208);
nor U26777 (N_26777,N_26331,N_26372);
and U26778 (N_26778,N_25601,N_25863);
nor U26779 (N_26779,N_25592,N_26184);
and U26780 (N_26780,N_25302,N_25213);
nor U26781 (N_26781,N_25974,N_25351);
xor U26782 (N_26782,N_25818,N_25563);
and U26783 (N_26783,N_25488,N_25954);
nor U26784 (N_26784,N_26116,N_25553);
nand U26785 (N_26785,N_26004,N_25308);
nand U26786 (N_26786,N_25880,N_26392);
and U26787 (N_26787,N_25576,N_25442);
xor U26788 (N_26788,N_25819,N_25802);
and U26789 (N_26789,N_26257,N_26072);
xor U26790 (N_26790,N_25725,N_25832);
or U26791 (N_26791,N_25610,N_26020);
or U26792 (N_26792,N_26028,N_25624);
nand U26793 (N_26793,N_26109,N_26156);
nand U26794 (N_26794,N_25706,N_25590);
xor U26795 (N_26795,N_26349,N_25604);
nor U26796 (N_26796,N_26163,N_25418);
xor U26797 (N_26797,N_26328,N_26307);
nand U26798 (N_26798,N_26215,N_25927);
nand U26799 (N_26799,N_25662,N_26223);
or U26800 (N_26800,N_25398,N_25256);
and U26801 (N_26801,N_25200,N_26325);
nand U26802 (N_26802,N_25754,N_25717);
and U26803 (N_26803,N_25641,N_26332);
xor U26804 (N_26804,N_25331,N_26204);
or U26805 (N_26805,N_25757,N_25304);
nand U26806 (N_26806,N_25611,N_25768);
or U26807 (N_26807,N_25468,N_25814);
nor U26808 (N_26808,N_25380,N_25852);
nor U26809 (N_26809,N_25798,N_26015);
nand U26810 (N_26810,N_25487,N_25274);
or U26811 (N_26811,N_26218,N_25720);
xnor U26812 (N_26812,N_26132,N_25632);
and U26813 (N_26813,N_25967,N_25979);
or U26814 (N_26814,N_25741,N_26157);
xor U26815 (N_26815,N_25337,N_25656);
nor U26816 (N_26816,N_25947,N_25244);
nor U26817 (N_26817,N_25560,N_25250);
and U26818 (N_26818,N_25215,N_26135);
and U26819 (N_26819,N_26191,N_25729);
and U26820 (N_26820,N_26219,N_25884);
and U26821 (N_26821,N_25510,N_25740);
and U26822 (N_26822,N_25498,N_26141);
or U26823 (N_26823,N_25678,N_26397);
or U26824 (N_26824,N_25598,N_25914);
nor U26825 (N_26825,N_25896,N_25221);
xnor U26826 (N_26826,N_25517,N_26075);
and U26827 (N_26827,N_26014,N_26335);
or U26828 (N_26828,N_25796,N_25445);
nand U26829 (N_26829,N_25799,N_25283);
xnor U26830 (N_26830,N_26050,N_26089);
or U26831 (N_26831,N_25233,N_26134);
or U26832 (N_26832,N_26305,N_25474);
xnor U26833 (N_26833,N_25605,N_25500);
nor U26834 (N_26834,N_26263,N_25712);
or U26835 (N_26835,N_25833,N_26047);
nand U26836 (N_26836,N_25251,N_25419);
and U26837 (N_26837,N_25746,N_26286);
nand U26838 (N_26838,N_26350,N_25582);
nand U26839 (N_26839,N_26357,N_25424);
nor U26840 (N_26840,N_25587,N_25303);
or U26841 (N_26841,N_26297,N_25575);
nand U26842 (N_26842,N_25609,N_25829);
nand U26843 (N_26843,N_26105,N_25511);
or U26844 (N_26844,N_26289,N_25937);
nand U26845 (N_26845,N_26019,N_26346);
xnor U26846 (N_26846,N_26383,N_25570);
nor U26847 (N_26847,N_25831,N_26282);
xor U26848 (N_26848,N_26288,N_25206);
or U26849 (N_26849,N_25899,N_25911);
nor U26850 (N_26850,N_26103,N_26008);
and U26851 (N_26851,N_26091,N_25803);
xnor U26852 (N_26852,N_26243,N_25558);
nand U26853 (N_26853,N_25834,N_25737);
and U26854 (N_26854,N_25242,N_25447);
nor U26855 (N_26855,N_26025,N_25435);
nand U26856 (N_26856,N_26186,N_26107);
and U26857 (N_26857,N_25962,N_25929);
and U26858 (N_26858,N_25426,N_26092);
or U26859 (N_26859,N_25540,N_25310);
and U26860 (N_26860,N_25423,N_25437);
and U26861 (N_26861,N_25309,N_26209);
xnor U26862 (N_26862,N_26041,N_25623);
and U26863 (N_26863,N_25436,N_26194);
or U26864 (N_26864,N_25502,N_25722);
xnor U26865 (N_26865,N_26327,N_25775);
or U26866 (N_26866,N_25277,N_25933);
nor U26867 (N_26867,N_25460,N_26140);
nor U26868 (N_26868,N_25868,N_26313);
nor U26869 (N_26869,N_25282,N_25249);
or U26870 (N_26870,N_25995,N_25541);
nand U26871 (N_26871,N_25354,N_25262);
xnor U26872 (N_26872,N_25730,N_26238);
xnor U26873 (N_26873,N_25821,N_25871);
nor U26874 (N_26874,N_25809,N_26002);
nor U26875 (N_26875,N_26083,N_25918);
or U26876 (N_26876,N_25861,N_25782);
xor U26877 (N_26877,N_25522,N_26287);
nand U26878 (N_26878,N_26123,N_25446);
nor U26879 (N_26879,N_25328,N_26212);
nor U26880 (N_26880,N_25403,N_26087);
nand U26881 (N_26881,N_25311,N_25898);
and U26882 (N_26882,N_25411,N_25410);
xor U26883 (N_26883,N_25513,N_25691);
nand U26884 (N_26884,N_25506,N_25841);
nor U26885 (N_26885,N_25902,N_25578);
nand U26886 (N_26886,N_25790,N_25901);
xnor U26887 (N_26887,N_25408,N_26396);
or U26888 (N_26888,N_25837,N_25597);
or U26889 (N_26889,N_25991,N_26032);
and U26890 (N_26890,N_25577,N_25941);
or U26891 (N_26891,N_26386,N_25557);
nor U26892 (N_26892,N_25716,N_26374);
nand U26893 (N_26893,N_25355,N_25417);
xnor U26894 (N_26894,N_25228,N_25220);
or U26895 (N_26895,N_25361,N_25372);
nor U26896 (N_26896,N_25823,N_26035);
xor U26897 (N_26897,N_25551,N_26211);
or U26898 (N_26898,N_26224,N_25543);
or U26899 (N_26899,N_26347,N_25348);
xor U26900 (N_26900,N_25583,N_25489);
nand U26901 (N_26901,N_26102,N_26039);
xor U26902 (N_26902,N_26060,N_26210);
nor U26903 (N_26903,N_25275,N_25950);
xnor U26904 (N_26904,N_25942,N_25387);
or U26905 (N_26905,N_25207,N_26205);
and U26906 (N_26906,N_26368,N_25810);
or U26907 (N_26907,N_26237,N_25495);
xnor U26908 (N_26908,N_25978,N_26387);
and U26909 (N_26909,N_25535,N_25855);
or U26910 (N_26910,N_26126,N_25456);
and U26911 (N_26911,N_25409,N_25710);
or U26912 (N_26912,N_25528,N_25492);
or U26913 (N_26913,N_25992,N_26234);
or U26914 (N_26914,N_25908,N_25567);
nor U26915 (N_26915,N_25438,N_25269);
nor U26916 (N_26916,N_26232,N_25857);
nor U26917 (N_26917,N_26208,N_25648);
nand U26918 (N_26918,N_26139,N_25324);
nand U26919 (N_26919,N_25562,N_26380);
nand U26920 (N_26920,N_25989,N_25879);
and U26921 (N_26921,N_25886,N_26122);
nand U26922 (N_26922,N_26178,N_25428);
and U26923 (N_26923,N_25923,N_26213);
and U26924 (N_26924,N_25836,N_25780);
or U26925 (N_26925,N_25964,N_25681);
nand U26926 (N_26926,N_25286,N_25556);
or U26927 (N_26927,N_25847,N_25356);
and U26928 (N_26928,N_26172,N_25862);
xnor U26929 (N_26929,N_25434,N_25966);
xnor U26930 (N_26930,N_25520,N_25531);
nor U26931 (N_26931,N_26129,N_25888);
and U26932 (N_26932,N_26128,N_25616);
or U26933 (N_26933,N_25476,N_25915);
and U26934 (N_26934,N_25670,N_25320);
nor U26935 (N_26935,N_25647,N_26319);
and U26936 (N_26936,N_26308,N_25931);
nor U26937 (N_26937,N_25776,N_25939);
and U26938 (N_26938,N_26001,N_25284);
or U26939 (N_26939,N_25561,N_26294);
nand U26940 (N_26940,N_25726,N_25216);
nand U26941 (N_26941,N_26049,N_26364);
or U26942 (N_26942,N_25874,N_25684);
nor U26943 (N_26943,N_25305,N_25986);
or U26944 (N_26944,N_25910,N_25366);
xor U26945 (N_26945,N_25665,N_25368);
nor U26946 (N_26946,N_26296,N_25376);
or U26947 (N_26947,N_26336,N_25976);
nor U26948 (N_26948,N_25892,N_26022);
nor U26949 (N_26949,N_25257,N_25464);
nand U26950 (N_26950,N_25773,N_26261);
or U26951 (N_26951,N_26166,N_25406);
and U26952 (N_26952,N_26064,N_26161);
nor U26953 (N_26953,N_25461,N_26398);
nor U26954 (N_26954,N_25633,N_25794);
and U26955 (N_26955,N_26059,N_26203);
nor U26956 (N_26956,N_25781,N_25238);
nor U26957 (N_26957,N_26148,N_25696);
or U26958 (N_26958,N_25672,N_25878);
nor U26959 (N_26959,N_26130,N_26222);
and U26960 (N_26960,N_25805,N_26240);
xnor U26961 (N_26961,N_25323,N_26221);
nand U26962 (N_26962,N_25344,N_25718);
xnor U26963 (N_26963,N_25393,N_25480);
xnor U26964 (N_26964,N_26362,N_25501);
nand U26965 (N_26965,N_25260,N_25734);
nor U26966 (N_26966,N_25596,N_25326);
nand U26967 (N_26967,N_25507,N_25638);
or U26968 (N_26968,N_25867,N_25518);
nor U26969 (N_26969,N_25835,N_26310);
or U26970 (N_26970,N_25639,N_26114);
nand U26971 (N_26971,N_25687,N_25536);
nand U26972 (N_26972,N_25585,N_26012);
or U26973 (N_26973,N_25702,N_25679);
xor U26974 (N_26974,N_25210,N_25807);
nor U26975 (N_26975,N_26106,N_26266);
xor U26976 (N_26976,N_26110,N_26030);
and U26977 (N_26977,N_25677,N_26192);
nand U26978 (N_26978,N_25748,N_25263);
xnor U26979 (N_26979,N_25245,N_25586);
nor U26980 (N_26980,N_26009,N_26216);
xnor U26981 (N_26981,N_25872,N_26324);
xor U26982 (N_26982,N_26045,N_26006);
nand U26983 (N_26983,N_26358,N_26021);
xnor U26984 (N_26984,N_25928,N_26333);
nand U26985 (N_26985,N_26225,N_25848);
nor U26986 (N_26986,N_26052,N_25728);
nand U26987 (N_26987,N_25971,N_26298);
nor U26988 (N_26988,N_25980,N_25804);
nor U26989 (N_26989,N_26196,N_25381);
or U26990 (N_26990,N_25682,N_25533);
nand U26991 (N_26991,N_25534,N_25882);
nand U26992 (N_26992,N_26146,N_26076);
and U26993 (N_26993,N_26262,N_26326);
nand U26994 (N_26994,N_26318,N_25642);
nor U26995 (N_26995,N_25719,N_25998);
nor U26996 (N_26996,N_26378,N_26095);
and U26997 (N_26997,N_25970,N_25285);
or U26998 (N_26998,N_25521,N_25844);
nor U26999 (N_26999,N_25612,N_26253);
nor U27000 (N_27000,N_26028,N_25234);
xnor U27001 (N_27001,N_26399,N_25972);
nand U27002 (N_27002,N_25462,N_25303);
nand U27003 (N_27003,N_25604,N_25496);
xnor U27004 (N_27004,N_25970,N_25244);
or U27005 (N_27005,N_25429,N_25548);
nand U27006 (N_27006,N_26364,N_25837);
nor U27007 (N_27007,N_25932,N_26377);
nor U27008 (N_27008,N_25415,N_26156);
xor U27009 (N_27009,N_26292,N_25628);
nand U27010 (N_27010,N_25278,N_25285);
nand U27011 (N_27011,N_25364,N_25623);
nor U27012 (N_27012,N_26082,N_25886);
nand U27013 (N_27013,N_26009,N_26283);
or U27014 (N_27014,N_25981,N_26096);
xnor U27015 (N_27015,N_26300,N_25830);
nor U27016 (N_27016,N_25521,N_25455);
xnor U27017 (N_27017,N_25702,N_25621);
and U27018 (N_27018,N_25592,N_25514);
or U27019 (N_27019,N_25649,N_25968);
nor U27020 (N_27020,N_26274,N_25264);
nor U27021 (N_27021,N_25980,N_25751);
nand U27022 (N_27022,N_25772,N_26111);
nand U27023 (N_27023,N_26300,N_26139);
and U27024 (N_27024,N_26005,N_25701);
xor U27025 (N_27025,N_26197,N_25264);
and U27026 (N_27026,N_25256,N_25713);
nor U27027 (N_27027,N_25974,N_26216);
nand U27028 (N_27028,N_25488,N_25437);
and U27029 (N_27029,N_25362,N_25494);
nor U27030 (N_27030,N_25256,N_25253);
xnor U27031 (N_27031,N_25472,N_25868);
and U27032 (N_27032,N_25577,N_26198);
or U27033 (N_27033,N_26102,N_26046);
or U27034 (N_27034,N_25389,N_25400);
nor U27035 (N_27035,N_26216,N_25347);
nand U27036 (N_27036,N_26346,N_25668);
xor U27037 (N_27037,N_26032,N_26290);
xor U27038 (N_27038,N_26062,N_25697);
xnor U27039 (N_27039,N_25241,N_25605);
nand U27040 (N_27040,N_25715,N_26146);
nand U27041 (N_27041,N_26011,N_25585);
and U27042 (N_27042,N_25810,N_25715);
and U27043 (N_27043,N_26244,N_25765);
or U27044 (N_27044,N_25268,N_26172);
nand U27045 (N_27045,N_25783,N_25818);
and U27046 (N_27046,N_26000,N_25659);
xnor U27047 (N_27047,N_26138,N_26024);
nand U27048 (N_27048,N_25965,N_26338);
and U27049 (N_27049,N_25213,N_25696);
and U27050 (N_27050,N_25600,N_25224);
and U27051 (N_27051,N_26114,N_25533);
nand U27052 (N_27052,N_25897,N_26139);
and U27053 (N_27053,N_25460,N_25501);
xnor U27054 (N_27054,N_25320,N_25875);
nor U27055 (N_27055,N_26334,N_25393);
xor U27056 (N_27056,N_25620,N_25997);
xnor U27057 (N_27057,N_26321,N_26282);
or U27058 (N_27058,N_26387,N_25943);
and U27059 (N_27059,N_25543,N_26111);
and U27060 (N_27060,N_25255,N_25542);
and U27061 (N_27061,N_26373,N_25634);
and U27062 (N_27062,N_26126,N_26274);
and U27063 (N_27063,N_25396,N_26146);
nand U27064 (N_27064,N_26300,N_25263);
nor U27065 (N_27065,N_25597,N_25257);
xor U27066 (N_27066,N_25354,N_25703);
or U27067 (N_27067,N_25977,N_25944);
nand U27068 (N_27068,N_25737,N_26159);
xnor U27069 (N_27069,N_25337,N_25865);
or U27070 (N_27070,N_26378,N_25354);
nand U27071 (N_27071,N_25921,N_25262);
nor U27072 (N_27072,N_26242,N_26155);
nand U27073 (N_27073,N_25753,N_25822);
and U27074 (N_27074,N_25522,N_26177);
nand U27075 (N_27075,N_26080,N_25876);
nand U27076 (N_27076,N_25346,N_25354);
nor U27077 (N_27077,N_25993,N_25237);
xnor U27078 (N_27078,N_26296,N_26123);
nand U27079 (N_27079,N_25637,N_25508);
nor U27080 (N_27080,N_25694,N_26065);
or U27081 (N_27081,N_25286,N_26029);
and U27082 (N_27082,N_25718,N_25594);
or U27083 (N_27083,N_25357,N_26032);
or U27084 (N_27084,N_26392,N_25465);
nor U27085 (N_27085,N_25442,N_26163);
xnor U27086 (N_27086,N_26177,N_25571);
nor U27087 (N_27087,N_25410,N_26045);
nand U27088 (N_27088,N_25892,N_25612);
and U27089 (N_27089,N_25574,N_26381);
and U27090 (N_27090,N_26270,N_26269);
xor U27091 (N_27091,N_25546,N_25962);
xor U27092 (N_27092,N_25955,N_26134);
nand U27093 (N_27093,N_26288,N_26124);
nand U27094 (N_27094,N_25429,N_26125);
and U27095 (N_27095,N_25222,N_25965);
xor U27096 (N_27096,N_25429,N_26397);
nand U27097 (N_27097,N_26113,N_25297);
xnor U27098 (N_27098,N_26256,N_26393);
nor U27099 (N_27099,N_25840,N_25847);
xor U27100 (N_27100,N_25598,N_25369);
and U27101 (N_27101,N_25698,N_25427);
and U27102 (N_27102,N_25906,N_25354);
nand U27103 (N_27103,N_25208,N_25853);
nor U27104 (N_27104,N_25694,N_25726);
nor U27105 (N_27105,N_25660,N_25250);
xor U27106 (N_27106,N_25637,N_25334);
or U27107 (N_27107,N_25594,N_26357);
nand U27108 (N_27108,N_26292,N_26102);
nand U27109 (N_27109,N_26160,N_25327);
nand U27110 (N_27110,N_25572,N_25215);
nand U27111 (N_27111,N_26266,N_25469);
and U27112 (N_27112,N_25933,N_26113);
xnor U27113 (N_27113,N_25742,N_25227);
nand U27114 (N_27114,N_26397,N_26138);
and U27115 (N_27115,N_26279,N_26289);
and U27116 (N_27116,N_26270,N_26028);
xor U27117 (N_27117,N_25456,N_25849);
xor U27118 (N_27118,N_25640,N_26051);
nand U27119 (N_27119,N_25874,N_25791);
nor U27120 (N_27120,N_26006,N_26284);
nand U27121 (N_27121,N_26042,N_26138);
xnor U27122 (N_27122,N_26131,N_25600);
or U27123 (N_27123,N_26112,N_25436);
or U27124 (N_27124,N_25341,N_26339);
xnor U27125 (N_27125,N_25946,N_25364);
nand U27126 (N_27126,N_25306,N_25957);
or U27127 (N_27127,N_25955,N_25416);
and U27128 (N_27128,N_25709,N_25789);
xor U27129 (N_27129,N_26108,N_25294);
xor U27130 (N_27130,N_25547,N_25757);
xor U27131 (N_27131,N_25642,N_25768);
and U27132 (N_27132,N_25951,N_25770);
or U27133 (N_27133,N_26098,N_25424);
or U27134 (N_27134,N_25576,N_25910);
nor U27135 (N_27135,N_25866,N_25978);
nor U27136 (N_27136,N_25766,N_25791);
nand U27137 (N_27137,N_25505,N_25949);
and U27138 (N_27138,N_25615,N_26005);
nor U27139 (N_27139,N_26224,N_26342);
or U27140 (N_27140,N_26391,N_25295);
or U27141 (N_27141,N_25700,N_26164);
xnor U27142 (N_27142,N_26239,N_25575);
xor U27143 (N_27143,N_25712,N_25658);
and U27144 (N_27144,N_25315,N_25760);
nor U27145 (N_27145,N_25655,N_26144);
nand U27146 (N_27146,N_25951,N_26381);
xor U27147 (N_27147,N_26224,N_25243);
or U27148 (N_27148,N_25222,N_25605);
or U27149 (N_27149,N_25675,N_25495);
or U27150 (N_27150,N_26220,N_25987);
nand U27151 (N_27151,N_26332,N_25737);
nor U27152 (N_27152,N_26190,N_26327);
xor U27153 (N_27153,N_25487,N_25328);
nor U27154 (N_27154,N_26072,N_26312);
nand U27155 (N_27155,N_26151,N_25572);
nor U27156 (N_27156,N_25639,N_25605);
nand U27157 (N_27157,N_25580,N_25955);
xor U27158 (N_27158,N_25912,N_26340);
xor U27159 (N_27159,N_25667,N_25509);
nand U27160 (N_27160,N_25633,N_26147);
xnor U27161 (N_27161,N_25878,N_25888);
nand U27162 (N_27162,N_25880,N_26259);
nor U27163 (N_27163,N_25624,N_26254);
nand U27164 (N_27164,N_25999,N_25538);
and U27165 (N_27165,N_25614,N_25661);
or U27166 (N_27166,N_25377,N_26304);
and U27167 (N_27167,N_25989,N_26016);
xor U27168 (N_27168,N_26315,N_26067);
nor U27169 (N_27169,N_26313,N_25610);
or U27170 (N_27170,N_26361,N_26208);
nor U27171 (N_27171,N_25557,N_26058);
xnor U27172 (N_27172,N_26183,N_26111);
nand U27173 (N_27173,N_26175,N_25499);
nand U27174 (N_27174,N_25976,N_25237);
nor U27175 (N_27175,N_25482,N_25901);
xor U27176 (N_27176,N_25820,N_25265);
nor U27177 (N_27177,N_25271,N_26258);
and U27178 (N_27178,N_25646,N_26176);
and U27179 (N_27179,N_26098,N_26232);
and U27180 (N_27180,N_25566,N_25724);
and U27181 (N_27181,N_26137,N_25487);
nor U27182 (N_27182,N_25400,N_26077);
and U27183 (N_27183,N_25274,N_25450);
nor U27184 (N_27184,N_25647,N_25238);
nor U27185 (N_27185,N_25349,N_26072);
nor U27186 (N_27186,N_26156,N_26119);
xnor U27187 (N_27187,N_26301,N_25973);
or U27188 (N_27188,N_25237,N_25978);
xor U27189 (N_27189,N_25736,N_25276);
and U27190 (N_27190,N_25545,N_25516);
or U27191 (N_27191,N_25504,N_26314);
and U27192 (N_27192,N_25415,N_25813);
xnor U27193 (N_27193,N_25978,N_26086);
or U27194 (N_27194,N_25485,N_25593);
or U27195 (N_27195,N_25418,N_25804);
and U27196 (N_27196,N_25437,N_25314);
nor U27197 (N_27197,N_26000,N_26154);
nand U27198 (N_27198,N_26375,N_25678);
nand U27199 (N_27199,N_25346,N_26303);
nand U27200 (N_27200,N_25313,N_25783);
and U27201 (N_27201,N_25287,N_25725);
nand U27202 (N_27202,N_25427,N_25766);
or U27203 (N_27203,N_25715,N_26361);
xnor U27204 (N_27204,N_25779,N_25277);
or U27205 (N_27205,N_25626,N_26327);
nor U27206 (N_27206,N_25830,N_25261);
or U27207 (N_27207,N_25675,N_26068);
or U27208 (N_27208,N_25970,N_25363);
nor U27209 (N_27209,N_25641,N_25352);
xor U27210 (N_27210,N_25829,N_25326);
nor U27211 (N_27211,N_25485,N_26374);
xor U27212 (N_27212,N_25387,N_26311);
or U27213 (N_27213,N_26331,N_25866);
xnor U27214 (N_27214,N_25731,N_25261);
and U27215 (N_27215,N_25460,N_25309);
nand U27216 (N_27216,N_25935,N_25537);
nor U27217 (N_27217,N_26260,N_26094);
nor U27218 (N_27218,N_25271,N_26391);
nand U27219 (N_27219,N_26296,N_25934);
nand U27220 (N_27220,N_25709,N_26395);
nand U27221 (N_27221,N_26122,N_25862);
and U27222 (N_27222,N_26354,N_26318);
and U27223 (N_27223,N_26090,N_26038);
or U27224 (N_27224,N_25834,N_25433);
and U27225 (N_27225,N_25929,N_25925);
and U27226 (N_27226,N_25648,N_26230);
and U27227 (N_27227,N_26009,N_25507);
xnor U27228 (N_27228,N_26179,N_25376);
xor U27229 (N_27229,N_25828,N_25717);
xnor U27230 (N_27230,N_26129,N_26130);
and U27231 (N_27231,N_25619,N_25492);
xor U27232 (N_27232,N_25638,N_25269);
xnor U27233 (N_27233,N_25722,N_26132);
nor U27234 (N_27234,N_25853,N_25806);
or U27235 (N_27235,N_26098,N_26257);
and U27236 (N_27236,N_25521,N_25504);
xnor U27237 (N_27237,N_25304,N_25262);
or U27238 (N_27238,N_25645,N_26127);
or U27239 (N_27239,N_26284,N_25221);
or U27240 (N_27240,N_25226,N_25781);
or U27241 (N_27241,N_25560,N_26134);
or U27242 (N_27242,N_25371,N_25260);
or U27243 (N_27243,N_25716,N_25938);
nand U27244 (N_27244,N_26242,N_25345);
or U27245 (N_27245,N_25383,N_25624);
and U27246 (N_27246,N_25570,N_26201);
and U27247 (N_27247,N_25874,N_25753);
nor U27248 (N_27248,N_25581,N_26291);
xor U27249 (N_27249,N_26378,N_26116);
xor U27250 (N_27250,N_25743,N_25887);
nor U27251 (N_27251,N_26256,N_25293);
nor U27252 (N_27252,N_26115,N_26169);
or U27253 (N_27253,N_25428,N_25706);
nand U27254 (N_27254,N_25507,N_25973);
nand U27255 (N_27255,N_25592,N_26078);
or U27256 (N_27256,N_25679,N_25386);
and U27257 (N_27257,N_25453,N_25448);
nand U27258 (N_27258,N_25989,N_26351);
nand U27259 (N_27259,N_25319,N_26076);
and U27260 (N_27260,N_26338,N_25711);
and U27261 (N_27261,N_25785,N_25692);
nand U27262 (N_27262,N_25715,N_25419);
and U27263 (N_27263,N_25698,N_25474);
or U27264 (N_27264,N_25449,N_25282);
or U27265 (N_27265,N_25240,N_26385);
and U27266 (N_27266,N_25980,N_25387);
or U27267 (N_27267,N_25832,N_26069);
or U27268 (N_27268,N_26146,N_25806);
nand U27269 (N_27269,N_25883,N_25649);
xnor U27270 (N_27270,N_26145,N_26381);
or U27271 (N_27271,N_25578,N_25204);
or U27272 (N_27272,N_26061,N_26137);
or U27273 (N_27273,N_26046,N_25959);
nor U27274 (N_27274,N_25541,N_26193);
or U27275 (N_27275,N_25296,N_25995);
nand U27276 (N_27276,N_26117,N_25585);
and U27277 (N_27277,N_26243,N_26150);
or U27278 (N_27278,N_25393,N_26210);
and U27279 (N_27279,N_25769,N_25476);
or U27280 (N_27280,N_26203,N_25442);
nand U27281 (N_27281,N_25246,N_26162);
or U27282 (N_27282,N_25802,N_25783);
nand U27283 (N_27283,N_25932,N_25953);
nor U27284 (N_27284,N_25954,N_25903);
or U27285 (N_27285,N_25639,N_25856);
or U27286 (N_27286,N_25490,N_25780);
nand U27287 (N_27287,N_26074,N_26382);
or U27288 (N_27288,N_25474,N_26121);
nand U27289 (N_27289,N_26361,N_26398);
and U27290 (N_27290,N_25962,N_26059);
and U27291 (N_27291,N_26269,N_26094);
nand U27292 (N_27292,N_25810,N_25615);
xor U27293 (N_27293,N_25519,N_25730);
xnor U27294 (N_27294,N_26201,N_26262);
nor U27295 (N_27295,N_25861,N_26087);
nand U27296 (N_27296,N_26217,N_25456);
nor U27297 (N_27297,N_25364,N_26301);
and U27298 (N_27298,N_26240,N_25639);
or U27299 (N_27299,N_25946,N_25273);
or U27300 (N_27300,N_26044,N_25236);
xnor U27301 (N_27301,N_25449,N_25387);
or U27302 (N_27302,N_25665,N_26160);
xor U27303 (N_27303,N_25896,N_26273);
nor U27304 (N_27304,N_25845,N_25933);
or U27305 (N_27305,N_26338,N_25700);
and U27306 (N_27306,N_26033,N_25555);
or U27307 (N_27307,N_25973,N_26288);
xnor U27308 (N_27308,N_25509,N_25504);
or U27309 (N_27309,N_26291,N_25322);
xor U27310 (N_27310,N_25749,N_25831);
nand U27311 (N_27311,N_25945,N_25849);
xnor U27312 (N_27312,N_26047,N_25514);
xor U27313 (N_27313,N_26224,N_26177);
nor U27314 (N_27314,N_26193,N_25344);
and U27315 (N_27315,N_26371,N_25713);
nand U27316 (N_27316,N_25714,N_25520);
nand U27317 (N_27317,N_26338,N_26204);
and U27318 (N_27318,N_25642,N_25965);
or U27319 (N_27319,N_25258,N_25980);
nor U27320 (N_27320,N_25830,N_25288);
and U27321 (N_27321,N_26313,N_25793);
nor U27322 (N_27322,N_26380,N_25306);
and U27323 (N_27323,N_25718,N_25813);
and U27324 (N_27324,N_25487,N_26184);
and U27325 (N_27325,N_26105,N_25832);
nand U27326 (N_27326,N_25523,N_25572);
nor U27327 (N_27327,N_26387,N_26290);
and U27328 (N_27328,N_26208,N_25544);
and U27329 (N_27329,N_26126,N_25206);
xnor U27330 (N_27330,N_26379,N_25357);
xor U27331 (N_27331,N_25499,N_26274);
and U27332 (N_27332,N_25714,N_26024);
or U27333 (N_27333,N_25870,N_25353);
or U27334 (N_27334,N_26249,N_25732);
xor U27335 (N_27335,N_25667,N_26182);
nor U27336 (N_27336,N_25329,N_25706);
and U27337 (N_27337,N_26104,N_26243);
nor U27338 (N_27338,N_25306,N_26170);
nand U27339 (N_27339,N_25516,N_25377);
or U27340 (N_27340,N_25305,N_25363);
or U27341 (N_27341,N_25867,N_26032);
nor U27342 (N_27342,N_25226,N_26020);
xnor U27343 (N_27343,N_25485,N_26071);
nand U27344 (N_27344,N_26295,N_25668);
xor U27345 (N_27345,N_26022,N_25327);
nor U27346 (N_27346,N_25577,N_26077);
xnor U27347 (N_27347,N_26384,N_25827);
nand U27348 (N_27348,N_26051,N_25851);
or U27349 (N_27349,N_25326,N_25953);
nand U27350 (N_27350,N_25650,N_25483);
or U27351 (N_27351,N_26250,N_26189);
nand U27352 (N_27352,N_26189,N_25936);
or U27353 (N_27353,N_25302,N_25465);
or U27354 (N_27354,N_26374,N_25231);
nor U27355 (N_27355,N_25977,N_25348);
and U27356 (N_27356,N_25681,N_25954);
xor U27357 (N_27357,N_25830,N_26286);
and U27358 (N_27358,N_25375,N_25766);
nand U27359 (N_27359,N_26045,N_26137);
and U27360 (N_27360,N_26211,N_26311);
nand U27361 (N_27361,N_25784,N_26103);
or U27362 (N_27362,N_25901,N_25981);
nand U27363 (N_27363,N_26100,N_26081);
nor U27364 (N_27364,N_25422,N_26302);
and U27365 (N_27365,N_25407,N_25351);
or U27366 (N_27366,N_26025,N_25353);
and U27367 (N_27367,N_26362,N_25441);
or U27368 (N_27368,N_26188,N_25533);
nor U27369 (N_27369,N_25432,N_25834);
nor U27370 (N_27370,N_25620,N_26398);
or U27371 (N_27371,N_26220,N_25453);
xor U27372 (N_27372,N_26222,N_25479);
xor U27373 (N_27373,N_26263,N_26010);
or U27374 (N_27374,N_25927,N_25910);
nor U27375 (N_27375,N_25283,N_25587);
xor U27376 (N_27376,N_26052,N_25817);
xor U27377 (N_27377,N_25913,N_26157);
nand U27378 (N_27378,N_25415,N_25753);
nor U27379 (N_27379,N_26101,N_26253);
nand U27380 (N_27380,N_26050,N_25785);
and U27381 (N_27381,N_25348,N_26364);
nand U27382 (N_27382,N_25764,N_25558);
xor U27383 (N_27383,N_25677,N_25663);
and U27384 (N_27384,N_25365,N_26332);
nor U27385 (N_27385,N_26256,N_25856);
and U27386 (N_27386,N_25992,N_25734);
xnor U27387 (N_27387,N_25403,N_25376);
and U27388 (N_27388,N_25610,N_25403);
and U27389 (N_27389,N_26167,N_25391);
and U27390 (N_27390,N_26320,N_26208);
and U27391 (N_27391,N_26200,N_25522);
or U27392 (N_27392,N_25698,N_25949);
xnor U27393 (N_27393,N_25362,N_25643);
nor U27394 (N_27394,N_26018,N_25483);
nor U27395 (N_27395,N_26027,N_25840);
nor U27396 (N_27396,N_25381,N_25735);
nor U27397 (N_27397,N_25803,N_25299);
nor U27398 (N_27398,N_25897,N_25508);
nor U27399 (N_27399,N_25219,N_26266);
nor U27400 (N_27400,N_25526,N_25733);
nor U27401 (N_27401,N_26066,N_25356);
xor U27402 (N_27402,N_26002,N_25825);
or U27403 (N_27403,N_25779,N_25398);
and U27404 (N_27404,N_25572,N_25810);
or U27405 (N_27405,N_25520,N_26216);
xor U27406 (N_27406,N_25551,N_26127);
nand U27407 (N_27407,N_25345,N_25703);
or U27408 (N_27408,N_25972,N_25696);
and U27409 (N_27409,N_26006,N_25691);
and U27410 (N_27410,N_25413,N_26105);
xor U27411 (N_27411,N_25699,N_25821);
nand U27412 (N_27412,N_25729,N_25267);
or U27413 (N_27413,N_26054,N_25246);
and U27414 (N_27414,N_26167,N_25308);
nand U27415 (N_27415,N_25614,N_25828);
or U27416 (N_27416,N_26042,N_25522);
or U27417 (N_27417,N_25575,N_26238);
and U27418 (N_27418,N_25949,N_26206);
nor U27419 (N_27419,N_25462,N_25844);
and U27420 (N_27420,N_25309,N_25638);
or U27421 (N_27421,N_26347,N_25311);
xnor U27422 (N_27422,N_26377,N_25919);
nand U27423 (N_27423,N_26269,N_26203);
xnor U27424 (N_27424,N_26078,N_25205);
xnor U27425 (N_27425,N_25271,N_26020);
and U27426 (N_27426,N_25711,N_25276);
xor U27427 (N_27427,N_25637,N_25322);
or U27428 (N_27428,N_26148,N_26153);
and U27429 (N_27429,N_25855,N_25286);
nor U27430 (N_27430,N_25256,N_26260);
or U27431 (N_27431,N_25362,N_26217);
nor U27432 (N_27432,N_26064,N_26343);
nand U27433 (N_27433,N_25764,N_25444);
or U27434 (N_27434,N_25445,N_25408);
xnor U27435 (N_27435,N_26257,N_25482);
and U27436 (N_27436,N_25627,N_26308);
nor U27437 (N_27437,N_26368,N_25448);
nand U27438 (N_27438,N_25496,N_26393);
or U27439 (N_27439,N_25650,N_26167);
xor U27440 (N_27440,N_25517,N_26319);
nand U27441 (N_27441,N_25277,N_26271);
or U27442 (N_27442,N_26305,N_25709);
nand U27443 (N_27443,N_26209,N_25840);
nor U27444 (N_27444,N_26321,N_26357);
nor U27445 (N_27445,N_25380,N_26180);
or U27446 (N_27446,N_26248,N_25911);
nand U27447 (N_27447,N_25782,N_25911);
xnor U27448 (N_27448,N_25636,N_25994);
and U27449 (N_27449,N_25869,N_25332);
xor U27450 (N_27450,N_25334,N_25933);
nor U27451 (N_27451,N_26319,N_25865);
and U27452 (N_27452,N_26033,N_25688);
nand U27453 (N_27453,N_26116,N_26369);
and U27454 (N_27454,N_26152,N_25519);
or U27455 (N_27455,N_25953,N_25727);
and U27456 (N_27456,N_25550,N_25225);
and U27457 (N_27457,N_26134,N_25232);
xor U27458 (N_27458,N_25716,N_25584);
nand U27459 (N_27459,N_26052,N_25350);
and U27460 (N_27460,N_25741,N_26224);
or U27461 (N_27461,N_25285,N_25941);
nor U27462 (N_27462,N_26065,N_26180);
nand U27463 (N_27463,N_25688,N_25637);
and U27464 (N_27464,N_25297,N_26390);
and U27465 (N_27465,N_25706,N_26047);
and U27466 (N_27466,N_25610,N_25318);
and U27467 (N_27467,N_26112,N_25573);
or U27468 (N_27468,N_25258,N_26178);
or U27469 (N_27469,N_25866,N_25276);
xor U27470 (N_27470,N_25920,N_26063);
and U27471 (N_27471,N_25284,N_25829);
or U27472 (N_27472,N_25773,N_25819);
xnor U27473 (N_27473,N_26297,N_26279);
and U27474 (N_27474,N_25207,N_26174);
or U27475 (N_27475,N_26206,N_25610);
and U27476 (N_27476,N_25986,N_25357);
nand U27477 (N_27477,N_25538,N_25669);
nand U27478 (N_27478,N_25912,N_26126);
or U27479 (N_27479,N_25877,N_26247);
nor U27480 (N_27480,N_25238,N_25250);
and U27481 (N_27481,N_26144,N_25439);
nand U27482 (N_27482,N_26365,N_25441);
and U27483 (N_27483,N_25253,N_25649);
and U27484 (N_27484,N_26100,N_25922);
xnor U27485 (N_27485,N_25573,N_26290);
and U27486 (N_27486,N_25326,N_25473);
and U27487 (N_27487,N_26224,N_25828);
xnor U27488 (N_27488,N_25917,N_26065);
nand U27489 (N_27489,N_25559,N_26265);
and U27490 (N_27490,N_26182,N_25991);
xor U27491 (N_27491,N_25904,N_25853);
and U27492 (N_27492,N_25590,N_25968);
xnor U27493 (N_27493,N_25602,N_25404);
or U27494 (N_27494,N_26219,N_25856);
or U27495 (N_27495,N_25445,N_26024);
and U27496 (N_27496,N_25790,N_25571);
and U27497 (N_27497,N_25453,N_25626);
xnor U27498 (N_27498,N_25524,N_26244);
nor U27499 (N_27499,N_25978,N_25705);
xor U27500 (N_27500,N_25948,N_25756);
nand U27501 (N_27501,N_26269,N_25971);
xor U27502 (N_27502,N_26220,N_26197);
or U27503 (N_27503,N_25709,N_25924);
or U27504 (N_27504,N_25304,N_25426);
nand U27505 (N_27505,N_25679,N_25957);
xnor U27506 (N_27506,N_25535,N_26307);
or U27507 (N_27507,N_25368,N_26358);
and U27508 (N_27508,N_25468,N_25351);
xnor U27509 (N_27509,N_25824,N_25625);
nand U27510 (N_27510,N_25586,N_25585);
nor U27511 (N_27511,N_25407,N_26017);
nor U27512 (N_27512,N_25725,N_25646);
or U27513 (N_27513,N_25527,N_26217);
nor U27514 (N_27514,N_25505,N_26118);
nor U27515 (N_27515,N_26121,N_25981);
or U27516 (N_27516,N_25849,N_25519);
nor U27517 (N_27517,N_25213,N_25306);
nor U27518 (N_27518,N_25214,N_26140);
and U27519 (N_27519,N_25422,N_25535);
nand U27520 (N_27520,N_26337,N_25669);
or U27521 (N_27521,N_25630,N_26098);
nor U27522 (N_27522,N_26199,N_25696);
or U27523 (N_27523,N_25772,N_25642);
nand U27524 (N_27524,N_25487,N_26290);
xnor U27525 (N_27525,N_25961,N_25643);
nor U27526 (N_27526,N_26371,N_25859);
or U27527 (N_27527,N_25463,N_25555);
and U27528 (N_27528,N_25548,N_26192);
and U27529 (N_27529,N_26114,N_26041);
or U27530 (N_27530,N_25781,N_26294);
nor U27531 (N_27531,N_25497,N_26136);
and U27532 (N_27532,N_25909,N_26008);
and U27533 (N_27533,N_25659,N_26115);
nand U27534 (N_27534,N_26034,N_25302);
and U27535 (N_27535,N_25729,N_25633);
and U27536 (N_27536,N_26295,N_25625);
nand U27537 (N_27537,N_26108,N_25709);
or U27538 (N_27538,N_25850,N_26024);
or U27539 (N_27539,N_25623,N_26179);
nor U27540 (N_27540,N_26395,N_26036);
and U27541 (N_27541,N_25776,N_25854);
xor U27542 (N_27542,N_25888,N_25681);
or U27543 (N_27543,N_26190,N_25918);
nand U27544 (N_27544,N_26300,N_25837);
xnor U27545 (N_27545,N_26338,N_25972);
nand U27546 (N_27546,N_25541,N_25969);
xor U27547 (N_27547,N_25851,N_25582);
and U27548 (N_27548,N_25907,N_26270);
or U27549 (N_27549,N_25417,N_25834);
nand U27550 (N_27550,N_26229,N_26350);
and U27551 (N_27551,N_26159,N_25899);
nor U27552 (N_27552,N_26207,N_25986);
or U27553 (N_27553,N_25830,N_25892);
xor U27554 (N_27554,N_26002,N_26349);
and U27555 (N_27555,N_25877,N_25746);
and U27556 (N_27556,N_25733,N_25233);
xnor U27557 (N_27557,N_25375,N_25287);
nor U27558 (N_27558,N_25663,N_25826);
and U27559 (N_27559,N_25939,N_26066);
and U27560 (N_27560,N_26162,N_26077);
xor U27561 (N_27561,N_26147,N_25913);
or U27562 (N_27562,N_25898,N_26211);
xor U27563 (N_27563,N_25772,N_26356);
nor U27564 (N_27564,N_25896,N_25314);
nand U27565 (N_27565,N_26359,N_25951);
or U27566 (N_27566,N_26181,N_25310);
nor U27567 (N_27567,N_25872,N_25817);
nand U27568 (N_27568,N_25246,N_25602);
nor U27569 (N_27569,N_25557,N_26327);
xnor U27570 (N_27570,N_25869,N_26353);
nand U27571 (N_27571,N_26061,N_25291);
nand U27572 (N_27572,N_25997,N_26113);
xnor U27573 (N_27573,N_26059,N_26053);
nand U27574 (N_27574,N_25839,N_25375);
and U27575 (N_27575,N_26306,N_25654);
or U27576 (N_27576,N_26149,N_25541);
nor U27577 (N_27577,N_25387,N_25564);
nor U27578 (N_27578,N_26299,N_25478);
or U27579 (N_27579,N_25961,N_25622);
nor U27580 (N_27580,N_26303,N_26096);
xor U27581 (N_27581,N_25496,N_25509);
xnor U27582 (N_27582,N_26344,N_25499);
or U27583 (N_27583,N_25636,N_25961);
or U27584 (N_27584,N_25555,N_25549);
nor U27585 (N_27585,N_26297,N_25930);
or U27586 (N_27586,N_25581,N_26327);
nor U27587 (N_27587,N_26059,N_25890);
or U27588 (N_27588,N_25736,N_26048);
and U27589 (N_27589,N_26374,N_25915);
and U27590 (N_27590,N_26247,N_26131);
nand U27591 (N_27591,N_25411,N_25449);
nand U27592 (N_27592,N_26037,N_25494);
xnor U27593 (N_27593,N_26294,N_25681);
xor U27594 (N_27594,N_25634,N_25934);
nor U27595 (N_27595,N_25500,N_26047);
and U27596 (N_27596,N_25358,N_25432);
nand U27597 (N_27597,N_25292,N_26250);
nor U27598 (N_27598,N_26057,N_25638);
nor U27599 (N_27599,N_26062,N_25340);
or U27600 (N_27600,N_26914,N_26850);
and U27601 (N_27601,N_26488,N_26954);
and U27602 (N_27602,N_27196,N_26896);
or U27603 (N_27603,N_26877,N_27498);
and U27604 (N_27604,N_27578,N_27456);
and U27605 (N_27605,N_26433,N_27470);
and U27606 (N_27606,N_27043,N_27049);
nand U27607 (N_27607,N_26884,N_27518);
nor U27608 (N_27608,N_27544,N_27213);
and U27609 (N_27609,N_26525,N_26645);
nand U27610 (N_27610,N_27262,N_27449);
and U27611 (N_27611,N_26978,N_27463);
xor U27612 (N_27612,N_27530,N_26431);
and U27613 (N_27613,N_27345,N_27417);
xnor U27614 (N_27614,N_27355,N_26744);
and U27615 (N_27615,N_26427,N_26554);
or U27616 (N_27616,N_27537,N_26933);
nand U27617 (N_27617,N_26802,N_27562);
xor U27618 (N_27618,N_27339,N_26632);
or U27619 (N_27619,N_27346,N_26757);
nor U27620 (N_27620,N_27200,N_26581);
nand U27621 (N_27621,N_27198,N_26718);
or U27622 (N_27622,N_26813,N_27121);
nor U27623 (N_27623,N_27547,N_27073);
or U27624 (N_27624,N_26668,N_27241);
and U27625 (N_27625,N_27065,N_26538);
and U27626 (N_27626,N_27304,N_27410);
nor U27627 (N_27627,N_27460,N_27014);
nor U27628 (N_27628,N_26919,N_26883);
nand U27629 (N_27629,N_27548,N_26417);
xnor U27630 (N_27630,N_26584,N_26780);
or U27631 (N_27631,N_27566,N_26456);
and U27632 (N_27632,N_27164,N_27273);
or U27633 (N_27633,N_26844,N_27114);
nor U27634 (N_27634,N_26922,N_26664);
nor U27635 (N_27635,N_26419,N_27507);
xnor U27636 (N_27636,N_27216,N_26586);
xnor U27637 (N_27637,N_27153,N_26736);
xor U27638 (N_27638,N_27592,N_26639);
or U27639 (N_27639,N_27349,N_27323);
xnor U27640 (N_27640,N_26528,N_26472);
nand U27641 (N_27641,N_27480,N_26480);
xor U27642 (N_27642,N_26868,N_27265);
or U27643 (N_27643,N_27158,N_26520);
and U27644 (N_27644,N_27524,N_27557);
or U27645 (N_27645,N_26734,N_26455);
xnor U27646 (N_27646,N_26517,N_26614);
xor U27647 (N_27647,N_27040,N_26847);
xor U27648 (N_27648,N_26557,N_26596);
and U27649 (N_27649,N_26934,N_26860);
or U27650 (N_27650,N_27327,N_27166);
xor U27651 (N_27651,N_26928,N_27443);
xor U27652 (N_27652,N_27174,N_27492);
and U27653 (N_27653,N_26826,N_27481);
or U27654 (N_27654,N_27512,N_27383);
and U27655 (N_27655,N_27084,N_26463);
or U27656 (N_27656,N_27585,N_27253);
nor U27657 (N_27657,N_26935,N_27430);
nand U27658 (N_27658,N_27280,N_26608);
nor U27659 (N_27659,N_27229,N_27154);
xnor U27660 (N_27660,N_26579,N_27337);
nand U27661 (N_27661,N_26949,N_27428);
xor U27662 (N_27662,N_27539,N_26406);
nor U27663 (N_27663,N_27057,N_27113);
nor U27664 (N_27664,N_26862,N_27161);
nand U27665 (N_27665,N_26763,N_26937);
nor U27666 (N_27666,N_27300,N_26749);
nand U27667 (N_27667,N_27266,N_27574);
nand U27668 (N_27668,N_26912,N_27187);
xor U27669 (N_27669,N_27434,N_26682);
nand U27670 (N_27670,N_26481,N_26485);
nor U27671 (N_27671,N_27311,N_26569);
xor U27672 (N_27672,N_27591,N_27450);
or U27673 (N_27673,N_27313,N_26953);
or U27674 (N_27674,N_27307,N_26651);
xor U27675 (N_27675,N_27499,N_26894);
nand U27676 (N_27676,N_26606,N_26719);
nand U27677 (N_27677,N_26773,N_27309);
and U27678 (N_27678,N_26574,N_26727);
and U27679 (N_27679,N_26701,N_26662);
nand U27680 (N_27680,N_26667,N_26654);
nand U27681 (N_27681,N_26439,N_26429);
nand U27682 (N_27682,N_27598,N_26938);
and U27683 (N_27683,N_26403,N_27199);
xnor U27684 (N_27684,N_27554,N_27396);
xnor U27685 (N_27685,N_27294,N_26505);
nor U27686 (N_27686,N_26856,N_27146);
nand U27687 (N_27687,N_27226,N_26723);
and U27688 (N_27688,N_26422,N_27124);
or U27689 (N_27689,N_26492,N_27320);
xnor U27690 (N_27690,N_27447,N_27052);
and U27691 (N_27691,N_27193,N_26550);
and U27692 (N_27692,N_27236,N_27206);
and U27693 (N_27693,N_27299,N_27155);
nand U27694 (N_27694,N_26986,N_26663);
or U27695 (N_27695,N_27485,N_27425);
and U27696 (N_27696,N_26991,N_26726);
nor U27697 (N_27697,N_26902,N_26426);
xor U27698 (N_27698,N_27330,N_27473);
and U27699 (N_27699,N_26687,N_27175);
nor U27700 (N_27700,N_27575,N_27017);
xnor U27701 (N_27701,N_27582,N_27493);
nor U27702 (N_27702,N_27092,N_27185);
xor U27703 (N_27703,N_26739,N_26743);
xnor U27704 (N_27704,N_27212,N_26781);
nor U27705 (N_27705,N_26612,N_27308);
nand U27706 (N_27706,N_26814,N_27532);
xor U27707 (N_27707,N_26600,N_26899);
nor U27708 (N_27708,N_27438,N_27469);
and U27709 (N_27709,N_26762,N_27517);
nor U27710 (N_27710,N_26836,N_26760);
nand U27711 (N_27711,N_27202,N_27271);
nor U27712 (N_27712,N_27244,N_26661);
nand U27713 (N_27713,N_26776,N_27415);
xor U27714 (N_27714,N_26904,N_26944);
and U27715 (N_27715,N_27409,N_27587);
and U27716 (N_27716,N_27569,N_26959);
and U27717 (N_27717,N_26696,N_27108);
and U27718 (N_27718,N_27044,N_27412);
nor U27719 (N_27719,N_27191,N_27468);
nor U27720 (N_27720,N_26804,N_27059);
xor U27721 (N_27721,N_27179,N_26437);
nand U27722 (N_27722,N_26909,N_27370);
and U27723 (N_27723,N_27351,N_27118);
nor U27724 (N_27724,N_27249,N_27208);
nor U27725 (N_27725,N_27018,N_26489);
xor U27726 (N_27726,N_26799,N_26445);
nand U27727 (N_27727,N_27382,N_27264);
or U27728 (N_27728,N_27426,N_27386);
or U27729 (N_27729,N_27560,N_26642);
xnor U27730 (N_27730,N_27007,N_26930);
and U27731 (N_27731,N_27501,N_26594);
xor U27732 (N_27732,N_27207,N_26578);
xnor U27733 (N_27733,N_26432,N_27344);
nor U27734 (N_27734,N_27322,N_27378);
nand U27735 (N_27735,N_26977,N_26857);
or U27736 (N_27736,N_27567,N_26607);
and U27737 (N_27737,N_27286,N_26895);
xnor U27738 (N_27738,N_27228,N_26777);
nand U27739 (N_27739,N_27004,N_27023);
nor U27740 (N_27740,N_26752,N_27270);
xnor U27741 (N_27741,N_26806,N_26646);
and U27742 (N_27742,N_27235,N_27522);
nor U27743 (N_27743,N_26533,N_26631);
nor U27744 (N_27744,N_26729,N_27488);
and U27745 (N_27745,N_27533,N_26716);
or U27746 (N_27746,N_27119,N_27197);
or U27747 (N_27747,N_26689,N_26995);
nand U27748 (N_27748,N_26989,N_27455);
and U27749 (N_27749,N_27534,N_27461);
nand U27750 (N_27750,N_26629,N_27060);
nand U27751 (N_27751,N_26573,N_27090);
or U27752 (N_27752,N_27291,N_27435);
nor U27753 (N_27753,N_27503,N_26658);
or U27754 (N_27754,N_27218,N_27366);
nor U27755 (N_27755,N_27094,N_26675);
nor U27756 (N_27756,N_27016,N_27494);
nand U27757 (N_27757,N_27462,N_26801);
nand U27758 (N_27758,N_26441,N_26873);
and U27759 (N_27759,N_26495,N_27359);
or U27760 (N_27760,N_26908,N_26459);
nor U27761 (N_27761,N_27105,N_27186);
nand U27762 (N_27762,N_26979,N_26917);
and U27763 (N_27763,N_27288,N_27422);
xor U27764 (N_27764,N_26807,N_26686);
xnor U27765 (N_27765,N_27545,N_27596);
or U27766 (N_27766,N_26731,N_26870);
xor U27767 (N_27767,N_26951,N_27203);
and U27768 (N_27768,N_26939,N_26575);
nand U27769 (N_27769,N_26706,N_26724);
nand U27770 (N_27770,N_26464,N_27506);
nand U27771 (N_27771,N_27163,N_26643);
or U27772 (N_27772,N_27131,N_27170);
nand U27773 (N_27773,N_27247,N_27472);
nor U27774 (N_27774,N_27325,N_26973);
xnor U27775 (N_27775,N_26747,N_27256);
or U27776 (N_27776,N_26601,N_27317);
or U27777 (N_27777,N_26774,N_26637);
nor U27778 (N_27778,N_27268,N_26741);
or U27779 (N_27779,N_26595,N_26451);
nand U27780 (N_27780,N_26821,N_26683);
xnor U27781 (N_27781,N_27275,N_26656);
nand U27782 (N_27782,N_27211,N_27348);
or U27783 (N_27783,N_27568,N_27022);
nand U27784 (N_27784,N_26698,N_26442);
and U27785 (N_27785,N_27593,N_26992);
nor U27786 (N_27786,N_26843,N_27306);
and U27787 (N_27787,N_26420,N_26404);
or U27788 (N_27788,N_26660,N_26770);
xor U27789 (N_27789,N_27096,N_26745);
nor U27790 (N_27790,N_26418,N_26925);
and U27791 (N_27791,N_26858,N_27579);
or U27792 (N_27792,N_26808,N_27448);
xor U27793 (N_27793,N_26571,N_27260);
nor U27794 (N_27794,N_26782,N_27089);
or U27795 (N_27795,N_26513,N_27282);
and U27796 (N_27796,N_27586,N_27132);
nand U27797 (N_27797,N_26544,N_27475);
xnor U27798 (N_27798,N_26630,N_27000);
and U27799 (N_27799,N_27254,N_27429);
nor U27800 (N_27800,N_27541,N_27402);
or U27801 (N_27801,N_26474,N_27451);
nor U27802 (N_27802,N_26748,N_26669);
or U27803 (N_27803,N_27332,N_26755);
or U27804 (N_27804,N_26691,N_27055);
xor U27805 (N_27805,N_27068,N_27230);
nor U27806 (N_27806,N_26604,N_26988);
xor U27807 (N_27807,N_27156,N_27053);
or U27808 (N_27808,N_26684,N_27357);
nor U27809 (N_27809,N_26620,N_27576);
nor U27810 (N_27810,N_26576,N_26876);
and U27811 (N_27811,N_27081,N_26649);
or U27812 (N_27812,N_27145,N_27246);
nor U27813 (N_27813,N_27437,N_26703);
nand U27814 (N_27814,N_26981,N_27599);
and U27815 (N_27815,N_26737,N_26623);
and U27816 (N_27816,N_27038,N_27571);
xor U27817 (N_27817,N_26446,N_26478);
xor U27818 (N_27818,N_27528,N_27025);
xnor U27819 (N_27819,N_27276,N_27008);
and U27820 (N_27820,N_26652,N_27142);
or U27821 (N_27821,N_27261,N_26511);
nand U27822 (N_27822,N_27381,N_26408);
and U27823 (N_27823,N_27086,N_26458);
xnor U27824 (N_27824,N_27367,N_26712);
or U27825 (N_27825,N_26761,N_26440);
nor U27826 (N_27826,N_26920,N_27459);
nand U27827 (N_27827,N_26583,N_27594);
nor U27828 (N_27828,N_26725,N_27223);
or U27829 (N_27829,N_27389,N_26779);
and U27830 (N_27830,N_27151,N_26592);
xor U27831 (N_27831,N_26966,N_27400);
xor U27832 (N_27832,N_27563,N_27103);
and U27833 (N_27833,N_27401,N_27336);
xnor U27834 (N_27834,N_26710,N_26657);
and U27835 (N_27835,N_27037,N_26428);
nor U27836 (N_27836,N_27172,N_27406);
xnor U27837 (N_27837,N_26674,N_26888);
nor U27838 (N_27838,N_26695,N_27178);
nor U27839 (N_27839,N_26536,N_27436);
or U27840 (N_27840,N_27183,N_26733);
nand U27841 (N_27841,N_27006,N_27267);
or U27842 (N_27842,N_26926,N_26628);
or U27843 (N_27843,N_26416,N_26722);
or U27844 (N_27844,N_27421,N_27075);
and U27845 (N_27845,N_27379,N_26769);
xnor U27846 (N_27846,N_26941,N_26816);
xnor U27847 (N_27847,N_26602,N_27516);
nand U27848 (N_27848,N_27141,N_27125);
nor U27849 (N_27849,N_27015,N_26906);
or U27850 (N_27850,N_27143,N_26792);
nand U27851 (N_27851,N_26615,N_27106);
or U27852 (N_27852,N_26508,N_26835);
or U27853 (N_27853,N_26950,N_27101);
nand U27854 (N_27854,N_27550,N_26443);
nor U27855 (N_27855,N_27529,N_26448);
xnor U27856 (N_27856,N_26984,N_26958);
nand U27857 (N_27857,N_26470,N_26855);
nand U27858 (N_27858,N_26924,N_27418);
or U27859 (N_27859,N_26491,N_27510);
and U27860 (N_27860,N_26570,N_26677);
and U27861 (N_27861,N_27478,N_26811);
nor U27862 (N_27862,N_27063,N_26700);
nor U27863 (N_27863,N_26540,N_26846);
or U27864 (N_27864,N_27058,N_26903);
nand U27865 (N_27865,N_27046,N_26982);
xnor U27866 (N_27866,N_27028,N_27444);
and U27867 (N_27867,N_27369,N_26539);
nand U27868 (N_27868,N_27149,N_27272);
or U27869 (N_27869,N_27215,N_27466);
and U27870 (N_27870,N_27021,N_26410);
xnor U27871 (N_27871,N_26956,N_26590);
nand U27872 (N_27872,N_27390,N_27589);
nand U27873 (N_27873,N_27511,N_27128);
nand U27874 (N_27874,N_26499,N_27420);
nor U27875 (N_27875,N_26787,N_27027);
or U27876 (N_27876,N_27210,N_26659);
or U27877 (N_27877,N_26940,N_26564);
nor U27878 (N_27878,N_26522,N_27521);
or U27879 (N_27879,N_26872,N_27490);
or U27880 (N_27880,N_26766,N_27546);
nor U27881 (N_27881,N_27252,N_26409);
xnor U27882 (N_27882,N_27077,N_26435);
nor U27883 (N_27883,N_27171,N_27117);
or U27884 (N_27884,N_26599,N_26845);
nor U27885 (N_27885,N_26778,N_27391);
or U27886 (N_27886,N_27150,N_26892);
and U27887 (N_27887,N_27380,N_27069);
and U27888 (N_27888,N_27441,N_27495);
and U27889 (N_27889,N_27479,N_26510);
nor U27890 (N_27890,N_26556,N_26972);
nand U27891 (N_27891,N_26795,N_26916);
and U27892 (N_27892,N_27375,N_26971);
nand U27893 (N_27893,N_26482,N_27255);
nor U27894 (N_27894,N_27220,N_26504);
nor U27895 (N_27895,N_27281,N_26962);
and U27896 (N_27896,N_26655,N_26771);
and U27897 (N_27897,N_26853,N_27312);
or U27898 (N_27898,N_26918,N_27347);
nor U27899 (N_27899,N_26534,N_26923);
and U27900 (N_27900,N_27561,N_26460);
and U27901 (N_27901,N_26775,N_26869);
and U27902 (N_27902,N_27167,N_26886);
and U27903 (N_27903,N_27147,N_27180);
or U27904 (N_27904,N_27368,N_27126);
nor U27905 (N_27905,N_26670,N_26530);
xor U27906 (N_27906,N_27338,N_27543);
or U27907 (N_27907,N_27595,N_27542);
xnor U27908 (N_27908,N_26679,N_27487);
and U27909 (N_27909,N_27413,N_26588);
nand U27910 (N_27910,N_26468,N_26751);
or U27911 (N_27911,N_26882,N_26688);
xor U27912 (N_27912,N_27583,N_26993);
or U27913 (N_27913,N_27283,N_27250);
nand U27914 (N_27914,N_27514,N_27284);
and U27915 (N_27915,N_27279,N_27572);
and U27916 (N_27916,N_27549,N_27064);
nand U27917 (N_27917,N_27240,N_26818);
nor U27918 (N_27918,N_26697,N_27361);
nor U27919 (N_27919,N_26673,N_26401);
or U27920 (N_27920,N_26735,N_27201);
xor U27921 (N_27921,N_26535,N_27169);
nor U27922 (N_27922,N_26598,N_26547);
nor U27923 (N_27923,N_26405,N_27245);
nor U27924 (N_27924,N_27237,N_26512);
xor U27925 (N_27925,N_26788,N_27019);
nand U27926 (N_27926,N_26822,N_26852);
nor U27927 (N_27927,N_27036,N_26503);
nand U27928 (N_27928,N_26627,N_26493);
xnor U27929 (N_27929,N_26466,N_26831);
nand U27930 (N_27930,N_26415,N_26929);
nor U27931 (N_27931,N_27477,N_26625);
or U27932 (N_27932,N_27474,N_26605);
nand U27933 (N_27933,N_26425,N_26653);
nand U27934 (N_27934,N_26562,N_27054);
nand U27935 (N_27935,N_27032,N_27165);
xor U27936 (N_27936,N_26692,N_27130);
nor U27937 (N_27937,N_26665,N_26497);
nand U27938 (N_27938,N_26915,N_26985);
or U27939 (N_27939,N_26825,N_26753);
xnor U27940 (N_27940,N_26681,N_26438);
nand U27941 (N_27941,N_27408,N_27520);
and U27942 (N_27942,N_26759,N_26402);
nand U27943 (N_27943,N_26568,N_27302);
nor U27944 (N_27944,N_26559,N_27024);
and U27945 (N_27945,N_26803,N_27500);
xor U27946 (N_27946,N_26449,N_27535);
nor U27947 (N_27947,N_27009,N_27373);
xnor U27948 (N_27948,N_26946,N_27050);
or U27949 (N_27949,N_26794,N_27452);
nand U27950 (N_27950,N_26819,N_26490);
or U27951 (N_27951,N_27352,N_26893);
and U27952 (N_27952,N_26476,N_27123);
or U27953 (N_27953,N_27134,N_27570);
and U27954 (N_27954,N_27305,N_26936);
xnor U27955 (N_27955,N_26975,N_27289);
xor U27956 (N_27956,N_27047,N_27177);
or U27957 (N_27957,N_27358,N_27397);
xor U27958 (N_27958,N_27353,N_26603);
xor U27959 (N_27959,N_26713,N_26514);
and U27960 (N_27960,N_27354,N_26859);
and U27961 (N_27961,N_26558,N_26577);
xor U27962 (N_27962,N_27467,N_26947);
nand U27963 (N_27963,N_27555,N_27588);
and U27964 (N_27964,N_27440,N_26638);
xnor U27965 (N_27965,N_26467,N_27465);
and U27966 (N_27966,N_26911,N_27527);
xnor U27967 (N_27967,N_27231,N_27098);
and U27968 (N_27968,N_26650,N_27301);
nand U27969 (N_27969,N_26720,N_27394);
xor U27970 (N_27970,N_27363,N_26943);
nand U27971 (N_27971,N_27597,N_26680);
nand U27972 (N_27972,N_27107,N_26509);
or U27973 (N_27973,N_27076,N_27251);
nor U27974 (N_27974,N_27135,N_27048);
and U27975 (N_27975,N_26672,N_27102);
and U27976 (N_27976,N_27026,N_27372);
nand U27977 (N_27977,N_26851,N_26864);
xnor U27978 (N_27978,N_26532,N_27136);
nor U27979 (N_27979,N_27439,N_27504);
nand U27980 (N_27980,N_26955,N_27427);
nor U27981 (N_27981,N_26832,N_26524);
or U27982 (N_27982,N_26848,N_26619);
xnor U27983 (N_27983,N_27340,N_26910);
nand U27984 (N_27984,N_27013,N_27335);
xnor U27985 (N_27985,N_26552,N_26411);
nand U27986 (N_27986,N_27297,N_26526);
and U27987 (N_27987,N_26541,N_27292);
xnor U27988 (N_27988,N_27293,N_27195);
and U27989 (N_27989,N_27398,N_26454);
and U27990 (N_27990,N_26580,N_27377);
or U27991 (N_27991,N_26507,N_27259);
nand U27992 (N_27992,N_27263,N_26473);
nor U27993 (N_27993,N_27062,N_26891);
xnor U27994 (N_27994,N_27031,N_26519);
nor U27995 (N_27995,N_27454,N_26897);
nand U27996 (N_27996,N_26863,N_26496);
or U27997 (N_27997,N_27219,N_26833);
or U27998 (N_27998,N_27115,N_27556);
nand U27999 (N_27999,N_27192,N_26900);
nor U28000 (N_28000,N_26756,N_26690);
nand U28001 (N_28001,N_26800,N_26715);
nand U28002 (N_28002,N_27221,N_27257);
nor U28003 (N_28003,N_27329,N_26593);
nor U28004 (N_28004,N_27039,N_26444);
nand U28005 (N_28005,N_27464,N_26502);
or U28006 (N_28006,N_27388,N_26462);
xnor U28007 (N_28007,N_26823,N_27278);
nor U28008 (N_28008,N_27148,N_27239);
and U28009 (N_28009,N_27416,N_27404);
or U28010 (N_28010,N_26622,N_26998);
xor U28011 (N_28011,N_27489,N_26815);
or U28012 (N_28012,N_27168,N_26987);
or U28013 (N_28013,N_27509,N_27122);
nor U28014 (N_28014,N_26527,N_27326);
nor U28015 (N_28015,N_27184,N_27314);
nor U28016 (N_28016,N_27233,N_26610);
nor U28017 (N_28017,N_26704,N_26702);
xor U28018 (N_28018,N_26500,N_27112);
nand U28019 (N_28019,N_26543,N_27395);
and U28020 (N_28020,N_26699,N_26830);
nand U28021 (N_28021,N_26561,N_27296);
and U28022 (N_28022,N_27424,N_27020);
nand U28023 (N_28023,N_27316,N_26783);
nand U28024 (N_28024,N_27225,N_27071);
xnor U28025 (N_28025,N_26790,N_26447);
and U28026 (N_28026,N_26732,N_26591);
xor U28027 (N_28027,N_26521,N_27190);
nor U28028 (N_28028,N_26913,N_27033);
nand U28029 (N_28029,N_27070,N_26636);
and U28030 (N_28030,N_27432,N_26791);
or U28031 (N_28031,N_26879,N_27573);
xor U28032 (N_28032,N_27111,N_26840);
and U28033 (N_28033,N_27277,N_26430);
nor U28034 (N_28034,N_27523,N_26764);
and U28035 (N_28035,N_27088,N_27011);
or U28036 (N_28036,N_27005,N_27310);
nor U28037 (N_28037,N_26400,N_27162);
or U28038 (N_28038,N_26621,N_26671);
and U28039 (N_28039,N_26611,N_26849);
nor U28040 (N_28040,N_27584,N_26738);
nand U28041 (N_28041,N_27222,N_26714);
nor U28042 (N_28042,N_26837,N_26767);
and U28043 (N_28043,N_26563,N_26980);
and U28044 (N_28044,N_26640,N_26878);
or U28045 (N_28045,N_26453,N_26957);
and U28046 (N_28046,N_26968,N_27100);
nand U28047 (N_28047,N_27129,N_27558);
and U28048 (N_28048,N_26880,N_26644);
or U28049 (N_28049,N_27341,N_26613);
nor U28050 (N_28050,N_27189,N_26553);
nor U28051 (N_28051,N_26785,N_27356);
nor U28052 (N_28052,N_27385,N_27496);
or U28053 (N_28053,N_27144,N_27333);
nor U28054 (N_28054,N_27003,N_27298);
nand U28055 (N_28055,N_27483,N_26865);
xor U28056 (N_28056,N_27453,N_26567);
or U28057 (N_28057,N_27238,N_26666);
nor U28058 (N_28058,N_26572,N_27224);
nor U28059 (N_28059,N_26952,N_26765);
and U28060 (N_28060,N_27095,N_27099);
nand U28061 (N_28061,N_26452,N_26494);
xor U28062 (N_28062,N_26963,N_27433);
xor U28063 (N_28063,N_27303,N_27067);
xnor U28064 (N_28064,N_26772,N_26875);
xor U28065 (N_28065,N_26498,N_27387);
or U28066 (N_28066,N_26817,N_26828);
xor U28067 (N_28067,N_26746,N_27525);
xor U28068 (N_28068,N_27319,N_27328);
xnor U28069 (N_28069,N_26990,N_26506);
or U28070 (N_28070,N_26555,N_26546);
nor U28071 (N_28071,N_27577,N_26932);
nand U28072 (N_28072,N_27414,N_27030);
and U28073 (N_28073,N_26471,N_27552);
nand U28074 (N_28074,N_27258,N_26901);
or U28075 (N_28075,N_27091,N_27565);
nor U28076 (N_28076,N_26708,N_27159);
nor U28077 (N_28077,N_26548,N_26589);
nor U28078 (N_28078,N_27034,N_26768);
and U28079 (N_28079,N_27157,N_27127);
nand U28080 (N_28080,N_26618,N_26413);
or U28081 (N_28081,N_26634,N_26529);
nand U28082 (N_28082,N_26711,N_26421);
xnor U28083 (N_28083,N_27376,N_27419);
nand U28084 (N_28084,N_27074,N_26709);
nand U28085 (N_28085,N_26931,N_26812);
and U28086 (N_28086,N_26565,N_27559);
or U28087 (N_28087,N_27133,N_26730);
nand U28088 (N_28088,N_27188,N_26997);
or U28089 (N_28089,N_26890,N_27140);
or U28090 (N_28090,N_27508,N_27362);
and U28091 (N_28091,N_27321,N_27085);
or U28092 (N_28092,N_27080,N_27083);
xor U28093 (N_28093,N_26585,N_26479);
and U28094 (N_28094,N_27384,N_27551);
nor U28095 (N_28095,N_26537,N_26945);
nor U28096 (N_28096,N_27110,N_27423);
or U28097 (N_28097,N_26624,N_27411);
and U28098 (N_28098,N_27079,N_27137);
or U28099 (N_28099,N_26867,N_26974);
and U28100 (N_28100,N_26810,N_27139);
and U28101 (N_28101,N_26647,N_26921);
nor U28102 (N_28102,N_27365,N_27502);
nor U28103 (N_28103,N_26983,N_26566);
nor U28104 (N_28104,N_27041,N_26881);
xor U28105 (N_28105,N_26827,N_26874);
or U28106 (N_28106,N_26633,N_27160);
or U28107 (N_28107,N_26842,N_27526);
and U28108 (N_28108,N_27072,N_27318);
xnor U28109 (N_28109,N_26805,N_26964);
or U28110 (N_28110,N_26797,N_27505);
and U28111 (N_28111,N_26518,N_27181);
nor U28112 (N_28112,N_27331,N_27553);
xnor U28113 (N_28113,N_27431,N_26798);
nand U28114 (N_28114,N_27486,N_26996);
xor U28115 (N_28115,N_26960,N_27343);
nand U28116 (N_28116,N_26898,N_26976);
or U28117 (N_28117,N_27078,N_26705);
nor U28118 (N_28118,N_27290,N_26970);
xor U28119 (N_28119,N_26861,N_27476);
xor U28120 (N_28120,N_27204,N_26616);
xor U28121 (N_28121,N_27051,N_27497);
xnor U28122 (N_28122,N_27471,N_27393);
nor U28123 (N_28123,N_27001,N_26809);
nor U28124 (N_28124,N_27029,N_27536);
nand U28125 (N_28125,N_27484,N_26969);
and U28126 (N_28126,N_26597,N_26871);
xor U28127 (N_28127,N_26641,N_26841);
or U28128 (N_28128,N_26407,N_26515);
nand U28129 (N_28129,N_27109,N_27360);
nand U28130 (N_28130,N_27182,N_26469);
nand U28131 (N_28131,N_27104,N_27061);
nor U28132 (N_28132,N_26786,N_27564);
and U28133 (N_28133,N_26961,N_26678);
and U28134 (N_28134,N_27035,N_26889);
nand U28135 (N_28135,N_27446,N_26728);
nand U28136 (N_28136,N_26587,N_26838);
xnor U28137 (N_28137,N_26483,N_26721);
xor U28138 (N_28138,N_27334,N_26626);
xnor U28139 (N_28139,N_27287,N_27087);
and U28140 (N_28140,N_27217,N_26758);
nor U28141 (N_28141,N_27350,N_27531);
and U28142 (N_28142,N_27392,N_26617);
nor U28143 (N_28143,N_26648,N_26465);
nand U28144 (N_28144,N_26523,N_26887);
nand U28145 (N_28145,N_27519,N_26412);
nand U28146 (N_28146,N_26907,N_26549);
or U28147 (N_28147,N_26707,N_27515);
nor U28148 (N_28148,N_27295,N_27513);
or U28149 (N_28149,N_26582,N_26885);
xor U28150 (N_28150,N_26414,N_26685);
nor U28151 (N_28151,N_27066,N_27364);
xor U28152 (N_28152,N_26531,N_26948);
and U28153 (N_28153,N_26999,N_27012);
and U28154 (N_28154,N_27445,N_26676);
and U28155 (N_28155,N_27120,N_26461);
or U28156 (N_28156,N_26484,N_26927);
or U28157 (N_28157,N_27315,N_27002);
nand U28158 (N_28158,N_27093,N_27045);
xor U28159 (N_28159,N_27580,N_27227);
xnor U28160 (N_28160,N_27371,N_27581);
nand U28161 (N_28161,N_26965,N_27209);
and U28162 (N_28162,N_26434,N_26450);
nand U28163 (N_28163,N_26820,N_27540);
or U28164 (N_28164,N_27234,N_26717);
xnor U28165 (N_28165,N_26551,N_26635);
or U28166 (N_28166,N_27269,N_26560);
nand U28167 (N_28167,N_26516,N_27590);
nor U28168 (N_28168,N_27403,N_26854);
or U28169 (N_28169,N_27491,N_26905);
nor U28170 (N_28170,N_26694,N_26834);
nor U28171 (N_28171,N_26793,N_26609);
nand U28172 (N_28172,N_27097,N_27152);
xnor U28173 (N_28173,N_27457,N_27138);
or U28174 (N_28174,N_27458,N_27274);
or U28175 (N_28175,N_27243,N_26423);
and U28176 (N_28176,N_27056,N_26542);
and U28177 (N_28177,N_26994,N_26487);
or U28178 (N_28178,N_27442,N_26545);
nand U28179 (N_28179,N_27205,N_27116);
and U28180 (N_28180,N_27194,N_27010);
nand U28181 (N_28181,N_26457,N_27176);
or U28182 (N_28182,N_26789,N_26424);
or U28183 (N_28183,N_26754,N_27405);
nand U28184 (N_28184,N_27538,N_26796);
or U28185 (N_28185,N_27407,N_27482);
and U28186 (N_28186,N_27242,N_27082);
or U28187 (N_28187,N_27232,N_26501);
nor U28188 (N_28188,N_26742,N_26740);
nor U28189 (N_28189,N_26866,N_26750);
nor U28190 (N_28190,N_27248,N_26693);
nand U28191 (N_28191,N_27324,N_26967);
xor U28192 (N_28192,N_26784,N_26477);
xor U28193 (N_28193,N_27374,N_27342);
nor U28194 (N_28194,N_27173,N_26942);
nand U28195 (N_28195,N_26829,N_27042);
nor U28196 (N_28196,N_27214,N_26475);
nand U28197 (N_28197,N_27399,N_26839);
or U28198 (N_28198,N_26486,N_26824);
nor U28199 (N_28199,N_26436,N_27285);
and U28200 (N_28200,N_27344,N_26499);
and U28201 (N_28201,N_27493,N_27199);
nand U28202 (N_28202,N_26881,N_27083);
nor U28203 (N_28203,N_27144,N_26832);
nand U28204 (N_28204,N_27248,N_27533);
or U28205 (N_28205,N_26973,N_27027);
and U28206 (N_28206,N_26452,N_26916);
nor U28207 (N_28207,N_26445,N_27567);
xor U28208 (N_28208,N_26852,N_27111);
or U28209 (N_28209,N_27462,N_27543);
nand U28210 (N_28210,N_26469,N_26947);
nand U28211 (N_28211,N_27503,N_26465);
and U28212 (N_28212,N_26400,N_26828);
nand U28213 (N_28213,N_27575,N_27247);
or U28214 (N_28214,N_26669,N_26784);
nand U28215 (N_28215,N_26437,N_26908);
or U28216 (N_28216,N_26976,N_27338);
xnor U28217 (N_28217,N_27423,N_27300);
nor U28218 (N_28218,N_27597,N_26423);
or U28219 (N_28219,N_27520,N_26570);
and U28220 (N_28220,N_27193,N_27371);
nor U28221 (N_28221,N_27020,N_26579);
xnor U28222 (N_28222,N_27579,N_27349);
nand U28223 (N_28223,N_27296,N_27058);
or U28224 (N_28224,N_27242,N_27073);
nand U28225 (N_28225,N_27179,N_27441);
nor U28226 (N_28226,N_26608,N_26708);
nand U28227 (N_28227,N_27407,N_27373);
nand U28228 (N_28228,N_26619,N_26908);
or U28229 (N_28229,N_26575,N_27159);
or U28230 (N_28230,N_26744,N_26555);
xor U28231 (N_28231,N_27289,N_27209);
or U28232 (N_28232,N_26863,N_26983);
xnor U28233 (N_28233,N_27222,N_26825);
nor U28234 (N_28234,N_27346,N_27493);
or U28235 (N_28235,N_27545,N_26946);
and U28236 (N_28236,N_26939,N_27015);
or U28237 (N_28237,N_27357,N_26625);
xnor U28238 (N_28238,N_26704,N_26643);
nand U28239 (N_28239,N_26869,N_26853);
and U28240 (N_28240,N_26550,N_26420);
nor U28241 (N_28241,N_26973,N_26440);
nor U28242 (N_28242,N_26596,N_26549);
nand U28243 (N_28243,N_26526,N_26897);
nand U28244 (N_28244,N_26603,N_27358);
xor U28245 (N_28245,N_27038,N_27155);
xnor U28246 (N_28246,N_27417,N_26868);
nand U28247 (N_28247,N_26460,N_27056);
xor U28248 (N_28248,N_26753,N_27257);
nor U28249 (N_28249,N_27162,N_26636);
nor U28250 (N_28250,N_27169,N_27186);
and U28251 (N_28251,N_27072,N_26950);
xor U28252 (N_28252,N_27513,N_26774);
and U28253 (N_28253,N_26927,N_27288);
nand U28254 (N_28254,N_26872,N_27171);
or U28255 (N_28255,N_26450,N_27247);
and U28256 (N_28256,N_26800,N_27056);
nand U28257 (N_28257,N_27248,N_26983);
nor U28258 (N_28258,N_27208,N_27308);
and U28259 (N_28259,N_27227,N_26696);
or U28260 (N_28260,N_27368,N_26788);
or U28261 (N_28261,N_27324,N_26737);
nor U28262 (N_28262,N_26567,N_27210);
nor U28263 (N_28263,N_27458,N_27474);
nand U28264 (N_28264,N_26606,N_27579);
nor U28265 (N_28265,N_27558,N_27184);
or U28266 (N_28266,N_27578,N_26893);
nand U28267 (N_28267,N_26905,N_27097);
nor U28268 (N_28268,N_27383,N_26677);
nor U28269 (N_28269,N_27583,N_27592);
and U28270 (N_28270,N_27548,N_27236);
nor U28271 (N_28271,N_27479,N_27489);
nand U28272 (N_28272,N_26418,N_27227);
and U28273 (N_28273,N_26679,N_27530);
nand U28274 (N_28274,N_26675,N_27255);
xnor U28275 (N_28275,N_26445,N_27391);
and U28276 (N_28276,N_26624,N_27204);
and U28277 (N_28277,N_27004,N_26901);
or U28278 (N_28278,N_27272,N_27223);
xor U28279 (N_28279,N_26416,N_26620);
and U28280 (N_28280,N_26555,N_27193);
nand U28281 (N_28281,N_26771,N_27212);
or U28282 (N_28282,N_27123,N_27005);
and U28283 (N_28283,N_26554,N_26531);
nand U28284 (N_28284,N_27386,N_26509);
nor U28285 (N_28285,N_26428,N_26784);
or U28286 (N_28286,N_27154,N_27425);
nand U28287 (N_28287,N_26739,N_26407);
nor U28288 (N_28288,N_26870,N_27589);
nor U28289 (N_28289,N_26572,N_26943);
nand U28290 (N_28290,N_27182,N_26904);
and U28291 (N_28291,N_27017,N_27407);
and U28292 (N_28292,N_26619,N_26643);
and U28293 (N_28293,N_27495,N_27425);
xnor U28294 (N_28294,N_26811,N_26455);
nand U28295 (N_28295,N_26450,N_27345);
nand U28296 (N_28296,N_27425,N_27382);
and U28297 (N_28297,N_26919,N_27310);
nor U28298 (N_28298,N_27237,N_27474);
nor U28299 (N_28299,N_26670,N_26985);
xor U28300 (N_28300,N_27222,N_26454);
or U28301 (N_28301,N_27252,N_27211);
and U28302 (N_28302,N_27372,N_27062);
xor U28303 (N_28303,N_26667,N_26808);
or U28304 (N_28304,N_27146,N_27008);
xnor U28305 (N_28305,N_27469,N_26434);
or U28306 (N_28306,N_27291,N_27525);
nand U28307 (N_28307,N_26664,N_26914);
and U28308 (N_28308,N_27295,N_26464);
nand U28309 (N_28309,N_27525,N_26688);
nand U28310 (N_28310,N_27574,N_27092);
or U28311 (N_28311,N_26675,N_26684);
or U28312 (N_28312,N_26647,N_27155);
or U28313 (N_28313,N_27250,N_26951);
or U28314 (N_28314,N_26985,N_27323);
and U28315 (N_28315,N_27170,N_27100);
or U28316 (N_28316,N_27164,N_26444);
nand U28317 (N_28317,N_26735,N_26950);
nand U28318 (N_28318,N_26971,N_27286);
or U28319 (N_28319,N_26675,N_27241);
and U28320 (N_28320,N_27452,N_26752);
nand U28321 (N_28321,N_26658,N_27082);
nand U28322 (N_28322,N_26444,N_26941);
or U28323 (N_28323,N_26436,N_26466);
nand U28324 (N_28324,N_27141,N_26410);
and U28325 (N_28325,N_27077,N_26412);
and U28326 (N_28326,N_27346,N_26474);
and U28327 (N_28327,N_26626,N_26630);
and U28328 (N_28328,N_26794,N_26664);
or U28329 (N_28329,N_27543,N_27261);
nor U28330 (N_28330,N_27459,N_27182);
and U28331 (N_28331,N_26644,N_27546);
or U28332 (N_28332,N_26943,N_26744);
xnor U28333 (N_28333,N_27327,N_27565);
xnor U28334 (N_28334,N_26654,N_27058);
and U28335 (N_28335,N_26655,N_27493);
nor U28336 (N_28336,N_26496,N_27081);
or U28337 (N_28337,N_27454,N_26551);
and U28338 (N_28338,N_26913,N_27431);
and U28339 (N_28339,N_27356,N_26843);
or U28340 (N_28340,N_26803,N_26618);
nor U28341 (N_28341,N_27091,N_26789);
xnor U28342 (N_28342,N_26963,N_27334);
nand U28343 (N_28343,N_27022,N_26737);
and U28344 (N_28344,N_27114,N_27179);
nor U28345 (N_28345,N_27251,N_26748);
nor U28346 (N_28346,N_27257,N_27189);
and U28347 (N_28347,N_27495,N_26474);
and U28348 (N_28348,N_27221,N_26774);
nand U28349 (N_28349,N_26579,N_27008);
nand U28350 (N_28350,N_26612,N_27585);
or U28351 (N_28351,N_26405,N_26443);
xor U28352 (N_28352,N_27133,N_26966);
nand U28353 (N_28353,N_26825,N_26416);
or U28354 (N_28354,N_27492,N_26586);
nand U28355 (N_28355,N_26702,N_26950);
or U28356 (N_28356,N_27225,N_26964);
or U28357 (N_28357,N_26947,N_27388);
xor U28358 (N_28358,N_26536,N_27115);
or U28359 (N_28359,N_26919,N_26892);
or U28360 (N_28360,N_27144,N_26843);
and U28361 (N_28361,N_27458,N_27101);
nor U28362 (N_28362,N_27434,N_27520);
or U28363 (N_28363,N_27267,N_26932);
nor U28364 (N_28364,N_26702,N_26687);
or U28365 (N_28365,N_26547,N_26831);
xor U28366 (N_28366,N_26938,N_26678);
or U28367 (N_28367,N_27377,N_27182);
nor U28368 (N_28368,N_27535,N_26854);
or U28369 (N_28369,N_27014,N_26883);
xor U28370 (N_28370,N_26950,N_27245);
and U28371 (N_28371,N_26794,N_27342);
and U28372 (N_28372,N_27268,N_26722);
nand U28373 (N_28373,N_27531,N_27325);
nor U28374 (N_28374,N_26924,N_27004);
nor U28375 (N_28375,N_27135,N_26557);
nand U28376 (N_28376,N_27528,N_26750);
nand U28377 (N_28377,N_27390,N_26531);
nand U28378 (N_28378,N_27119,N_27085);
and U28379 (N_28379,N_27117,N_27124);
nand U28380 (N_28380,N_27293,N_27258);
or U28381 (N_28381,N_27553,N_26520);
nor U28382 (N_28382,N_26949,N_26817);
nand U28383 (N_28383,N_27175,N_26975);
or U28384 (N_28384,N_27087,N_26902);
xor U28385 (N_28385,N_26650,N_26522);
nor U28386 (N_28386,N_26641,N_26774);
and U28387 (N_28387,N_27411,N_27117);
or U28388 (N_28388,N_26611,N_26834);
or U28389 (N_28389,N_27154,N_27595);
and U28390 (N_28390,N_26556,N_27287);
nand U28391 (N_28391,N_27276,N_26787);
or U28392 (N_28392,N_27436,N_27153);
xor U28393 (N_28393,N_26908,N_26478);
xnor U28394 (N_28394,N_26995,N_26775);
and U28395 (N_28395,N_26450,N_26428);
xnor U28396 (N_28396,N_27251,N_27418);
and U28397 (N_28397,N_27130,N_26652);
xor U28398 (N_28398,N_27405,N_27532);
and U28399 (N_28399,N_26705,N_27134);
or U28400 (N_28400,N_27099,N_26413);
and U28401 (N_28401,N_26533,N_26907);
xnor U28402 (N_28402,N_27182,N_26513);
and U28403 (N_28403,N_27114,N_26633);
and U28404 (N_28404,N_26453,N_27129);
nor U28405 (N_28405,N_26451,N_27291);
xnor U28406 (N_28406,N_26599,N_27324);
xor U28407 (N_28407,N_27063,N_27485);
xnor U28408 (N_28408,N_26683,N_27057);
xnor U28409 (N_28409,N_27171,N_27021);
xnor U28410 (N_28410,N_26535,N_27243);
nand U28411 (N_28411,N_26778,N_26907);
xor U28412 (N_28412,N_26418,N_26735);
xnor U28413 (N_28413,N_27471,N_27419);
or U28414 (N_28414,N_26780,N_26619);
or U28415 (N_28415,N_27283,N_26801);
or U28416 (N_28416,N_26427,N_26594);
nand U28417 (N_28417,N_26540,N_26704);
or U28418 (N_28418,N_26557,N_26653);
nor U28419 (N_28419,N_26874,N_26763);
nand U28420 (N_28420,N_27241,N_26890);
nand U28421 (N_28421,N_27187,N_27288);
nand U28422 (N_28422,N_26725,N_27199);
and U28423 (N_28423,N_26647,N_26744);
xor U28424 (N_28424,N_27046,N_27171);
xor U28425 (N_28425,N_27133,N_27253);
or U28426 (N_28426,N_26685,N_27069);
and U28427 (N_28427,N_27259,N_27462);
and U28428 (N_28428,N_27226,N_26648);
nand U28429 (N_28429,N_26777,N_26663);
and U28430 (N_28430,N_27550,N_27227);
or U28431 (N_28431,N_26774,N_26741);
and U28432 (N_28432,N_26545,N_26948);
xnor U28433 (N_28433,N_27414,N_26446);
xnor U28434 (N_28434,N_27270,N_26444);
nor U28435 (N_28435,N_27181,N_26720);
nand U28436 (N_28436,N_26648,N_27243);
xor U28437 (N_28437,N_26419,N_26440);
xnor U28438 (N_28438,N_27356,N_26657);
nand U28439 (N_28439,N_27432,N_26761);
xor U28440 (N_28440,N_26834,N_27476);
and U28441 (N_28441,N_27466,N_26676);
and U28442 (N_28442,N_27435,N_27013);
and U28443 (N_28443,N_26491,N_26444);
nor U28444 (N_28444,N_26914,N_26752);
and U28445 (N_28445,N_27082,N_27106);
xor U28446 (N_28446,N_26422,N_27382);
nor U28447 (N_28447,N_26647,N_26823);
nand U28448 (N_28448,N_27385,N_26710);
nand U28449 (N_28449,N_27352,N_27413);
xnor U28450 (N_28450,N_27348,N_26437);
or U28451 (N_28451,N_26943,N_27471);
and U28452 (N_28452,N_26765,N_27167);
and U28453 (N_28453,N_27489,N_26496);
xnor U28454 (N_28454,N_26872,N_27352);
nand U28455 (N_28455,N_27300,N_27312);
or U28456 (N_28456,N_27542,N_27307);
nor U28457 (N_28457,N_27452,N_27302);
nand U28458 (N_28458,N_27252,N_27558);
xor U28459 (N_28459,N_27420,N_27255);
and U28460 (N_28460,N_27437,N_27166);
and U28461 (N_28461,N_27498,N_26577);
nor U28462 (N_28462,N_26917,N_26629);
nand U28463 (N_28463,N_27559,N_27335);
or U28464 (N_28464,N_27566,N_26883);
nor U28465 (N_28465,N_27520,N_27397);
and U28466 (N_28466,N_26990,N_26594);
xnor U28467 (N_28467,N_26639,N_26594);
xnor U28468 (N_28468,N_27096,N_26668);
xor U28469 (N_28469,N_27288,N_26761);
nand U28470 (N_28470,N_27460,N_26927);
and U28471 (N_28471,N_26827,N_27512);
nand U28472 (N_28472,N_27127,N_26765);
and U28473 (N_28473,N_27424,N_27284);
xor U28474 (N_28474,N_27045,N_27260);
xnor U28475 (N_28475,N_27100,N_26985);
xnor U28476 (N_28476,N_27436,N_26585);
xor U28477 (N_28477,N_27586,N_27098);
or U28478 (N_28478,N_26457,N_27437);
and U28479 (N_28479,N_27545,N_27169);
xor U28480 (N_28480,N_26664,N_26565);
nand U28481 (N_28481,N_26712,N_26857);
or U28482 (N_28482,N_26903,N_26602);
and U28483 (N_28483,N_27282,N_27196);
xnor U28484 (N_28484,N_26970,N_26521);
and U28485 (N_28485,N_26910,N_26833);
nor U28486 (N_28486,N_26801,N_27409);
and U28487 (N_28487,N_27437,N_27572);
or U28488 (N_28488,N_27249,N_27423);
xnor U28489 (N_28489,N_27106,N_26523);
xnor U28490 (N_28490,N_27569,N_27147);
or U28491 (N_28491,N_26831,N_27063);
or U28492 (N_28492,N_27184,N_26561);
or U28493 (N_28493,N_27149,N_26997);
and U28494 (N_28494,N_26481,N_26534);
xor U28495 (N_28495,N_27469,N_27366);
nand U28496 (N_28496,N_26533,N_26701);
nand U28497 (N_28497,N_27569,N_27376);
nor U28498 (N_28498,N_27035,N_27573);
nand U28499 (N_28499,N_26446,N_27367);
nand U28500 (N_28500,N_27388,N_26564);
and U28501 (N_28501,N_26637,N_26715);
nand U28502 (N_28502,N_26757,N_26937);
xnor U28503 (N_28503,N_27012,N_27096);
or U28504 (N_28504,N_26567,N_27447);
nand U28505 (N_28505,N_27491,N_27347);
or U28506 (N_28506,N_27029,N_26551);
nand U28507 (N_28507,N_27024,N_27193);
nand U28508 (N_28508,N_26880,N_26539);
nor U28509 (N_28509,N_26718,N_26944);
and U28510 (N_28510,N_27081,N_26517);
nor U28511 (N_28511,N_26506,N_27053);
nand U28512 (N_28512,N_26662,N_26611);
and U28513 (N_28513,N_26932,N_27072);
nand U28514 (N_28514,N_27226,N_27248);
nand U28515 (N_28515,N_26689,N_27519);
and U28516 (N_28516,N_26650,N_26941);
xnor U28517 (N_28517,N_26910,N_26440);
nor U28518 (N_28518,N_27338,N_26694);
or U28519 (N_28519,N_26521,N_27185);
xnor U28520 (N_28520,N_26893,N_26597);
xnor U28521 (N_28521,N_27235,N_27085);
xnor U28522 (N_28522,N_27449,N_27088);
and U28523 (N_28523,N_26785,N_26796);
or U28524 (N_28524,N_26993,N_26556);
and U28525 (N_28525,N_26699,N_27364);
nor U28526 (N_28526,N_27469,N_26825);
xnor U28527 (N_28527,N_27540,N_27356);
and U28528 (N_28528,N_27317,N_26592);
nor U28529 (N_28529,N_27135,N_27216);
or U28530 (N_28530,N_26750,N_26730);
and U28531 (N_28531,N_27041,N_26610);
xor U28532 (N_28532,N_27180,N_26488);
xor U28533 (N_28533,N_27140,N_27036);
xnor U28534 (N_28534,N_26920,N_27023);
nor U28535 (N_28535,N_26929,N_27259);
and U28536 (N_28536,N_27174,N_27035);
or U28537 (N_28537,N_27084,N_26934);
xor U28538 (N_28538,N_26863,N_27128);
nor U28539 (N_28539,N_26603,N_26670);
xnor U28540 (N_28540,N_26997,N_26786);
and U28541 (N_28541,N_26617,N_26683);
nor U28542 (N_28542,N_27551,N_26491);
nand U28543 (N_28543,N_26891,N_26467);
nor U28544 (N_28544,N_27318,N_26635);
or U28545 (N_28545,N_27082,N_27414);
xnor U28546 (N_28546,N_26744,N_26616);
xor U28547 (N_28547,N_26919,N_27586);
nor U28548 (N_28548,N_26530,N_26628);
nor U28549 (N_28549,N_26699,N_27295);
xnor U28550 (N_28550,N_27138,N_26733);
nor U28551 (N_28551,N_27452,N_27569);
nor U28552 (N_28552,N_26768,N_26977);
xnor U28553 (N_28553,N_26684,N_27542);
nor U28554 (N_28554,N_26524,N_27152);
nand U28555 (N_28555,N_26603,N_27136);
nor U28556 (N_28556,N_26981,N_27475);
or U28557 (N_28557,N_26943,N_26989);
nand U28558 (N_28558,N_27347,N_26577);
and U28559 (N_28559,N_26956,N_26684);
nand U28560 (N_28560,N_27266,N_26685);
nand U28561 (N_28561,N_26786,N_26989);
nor U28562 (N_28562,N_26669,N_26698);
or U28563 (N_28563,N_26824,N_27184);
nor U28564 (N_28564,N_26988,N_26738);
and U28565 (N_28565,N_26577,N_27553);
nand U28566 (N_28566,N_27014,N_27287);
nand U28567 (N_28567,N_26898,N_27191);
nor U28568 (N_28568,N_27097,N_26434);
xnor U28569 (N_28569,N_26503,N_26582);
and U28570 (N_28570,N_27035,N_26730);
and U28571 (N_28571,N_27497,N_26865);
or U28572 (N_28572,N_26949,N_27150);
nor U28573 (N_28573,N_27292,N_26659);
xnor U28574 (N_28574,N_26817,N_26954);
xnor U28575 (N_28575,N_26993,N_26877);
or U28576 (N_28576,N_27001,N_27477);
xnor U28577 (N_28577,N_26599,N_26502);
xnor U28578 (N_28578,N_27149,N_26571);
xor U28579 (N_28579,N_26840,N_27073);
xor U28580 (N_28580,N_27354,N_26795);
xor U28581 (N_28581,N_26766,N_26860);
nand U28582 (N_28582,N_26984,N_27311);
and U28583 (N_28583,N_27409,N_27075);
xnor U28584 (N_28584,N_27119,N_26474);
and U28585 (N_28585,N_27508,N_26922);
nand U28586 (N_28586,N_27557,N_26698);
xnor U28587 (N_28587,N_27293,N_27150);
nand U28588 (N_28588,N_26679,N_27544);
xnor U28589 (N_28589,N_26829,N_27374);
nor U28590 (N_28590,N_26841,N_26410);
and U28591 (N_28591,N_27376,N_27460);
or U28592 (N_28592,N_26526,N_27430);
xor U28593 (N_28593,N_27567,N_26829);
xnor U28594 (N_28594,N_27396,N_27580);
nand U28595 (N_28595,N_27255,N_26446);
nor U28596 (N_28596,N_26728,N_26783);
or U28597 (N_28597,N_27178,N_27428);
or U28598 (N_28598,N_27083,N_26765);
and U28599 (N_28599,N_27127,N_27038);
xnor U28600 (N_28600,N_26922,N_27163);
nor U28601 (N_28601,N_26864,N_26849);
xnor U28602 (N_28602,N_27052,N_27481);
and U28603 (N_28603,N_27213,N_26558);
and U28604 (N_28604,N_27309,N_27444);
nor U28605 (N_28605,N_27146,N_26667);
xor U28606 (N_28606,N_27006,N_26756);
nand U28607 (N_28607,N_26934,N_27295);
xor U28608 (N_28608,N_26509,N_27398);
xor U28609 (N_28609,N_27426,N_27360);
nor U28610 (N_28610,N_26559,N_26822);
or U28611 (N_28611,N_27307,N_26954);
or U28612 (N_28612,N_26477,N_27304);
and U28613 (N_28613,N_27241,N_26416);
and U28614 (N_28614,N_26659,N_26761);
nor U28615 (N_28615,N_27427,N_26975);
or U28616 (N_28616,N_26782,N_26414);
xor U28617 (N_28617,N_27054,N_26485);
and U28618 (N_28618,N_27002,N_26609);
and U28619 (N_28619,N_27205,N_27139);
nor U28620 (N_28620,N_27101,N_26895);
or U28621 (N_28621,N_26458,N_26783);
nand U28622 (N_28622,N_27048,N_27032);
xor U28623 (N_28623,N_27365,N_26957);
or U28624 (N_28624,N_27317,N_26452);
and U28625 (N_28625,N_26435,N_26997);
nor U28626 (N_28626,N_27452,N_27024);
nand U28627 (N_28627,N_27290,N_27064);
nand U28628 (N_28628,N_27554,N_27192);
nor U28629 (N_28629,N_26502,N_26415);
and U28630 (N_28630,N_26792,N_26996);
nand U28631 (N_28631,N_27392,N_27449);
and U28632 (N_28632,N_26650,N_27570);
nand U28633 (N_28633,N_27384,N_27344);
nand U28634 (N_28634,N_27229,N_27456);
nor U28635 (N_28635,N_26606,N_27429);
xnor U28636 (N_28636,N_27558,N_27412);
nand U28637 (N_28637,N_26896,N_26737);
xor U28638 (N_28638,N_27043,N_26484);
and U28639 (N_28639,N_26524,N_27046);
and U28640 (N_28640,N_26938,N_27125);
xnor U28641 (N_28641,N_26914,N_27143);
nand U28642 (N_28642,N_26985,N_27274);
xor U28643 (N_28643,N_27027,N_26518);
nor U28644 (N_28644,N_26885,N_27534);
nor U28645 (N_28645,N_27125,N_27230);
nor U28646 (N_28646,N_26486,N_26895);
nor U28647 (N_28647,N_27312,N_26531);
nor U28648 (N_28648,N_26903,N_27266);
xnor U28649 (N_28649,N_26748,N_26403);
nand U28650 (N_28650,N_26708,N_27214);
nor U28651 (N_28651,N_27203,N_26861);
nand U28652 (N_28652,N_27523,N_27017);
nor U28653 (N_28653,N_27197,N_27474);
nand U28654 (N_28654,N_26540,N_27062);
and U28655 (N_28655,N_27514,N_27343);
or U28656 (N_28656,N_26692,N_27528);
nor U28657 (N_28657,N_27352,N_27120);
nand U28658 (N_28658,N_27231,N_27457);
nand U28659 (N_28659,N_26618,N_27210);
and U28660 (N_28660,N_27371,N_27414);
xnor U28661 (N_28661,N_26854,N_27461);
nor U28662 (N_28662,N_26859,N_27427);
nor U28663 (N_28663,N_27189,N_26585);
or U28664 (N_28664,N_26881,N_27317);
nor U28665 (N_28665,N_26560,N_26533);
xnor U28666 (N_28666,N_26508,N_26744);
nand U28667 (N_28667,N_27458,N_26686);
xnor U28668 (N_28668,N_26552,N_27166);
or U28669 (N_28669,N_26965,N_27365);
or U28670 (N_28670,N_26686,N_27468);
xor U28671 (N_28671,N_26626,N_26789);
xor U28672 (N_28672,N_27327,N_26536);
nor U28673 (N_28673,N_26938,N_27582);
nand U28674 (N_28674,N_26763,N_26487);
and U28675 (N_28675,N_27431,N_26776);
nand U28676 (N_28676,N_26854,N_26719);
xnor U28677 (N_28677,N_27176,N_27510);
nand U28678 (N_28678,N_26636,N_26562);
and U28679 (N_28679,N_27246,N_27212);
or U28680 (N_28680,N_26416,N_27268);
nand U28681 (N_28681,N_26947,N_26420);
nand U28682 (N_28682,N_26691,N_26788);
and U28683 (N_28683,N_26737,N_26719);
and U28684 (N_28684,N_27128,N_26588);
nand U28685 (N_28685,N_27130,N_27593);
and U28686 (N_28686,N_27386,N_26507);
nand U28687 (N_28687,N_26793,N_26427);
nor U28688 (N_28688,N_26573,N_26925);
xnor U28689 (N_28689,N_27115,N_27249);
nand U28690 (N_28690,N_26848,N_26618);
nand U28691 (N_28691,N_27552,N_26621);
nor U28692 (N_28692,N_26877,N_26986);
and U28693 (N_28693,N_27293,N_26695);
or U28694 (N_28694,N_27307,N_27048);
nor U28695 (N_28695,N_26775,N_26904);
xnor U28696 (N_28696,N_26501,N_26595);
nor U28697 (N_28697,N_27030,N_26978);
and U28698 (N_28698,N_26766,N_27232);
or U28699 (N_28699,N_27062,N_27488);
nor U28700 (N_28700,N_27000,N_27409);
nand U28701 (N_28701,N_27065,N_27004);
nor U28702 (N_28702,N_27253,N_27231);
and U28703 (N_28703,N_27273,N_26841);
xor U28704 (N_28704,N_26477,N_26561);
nor U28705 (N_28705,N_26760,N_27513);
nand U28706 (N_28706,N_27323,N_27222);
or U28707 (N_28707,N_26512,N_27220);
or U28708 (N_28708,N_27241,N_26904);
nor U28709 (N_28709,N_26667,N_26513);
nor U28710 (N_28710,N_27094,N_26632);
xnor U28711 (N_28711,N_27092,N_26732);
or U28712 (N_28712,N_27099,N_27503);
nor U28713 (N_28713,N_26998,N_27374);
nand U28714 (N_28714,N_27568,N_26405);
and U28715 (N_28715,N_27079,N_26588);
nand U28716 (N_28716,N_27077,N_26603);
and U28717 (N_28717,N_27127,N_27005);
xor U28718 (N_28718,N_27234,N_26994);
xor U28719 (N_28719,N_27434,N_26419);
and U28720 (N_28720,N_27016,N_27036);
nor U28721 (N_28721,N_27126,N_26569);
nor U28722 (N_28722,N_26748,N_26406);
nor U28723 (N_28723,N_26505,N_26953);
xor U28724 (N_28724,N_27488,N_27376);
and U28725 (N_28725,N_26705,N_27366);
nand U28726 (N_28726,N_27537,N_26591);
nor U28727 (N_28727,N_26943,N_27525);
or U28728 (N_28728,N_27487,N_26821);
or U28729 (N_28729,N_27081,N_27481);
nor U28730 (N_28730,N_26441,N_26950);
or U28731 (N_28731,N_26960,N_26666);
xor U28732 (N_28732,N_27361,N_26624);
and U28733 (N_28733,N_26798,N_27246);
or U28734 (N_28734,N_26921,N_27052);
nor U28735 (N_28735,N_27141,N_27215);
and U28736 (N_28736,N_27481,N_26739);
nor U28737 (N_28737,N_27587,N_26657);
nor U28738 (N_28738,N_26457,N_27115);
or U28739 (N_28739,N_27006,N_26766);
nand U28740 (N_28740,N_26601,N_26699);
nand U28741 (N_28741,N_26866,N_27104);
nand U28742 (N_28742,N_27060,N_27489);
and U28743 (N_28743,N_27163,N_27331);
and U28744 (N_28744,N_27511,N_26893);
or U28745 (N_28745,N_27224,N_26930);
xnor U28746 (N_28746,N_26638,N_26929);
and U28747 (N_28747,N_26938,N_27370);
or U28748 (N_28748,N_27089,N_27238);
or U28749 (N_28749,N_27159,N_26534);
xor U28750 (N_28750,N_26600,N_26528);
nor U28751 (N_28751,N_27150,N_26482);
nand U28752 (N_28752,N_26549,N_26646);
or U28753 (N_28753,N_27024,N_26754);
xor U28754 (N_28754,N_27530,N_26503);
or U28755 (N_28755,N_26989,N_27539);
xnor U28756 (N_28756,N_26719,N_26736);
or U28757 (N_28757,N_26677,N_27469);
xor U28758 (N_28758,N_26461,N_27304);
and U28759 (N_28759,N_27231,N_27293);
and U28760 (N_28760,N_26479,N_27506);
and U28761 (N_28761,N_26708,N_27336);
xnor U28762 (N_28762,N_27500,N_27174);
nand U28763 (N_28763,N_26468,N_27511);
or U28764 (N_28764,N_26977,N_27209);
and U28765 (N_28765,N_26860,N_26582);
xor U28766 (N_28766,N_26816,N_26451);
nand U28767 (N_28767,N_26803,N_27521);
and U28768 (N_28768,N_26997,N_27042);
nand U28769 (N_28769,N_27264,N_26563);
xnor U28770 (N_28770,N_26996,N_27017);
nor U28771 (N_28771,N_26431,N_27425);
and U28772 (N_28772,N_27344,N_27466);
xnor U28773 (N_28773,N_27244,N_27116);
nor U28774 (N_28774,N_27408,N_27157);
xor U28775 (N_28775,N_27255,N_26721);
nor U28776 (N_28776,N_27343,N_27353);
or U28777 (N_28777,N_26506,N_26417);
nor U28778 (N_28778,N_26544,N_27221);
nand U28779 (N_28779,N_27034,N_27195);
nor U28780 (N_28780,N_26894,N_26881);
and U28781 (N_28781,N_27183,N_26977);
nor U28782 (N_28782,N_26691,N_26480);
xor U28783 (N_28783,N_26889,N_26813);
and U28784 (N_28784,N_26802,N_27329);
xor U28785 (N_28785,N_27134,N_26558);
xor U28786 (N_28786,N_27296,N_26733);
nand U28787 (N_28787,N_27258,N_27537);
nor U28788 (N_28788,N_26459,N_26868);
xnor U28789 (N_28789,N_27489,N_26813);
or U28790 (N_28790,N_26471,N_26924);
xor U28791 (N_28791,N_27083,N_26786);
xnor U28792 (N_28792,N_27064,N_26594);
nor U28793 (N_28793,N_26637,N_27105);
and U28794 (N_28794,N_26596,N_27160);
and U28795 (N_28795,N_26708,N_26952);
or U28796 (N_28796,N_26446,N_26873);
and U28797 (N_28797,N_27226,N_27384);
and U28798 (N_28798,N_26963,N_27512);
nor U28799 (N_28799,N_26416,N_26449);
xnor U28800 (N_28800,N_28646,N_28330);
or U28801 (N_28801,N_28064,N_28675);
and U28802 (N_28802,N_27901,N_28732);
nand U28803 (N_28803,N_27922,N_28766);
and U28804 (N_28804,N_28385,N_27786);
nor U28805 (N_28805,N_28116,N_27731);
xnor U28806 (N_28806,N_28166,N_27938);
nand U28807 (N_28807,N_27788,N_28018);
or U28808 (N_28808,N_28053,N_28102);
nand U28809 (N_28809,N_28659,N_28419);
or U28810 (N_28810,N_28208,N_27750);
or U28811 (N_28811,N_28325,N_28606);
or U28812 (N_28812,N_28788,N_27666);
nand U28813 (N_28813,N_27821,N_28504);
xnor U28814 (N_28814,N_28148,N_28192);
xnor U28815 (N_28815,N_27815,N_27622);
xor U28816 (N_28816,N_27921,N_28787);
xor U28817 (N_28817,N_27974,N_28292);
or U28818 (N_28818,N_28439,N_28351);
xnor U28819 (N_28819,N_27771,N_28026);
xor U28820 (N_28820,N_28489,N_28366);
nor U28821 (N_28821,N_27682,N_27784);
and U28822 (N_28822,N_28099,N_28476);
nor U28823 (N_28823,N_27691,N_28238);
xor U28824 (N_28824,N_28127,N_27793);
or U28825 (N_28825,N_27842,N_28161);
xnor U28826 (N_28826,N_27669,N_28651);
xnor U28827 (N_28827,N_28394,N_27678);
and U28828 (N_28828,N_27768,N_28700);
xor U28829 (N_28829,N_28584,N_28591);
nand U28830 (N_28830,N_28557,N_28478);
and U28831 (N_28831,N_28631,N_28400);
or U28832 (N_28832,N_28185,N_28249);
or U28833 (N_28833,N_28550,N_28129);
xor U28834 (N_28834,N_28364,N_27916);
xnor U28835 (N_28835,N_28746,N_27765);
or U28836 (N_28836,N_27713,N_28067);
or U28837 (N_28837,N_27726,N_27871);
or U28838 (N_28838,N_28272,N_28620);
nand U28839 (N_28839,N_28341,N_28475);
nand U28840 (N_28840,N_27639,N_27830);
or U28841 (N_28841,N_28072,N_28637);
or U28842 (N_28842,N_28309,N_27658);
xor U28843 (N_28843,N_27787,N_28375);
or U28844 (N_28844,N_27603,N_27987);
and U28845 (N_28845,N_28623,N_28568);
or U28846 (N_28846,N_27655,N_27849);
nand U28847 (N_28847,N_28462,N_27873);
nand U28848 (N_28848,N_28164,N_28432);
xor U28849 (N_28849,N_28368,N_28149);
nor U28850 (N_28850,N_27758,N_28514);
nand U28851 (N_28851,N_28434,N_27613);
or U28852 (N_28852,N_27948,N_28312);
xor U28853 (N_28853,N_27918,N_27944);
nand U28854 (N_28854,N_28370,N_28662);
nor U28855 (N_28855,N_28636,N_27915);
nand U28856 (N_28856,N_28595,N_28590);
or U28857 (N_28857,N_27970,N_28046);
and U28858 (N_28858,N_28305,N_27611);
or U28859 (N_28859,N_27646,N_27863);
nand U28860 (N_28860,N_27879,N_27618);
or U28861 (N_28861,N_28730,N_27664);
nor U28862 (N_28862,N_28790,N_27614);
and U28863 (N_28863,N_28290,N_28331);
nand U28864 (N_28864,N_28182,N_27656);
xnor U28865 (N_28865,N_27814,N_28545);
or U28866 (N_28866,N_28034,N_27952);
or U28867 (N_28867,N_28795,N_28177);
nand U28868 (N_28868,N_27660,N_28684);
and U28869 (N_28869,N_28772,N_28665);
and U28870 (N_28870,N_27962,N_27757);
or U28871 (N_28871,N_28578,N_28227);
or U28872 (N_28872,N_28598,N_28791);
nor U28873 (N_28873,N_28390,N_27616);
or U28874 (N_28874,N_28650,N_27817);
nand U28875 (N_28875,N_27882,N_27960);
or U28876 (N_28876,N_28518,N_27846);
xor U28877 (N_28877,N_28410,N_28525);
nor U28878 (N_28878,N_27967,N_27973);
nand U28879 (N_28879,N_28090,N_27700);
nand U28880 (N_28880,N_28200,N_28387);
or U28881 (N_28881,N_28126,N_27902);
xor U28882 (N_28882,N_27790,N_28193);
or U28883 (N_28883,N_27626,N_28115);
xnor U28884 (N_28884,N_28245,N_28376);
nand U28885 (N_28885,N_28444,N_28445);
nand U28886 (N_28886,N_28477,N_28248);
or U28887 (N_28887,N_27752,N_28757);
or U28888 (N_28888,N_27883,N_27694);
and U28889 (N_28889,N_27612,N_28269);
xor U28890 (N_28890,N_28288,N_27601);
and U28891 (N_28891,N_28332,N_28609);
xor U28892 (N_28892,N_27703,N_28002);
xnor U28893 (N_28893,N_28567,N_27699);
nor U28894 (N_28894,N_28213,N_27940);
or U28895 (N_28895,N_28028,N_28397);
or U28896 (N_28896,N_27839,N_27898);
nand U28897 (N_28897,N_28508,N_27670);
nand U28898 (N_28898,N_28784,N_28315);
nor U28899 (N_28899,N_27744,N_27761);
and U28900 (N_28900,N_28393,N_28635);
and U28901 (N_28901,N_28740,N_28306);
or U28902 (N_28902,N_28079,N_28284);
nor U28903 (N_28903,N_28076,N_28451);
and U28904 (N_28904,N_27980,N_27982);
xnor U28905 (N_28905,N_27759,N_27939);
and U28906 (N_28906,N_28293,N_28660);
xor U28907 (N_28907,N_28159,N_27629);
xnor U28908 (N_28908,N_28179,N_27766);
nor U28909 (N_28909,N_28274,N_28664);
nand U28910 (N_28910,N_28524,N_28541);
nand U28911 (N_28911,N_27826,N_28174);
or U28912 (N_28912,N_27755,N_28198);
or U28913 (N_28913,N_28041,N_28285);
nor U28914 (N_28914,N_27977,N_28407);
xnor U28915 (N_28915,N_28307,N_28367);
nor U28916 (N_28916,N_28782,N_27868);
and U28917 (N_28917,N_28141,N_27850);
nand U28918 (N_28918,N_28236,N_28059);
nand U28919 (N_28919,N_28256,N_27874);
nand U28920 (N_28920,N_27679,N_28764);
nor U28921 (N_28921,N_28362,N_28629);
or U28922 (N_28922,N_27742,N_27932);
nor U28923 (N_28923,N_28391,N_28701);
and U28924 (N_28924,N_27647,N_27609);
nor U28925 (N_28925,N_27734,N_28075);
and U28926 (N_28926,N_27870,N_28011);
nand U28927 (N_28927,N_28570,N_28589);
nor U28928 (N_28928,N_27667,N_28638);
nor U28929 (N_28929,N_27966,N_27866);
or U28930 (N_28930,N_27756,N_28258);
nor U28931 (N_28931,N_27896,N_28142);
xnor U28932 (N_28932,N_28277,N_28374);
or U28933 (N_28933,N_27828,N_28729);
or U28934 (N_28934,N_28178,N_28043);
nor U28935 (N_28935,N_28054,N_28440);
or U28936 (N_28936,N_28280,N_27968);
xnor U28937 (N_28937,N_27843,N_28247);
or U28938 (N_28938,N_28540,N_27941);
nor U28939 (N_28939,N_28505,N_28798);
xnor U28940 (N_28940,N_28209,N_28077);
and U28941 (N_28941,N_27727,N_28340);
nor U28942 (N_28942,N_27781,N_28671);
and U28943 (N_28943,N_28088,N_28024);
xor U28944 (N_28944,N_28435,N_27858);
xor U28945 (N_28945,N_28255,N_27988);
xnor U28946 (N_28946,N_28719,N_27947);
and U28947 (N_28947,N_27957,N_27897);
or U28948 (N_28948,N_27976,N_28747);
or U28949 (N_28949,N_28260,N_28743);
or U28950 (N_28950,N_27894,N_27906);
nor U28951 (N_28951,N_28345,N_28372);
or U28952 (N_28952,N_28128,N_27762);
nor U28953 (N_28953,N_28217,N_28109);
nand U28954 (N_28954,N_28493,N_27723);
nor U28955 (N_28955,N_28282,N_28682);
nand U28956 (N_28956,N_27773,N_27869);
nor U28957 (N_28957,N_28089,N_27841);
or U28958 (N_28958,N_28082,N_28032);
nor U28959 (N_28959,N_27711,N_28436);
nor U28960 (N_28960,N_28399,N_28555);
xnor U28961 (N_28961,N_28441,N_28634);
nor U28962 (N_28962,N_28071,N_27619);
and U28963 (N_28963,N_28098,N_28287);
and U28964 (N_28964,N_28744,N_27692);
or U28965 (N_28965,N_28145,N_28420);
nand U28966 (N_28966,N_28537,N_28443);
xor U28967 (N_28967,N_28106,N_28146);
nand U28968 (N_28968,N_28551,N_28723);
nor U28969 (N_28969,N_28749,N_28528);
or U28970 (N_28970,N_28699,N_28031);
and U28971 (N_28971,N_28498,N_28728);
and U28972 (N_28972,N_28733,N_28379);
nand U28973 (N_28973,N_28753,N_28383);
and U28974 (N_28974,N_28409,N_28482);
nor U28975 (N_28975,N_28668,N_27854);
nor U28976 (N_28976,N_28311,N_28742);
xor U28977 (N_28977,N_27684,N_28377);
nand U28978 (N_28978,N_27764,N_28454);
nor U28979 (N_28979,N_27736,N_28333);
or U28980 (N_28980,N_28632,N_28422);
nor U28981 (N_28981,N_28763,N_28074);
or U28982 (N_28982,N_28020,N_28676);
xor U28983 (N_28983,N_28052,N_28512);
nor U28984 (N_28984,N_27845,N_27714);
and U28985 (N_28985,N_27641,N_28007);
or U28986 (N_28986,N_28327,N_28658);
xnor U28987 (N_28987,N_28471,N_28726);
or U28988 (N_28988,N_27607,N_28424);
and U28989 (N_28989,N_27783,N_28428);
or U28990 (N_28990,N_28736,N_27633);
or U28991 (N_28991,N_27949,N_28796);
nand U28992 (N_28992,N_28547,N_27649);
xor U28993 (N_28993,N_28770,N_28196);
nor U28994 (N_28994,N_28479,N_28014);
nor U28995 (N_28995,N_28497,N_28158);
and U28996 (N_28996,N_27877,N_27677);
xnor U28997 (N_28997,N_27665,N_28692);
xnor U28998 (N_28998,N_27753,N_28470);
xnor U28999 (N_28999,N_27958,N_27777);
nor U29000 (N_29000,N_27946,N_27965);
or U29001 (N_29001,N_28343,N_28016);
or U29002 (N_29002,N_27867,N_27640);
nand U29003 (N_29003,N_27981,N_28688);
xnor U29004 (N_29004,N_28310,N_28322);
nor U29005 (N_29005,N_27803,N_28473);
nand U29006 (N_29006,N_27943,N_28681);
or U29007 (N_29007,N_27878,N_28097);
or U29008 (N_29008,N_27747,N_28040);
and U29009 (N_29009,N_28725,N_28360);
xnor U29010 (N_29010,N_27994,N_27698);
or U29011 (N_29011,N_28622,N_28502);
and U29012 (N_29012,N_28022,N_27820);
xnor U29013 (N_29013,N_28296,N_28495);
nor U29014 (N_29014,N_28147,N_28600);
nor U29015 (N_29015,N_28122,N_27709);
nand U29016 (N_29016,N_28205,N_27913);
xnor U29017 (N_29017,N_28013,N_27637);
nor U29018 (N_29018,N_28242,N_28101);
xnor U29019 (N_29019,N_27903,N_28438);
and U29020 (N_29020,N_28610,N_28318);
nor U29021 (N_29021,N_27978,N_28580);
and U29022 (N_29022,N_27673,N_28170);
xor U29023 (N_29023,N_27663,N_28500);
nor U29024 (N_29024,N_27717,N_28063);
nand U29025 (N_29025,N_28469,N_28133);
xnor U29026 (N_29026,N_28652,N_28369);
and U29027 (N_29027,N_27721,N_27780);
nand U29028 (N_29028,N_27975,N_28546);
and U29029 (N_29029,N_28000,N_27865);
and U29030 (N_29030,N_28472,N_28095);
nor U29031 (N_29031,N_27862,N_28211);
nor U29032 (N_29032,N_28587,N_28281);
nor U29033 (N_29033,N_28301,N_27991);
and U29034 (N_29034,N_28283,N_27895);
xnor U29035 (N_29035,N_28207,N_28056);
and U29036 (N_29036,N_28669,N_27620);
nor U29037 (N_29037,N_27886,N_28357);
xor U29038 (N_29038,N_27890,N_27838);
or U29039 (N_29039,N_28427,N_28769);
or U29040 (N_29040,N_28153,N_28690);
nand U29041 (N_29041,N_28503,N_27628);
xnor U29042 (N_29042,N_28299,N_28703);
or U29043 (N_29043,N_27652,N_28481);
or U29044 (N_29044,N_28752,N_27674);
nor U29045 (N_29045,N_28065,N_27995);
or U29046 (N_29046,N_28751,N_28253);
and U29047 (N_29047,N_28674,N_27724);
or U29048 (N_29048,N_28694,N_28237);
nor U29049 (N_29049,N_28756,N_28492);
xnor U29050 (N_29050,N_28416,N_27625);
nand U29051 (N_29051,N_28015,N_28354);
and U29052 (N_29052,N_28349,N_27951);
xnor U29053 (N_29053,N_28317,N_28405);
or U29054 (N_29054,N_28696,N_28779);
nor U29055 (N_29055,N_27608,N_28686);
nor U29056 (N_29056,N_27855,N_28533);
or U29057 (N_29057,N_28566,N_28244);
and U29058 (N_29058,N_27707,N_27754);
or U29059 (N_29059,N_27937,N_28712);
and U29060 (N_29060,N_28175,N_28713);
or U29061 (N_29061,N_27778,N_28176);
nor U29062 (N_29062,N_27831,N_28654);
nand U29063 (N_29063,N_28768,N_27840);
and U29064 (N_29064,N_27800,N_28656);
and U29065 (N_29065,N_28113,N_28395);
nor U29066 (N_29066,N_28335,N_28507);
or U29067 (N_29067,N_28216,N_27893);
nor U29068 (N_29068,N_27688,N_27719);
xor U29069 (N_29069,N_28794,N_28655);
xor U29070 (N_29070,N_27749,N_27972);
or U29071 (N_29071,N_28775,N_28418);
nand U29072 (N_29072,N_27774,N_28573);
xnor U29073 (N_29073,N_28136,N_28644);
nand U29074 (N_29074,N_28388,N_27885);
and U29075 (N_29075,N_28398,N_28510);
nand U29076 (N_29076,N_27739,N_27805);
or U29077 (N_29077,N_27942,N_27776);
nand U29078 (N_29078,N_28093,N_28214);
xor U29079 (N_29079,N_28496,N_28218);
and U29080 (N_29080,N_28561,N_28488);
or U29081 (N_29081,N_27680,N_28384);
xor U29082 (N_29082,N_28336,N_28544);
xor U29083 (N_29083,N_28588,N_28358);
nor U29084 (N_29084,N_28552,N_28618);
or U29085 (N_29085,N_28104,N_28767);
xor U29086 (N_29086,N_28259,N_27853);
and U29087 (N_29087,N_28371,N_28118);
nand U29088 (N_29088,N_28137,N_27889);
and U29089 (N_29089,N_28163,N_28778);
nor U29090 (N_29090,N_28008,N_27892);
nor U29091 (N_29091,N_28215,N_27745);
or U29092 (N_29092,N_28091,N_28263);
nand U29093 (N_29093,N_28162,N_28268);
and U29094 (N_29094,N_27971,N_27811);
or U29095 (N_29095,N_28267,N_28680);
nand U29096 (N_29096,N_28792,N_28594);
xor U29097 (N_29097,N_28017,N_28107);
xnor U29098 (N_29098,N_27634,N_28585);
nand U29099 (N_29099,N_28643,N_28710);
nor U29100 (N_29100,N_28225,N_28707);
nor U29101 (N_29101,N_28621,N_28604);
or U29102 (N_29102,N_28607,N_27746);
nor U29103 (N_29103,N_28019,N_27763);
or U29104 (N_29104,N_28401,N_27998);
xor U29105 (N_29105,N_27806,N_27775);
nor U29106 (N_29106,N_27685,N_28363);
or U29107 (N_29107,N_28799,N_27624);
xor U29108 (N_29108,N_27675,N_27769);
nand U29109 (N_29109,N_28139,N_28716);
nand U29110 (N_29110,N_28641,N_28734);
or U29111 (N_29111,N_27956,N_28157);
xnor U29112 (N_29112,N_27671,N_28023);
nand U29113 (N_29113,N_28191,N_28037);
nand U29114 (N_29114,N_27911,N_28073);
nor U29115 (N_29115,N_27955,N_28464);
or U29116 (N_29116,N_28184,N_27837);
nor U29117 (N_29117,N_27743,N_28529);
or U29118 (N_29118,N_27600,N_28415);
xnor U29119 (N_29119,N_28199,N_28291);
nor U29120 (N_29120,N_28001,N_28110);
xor U29121 (N_29121,N_28563,N_28152);
and U29122 (N_29122,N_28169,N_28564);
or U29123 (N_29123,N_28261,N_28691);
nand U29124 (N_29124,N_28061,N_27887);
and U29125 (N_29125,N_28144,N_28648);
nor U29126 (N_29126,N_28738,N_27996);
or U29127 (N_29127,N_28316,N_28038);
or U29128 (N_29128,N_27836,N_28273);
xor U29129 (N_29129,N_27930,N_28289);
nand U29130 (N_29130,N_28516,N_28339);
nor U29131 (N_29131,N_28513,N_28134);
or U29132 (N_29132,N_28754,N_28295);
xnor U29133 (N_29133,N_28569,N_28797);
and U29134 (N_29134,N_28762,N_28173);
or U29135 (N_29135,N_28532,N_28069);
xor U29136 (N_29136,N_27728,N_27621);
nand U29137 (N_29137,N_27861,N_28484);
nand U29138 (N_29138,N_28560,N_27804);
and U29139 (N_29139,N_28096,N_28592);
nand U29140 (N_29140,N_28718,N_27884);
xnor U29141 (N_29141,N_27789,N_27760);
nand U29142 (N_29142,N_28086,N_28042);
xor U29143 (N_29143,N_28130,N_27662);
or U29144 (N_29144,N_28735,N_28755);
nor U29145 (N_29145,N_28265,N_28414);
or U29146 (N_29146,N_28765,N_28683);
xnor U29147 (N_29147,N_28499,N_28771);
and U29148 (N_29148,N_27704,N_27710);
nand U29149 (N_29149,N_27876,N_28534);
nor U29150 (N_29150,N_28466,N_27827);
nand U29151 (N_29151,N_28112,N_27857);
nor U29152 (N_29152,N_28527,N_28006);
nand U29153 (N_29153,N_28297,N_28189);
nand U29154 (N_29154,N_28050,N_28353);
and U29155 (N_29155,N_28346,N_27912);
or U29156 (N_29156,N_27693,N_27833);
and U29157 (N_29157,N_27792,N_28204);
xnor U29158 (N_29158,N_27963,N_28012);
xor U29159 (N_29159,N_28522,N_28119);
nor U29160 (N_29160,N_27636,N_28223);
xor U29161 (N_29161,N_28328,N_28761);
or U29162 (N_29162,N_28165,N_27825);
nor U29163 (N_29163,N_28373,N_28143);
xor U29164 (N_29164,N_28549,N_28640);
or U29165 (N_29165,N_27794,N_28461);
nand U29166 (N_29166,N_28760,N_27954);
xor U29167 (N_29167,N_28612,N_28603);
xor U29168 (N_29168,N_28233,N_28188);
or U29169 (N_29169,N_28448,N_28080);
and U29170 (N_29170,N_28647,N_28087);
or U29171 (N_29171,N_28487,N_28672);
xnor U29172 (N_29172,N_27829,N_28490);
xor U29173 (N_29173,N_27610,N_28727);
xor U29174 (N_29174,N_27690,N_28705);
or U29175 (N_29175,N_28168,N_28463);
nand U29176 (N_29176,N_28465,N_27785);
nand U29177 (N_29177,N_28323,N_27986);
and U29178 (N_29178,N_28467,N_28459);
or U29179 (N_29179,N_27999,N_28220);
and U29180 (N_29180,N_27651,N_27899);
or U29181 (N_29181,N_28523,N_28536);
nand U29182 (N_29182,N_28206,N_28412);
and U29183 (N_29183,N_28642,N_28491);
or U29184 (N_29184,N_28085,N_27832);
or U29185 (N_29185,N_28049,N_28679);
nor U29186 (N_29186,N_28628,N_28081);
nand U29187 (N_29187,N_28124,N_28486);
xor U29188 (N_29188,N_28396,N_27659);
xnor U29189 (N_29189,N_27720,N_28447);
xor U29190 (N_29190,N_28449,N_28203);
or U29191 (N_29191,N_28270,N_27819);
and U29192 (N_29192,N_27779,N_27772);
nor U29193 (N_29193,N_27824,N_28667);
xnor U29194 (N_29194,N_28653,N_28748);
and U29195 (N_29195,N_28442,N_28121);
xor U29196 (N_29196,N_27696,N_28553);
nor U29197 (N_29197,N_27798,N_28117);
nand U29198 (N_29198,N_28741,N_28111);
and U29199 (N_29199,N_27891,N_27702);
and U29200 (N_29200,N_27969,N_28271);
nand U29201 (N_29201,N_28708,N_28302);
and U29202 (N_29202,N_28501,N_28078);
or U29203 (N_29203,N_28721,N_28224);
nand U29204 (N_29204,N_27751,N_28229);
nand U29205 (N_29205,N_28123,N_28685);
nand U29206 (N_29206,N_28036,N_27935);
or U29207 (N_29207,N_27695,N_28344);
and U29208 (N_29208,N_28724,N_28559);
xnor U29209 (N_29209,N_28565,N_28314);
and U29210 (N_29210,N_27844,N_28381);
and U29211 (N_29211,N_28254,N_28717);
xnor U29212 (N_29212,N_27919,N_27617);
nor U29213 (N_29213,N_28337,N_28630);
or U29214 (N_29214,N_28714,N_28114);
nand U29215 (N_29215,N_28251,N_28276);
nand U29216 (N_29216,N_28252,N_28677);
nand U29217 (N_29217,N_28355,N_28558);
nand U29218 (N_29218,N_27705,N_27997);
nor U29219 (N_29219,N_28731,N_28404);
nand U29220 (N_29220,N_28180,N_28300);
and U29221 (N_29221,N_27936,N_27643);
and U29222 (N_29222,N_28108,N_27644);
or U29223 (N_29223,N_28776,N_27993);
nand U29224 (N_29224,N_27602,N_28408);
xnor U29225 (N_29225,N_28392,N_27979);
nor U29226 (N_29226,N_27905,N_28693);
xnor U29227 (N_29227,N_28201,N_28321);
or U29228 (N_29228,N_28530,N_27737);
xnor U29229 (N_29229,N_27964,N_28380);
nor U29230 (N_29230,N_28548,N_28455);
and U29231 (N_29231,N_27741,N_28167);
xor U29232 (N_29232,N_28181,N_27928);
or U29233 (N_29233,N_27847,N_27851);
nor U29234 (N_29234,N_27689,N_28055);
and U29235 (N_29235,N_28021,N_28615);
xnor U29236 (N_29236,N_27668,N_28172);
and U29237 (N_29237,N_28720,N_28485);
nand U29238 (N_29238,N_28202,N_28103);
and U29239 (N_29239,N_27910,N_28083);
xnor U29240 (N_29240,N_28406,N_28626);
xnor U29241 (N_29241,N_28758,N_28062);
xnor U29242 (N_29242,N_28231,N_27722);
xor U29243 (N_29243,N_28030,N_28556);
nor U29244 (N_29244,N_28773,N_27807);
and U29245 (N_29245,N_28697,N_28579);
xor U29246 (N_29246,N_28342,N_27835);
nor U29247 (N_29247,N_28539,N_28460);
nor U29248 (N_29248,N_27926,N_27796);
nor U29249 (N_29249,N_28275,N_27816);
xnor U29250 (N_29250,N_27716,N_28279);
or U29251 (N_29251,N_28739,N_27657);
nor U29252 (N_29252,N_28135,N_28437);
nor U29253 (N_29253,N_27797,N_27923);
or U29254 (N_29254,N_28576,N_28232);
or U29255 (N_29255,N_28657,N_27606);
xor U29256 (N_29256,N_28230,N_28010);
or U29257 (N_29257,N_28538,N_28386);
nor U29258 (N_29258,N_28389,N_27638);
and U29259 (N_29259,N_28750,N_27852);
and U29260 (N_29260,N_27795,N_28094);
and U29261 (N_29261,N_28264,N_28783);
xor U29262 (N_29262,N_28303,N_28190);
and U29263 (N_29263,N_28150,N_28045);
nor U29264 (N_29264,N_28421,N_28572);
or U29265 (N_29265,N_28352,N_28066);
and U29266 (N_29266,N_27791,N_28221);
nor U29267 (N_29267,N_28212,N_28446);
xor U29268 (N_29268,N_27875,N_27950);
nand U29269 (N_29269,N_28480,N_28411);
and U29270 (N_29270,N_28571,N_28526);
xor U29271 (N_29271,N_28005,N_28348);
nor U29272 (N_29272,N_28715,N_28057);
nand U29273 (N_29273,N_27770,N_27605);
nand U29274 (N_29274,N_27813,N_28509);
nand U29275 (N_29275,N_28417,N_28687);
or U29276 (N_29276,N_28160,N_28613);
or U29277 (N_29277,N_28698,N_28187);
nand U29278 (N_29278,N_28639,N_27888);
nor U29279 (N_29279,N_27907,N_28625);
nand U29280 (N_29280,N_28780,N_28068);
nor U29281 (N_29281,N_28239,N_28793);
or U29282 (N_29282,N_28619,N_28186);
nand U29283 (N_29283,N_27859,N_28356);
or U29284 (N_29284,N_27653,N_28709);
and U29285 (N_29285,N_28483,N_27706);
and U29286 (N_29286,N_27934,N_28131);
or U29287 (N_29287,N_27945,N_28575);
nand U29288 (N_29288,N_28611,N_28210);
xnor U29289 (N_29289,N_28608,N_27929);
xor U29290 (N_29290,N_27992,N_28474);
or U29291 (N_29291,N_27648,N_28058);
and U29292 (N_29292,N_28689,N_28235);
or U29293 (N_29293,N_28308,N_28661);
and U29294 (N_29294,N_28453,N_28044);
xor U29295 (N_29295,N_27848,N_27687);
nand U29296 (N_29296,N_28704,N_28228);
nor U29297 (N_29297,N_28781,N_27799);
nand U29298 (N_29298,N_27701,N_27642);
or U29299 (N_29299,N_27990,N_27959);
nand U29300 (N_29300,N_27984,N_28100);
and U29301 (N_29301,N_28313,N_28402);
or U29302 (N_29302,N_28673,N_28154);
or U29303 (N_29303,N_27818,N_27802);
xor U29304 (N_29304,N_27672,N_28304);
or U29305 (N_29305,N_28431,N_28234);
or U29306 (N_29306,N_28194,N_28711);
or U29307 (N_29307,N_28033,N_28450);
nand U29308 (N_29308,N_28140,N_27715);
and U29309 (N_29309,N_28378,N_28350);
xnor U29310 (N_29310,N_27733,N_28365);
or U29311 (N_29311,N_28298,N_27908);
xor U29312 (N_29312,N_27931,N_27630);
or U29313 (N_29313,N_28706,N_28125);
nor U29314 (N_29314,N_27983,N_28226);
nor U29315 (N_29315,N_28759,N_27933);
xor U29316 (N_29316,N_28241,N_27808);
nor U29317 (N_29317,N_27729,N_28009);
nand U29318 (N_29318,N_27961,N_27920);
and U29319 (N_29319,N_28542,N_28666);
nand U29320 (N_29320,N_27718,N_27927);
nand U29321 (N_29321,N_28602,N_28624);
nor U29322 (N_29322,N_28777,N_27604);
and U29323 (N_29323,N_28039,N_28070);
nand U29324 (N_29324,N_27697,N_27881);
nor U29325 (N_29325,N_27681,N_28517);
nand U29326 (N_29326,N_28737,N_28329);
xor U29327 (N_29327,N_28266,N_28785);
nor U29328 (N_29328,N_28645,N_28581);
xnor U29329 (N_29329,N_28151,N_27732);
nor U29330 (N_29330,N_27635,N_28452);
and U29331 (N_29331,N_28456,N_28678);
or U29332 (N_29332,N_28543,N_27953);
nand U29333 (N_29333,N_28048,N_27914);
nand U29334 (N_29334,N_28593,N_28430);
xor U29335 (N_29335,N_27615,N_28084);
or U29336 (N_29336,N_28347,N_28092);
xor U29337 (N_29337,N_28670,N_28171);
xnor U29338 (N_29338,N_28695,N_27661);
or U29339 (N_29339,N_28222,N_27872);
nor U29340 (N_29340,N_28601,N_28745);
xor U29341 (N_29341,N_27725,N_28663);
and U29342 (N_29342,N_28531,N_27740);
xor U29343 (N_29343,N_28278,N_28324);
nor U29344 (N_29344,N_28722,N_28361);
nor U29345 (N_29345,N_28511,N_27631);
nor U29346 (N_29346,N_28520,N_28240);
xor U29347 (N_29347,N_27654,N_28195);
and U29348 (N_29348,N_27708,N_28633);
xor U29349 (N_29349,N_28617,N_28197);
nand U29350 (N_29350,N_28562,N_27985);
nor U29351 (N_29351,N_27730,N_28003);
xnor U29352 (N_29352,N_27812,N_27900);
xor U29353 (N_29353,N_28334,N_28425);
nand U29354 (N_29354,N_28359,N_28286);
nor U29355 (N_29355,N_27686,N_28338);
nand U29356 (N_29356,N_27834,N_28025);
nor U29357 (N_29357,N_28138,N_28320);
xnor U29358 (N_29358,N_28246,N_28035);
xnor U29359 (N_29359,N_28243,N_28433);
or U29360 (N_29360,N_28535,N_27810);
nand U29361 (N_29361,N_28786,N_27782);
nor U29362 (N_29362,N_28521,N_28605);
nor U29363 (N_29363,N_28426,N_27904);
or U29364 (N_29364,N_27856,N_27645);
xnor U29365 (N_29365,N_28027,N_28047);
xor U29366 (N_29366,N_28120,N_28789);
xor U29367 (N_29367,N_28515,N_27924);
and U29368 (N_29368,N_27864,N_27880);
nor U29369 (N_29369,N_28156,N_28614);
or U29370 (N_29370,N_27860,N_28574);
nor U29371 (N_29371,N_28423,N_28219);
nand U29372 (N_29372,N_28132,N_27683);
and U29373 (N_29373,N_27712,N_27632);
and U29374 (N_29374,N_27989,N_27823);
or U29375 (N_29375,N_28413,N_28577);
xnor U29376 (N_29376,N_27925,N_28029);
nor U29377 (N_29377,N_27735,N_28596);
nand U29378 (N_29378,N_28060,N_28582);
nand U29379 (N_29379,N_28597,N_28429);
nand U29380 (N_29380,N_28250,N_27909);
nor U29381 (N_29381,N_28294,N_27822);
xnor U29382 (N_29382,N_27767,N_28105);
nor U29383 (N_29383,N_28506,N_27676);
nand U29384 (N_29384,N_27748,N_27809);
nor U29385 (N_29385,N_28458,N_28774);
or U29386 (N_29386,N_28262,N_28702);
nand U29387 (N_29387,N_28616,N_28155);
and U29388 (N_29388,N_27738,N_28257);
xnor U29389 (N_29389,N_27801,N_28468);
and U29390 (N_29390,N_28183,N_28519);
nand U29391 (N_29391,N_28586,N_27627);
nor U29392 (N_29392,N_28583,N_28319);
nor U29393 (N_29393,N_28051,N_28554);
nor U29394 (N_29394,N_28382,N_28599);
and U29395 (N_29395,N_28627,N_27917);
nand U29396 (N_29396,N_28649,N_27650);
nand U29397 (N_29397,N_28457,N_28004);
nor U29398 (N_29398,N_28403,N_27623);
and U29399 (N_29399,N_28494,N_28326);
nor U29400 (N_29400,N_28292,N_28542);
and U29401 (N_29401,N_28757,N_28214);
or U29402 (N_29402,N_28404,N_27678);
xor U29403 (N_29403,N_28429,N_27785);
and U29404 (N_29404,N_27964,N_28211);
and U29405 (N_29405,N_28771,N_28206);
and U29406 (N_29406,N_28231,N_28024);
and U29407 (N_29407,N_28724,N_27634);
xor U29408 (N_29408,N_28057,N_27872);
nor U29409 (N_29409,N_28795,N_28142);
nand U29410 (N_29410,N_28590,N_28239);
nand U29411 (N_29411,N_27609,N_28540);
nand U29412 (N_29412,N_28231,N_28318);
nand U29413 (N_29413,N_28038,N_28598);
and U29414 (N_29414,N_28232,N_27780);
nand U29415 (N_29415,N_28280,N_28311);
xor U29416 (N_29416,N_27883,N_28467);
nor U29417 (N_29417,N_28182,N_28649);
or U29418 (N_29418,N_28792,N_28352);
nand U29419 (N_29419,N_28693,N_27612);
nor U29420 (N_29420,N_28479,N_28107);
and U29421 (N_29421,N_27830,N_28746);
nand U29422 (N_29422,N_28540,N_28658);
and U29423 (N_29423,N_28783,N_28665);
and U29424 (N_29424,N_28000,N_27867);
xnor U29425 (N_29425,N_28493,N_28110);
nand U29426 (N_29426,N_28785,N_28786);
and U29427 (N_29427,N_28546,N_27687);
nor U29428 (N_29428,N_27992,N_28455);
nand U29429 (N_29429,N_27902,N_28757);
nand U29430 (N_29430,N_28159,N_28433);
or U29431 (N_29431,N_28588,N_28305);
xnor U29432 (N_29432,N_28100,N_28484);
nor U29433 (N_29433,N_27638,N_28742);
nor U29434 (N_29434,N_28310,N_28214);
nand U29435 (N_29435,N_28279,N_28469);
xnor U29436 (N_29436,N_27942,N_27664);
xnor U29437 (N_29437,N_27817,N_28648);
xor U29438 (N_29438,N_28457,N_27657);
nand U29439 (N_29439,N_28246,N_28102);
nor U29440 (N_29440,N_27930,N_28305);
nor U29441 (N_29441,N_28558,N_28131);
or U29442 (N_29442,N_28024,N_27917);
nand U29443 (N_29443,N_28606,N_28741);
nand U29444 (N_29444,N_28505,N_28429);
or U29445 (N_29445,N_27691,N_27836);
and U29446 (N_29446,N_28150,N_28120);
or U29447 (N_29447,N_28699,N_27865);
nor U29448 (N_29448,N_27757,N_28135);
xor U29449 (N_29449,N_28288,N_28652);
nand U29450 (N_29450,N_28582,N_28109);
and U29451 (N_29451,N_28113,N_27714);
nand U29452 (N_29452,N_27761,N_27925);
or U29453 (N_29453,N_27865,N_28721);
xor U29454 (N_29454,N_28035,N_28406);
xor U29455 (N_29455,N_28556,N_27848);
nor U29456 (N_29456,N_27844,N_28066);
nand U29457 (N_29457,N_27723,N_27708);
nand U29458 (N_29458,N_28095,N_28102);
nand U29459 (N_29459,N_27830,N_27854);
nand U29460 (N_29460,N_28538,N_28312);
and U29461 (N_29461,N_28551,N_28078);
xnor U29462 (N_29462,N_28496,N_28077);
nor U29463 (N_29463,N_28085,N_27704);
and U29464 (N_29464,N_28104,N_28409);
nor U29465 (N_29465,N_28395,N_27890);
nand U29466 (N_29466,N_27947,N_28678);
xor U29467 (N_29467,N_28525,N_28284);
or U29468 (N_29468,N_28524,N_28095);
nor U29469 (N_29469,N_28329,N_28142);
nor U29470 (N_29470,N_27923,N_27910);
or U29471 (N_29471,N_28752,N_28039);
or U29472 (N_29472,N_28084,N_28247);
and U29473 (N_29473,N_28331,N_28093);
and U29474 (N_29474,N_27943,N_28599);
xor U29475 (N_29475,N_28122,N_28776);
or U29476 (N_29476,N_28416,N_28266);
xor U29477 (N_29477,N_27737,N_28544);
and U29478 (N_29478,N_28354,N_28063);
nand U29479 (N_29479,N_27750,N_27960);
and U29480 (N_29480,N_27918,N_27608);
and U29481 (N_29481,N_28470,N_28728);
nor U29482 (N_29482,N_28023,N_28444);
and U29483 (N_29483,N_28231,N_27613);
xor U29484 (N_29484,N_27963,N_27825);
or U29485 (N_29485,N_27819,N_28319);
and U29486 (N_29486,N_28374,N_27692);
or U29487 (N_29487,N_27697,N_28493);
and U29488 (N_29488,N_28089,N_27850);
nand U29489 (N_29489,N_28266,N_28323);
and U29490 (N_29490,N_28312,N_27870);
xnor U29491 (N_29491,N_28270,N_27907);
and U29492 (N_29492,N_28793,N_27930);
nor U29493 (N_29493,N_27886,N_28476);
and U29494 (N_29494,N_28347,N_28574);
nand U29495 (N_29495,N_27839,N_28675);
xnor U29496 (N_29496,N_28556,N_27987);
nor U29497 (N_29497,N_28748,N_27757);
and U29498 (N_29498,N_27883,N_27906);
xnor U29499 (N_29499,N_28573,N_28268);
and U29500 (N_29500,N_28328,N_28554);
nor U29501 (N_29501,N_28124,N_27700);
or U29502 (N_29502,N_28084,N_28185);
or U29503 (N_29503,N_27810,N_27645);
and U29504 (N_29504,N_28458,N_28171);
and U29505 (N_29505,N_28789,N_28629);
or U29506 (N_29506,N_28165,N_28317);
xor U29507 (N_29507,N_28245,N_28279);
xnor U29508 (N_29508,N_28787,N_28686);
nand U29509 (N_29509,N_28161,N_28396);
or U29510 (N_29510,N_27881,N_27739);
and U29511 (N_29511,N_28411,N_28484);
or U29512 (N_29512,N_28675,N_28692);
xor U29513 (N_29513,N_28660,N_28051);
and U29514 (N_29514,N_28628,N_27910);
or U29515 (N_29515,N_28036,N_28606);
and U29516 (N_29516,N_27846,N_28361);
nor U29517 (N_29517,N_28088,N_28433);
or U29518 (N_29518,N_28584,N_27856);
xor U29519 (N_29519,N_27732,N_28077);
nor U29520 (N_29520,N_28486,N_28653);
nor U29521 (N_29521,N_28770,N_28327);
nor U29522 (N_29522,N_28079,N_27622);
or U29523 (N_29523,N_28055,N_27999);
and U29524 (N_29524,N_27634,N_27753);
or U29525 (N_29525,N_28336,N_28027);
and U29526 (N_29526,N_28765,N_28150);
xor U29527 (N_29527,N_28131,N_27735);
nand U29528 (N_29528,N_28104,N_27912);
nand U29529 (N_29529,N_28682,N_27759);
nand U29530 (N_29530,N_27766,N_28151);
and U29531 (N_29531,N_27932,N_27615);
or U29532 (N_29532,N_27623,N_28555);
xnor U29533 (N_29533,N_28593,N_28347);
nor U29534 (N_29534,N_28480,N_27931);
nor U29535 (N_29535,N_27970,N_27961);
and U29536 (N_29536,N_28405,N_28646);
and U29537 (N_29537,N_28169,N_28532);
and U29538 (N_29538,N_28367,N_28571);
nor U29539 (N_29539,N_28170,N_27695);
or U29540 (N_29540,N_28410,N_28143);
xor U29541 (N_29541,N_28565,N_28350);
or U29542 (N_29542,N_27827,N_28623);
nand U29543 (N_29543,N_27854,N_27931);
nor U29544 (N_29544,N_27752,N_28450);
xor U29545 (N_29545,N_28299,N_27696);
and U29546 (N_29546,N_28170,N_27739);
nor U29547 (N_29547,N_27767,N_28352);
nand U29548 (N_29548,N_27891,N_28210);
or U29549 (N_29549,N_27703,N_27971);
xnor U29550 (N_29550,N_28213,N_28185);
and U29551 (N_29551,N_28680,N_28715);
xor U29552 (N_29552,N_28729,N_28703);
nand U29553 (N_29553,N_27897,N_28290);
nand U29554 (N_29554,N_27848,N_28550);
nor U29555 (N_29555,N_28379,N_28591);
nand U29556 (N_29556,N_28315,N_28390);
and U29557 (N_29557,N_28111,N_27830);
nor U29558 (N_29558,N_27634,N_28386);
nor U29559 (N_29559,N_28509,N_28727);
and U29560 (N_29560,N_28070,N_28742);
nor U29561 (N_29561,N_28252,N_28726);
xor U29562 (N_29562,N_27997,N_27987);
and U29563 (N_29563,N_28604,N_28458);
xnor U29564 (N_29564,N_28708,N_28697);
xor U29565 (N_29565,N_28789,N_27922);
xor U29566 (N_29566,N_27605,N_27628);
nor U29567 (N_29567,N_27603,N_28091);
nor U29568 (N_29568,N_28127,N_27726);
or U29569 (N_29569,N_28656,N_28338);
nand U29570 (N_29570,N_28339,N_28078);
and U29571 (N_29571,N_27970,N_27812);
nand U29572 (N_29572,N_27652,N_27663);
or U29573 (N_29573,N_28212,N_28041);
or U29574 (N_29574,N_27939,N_27848);
xnor U29575 (N_29575,N_28087,N_27863);
xor U29576 (N_29576,N_27645,N_28676);
and U29577 (N_29577,N_28734,N_27735);
xnor U29578 (N_29578,N_28179,N_28057);
nand U29579 (N_29579,N_27977,N_28245);
or U29580 (N_29580,N_28511,N_28119);
nand U29581 (N_29581,N_28314,N_28087);
xnor U29582 (N_29582,N_27606,N_27753);
and U29583 (N_29583,N_27917,N_28602);
nand U29584 (N_29584,N_28225,N_27734);
xor U29585 (N_29585,N_28354,N_27850);
and U29586 (N_29586,N_28288,N_28498);
xor U29587 (N_29587,N_28635,N_28411);
nand U29588 (N_29588,N_27871,N_27685);
or U29589 (N_29589,N_27698,N_27617);
or U29590 (N_29590,N_27852,N_28289);
xor U29591 (N_29591,N_28686,N_28437);
nor U29592 (N_29592,N_28374,N_28193);
or U29593 (N_29593,N_28285,N_28303);
nand U29594 (N_29594,N_27635,N_28048);
nand U29595 (N_29595,N_28047,N_28340);
and U29596 (N_29596,N_28645,N_27908);
xor U29597 (N_29597,N_28475,N_28789);
and U29598 (N_29598,N_27896,N_28731);
nor U29599 (N_29599,N_28724,N_28741);
xnor U29600 (N_29600,N_28095,N_28308);
nand U29601 (N_29601,N_28320,N_27767);
nor U29602 (N_29602,N_28368,N_28458);
and U29603 (N_29603,N_28389,N_27801);
nand U29604 (N_29604,N_27859,N_28199);
nand U29605 (N_29605,N_28729,N_28573);
and U29606 (N_29606,N_28333,N_28731);
and U29607 (N_29607,N_27923,N_27976);
xnor U29608 (N_29608,N_27729,N_28043);
and U29609 (N_29609,N_28267,N_28178);
nand U29610 (N_29610,N_28214,N_28794);
nor U29611 (N_29611,N_28658,N_27615);
and U29612 (N_29612,N_28480,N_28113);
and U29613 (N_29613,N_28526,N_28523);
nand U29614 (N_29614,N_28610,N_28399);
or U29615 (N_29615,N_27849,N_27806);
xor U29616 (N_29616,N_28677,N_28701);
nand U29617 (N_29617,N_28735,N_28309);
and U29618 (N_29618,N_27753,N_28389);
or U29619 (N_29619,N_28797,N_27628);
or U29620 (N_29620,N_27736,N_28386);
nor U29621 (N_29621,N_28326,N_28055);
nand U29622 (N_29622,N_28487,N_28749);
nand U29623 (N_29623,N_27731,N_27615);
and U29624 (N_29624,N_28719,N_28029);
nand U29625 (N_29625,N_28518,N_27837);
and U29626 (N_29626,N_28157,N_27763);
and U29627 (N_29627,N_28798,N_28508);
nor U29628 (N_29628,N_27894,N_28429);
xnor U29629 (N_29629,N_27618,N_28129);
xnor U29630 (N_29630,N_28257,N_28565);
nand U29631 (N_29631,N_28779,N_28679);
or U29632 (N_29632,N_27774,N_27844);
nand U29633 (N_29633,N_27754,N_27682);
or U29634 (N_29634,N_27892,N_28064);
or U29635 (N_29635,N_28741,N_27693);
nor U29636 (N_29636,N_27694,N_28645);
and U29637 (N_29637,N_28739,N_27748);
nand U29638 (N_29638,N_28718,N_28748);
and U29639 (N_29639,N_27655,N_28186);
and U29640 (N_29640,N_28048,N_28208);
xor U29641 (N_29641,N_28145,N_28286);
and U29642 (N_29642,N_27633,N_27935);
nand U29643 (N_29643,N_27730,N_27884);
xor U29644 (N_29644,N_28779,N_28066);
nor U29645 (N_29645,N_27905,N_28411);
nor U29646 (N_29646,N_28099,N_28014);
or U29647 (N_29647,N_27905,N_28645);
nand U29648 (N_29648,N_28306,N_28036);
nand U29649 (N_29649,N_28141,N_27648);
or U29650 (N_29650,N_28440,N_28055);
nor U29651 (N_29651,N_28149,N_28164);
and U29652 (N_29652,N_28387,N_28172);
nor U29653 (N_29653,N_28296,N_28477);
nand U29654 (N_29654,N_28222,N_28118);
or U29655 (N_29655,N_28682,N_27868);
nand U29656 (N_29656,N_28197,N_28655);
and U29657 (N_29657,N_28505,N_28717);
nor U29658 (N_29658,N_28229,N_27707);
or U29659 (N_29659,N_28463,N_27618);
xnor U29660 (N_29660,N_28476,N_28658);
and U29661 (N_29661,N_27977,N_28191);
xnor U29662 (N_29662,N_27601,N_28728);
and U29663 (N_29663,N_28608,N_28797);
and U29664 (N_29664,N_28131,N_27703);
nand U29665 (N_29665,N_28707,N_28435);
xor U29666 (N_29666,N_28741,N_28337);
nand U29667 (N_29667,N_27849,N_28696);
nor U29668 (N_29668,N_27889,N_27607);
or U29669 (N_29669,N_28763,N_28791);
nand U29670 (N_29670,N_27910,N_27758);
and U29671 (N_29671,N_27746,N_28027);
and U29672 (N_29672,N_28494,N_28378);
nand U29673 (N_29673,N_28678,N_28112);
and U29674 (N_29674,N_28722,N_28763);
nor U29675 (N_29675,N_27601,N_28704);
nand U29676 (N_29676,N_28484,N_27724);
and U29677 (N_29677,N_27899,N_28062);
nor U29678 (N_29678,N_28077,N_28772);
and U29679 (N_29679,N_28179,N_28089);
nand U29680 (N_29680,N_27605,N_27643);
and U29681 (N_29681,N_28067,N_28103);
xnor U29682 (N_29682,N_28764,N_28372);
nand U29683 (N_29683,N_28574,N_28395);
and U29684 (N_29684,N_27797,N_28673);
nand U29685 (N_29685,N_27793,N_27997);
xnor U29686 (N_29686,N_28564,N_28358);
or U29687 (N_29687,N_28399,N_28250);
nor U29688 (N_29688,N_27606,N_28590);
and U29689 (N_29689,N_27654,N_28537);
nand U29690 (N_29690,N_28383,N_28403);
nand U29691 (N_29691,N_27818,N_28650);
xor U29692 (N_29692,N_28490,N_27656);
and U29693 (N_29693,N_27996,N_28239);
nor U29694 (N_29694,N_28460,N_27929);
or U29695 (N_29695,N_28380,N_27770);
nor U29696 (N_29696,N_28434,N_28431);
nand U29697 (N_29697,N_28689,N_27724);
nand U29698 (N_29698,N_28199,N_27808);
nand U29699 (N_29699,N_28556,N_28136);
nor U29700 (N_29700,N_28736,N_28283);
and U29701 (N_29701,N_28316,N_28294);
nor U29702 (N_29702,N_27903,N_28065);
xnor U29703 (N_29703,N_28684,N_27902);
nand U29704 (N_29704,N_28663,N_28119);
nand U29705 (N_29705,N_27797,N_28292);
xor U29706 (N_29706,N_28467,N_28475);
xor U29707 (N_29707,N_28445,N_28129);
nor U29708 (N_29708,N_28251,N_28201);
and U29709 (N_29709,N_28660,N_28745);
nor U29710 (N_29710,N_27634,N_27892);
and U29711 (N_29711,N_28581,N_27624);
xnor U29712 (N_29712,N_28022,N_28477);
xnor U29713 (N_29713,N_28239,N_27797);
xnor U29714 (N_29714,N_28593,N_28060);
nand U29715 (N_29715,N_27738,N_27990);
xor U29716 (N_29716,N_28620,N_28209);
nand U29717 (N_29717,N_28713,N_28273);
and U29718 (N_29718,N_28370,N_27716);
and U29719 (N_29719,N_28662,N_28054);
nand U29720 (N_29720,N_28473,N_27688);
and U29721 (N_29721,N_27699,N_27647);
or U29722 (N_29722,N_27655,N_28667);
or U29723 (N_29723,N_28489,N_28438);
nor U29724 (N_29724,N_28678,N_28679);
nand U29725 (N_29725,N_28096,N_27813);
or U29726 (N_29726,N_27789,N_27737);
or U29727 (N_29727,N_28352,N_28482);
and U29728 (N_29728,N_28062,N_27914);
nor U29729 (N_29729,N_28778,N_28372);
nor U29730 (N_29730,N_27929,N_27850);
nand U29731 (N_29731,N_28125,N_28133);
nor U29732 (N_29732,N_27921,N_28141);
or U29733 (N_29733,N_28567,N_28461);
or U29734 (N_29734,N_28590,N_28428);
and U29735 (N_29735,N_28042,N_28546);
xnor U29736 (N_29736,N_27810,N_27833);
and U29737 (N_29737,N_28716,N_27848);
nand U29738 (N_29738,N_28691,N_28662);
and U29739 (N_29739,N_28603,N_27752);
or U29740 (N_29740,N_27695,N_28267);
or U29741 (N_29741,N_27754,N_27739);
nor U29742 (N_29742,N_27836,N_27656);
nand U29743 (N_29743,N_28144,N_28709);
xnor U29744 (N_29744,N_27913,N_28408);
xnor U29745 (N_29745,N_28228,N_28619);
nand U29746 (N_29746,N_28410,N_28038);
nand U29747 (N_29747,N_28182,N_28189);
or U29748 (N_29748,N_28788,N_28666);
or U29749 (N_29749,N_27765,N_28756);
nand U29750 (N_29750,N_28330,N_28384);
nor U29751 (N_29751,N_28704,N_28335);
xnor U29752 (N_29752,N_28486,N_28602);
or U29753 (N_29753,N_28422,N_28397);
nand U29754 (N_29754,N_28207,N_27992);
xnor U29755 (N_29755,N_28222,N_27659);
nand U29756 (N_29756,N_28487,N_28361);
nor U29757 (N_29757,N_28068,N_28132);
xor U29758 (N_29758,N_28596,N_28660);
and U29759 (N_29759,N_27855,N_28682);
nand U29760 (N_29760,N_28119,N_27620);
or U29761 (N_29761,N_28633,N_27824);
nand U29762 (N_29762,N_28288,N_28265);
or U29763 (N_29763,N_27973,N_27993);
nand U29764 (N_29764,N_28566,N_28018);
or U29765 (N_29765,N_28779,N_28063);
and U29766 (N_29766,N_28754,N_27701);
nor U29767 (N_29767,N_27738,N_28347);
and U29768 (N_29768,N_27636,N_28072);
and U29769 (N_29769,N_27607,N_28019);
nor U29770 (N_29770,N_27815,N_28099);
xnor U29771 (N_29771,N_28621,N_27961);
and U29772 (N_29772,N_28519,N_27642);
nand U29773 (N_29773,N_28118,N_28281);
xnor U29774 (N_29774,N_28342,N_28588);
or U29775 (N_29775,N_27827,N_28339);
and U29776 (N_29776,N_28307,N_28255);
nor U29777 (N_29777,N_28053,N_28465);
or U29778 (N_29778,N_28401,N_27895);
nand U29779 (N_29779,N_27828,N_28290);
xnor U29780 (N_29780,N_28354,N_28029);
or U29781 (N_29781,N_27943,N_28657);
nand U29782 (N_29782,N_28771,N_27850);
xnor U29783 (N_29783,N_28578,N_28210);
nand U29784 (N_29784,N_28325,N_28024);
nor U29785 (N_29785,N_28170,N_27995);
and U29786 (N_29786,N_28472,N_28467);
and U29787 (N_29787,N_28609,N_27788);
and U29788 (N_29788,N_28777,N_28128);
or U29789 (N_29789,N_28630,N_28578);
nand U29790 (N_29790,N_28391,N_28414);
xnor U29791 (N_29791,N_28577,N_27950);
and U29792 (N_29792,N_28663,N_28382);
and U29793 (N_29793,N_28778,N_28373);
or U29794 (N_29794,N_28679,N_28791);
nor U29795 (N_29795,N_28275,N_27756);
and U29796 (N_29796,N_27985,N_27754);
and U29797 (N_29797,N_28211,N_27612);
nor U29798 (N_29798,N_27622,N_28062);
nand U29799 (N_29799,N_27992,N_28538);
xnor U29800 (N_29800,N_27733,N_28530);
xnor U29801 (N_29801,N_28202,N_27999);
or U29802 (N_29802,N_28569,N_28781);
or U29803 (N_29803,N_28101,N_27978);
and U29804 (N_29804,N_28244,N_28778);
xor U29805 (N_29805,N_28112,N_27616);
nand U29806 (N_29806,N_28548,N_27901);
and U29807 (N_29807,N_27876,N_28230);
and U29808 (N_29808,N_27919,N_28683);
xnor U29809 (N_29809,N_28400,N_28236);
or U29810 (N_29810,N_27628,N_28513);
and U29811 (N_29811,N_28065,N_28249);
xnor U29812 (N_29812,N_27620,N_28069);
xor U29813 (N_29813,N_28366,N_28202);
nor U29814 (N_29814,N_27779,N_27824);
nor U29815 (N_29815,N_27745,N_27866);
xor U29816 (N_29816,N_28626,N_28499);
and U29817 (N_29817,N_27869,N_28768);
and U29818 (N_29818,N_27680,N_27853);
or U29819 (N_29819,N_28134,N_28276);
nand U29820 (N_29820,N_28680,N_27753);
xnor U29821 (N_29821,N_27925,N_27704);
nand U29822 (N_29822,N_27692,N_27940);
nor U29823 (N_29823,N_27891,N_27873);
xor U29824 (N_29824,N_28483,N_27620);
nand U29825 (N_29825,N_28540,N_28404);
and U29826 (N_29826,N_28502,N_27642);
nor U29827 (N_29827,N_28277,N_28716);
nor U29828 (N_29828,N_28384,N_27745);
xor U29829 (N_29829,N_27678,N_27861);
nor U29830 (N_29830,N_27716,N_27697);
nand U29831 (N_29831,N_27729,N_28318);
nor U29832 (N_29832,N_28608,N_27732);
nand U29833 (N_29833,N_28563,N_28346);
nand U29834 (N_29834,N_28432,N_28095);
nor U29835 (N_29835,N_28449,N_27830);
xor U29836 (N_29836,N_28633,N_28006);
or U29837 (N_29837,N_27746,N_27931);
or U29838 (N_29838,N_28221,N_28740);
or U29839 (N_29839,N_28303,N_27704);
xor U29840 (N_29840,N_28525,N_28201);
nor U29841 (N_29841,N_28091,N_28041);
nand U29842 (N_29842,N_28191,N_28479);
xor U29843 (N_29843,N_28454,N_27878);
nand U29844 (N_29844,N_28377,N_28137);
nor U29845 (N_29845,N_28517,N_27845);
xnor U29846 (N_29846,N_28003,N_27669);
and U29847 (N_29847,N_28040,N_28080);
nor U29848 (N_29848,N_27998,N_27961);
nand U29849 (N_29849,N_28729,N_28099);
or U29850 (N_29850,N_28133,N_28457);
nand U29851 (N_29851,N_27654,N_28564);
nor U29852 (N_29852,N_28460,N_27981);
and U29853 (N_29853,N_28754,N_28451);
nand U29854 (N_29854,N_27837,N_27670);
xnor U29855 (N_29855,N_27802,N_28026);
or U29856 (N_29856,N_28741,N_28608);
and U29857 (N_29857,N_27621,N_28143);
nand U29858 (N_29858,N_28126,N_27634);
xnor U29859 (N_29859,N_27686,N_28356);
or U29860 (N_29860,N_27922,N_27666);
and U29861 (N_29861,N_28396,N_28329);
xnor U29862 (N_29862,N_28028,N_28499);
or U29863 (N_29863,N_28236,N_28609);
and U29864 (N_29864,N_28787,N_27635);
nor U29865 (N_29865,N_28766,N_28751);
or U29866 (N_29866,N_28048,N_28035);
or U29867 (N_29867,N_28532,N_27845);
and U29868 (N_29868,N_28018,N_28513);
or U29869 (N_29869,N_27875,N_28221);
nand U29870 (N_29870,N_28526,N_28281);
or U29871 (N_29871,N_28739,N_28042);
or U29872 (N_29872,N_28796,N_28112);
xor U29873 (N_29873,N_28330,N_28334);
xnor U29874 (N_29874,N_28221,N_28787);
xor U29875 (N_29875,N_27607,N_28703);
and U29876 (N_29876,N_28316,N_28660);
nand U29877 (N_29877,N_28148,N_27676);
or U29878 (N_29878,N_28051,N_28440);
or U29879 (N_29879,N_28336,N_28006);
nor U29880 (N_29880,N_28193,N_27636);
nor U29881 (N_29881,N_28718,N_27950);
nor U29882 (N_29882,N_28506,N_28702);
xor U29883 (N_29883,N_28537,N_28172);
nand U29884 (N_29884,N_28060,N_28015);
xor U29885 (N_29885,N_28585,N_28567);
xor U29886 (N_29886,N_28283,N_28323);
nand U29887 (N_29887,N_28465,N_27661);
or U29888 (N_29888,N_28385,N_27628);
or U29889 (N_29889,N_27610,N_27863);
nor U29890 (N_29890,N_28189,N_27803);
xnor U29891 (N_29891,N_28517,N_27817);
nor U29892 (N_29892,N_28749,N_28393);
and U29893 (N_29893,N_28094,N_27952);
nor U29894 (N_29894,N_28297,N_28721);
or U29895 (N_29895,N_27602,N_28101);
nor U29896 (N_29896,N_28773,N_27957);
xnor U29897 (N_29897,N_28488,N_28036);
and U29898 (N_29898,N_28058,N_28159);
xor U29899 (N_29899,N_27703,N_27821);
and U29900 (N_29900,N_28157,N_27911);
xor U29901 (N_29901,N_27925,N_28200);
or U29902 (N_29902,N_28157,N_28343);
nand U29903 (N_29903,N_28796,N_28452);
or U29904 (N_29904,N_28521,N_28249);
xor U29905 (N_29905,N_27774,N_28320);
nor U29906 (N_29906,N_28544,N_27619);
and U29907 (N_29907,N_28387,N_28789);
or U29908 (N_29908,N_28013,N_28386);
nor U29909 (N_29909,N_27897,N_27947);
xor U29910 (N_29910,N_28231,N_28360);
xor U29911 (N_29911,N_28659,N_28091);
nand U29912 (N_29912,N_28509,N_27626);
nand U29913 (N_29913,N_28071,N_28184);
or U29914 (N_29914,N_27824,N_27882);
nand U29915 (N_29915,N_28688,N_28403);
and U29916 (N_29916,N_28164,N_28324);
xnor U29917 (N_29917,N_28001,N_28506);
xor U29918 (N_29918,N_27712,N_28697);
and U29919 (N_29919,N_28344,N_28760);
nor U29920 (N_29920,N_27945,N_28681);
nand U29921 (N_29921,N_28512,N_28286);
nor U29922 (N_29922,N_27729,N_27733);
nand U29923 (N_29923,N_27968,N_28224);
or U29924 (N_29924,N_28522,N_27683);
nor U29925 (N_29925,N_28435,N_28089);
and U29926 (N_29926,N_27846,N_28484);
and U29927 (N_29927,N_27782,N_28659);
xnor U29928 (N_29928,N_28222,N_28471);
or U29929 (N_29929,N_27828,N_28274);
or U29930 (N_29930,N_28270,N_27856);
and U29931 (N_29931,N_28305,N_28392);
or U29932 (N_29932,N_28315,N_27865);
xnor U29933 (N_29933,N_27726,N_28574);
nand U29934 (N_29934,N_28349,N_28724);
nand U29935 (N_29935,N_28519,N_27819);
nor U29936 (N_29936,N_28361,N_27915);
nor U29937 (N_29937,N_27776,N_28560);
xor U29938 (N_29938,N_28175,N_28387);
nand U29939 (N_29939,N_28231,N_28470);
nand U29940 (N_29940,N_27675,N_28076);
nand U29941 (N_29941,N_27777,N_27951);
or U29942 (N_29942,N_27841,N_27972);
nand U29943 (N_29943,N_28398,N_28225);
nand U29944 (N_29944,N_27942,N_27812);
and U29945 (N_29945,N_27886,N_28158);
nor U29946 (N_29946,N_28437,N_27837);
or U29947 (N_29947,N_28275,N_28256);
nand U29948 (N_29948,N_28381,N_28023);
xor U29949 (N_29949,N_27671,N_28451);
or U29950 (N_29950,N_28256,N_27883);
and U29951 (N_29951,N_28119,N_27864);
nor U29952 (N_29952,N_27879,N_28579);
nand U29953 (N_29953,N_27800,N_27705);
nor U29954 (N_29954,N_28066,N_28008);
nand U29955 (N_29955,N_28038,N_27906);
or U29956 (N_29956,N_28431,N_27855);
xor U29957 (N_29957,N_28663,N_27967);
nor U29958 (N_29958,N_28135,N_27735);
or U29959 (N_29959,N_28644,N_28587);
xnor U29960 (N_29960,N_28644,N_27810);
xor U29961 (N_29961,N_27880,N_27982);
xnor U29962 (N_29962,N_28095,N_27804);
xor U29963 (N_29963,N_27688,N_28238);
nor U29964 (N_29964,N_28381,N_28277);
xnor U29965 (N_29965,N_28521,N_28333);
and U29966 (N_29966,N_27713,N_27677);
or U29967 (N_29967,N_28095,N_28596);
nor U29968 (N_29968,N_28518,N_28222);
and U29969 (N_29969,N_28440,N_28243);
nor U29970 (N_29970,N_28565,N_28306);
nand U29971 (N_29971,N_28398,N_27669);
nand U29972 (N_29972,N_27706,N_28751);
xnor U29973 (N_29973,N_28480,N_27756);
nor U29974 (N_29974,N_28385,N_28236);
or U29975 (N_29975,N_28610,N_27698);
nand U29976 (N_29976,N_28371,N_28102);
nor U29977 (N_29977,N_28259,N_28049);
nor U29978 (N_29978,N_28329,N_27928);
nand U29979 (N_29979,N_27675,N_28537);
and U29980 (N_29980,N_27961,N_28712);
and U29981 (N_29981,N_27719,N_28405);
xor U29982 (N_29982,N_27994,N_28148);
nor U29983 (N_29983,N_28150,N_28506);
or U29984 (N_29984,N_27918,N_28074);
nor U29985 (N_29985,N_28082,N_28168);
nor U29986 (N_29986,N_27881,N_27969);
nor U29987 (N_29987,N_27641,N_28023);
nand U29988 (N_29988,N_28723,N_27727);
nand U29989 (N_29989,N_28607,N_28727);
nor U29990 (N_29990,N_27889,N_28169);
nand U29991 (N_29991,N_28428,N_28235);
nor U29992 (N_29992,N_28494,N_28125);
and U29993 (N_29993,N_28736,N_28621);
and U29994 (N_29994,N_27994,N_28206);
nand U29995 (N_29995,N_28613,N_28447);
and U29996 (N_29996,N_28610,N_28604);
nor U29997 (N_29997,N_28725,N_28665);
and U29998 (N_29998,N_28505,N_28096);
xor U29999 (N_29999,N_27805,N_27615);
xnor UO_0 (O_0,N_28847,N_29509);
and UO_1 (O_1,N_29408,N_29203);
nand UO_2 (O_2,N_28991,N_29834);
nor UO_3 (O_3,N_29751,N_29764);
nor UO_4 (O_4,N_29972,N_29132);
and UO_5 (O_5,N_28875,N_29676);
nor UO_6 (O_6,N_29853,N_29713);
nor UO_7 (O_7,N_29877,N_29559);
xor UO_8 (O_8,N_29033,N_29224);
and UO_9 (O_9,N_29611,N_29695);
xnor UO_10 (O_10,N_29083,N_29650);
or UO_11 (O_11,N_29534,N_29946);
and UO_12 (O_12,N_29384,N_29626);
nand UO_13 (O_13,N_29291,N_29304);
nand UO_14 (O_14,N_29953,N_29613);
nor UO_15 (O_15,N_29097,N_29682);
nand UO_16 (O_16,N_29598,N_28965);
nor UO_17 (O_17,N_29010,N_29423);
nor UO_18 (O_18,N_29466,N_28812);
xor UO_19 (O_19,N_29893,N_29225);
nor UO_20 (O_20,N_29744,N_29388);
or UO_21 (O_21,N_28859,N_29678);
or UO_22 (O_22,N_29298,N_29257);
or UO_23 (O_23,N_28919,N_29757);
nand UO_24 (O_24,N_29400,N_29206);
nand UO_25 (O_25,N_29440,N_29797);
and UO_26 (O_26,N_29443,N_29868);
nand UO_27 (O_27,N_28878,N_29831);
nand UO_28 (O_28,N_29560,N_29832);
nand UO_29 (O_29,N_29036,N_29507);
nor UO_30 (O_30,N_29873,N_29147);
nand UO_31 (O_31,N_28906,N_29951);
and UO_32 (O_32,N_28876,N_29092);
or UO_33 (O_33,N_29639,N_29102);
and UO_34 (O_34,N_29374,N_29531);
and UO_35 (O_35,N_29821,N_29745);
xor UO_36 (O_36,N_29251,N_28846);
nand UO_37 (O_37,N_29095,N_29841);
nor UO_38 (O_38,N_29530,N_28999);
nand UO_39 (O_39,N_29334,N_29077);
and UO_40 (O_40,N_29982,N_28888);
or UO_41 (O_41,N_29281,N_29902);
xnor UO_42 (O_42,N_28980,N_29199);
xnor UO_43 (O_43,N_29746,N_29414);
nand UO_44 (O_44,N_29546,N_28836);
or UO_45 (O_45,N_29581,N_29798);
nor UO_46 (O_46,N_29526,N_29485);
xor UO_47 (O_47,N_29382,N_29362);
nand UO_48 (O_48,N_29794,N_29048);
and UO_49 (O_49,N_29429,N_28867);
nand UO_50 (O_50,N_29035,N_29570);
or UO_51 (O_51,N_29996,N_29136);
nand UO_52 (O_52,N_29652,N_28938);
nor UO_53 (O_53,N_29365,N_29282);
nand UO_54 (O_54,N_29568,N_28889);
nor UO_55 (O_55,N_29645,N_29265);
xor UO_56 (O_56,N_28863,N_29619);
nor UO_57 (O_57,N_29002,N_29891);
nor UO_58 (O_58,N_29909,N_29532);
and UO_59 (O_59,N_29974,N_29734);
xor UO_60 (O_60,N_29822,N_28964);
nor UO_61 (O_61,N_29890,N_29514);
xor UO_62 (O_62,N_29826,N_29828);
or UO_63 (O_63,N_29226,N_28858);
or UO_64 (O_64,N_28913,N_29066);
nor UO_65 (O_65,N_29180,N_29958);
and UO_66 (O_66,N_29620,N_29335);
or UO_67 (O_67,N_28860,N_29741);
nor UO_68 (O_68,N_29005,N_29484);
nand UO_69 (O_69,N_29571,N_29394);
and UO_70 (O_70,N_28985,N_29163);
or UO_71 (O_71,N_29276,N_28885);
and UO_72 (O_72,N_28877,N_29270);
or UO_73 (O_73,N_29245,N_29959);
or UO_74 (O_74,N_29081,N_29451);
nand UO_75 (O_75,N_29082,N_28924);
and UO_76 (O_76,N_29504,N_29707);
nor UO_77 (O_77,N_28987,N_29855);
or UO_78 (O_78,N_29787,N_29754);
xnor UO_79 (O_79,N_29173,N_29896);
and UO_80 (O_80,N_28920,N_29973);
and UO_81 (O_81,N_28855,N_28975);
or UO_82 (O_82,N_29632,N_29904);
nor UO_83 (O_83,N_29494,N_29627);
nand UO_84 (O_84,N_29887,N_29486);
or UO_85 (O_85,N_29849,N_29729);
nor UO_86 (O_86,N_28970,N_29455);
nor UO_87 (O_87,N_28838,N_29057);
or UO_88 (O_88,N_29715,N_29011);
and UO_89 (O_89,N_29567,N_29814);
nand UO_90 (O_90,N_28911,N_29330);
or UO_91 (O_91,N_29178,N_29720);
and UO_92 (O_92,N_29123,N_29047);
and UO_93 (O_93,N_29943,N_29847);
xor UO_94 (O_94,N_29127,N_29419);
nand UO_95 (O_95,N_29422,N_29901);
or UO_96 (O_96,N_29612,N_29234);
and UO_97 (O_97,N_29587,N_29886);
xor UO_98 (O_98,N_28990,N_29774);
nor UO_99 (O_99,N_29080,N_29802);
and UO_100 (O_100,N_29054,N_29478);
nor UO_101 (O_101,N_29302,N_29823);
nor UO_102 (O_102,N_29447,N_28822);
and UO_103 (O_103,N_29964,N_29583);
nor UO_104 (O_104,N_29370,N_28946);
nor UO_105 (O_105,N_29777,N_28800);
and UO_106 (O_106,N_29029,N_28806);
nor UO_107 (O_107,N_28997,N_29174);
nand UO_108 (O_108,N_29194,N_29815);
nor UO_109 (O_109,N_28949,N_29043);
nor UO_110 (O_110,N_29966,N_29692);
nand UO_111 (O_111,N_28894,N_29089);
nand UO_112 (O_112,N_29806,N_29109);
and UO_113 (O_113,N_29211,N_29143);
nor UO_114 (O_114,N_29771,N_28971);
xnor UO_115 (O_115,N_29062,N_29128);
and UO_116 (O_116,N_29091,N_28879);
nor UO_117 (O_117,N_28998,N_29268);
nand UO_118 (O_118,N_28861,N_29730);
nor UO_119 (O_119,N_29607,N_29329);
or UO_120 (O_120,N_29412,N_29284);
and UO_121 (O_121,N_29100,N_29851);
and UO_122 (O_122,N_29196,N_29125);
and UO_123 (O_123,N_29117,N_29702);
and UO_124 (O_124,N_29905,N_29333);
and UO_125 (O_125,N_29610,N_29320);
nor UO_126 (O_126,N_28815,N_29596);
and UO_127 (O_127,N_28969,N_29050);
nand UO_128 (O_128,N_29808,N_29157);
xnor UO_129 (O_129,N_29616,N_29044);
xnor UO_130 (O_130,N_28940,N_29471);
or UO_131 (O_131,N_29110,N_29498);
nand UO_132 (O_132,N_29253,N_28852);
nor UO_133 (O_133,N_29190,N_29885);
and UO_134 (O_134,N_29848,N_29437);
and UO_135 (O_135,N_29899,N_29218);
xor UO_136 (O_136,N_29236,N_29643);
nor UO_137 (O_137,N_29034,N_29032);
nor UO_138 (O_138,N_29854,N_29398);
and UO_139 (O_139,N_29459,N_29759);
nor UO_140 (O_140,N_28891,N_29013);
nand UO_141 (O_141,N_29415,N_29309);
nor UO_142 (O_142,N_29508,N_29728);
nor UO_143 (O_143,N_29867,N_29331);
nor UO_144 (O_144,N_28962,N_29263);
or UO_145 (O_145,N_29202,N_29748);
nand UO_146 (O_146,N_29111,N_28881);
nand UO_147 (O_147,N_29718,N_29184);
nor UO_148 (O_148,N_29181,N_29703);
or UO_149 (O_149,N_29468,N_29765);
nand UO_150 (O_150,N_29602,N_28909);
xor UO_151 (O_151,N_29090,N_29781);
nor UO_152 (O_152,N_28939,N_29279);
and UO_153 (O_153,N_29146,N_29906);
and UO_154 (O_154,N_29927,N_28902);
and UO_155 (O_155,N_29475,N_29058);
xnor UO_156 (O_156,N_29142,N_29294);
nand UO_157 (O_157,N_28937,N_29881);
xnor UO_158 (O_158,N_29863,N_29235);
and UO_159 (O_159,N_29971,N_29326);
nand UO_160 (O_160,N_29617,N_29898);
and UO_161 (O_161,N_29552,N_28887);
or UO_162 (O_162,N_29576,N_29244);
xnor UO_163 (O_163,N_29723,N_29633);
or UO_164 (O_164,N_29297,N_29363);
xnor UO_165 (O_165,N_29489,N_29230);
and UO_166 (O_166,N_29555,N_29920);
and UO_167 (O_167,N_29843,N_29420);
and UO_168 (O_168,N_29457,N_29053);
xnor UO_169 (O_169,N_29937,N_29183);
and UO_170 (O_170,N_29837,N_29207);
xnor UO_171 (O_171,N_29697,N_29264);
or UO_172 (O_172,N_29046,N_29239);
xnor UO_173 (O_173,N_29708,N_28843);
and UO_174 (O_174,N_29932,N_29139);
xnor UO_175 (O_175,N_29663,N_29767);
nor UO_176 (O_176,N_29287,N_29689);
and UO_177 (O_177,N_28810,N_29594);
or UO_178 (O_178,N_29205,N_29929);
or UO_179 (O_179,N_29481,N_29908);
or UO_180 (O_180,N_29246,N_29373);
nor UO_181 (O_181,N_29208,N_29738);
nand UO_182 (O_182,N_29719,N_29160);
nand UO_183 (O_183,N_29223,N_28947);
and UO_184 (O_184,N_29068,N_29193);
nand UO_185 (O_185,N_29789,N_29548);
nor UO_186 (O_186,N_28831,N_29733);
nor UO_187 (O_187,N_29684,N_29303);
nand UO_188 (O_188,N_29687,N_28827);
or UO_189 (O_189,N_29773,N_29170);
nand UO_190 (O_190,N_28988,N_29332);
and UO_191 (O_191,N_28842,N_29416);
nand UO_192 (O_192,N_29176,N_29118);
and UO_193 (O_193,N_29300,N_29115);
nand UO_194 (O_194,N_29024,N_29483);
nand UO_195 (O_195,N_29769,N_28825);
and UO_196 (O_196,N_29661,N_29712);
or UO_197 (O_197,N_29753,N_29391);
or UO_198 (O_198,N_29878,N_29623);
xor UO_199 (O_199,N_29800,N_29477);
or UO_200 (O_200,N_29368,N_29574);
or UO_201 (O_201,N_29149,N_29856);
and UO_202 (O_202,N_29052,N_29827);
or UO_203 (O_203,N_29059,N_29677);
nor UO_204 (O_204,N_29116,N_28963);
nand UO_205 (O_205,N_29683,N_28829);
or UO_206 (O_206,N_29659,N_29254);
or UO_207 (O_207,N_29228,N_29638);
nand UO_208 (O_208,N_29523,N_29406);
or UO_209 (O_209,N_29563,N_29780);
or UO_210 (O_210,N_29519,N_29130);
nor UO_211 (O_211,N_29410,N_29811);
and UO_212 (O_212,N_29315,N_29954);
and UO_213 (O_213,N_29114,N_29538);
nor UO_214 (O_214,N_29094,N_29355);
nand UO_215 (O_215,N_29680,N_28958);
nor UO_216 (O_216,N_29872,N_28922);
nand UO_217 (O_217,N_29182,N_28833);
nor UO_218 (O_218,N_29956,N_29924);
nand UO_219 (O_219,N_29188,N_29405);
xor UO_220 (O_220,N_29278,N_29679);
or UO_221 (O_221,N_29987,N_29935);
nor UO_222 (O_222,N_28948,N_29995);
nor UO_223 (O_223,N_29894,N_29113);
nand UO_224 (O_224,N_29869,N_29942);
or UO_225 (O_225,N_29989,N_29283);
nor UO_226 (O_226,N_29600,N_28844);
nand UO_227 (O_227,N_29487,N_29380);
nand UO_228 (O_228,N_28989,N_29865);
nand UO_229 (O_229,N_29700,N_28932);
nand UO_230 (O_230,N_29641,N_28943);
nand UO_231 (O_231,N_29280,N_29322);
and UO_232 (O_232,N_29325,N_29941);
nand UO_233 (O_233,N_29018,N_29866);
nor UO_234 (O_234,N_29615,N_29686);
xor UO_235 (O_235,N_29274,N_29007);
nand UO_236 (O_236,N_28934,N_29582);
nand UO_237 (O_237,N_29969,N_29262);
nor UO_238 (O_238,N_29662,N_29249);
and UO_239 (O_239,N_29540,N_29536);
nand UO_240 (O_240,N_29096,N_29028);
xnor UO_241 (O_241,N_29148,N_29553);
nor UO_242 (O_242,N_29810,N_29004);
or UO_243 (O_243,N_29772,N_29624);
nand UO_244 (O_244,N_29649,N_29690);
nand UO_245 (O_245,N_29296,N_29622);
and UO_246 (O_246,N_29482,N_28923);
or UO_247 (O_247,N_29448,N_29469);
and UO_248 (O_248,N_29474,N_28873);
and UO_249 (O_249,N_29817,N_29016);
or UO_250 (O_250,N_29786,N_29835);
nand UO_251 (O_251,N_29704,N_29232);
nand UO_252 (O_252,N_29586,N_29880);
xnor UO_253 (O_253,N_29916,N_29785);
nand UO_254 (O_254,N_29913,N_29436);
xnor UO_255 (O_255,N_29820,N_29162);
and UO_256 (O_256,N_28978,N_29324);
nand UO_257 (O_257,N_29926,N_29430);
or UO_258 (O_258,N_29840,N_29884);
nor UO_259 (O_259,N_29860,N_29306);
xor UO_260 (O_260,N_29575,N_29545);
nand UO_261 (O_261,N_29731,N_29051);
and UO_262 (O_262,N_29403,N_29566);
nand UO_263 (O_263,N_29497,N_29356);
nand UO_264 (O_264,N_29621,N_28897);
and UO_265 (O_265,N_29227,N_28950);
nor UO_266 (O_266,N_29165,N_29818);
and UO_267 (O_267,N_29241,N_29983);
nand UO_268 (O_268,N_29914,N_28935);
or UO_269 (O_269,N_29669,N_29431);
nand UO_270 (O_270,N_29931,N_28851);
xnor UO_271 (O_271,N_29985,N_29727);
nor UO_272 (O_272,N_29522,N_29348);
and UO_273 (O_273,N_29075,N_28821);
or UO_274 (O_274,N_29385,N_29897);
nand UO_275 (O_275,N_29701,N_29614);
and UO_276 (O_276,N_29413,N_29945);
nand UO_277 (O_277,N_29328,N_29783);
nor UO_278 (O_278,N_29175,N_29336);
and UO_279 (O_279,N_29131,N_29017);
and UO_280 (O_280,N_28979,N_29544);
and UO_281 (O_281,N_29503,N_29625);
nor UO_282 (O_282,N_29829,N_28864);
nor UO_283 (O_283,N_29337,N_29883);
or UO_284 (O_284,N_29397,N_29518);
nor UO_285 (O_285,N_28868,N_29573);
and UO_286 (O_286,N_29952,N_28899);
xnor UO_287 (O_287,N_29072,N_29516);
nand UO_288 (O_288,N_29637,N_29305);
xor UO_289 (O_289,N_29960,N_29763);
nor UO_290 (O_290,N_29045,N_29271);
and UO_291 (O_291,N_29238,N_29535);
and UO_292 (O_292,N_29502,N_29630);
or UO_293 (O_293,N_29709,N_29351);
xor UO_294 (O_294,N_29340,N_29495);
and UO_295 (O_295,N_29838,N_29458);
and UO_296 (O_296,N_29001,N_29079);
nor UO_297 (O_297,N_29316,N_29361);
xnor UO_298 (O_298,N_29543,N_29980);
nor UO_299 (O_299,N_29377,N_29961);
and UO_300 (O_300,N_29673,N_29938);
xor UO_301 (O_301,N_29845,N_29439);
or UO_302 (O_302,N_29766,N_29376);
nor UO_303 (O_303,N_28931,N_29667);
and UO_304 (O_304,N_28910,N_29722);
nand UO_305 (O_305,N_28872,N_29120);
and UO_306 (O_306,N_29360,N_29512);
or UO_307 (O_307,N_29452,N_28995);
xnor UO_308 (O_308,N_29014,N_29450);
or UO_309 (O_309,N_29156,N_29876);
or UO_310 (O_310,N_29842,N_29949);
xor UO_311 (O_311,N_29461,N_29572);
nand UO_312 (O_312,N_29456,N_29978);
nor UO_313 (O_313,N_29212,N_29145);
nand UO_314 (O_314,N_28870,N_29237);
or UO_315 (O_315,N_28862,N_29022);
and UO_316 (O_316,N_29747,N_28996);
or UO_317 (O_317,N_28993,N_29634);
nor UO_318 (O_318,N_29019,N_29220);
or UO_319 (O_319,N_29387,N_29349);
nand UO_320 (O_320,N_29069,N_29442);
xnor UO_321 (O_321,N_29597,N_29915);
nor UO_322 (O_322,N_29446,N_29493);
and UO_323 (O_323,N_29060,N_29647);
and UO_324 (O_324,N_29830,N_28884);
or UO_325 (O_325,N_29318,N_29171);
nand UO_326 (O_326,N_28941,N_29386);
nand UO_327 (O_327,N_28837,N_28882);
or UO_328 (O_328,N_29912,N_29476);
or UO_329 (O_329,N_28820,N_29026);
or UO_330 (O_330,N_28928,N_29740);
nand UO_331 (O_331,N_29520,N_29788);
or UO_332 (O_332,N_29399,N_29108);
or UO_333 (O_333,N_28925,N_28826);
xnor UO_334 (O_334,N_29168,N_29882);
nand UO_335 (O_335,N_28866,N_29591);
nand UO_336 (O_336,N_29401,N_29112);
nand UO_337 (O_337,N_29976,N_28956);
nand UO_338 (O_338,N_29651,N_29939);
and UO_339 (O_339,N_28982,N_29642);
or UO_340 (O_340,N_28814,N_28967);
nand UO_341 (O_341,N_29067,N_29584);
nand UO_342 (O_342,N_29565,N_28957);
or UO_343 (O_343,N_29344,N_29592);
nor UO_344 (O_344,N_29164,N_29658);
nor UO_345 (O_345,N_29934,N_29608);
xnor UO_346 (O_346,N_29345,N_29585);
or UO_347 (O_347,N_29233,N_29970);
nor UO_348 (O_348,N_29674,N_29813);
nand UO_349 (O_349,N_29628,N_29445);
or UO_350 (O_350,N_29252,N_29737);
nand UO_351 (O_351,N_28966,N_29242);
nor UO_352 (O_352,N_29295,N_28968);
or UO_353 (O_353,N_29857,N_29392);
or UO_354 (O_354,N_28901,N_29790);
xnor UO_355 (O_355,N_28936,N_28840);
and UO_356 (O_356,N_28811,N_29463);
or UO_357 (O_357,N_28803,N_29402);
and UO_358 (O_358,N_29243,N_29037);
xnor UO_359 (O_359,N_29369,N_29743);
xnor UO_360 (O_360,N_29441,N_29874);
and UO_361 (O_361,N_29782,N_29214);
and UO_362 (O_362,N_29870,N_29438);
and UO_363 (O_363,N_29105,N_29308);
nor UO_364 (O_364,N_29159,N_29152);
nor UO_365 (O_365,N_29354,N_29825);
xnor UO_366 (O_366,N_29101,N_29008);
or UO_367 (O_367,N_29672,N_28933);
nor UO_368 (O_368,N_29685,N_29462);
nor UO_369 (O_369,N_29735,N_29185);
and UO_370 (O_370,N_29928,N_29124);
or UO_371 (O_371,N_29041,N_29770);
xnor UO_372 (O_372,N_29103,N_29085);
or UO_373 (O_373,N_29460,N_29524);
nand UO_374 (O_374,N_29421,N_29266);
nor UO_375 (O_375,N_29562,N_29107);
and UO_376 (O_376,N_29595,N_29210);
and UO_377 (O_377,N_29525,N_29706);
xor UO_378 (O_378,N_29824,N_29605);
or UO_379 (O_379,N_29779,N_29694);
or UO_380 (O_380,N_29580,N_29528);
nand UO_381 (O_381,N_29106,N_29809);
xor UO_382 (O_382,N_29064,N_29569);
nor UO_383 (O_383,N_29795,N_29846);
xnor UO_384 (O_384,N_28930,N_29646);
and UO_385 (O_385,N_29167,N_29589);
and UO_386 (O_386,N_29258,N_29819);
nand UO_387 (O_387,N_29093,N_29907);
and UO_388 (O_388,N_29327,N_29470);
or UO_389 (O_389,N_29343,N_29098);
and UO_390 (O_390,N_29601,N_29892);
xor UO_391 (O_391,N_29323,N_29895);
and UO_392 (O_392,N_29670,N_29812);
or UO_393 (O_393,N_28908,N_29381);
nor UO_394 (O_394,N_29705,N_29997);
and UO_395 (O_395,N_28849,N_28942);
and UO_396 (O_396,N_29861,N_29259);
and UO_397 (O_397,N_28916,N_29711);
nor UO_398 (O_398,N_29191,N_29505);
nor UO_399 (O_399,N_29578,N_29134);
nor UO_400 (O_400,N_29395,N_29862);
or UO_401 (O_401,N_29169,N_29635);
or UO_402 (O_402,N_29691,N_29515);
nor UO_403 (O_403,N_28834,N_29921);
and UO_404 (O_404,N_29158,N_29752);
nand UO_405 (O_405,N_28973,N_29629);
or UO_406 (O_406,N_29500,N_29358);
nand UO_407 (O_407,N_29427,N_29129);
xnor UO_408 (O_408,N_29078,N_29247);
xnor UO_409 (O_409,N_29962,N_29293);
and UO_410 (O_410,N_29074,N_29285);
xnor UO_411 (O_411,N_29491,N_28892);
xnor UO_412 (O_412,N_29999,N_29453);
and UO_413 (O_413,N_28816,N_29286);
xor UO_414 (O_414,N_28976,N_29076);
and UO_415 (O_415,N_29721,N_29301);
or UO_416 (O_416,N_29341,N_29424);
and UO_417 (O_417,N_29732,N_29119);
xnor UO_418 (O_418,N_29796,N_28984);
or UO_419 (O_419,N_29166,N_28954);
and UO_420 (O_420,N_29219,N_28808);
nand UO_421 (O_421,N_29137,N_29099);
and UO_422 (O_422,N_29768,N_28893);
and UO_423 (O_423,N_29858,N_28927);
nor UO_424 (O_424,N_29556,N_29981);
or UO_425 (O_425,N_29390,N_29955);
xor UO_426 (O_426,N_29725,N_29359);
or UO_427 (O_427,N_29903,N_29599);
or UO_428 (O_428,N_28857,N_28994);
or UO_429 (O_429,N_29135,N_29389);
xnor UO_430 (O_430,N_29984,N_28917);
nand UO_431 (O_431,N_29240,N_28845);
xnor UO_432 (O_432,N_29087,N_29371);
nand UO_433 (O_433,N_29488,N_29027);
or UO_434 (O_434,N_29664,N_29290);
and UO_435 (O_435,N_29133,N_29267);
and UO_436 (O_436,N_29396,N_29852);
xnor UO_437 (O_437,N_29307,N_29049);
and UO_438 (O_438,N_28914,N_29760);
nor UO_439 (O_439,N_29009,N_28848);
nor UO_440 (O_440,N_29991,N_29222);
xor UO_441 (O_441,N_29272,N_29221);
and UO_442 (O_442,N_29065,N_29204);
and UO_443 (O_443,N_29198,N_29698);
nand UO_444 (O_444,N_29189,N_29350);
and UO_445 (O_445,N_29784,N_29417);
xnor UO_446 (O_446,N_29186,N_28915);
nand UO_447 (O_447,N_29418,N_29261);
or UO_448 (O_448,N_29804,N_29364);
nor UO_449 (O_449,N_29038,N_28992);
and UO_450 (O_450,N_29816,N_29724);
nand UO_451 (O_451,N_29444,N_29648);
nand UO_452 (O_452,N_29803,N_29040);
or UO_453 (O_453,N_29464,N_29758);
and UO_454 (O_454,N_29947,N_29940);
xor UO_455 (O_455,N_28839,N_28819);
nor UO_456 (O_456,N_29910,N_29521);
and UO_457 (O_457,N_29558,N_29229);
or UO_458 (O_458,N_29353,N_29668);
or UO_459 (O_459,N_29346,N_28805);
xor UO_460 (O_460,N_29352,N_29750);
or UO_461 (O_461,N_29590,N_29762);
nor UO_462 (O_462,N_28926,N_29126);
xnor UO_463 (O_463,N_29655,N_29310);
or UO_464 (O_464,N_29404,N_29998);
xnor UO_465 (O_465,N_29968,N_28853);
and UO_466 (O_466,N_29151,N_29375);
or UO_467 (O_467,N_28865,N_29653);
nand UO_468 (O_468,N_29177,N_29000);
nor UO_469 (O_469,N_29948,N_29844);
nand UO_470 (O_470,N_29577,N_29688);
and UO_471 (O_471,N_28907,N_29542);
nor UO_472 (O_472,N_29339,N_29084);
or UO_473 (O_473,N_29209,N_28830);
and UO_474 (O_474,N_29990,N_29187);
xor UO_475 (O_475,N_29693,N_29506);
xor UO_476 (O_476,N_29644,N_29088);
or UO_477 (O_477,N_29312,N_28804);
xor UO_478 (O_478,N_29031,N_28886);
nand UO_479 (O_479,N_28944,N_29435);
and UO_480 (O_480,N_29288,N_29911);
nor UO_481 (O_481,N_29925,N_29965);
nor UO_482 (O_482,N_29666,N_29490);
xor UO_483 (O_483,N_28802,N_29755);
nand UO_484 (O_484,N_29710,N_29042);
nor UO_485 (O_485,N_28824,N_29761);
and UO_486 (O_486,N_29510,N_29776);
nand UO_487 (O_487,N_29260,N_29020);
or UO_488 (O_488,N_29023,N_29273);
xnor UO_489 (O_489,N_29003,N_29492);
nand UO_490 (O_490,N_29918,N_29372);
or UO_491 (O_491,N_29172,N_29338);
nor UO_492 (O_492,N_28817,N_29871);
or UO_493 (O_493,N_29833,N_29529);
and UO_494 (O_494,N_29393,N_29025);
xor UO_495 (O_495,N_29055,N_29917);
and UO_496 (O_496,N_29665,N_28900);
or UO_497 (O_497,N_29063,N_29606);
nor UO_498 (O_498,N_29879,N_29933);
xnor UO_499 (O_499,N_29292,N_28904);
and UO_500 (O_500,N_29311,N_29467);
and UO_501 (O_501,N_29603,N_29141);
nand UO_502 (O_502,N_29756,N_29342);
and UO_503 (O_503,N_29936,N_29383);
xnor UO_504 (O_504,N_29407,N_29378);
and UO_505 (O_505,N_28929,N_29967);
nor UO_506 (O_506,N_28828,N_28977);
xor UO_507 (O_507,N_29511,N_29850);
or UO_508 (O_508,N_28809,N_29631);
xnor UO_509 (O_509,N_29944,N_29775);
nor UO_510 (O_510,N_29749,N_29919);
nor UO_511 (O_511,N_28959,N_28850);
or UO_512 (O_512,N_29714,N_29006);
or UO_513 (O_513,N_29992,N_28801);
nor UO_514 (O_514,N_29930,N_29561);
xor UO_515 (O_515,N_29366,N_28918);
xor UO_516 (O_516,N_29979,N_29805);
and UO_517 (O_517,N_29922,N_28823);
or UO_518 (O_518,N_29657,N_29357);
or UO_519 (O_519,N_29231,N_29299);
xor UO_520 (O_520,N_29277,N_29636);
or UO_521 (O_521,N_29379,N_29550);
or UO_522 (O_522,N_29604,N_29537);
nor UO_523 (O_523,N_29593,N_29201);
or UO_524 (O_524,N_29950,N_29217);
nor UO_525 (O_525,N_29654,N_28972);
and UO_526 (O_526,N_29071,N_29155);
nor UO_527 (O_527,N_28871,N_29140);
nor UO_528 (O_528,N_29859,N_29426);
nor UO_529 (O_529,N_29889,N_29454);
and UO_530 (O_530,N_28952,N_29541);
nand UO_531 (O_531,N_29793,N_29433);
and UO_532 (O_532,N_28986,N_29192);
nor UO_533 (O_533,N_29144,N_29197);
nand UO_534 (O_534,N_29480,N_28890);
nand UO_535 (O_535,N_28905,N_29256);
nor UO_536 (O_536,N_29314,N_28981);
nor UO_537 (O_537,N_29215,N_29030);
xnor UO_538 (O_538,N_29900,N_29216);
and UO_539 (O_539,N_29449,N_29660);
nor UO_540 (O_540,N_29289,N_28903);
xnor UO_541 (O_541,N_29425,N_29432);
or UO_542 (O_542,N_28898,N_28880);
nand UO_543 (O_543,N_29347,N_29472);
nand UO_544 (O_544,N_29021,N_29957);
nand UO_545 (O_545,N_29640,N_29618);
and UO_546 (O_546,N_29195,N_29656);
nand UO_547 (O_547,N_28912,N_29836);
nor UO_548 (O_548,N_29675,N_29994);
nor UO_549 (O_549,N_29513,N_28961);
nor UO_550 (O_550,N_29736,N_28807);
and UO_551 (O_551,N_29517,N_29864);
xnor UO_552 (O_552,N_29250,N_29012);
xor UO_553 (O_553,N_29161,N_29564);
nand UO_554 (O_554,N_29121,N_28869);
nand UO_555 (O_555,N_29015,N_29056);
xnor UO_556 (O_556,N_29248,N_29367);
xor UO_557 (O_557,N_29717,N_29547);
nand UO_558 (O_558,N_28874,N_29138);
or UO_559 (O_559,N_29200,N_29179);
and UO_560 (O_560,N_29791,N_29434);
or UO_561 (O_561,N_29681,N_29039);
xor UO_562 (O_562,N_29742,N_29739);
nor UO_563 (O_563,N_28951,N_29671);
xor UO_564 (O_564,N_28953,N_29255);
nand UO_565 (O_565,N_29479,N_29551);
nor UO_566 (O_566,N_29465,N_29533);
xnor UO_567 (O_567,N_29213,N_28921);
nand UO_568 (O_568,N_29070,N_28835);
xnor UO_569 (O_569,N_28955,N_29104);
nor UO_570 (O_570,N_29557,N_28945);
or UO_571 (O_571,N_28854,N_28832);
nand UO_572 (O_572,N_29986,N_29588);
and UO_573 (O_573,N_29579,N_28974);
xor UO_574 (O_574,N_28813,N_29801);
xnor UO_575 (O_575,N_29319,N_29609);
and UO_576 (O_576,N_29496,N_28818);
and UO_577 (O_577,N_29269,N_29792);
xor UO_578 (O_578,N_29778,N_29122);
or UO_579 (O_579,N_29499,N_29153);
nor UO_580 (O_580,N_29473,N_28896);
xor UO_581 (O_581,N_29799,N_29086);
xor UO_582 (O_582,N_29317,N_29716);
xnor UO_583 (O_583,N_29411,N_29549);
or UO_584 (O_584,N_28841,N_29539);
xor UO_585 (O_585,N_29839,N_29988);
and UO_586 (O_586,N_28960,N_29409);
and UO_587 (O_587,N_28856,N_29875);
and UO_588 (O_588,N_29154,N_29073);
nor UO_589 (O_589,N_28983,N_29699);
nor UO_590 (O_590,N_29275,N_29321);
xor UO_591 (O_591,N_28895,N_29993);
xnor UO_592 (O_592,N_29975,N_29888);
nand UO_593 (O_593,N_28883,N_29150);
xor UO_594 (O_594,N_29923,N_29807);
or UO_595 (O_595,N_29428,N_29061);
xnor UO_596 (O_596,N_29977,N_29527);
or UO_597 (O_597,N_29554,N_29963);
or UO_598 (O_598,N_29313,N_29726);
and UO_599 (O_599,N_29501,N_29696);
nor UO_600 (O_600,N_29701,N_29527);
and UO_601 (O_601,N_28817,N_29558);
nor UO_602 (O_602,N_29614,N_29199);
nor UO_603 (O_603,N_29070,N_28825);
nand UO_604 (O_604,N_29989,N_29616);
and UO_605 (O_605,N_29556,N_29630);
and UO_606 (O_606,N_29499,N_29995);
or UO_607 (O_607,N_29392,N_28826);
or UO_608 (O_608,N_28895,N_28828);
nand UO_609 (O_609,N_28843,N_29627);
and UO_610 (O_610,N_29151,N_29146);
or UO_611 (O_611,N_28801,N_29407);
or UO_612 (O_612,N_29732,N_29454);
and UO_613 (O_613,N_29047,N_29316);
xor UO_614 (O_614,N_29369,N_29572);
or UO_615 (O_615,N_29919,N_29351);
xor UO_616 (O_616,N_29349,N_29275);
nor UO_617 (O_617,N_28887,N_29040);
and UO_618 (O_618,N_29991,N_29746);
or UO_619 (O_619,N_28964,N_29738);
xnor UO_620 (O_620,N_28812,N_29608);
and UO_621 (O_621,N_29909,N_29258);
xor UO_622 (O_622,N_28882,N_29803);
and UO_623 (O_623,N_29157,N_29190);
nor UO_624 (O_624,N_29043,N_29963);
nand UO_625 (O_625,N_29019,N_29267);
or UO_626 (O_626,N_29741,N_29163);
xor UO_627 (O_627,N_29518,N_29958);
or UO_628 (O_628,N_29344,N_29101);
nor UO_629 (O_629,N_29932,N_28879);
and UO_630 (O_630,N_29849,N_29297);
or UO_631 (O_631,N_29999,N_29920);
and UO_632 (O_632,N_29292,N_29596);
nor UO_633 (O_633,N_28857,N_29499);
xor UO_634 (O_634,N_28875,N_29808);
nor UO_635 (O_635,N_29933,N_29877);
nor UO_636 (O_636,N_29728,N_29898);
and UO_637 (O_637,N_29132,N_29723);
nand UO_638 (O_638,N_29670,N_29210);
and UO_639 (O_639,N_29678,N_29540);
nand UO_640 (O_640,N_29742,N_29230);
or UO_641 (O_641,N_29393,N_28857);
nor UO_642 (O_642,N_29797,N_29439);
and UO_643 (O_643,N_29745,N_29068);
xnor UO_644 (O_644,N_28800,N_29631);
or UO_645 (O_645,N_29216,N_29249);
and UO_646 (O_646,N_29556,N_29860);
nand UO_647 (O_647,N_29829,N_29241);
and UO_648 (O_648,N_28971,N_29409);
or UO_649 (O_649,N_29914,N_29150);
or UO_650 (O_650,N_29119,N_28907);
or UO_651 (O_651,N_29326,N_29989);
xnor UO_652 (O_652,N_29101,N_28908);
and UO_653 (O_653,N_29604,N_29961);
nor UO_654 (O_654,N_29065,N_29246);
xnor UO_655 (O_655,N_29067,N_29437);
and UO_656 (O_656,N_29462,N_29246);
nand UO_657 (O_657,N_29945,N_29414);
nor UO_658 (O_658,N_29686,N_28905);
and UO_659 (O_659,N_29282,N_29442);
or UO_660 (O_660,N_29287,N_28853);
or UO_661 (O_661,N_29611,N_29008);
or UO_662 (O_662,N_28968,N_29276);
nand UO_663 (O_663,N_29636,N_29040);
or UO_664 (O_664,N_29611,N_28926);
or UO_665 (O_665,N_29512,N_29169);
and UO_666 (O_666,N_28802,N_29318);
xor UO_667 (O_667,N_29047,N_29084);
xnor UO_668 (O_668,N_28939,N_28988);
nor UO_669 (O_669,N_29134,N_29815);
or UO_670 (O_670,N_29496,N_29647);
and UO_671 (O_671,N_29877,N_29111);
nand UO_672 (O_672,N_29517,N_29073);
xnor UO_673 (O_673,N_29129,N_29957);
nand UO_674 (O_674,N_29032,N_29076);
and UO_675 (O_675,N_29036,N_28972);
and UO_676 (O_676,N_29046,N_29637);
and UO_677 (O_677,N_29838,N_29017);
and UO_678 (O_678,N_29312,N_29360);
or UO_679 (O_679,N_29404,N_29776);
nor UO_680 (O_680,N_29151,N_29603);
nor UO_681 (O_681,N_29438,N_29901);
nand UO_682 (O_682,N_29560,N_29092);
xnor UO_683 (O_683,N_29550,N_29131);
xor UO_684 (O_684,N_28970,N_29496);
xor UO_685 (O_685,N_29383,N_29870);
or UO_686 (O_686,N_28841,N_28800);
nand UO_687 (O_687,N_29776,N_29018);
nand UO_688 (O_688,N_29668,N_29197);
and UO_689 (O_689,N_29259,N_28962);
xnor UO_690 (O_690,N_28808,N_29152);
nor UO_691 (O_691,N_29373,N_29064);
xnor UO_692 (O_692,N_29443,N_28940);
xor UO_693 (O_693,N_29547,N_29886);
xnor UO_694 (O_694,N_29420,N_28813);
nand UO_695 (O_695,N_28971,N_29378);
xor UO_696 (O_696,N_29258,N_29665);
nor UO_697 (O_697,N_29228,N_29557);
or UO_698 (O_698,N_29181,N_28869);
xnor UO_699 (O_699,N_28949,N_29408);
or UO_700 (O_700,N_29709,N_29242);
and UO_701 (O_701,N_29729,N_29273);
xnor UO_702 (O_702,N_29137,N_29229);
nand UO_703 (O_703,N_29151,N_29824);
xnor UO_704 (O_704,N_28950,N_28980);
and UO_705 (O_705,N_29950,N_29045);
xnor UO_706 (O_706,N_29049,N_29487);
and UO_707 (O_707,N_28847,N_29673);
nand UO_708 (O_708,N_29312,N_29796);
nand UO_709 (O_709,N_29215,N_29641);
xnor UO_710 (O_710,N_28907,N_29203);
nor UO_711 (O_711,N_29204,N_29802);
xnor UO_712 (O_712,N_29137,N_29711);
or UO_713 (O_713,N_29980,N_29413);
nor UO_714 (O_714,N_29104,N_29000);
and UO_715 (O_715,N_29816,N_29760);
nor UO_716 (O_716,N_29283,N_29655);
nand UO_717 (O_717,N_28903,N_29366);
or UO_718 (O_718,N_29832,N_29062);
xor UO_719 (O_719,N_29952,N_29015);
xnor UO_720 (O_720,N_29841,N_29893);
or UO_721 (O_721,N_28892,N_29196);
and UO_722 (O_722,N_29261,N_29175);
nor UO_723 (O_723,N_29396,N_29528);
nor UO_724 (O_724,N_29138,N_29101);
nor UO_725 (O_725,N_29973,N_29600);
and UO_726 (O_726,N_28878,N_29721);
nand UO_727 (O_727,N_29244,N_29686);
nand UO_728 (O_728,N_29880,N_28810);
nand UO_729 (O_729,N_28937,N_29751);
and UO_730 (O_730,N_29666,N_29616);
or UO_731 (O_731,N_29349,N_29057);
and UO_732 (O_732,N_29282,N_29656);
or UO_733 (O_733,N_29384,N_28884);
and UO_734 (O_734,N_29785,N_29519);
nor UO_735 (O_735,N_29721,N_29268);
nand UO_736 (O_736,N_29850,N_29545);
and UO_737 (O_737,N_29261,N_29139);
xor UO_738 (O_738,N_28842,N_29440);
and UO_739 (O_739,N_28886,N_29338);
nor UO_740 (O_740,N_29193,N_29419);
xnor UO_741 (O_741,N_29454,N_29497);
nor UO_742 (O_742,N_29357,N_29730);
nand UO_743 (O_743,N_29380,N_29038);
and UO_744 (O_744,N_29934,N_29666);
or UO_745 (O_745,N_28856,N_29534);
and UO_746 (O_746,N_29817,N_29799);
nand UO_747 (O_747,N_29374,N_29582);
nand UO_748 (O_748,N_29947,N_29662);
xnor UO_749 (O_749,N_28878,N_29193);
and UO_750 (O_750,N_29239,N_28866);
and UO_751 (O_751,N_29207,N_29660);
nand UO_752 (O_752,N_29689,N_29547);
and UO_753 (O_753,N_29098,N_29353);
nand UO_754 (O_754,N_29611,N_29851);
xnor UO_755 (O_755,N_29555,N_29185);
xor UO_756 (O_756,N_29789,N_28810);
xnor UO_757 (O_757,N_28905,N_28953);
nand UO_758 (O_758,N_29708,N_29699);
or UO_759 (O_759,N_29466,N_28903);
xnor UO_760 (O_760,N_29315,N_29336);
and UO_761 (O_761,N_29294,N_29090);
or UO_762 (O_762,N_28967,N_29541);
or UO_763 (O_763,N_29521,N_29050);
and UO_764 (O_764,N_29704,N_29116);
and UO_765 (O_765,N_29713,N_29217);
nand UO_766 (O_766,N_28878,N_29753);
and UO_767 (O_767,N_29858,N_29103);
or UO_768 (O_768,N_29232,N_29822);
or UO_769 (O_769,N_29840,N_29798);
or UO_770 (O_770,N_29491,N_29278);
nand UO_771 (O_771,N_29552,N_29789);
xnor UO_772 (O_772,N_28820,N_29217);
nor UO_773 (O_773,N_29673,N_29552);
or UO_774 (O_774,N_29254,N_29302);
and UO_775 (O_775,N_29506,N_29106);
and UO_776 (O_776,N_29923,N_29005);
and UO_777 (O_777,N_29828,N_29937);
xor UO_778 (O_778,N_29592,N_29342);
nor UO_779 (O_779,N_29312,N_28898);
nor UO_780 (O_780,N_29368,N_29742);
nand UO_781 (O_781,N_29237,N_29265);
nand UO_782 (O_782,N_28875,N_29268);
nand UO_783 (O_783,N_28905,N_28896);
and UO_784 (O_784,N_29996,N_29062);
or UO_785 (O_785,N_29452,N_29588);
xnor UO_786 (O_786,N_29220,N_29512);
or UO_787 (O_787,N_29347,N_29078);
nor UO_788 (O_788,N_29560,N_28957);
xnor UO_789 (O_789,N_28919,N_28909);
or UO_790 (O_790,N_29661,N_29268);
nor UO_791 (O_791,N_29703,N_29478);
nor UO_792 (O_792,N_29581,N_29303);
nor UO_793 (O_793,N_29250,N_29519);
nand UO_794 (O_794,N_29099,N_29035);
and UO_795 (O_795,N_29403,N_29367);
xor UO_796 (O_796,N_28969,N_29011);
nand UO_797 (O_797,N_29493,N_29841);
or UO_798 (O_798,N_29999,N_29175);
xor UO_799 (O_799,N_29406,N_28863);
and UO_800 (O_800,N_29640,N_29328);
xor UO_801 (O_801,N_29494,N_29468);
nor UO_802 (O_802,N_29626,N_29465);
or UO_803 (O_803,N_29134,N_29897);
or UO_804 (O_804,N_29643,N_29696);
nor UO_805 (O_805,N_29812,N_29399);
nor UO_806 (O_806,N_29977,N_29031);
or UO_807 (O_807,N_29311,N_29972);
xnor UO_808 (O_808,N_29917,N_29565);
xor UO_809 (O_809,N_29954,N_28946);
xor UO_810 (O_810,N_29805,N_29062);
and UO_811 (O_811,N_29132,N_29948);
xor UO_812 (O_812,N_29113,N_29849);
nor UO_813 (O_813,N_29256,N_29012);
or UO_814 (O_814,N_28928,N_29645);
nor UO_815 (O_815,N_29356,N_29477);
nand UO_816 (O_816,N_29349,N_29127);
and UO_817 (O_817,N_29822,N_29292);
and UO_818 (O_818,N_29330,N_29680);
and UO_819 (O_819,N_29099,N_29613);
or UO_820 (O_820,N_29604,N_28947);
and UO_821 (O_821,N_28953,N_29038);
xnor UO_822 (O_822,N_29504,N_29438);
nand UO_823 (O_823,N_29149,N_29219);
or UO_824 (O_824,N_29836,N_28986);
and UO_825 (O_825,N_28850,N_28839);
nor UO_826 (O_826,N_29412,N_28984);
nor UO_827 (O_827,N_29409,N_29815);
nand UO_828 (O_828,N_29825,N_29358);
or UO_829 (O_829,N_29467,N_28895);
or UO_830 (O_830,N_29473,N_29344);
xnor UO_831 (O_831,N_29519,N_29415);
nor UO_832 (O_832,N_29489,N_29971);
xor UO_833 (O_833,N_29990,N_29310);
and UO_834 (O_834,N_29994,N_29349);
xnor UO_835 (O_835,N_29737,N_29136);
or UO_836 (O_836,N_28965,N_29743);
or UO_837 (O_837,N_29930,N_29802);
or UO_838 (O_838,N_29224,N_28931);
or UO_839 (O_839,N_29511,N_29800);
and UO_840 (O_840,N_29499,N_28809);
xnor UO_841 (O_841,N_29371,N_29661);
and UO_842 (O_842,N_29245,N_29850);
and UO_843 (O_843,N_29665,N_29129);
nor UO_844 (O_844,N_29712,N_29553);
and UO_845 (O_845,N_29931,N_29541);
nor UO_846 (O_846,N_29657,N_29773);
nor UO_847 (O_847,N_29651,N_29620);
and UO_848 (O_848,N_29980,N_29120);
xnor UO_849 (O_849,N_28948,N_29867);
and UO_850 (O_850,N_29396,N_29957);
nor UO_851 (O_851,N_29080,N_29289);
or UO_852 (O_852,N_29581,N_29583);
and UO_853 (O_853,N_29393,N_29724);
nor UO_854 (O_854,N_29686,N_29894);
and UO_855 (O_855,N_29629,N_29981);
nand UO_856 (O_856,N_29812,N_28856);
nor UO_857 (O_857,N_29330,N_29458);
nand UO_858 (O_858,N_29694,N_29696);
nor UO_859 (O_859,N_29073,N_29661);
or UO_860 (O_860,N_29111,N_29589);
nor UO_861 (O_861,N_28942,N_29064);
and UO_862 (O_862,N_29581,N_29148);
or UO_863 (O_863,N_29188,N_29010);
or UO_864 (O_864,N_29146,N_29073);
or UO_865 (O_865,N_29924,N_29543);
nor UO_866 (O_866,N_29869,N_29652);
and UO_867 (O_867,N_29271,N_29605);
nand UO_868 (O_868,N_28930,N_28997);
or UO_869 (O_869,N_29490,N_29870);
nor UO_870 (O_870,N_29025,N_29178);
nand UO_871 (O_871,N_29478,N_29160);
xnor UO_872 (O_872,N_29281,N_29068);
or UO_873 (O_873,N_29184,N_28888);
nor UO_874 (O_874,N_29937,N_29565);
nand UO_875 (O_875,N_29353,N_29956);
nor UO_876 (O_876,N_29906,N_29371);
and UO_877 (O_877,N_29417,N_29650);
nor UO_878 (O_878,N_29824,N_29342);
xnor UO_879 (O_879,N_29611,N_29869);
nor UO_880 (O_880,N_29580,N_29345);
nor UO_881 (O_881,N_29993,N_29329);
or UO_882 (O_882,N_29526,N_29122);
nand UO_883 (O_883,N_29542,N_29792);
xor UO_884 (O_884,N_29547,N_28938);
and UO_885 (O_885,N_29199,N_29800);
and UO_886 (O_886,N_29995,N_29860);
nand UO_887 (O_887,N_29273,N_28892);
nand UO_888 (O_888,N_29818,N_28883);
nor UO_889 (O_889,N_28944,N_29465);
nor UO_890 (O_890,N_29418,N_29431);
nand UO_891 (O_891,N_29132,N_28906);
or UO_892 (O_892,N_29951,N_29409);
nand UO_893 (O_893,N_29822,N_28866);
xnor UO_894 (O_894,N_29633,N_28906);
nand UO_895 (O_895,N_28920,N_29280);
nor UO_896 (O_896,N_29879,N_29387);
or UO_897 (O_897,N_29283,N_29203);
and UO_898 (O_898,N_29625,N_29449);
and UO_899 (O_899,N_28980,N_29581);
or UO_900 (O_900,N_29536,N_29313);
nor UO_901 (O_901,N_29620,N_28987);
nand UO_902 (O_902,N_28872,N_29790);
or UO_903 (O_903,N_29145,N_29122);
xor UO_904 (O_904,N_29984,N_29961);
and UO_905 (O_905,N_28823,N_29189);
xnor UO_906 (O_906,N_29345,N_29055);
nand UO_907 (O_907,N_29316,N_28809);
xnor UO_908 (O_908,N_29534,N_29223);
xnor UO_909 (O_909,N_29058,N_28917);
xor UO_910 (O_910,N_29942,N_29288);
or UO_911 (O_911,N_29171,N_29529);
nand UO_912 (O_912,N_29271,N_28928);
nand UO_913 (O_913,N_29300,N_29634);
or UO_914 (O_914,N_29709,N_29649);
or UO_915 (O_915,N_29294,N_29840);
and UO_916 (O_916,N_29630,N_29453);
nand UO_917 (O_917,N_29416,N_29979);
xor UO_918 (O_918,N_29838,N_29524);
and UO_919 (O_919,N_29331,N_28819);
and UO_920 (O_920,N_29465,N_29028);
and UO_921 (O_921,N_29412,N_29726);
nor UO_922 (O_922,N_29119,N_29944);
and UO_923 (O_923,N_29058,N_29523);
and UO_924 (O_924,N_29672,N_29015);
nand UO_925 (O_925,N_29785,N_29823);
xor UO_926 (O_926,N_29484,N_29994);
nand UO_927 (O_927,N_29158,N_29465);
nor UO_928 (O_928,N_29894,N_28940);
or UO_929 (O_929,N_28977,N_29827);
nor UO_930 (O_930,N_29448,N_28920);
nand UO_931 (O_931,N_28979,N_29838);
or UO_932 (O_932,N_29378,N_29405);
xnor UO_933 (O_933,N_28977,N_29624);
and UO_934 (O_934,N_29884,N_29489);
nand UO_935 (O_935,N_29601,N_29835);
or UO_936 (O_936,N_29333,N_29236);
or UO_937 (O_937,N_29252,N_28801);
xnor UO_938 (O_938,N_29457,N_28911);
nor UO_939 (O_939,N_29996,N_29138);
or UO_940 (O_940,N_28883,N_28806);
or UO_941 (O_941,N_29643,N_29795);
or UO_942 (O_942,N_29861,N_29828);
and UO_943 (O_943,N_29229,N_29388);
xnor UO_944 (O_944,N_29508,N_29399);
and UO_945 (O_945,N_29969,N_29832);
and UO_946 (O_946,N_29413,N_29910);
nand UO_947 (O_947,N_29359,N_28818);
xnor UO_948 (O_948,N_28834,N_29665);
xor UO_949 (O_949,N_29764,N_29707);
or UO_950 (O_950,N_29743,N_29589);
or UO_951 (O_951,N_29281,N_28902);
or UO_952 (O_952,N_28884,N_29097);
or UO_953 (O_953,N_29852,N_28954);
and UO_954 (O_954,N_29288,N_29602);
and UO_955 (O_955,N_29202,N_29425);
and UO_956 (O_956,N_29845,N_29172);
xnor UO_957 (O_957,N_28918,N_29187);
and UO_958 (O_958,N_29429,N_29509);
xnor UO_959 (O_959,N_29467,N_29769);
nor UO_960 (O_960,N_29064,N_29112);
nand UO_961 (O_961,N_29258,N_29117);
xor UO_962 (O_962,N_29652,N_29925);
and UO_963 (O_963,N_29847,N_29992);
nor UO_964 (O_964,N_29009,N_29291);
nor UO_965 (O_965,N_28982,N_29389);
or UO_966 (O_966,N_29035,N_29870);
nor UO_967 (O_967,N_29627,N_29610);
or UO_968 (O_968,N_29724,N_29285);
or UO_969 (O_969,N_29804,N_29991);
nor UO_970 (O_970,N_29846,N_29593);
nor UO_971 (O_971,N_29569,N_28941);
or UO_972 (O_972,N_29481,N_29047);
and UO_973 (O_973,N_29721,N_29845);
and UO_974 (O_974,N_29583,N_29239);
xor UO_975 (O_975,N_29275,N_29616);
and UO_976 (O_976,N_28981,N_29988);
xnor UO_977 (O_977,N_29520,N_29374);
nor UO_978 (O_978,N_28820,N_29287);
nor UO_979 (O_979,N_29549,N_29917);
nand UO_980 (O_980,N_29556,N_29294);
nand UO_981 (O_981,N_29637,N_29122);
or UO_982 (O_982,N_29876,N_29177);
or UO_983 (O_983,N_28891,N_28944);
xnor UO_984 (O_984,N_29347,N_29637);
or UO_985 (O_985,N_29262,N_29371);
nand UO_986 (O_986,N_28901,N_28810);
nand UO_987 (O_987,N_29041,N_29869);
or UO_988 (O_988,N_29200,N_29901);
and UO_989 (O_989,N_29261,N_28850);
or UO_990 (O_990,N_29454,N_29979);
xnor UO_991 (O_991,N_29820,N_28876);
nand UO_992 (O_992,N_28945,N_28811);
and UO_993 (O_993,N_29730,N_29905);
or UO_994 (O_994,N_29930,N_28831);
nand UO_995 (O_995,N_29407,N_29984);
nor UO_996 (O_996,N_29483,N_29373);
nand UO_997 (O_997,N_29699,N_29281);
or UO_998 (O_998,N_29954,N_29567);
or UO_999 (O_999,N_29861,N_29895);
or UO_1000 (O_1000,N_28807,N_29433);
nor UO_1001 (O_1001,N_29551,N_29020);
xor UO_1002 (O_1002,N_29310,N_28998);
or UO_1003 (O_1003,N_29246,N_29411);
xnor UO_1004 (O_1004,N_29830,N_29905);
nand UO_1005 (O_1005,N_29891,N_29058);
nor UO_1006 (O_1006,N_29488,N_29133);
nand UO_1007 (O_1007,N_28802,N_29744);
or UO_1008 (O_1008,N_29304,N_29912);
xnor UO_1009 (O_1009,N_29781,N_29862);
nand UO_1010 (O_1010,N_29487,N_29354);
or UO_1011 (O_1011,N_28915,N_29223);
nor UO_1012 (O_1012,N_29662,N_29057);
nand UO_1013 (O_1013,N_29408,N_29469);
and UO_1014 (O_1014,N_29726,N_29216);
nor UO_1015 (O_1015,N_29576,N_29912);
xor UO_1016 (O_1016,N_29867,N_29221);
nand UO_1017 (O_1017,N_28855,N_29610);
and UO_1018 (O_1018,N_28879,N_29089);
xor UO_1019 (O_1019,N_29622,N_29558);
nor UO_1020 (O_1020,N_28912,N_28805);
or UO_1021 (O_1021,N_28920,N_29901);
or UO_1022 (O_1022,N_29049,N_29409);
or UO_1023 (O_1023,N_29903,N_29927);
and UO_1024 (O_1024,N_28980,N_29896);
xor UO_1025 (O_1025,N_29295,N_29304);
nor UO_1026 (O_1026,N_29662,N_29985);
nand UO_1027 (O_1027,N_29207,N_28808);
nor UO_1028 (O_1028,N_29720,N_29703);
and UO_1029 (O_1029,N_29501,N_29686);
or UO_1030 (O_1030,N_29138,N_29171);
and UO_1031 (O_1031,N_28839,N_29861);
or UO_1032 (O_1032,N_29124,N_28894);
xnor UO_1033 (O_1033,N_29704,N_28857);
and UO_1034 (O_1034,N_29527,N_29053);
nor UO_1035 (O_1035,N_29709,N_29277);
xor UO_1036 (O_1036,N_29664,N_29724);
nand UO_1037 (O_1037,N_29881,N_29399);
nand UO_1038 (O_1038,N_29735,N_29465);
xnor UO_1039 (O_1039,N_29499,N_29714);
or UO_1040 (O_1040,N_28958,N_29495);
nor UO_1041 (O_1041,N_29699,N_29524);
xor UO_1042 (O_1042,N_29408,N_29688);
nand UO_1043 (O_1043,N_29893,N_29686);
xor UO_1044 (O_1044,N_29648,N_29941);
or UO_1045 (O_1045,N_28913,N_28826);
and UO_1046 (O_1046,N_28838,N_29142);
and UO_1047 (O_1047,N_29337,N_29084);
nor UO_1048 (O_1048,N_29508,N_29623);
and UO_1049 (O_1049,N_29925,N_29015);
and UO_1050 (O_1050,N_29558,N_29525);
nor UO_1051 (O_1051,N_29809,N_28984);
and UO_1052 (O_1052,N_28841,N_29464);
xor UO_1053 (O_1053,N_29862,N_29227);
nor UO_1054 (O_1054,N_29174,N_28972);
nor UO_1055 (O_1055,N_29831,N_29294);
and UO_1056 (O_1056,N_29022,N_28942);
and UO_1057 (O_1057,N_29846,N_28913);
and UO_1058 (O_1058,N_29645,N_29658);
and UO_1059 (O_1059,N_29884,N_28867);
or UO_1060 (O_1060,N_29856,N_29193);
nor UO_1061 (O_1061,N_28922,N_29290);
and UO_1062 (O_1062,N_29903,N_29262);
xnor UO_1063 (O_1063,N_29956,N_29511);
or UO_1064 (O_1064,N_29606,N_29171);
xnor UO_1065 (O_1065,N_29905,N_29996);
and UO_1066 (O_1066,N_29925,N_29191);
or UO_1067 (O_1067,N_29608,N_29840);
nor UO_1068 (O_1068,N_29343,N_29127);
or UO_1069 (O_1069,N_29520,N_28960);
xor UO_1070 (O_1070,N_29083,N_29134);
or UO_1071 (O_1071,N_29237,N_29873);
and UO_1072 (O_1072,N_29898,N_29084);
xnor UO_1073 (O_1073,N_28886,N_29028);
or UO_1074 (O_1074,N_29475,N_29599);
nor UO_1075 (O_1075,N_29933,N_29618);
and UO_1076 (O_1076,N_29237,N_28986);
and UO_1077 (O_1077,N_29318,N_29595);
and UO_1078 (O_1078,N_29819,N_29862);
and UO_1079 (O_1079,N_29168,N_29183);
or UO_1080 (O_1080,N_29820,N_28831);
nand UO_1081 (O_1081,N_29619,N_29901);
or UO_1082 (O_1082,N_29010,N_28900);
nor UO_1083 (O_1083,N_29569,N_29330);
nor UO_1084 (O_1084,N_29607,N_28954);
nand UO_1085 (O_1085,N_28827,N_29530);
and UO_1086 (O_1086,N_29974,N_29534);
or UO_1087 (O_1087,N_28829,N_28851);
nor UO_1088 (O_1088,N_29569,N_29266);
xnor UO_1089 (O_1089,N_28813,N_29040);
and UO_1090 (O_1090,N_29645,N_29936);
nand UO_1091 (O_1091,N_29886,N_28924);
nand UO_1092 (O_1092,N_29602,N_28940);
nand UO_1093 (O_1093,N_29479,N_29523);
nor UO_1094 (O_1094,N_29738,N_29818);
nand UO_1095 (O_1095,N_29263,N_29165);
xor UO_1096 (O_1096,N_29407,N_29228);
and UO_1097 (O_1097,N_29568,N_29162);
nand UO_1098 (O_1098,N_29819,N_29736);
and UO_1099 (O_1099,N_29633,N_29387);
and UO_1100 (O_1100,N_29604,N_29682);
nor UO_1101 (O_1101,N_28867,N_28820);
nor UO_1102 (O_1102,N_29024,N_29265);
xor UO_1103 (O_1103,N_29613,N_28819);
and UO_1104 (O_1104,N_29928,N_29584);
and UO_1105 (O_1105,N_29697,N_29295);
nor UO_1106 (O_1106,N_29657,N_29355);
nand UO_1107 (O_1107,N_29062,N_29392);
nand UO_1108 (O_1108,N_29677,N_29552);
nor UO_1109 (O_1109,N_29226,N_29935);
nor UO_1110 (O_1110,N_29151,N_29499);
or UO_1111 (O_1111,N_29660,N_29326);
xnor UO_1112 (O_1112,N_29575,N_28878);
nor UO_1113 (O_1113,N_28907,N_29648);
or UO_1114 (O_1114,N_29835,N_28815);
nand UO_1115 (O_1115,N_29171,N_29672);
nand UO_1116 (O_1116,N_29397,N_29648);
xor UO_1117 (O_1117,N_28908,N_28832);
nor UO_1118 (O_1118,N_29543,N_28930);
xnor UO_1119 (O_1119,N_29392,N_29584);
xnor UO_1120 (O_1120,N_29612,N_29368);
or UO_1121 (O_1121,N_29009,N_29447);
and UO_1122 (O_1122,N_29171,N_29494);
nor UO_1123 (O_1123,N_28902,N_28836);
xor UO_1124 (O_1124,N_28852,N_29405);
nand UO_1125 (O_1125,N_29234,N_29398);
or UO_1126 (O_1126,N_29258,N_29244);
xor UO_1127 (O_1127,N_29275,N_29323);
nor UO_1128 (O_1128,N_29380,N_29122);
nor UO_1129 (O_1129,N_29038,N_29106);
xnor UO_1130 (O_1130,N_29065,N_29955);
nand UO_1131 (O_1131,N_29552,N_29593);
xnor UO_1132 (O_1132,N_29920,N_28804);
or UO_1133 (O_1133,N_29573,N_29341);
xor UO_1134 (O_1134,N_29620,N_29266);
or UO_1135 (O_1135,N_29694,N_29697);
nor UO_1136 (O_1136,N_28841,N_29570);
and UO_1137 (O_1137,N_29514,N_29589);
nor UO_1138 (O_1138,N_29159,N_29657);
nor UO_1139 (O_1139,N_29798,N_29685);
or UO_1140 (O_1140,N_29547,N_29240);
or UO_1141 (O_1141,N_29361,N_29770);
or UO_1142 (O_1142,N_29856,N_29058);
and UO_1143 (O_1143,N_29840,N_29198);
and UO_1144 (O_1144,N_28953,N_29936);
xor UO_1145 (O_1145,N_29590,N_29262);
xor UO_1146 (O_1146,N_29504,N_29452);
and UO_1147 (O_1147,N_29076,N_29044);
nand UO_1148 (O_1148,N_29592,N_29240);
and UO_1149 (O_1149,N_29000,N_28804);
xor UO_1150 (O_1150,N_28961,N_29774);
nand UO_1151 (O_1151,N_29289,N_29805);
xor UO_1152 (O_1152,N_29712,N_28809);
and UO_1153 (O_1153,N_29359,N_29523);
nor UO_1154 (O_1154,N_29801,N_29415);
xnor UO_1155 (O_1155,N_29669,N_29560);
and UO_1156 (O_1156,N_29948,N_29392);
nor UO_1157 (O_1157,N_29633,N_29394);
xnor UO_1158 (O_1158,N_28908,N_29079);
and UO_1159 (O_1159,N_29189,N_29745);
nor UO_1160 (O_1160,N_29647,N_29129);
or UO_1161 (O_1161,N_28977,N_29094);
nor UO_1162 (O_1162,N_29277,N_29725);
and UO_1163 (O_1163,N_29550,N_29048);
nor UO_1164 (O_1164,N_29803,N_28812);
xnor UO_1165 (O_1165,N_28929,N_29214);
and UO_1166 (O_1166,N_29541,N_29461);
nor UO_1167 (O_1167,N_29321,N_29038);
or UO_1168 (O_1168,N_29880,N_29578);
nand UO_1169 (O_1169,N_29664,N_28853);
and UO_1170 (O_1170,N_29753,N_29220);
nor UO_1171 (O_1171,N_29158,N_29052);
and UO_1172 (O_1172,N_29286,N_29029);
nand UO_1173 (O_1173,N_28908,N_29789);
xor UO_1174 (O_1174,N_29796,N_29941);
nor UO_1175 (O_1175,N_29221,N_29820);
xor UO_1176 (O_1176,N_29345,N_29853);
or UO_1177 (O_1177,N_29735,N_28839);
nor UO_1178 (O_1178,N_29920,N_29480);
and UO_1179 (O_1179,N_29836,N_29817);
and UO_1180 (O_1180,N_29107,N_29971);
nor UO_1181 (O_1181,N_29271,N_29868);
and UO_1182 (O_1182,N_28841,N_29194);
or UO_1183 (O_1183,N_29537,N_29046);
nand UO_1184 (O_1184,N_29446,N_29735);
xor UO_1185 (O_1185,N_29637,N_29648);
xnor UO_1186 (O_1186,N_29467,N_29279);
nor UO_1187 (O_1187,N_29832,N_28957);
and UO_1188 (O_1188,N_29099,N_28871);
or UO_1189 (O_1189,N_29011,N_29343);
and UO_1190 (O_1190,N_29999,N_28869);
nand UO_1191 (O_1191,N_29590,N_29076);
xnor UO_1192 (O_1192,N_29947,N_28816);
xnor UO_1193 (O_1193,N_29788,N_28995);
and UO_1194 (O_1194,N_29607,N_29024);
and UO_1195 (O_1195,N_29656,N_29314);
or UO_1196 (O_1196,N_29498,N_29892);
nor UO_1197 (O_1197,N_29566,N_29726);
nor UO_1198 (O_1198,N_29450,N_29397);
and UO_1199 (O_1199,N_29916,N_28827);
nand UO_1200 (O_1200,N_29402,N_29152);
xnor UO_1201 (O_1201,N_29631,N_28975);
nor UO_1202 (O_1202,N_29430,N_29391);
xnor UO_1203 (O_1203,N_28879,N_29866);
or UO_1204 (O_1204,N_28909,N_29949);
nor UO_1205 (O_1205,N_28826,N_28923);
or UO_1206 (O_1206,N_29174,N_29158);
or UO_1207 (O_1207,N_29122,N_29311);
xnor UO_1208 (O_1208,N_29290,N_28914);
nand UO_1209 (O_1209,N_29210,N_29063);
or UO_1210 (O_1210,N_29173,N_29903);
or UO_1211 (O_1211,N_29327,N_29818);
nor UO_1212 (O_1212,N_29447,N_29873);
or UO_1213 (O_1213,N_29612,N_28976);
nor UO_1214 (O_1214,N_29985,N_29344);
nor UO_1215 (O_1215,N_29504,N_29506);
and UO_1216 (O_1216,N_29764,N_29012);
or UO_1217 (O_1217,N_28824,N_29622);
or UO_1218 (O_1218,N_29734,N_29479);
or UO_1219 (O_1219,N_29488,N_29512);
or UO_1220 (O_1220,N_29119,N_29940);
or UO_1221 (O_1221,N_29567,N_29079);
nor UO_1222 (O_1222,N_29086,N_28811);
and UO_1223 (O_1223,N_29081,N_29776);
nor UO_1224 (O_1224,N_29931,N_29665);
nor UO_1225 (O_1225,N_29380,N_28885);
nand UO_1226 (O_1226,N_29449,N_29509);
nand UO_1227 (O_1227,N_28923,N_29168);
nand UO_1228 (O_1228,N_29597,N_29846);
xnor UO_1229 (O_1229,N_29303,N_29886);
or UO_1230 (O_1230,N_29355,N_29366);
nand UO_1231 (O_1231,N_29869,N_29695);
nand UO_1232 (O_1232,N_29157,N_29481);
or UO_1233 (O_1233,N_29148,N_29726);
xnor UO_1234 (O_1234,N_29929,N_29788);
xor UO_1235 (O_1235,N_29087,N_29329);
nor UO_1236 (O_1236,N_29299,N_29261);
xor UO_1237 (O_1237,N_28919,N_28947);
nand UO_1238 (O_1238,N_29432,N_29453);
nand UO_1239 (O_1239,N_29496,N_29790);
xnor UO_1240 (O_1240,N_29117,N_29320);
xor UO_1241 (O_1241,N_29655,N_29222);
or UO_1242 (O_1242,N_29502,N_29684);
and UO_1243 (O_1243,N_29415,N_28886);
or UO_1244 (O_1244,N_29845,N_28886);
nor UO_1245 (O_1245,N_29689,N_29377);
or UO_1246 (O_1246,N_29657,N_29181);
and UO_1247 (O_1247,N_29490,N_29806);
xnor UO_1248 (O_1248,N_29347,N_29495);
nand UO_1249 (O_1249,N_29137,N_29273);
xor UO_1250 (O_1250,N_29335,N_29333);
or UO_1251 (O_1251,N_29608,N_29092);
xor UO_1252 (O_1252,N_29407,N_29076);
or UO_1253 (O_1253,N_29888,N_29478);
or UO_1254 (O_1254,N_29533,N_29520);
and UO_1255 (O_1255,N_29222,N_29449);
and UO_1256 (O_1256,N_29169,N_28830);
and UO_1257 (O_1257,N_29884,N_29805);
and UO_1258 (O_1258,N_28844,N_29018);
or UO_1259 (O_1259,N_29810,N_29170);
xnor UO_1260 (O_1260,N_28880,N_29898);
or UO_1261 (O_1261,N_29976,N_29585);
nand UO_1262 (O_1262,N_28927,N_29741);
xor UO_1263 (O_1263,N_29665,N_29310);
nand UO_1264 (O_1264,N_29727,N_29689);
nor UO_1265 (O_1265,N_29411,N_29143);
xnor UO_1266 (O_1266,N_29322,N_29319);
and UO_1267 (O_1267,N_29602,N_29370);
and UO_1268 (O_1268,N_29638,N_29834);
nand UO_1269 (O_1269,N_29223,N_29915);
xnor UO_1270 (O_1270,N_29022,N_29219);
nor UO_1271 (O_1271,N_29489,N_29799);
or UO_1272 (O_1272,N_28872,N_29331);
xor UO_1273 (O_1273,N_29208,N_29319);
nand UO_1274 (O_1274,N_29547,N_28876);
nand UO_1275 (O_1275,N_29408,N_29338);
or UO_1276 (O_1276,N_28843,N_29976);
nand UO_1277 (O_1277,N_29213,N_29459);
and UO_1278 (O_1278,N_29400,N_29225);
nor UO_1279 (O_1279,N_29021,N_29456);
or UO_1280 (O_1280,N_28998,N_29418);
xor UO_1281 (O_1281,N_29106,N_29431);
nor UO_1282 (O_1282,N_29792,N_28949);
or UO_1283 (O_1283,N_29927,N_29936);
nor UO_1284 (O_1284,N_29541,N_29870);
nor UO_1285 (O_1285,N_29033,N_29238);
xnor UO_1286 (O_1286,N_29780,N_29974);
xor UO_1287 (O_1287,N_29044,N_29163);
xor UO_1288 (O_1288,N_29324,N_29493);
xor UO_1289 (O_1289,N_29706,N_29508);
nand UO_1290 (O_1290,N_28893,N_28938);
and UO_1291 (O_1291,N_29930,N_29546);
and UO_1292 (O_1292,N_28823,N_29061);
or UO_1293 (O_1293,N_28932,N_29006);
nand UO_1294 (O_1294,N_29180,N_29139);
and UO_1295 (O_1295,N_29892,N_29740);
nor UO_1296 (O_1296,N_29182,N_29790);
nand UO_1297 (O_1297,N_29335,N_29656);
or UO_1298 (O_1298,N_29287,N_29761);
nor UO_1299 (O_1299,N_29112,N_29951);
nand UO_1300 (O_1300,N_29144,N_29670);
and UO_1301 (O_1301,N_29519,N_29827);
and UO_1302 (O_1302,N_29437,N_29753);
and UO_1303 (O_1303,N_29663,N_29975);
nand UO_1304 (O_1304,N_29682,N_29711);
nor UO_1305 (O_1305,N_29072,N_29057);
or UO_1306 (O_1306,N_28993,N_29030);
xor UO_1307 (O_1307,N_29370,N_29631);
nand UO_1308 (O_1308,N_29790,N_29005);
xor UO_1309 (O_1309,N_29125,N_29284);
xnor UO_1310 (O_1310,N_28807,N_29416);
xor UO_1311 (O_1311,N_29282,N_29119);
xnor UO_1312 (O_1312,N_29607,N_29909);
xor UO_1313 (O_1313,N_29174,N_29302);
nor UO_1314 (O_1314,N_29764,N_29052);
xnor UO_1315 (O_1315,N_29893,N_29502);
nor UO_1316 (O_1316,N_29657,N_29115);
nor UO_1317 (O_1317,N_29809,N_29489);
and UO_1318 (O_1318,N_29056,N_29897);
or UO_1319 (O_1319,N_29780,N_29436);
or UO_1320 (O_1320,N_29982,N_28890);
nor UO_1321 (O_1321,N_29509,N_29475);
nand UO_1322 (O_1322,N_29095,N_29171);
xnor UO_1323 (O_1323,N_29157,N_29958);
or UO_1324 (O_1324,N_29545,N_29501);
xnor UO_1325 (O_1325,N_29917,N_29078);
nand UO_1326 (O_1326,N_29711,N_29700);
nand UO_1327 (O_1327,N_29835,N_29881);
nor UO_1328 (O_1328,N_29717,N_29817);
nor UO_1329 (O_1329,N_29268,N_29064);
nor UO_1330 (O_1330,N_29189,N_29696);
nor UO_1331 (O_1331,N_29871,N_28961);
and UO_1332 (O_1332,N_28838,N_29977);
and UO_1333 (O_1333,N_29628,N_29527);
and UO_1334 (O_1334,N_29037,N_28868);
nand UO_1335 (O_1335,N_29467,N_29482);
and UO_1336 (O_1336,N_28968,N_28880);
and UO_1337 (O_1337,N_29267,N_29604);
xnor UO_1338 (O_1338,N_29020,N_29979);
xor UO_1339 (O_1339,N_29163,N_29368);
nor UO_1340 (O_1340,N_28948,N_28934);
xor UO_1341 (O_1341,N_29166,N_29031);
or UO_1342 (O_1342,N_29884,N_29051);
nor UO_1343 (O_1343,N_29660,N_29511);
and UO_1344 (O_1344,N_29047,N_29615);
nor UO_1345 (O_1345,N_29753,N_29919);
and UO_1346 (O_1346,N_29699,N_29522);
nand UO_1347 (O_1347,N_29359,N_29779);
or UO_1348 (O_1348,N_28885,N_29768);
and UO_1349 (O_1349,N_29143,N_29182);
nand UO_1350 (O_1350,N_29619,N_29159);
or UO_1351 (O_1351,N_29205,N_29780);
and UO_1352 (O_1352,N_29399,N_29470);
nor UO_1353 (O_1353,N_29384,N_28988);
xor UO_1354 (O_1354,N_29121,N_29885);
nor UO_1355 (O_1355,N_29308,N_29992);
and UO_1356 (O_1356,N_29140,N_29072);
nor UO_1357 (O_1357,N_29903,N_28852);
or UO_1358 (O_1358,N_29007,N_29383);
xor UO_1359 (O_1359,N_29327,N_29336);
and UO_1360 (O_1360,N_29366,N_28933);
nor UO_1361 (O_1361,N_29888,N_29943);
and UO_1362 (O_1362,N_28875,N_29384);
nand UO_1363 (O_1363,N_28830,N_29793);
and UO_1364 (O_1364,N_29392,N_28807);
nand UO_1365 (O_1365,N_29574,N_29999);
nor UO_1366 (O_1366,N_28883,N_29145);
and UO_1367 (O_1367,N_29449,N_29337);
nand UO_1368 (O_1368,N_29841,N_29258);
and UO_1369 (O_1369,N_29706,N_29689);
xnor UO_1370 (O_1370,N_29265,N_29386);
or UO_1371 (O_1371,N_29514,N_29096);
and UO_1372 (O_1372,N_29693,N_29332);
nand UO_1373 (O_1373,N_29396,N_29896);
or UO_1374 (O_1374,N_29367,N_29353);
nor UO_1375 (O_1375,N_29285,N_29798);
xnor UO_1376 (O_1376,N_29269,N_29085);
or UO_1377 (O_1377,N_29533,N_29281);
and UO_1378 (O_1378,N_29974,N_28836);
and UO_1379 (O_1379,N_29813,N_28891);
xnor UO_1380 (O_1380,N_29659,N_28977);
xnor UO_1381 (O_1381,N_29923,N_28842);
and UO_1382 (O_1382,N_29012,N_29356);
nand UO_1383 (O_1383,N_29341,N_29329);
xor UO_1384 (O_1384,N_29669,N_29737);
xor UO_1385 (O_1385,N_29808,N_29974);
or UO_1386 (O_1386,N_29861,N_29316);
or UO_1387 (O_1387,N_29636,N_29598);
or UO_1388 (O_1388,N_29420,N_29697);
nand UO_1389 (O_1389,N_29811,N_28998);
xor UO_1390 (O_1390,N_29421,N_28942);
and UO_1391 (O_1391,N_29104,N_28882);
or UO_1392 (O_1392,N_29017,N_28871);
xor UO_1393 (O_1393,N_29545,N_29257);
and UO_1394 (O_1394,N_29014,N_29735);
xnor UO_1395 (O_1395,N_28817,N_29152);
nor UO_1396 (O_1396,N_29640,N_29966);
or UO_1397 (O_1397,N_29948,N_29860);
or UO_1398 (O_1398,N_29151,N_28821);
xnor UO_1399 (O_1399,N_29650,N_29675);
and UO_1400 (O_1400,N_29093,N_29876);
nor UO_1401 (O_1401,N_29428,N_29260);
or UO_1402 (O_1402,N_29335,N_29986);
nor UO_1403 (O_1403,N_29961,N_29785);
and UO_1404 (O_1404,N_29802,N_29189);
or UO_1405 (O_1405,N_29266,N_29092);
nor UO_1406 (O_1406,N_28950,N_29024);
xnor UO_1407 (O_1407,N_29434,N_29254);
and UO_1408 (O_1408,N_29578,N_29485);
xor UO_1409 (O_1409,N_29444,N_29245);
nand UO_1410 (O_1410,N_29685,N_29489);
nor UO_1411 (O_1411,N_29111,N_29279);
and UO_1412 (O_1412,N_29500,N_29448);
and UO_1413 (O_1413,N_29853,N_29398);
nor UO_1414 (O_1414,N_28970,N_29658);
nor UO_1415 (O_1415,N_29495,N_29720);
nand UO_1416 (O_1416,N_28849,N_29590);
nand UO_1417 (O_1417,N_29168,N_29427);
nand UO_1418 (O_1418,N_29677,N_29370);
nor UO_1419 (O_1419,N_29129,N_29292);
nand UO_1420 (O_1420,N_29169,N_29560);
nor UO_1421 (O_1421,N_29266,N_29573);
nand UO_1422 (O_1422,N_29770,N_29333);
or UO_1423 (O_1423,N_28960,N_29192);
or UO_1424 (O_1424,N_29672,N_29242);
or UO_1425 (O_1425,N_29149,N_29227);
nor UO_1426 (O_1426,N_29500,N_29542);
nor UO_1427 (O_1427,N_29081,N_28936);
and UO_1428 (O_1428,N_29920,N_28904);
xor UO_1429 (O_1429,N_29591,N_29736);
xor UO_1430 (O_1430,N_29423,N_29498);
or UO_1431 (O_1431,N_29643,N_29405);
or UO_1432 (O_1432,N_29230,N_29227);
or UO_1433 (O_1433,N_29683,N_29890);
and UO_1434 (O_1434,N_29355,N_29194);
xnor UO_1435 (O_1435,N_29860,N_29078);
nor UO_1436 (O_1436,N_29802,N_28935);
and UO_1437 (O_1437,N_29200,N_29974);
or UO_1438 (O_1438,N_29392,N_29621);
nand UO_1439 (O_1439,N_29478,N_29140);
nor UO_1440 (O_1440,N_29557,N_29115);
or UO_1441 (O_1441,N_29489,N_29479);
nor UO_1442 (O_1442,N_29812,N_29814);
nor UO_1443 (O_1443,N_29288,N_29603);
and UO_1444 (O_1444,N_29042,N_28852);
or UO_1445 (O_1445,N_29141,N_28848);
and UO_1446 (O_1446,N_28919,N_29926);
nand UO_1447 (O_1447,N_28920,N_29561);
xor UO_1448 (O_1448,N_29192,N_29389);
xor UO_1449 (O_1449,N_29683,N_29490);
and UO_1450 (O_1450,N_29659,N_29789);
nand UO_1451 (O_1451,N_29681,N_29728);
or UO_1452 (O_1452,N_29583,N_29039);
nand UO_1453 (O_1453,N_29126,N_29557);
and UO_1454 (O_1454,N_29511,N_29047);
and UO_1455 (O_1455,N_29745,N_29165);
xor UO_1456 (O_1456,N_29481,N_28897);
xnor UO_1457 (O_1457,N_29912,N_28872);
nand UO_1458 (O_1458,N_29103,N_29810);
nand UO_1459 (O_1459,N_29004,N_29326);
and UO_1460 (O_1460,N_29611,N_29129);
xnor UO_1461 (O_1461,N_29420,N_28912);
nand UO_1462 (O_1462,N_29217,N_29896);
and UO_1463 (O_1463,N_28854,N_29682);
and UO_1464 (O_1464,N_29337,N_28836);
nand UO_1465 (O_1465,N_29530,N_28985);
nand UO_1466 (O_1466,N_29833,N_28877);
nor UO_1467 (O_1467,N_29405,N_29759);
or UO_1468 (O_1468,N_29655,N_29965);
xor UO_1469 (O_1469,N_29955,N_29938);
xor UO_1470 (O_1470,N_29970,N_29088);
and UO_1471 (O_1471,N_29358,N_29398);
nor UO_1472 (O_1472,N_29340,N_29636);
nor UO_1473 (O_1473,N_29656,N_29408);
nand UO_1474 (O_1474,N_29356,N_29567);
xnor UO_1475 (O_1475,N_29894,N_29959);
nor UO_1476 (O_1476,N_29527,N_28889);
xnor UO_1477 (O_1477,N_29241,N_29268);
and UO_1478 (O_1478,N_29536,N_28858);
xnor UO_1479 (O_1479,N_29657,N_29012);
nor UO_1480 (O_1480,N_29381,N_29333);
and UO_1481 (O_1481,N_29270,N_29805);
nor UO_1482 (O_1482,N_29901,N_29958);
or UO_1483 (O_1483,N_29301,N_29043);
or UO_1484 (O_1484,N_29904,N_28847);
or UO_1485 (O_1485,N_29035,N_29604);
or UO_1486 (O_1486,N_29038,N_29168);
xnor UO_1487 (O_1487,N_29717,N_29453);
and UO_1488 (O_1488,N_29199,N_29257);
and UO_1489 (O_1489,N_28826,N_29657);
nor UO_1490 (O_1490,N_29739,N_28986);
and UO_1491 (O_1491,N_29322,N_29432);
nor UO_1492 (O_1492,N_29726,N_29634);
nand UO_1493 (O_1493,N_28845,N_29270);
xnor UO_1494 (O_1494,N_29241,N_29222);
and UO_1495 (O_1495,N_29038,N_29167);
nor UO_1496 (O_1496,N_29780,N_29658);
xnor UO_1497 (O_1497,N_29108,N_29000);
or UO_1498 (O_1498,N_28924,N_29133);
or UO_1499 (O_1499,N_29244,N_28853);
xnor UO_1500 (O_1500,N_29144,N_29344);
nand UO_1501 (O_1501,N_29266,N_29242);
nand UO_1502 (O_1502,N_29565,N_29485);
or UO_1503 (O_1503,N_29670,N_29572);
or UO_1504 (O_1504,N_29698,N_28802);
nor UO_1505 (O_1505,N_29262,N_29126);
xnor UO_1506 (O_1506,N_29014,N_29050);
xnor UO_1507 (O_1507,N_28976,N_29221);
and UO_1508 (O_1508,N_29442,N_29024);
nor UO_1509 (O_1509,N_29116,N_28885);
nor UO_1510 (O_1510,N_29656,N_29788);
xnor UO_1511 (O_1511,N_28838,N_29061);
nand UO_1512 (O_1512,N_29106,N_28897);
and UO_1513 (O_1513,N_29185,N_29151);
nand UO_1514 (O_1514,N_29896,N_29491);
nor UO_1515 (O_1515,N_29343,N_29221);
xor UO_1516 (O_1516,N_28835,N_29804);
nand UO_1517 (O_1517,N_29865,N_28866);
and UO_1518 (O_1518,N_29369,N_28829);
nand UO_1519 (O_1519,N_29853,N_29457);
or UO_1520 (O_1520,N_29011,N_29712);
nor UO_1521 (O_1521,N_28882,N_29583);
xor UO_1522 (O_1522,N_29015,N_29860);
nand UO_1523 (O_1523,N_29935,N_28963);
or UO_1524 (O_1524,N_29346,N_28904);
xor UO_1525 (O_1525,N_29380,N_29068);
xor UO_1526 (O_1526,N_29456,N_29362);
xor UO_1527 (O_1527,N_29495,N_29472);
xor UO_1528 (O_1528,N_29199,N_29703);
or UO_1529 (O_1529,N_29926,N_29916);
nand UO_1530 (O_1530,N_29672,N_28974);
or UO_1531 (O_1531,N_29660,N_29590);
nand UO_1532 (O_1532,N_29790,N_29991);
nor UO_1533 (O_1533,N_28973,N_29619);
or UO_1534 (O_1534,N_29128,N_28816);
xor UO_1535 (O_1535,N_29692,N_29981);
and UO_1536 (O_1536,N_29042,N_29305);
xnor UO_1537 (O_1537,N_29556,N_29824);
nand UO_1538 (O_1538,N_29965,N_29203);
and UO_1539 (O_1539,N_28903,N_29888);
nand UO_1540 (O_1540,N_29954,N_29483);
or UO_1541 (O_1541,N_28875,N_29639);
and UO_1542 (O_1542,N_29014,N_29603);
or UO_1543 (O_1543,N_29794,N_29212);
and UO_1544 (O_1544,N_29901,N_28956);
or UO_1545 (O_1545,N_29524,N_28800);
or UO_1546 (O_1546,N_29719,N_29723);
nand UO_1547 (O_1547,N_29287,N_29259);
xor UO_1548 (O_1548,N_29161,N_29106);
and UO_1549 (O_1549,N_29049,N_29136);
or UO_1550 (O_1550,N_29332,N_29398);
nor UO_1551 (O_1551,N_28886,N_29126);
or UO_1552 (O_1552,N_29926,N_29260);
or UO_1553 (O_1553,N_29639,N_29516);
xor UO_1554 (O_1554,N_29864,N_29000);
nor UO_1555 (O_1555,N_29789,N_29440);
or UO_1556 (O_1556,N_29631,N_29688);
nor UO_1557 (O_1557,N_29450,N_29610);
and UO_1558 (O_1558,N_29636,N_29611);
xnor UO_1559 (O_1559,N_28860,N_29252);
xor UO_1560 (O_1560,N_29054,N_29929);
nand UO_1561 (O_1561,N_29963,N_29810);
xnor UO_1562 (O_1562,N_29040,N_29517);
or UO_1563 (O_1563,N_29478,N_28911);
nor UO_1564 (O_1564,N_29364,N_28982);
xor UO_1565 (O_1565,N_29784,N_29535);
xnor UO_1566 (O_1566,N_28867,N_28979);
and UO_1567 (O_1567,N_29320,N_29644);
nor UO_1568 (O_1568,N_29950,N_29171);
or UO_1569 (O_1569,N_28826,N_29248);
nor UO_1570 (O_1570,N_28898,N_29808);
and UO_1571 (O_1571,N_29831,N_29087);
nand UO_1572 (O_1572,N_29292,N_29555);
or UO_1573 (O_1573,N_29605,N_29061);
or UO_1574 (O_1574,N_29566,N_28835);
or UO_1575 (O_1575,N_29549,N_29598);
xnor UO_1576 (O_1576,N_29478,N_29585);
xnor UO_1577 (O_1577,N_29079,N_29171);
nor UO_1578 (O_1578,N_29904,N_29292);
or UO_1579 (O_1579,N_29282,N_29175);
and UO_1580 (O_1580,N_29853,N_28966);
nand UO_1581 (O_1581,N_29621,N_29847);
nor UO_1582 (O_1582,N_28916,N_28825);
or UO_1583 (O_1583,N_29962,N_29513);
xor UO_1584 (O_1584,N_28985,N_28958);
nand UO_1585 (O_1585,N_28885,N_29488);
xnor UO_1586 (O_1586,N_29837,N_29825);
and UO_1587 (O_1587,N_29002,N_29640);
or UO_1588 (O_1588,N_29628,N_29635);
xnor UO_1589 (O_1589,N_29029,N_29960);
nand UO_1590 (O_1590,N_29976,N_29675);
nor UO_1591 (O_1591,N_29485,N_29791);
or UO_1592 (O_1592,N_29783,N_29163);
xnor UO_1593 (O_1593,N_28871,N_29660);
nand UO_1594 (O_1594,N_29716,N_29291);
and UO_1595 (O_1595,N_29548,N_29461);
nor UO_1596 (O_1596,N_28999,N_29818);
nand UO_1597 (O_1597,N_29686,N_28835);
nand UO_1598 (O_1598,N_29611,N_29328);
nand UO_1599 (O_1599,N_29285,N_29491);
xnor UO_1600 (O_1600,N_28980,N_29742);
xor UO_1601 (O_1601,N_29247,N_29228);
nand UO_1602 (O_1602,N_29755,N_29867);
nand UO_1603 (O_1603,N_29933,N_28811);
xor UO_1604 (O_1604,N_29610,N_29134);
xor UO_1605 (O_1605,N_29243,N_29071);
or UO_1606 (O_1606,N_29808,N_29207);
nor UO_1607 (O_1607,N_29856,N_29607);
or UO_1608 (O_1608,N_29613,N_29574);
and UO_1609 (O_1609,N_29780,N_29041);
and UO_1610 (O_1610,N_29941,N_29966);
and UO_1611 (O_1611,N_29665,N_29210);
or UO_1612 (O_1612,N_29233,N_29059);
or UO_1613 (O_1613,N_29491,N_29735);
nand UO_1614 (O_1614,N_29745,N_29790);
xnor UO_1615 (O_1615,N_29714,N_29198);
nor UO_1616 (O_1616,N_29480,N_29988);
and UO_1617 (O_1617,N_29569,N_29728);
nor UO_1618 (O_1618,N_29094,N_29065);
nand UO_1619 (O_1619,N_29966,N_29504);
and UO_1620 (O_1620,N_29535,N_28984);
xnor UO_1621 (O_1621,N_29636,N_29895);
xnor UO_1622 (O_1622,N_28950,N_28800);
nor UO_1623 (O_1623,N_29947,N_28931);
nand UO_1624 (O_1624,N_28834,N_28928);
nand UO_1625 (O_1625,N_28804,N_29014);
nor UO_1626 (O_1626,N_29038,N_29963);
nand UO_1627 (O_1627,N_29483,N_29984);
nor UO_1628 (O_1628,N_29353,N_29610);
and UO_1629 (O_1629,N_28897,N_28950);
or UO_1630 (O_1630,N_29117,N_29915);
xnor UO_1631 (O_1631,N_29808,N_28886);
or UO_1632 (O_1632,N_29092,N_29042);
nor UO_1633 (O_1633,N_29831,N_29342);
and UO_1634 (O_1634,N_29277,N_29653);
xor UO_1635 (O_1635,N_28817,N_28997);
nor UO_1636 (O_1636,N_28979,N_29926);
and UO_1637 (O_1637,N_29998,N_29377);
nor UO_1638 (O_1638,N_28843,N_29550);
or UO_1639 (O_1639,N_29877,N_29607);
or UO_1640 (O_1640,N_29960,N_29448);
or UO_1641 (O_1641,N_29722,N_29979);
or UO_1642 (O_1642,N_29253,N_29418);
and UO_1643 (O_1643,N_29132,N_29728);
or UO_1644 (O_1644,N_28900,N_29130);
nor UO_1645 (O_1645,N_29637,N_29585);
nor UO_1646 (O_1646,N_29796,N_29681);
nor UO_1647 (O_1647,N_29233,N_29825);
nand UO_1648 (O_1648,N_29668,N_29727);
nand UO_1649 (O_1649,N_29738,N_29160);
or UO_1650 (O_1650,N_28863,N_29319);
and UO_1651 (O_1651,N_29306,N_29909);
or UO_1652 (O_1652,N_29817,N_29821);
nand UO_1653 (O_1653,N_29916,N_29320);
or UO_1654 (O_1654,N_29731,N_29639);
nand UO_1655 (O_1655,N_29249,N_29714);
xnor UO_1656 (O_1656,N_28847,N_29829);
or UO_1657 (O_1657,N_29657,N_29518);
xor UO_1658 (O_1658,N_29827,N_29613);
xnor UO_1659 (O_1659,N_29410,N_28954);
xnor UO_1660 (O_1660,N_29883,N_29984);
xor UO_1661 (O_1661,N_29805,N_29830);
nor UO_1662 (O_1662,N_29163,N_29184);
xnor UO_1663 (O_1663,N_28826,N_29963);
and UO_1664 (O_1664,N_29089,N_29954);
nor UO_1665 (O_1665,N_29167,N_29365);
xnor UO_1666 (O_1666,N_29771,N_29963);
nand UO_1667 (O_1667,N_29904,N_29970);
or UO_1668 (O_1668,N_28945,N_29646);
nor UO_1669 (O_1669,N_28929,N_29286);
nor UO_1670 (O_1670,N_29593,N_28873);
or UO_1671 (O_1671,N_29591,N_29208);
nor UO_1672 (O_1672,N_29883,N_29418);
and UO_1673 (O_1673,N_28955,N_29942);
xnor UO_1674 (O_1674,N_29838,N_29571);
and UO_1675 (O_1675,N_28918,N_29854);
or UO_1676 (O_1676,N_29787,N_29435);
or UO_1677 (O_1677,N_29220,N_29067);
or UO_1678 (O_1678,N_29405,N_29107);
or UO_1679 (O_1679,N_29571,N_29638);
nor UO_1680 (O_1680,N_29393,N_28807);
or UO_1681 (O_1681,N_29449,N_29168);
nor UO_1682 (O_1682,N_29757,N_28984);
nand UO_1683 (O_1683,N_29996,N_29499);
or UO_1684 (O_1684,N_29194,N_29712);
nand UO_1685 (O_1685,N_29995,N_29082);
and UO_1686 (O_1686,N_28997,N_29272);
nor UO_1687 (O_1687,N_29699,N_29757);
nor UO_1688 (O_1688,N_29122,N_29867);
xnor UO_1689 (O_1689,N_29247,N_29951);
xnor UO_1690 (O_1690,N_28987,N_29384);
nor UO_1691 (O_1691,N_29314,N_29504);
nor UO_1692 (O_1692,N_29885,N_29951);
nor UO_1693 (O_1693,N_28988,N_29955);
and UO_1694 (O_1694,N_28869,N_29843);
nor UO_1695 (O_1695,N_29573,N_29712);
or UO_1696 (O_1696,N_29536,N_29626);
nand UO_1697 (O_1697,N_29620,N_29389);
xor UO_1698 (O_1698,N_29718,N_29886);
or UO_1699 (O_1699,N_29178,N_28856);
or UO_1700 (O_1700,N_29139,N_28924);
nand UO_1701 (O_1701,N_29382,N_29412);
nor UO_1702 (O_1702,N_29528,N_29015);
and UO_1703 (O_1703,N_28973,N_29581);
and UO_1704 (O_1704,N_29013,N_29972);
xor UO_1705 (O_1705,N_29351,N_29322);
or UO_1706 (O_1706,N_29250,N_28973);
xnor UO_1707 (O_1707,N_29928,N_29753);
nor UO_1708 (O_1708,N_29770,N_28856);
xnor UO_1709 (O_1709,N_29788,N_29119);
nand UO_1710 (O_1710,N_28948,N_29709);
nor UO_1711 (O_1711,N_29414,N_29738);
xor UO_1712 (O_1712,N_29512,N_29193);
and UO_1713 (O_1713,N_29922,N_29503);
or UO_1714 (O_1714,N_29477,N_29999);
nor UO_1715 (O_1715,N_29009,N_29204);
xnor UO_1716 (O_1716,N_29841,N_29802);
nor UO_1717 (O_1717,N_29443,N_29100);
or UO_1718 (O_1718,N_29568,N_29813);
nand UO_1719 (O_1719,N_29601,N_29239);
and UO_1720 (O_1720,N_29673,N_29433);
nand UO_1721 (O_1721,N_29867,N_29160);
nand UO_1722 (O_1722,N_29289,N_29331);
and UO_1723 (O_1723,N_29454,N_29993);
and UO_1724 (O_1724,N_29732,N_29504);
and UO_1725 (O_1725,N_29055,N_29342);
nor UO_1726 (O_1726,N_29686,N_28971);
nand UO_1727 (O_1727,N_28999,N_29077);
and UO_1728 (O_1728,N_29332,N_29133);
nor UO_1729 (O_1729,N_29844,N_29313);
or UO_1730 (O_1730,N_29957,N_29310);
nor UO_1731 (O_1731,N_29685,N_29776);
nand UO_1732 (O_1732,N_29654,N_29143);
and UO_1733 (O_1733,N_28859,N_29628);
and UO_1734 (O_1734,N_28895,N_29683);
xor UO_1735 (O_1735,N_29885,N_29636);
nand UO_1736 (O_1736,N_29931,N_29051);
and UO_1737 (O_1737,N_29329,N_29948);
or UO_1738 (O_1738,N_29478,N_29890);
or UO_1739 (O_1739,N_28889,N_29185);
xnor UO_1740 (O_1740,N_29003,N_29503);
nor UO_1741 (O_1741,N_28946,N_28999);
and UO_1742 (O_1742,N_29836,N_29543);
or UO_1743 (O_1743,N_28858,N_29043);
or UO_1744 (O_1744,N_29789,N_29101);
nor UO_1745 (O_1745,N_29292,N_29512);
nor UO_1746 (O_1746,N_29838,N_29063);
xnor UO_1747 (O_1747,N_29705,N_29214);
nor UO_1748 (O_1748,N_29204,N_28845);
and UO_1749 (O_1749,N_29348,N_29428);
nor UO_1750 (O_1750,N_28923,N_29399);
or UO_1751 (O_1751,N_29984,N_29171);
nand UO_1752 (O_1752,N_29148,N_29014);
nor UO_1753 (O_1753,N_29750,N_29405);
or UO_1754 (O_1754,N_29747,N_29969);
xnor UO_1755 (O_1755,N_28954,N_29276);
and UO_1756 (O_1756,N_29816,N_28929);
xnor UO_1757 (O_1757,N_29173,N_29006);
or UO_1758 (O_1758,N_29718,N_29306);
and UO_1759 (O_1759,N_29244,N_29362);
or UO_1760 (O_1760,N_29269,N_29460);
nand UO_1761 (O_1761,N_29644,N_29782);
nor UO_1762 (O_1762,N_28990,N_29824);
or UO_1763 (O_1763,N_29365,N_29395);
nand UO_1764 (O_1764,N_29102,N_29045);
or UO_1765 (O_1765,N_29577,N_29006);
and UO_1766 (O_1766,N_29083,N_29345);
and UO_1767 (O_1767,N_29859,N_28862);
or UO_1768 (O_1768,N_29371,N_29968);
and UO_1769 (O_1769,N_29154,N_29507);
xor UO_1770 (O_1770,N_29284,N_29041);
xor UO_1771 (O_1771,N_29267,N_29762);
nor UO_1772 (O_1772,N_29924,N_29815);
and UO_1773 (O_1773,N_29644,N_29923);
xor UO_1774 (O_1774,N_28964,N_29577);
or UO_1775 (O_1775,N_29771,N_29554);
xor UO_1776 (O_1776,N_28910,N_29391);
xnor UO_1777 (O_1777,N_29609,N_29007);
nor UO_1778 (O_1778,N_29572,N_28970);
and UO_1779 (O_1779,N_29199,N_29778);
and UO_1780 (O_1780,N_29564,N_29722);
nor UO_1781 (O_1781,N_29025,N_29283);
nor UO_1782 (O_1782,N_29283,N_29831);
nor UO_1783 (O_1783,N_29093,N_29753);
xnor UO_1784 (O_1784,N_29708,N_29471);
or UO_1785 (O_1785,N_29264,N_29633);
or UO_1786 (O_1786,N_28981,N_29544);
xor UO_1787 (O_1787,N_29855,N_28817);
nand UO_1788 (O_1788,N_28815,N_28801);
or UO_1789 (O_1789,N_28845,N_28859);
nor UO_1790 (O_1790,N_29980,N_29165);
nand UO_1791 (O_1791,N_29277,N_29519);
and UO_1792 (O_1792,N_29331,N_29512);
xor UO_1793 (O_1793,N_29806,N_28972);
nor UO_1794 (O_1794,N_29188,N_29745);
or UO_1795 (O_1795,N_29613,N_29899);
nor UO_1796 (O_1796,N_29188,N_29083);
and UO_1797 (O_1797,N_29220,N_29331);
nand UO_1798 (O_1798,N_29620,N_29175);
nand UO_1799 (O_1799,N_29847,N_29301);
xor UO_1800 (O_1800,N_29205,N_29758);
nand UO_1801 (O_1801,N_29465,N_29386);
nor UO_1802 (O_1802,N_29012,N_29471);
or UO_1803 (O_1803,N_29176,N_29022);
xor UO_1804 (O_1804,N_29457,N_28980);
nor UO_1805 (O_1805,N_28880,N_29942);
nand UO_1806 (O_1806,N_29533,N_29188);
xor UO_1807 (O_1807,N_29409,N_28851);
nor UO_1808 (O_1808,N_29790,N_29192);
or UO_1809 (O_1809,N_28945,N_29469);
xnor UO_1810 (O_1810,N_29870,N_29376);
or UO_1811 (O_1811,N_29794,N_29626);
xnor UO_1812 (O_1812,N_29942,N_29627);
nand UO_1813 (O_1813,N_29977,N_29711);
nand UO_1814 (O_1814,N_29541,N_29720);
nor UO_1815 (O_1815,N_29398,N_29933);
xor UO_1816 (O_1816,N_29659,N_29486);
nor UO_1817 (O_1817,N_29330,N_29800);
xnor UO_1818 (O_1818,N_29544,N_29557);
or UO_1819 (O_1819,N_29651,N_29358);
or UO_1820 (O_1820,N_29146,N_28850);
xnor UO_1821 (O_1821,N_29258,N_29073);
nand UO_1822 (O_1822,N_29960,N_28907);
and UO_1823 (O_1823,N_29484,N_29512);
and UO_1824 (O_1824,N_29692,N_28895);
and UO_1825 (O_1825,N_29934,N_29041);
and UO_1826 (O_1826,N_29672,N_29480);
or UO_1827 (O_1827,N_28928,N_29283);
xnor UO_1828 (O_1828,N_29010,N_29341);
and UO_1829 (O_1829,N_29146,N_28822);
xnor UO_1830 (O_1830,N_29831,N_29490);
or UO_1831 (O_1831,N_28922,N_29086);
xnor UO_1832 (O_1832,N_29214,N_29945);
nor UO_1833 (O_1833,N_29809,N_28999);
nor UO_1834 (O_1834,N_29257,N_28999);
nand UO_1835 (O_1835,N_28905,N_29197);
or UO_1836 (O_1836,N_29992,N_29516);
nand UO_1837 (O_1837,N_29360,N_29382);
and UO_1838 (O_1838,N_28868,N_29999);
xnor UO_1839 (O_1839,N_29357,N_28843);
or UO_1840 (O_1840,N_29830,N_29061);
nor UO_1841 (O_1841,N_29959,N_29101);
nand UO_1842 (O_1842,N_29263,N_29788);
or UO_1843 (O_1843,N_29979,N_28949);
xnor UO_1844 (O_1844,N_29114,N_29853);
nor UO_1845 (O_1845,N_29151,N_29866);
and UO_1846 (O_1846,N_29488,N_29769);
or UO_1847 (O_1847,N_29241,N_28921);
or UO_1848 (O_1848,N_29703,N_29868);
xor UO_1849 (O_1849,N_29020,N_29728);
nand UO_1850 (O_1850,N_28889,N_29329);
nor UO_1851 (O_1851,N_29519,N_29690);
nand UO_1852 (O_1852,N_29244,N_29755);
nand UO_1853 (O_1853,N_29079,N_29031);
nor UO_1854 (O_1854,N_29929,N_29216);
and UO_1855 (O_1855,N_29459,N_28906);
xor UO_1856 (O_1856,N_29290,N_29928);
and UO_1857 (O_1857,N_29372,N_28994);
nand UO_1858 (O_1858,N_29086,N_29640);
nand UO_1859 (O_1859,N_29001,N_29830);
or UO_1860 (O_1860,N_29822,N_29101);
or UO_1861 (O_1861,N_29732,N_29445);
xor UO_1862 (O_1862,N_29077,N_29459);
or UO_1863 (O_1863,N_29044,N_29082);
xnor UO_1864 (O_1864,N_29046,N_29858);
nor UO_1865 (O_1865,N_29320,N_29229);
or UO_1866 (O_1866,N_29081,N_29086);
nor UO_1867 (O_1867,N_29131,N_29704);
nor UO_1868 (O_1868,N_29252,N_29694);
nor UO_1869 (O_1869,N_29124,N_29817);
or UO_1870 (O_1870,N_29455,N_29248);
nor UO_1871 (O_1871,N_29325,N_28824);
and UO_1872 (O_1872,N_29737,N_29502);
and UO_1873 (O_1873,N_29194,N_29134);
nor UO_1874 (O_1874,N_29385,N_28946);
nand UO_1875 (O_1875,N_28993,N_29663);
nor UO_1876 (O_1876,N_28920,N_29477);
and UO_1877 (O_1877,N_28994,N_29537);
nor UO_1878 (O_1878,N_28845,N_29338);
nor UO_1879 (O_1879,N_28963,N_29458);
nand UO_1880 (O_1880,N_28974,N_29231);
or UO_1881 (O_1881,N_29467,N_29549);
nor UO_1882 (O_1882,N_29808,N_29033);
nor UO_1883 (O_1883,N_29712,N_28890);
nor UO_1884 (O_1884,N_29757,N_29125);
and UO_1885 (O_1885,N_28941,N_29229);
xor UO_1886 (O_1886,N_29737,N_29862);
nor UO_1887 (O_1887,N_29975,N_29998);
and UO_1888 (O_1888,N_29820,N_28907);
nor UO_1889 (O_1889,N_29138,N_29431);
nor UO_1890 (O_1890,N_29166,N_28887);
and UO_1891 (O_1891,N_29027,N_29435);
nor UO_1892 (O_1892,N_28836,N_29184);
and UO_1893 (O_1893,N_29123,N_29437);
nor UO_1894 (O_1894,N_29643,N_29616);
nor UO_1895 (O_1895,N_29374,N_29478);
nor UO_1896 (O_1896,N_28886,N_29204);
or UO_1897 (O_1897,N_29400,N_28991);
or UO_1898 (O_1898,N_29182,N_29836);
xor UO_1899 (O_1899,N_28860,N_29843);
nand UO_1900 (O_1900,N_29142,N_29355);
nor UO_1901 (O_1901,N_28947,N_29368);
nor UO_1902 (O_1902,N_29380,N_29316);
and UO_1903 (O_1903,N_28863,N_29750);
nand UO_1904 (O_1904,N_29370,N_29206);
nor UO_1905 (O_1905,N_29915,N_29282);
xor UO_1906 (O_1906,N_28901,N_29504);
xor UO_1907 (O_1907,N_29315,N_29276);
nor UO_1908 (O_1908,N_28897,N_29050);
xor UO_1909 (O_1909,N_29809,N_28941);
or UO_1910 (O_1910,N_29088,N_29694);
and UO_1911 (O_1911,N_29245,N_29087);
nor UO_1912 (O_1912,N_28992,N_29499);
nand UO_1913 (O_1913,N_29335,N_29685);
xnor UO_1914 (O_1914,N_29125,N_29887);
xnor UO_1915 (O_1915,N_29784,N_29677);
nand UO_1916 (O_1916,N_29401,N_28835);
nor UO_1917 (O_1917,N_28895,N_29757);
xor UO_1918 (O_1918,N_29836,N_29787);
or UO_1919 (O_1919,N_28958,N_29034);
xor UO_1920 (O_1920,N_28820,N_29649);
and UO_1921 (O_1921,N_29682,N_29746);
xnor UO_1922 (O_1922,N_29802,N_29478);
xnor UO_1923 (O_1923,N_29617,N_29442);
xnor UO_1924 (O_1924,N_29706,N_29237);
and UO_1925 (O_1925,N_29211,N_29217);
or UO_1926 (O_1926,N_29822,N_29785);
or UO_1927 (O_1927,N_28803,N_29548);
or UO_1928 (O_1928,N_28996,N_28862);
and UO_1929 (O_1929,N_29967,N_29529);
nor UO_1930 (O_1930,N_29551,N_29988);
xor UO_1931 (O_1931,N_29461,N_29084);
nor UO_1932 (O_1932,N_29616,N_29387);
or UO_1933 (O_1933,N_29628,N_29384);
nand UO_1934 (O_1934,N_29346,N_29152);
xor UO_1935 (O_1935,N_28841,N_29932);
nand UO_1936 (O_1936,N_29587,N_29668);
nand UO_1937 (O_1937,N_29666,N_28852);
nor UO_1938 (O_1938,N_28908,N_29043);
nor UO_1939 (O_1939,N_29628,N_29205);
nand UO_1940 (O_1940,N_29904,N_29725);
xnor UO_1941 (O_1941,N_29495,N_28984);
or UO_1942 (O_1942,N_29853,N_29912);
or UO_1943 (O_1943,N_29787,N_28877);
xnor UO_1944 (O_1944,N_29845,N_29330);
or UO_1945 (O_1945,N_28908,N_28913);
xnor UO_1946 (O_1946,N_29777,N_29818);
xor UO_1947 (O_1947,N_29125,N_29722);
and UO_1948 (O_1948,N_28830,N_29584);
or UO_1949 (O_1949,N_29548,N_29598);
and UO_1950 (O_1950,N_29976,N_29075);
xnor UO_1951 (O_1951,N_29895,N_29103);
nand UO_1952 (O_1952,N_28935,N_29660);
and UO_1953 (O_1953,N_28851,N_29527);
or UO_1954 (O_1954,N_29955,N_29856);
nand UO_1955 (O_1955,N_29237,N_28806);
or UO_1956 (O_1956,N_29329,N_29365);
and UO_1957 (O_1957,N_28965,N_29377);
xor UO_1958 (O_1958,N_29925,N_29507);
and UO_1959 (O_1959,N_28908,N_29339);
xor UO_1960 (O_1960,N_29967,N_28916);
nand UO_1961 (O_1961,N_29906,N_29858);
xor UO_1962 (O_1962,N_29899,N_29727);
nor UO_1963 (O_1963,N_29411,N_29270);
nand UO_1964 (O_1964,N_28928,N_28889);
or UO_1965 (O_1965,N_28919,N_29829);
nand UO_1966 (O_1966,N_29407,N_29199);
xor UO_1967 (O_1967,N_29949,N_29761);
nand UO_1968 (O_1968,N_29573,N_29702);
nand UO_1969 (O_1969,N_29032,N_29911);
nand UO_1970 (O_1970,N_28867,N_28895);
nand UO_1971 (O_1971,N_29500,N_29466);
and UO_1972 (O_1972,N_29790,N_29083);
nand UO_1973 (O_1973,N_29919,N_29497);
and UO_1974 (O_1974,N_29564,N_29831);
and UO_1975 (O_1975,N_29052,N_29877);
or UO_1976 (O_1976,N_28867,N_29482);
nand UO_1977 (O_1977,N_29723,N_29720);
xnor UO_1978 (O_1978,N_29486,N_29271);
xnor UO_1979 (O_1979,N_29368,N_29812);
nand UO_1980 (O_1980,N_29276,N_28848);
nor UO_1981 (O_1981,N_28998,N_29189);
xor UO_1982 (O_1982,N_28949,N_29608);
and UO_1983 (O_1983,N_29154,N_29382);
xor UO_1984 (O_1984,N_29442,N_28861);
nor UO_1985 (O_1985,N_29897,N_29034);
nand UO_1986 (O_1986,N_29569,N_29160);
and UO_1987 (O_1987,N_29690,N_29948);
or UO_1988 (O_1988,N_29923,N_29983);
nand UO_1989 (O_1989,N_29020,N_29200);
or UO_1990 (O_1990,N_29889,N_29173);
and UO_1991 (O_1991,N_29583,N_29944);
xnor UO_1992 (O_1992,N_29803,N_29331);
nor UO_1993 (O_1993,N_29734,N_28974);
and UO_1994 (O_1994,N_28866,N_28878);
nand UO_1995 (O_1995,N_29799,N_29843);
nor UO_1996 (O_1996,N_29410,N_28872);
and UO_1997 (O_1997,N_29077,N_28839);
and UO_1998 (O_1998,N_29758,N_29683);
nor UO_1999 (O_1999,N_29298,N_29788);
nand UO_2000 (O_2000,N_29535,N_29190);
nand UO_2001 (O_2001,N_29842,N_29955);
xnor UO_2002 (O_2002,N_28956,N_29248);
nand UO_2003 (O_2003,N_29846,N_29663);
or UO_2004 (O_2004,N_29346,N_29020);
nand UO_2005 (O_2005,N_28873,N_29824);
or UO_2006 (O_2006,N_29029,N_28985);
xnor UO_2007 (O_2007,N_29670,N_29243);
xnor UO_2008 (O_2008,N_29505,N_29563);
and UO_2009 (O_2009,N_29681,N_29250);
nor UO_2010 (O_2010,N_29468,N_29675);
nor UO_2011 (O_2011,N_28977,N_29009);
and UO_2012 (O_2012,N_29627,N_29045);
or UO_2013 (O_2013,N_28959,N_29758);
and UO_2014 (O_2014,N_29201,N_29064);
or UO_2015 (O_2015,N_29080,N_29902);
or UO_2016 (O_2016,N_28820,N_28832);
nor UO_2017 (O_2017,N_29618,N_29521);
nor UO_2018 (O_2018,N_28942,N_29923);
or UO_2019 (O_2019,N_29824,N_29062);
xor UO_2020 (O_2020,N_28957,N_29802);
xnor UO_2021 (O_2021,N_28880,N_29424);
nand UO_2022 (O_2022,N_29042,N_28896);
or UO_2023 (O_2023,N_29945,N_29732);
and UO_2024 (O_2024,N_29729,N_29880);
and UO_2025 (O_2025,N_29208,N_28899);
and UO_2026 (O_2026,N_28939,N_29847);
nand UO_2027 (O_2027,N_29869,N_29838);
nor UO_2028 (O_2028,N_29034,N_29601);
and UO_2029 (O_2029,N_29807,N_28856);
xor UO_2030 (O_2030,N_29886,N_29524);
and UO_2031 (O_2031,N_29040,N_29976);
xnor UO_2032 (O_2032,N_29842,N_29853);
nand UO_2033 (O_2033,N_28864,N_29244);
xnor UO_2034 (O_2034,N_29933,N_29814);
or UO_2035 (O_2035,N_29592,N_29508);
or UO_2036 (O_2036,N_29911,N_29112);
nor UO_2037 (O_2037,N_29676,N_29930);
nor UO_2038 (O_2038,N_29559,N_29473);
nand UO_2039 (O_2039,N_29952,N_28809);
or UO_2040 (O_2040,N_29403,N_29299);
xnor UO_2041 (O_2041,N_28866,N_29768);
xor UO_2042 (O_2042,N_29512,N_29660);
nand UO_2043 (O_2043,N_29596,N_29283);
and UO_2044 (O_2044,N_29451,N_29733);
nor UO_2045 (O_2045,N_28826,N_29821);
nor UO_2046 (O_2046,N_29602,N_29263);
nor UO_2047 (O_2047,N_28845,N_29756);
or UO_2048 (O_2048,N_29280,N_29165);
or UO_2049 (O_2049,N_29543,N_29494);
xnor UO_2050 (O_2050,N_29202,N_29418);
and UO_2051 (O_2051,N_29598,N_29434);
xnor UO_2052 (O_2052,N_28990,N_29143);
nand UO_2053 (O_2053,N_29509,N_29117);
nand UO_2054 (O_2054,N_29813,N_28849);
and UO_2055 (O_2055,N_29495,N_29386);
nor UO_2056 (O_2056,N_29508,N_28855);
nand UO_2057 (O_2057,N_29702,N_28981);
nor UO_2058 (O_2058,N_29556,N_29688);
nand UO_2059 (O_2059,N_29245,N_29933);
nor UO_2060 (O_2060,N_29216,N_29973);
or UO_2061 (O_2061,N_29976,N_29837);
or UO_2062 (O_2062,N_29180,N_29869);
nor UO_2063 (O_2063,N_29337,N_29871);
nor UO_2064 (O_2064,N_29351,N_29825);
nand UO_2065 (O_2065,N_29320,N_28823);
and UO_2066 (O_2066,N_29800,N_28859);
xor UO_2067 (O_2067,N_29171,N_28924);
nor UO_2068 (O_2068,N_29448,N_29670);
or UO_2069 (O_2069,N_28828,N_28900);
nand UO_2070 (O_2070,N_29192,N_29778);
nor UO_2071 (O_2071,N_29837,N_29167);
nand UO_2072 (O_2072,N_29543,N_29833);
xor UO_2073 (O_2073,N_29589,N_29122);
or UO_2074 (O_2074,N_29740,N_29574);
nor UO_2075 (O_2075,N_28955,N_29922);
nor UO_2076 (O_2076,N_29773,N_29440);
nor UO_2077 (O_2077,N_29862,N_29969);
and UO_2078 (O_2078,N_29219,N_29352);
xnor UO_2079 (O_2079,N_29596,N_29197);
xnor UO_2080 (O_2080,N_29286,N_29925);
or UO_2081 (O_2081,N_29941,N_29063);
nand UO_2082 (O_2082,N_29738,N_28865);
or UO_2083 (O_2083,N_28918,N_28822);
nor UO_2084 (O_2084,N_29105,N_29343);
and UO_2085 (O_2085,N_29011,N_29176);
and UO_2086 (O_2086,N_29033,N_29479);
nand UO_2087 (O_2087,N_28948,N_29195);
xnor UO_2088 (O_2088,N_29155,N_29391);
and UO_2089 (O_2089,N_29117,N_28967);
xnor UO_2090 (O_2090,N_29135,N_29128);
nand UO_2091 (O_2091,N_29016,N_29960);
xnor UO_2092 (O_2092,N_28959,N_29005);
xor UO_2093 (O_2093,N_28956,N_29117);
nand UO_2094 (O_2094,N_29250,N_29452);
or UO_2095 (O_2095,N_29130,N_29244);
xnor UO_2096 (O_2096,N_29591,N_29862);
nand UO_2097 (O_2097,N_29321,N_29714);
nor UO_2098 (O_2098,N_28837,N_29326);
xor UO_2099 (O_2099,N_29627,N_28806);
or UO_2100 (O_2100,N_28942,N_29948);
xnor UO_2101 (O_2101,N_29480,N_29117);
nand UO_2102 (O_2102,N_29143,N_29094);
and UO_2103 (O_2103,N_29384,N_29072);
nand UO_2104 (O_2104,N_29585,N_29816);
xor UO_2105 (O_2105,N_29937,N_29992);
xor UO_2106 (O_2106,N_29939,N_29143);
or UO_2107 (O_2107,N_29975,N_29976);
nor UO_2108 (O_2108,N_29690,N_29029);
nand UO_2109 (O_2109,N_29139,N_29867);
xor UO_2110 (O_2110,N_29666,N_29094);
and UO_2111 (O_2111,N_29989,N_28975);
xor UO_2112 (O_2112,N_29607,N_29688);
or UO_2113 (O_2113,N_29111,N_29616);
xnor UO_2114 (O_2114,N_28826,N_29873);
and UO_2115 (O_2115,N_29674,N_29779);
and UO_2116 (O_2116,N_29300,N_29485);
nor UO_2117 (O_2117,N_28983,N_29185);
xor UO_2118 (O_2118,N_29971,N_29998);
nand UO_2119 (O_2119,N_29028,N_29222);
or UO_2120 (O_2120,N_29794,N_29395);
xnor UO_2121 (O_2121,N_29387,N_28911);
or UO_2122 (O_2122,N_29146,N_29136);
xnor UO_2123 (O_2123,N_29662,N_28893);
nand UO_2124 (O_2124,N_29807,N_29212);
and UO_2125 (O_2125,N_29309,N_29538);
nor UO_2126 (O_2126,N_29606,N_29909);
xnor UO_2127 (O_2127,N_29446,N_29823);
nor UO_2128 (O_2128,N_29933,N_29472);
and UO_2129 (O_2129,N_29242,N_29959);
nand UO_2130 (O_2130,N_29994,N_29161);
xor UO_2131 (O_2131,N_29076,N_29846);
nor UO_2132 (O_2132,N_29431,N_29523);
nand UO_2133 (O_2133,N_29917,N_28958);
nand UO_2134 (O_2134,N_29865,N_29576);
nand UO_2135 (O_2135,N_29479,N_29806);
nor UO_2136 (O_2136,N_28896,N_29475);
nand UO_2137 (O_2137,N_29757,N_29726);
nand UO_2138 (O_2138,N_29241,N_29300);
nand UO_2139 (O_2139,N_29732,N_29601);
or UO_2140 (O_2140,N_29102,N_29525);
and UO_2141 (O_2141,N_29811,N_29115);
xor UO_2142 (O_2142,N_29312,N_29449);
xnor UO_2143 (O_2143,N_29339,N_29517);
and UO_2144 (O_2144,N_29155,N_29583);
nand UO_2145 (O_2145,N_29455,N_28861);
xnor UO_2146 (O_2146,N_29036,N_29188);
or UO_2147 (O_2147,N_29074,N_29044);
nand UO_2148 (O_2148,N_29896,N_29474);
and UO_2149 (O_2149,N_29242,N_29907);
and UO_2150 (O_2150,N_29742,N_29288);
and UO_2151 (O_2151,N_29979,N_29840);
and UO_2152 (O_2152,N_29686,N_29055);
xnor UO_2153 (O_2153,N_29545,N_28820);
xnor UO_2154 (O_2154,N_28904,N_29787);
nor UO_2155 (O_2155,N_29873,N_29693);
and UO_2156 (O_2156,N_29823,N_29843);
xnor UO_2157 (O_2157,N_29687,N_29926);
or UO_2158 (O_2158,N_29909,N_29901);
or UO_2159 (O_2159,N_29105,N_29256);
nand UO_2160 (O_2160,N_29344,N_29254);
and UO_2161 (O_2161,N_29275,N_29520);
and UO_2162 (O_2162,N_29510,N_29223);
and UO_2163 (O_2163,N_29589,N_29842);
or UO_2164 (O_2164,N_29289,N_29555);
nor UO_2165 (O_2165,N_28827,N_29679);
xnor UO_2166 (O_2166,N_29087,N_29136);
xnor UO_2167 (O_2167,N_29112,N_29854);
and UO_2168 (O_2168,N_29277,N_29340);
nor UO_2169 (O_2169,N_28859,N_29090);
nor UO_2170 (O_2170,N_29878,N_29648);
nor UO_2171 (O_2171,N_29353,N_29036);
nor UO_2172 (O_2172,N_29810,N_29685);
or UO_2173 (O_2173,N_29440,N_29568);
or UO_2174 (O_2174,N_29825,N_28844);
or UO_2175 (O_2175,N_29973,N_29564);
xnor UO_2176 (O_2176,N_29233,N_29229);
or UO_2177 (O_2177,N_29489,N_29731);
nand UO_2178 (O_2178,N_29481,N_29393);
and UO_2179 (O_2179,N_29909,N_29255);
and UO_2180 (O_2180,N_29998,N_29718);
and UO_2181 (O_2181,N_29160,N_29186);
nor UO_2182 (O_2182,N_28849,N_29383);
nand UO_2183 (O_2183,N_29992,N_29791);
or UO_2184 (O_2184,N_29810,N_28927);
nor UO_2185 (O_2185,N_29192,N_29417);
or UO_2186 (O_2186,N_29596,N_29625);
nor UO_2187 (O_2187,N_29782,N_28985);
or UO_2188 (O_2188,N_29696,N_29620);
nand UO_2189 (O_2189,N_28953,N_28901);
nor UO_2190 (O_2190,N_29650,N_29317);
or UO_2191 (O_2191,N_29046,N_29010);
nor UO_2192 (O_2192,N_29524,N_29188);
nor UO_2193 (O_2193,N_29866,N_29490);
nor UO_2194 (O_2194,N_29483,N_28983);
nor UO_2195 (O_2195,N_29844,N_29259);
and UO_2196 (O_2196,N_29408,N_29344);
or UO_2197 (O_2197,N_28962,N_29947);
or UO_2198 (O_2198,N_29393,N_29343);
nor UO_2199 (O_2199,N_29190,N_29715);
xor UO_2200 (O_2200,N_29272,N_29413);
nor UO_2201 (O_2201,N_29925,N_29534);
nand UO_2202 (O_2202,N_29612,N_29308);
and UO_2203 (O_2203,N_29668,N_29128);
xnor UO_2204 (O_2204,N_29653,N_29233);
xnor UO_2205 (O_2205,N_29120,N_29579);
nor UO_2206 (O_2206,N_29234,N_29716);
and UO_2207 (O_2207,N_29143,N_29368);
and UO_2208 (O_2208,N_29173,N_29462);
or UO_2209 (O_2209,N_29864,N_29156);
and UO_2210 (O_2210,N_29087,N_29715);
xnor UO_2211 (O_2211,N_29214,N_29021);
nor UO_2212 (O_2212,N_29643,N_29688);
nor UO_2213 (O_2213,N_29906,N_29260);
and UO_2214 (O_2214,N_29313,N_29191);
xor UO_2215 (O_2215,N_29822,N_29881);
nor UO_2216 (O_2216,N_28991,N_29111);
xnor UO_2217 (O_2217,N_29757,N_29579);
nor UO_2218 (O_2218,N_29408,N_29089);
nor UO_2219 (O_2219,N_29239,N_28833);
nor UO_2220 (O_2220,N_29974,N_29834);
or UO_2221 (O_2221,N_28875,N_28942);
or UO_2222 (O_2222,N_28916,N_29494);
nand UO_2223 (O_2223,N_29577,N_29966);
nand UO_2224 (O_2224,N_29588,N_29668);
and UO_2225 (O_2225,N_29004,N_29337);
xor UO_2226 (O_2226,N_29864,N_29196);
xnor UO_2227 (O_2227,N_29803,N_28893);
and UO_2228 (O_2228,N_29701,N_29946);
xor UO_2229 (O_2229,N_28912,N_29150);
nand UO_2230 (O_2230,N_29638,N_29179);
or UO_2231 (O_2231,N_29122,N_29314);
and UO_2232 (O_2232,N_29565,N_29628);
nand UO_2233 (O_2233,N_29071,N_29818);
and UO_2234 (O_2234,N_29318,N_29462);
and UO_2235 (O_2235,N_29820,N_28919);
nor UO_2236 (O_2236,N_28954,N_29600);
nand UO_2237 (O_2237,N_29895,N_29275);
and UO_2238 (O_2238,N_29412,N_29437);
nand UO_2239 (O_2239,N_29578,N_29697);
nor UO_2240 (O_2240,N_28995,N_29891);
or UO_2241 (O_2241,N_28801,N_29685);
nor UO_2242 (O_2242,N_29362,N_28989);
nand UO_2243 (O_2243,N_28987,N_29203);
nor UO_2244 (O_2244,N_29273,N_29215);
or UO_2245 (O_2245,N_28898,N_29947);
xor UO_2246 (O_2246,N_28906,N_29934);
nand UO_2247 (O_2247,N_29397,N_29981);
or UO_2248 (O_2248,N_29642,N_29985);
xor UO_2249 (O_2249,N_29503,N_29990);
nor UO_2250 (O_2250,N_29037,N_28851);
xnor UO_2251 (O_2251,N_29791,N_28917);
nand UO_2252 (O_2252,N_29830,N_28829);
or UO_2253 (O_2253,N_29818,N_29863);
and UO_2254 (O_2254,N_29664,N_29457);
xnor UO_2255 (O_2255,N_29164,N_29327);
xor UO_2256 (O_2256,N_29428,N_28897);
nor UO_2257 (O_2257,N_29480,N_29152);
xnor UO_2258 (O_2258,N_29464,N_29692);
nand UO_2259 (O_2259,N_29503,N_29327);
xnor UO_2260 (O_2260,N_29875,N_29601);
nor UO_2261 (O_2261,N_28806,N_29904);
nor UO_2262 (O_2262,N_28991,N_29762);
or UO_2263 (O_2263,N_29974,N_29264);
xor UO_2264 (O_2264,N_29797,N_29071);
nand UO_2265 (O_2265,N_29722,N_29119);
xnor UO_2266 (O_2266,N_29506,N_29782);
and UO_2267 (O_2267,N_29544,N_29956);
nand UO_2268 (O_2268,N_29692,N_29183);
xor UO_2269 (O_2269,N_29734,N_29383);
and UO_2270 (O_2270,N_28988,N_29559);
nor UO_2271 (O_2271,N_29737,N_29587);
nand UO_2272 (O_2272,N_29445,N_29925);
nor UO_2273 (O_2273,N_29495,N_29432);
nor UO_2274 (O_2274,N_29831,N_29279);
and UO_2275 (O_2275,N_29297,N_28910);
and UO_2276 (O_2276,N_29265,N_29261);
nor UO_2277 (O_2277,N_29526,N_29478);
xnor UO_2278 (O_2278,N_29352,N_28858);
nand UO_2279 (O_2279,N_29144,N_28810);
nor UO_2280 (O_2280,N_28856,N_29845);
or UO_2281 (O_2281,N_29644,N_29085);
xnor UO_2282 (O_2282,N_29945,N_29545);
and UO_2283 (O_2283,N_29216,N_29369);
nand UO_2284 (O_2284,N_28810,N_28904);
xor UO_2285 (O_2285,N_29323,N_29522);
nor UO_2286 (O_2286,N_28840,N_28877);
xor UO_2287 (O_2287,N_29803,N_29504);
or UO_2288 (O_2288,N_29559,N_29099);
and UO_2289 (O_2289,N_29791,N_28985);
and UO_2290 (O_2290,N_29906,N_29370);
nor UO_2291 (O_2291,N_29357,N_29254);
nand UO_2292 (O_2292,N_29021,N_29136);
or UO_2293 (O_2293,N_29848,N_28865);
nand UO_2294 (O_2294,N_28840,N_28891);
nor UO_2295 (O_2295,N_28986,N_29967);
and UO_2296 (O_2296,N_29338,N_29656);
xor UO_2297 (O_2297,N_28857,N_29538);
nor UO_2298 (O_2298,N_29966,N_29594);
xnor UO_2299 (O_2299,N_29358,N_29750);
nand UO_2300 (O_2300,N_29569,N_29553);
and UO_2301 (O_2301,N_29870,N_29768);
nor UO_2302 (O_2302,N_29118,N_29754);
nand UO_2303 (O_2303,N_29171,N_29709);
and UO_2304 (O_2304,N_29681,N_29257);
xor UO_2305 (O_2305,N_29446,N_28912);
nand UO_2306 (O_2306,N_29799,N_29815);
nor UO_2307 (O_2307,N_29316,N_29018);
nand UO_2308 (O_2308,N_29863,N_29905);
nor UO_2309 (O_2309,N_29236,N_29652);
or UO_2310 (O_2310,N_29418,N_29005);
and UO_2311 (O_2311,N_29161,N_28997);
and UO_2312 (O_2312,N_29462,N_29977);
or UO_2313 (O_2313,N_29160,N_29559);
and UO_2314 (O_2314,N_29473,N_29953);
or UO_2315 (O_2315,N_29716,N_29604);
or UO_2316 (O_2316,N_29244,N_29088);
or UO_2317 (O_2317,N_29102,N_29168);
nand UO_2318 (O_2318,N_29695,N_29663);
and UO_2319 (O_2319,N_28866,N_29338);
nand UO_2320 (O_2320,N_28882,N_29676);
nor UO_2321 (O_2321,N_28925,N_28821);
nor UO_2322 (O_2322,N_29913,N_29274);
and UO_2323 (O_2323,N_29135,N_29924);
and UO_2324 (O_2324,N_29180,N_28831);
nand UO_2325 (O_2325,N_29036,N_29085);
xor UO_2326 (O_2326,N_29552,N_29387);
and UO_2327 (O_2327,N_29482,N_29701);
or UO_2328 (O_2328,N_28896,N_29810);
nor UO_2329 (O_2329,N_29700,N_29584);
and UO_2330 (O_2330,N_29095,N_29446);
and UO_2331 (O_2331,N_29349,N_29974);
or UO_2332 (O_2332,N_29161,N_29447);
and UO_2333 (O_2333,N_29360,N_29714);
or UO_2334 (O_2334,N_29856,N_29036);
or UO_2335 (O_2335,N_29468,N_29543);
and UO_2336 (O_2336,N_29253,N_28899);
or UO_2337 (O_2337,N_29789,N_29819);
and UO_2338 (O_2338,N_29711,N_28975);
nand UO_2339 (O_2339,N_29405,N_29180);
and UO_2340 (O_2340,N_29803,N_29862);
xor UO_2341 (O_2341,N_29057,N_29202);
xor UO_2342 (O_2342,N_29647,N_29822);
xor UO_2343 (O_2343,N_29458,N_29359);
xnor UO_2344 (O_2344,N_29137,N_28832);
nor UO_2345 (O_2345,N_29031,N_29421);
nand UO_2346 (O_2346,N_29450,N_28897);
nor UO_2347 (O_2347,N_29436,N_29141);
nor UO_2348 (O_2348,N_29470,N_28926);
and UO_2349 (O_2349,N_29389,N_29261);
or UO_2350 (O_2350,N_29327,N_29134);
nor UO_2351 (O_2351,N_28997,N_29026);
or UO_2352 (O_2352,N_29848,N_28978);
nor UO_2353 (O_2353,N_28951,N_29788);
nor UO_2354 (O_2354,N_29885,N_29444);
or UO_2355 (O_2355,N_29009,N_28882);
nand UO_2356 (O_2356,N_29357,N_29039);
nand UO_2357 (O_2357,N_28828,N_29758);
nor UO_2358 (O_2358,N_28875,N_29658);
nand UO_2359 (O_2359,N_29619,N_29672);
and UO_2360 (O_2360,N_28871,N_29158);
nor UO_2361 (O_2361,N_29605,N_29115);
nand UO_2362 (O_2362,N_29160,N_29831);
or UO_2363 (O_2363,N_28876,N_29252);
nor UO_2364 (O_2364,N_29909,N_29581);
nand UO_2365 (O_2365,N_29337,N_28927);
or UO_2366 (O_2366,N_29151,N_29752);
nor UO_2367 (O_2367,N_29134,N_28876);
xnor UO_2368 (O_2368,N_29137,N_29515);
xor UO_2369 (O_2369,N_29185,N_29664);
nor UO_2370 (O_2370,N_29021,N_29038);
or UO_2371 (O_2371,N_29454,N_29747);
or UO_2372 (O_2372,N_29193,N_29159);
xnor UO_2373 (O_2373,N_29472,N_29199);
nand UO_2374 (O_2374,N_29257,N_28962);
nand UO_2375 (O_2375,N_29211,N_29059);
nand UO_2376 (O_2376,N_28964,N_28876);
nor UO_2377 (O_2377,N_29986,N_29267);
nand UO_2378 (O_2378,N_29743,N_29136);
and UO_2379 (O_2379,N_29488,N_29837);
nand UO_2380 (O_2380,N_29551,N_29250);
or UO_2381 (O_2381,N_29991,N_29271);
nand UO_2382 (O_2382,N_29857,N_29718);
and UO_2383 (O_2383,N_29166,N_29383);
nor UO_2384 (O_2384,N_29660,N_29582);
nand UO_2385 (O_2385,N_29164,N_28977);
xnor UO_2386 (O_2386,N_29178,N_28932);
nor UO_2387 (O_2387,N_29658,N_29356);
xor UO_2388 (O_2388,N_29949,N_28914);
nor UO_2389 (O_2389,N_29803,N_29375);
and UO_2390 (O_2390,N_29597,N_29107);
nand UO_2391 (O_2391,N_29072,N_29125);
or UO_2392 (O_2392,N_29159,N_29801);
and UO_2393 (O_2393,N_29416,N_29760);
nand UO_2394 (O_2394,N_29065,N_28910);
xnor UO_2395 (O_2395,N_29286,N_29273);
or UO_2396 (O_2396,N_29829,N_28828);
nor UO_2397 (O_2397,N_29982,N_29894);
and UO_2398 (O_2398,N_29608,N_28826);
nand UO_2399 (O_2399,N_29992,N_29254);
nand UO_2400 (O_2400,N_29570,N_29152);
and UO_2401 (O_2401,N_29408,N_29240);
nand UO_2402 (O_2402,N_29085,N_29066);
or UO_2403 (O_2403,N_29069,N_28832);
or UO_2404 (O_2404,N_28977,N_29674);
nand UO_2405 (O_2405,N_29282,N_29129);
nand UO_2406 (O_2406,N_29322,N_28834);
nor UO_2407 (O_2407,N_29454,N_29109);
or UO_2408 (O_2408,N_29245,N_29240);
or UO_2409 (O_2409,N_29453,N_28981);
nor UO_2410 (O_2410,N_29023,N_29404);
nand UO_2411 (O_2411,N_28823,N_28867);
or UO_2412 (O_2412,N_29460,N_28976);
nand UO_2413 (O_2413,N_28836,N_29989);
nor UO_2414 (O_2414,N_29948,N_29414);
nor UO_2415 (O_2415,N_29180,N_29349);
xor UO_2416 (O_2416,N_29779,N_29130);
nor UO_2417 (O_2417,N_29637,N_29536);
nand UO_2418 (O_2418,N_29704,N_28854);
xnor UO_2419 (O_2419,N_29394,N_29519);
or UO_2420 (O_2420,N_29776,N_29956);
xnor UO_2421 (O_2421,N_29808,N_29688);
or UO_2422 (O_2422,N_29252,N_29364);
or UO_2423 (O_2423,N_28966,N_28950);
or UO_2424 (O_2424,N_28832,N_29054);
or UO_2425 (O_2425,N_29163,N_29820);
or UO_2426 (O_2426,N_29838,N_29105);
nor UO_2427 (O_2427,N_29560,N_29792);
xnor UO_2428 (O_2428,N_29161,N_29694);
nor UO_2429 (O_2429,N_29647,N_28964);
nand UO_2430 (O_2430,N_29455,N_29299);
xnor UO_2431 (O_2431,N_29275,N_29991);
or UO_2432 (O_2432,N_29636,N_29131);
nor UO_2433 (O_2433,N_29168,N_29317);
nor UO_2434 (O_2434,N_29864,N_29958);
nand UO_2435 (O_2435,N_29348,N_29884);
nor UO_2436 (O_2436,N_29402,N_29178);
nand UO_2437 (O_2437,N_29965,N_29598);
or UO_2438 (O_2438,N_29999,N_29499);
xor UO_2439 (O_2439,N_28997,N_29234);
or UO_2440 (O_2440,N_29189,N_29955);
nand UO_2441 (O_2441,N_29983,N_29986);
nor UO_2442 (O_2442,N_28853,N_29022);
nor UO_2443 (O_2443,N_29103,N_29029);
nand UO_2444 (O_2444,N_29933,N_29905);
nor UO_2445 (O_2445,N_29848,N_29062);
or UO_2446 (O_2446,N_29294,N_29361);
nand UO_2447 (O_2447,N_28805,N_29554);
or UO_2448 (O_2448,N_29174,N_28866);
or UO_2449 (O_2449,N_29880,N_29341);
nor UO_2450 (O_2450,N_29169,N_29501);
xor UO_2451 (O_2451,N_29144,N_29323);
or UO_2452 (O_2452,N_29151,N_29903);
and UO_2453 (O_2453,N_28945,N_29965);
nor UO_2454 (O_2454,N_29116,N_29850);
nor UO_2455 (O_2455,N_29845,N_29833);
xor UO_2456 (O_2456,N_29330,N_28976);
nand UO_2457 (O_2457,N_29799,N_29267);
nor UO_2458 (O_2458,N_29837,N_28865);
nor UO_2459 (O_2459,N_29664,N_29227);
xor UO_2460 (O_2460,N_29318,N_29532);
and UO_2461 (O_2461,N_29240,N_29798);
and UO_2462 (O_2462,N_29169,N_29232);
and UO_2463 (O_2463,N_29226,N_29371);
and UO_2464 (O_2464,N_29529,N_29745);
nor UO_2465 (O_2465,N_29269,N_29983);
nor UO_2466 (O_2466,N_29400,N_29434);
nor UO_2467 (O_2467,N_29649,N_29972);
nand UO_2468 (O_2468,N_29727,N_28976);
xor UO_2469 (O_2469,N_29479,N_29821);
and UO_2470 (O_2470,N_29404,N_29005);
and UO_2471 (O_2471,N_29072,N_29584);
nand UO_2472 (O_2472,N_29753,N_29370);
and UO_2473 (O_2473,N_29442,N_29352);
nor UO_2474 (O_2474,N_29906,N_29384);
and UO_2475 (O_2475,N_29119,N_28824);
or UO_2476 (O_2476,N_29460,N_28979);
nor UO_2477 (O_2477,N_29668,N_29608);
and UO_2478 (O_2478,N_29212,N_29615);
or UO_2479 (O_2479,N_29290,N_29627);
and UO_2480 (O_2480,N_29767,N_29630);
or UO_2481 (O_2481,N_29144,N_29862);
and UO_2482 (O_2482,N_28932,N_29615);
and UO_2483 (O_2483,N_29986,N_29277);
and UO_2484 (O_2484,N_28977,N_29569);
and UO_2485 (O_2485,N_29161,N_29904);
nand UO_2486 (O_2486,N_29589,N_29924);
nand UO_2487 (O_2487,N_29326,N_29650);
nor UO_2488 (O_2488,N_29228,N_29316);
and UO_2489 (O_2489,N_29931,N_29389);
xnor UO_2490 (O_2490,N_29942,N_29557);
nand UO_2491 (O_2491,N_29906,N_29466);
or UO_2492 (O_2492,N_29637,N_29988);
xor UO_2493 (O_2493,N_29211,N_29714);
or UO_2494 (O_2494,N_29182,N_29966);
and UO_2495 (O_2495,N_29085,N_28888);
nor UO_2496 (O_2496,N_29249,N_29226);
or UO_2497 (O_2497,N_29909,N_29322);
nand UO_2498 (O_2498,N_29718,N_29644);
or UO_2499 (O_2499,N_29172,N_29100);
or UO_2500 (O_2500,N_28839,N_29442);
or UO_2501 (O_2501,N_28942,N_29074);
or UO_2502 (O_2502,N_29951,N_28905);
nor UO_2503 (O_2503,N_29891,N_28934);
and UO_2504 (O_2504,N_29808,N_29497);
and UO_2505 (O_2505,N_29763,N_29690);
xnor UO_2506 (O_2506,N_28835,N_29302);
xor UO_2507 (O_2507,N_29243,N_29097);
nand UO_2508 (O_2508,N_29619,N_29606);
nor UO_2509 (O_2509,N_29621,N_29006);
xnor UO_2510 (O_2510,N_29350,N_29805);
and UO_2511 (O_2511,N_29617,N_29706);
or UO_2512 (O_2512,N_29517,N_29381);
xnor UO_2513 (O_2513,N_28956,N_29541);
nand UO_2514 (O_2514,N_28998,N_29281);
and UO_2515 (O_2515,N_29453,N_29379);
or UO_2516 (O_2516,N_29212,N_29127);
or UO_2517 (O_2517,N_29795,N_29782);
nor UO_2518 (O_2518,N_29460,N_29328);
nor UO_2519 (O_2519,N_29328,N_29671);
nand UO_2520 (O_2520,N_29272,N_29376);
nand UO_2521 (O_2521,N_29346,N_29455);
and UO_2522 (O_2522,N_29865,N_29006);
nand UO_2523 (O_2523,N_29240,N_29402);
nand UO_2524 (O_2524,N_29585,N_29103);
nor UO_2525 (O_2525,N_29859,N_29050);
and UO_2526 (O_2526,N_29285,N_29052);
or UO_2527 (O_2527,N_29586,N_29873);
xor UO_2528 (O_2528,N_29062,N_28912);
nor UO_2529 (O_2529,N_29773,N_29902);
nor UO_2530 (O_2530,N_29382,N_29160);
or UO_2531 (O_2531,N_29614,N_29737);
xnor UO_2532 (O_2532,N_29859,N_29950);
xnor UO_2533 (O_2533,N_29180,N_29520);
or UO_2534 (O_2534,N_29587,N_29130);
and UO_2535 (O_2535,N_28818,N_29894);
or UO_2536 (O_2536,N_29866,N_29269);
or UO_2537 (O_2537,N_29047,N_29945);
xor UO_2538 (O_2538,N_29297,N_29459);
nand UO_2539 (O_2539,N_29913,N_29586);
and UO_2540 (O_2540,N_29446,N_29897);
nand UO_2541 (O_2541,N_29283,N_28929);
nor UO_2542 (O_2542,N_29969,N_29441);
or UO_2543 (O_2543,N_29730,N_29296);
nor UO_2544 (O_2544,N_29970,N_28812);
or UO_2545 (O_2545,N_29069,N_29577);
nand UO_2546 (O_2546,N_29883,N_29145);
nor UO_2547 (O_2547,N_29168,N_29149);
nor UO_2548 (O_2548,N_29469,N_29905);
or UO_2549 (O_2549,N_28827,N_29387);
or UO_2550 (O_2550,N_29072,N_29664);
xor UO_2551 (O_2551,N_29886,N_29287);
xnor UO_2552 (O_2552,N_29668,N_29152);
xnor UO_2553 (O_2553,N_29672,N_29478);
nand UO_2554 (O_2554,N_29494,N_29134);
nand UO_2555 (O_2555,N_29742,N_28897);
nor UO_2556 (O_2556,N_29754,N_29220);
xor UO_2557 (O_2557,N_29762,N_29940);
xnor UO_2558 (O_2558,N_29489,N_29106);
nor UO_2559 (O_2559,N_29356,N_29493);
nor UO_2560 (O_2560,N_29400,N_28849);
nand UO_2561 (O_2561,N_28898,N_29907);
nor UO_2562 (O_2562,N_28837,N_29065);
nor UO_2563 (O_2563,N_28883,N_29135);
nor UO_2564 (O_2564,N_29640,N_29177);
nor UO_2565 (O_2565,N_29680,N_29217);
nor UO_2566 (O_2566,N_29788,N_29718);
and UO_2567 (O_2567,N_29445,N_28941);
and UO_2568 (O_2568,N_29171,N_28828);
nor UO_2569 (O_2569,N_29169,N_29874);
nor UO_2570 (O_2570,N_28946,N_29576);
nor UO_2571 (O_2571,N_29312,N_29873);
xnor UO_2572 (O_2572,N_28826,N_28805);
nor UO_2573 (O_2573,N_29147,N_29018);
xnor UO_2574 (O_2574,N_28904,N_29665);
nand UO_2575 (O_2575,N_29262,N_29217);
or UO_2576 (O_2576,N_29430,N_29720);
xnor UO_2577 (O_2577,N_28946,N_29587);
or UO_2578 (O_2578,N_28964,N_29461);
nand UO_2579 (O_2579,N_29980,N_29532);
or UO_2580 (O_2580,N_29416,N_29474);
and UO_2581 (O_2581,N_29918,N_29848);
or UO_2582 (O_2582,N_29334,N_29800);
or UO_2583 (O_2583,N_28880,N_29466);
nand UO_2584 (O_2584,N_29641,N_29549);
xor UO_2585 (O_2585,N_29628,N_29408);
xnor UO_2586 (O_2586,N_29649,N_29609);
and UO_2587 (O_2587,N_29104,N_29495);
or UO_2588 (O_2588,N_29824,N_29846);
xor UO_2589 (O_2589,N_28948,N_29806);
xnor UO_2590 (O_2590,N_29400,N_29150);
nand UO_2591 (O_2591,N_29081,N_29984);
nor UO_2592 (O_2592,N_28804,N_28821);
and UO_2593 (O_2593,N_29378,N_28949);
or UO_2594 (O_2594,N_29770,N_29975);
nand UO_2595 (O_2595,N_29392,N_29318);
xnor UO_2596 (O_2596,N_29349,N_29554);
or UO_2597 (O_2597,N_29399,N_28875);
xnor UO_2598 (O_2598,N_29614,N_29152);
or UO_2599 (O_2599,N_29805,N_29835);
nand UO_2600 (O_2600,N_29996,N_29170);
xor UO_2601 (O_2601,N_29169,N_29085);
and UO_2602 (O_2602,N_29720,N_29034);
or UO_2603 (O_2603,N_29380,N_29917);
nor UO_2604 (O_2604,N_29027,N_29373);
or UO_2605 (O_2605,N_29910,N_29916);
nand UO_2606 (O_2606,N_29794,N_29434);
xnor UO_2607 (O_2607,N_29185,N_29169);
or UO_2608 (O_2608,N_29699,N_29422);
xor UO_2609 (O_2609,N_29945,N_29976);
nand UO_2610 (O_2610,N_29992,N_28835);
and UO_2611 (O_2611,N_29930,N_29201);
nand UO_2612 (O_2612,N_29888,N_29864);
nand UO_2613 (O_2613,N_29564,N_29594);
or UO_2614 (O_2614,N_29433,N_29893);
xor UO_2615 (O_2615,N_29435,N_28829);
and UO_2616 (O_2616,N_28822,N_28920);
and UO_2617 (O_2617,N_29690,N_29953);
and UO_2618 (O_2618,N_29178,N_28904);
or UO_2619 (O_2619,N_29163,N_29750);
xnor UO_2620 (O_2620,N_29996,N_28965);
and UO_2621 (O_2621,N_29342,N_29610);
or UO_2622 (O_2622,N_29515,N_29319);
nand UO_2623 (O_2623,N_29641,N_29319);
xor UO_2624 (O_2624,N_28807,N_29727);
xor UO_2625 (O_2625,N_28822,N_29755);
nor UO_2626 (O_2626,N_29035,N_28853);
xnor UO_2627 (O_2627,N_29131,N_29482);
xor UO_2628 (O_2628,N_29707,N_29555);
nand UO_2629 (O_2629,N_29873,N_29352);
nor UO_2630 (O_2630,N_29070,N_29543);
or UO_2631 (O_2631,N_29189,N_28907);
nor UO_2632 (O_2632,N_29886,N_29347);
and UO_2633 (O_2633,N_29189,N_29687);
or UO_2634 (O_2634,N_29712,N_29461);
xnor UO_2635 (O_2635,N_29682,N_29769);
nand UO_2636 (O_2636,N_29324,N_29873);
and UO_2637 (O_2637,N_29200,N_29565);
and UO_2638 (O_2638,N_29473,N_29736);
nand UO_2639 (O_2639,N_29071,N_29483);
nand UO_2640 (O_2640,N_29972,N_28844);
xnor UO_2641 (O_2641,N_29941,N_28932);
nand UO_2642 (O_2642,N_29526,N_29123);
or UO_2643 (O_2643,N_29043,N_29542);
or UO_2644 (O_2644,N_29811,N_29985);
or UO_2645 (O_2645,N_29692,N_29818);
and UO_2646 (O_2646,N_29889,N_29965);
nand UO_2647 (O_2647,N_29652,N_29422);
and UO_2648 (O_2648,N_29688,N_29152);
nor UO_2649 (O_2649,N_29231,N_28907);
xnor UO_2650 (O_2650,N_29610,N_29523);
nor UO_2651 (O_2651,N_29611,N_28831);
nor UO_2652 (O_2652,N_29498,N_29856);
or UO_2653 (O_2653,N_29827,N_29899);
nor UO_2654 (O_2654,N_29703,N_29905);
or UO_2655 (O_2655,N_29016,N_29010);
nor UO_2656 (O_2656,N_29813,N_29975);
nand UO_2657 (O_2657,N_28852,N_29971);
xor UO_2658 (O_2658,N_29765,N_29005);
or UO_2659 (O_2659,N_29613,N_29750);
nor UO_2660 (O_2660,N_29680,N_28944);
nand UO_2661 (O_2661,N_29839,N_28949);
nand UO_2662 (O_2662,N_29331,N_29680);
xnor UO_2663 (O_2663,N_29161,N_28889);
or UO_2664 (O_2664,N_28950,N_28948);
and UO_2665 (O_2665,N_29167,N_29653);
or UO_2666 (O_2666,N_29730,N_28982);
nor UO_2667 (O_2667,N_28960,N_29880);
nand UO_2668 (O_2668,N_29477,N_29177);
nor UO_2669 (O_2669,N_29968,N_29637);
and UO_2670 (O_2670,N_29600,N_29030);
and UO_2671 (O_2671,N_29852,N_29316);
nor UO_2672 (O_2672,N_29443,N_29235);
and UO_2673 (O_2673,N_29468,N_28821);
nand UO_2674 (O_2674,N_29487,N_29161);
or UO_2675 (O_2675,N_29236,N_29293);
or UO_2676 (O_2676,N_29206,N_28990);
xor UO_2677 (O_2677,N_29600,N_28919);
xnor UO_2678 (O_2678,N_29604,N_29646);
nor UO_2679 (O_2679,N_29197,N_28918);
or UO_2680 (O_2680,N_29414,N_29185);
or UO_2681 (O_2681,N_29923,N_29186);
and UO_2682 (O_2682,N_29193,N_29627);
and UO_2683 (O_2683,N_28826,N_29448);
nand UO_2684 (O_2684,N_29903,N_29253);
and UO_2685 (O_2685,N_29697,N_29020);
and UO_2686 (O_2686,N_28845,N_29827);
or UO_2687 (O_2687,N_28896,N_29064);
nor UO_2688 (O_2688,N_28921,N_28881);
nand UO_2689 (O_2689,N_29375,N_29308);
nor UO_2690 (O_2690,N_28810,N_29555);
nor UO_2691 (O_2691,N_29431,N_29185);
xnor UO_2692 (O_2692,N_28833,N_28931);
xnor UO_2693 (O_2693,N_28904,N_29934);
nor UO_2694 (O_2694,N_29448,N_28995);
and UO_2695 (O_2695,N_29272,N_28897);
nor UO_2696 (O_2696,N_28819,N_29585);
xor UO_2697 (O_2697,N_29978,N_29438);
xnor UO_2698 (O_2698,N_29311,N_29075);
nor UO_2699 (O_2699,N_29409,N_29084);
nor UO_2700 (O_2700,N_29759,N_29214);
nand UO_2701 (O_2701,N_29586,N_29961);
xor UO_2702 (O_2702,N_29753,N_29995);
nor UO_2703 (O_2703,N_29194,N_29145);
xnor UO_2704 (O_2704,N_29645,N_29806);
nand UO_2705 (O_2705,N_29157,N_29509);
nand UO_2706 (O_2706,N_29221,N_28968);
nor UO_2707 (O_2707,N_29804,N_29474);
nor UO_2708 (O_2708,N_29501,N_29275);
nor UO_2709 (O_2709,N_28809,N_29286);
nor UO_2710 (O_2710,N_28945,N_28934);
nor UO_2711 (O_2711,N_28924,N_29008);
nand UO_2712 (O_2712,N_29624,N_28905);
nor UO_2713 (O_2713,N_29744,N_29743);
or UO_2714 (O_2714,N_29078,N_29794);
nand UO_2715 (O_2715,N_29234,N_28899);
or UO_2716 (O_2716,N_28895,N_29751);
nand UO_2717 (O_2717,N_29348,N_29501);
or UO_2718 (O_2718,N_29138,N_29744);
and UO_2719 (O_2719,N_28955,N_29760);
xnor UO_2720 (O_2720,N_29169,N_28888);
and UO_2721 (O_2721,N_29517,N_28805);
and UO_2722 (O_2722,N_29446,N_29451);
or UO_2723 (O_2723,N_29528,N_29877);
nand UO_2724 (O_2724,N_29562,N_29951);
nand UO_2725 (O_2725,N_28993,N_29566);
nand UO_2726 (O_2726,N_29494,N_28864);
nor UO_2727 (O_2727,N_29459,N_29645);
nor UO_2728 (O_2728,N_29579,N_29826);
nand UO_2729 (O_2729,N_29926,N_28909);
xnor UO_2730 (O_2730,N_29345,N_29782);
and UO_2731 (O_2731,N_29127,N_28909);
or UO_2732 (O_2732,N_28880,N_29750);
xnor UO_2733 (O_2733,N_29257,N_29431);
nand UO_2734 (O_2734,N_29882,N_29125);
nand UO_2735 (O_2735,N_28847,N_29681);
xor UO_2736 (O_2736,N_29241,N_29874);
nand UO_2737 (O_2737,N_29631,N_29654);
or UO_2738 (O_2738,N_29942,N_29251);
nand UO_2739 (O_2739,N_29086,N_29496);
nand UO_2740 (O_2740,N_29911,N_28860);
xnor UO_2741 (O_2741,N_28971,N_29981);
nand UO_2742 (O_2742,N_28922,N_29863);
nand UO_2743 (O_2743,N_28822,N_29606);
nor UO_2744 (O_2744,N_29176,N_28978);
or UO_2745 (O_2745,N_29375,N_29922);
and UO_2746 (O_2746,N_29970,N_29156);
nor UO_2747 (O_2747,N_29515,N_29283);
nand UO_2748 (O_2748,N_28878,N_29398);
or UO_2749 (O_2749,N_28837,N_29394);
nor UO_2750 (O_2750,N_29309,N_29661);
nor UO_2751 (O_2751,N_29419,N_29801);
nor UO_2752 (O_2752,N_29115,N_29982);
and UO_2753 (O_2753,N_29201,N_29723);
or UO_2754 (O_2754,N_29937,N_29194);
xnor UO_2755 (O_2755,N_29125,N_29242);
and UO_2756 (O_2756,N_29595,N_28842);
xor UO_2757 (O_2757,N_29009,N_28838);
or UO_2758 (O_2758,N_28966,N_29972);
nand UO_2759 (O_2759,N_29609,N_29848);
and UO_2760 (O_2760,N_29810,N_28869);
and UO_2761 (O_2761,N_29831,N_29101);
or UO_2762 (O_2762,N_29491,N_29612);
nor UO_2763 (O_2763,N_29920,N_29470);
or UO_2764 (O_2764,N_29657,N_29922);
nor UO_2765 (O_2765,N_29983,N_29239);
nor UO_2766 (O_2766,N_29075,N_29407);
and UO_2767 (O_2767,N_29566,N_29546);
xor UO_2768 (O_2768,N_29400,N_29556);
nor UO_2769 (O_2769,N_29413,N_29617);
nor UO_2770 (O_2770,N_29012,N_29627);
nor UO_2771 (O_2771,N_29121,N_29579);
nand UO_2772 (O_2772,N_29877,N_29787);
nor UO_2773 (O_2773,N_29148,N_29879);
xnor UO_2774 (O_2774,N_29851,N_29644);
and UO_2775 (O_2775,N_29112,N_29264);
or UO_2776 (O_2776,N_29141,N_28812);
and UO_2777 (O_2777,N_29872,N_29349);
nand UO_2778 (O_2778,N_29116,N_29483);
xnor UO_2779 (O_2779,N_29265,N_29481);
nor UO_2780 (O_2780,N_29816,N_29509);
and UO_2781 (O_2781,N_29602,N_29643);
nor UO_2782 (O_2782,N_29208,N_29967);
nor UO_2783 (O_2783,N_29775,N_29450);
nand UO_2784 (O_2784,N_28876,N_28801);
or UO_2785 (O_2785,N_29920,N_29240);
and UO_2786 (O_2786,N_29437,N_29249);
xor UO_2787 (O_2787,N_29966,N_29530);
xor UO_2788 (O_2788,N_29893,N_29317);
or UO_2789 (O_2789,N_29358,N_29738);
and UO_2790 (O_2790,N_29767,N_29594);
xnor UO_2791 (O_2791,N_29537,N_29495);
nor UO_2792 (O_2792,N_28864,N_29934);
or UO_2793 (O_2793,N_29955,N_29968);
nand UO_2794 (O_2794,N_29905,N_29494);
nand UO_2795 (O_2795,N_28944,N_29977);
xnor UO_2796 (O_2796,N_29311,N_29553);
and UO_2797 (O_2797,N_29086,N_29520);
xor UO_2798 (O_2798,N_29102,N_29818);
nand UO_2799 (O_2799,N_29669,N_29138);
or UO_2800 (O_2800,N_29483,N_29129);
xnor UO_2801 (O_2801,N_28825,N_29025);
nor UO_2802 (O_2802,N_29157,N_29715);
nor UO_2803 (O_2803,N_29741,N_29069);
nand UO_2804 (O_2804,N_29163,N_29338);
nand UO_2805 (O_2805,N_29555,N_29168);
and UO_2806 (O_2806,N_29927,N_29176);
nor UO_2807 (O_2807,N_28885,N_29258);
and UO_2808 (O_2808,N_29646,N_29751);
nor UO_2809 (O_2809,N_29497,N_29104);
nand UO_2810 (O_2810,N_29803,N_29451);
nand UO_2811 (O_2811,N_29635,N_29857);
or UO_2812 (O_2812,N_29575,N_28961);
nor UO_2813 (O_2813,N_29008,N_29001);
and UO_2814 (O_2814,N_29535,N_29039);
nand UO_2815 (O_2815,N_29001,N_29142);
or UO_2816 (O_2816,N_29147,N_28989);
and UO_2817 (O_2817,N_29741,N_29497);
or UO_2818 (O_2818,N_29018,N_29852);
nand UO_2819 (O_2819,N_29144,N_29244);
or UO_2820 (O_2820,N_29033,N_29376);
xnor UO_2821 (O_2821,N_29509,N_28936);
nand UO_2822 (O_2822,N_29901,N_29937);
nand UO_2823 (O_2823,N_29234,N_28883);
nand UO_2824 (O_2824,N_29942,N_28935);
or UO_2825 (O_2825,N_29269,N_29812);
xor UO_2826 (O_2826,N_28978,N_29778);
and UO_2827 (O_2827,N_29344,N_29480);
or UO_2828 (O_2828,N_29236,N_29059);
nand UO_2829 (O_2829,N_29890,N_28839);
or UO_2830 (O_2830,N_29320,N_29334);
xnor UO_2831 (O_2831,N_29480,N_29822);
nand UO_2832 (O_2832,N_29235,N_29381);
nand UO_2833 (O_2833,N_29475,N_29434);
nor UO_2834 (O_2834,N_29121,N_28865);
or UO_2835 (O_2835,N_29317,N_29244);
nand UO_2836 (O_2836,N_29962,N_29251);
and UO_2837 (O_2837,N_28906,N_29040);
xor UO_2838 (O_2838,N_29683,N_29054);
nand UO_2839 (O_2839,N_29271,N_29536);
and UO_2840 (O_2840,N_29078,N_28854);
nor UO_2841 (O_2841,N_29592,N_29611);
nor UO_2842 (O_2842,N_29902,N_29000);
nor UO_2843 (O_2843,N_29059,N_29293);
nand UO_2844 (O_2844,N_29369,N_29388);
xnor UO_2845 (O_2845,N_29273,N_29650);
or UO_2846 (O_2846,N_29378,N_29733);
xor UO_2847 (O_2847,N_29163,N_29023);
nand UO_2848 (O_2848,N_29806,N_29261);
nor UO_2849 (O_2849,N_29679,N_28829);
nor UO_2850 (O_2850,N_29395,N_29798);
and UO_2851 (O_2851,N_29611,N_29326);
nand UO_2852 (O_2852,N_29486,N_29325);
or UO_2853 (O_2853,N_29818,N_28967);
or UO_2854 (O_2854,N_29080,N_29033);
or UO_2855 (O_2855,N_29030,N_29441);
nor UO_2856 (O_2856,N_29813,N_29765);
or UO_2857 (O_2857,N_29059,N_29523);
or UO_2858 (O_2858,N_29700,N_29113);
and UO_2859 (O_2859,N_29708,N_29772);
or UO_2860 (O_2860,N_29944,N_29261);
xnor UO_2861 (O_2861,N_29089,N_29526);
and UO_2862 (O_2862,N_29202,N_29912);
or UO_2863 (O_2863,N_29286,N_29119);
nand UO_2864 (O_2864,N_29760,N_29115);
and UO_2865 (O_2865,N_29131,N_29569);
nand UO_2866 (O_2866,N_28876,N_28883);
nand UO_2867 (O_2867,N_29227,N_29659);
or UO_2868 (O_2868,N_29223,N_29272);
and UO_2869 (O_2869,N_29708,N_29743);
nand UO_2870 (O_2870,N_29454,N_29962);
nor UO_2871 (O_2871,N_29718,N_29372);
xnor UO_2872 (O_2872,N_28905,N_29224);
nand UO_2873 (O_2873,N_29740,N_29824);
xnor UO_2874 (O_2874,N_29393,N_28966);
xor UO_2875 (O_2875,N_28897,N_29735);
nor UO_2876 (O_2876,N_29474,N_29466);
or UO_2877 (O_2877,N_29797,N_29118);
xor UO_2878 (O_2878,N_29946,N_29463);
or UO_2879 (O_2879,N_28951,N_29535);
xnor UO_2880 (O_2880,N_29184,N_29563);
or UO_2881 (O_2881,N_29201,N_29395);
xnor UO_2882 (O_2882,N_28908,N_29353);
nand UO_2883 (O_2883,N_29636,N_28840);
or UO_2884 (O_2884,N_29788,N_29541);
nand UO_2885 (O_2885,N_29648,N_29113);
or UO_2886 (O_2886,N_29257,N_29172);
xor UO_2887 (O_2887,N_29669,N_29622);
and UO_2888 (O_2888,N_29113,N_29116);
xor UO_2889 (O_2889,N_29570,N_29322);
xor UO_2890 (O_2890,N_29467,N_29474);
and UO_2891 (O_2891,N_29703,N_28885);
nor UO_2892 (O_2892,N_28971,N_29700);
xor UO_2893 (O_2893,N_29616,N_29540);
xor UO_2894 (O_2894,N_29404,N_29347);
xnor UO_2895 (O_2895,N_29712,N_29977);
or UO_2896 (O_2896,N_29003,N_29520);
nand UO_2897 (O_2897,N_29880,N_28995);
nor UO_2898 (O_2898,N_29635,N_29203);
and UO_2899 (O_2899,N_29180,N_29841);
nand UO_2900 (O_2900,N_29163,N_29459);
xor UO_2901 (O_2901,N_29278,N_28854);
nand UO_2902 (O_2902,N_29981,N_29988);
or UO_2903 (O_2903,N_29524,N_29355);
nand UO_2904 (O_2904,N_29814,N_28902);
nand UO_2905 (O_2905,N_29059,N_29714);
and UO_2906 (O_2906,N_28804,N_29957);
nand UO_2907 (O_2907,N_29882,N_29625);
nand UO_2908 (O_2908,N_29587,N_29930);
or UO_2909 (O_2909,N_29587,N_29971);
or UO_2910 (O_2910,N_29593,N_29924);
nor UO_2911 (O_2911,N_29571,N_29461);
xor UO_2912 (O_2912,N_28809,N_29319);
nor UO_2913 (O_2913,N_28913,N_29441);
nor UO_2914 (O_2914,N_29495,N_29642);
or UO_2915 (O_2915,N_29692,N_29065);
or UO_2916 (O_2916,N_29423,N_29932);
nor UO_2917 (O_2917,N_28919,N_29365);
xor UO_2918 (O_2918,N_29155,N_29979);
nor UO_2919 (O_2919,N_28845,N_29090);
xor UO_2920 (O_2920,N_28870,N_29716);
nand UO_2921 (O_2921,N_29104,N_29890);
or UO_2922 (O_2922,N_29723,N_29465);
and UO_2923 (O_2923,N_29153,N_29567);
xnor UO_2924 (O_2924,N_29597,N_29938);
or UO_2925 (O_2925,N_29042,N_29280);
xor UO_2926 (O_2926,N_28860,N_29994);
nor UO_2927 (O_2927,N_29742,N_29792);
xor UO_2928 (O_2928,N_28964,N_29175);
or UO_2929 (O_2929,N_29575,N_28944);
nor UO_2930 (O_2930,N_28993,N_29868);
nor UO_2931 (O_2931,N_29539,N_29788);
xnor UO_2932 (O_2932,N_29987,N_29840);
nor UO_2933 (O_2933,N_28912,N_29052);
nand UO_2934 (O_2934,N_28991,N_29939);
nor UO_2935 (O_2935,N_29888,N_29177);
nand UO_2936 (O_2936,N_29779,N_29302);
and UO_2937 (O_2937,N_29527,N_29742);
xnor UO_2938 (O_2938,N_28978,N_29030);
nor UO_2939 (O_2939,N_29153,N_29444);
nand UO_2940 (O_2940,N_28999,N_29199);
or UO_2941 (O_2941,N_28888,N_29320);
nor UO_2942 (O_2942,N_29212,N_28857);
xor UO_2943 (O_2943,N_29750,N_29340);
xnor UO_2944 (O_2944,N_29326,N_29228);
or UO_2945 (O_2945,N_28814,N_29814);
and UO_2946 (O_2946,N_29076,N_29707);
nand UO_2947 (O_2947,N_29376,N_29831);
or UO_2948 (O_2948,N_28946,N_29636);
xnor UO_2949 (O_2949,N_29333,N_28983);
and UO_2950 (O_2950,N_29590,N_29567);
nand UO_2951 (O_2951,N_29463,N_29164);
nor UO_2952 (O_2952,N_29365,N_29732);
and UO_2953 (O_2953,N_29072,N_28966);
nor UO_2954 (O_2954,N_28838,N_29464);
and UO_2955 (O_2955,N_29299,N_29392);
or UO_2956 (O_2956,N_29366,N_29602);
and UO_2957 (O_2957,N_29109,N_29424);
nand UO_2958 (O_2958,N_29452,N_28810);
nand UO_2959 (O_2959,N_29251,N_29372);
xnor UO_2960 (O_2960,N_29114,N_29953);
and UO_2961 (O_2961,N_29940,N_29563);
and UO_2962 (O_2962,N_29653,N_29365);
and UO_2963 (O_2963,N_28959,N_29781);
nand UO_2964 (O_2964,N_29526,N_29350);
xnor UO_2965 (O_2965,N_29261,N_29216);
and UO_2966 (O_2966,N_29311,N_29624);
or UO_2967 (O_2967,N_29859,N_29190);
xor UO_2968 (O_2968,N_29489,N_29650);
nand UO_2969 (O_2969,N_29666,N_28819);
and UO_2970 (O_2970,N_29696,N_28818);
or UO_2971 (O_2971,N_29108,N_29978);
and UO_2972 (O_2972,N_29868,N_29533);
and UO_2973 (O_2973,N_29398,N_29270);
xor UO_2974 (O_2974,N_29918,N_28873);
nand UO_2975 (O_2975,N_29067,N_29645);
and UO_2976 (O_2976,N_29753,N_29650);
nand UO_2977 (O_2977,N_29635,N_28831);
and UO_2978 (O_2978,N_29877,N_29629);
nor UO_2979 (O_2979,N_28828,N_28964);
nor UO_2980 (O_2980,N_29983,N_29584);
nand UO_2981 (O_2981,N_29983,N_29950);
and UO_2982 (O_2982,N_29746,N_29586);
nand UO_2983 (O_2983,N_29890,N_29817);
nor UO_2984 (O_2984,N_29232,N_29599);
or UO_2985 (O_2985,N_28984,N_29970);
or UO_2986 (O_2986,N_28800,N_29075);
nand UO_2987 (O_2987,N_29992,N_28817);
nor UO_2988 (O_2988,N_29332,N_28858);
nor UO_2989 (O_2989,N_29075,N_29957);
and UO_2990 (O_2990,N_29216,N_29296);
and UO_2991 (O_2991,N_29684,N_29742);
or UO_2992 (O_2992,N_29957,N_29573);
nand UO_2993 (O_2993,N_29247,N_28968);
xor UO_2994 (O_2994,N_29058,N_29378);
and UO_2995 (O_2995,N_29756,N_28891);
nor UO_2996 (O_2996,N_29115,N_29230);
or UO_2997 (O_2997,N_29101,N_29365);
or UO_2998 (O_2998,N_29720,N_29591);
nand UO_2999 (O_2999,N_28952,N_29022);
nor UO_3000 (O_3000,N_29750,N_28881);
nor UO_3001 (O_3001,N_29257,N_29255);
nand UO_3002 (O_3002,N_29717,N_29968);
nor UO_3003 (O_3003,N_29106,N_29829);
and UO_3004 (O_3004,N_28803,N_29923);
or UO_3005 (O_3005,N_28937,N_29607);
xnor UO_3006 (O_3006,N_29059,N_29163);
nand UO_3007 (O_3007,N_29485,N_29473);
nor UO_3008 (O_3008,N_29164,N_29711);
xor UO_3009 (O_3009,N_29782,N_29423);
xor UO_3010 (O_3010,N_29608,N_29116);
nand UO_3011 (O_3011,N_29455,N_29588);
nor UO_3012 (O_3012,N_29803,N_29869);
xnor UO_3013 (O_3013,N_29418,N_29071);
nand UO_3014 (O_3014,N_29307,N_29134);
xor UO_3015 (O_3015,N_29606,N_28956);
nor UO_3016 (O_3016,N_29699,N_29225);
nor UO_3017 (O_3017,N_29439,N_29780);
or UO_3018 (O_3018,N_29543,N_29567);
nand UO_3019 (O_3019,N_29030,N_28822);
nor UO_3020 (O_3020,N_29917,N_29582);
nor UO_3021 (O_3021,N_29794,N_29448);
nand UO_3022 (O_3022,N_28871,N_28827);
nand UO_3023 (O_3023,N_29211,N_29220);
nor UO_3024 (O_3024,N_29517,N_28875);
or UO_3025 (O_3025,N_29667,N_29520);
nor UO_3026 (O_3026,N_29281,N_29634);
nand UO_3027 (O_3027,N_29899,N_29631);
nor UO_3028 (O_3028,N_29142,N_29534);
or UO_3029 (O_3029,N_29654,N_28890);
nor UO_3030 (O_3030,N_29059,N_28909);
or UO_3031 (O_3031,N_29458,N_29674);
nand UO_3032 (O_3032,N_29067,N_29203);
nor UO_3033 (O_3033,N_29184,N_29263);
or UO_3034 (O_3034,N_28893,N_29115);
and UO_3035 (O_3035,N_29518,N_29318);
nand UO_3036 (O_3036,N_29424,N_29379);
nor UO_3037 (O_3037,N_29768,N_29425);
xnor UO_3038 (O_3038,N_29905,N_29411);
and UO_3039 (O_3039,N_29112,N_29754);
nand UO_3040 (O_3040,N_29959,N_28993);
nand UO_3041 (O_3041,N_29633,N_29966);
or UO_3042 (O_3042,N_29932,N_29772);
xnor UO_3043 (O_3043,N_29834,N_29855);
xnor UO_3044 (O_3044,N_29565,N_29539);
or UO_3045 (O_3045,N_29421,N_29480);
nor UO_3046 (O_3046,N_29449,N_29135);
xor UO_3047 (O_3047,N_29368,N_28924);
nor UO_3048 (O_3048,N_28836,N_29442);
or UO_3049 (O_3049,N_29411,N_29501);
nand UO_3050 (O_3050,N_29422,N_29764);
and UO_3051 (O_3051,N_29562,N_28981);
xnor UO_3052 (O_3052,N_29850,N_29471);
nand UO_3053 (O_3053,N_29507,N_29256);
nor UO_3054 (O_3054,N_29210,N_29339);
xor UO_3055 (O_3055,N_29531,N_29164);
and UO_3056 (O_3056,N_29708,N_29530);
nand UO_3057 (O_3057,N_29697,N_29114);
and UO_3058 (O_3058,N_29538,N_28886);
nand UO_3059 (O_3059,N_28940,N_29206);
and UO_3060 (O_3060,N_29194,N_28928);
nand UO_3061 (O_3061,N_29342,N_29728);
and UO_3062 (O_3062,N_29535,N_29151);
or UO_3063 (O_3063,N_29497,N_28881);
or UO_3064 (O_3064,N_29316,N_29031);
or UO_3065 (O_3065,N_28986,N_29235);
xnor UO_3066 (O_3066,N_29341,N_29289);
nor UO_3067 (O_3067,N_29209,N_29247);
and UO_3068 (O_3068,N_29219,N_29882);
nor UO_3069 (O_3069,N_28958,N_29642);
nor UO_3070 (O_3070,N_29609,N_28999);
xor UO_3071 (O_3071,N_29401,N_29574);
or UO_3072 (O_3072,N_29867,N_29520);
xor UO_3073 (O_3073,N_28929,N_28810);
nor UO_3074 (O_3074,N_29591,N_29896);
and UO_3075 (O_3075,N_28924,N_29522);
nand UO_3076 (O_3076,N_29117,N_29856);
xor UO_3077 (O_3077,N_29902,N_29032);
nor UO_3078 (O_3078,N_29576,N_29568);
nor UO_3079 (O_3079,N_28831,N_29758);
xnor UO_3080 (O_3080,N_28829,N_29686);
and UO_3081 (O_3081,N_29357,N_29199);
and UO_3082 (O_3082,N_29781,N_28943);
xor UO_3083 (O_3083,N_29863,N_28852);
or UO_3084 (O_3084,N_29417,N_28824);
nand UO_3085 (O_3085,N_29025,N_29695);
or UO_3086 (O_3086,N_29489,N_29035);
and UO_3087 (O_3087,N_29542,N_29798);
or UO_3088 (O_3088,N_28804,N_29106);
xnor UO_3089 (O_3089,N_29052,N_29368);
nand UO_3090 (O_3090,N_28825,N_29601);
or UO_3091 (O_3091,N_29686,N_29871);
nor UO_3092 (O_3092,N_29079,N_29885);
and UO_3093 (O_3093,N_29048,N_29037);
xnor UO_3094 (O_3094,N_29736,N_29202);
nand UO_3095 (O_3095,N_29268,N_29486);
or UO_3096 (O_3096,N_28816,N_29682);
and UO_3097 (O_3097,N_29585,N_29629);
nor UO_3098 (O_3098,N_29949,N_29223);
xor UO_3099 (O_3099,N_29047,N_29124);
xor UO_3100 (O_3100,N_29298,N_29937);
nand UO_3101 (O_3101,N_29172,N_29900);
and UO_3102 (O_3102,N_28832,N_29569);
or UO_3103 (O_3103,N_29257,N_29992);
nand UO_3104 (O_3104,N_29346,N_29641);
nand UO_3105 (O_3105,N_29668,N_28858);
nand UO_3106 (O_3106,N_29989,N_29364);
and UO_3107 (O_3107,N_28970,N_29791);
nand UO_3108 (O_3108,N_29793,N_29469);
xor UO_3109 (O_3109,N_29399,N_29314);
nand UO_3110 (O_3110,N_29497,N_29864);
or UO_3111 (O_3111,N_29830,N_29381);
and UO_3112 (O_3112,N_29892,N_29530);
nor UO_3113 (O_3113,N_29213,N_29709);
nand UO_3114 (O_3114,N_29008,N_29977);
nor UO_3115 (O_3115,N_29450,N_29967);
and UO_3116 (O_3116,N_28993,N_28946);
or UO_3117 (O_3117,N_29071,N_29920);
and UO_3118 (O_3118,N_29708,N_29918);
or UO_3119 (O_3119,N_29203,N_29536);
and UO_3120 (O_3120,N_29794,N_29874);
nand UO_3121 (O_3121,N_29968,N_29259);
or UO_3122 (O_3122,N_29840,N_29792);
xor UO_3123 (O_3123,N_29292,N_29094);
xor UO_3124 (O_3124,N_29754,N_28977);
nor UO_3125 (O_3125,N_29331,N_29495);
or UO_3126 (O_3126,N_29712,N_29508);
and UO_3127 (O_3127,N_29411,N_29153);
or UO_3128 (O_3128,N_29445,N_29766);
nor UO_3129 (O_3129,N_29627,N_29751);
nor UO_3130 (O_3130,N_29932,N_29323);
or UO_3131 (O_3131,N_29613,N_29270);
xnor UO_3132 (O_3132,N_29928,N_29332);
or UO_3133 (O_3133,N_28838,N_29198);
or UO_3134 (O_3134,N_29393,N_29297);
and UO_3135 (O_3135,N_29974,N_29374);
nor UO_3136 (O_3136,N_29816,N_29529);
nand UO_3137 (O_3137,N_29929,N_29240);
xnor UO_3138 (O_3138,N_29975,N_29030);
or UO_3139 (O_3139,N_29062,N_29142);
nand UO_3140 (O_3140,N_28829,N_29017);
nor UO_3141 (O_3141,N_29634,N_29169);
or UO_3142 (O_3142,N_29625,N_29697);
or UO_3143 (O_3143,N_28948,N_28936);
nor UO_3144 (O_3144,N_29418,N_29320);
nor UO_3145 (O_3145,N_29229,N_29685);
and UO_3146 (O_3146,N_29611,N_29899);
nand UO_3147 (O_3147,N_29318,N_28831);
or UO_3148 (O_3148,N_29075,N_29673);
or UO_3149 (O_3149,N_29668,N_29822);
nor UO_3150 (O_3150,N_28816,N_28914);
and UO_3151 (O_3151,N_29626,N_29387);
and UO_3152 (O_3152,N_29219,N_29902);
or UO_3153 (O_3153,N_28806,N_29909);
nand UO_3154 (O_3154,N_28845,N_29837);
and UO_3155 (O_3155,N_29686,N_29517);
nand UO_3156 (O_3156,N_29819,N_28982);
nor UO_3157 (O_3157,N_29879,N_29715);
xor UO_3158 (O_3158,N_29242,N_29479);
and UO_3159 (O_3159,N_29249,N_29165);
and UO_3160 (O_3160,N_29913,N_29433);
nor UO_3161 (O_3161,N_29097,N_29579);
xor UO_3162 (O_3162,N_29726,N_28987);
nor UO_3163 (O_3163,N_29786,N_29854);
xor UO_3164 (O_3164,N_29506,N_29231);
or UO_3165 (O_3165,N_29683,N_29359);
xnor UO_3166 (O_3166,N_29868,N_29953);
or UO_3167 (O_3167,N_29066,N_29444);
nand UO_3168 (O_3168,N_29425,N_29928);
xnor UO_3169 (O_3169,N_29908,N_28843);
xnor UO_3170 (O_3170,N_28823,N_29217);
or UO_3171 (O_3171,N_29412,N_29112);
and UO_3172 (O_3172,N_29381,N_29294);
or UO_3173 (O_3173,N_29146,N_29153);
xnor UO_3174 (O_3174,N_29613,N_28950);
and UO_3175 (O_3175,N_28888,N_29927);
xnor UO_3176 (O_3176,N_28835,N_29671);
nand UO_3177 (O_3177,N_28846,N_29630);
nand UO_3178 (O_3178,N_29101,N_28837);
nand UO_3179 (O_3179,N_29737,N_29730);
nor UO_3180 (O_3180,N_29456,N_29895);
xnor UO_3181 (O_3181,N_29449,N_29255);
xnor UO_3182 (O_3182,N_29500,N_29867);
or UO_3183 (O_3183,N_29875,N_29703);
or UO_3184 (O_3184,N_29745,N_29351);
xor UO_3185 (O_3185,N_28917,N_28831);
xor UO_3186 (O_3186,N_28987,N_29428);
or UO_3187 (O_3187,N_29398,N_29992);
or UO_3188 (O_3188,N_29467,N_29437);
and UO_3189 (O_3189,N_29337,N_29093);
nor UO_3190 (O_3190,N_29056,N_29423);
xor UO_3191 (O_3191,N_29098,N_28928);
or UO_3192 (O_3192,N_29729,N_29960);
nor UO_3193 (O_3193,N_29040,N_29076);
nor UO_3194 (O_3194,N_29924,N_28840);
and UO_3195 (O_3195,N_29196,N_29855);
and UO_3196 (O_3196,N_29262,N_29070);
xor UO_3197 (O_3197,N_29590,N_28925);
xnor UO_3198 (O_3198,N_29597,N_29144);
or UO_3199 (O_3199,N_28854,N_29953);
or UO_3200 (O_3200,N_28879,N_29985);
nor UO_3201 (O_3201,N_29727,N_29060);
nand UO_3202 (O_3202,N_29895,N_29215);
and UO_3203 (O_3203,N_29829,N_29172);
and UO_3204 (O_3204,N_28876,N_29683);
xor UO_3205 (O_3205,N_29366,N_28804);
xnor UO_3206 (O_3206,N_29417,N_29766);
or UO_3207 (O_3207,N_29307,N_29486);
and UO_3208 (O_3208,N_29909,N_29714);
and UO_3209 (O_3209,N_28937,N_28844);
or UO_3210 (O_3210,N_29775,N_28941);
xor UO_3211 (O_3211,N_29358,N_29677);
nand UO_3212 (O_3212,N_29308,N_28863);
nor UO_3213 (O_3213,N_29380,N_29906);
nand UO_3214 (O_3214,N_29253,N_29212);
or UO_3215 (O_3215,N_28866,N_28815);
nand UO_3216 (O_3216,N_29807,N_29627);
or UO_3217 (O_3217,N_29737,N_29358);
nand UO_3218 (O_3218,N_29711,N_28847);
or UO_3219 (O_3219,N_29917,N_29941);
nor UO_3220 (O_3220,N_29591,N_29013);
or UO_3221 (O_3221,N_29104,N_29702);
and UO_3222 (O_3222,N_28813,N_29958);
nor UO_3223 (O_3223,N_29935,N_28927);
xor UO_3224 (O_3224,N_29535,N_29830);
or UO_3225 (O_3225,N_29989,N_29752);
xnor UO_3226 (O_3226,N_29697,N_29514);
nand UO_3227 (O_3227,N_29733,N_29580);
xnor UO_3228 (O_3228,N_29532,N_28955);
or UO_3229 (O_3229,N_29355,N_28980);
and UO_3230 (O_3230,N_29057,N_29076);
and UO_3231 (O_3231,N_29803,N_29455);
nor UO_3232 (O_3232,N_29113,N_29749);
and UO_3233 (O_3233,N_29655,N_29932);
and UO_3234 (O_3234,N_29831,N_29566);
nor UO_3235 (O_3235,N_29062,N_29933);
or UO_3236 (O_3236,N_29180,N_28862);
nor UO_3237 (O_3237,N_29358,N_29368);
xor UO_3238 (O_3238,N_29493,N_29415);
nor UO_3239 (O_3239,N_29258,N_29367);
and UO_3240 (O_3240,N_29010,N_29025);
xnor UO_3241 (O_3241,N_29746,N_29269);
nor UO_3242 (O_3242,N_29425,N_29756);
and UO_3243 (O_3243,N_29609,N_29853);
and UO_3244 (O_3244,N_29706,N_29754);
xor UO_3245 (O_3245,N_29844,N_28806);
xor UO_3246 (O_3246,N_28966,N_28911);
or UO_3247 (O_3247,N_29763,N_28868);
nor UO_3248 (O_3248,N_29698,N_29376);
and UO_3249 (O_3249,N_29322,N_29105);
xor UO_3250 (O_3250,N_29880,N_29741);
or UO_3251 (O_3251,N_29841,N_29160);
nand UO_3252 (O_3252,N_29671,N_29997);
nand UO_3253 (O_3253,N_28932,N_29650);
nor UO_3254 (O_3254,N_28886,N_29438);
nor UO_3255 (O_3255,N_28877,N_29216);
or UO_3256 (O_3256,N_29441,N_29577);
nor UO_3257 (O_3257,N_28846,N_29810);
and UO_3258 (O_3258,N_29258,N_29254);
and UO_3259 (O_3259,N_28829,N_29061);
nor UO_3260 (O_3260,N_29219,N_29710);
nor UO_3261 (O_3261,N_29322,N_28844);
and UO_3262 (O_3262,N_28974,N_29253);
nor UO_3263 (O_3263,N_28996,N_29018);
or UO_3264 (O_3264,N_28883,N_28839);
nand UO_3265 (O_3265,N_29552,N_29157);
xnor UO_3266 (O_3266,N_29219,N_29198);
nand UO_3267 (O_3267,N_28940,N_29074);
nand UO_3268 (O_3268,N_29495,N_28963);
nor UO_3269 (O_3269,N_29389,N_29648);
nor UO_3270 (O_3270,N_29441,N_29593);
xor UO_3271 (O_3271,N_29317,N_29840);
or UO_3272 (O_3272,N_29357,N_29715);
nand UO_3273 (O_3273,N_29854,N_29658);
xor UO_3274 (O_3274,N_29126,N_29128);
and UO_3275 (O_3275,N_28898,N_29727);
or UO_3276 (O_3276,N_29195,N_29325);
xor UO_3277 (O_3277,N_29833,N_29390);
and UO_3278 (O_3278,N_29236,N_29184);
xor UO_3279 (O_3279,N_29818,N_28915);
nand UO_3280 (O_3280,N_29703,N_29250);
xor UO_3281 (O_3281,N_29249,N_29883);
and UO_3282 (O_3282,N_28940,N_29023);
nor UO_3283 (O_3283,N_29065,N_29630);
or UO_3284 (O_3284,N_29263,N_29121);
xor UO_3285 (O_3285,N_29966,N_29889);
and UO_3286 (O_3286,N_29041,N_28879);
nand UO_3287 (O_3287,N_29031,N_29763);
nand UO_3288 (O_3288,N_29822,N_29497);
xor UO_3289 (O_3289,N_29686,N_28873);
xnor UO_3290 (O_3290,N_29703,N_29438);
xnor UO_3291 (O_3291,N_29735,N_29714);
nor UO_3292 (O_3292,N_29109,N_29056);
or UO_3293 (O_3293,N_29752,N_28951);
nor UO_3294 (O_3294,N_29102,N_29833);
or UO_3295 (O_3295,N_29719,N_29308);
xnor UO_3296 (O_3296,N_29449,N_29981);
xnor UO_3297 (O_3297,N_29636,N_29896);
xnor UO_3298 (O_3298,N_29186,N_29495);
or UO_3299 (O_3299,N_29784,N_29813);
xnor UO_3300 (O_3300,N_29706,N_29047);
xor UO_3301 (O_3301,N_29350,N_29036);
or UO_3302 (O_3302,N_29608,N_29378);
nor UO_3303 (O_3303,N_29510,N_29648);
and UO_3304 (O_3304,N_28823,N_29231);
or UO_3305 (O_3305,N_29849,N_29201);
and UO_3306 (O_3306,N_29473,N_29846);
nor UO_3307 (O_3307,N_29870,N_29791);
and UO_3308 (O_3308,N_29724,N_29207);
or UO_3309 (O_3309,N_29059,N_28908);
xnor UO_3310 (O_3310,N_29500,N_29606);
nor UO_3311 (O_3311,N_29627,N_29779);
nand UO_3312 (O_3312,N_28945,N_28881);
xor UO_3313 (O_3313,N_29004,N_28999);
nand UO_3314 (O_3314,N_29938,N_29470);
nor UO_3315 (O_3315,N_29182,N_29612);
or UO_3316 (O_3316,N_29526,N_28898);
and UO_3317 (O_3317,N_28876,N_28979);
and UO_3318 (O_3318,N_29637,N_28984);
nor UO_3319 (O_3319,N_29772,N_29805);
xor UO_3320 (O_3320,N_28967,N_29349);
xor UO_3321 (O_3321,N_29106,N_28995);
xnor UO_3322 (O_3322,N_29968,N_29678);
or UO_3323 (O_3323,N_28870,N_29148);
xor UO_3324 (O_3324,N_29861,N_29091);
nand UO_3325 (O_3325,N_29923,N_29234);
or UO_3326 (O_3326,N_29742,N_29194);
and UO_3327 (O_3327,N_29431,N_29059);
or UO_3328 (O_3328,N_29834,N_29007);
and UO_3329 (O_3329,N_29926,N_29136);
or UO_3330 (O_3330,N_29075,N_28822);
xnor UO_3331 (O_3331,N_28950,N_29660);
nand UO_3332 (O_3332,N_29689,N_29083);
or UO_3333 (O_3333,N_29984,N_29954);
xor UO_3334 (O_3334,N_28951,N_28827);
and UO_3335 (O_3335,N_28981,N_29166);
nor UO_3336 (O_3336,N_29028,N_29296);
xnor UO_3337 (O_3337,N_29145,N_29343);
or UO_3338 (O_3338,N_29028,N_29753);
xnor UO_3339 (O_3339,N_29566,N_28936);
and UO_3340 (O_3340,N_29436,N_29358);
or UO_3341 (O_3341,N_29670,N_29708);
nand UO_3342 (O_3342,N_29604,N_29556);
and UO_3343 (O_3343,N_29515,N_29974);
nand UO_3344 (O_3344,N_29069,N_29544);
or UO_3345 (O_3345,N_29397,N_29666);
and UO_3346 (O_3346,N_29450,N_29818);
or UO_3347 (O_3347,N_29387,N_29911);
xor UO_3348 (O_3348,N_29100,N_29572);
and UO_3349 (O_3349,N_28931,N_29860);
xor UO_3350 (O_3350,N_28881,N_29521);
and UO_3351 (O_3351,N_29949,N_29166);
xor UO_3352 (O_3352,N_29959,N_29338);
and UO_3353 (O_3353,N_29752,N_29300);
xor UO_3354 (O_3354,N_29187,N_28826);
nor UO_3355 (O_3355,N_28987,N_29939);
xnor UO_3356 (O_3356,N_29855,N_28878);
xnor UO_3357 (O_3357,N_29848,N_29418);
nand UO_3358 (O_3358,N_29526,N_29027);
or UO_3359 (O_3359,N_29823,N_29764);
nand UO_3360 (O_3360,N_29414,N_29784);
nand UO_3361 (O_3361,N_29829,N_28958);
nand UO_3362 (O_3362,N_29659,N_29080);
nand UO_3363 (O_3363,N_29019,N_29475);
or UO_3364 (O_3364,N_28986,N_29215);
nand UO_3365 (O_3365,N_29028,N_29655);
nor UO_3366 (O_3366,N_29361,N_29152);
or UO_3367 (O_3367,N_28974,N_29837);
nor UO_3368 (O_3368,N_28825,N_29343);
or UO_3369 (O_3369,N_29604,N_29683);
and UO_3370 (O_3370,N_29691,N_29289);
nand UO_3371 (O_3371,N_28936,N_29236);
nand UO_3372 (O_3372,N_29714,N_29658);
and UO_3373 (O_3373,N_28910,N_29007);
xor UO_3374 (O_3374,N_29666,N_28804);
xnor UO_3375 (O_3375,N_29471,N_29661);
or UO_3376 (O_3376,N_29432,N_29919);
nor UO_3377 (O_3377,N_29129,N_29585);
nor UO_3378 (O_3378,N_29701,N_29024);
nand UO_3379 (O_3379,N_28882,N_29476);
and UO_3380 (O_3380,N_29825,N_29660);
xor UO_3381 (O_3381,N_29885,N_29918);
and UO_3382 (O_3382,N_29478,N_29096);
nand UO_3383 (O_3383,N_29333,N_29277);
and UO_3384 (O_3384,N_29443,N_29812);
and UO_3385 (O_3385,N_29710,N_29527);
xor UO_3386 (O_3386,N_29998,N_29713);
nand UO_3387 (O_3387,N_29306,N_28995);
or UO_3388 (O_3388,N_29802,N_29813);
nor UO_3389 (O_3389,N_29405,N_29530);
or UO_3390 (O_3390,N_29694,N_29603);
and UO_3391 (O_3391,N_29648,N_29885);
xor UO_3392 (O_3392,N_28826,N_29009);
nand UO_3393 (O_3393,N_28994,N_28970);
xnor UO_3394 (O_3394,N_28840,N_29531);
and UO_3395 (O_3395,N_29347,N_29601);
xor UO_3396 (O_3396,N_29523,N_29986);
and UO_3397 (O_3397,N_29424,N_29296);
nand UO_3398 (O_3398,N_29102,N_29696);
nand UO_3399 (O_3399,N_29694,N_29126);
and UO_3400 (O_3400,N_28837,N_29180);
xor UO_3401 (O_3401,N_29153,N_28986);
and UO_3402 (O_3402,N_29405,N_29885);
and UO_3403 (O_3403,N_29202,N_29946);
and UO_3404 (O_3404,N_29057,N_28949);
and UO_3405 (O_3405,N_28983,N_28802);
xor UO_3406 (O_3406,N_29145,N_29544);
nor UO_3407 (O_3407,N_29793,N_29897);
nand UO_3408 (O_3408,N_29995,N_29994);
nor UO_3409 (O_3409,N_29372,N_29997);
and UO_3410 (O_3410,N_29577,N_29026);
xor UO_3411 (O_3411,N_29543,N_29945);
or UO_3412 (O_3412,N_28805,N_29005);
or UO_3413 (O_3413,N_28869,N_29318);
nor UO_3414 (O_3414,N_29885,N_29872);
and UO_3415 (O_3415,N_29061,N_29981);
nor UO_3416 (O_3416,N_29411,N_28930);
or UO_3417 (O_3417,N_29823,N_29176);
xor UO_3418 (O_3418,N_29396,N_29566);
and UO_3419 (O_3419,N_28931,N_29980);
xor UO_3420 (O_3420,N_28973,N_29817);
nor UO_3421 (O_3421,N_29367,N_29881);
nor UO_3422 (O_3422,N_29668,N_29055);
nand UO_3423 (O_3423,N_28976,N_29026);
or UO_3424 (O_3424,N_28990,N_29385);
nand UO_3425 (O_3425,N_29529,N_29940);
nor UO_3426 (O_3426,N_29570,N_29319);
nor UO_3427 (O_3427,N_29435,N_29313);
xnor UO_3428 (O_3428,N_28912,N_29876);
nor UO_3429 (O_3429,N_28882,N_28849);
and UO_3430 (O_3430,N_29714,N_29664);
nor UO_3431 (O_3431,N_29290,N_29321);
nand UO_3432 (O_3432,N_29920,N_28985);
nand UO_3433 (O_3433,N_29965,N_29644);
xnor UO_3434 (O_3434,N_29200,N_29801);
xnor UO_3435 (O_3435,N_29289,N_29454);
nand UO_3436 (O_3436,N_29761,N_29454);
xnor UO_3437 (O_3437,N_29762,N_29799);
nand UO_3438 (O_3438,N_29827,N_29237);
nand UO_3439 (O_3439,N_29172,N_29470);
or UO_3440 (O_3440,N_29007,N_29210);
or UO_3441 (O_3441,N_29993,N_29840);
and UO_3442 (O_3442,N_29938,N_29484);
nand UO_3443 (O_3443,N_28880,N_29664);
xor UO_3444 (O_3444,N_28810,N_29021);
nor UO_3445 (O_3445,N_29515,N_29291);
or UO_3446 (O_3446,N_28817,N_29677);
and UO_3447 (O_3447,N_29844,N_28893);
nor UO_3448 (O_3448,N_28890,N_29445);
and UO_3449 (O_3449,N_29268,N_29410);
and UO_3450 (O_3450,N_29035,N_29958);
and UO_3451 (O_3451,N_29753,N_29629);
and UO_3452 (O_3452,N_29526,N_29472);
nor UO_3453 (O_3453,N_29845,N_29686);
nor UO_3454 (O_3454,N_28923,N_29201);
or UO_3455 (O_3455,N_29014,N_28884);
and UO_3456 (O_3456,N_29624,N_29715);
xnor UO_3457 (O_3457,N_29470,N_29275);
nand UO_3458 (O_3458,N_29689,N_29407);
and UO_3459 (O_3459,N_29877,N_29918);
and UO_3460 (O_3460,N_29704,N_28977);
nand UO_3461 (O_3461,N_29222,N_29366);
and UO_3462 (O_3462,N_29702,N_29808);
and UO_3463 (O_3463,N_29194,N_29056);
nand UO_3464 (O_3464,N_29376,N_29628);
nor UO_3465 (O_3465,N_28901,N_29107);
nor UO_3466 (O_3466,N_28946,N_29675);
nand UO_3467 (O_3467,N_29883,N_28944);
nand UO_3468 (O_3468,N_29285,N_28865);
nor UO_3469 (O_3469,N_29449,N_29476);
and UO_3470 (O_3470,N_29575,N_29840);
or UO_3471 (O_3471,N_29692,N_29994);
nor UO_3472 (O_3472,N_29540,N_29079);
and UO_3473 (O_3473,N_28813,N_29278);
nand UO_3474 (O_3474,N_29787,N_28866);
nor UO_3475 (O_3475,N_29771,N_29169);
nor UO_3476 (O_3476,N_29340,N_29308);
xor UO_3477 (O_3477,N_29422,N_29660);
xnor UO_3478 (O_3478,N_28966,N_29340);
xnor UO_3479 (O_3479,N_29637,N_29963);
nand UO_3480 (O_3480,N_29928,N_29790);
xnor UO_3481 (O_3481,N_29938,N_29648);
xor UO_3482 (O_3482,N_29787,N_29688);
or UO_3483 (O_3483,N_29236,N_29218);
xor UO_3484 (O_3484,N_29882,N_28924);
or UO_3485 (O_3485,N_29389,N_29102);
nand UO_3486 (O_3486,N_29410,N_28955);
xor UO_3487 (O_3487,N_29292,N_29585);
or UO_3488 (O_3488,N_29584,N_29172);
and UO_3489 (O_3489,N_29218,N_29557);
xor UO_3490 (O_3490,N_29256,N_29598);
nor UO_3491 (O_3491,N_29403,N_28860);
nor UO_3492 (O_3492,N_29294,N_28943);
xnor UO_3493 (O_3493,N_29530,N_29200);
nand UO_3494 (O_3494,N_29373,N_29822);
xor UO_3495 (O_3495,N_28883,N_29401);
and UO_3496 (O_3496,N_28976,N_29358);
nand UO_3497 (O_3497,N_29190,N_29772);
nand UO_3498 (O_3498,N_29806,N_29614);
or UO_3499 (O_3499,N_29975,N_28907);
endmodule