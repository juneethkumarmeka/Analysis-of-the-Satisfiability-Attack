module basic_500_3000_500_60_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_468,In_47);
and U1 (N_1,In_308,In_173);
nor U2 (N_2,In_226,In_63);
or U3 (N_3,In_96,In_236);
nand U4 (N_4,In_478,In_156);
and U5 (N_5,In_209,In_348);
nand U6 (N_6,In_303,In_329);
or U7 (N_7,In_427,In_229);
or U8 (N_8,In_79,In_328);
nand U9 (N_9,In_385,In_284);
nand U10 (N_10,In_126,In_71);
nand U11 (N_11,In_208,In_278);
and U12 (N_12,In_492,In_86);
nand U13 (N_13,In_80,In_424);
and U14 (N_14,In_186,In_50);
or U15 (N_15,In_318,In_325);
or U16 (N_16,In_399,In_405);
or U17 (N_17,In_457,In_392);
and U18 (N_18,In_109,In_233);
and U19 (N_19,In_432,In_205);
and U20 (N_20,In_360,In_3);
and U21 (N_21,In_351,In_148);
nand U22 (N_22,In_43,In_41);
nor U23 (N_23,In_95,In_476);
nor U24 (N_24,In_197,In_112);
and U25 (N_25,In_474,In_172);
nand U26 (N_26,In_435,In_398);
or U27 (N_27,In_304,In_55);
or U28 (N_28,In_422,In_184);
and U29 (N_29,In_106,In_0);
nand U30 (N_30,In_370,In_389);
or U31 (N_31,In_105,In_78);
nor U32 (N_32,In_253,In_242);
nand U33 (N_33,In_54,In_271);
nand U34 (N_34,In_85,In_157);
nand U35 (N_35,In_280,In_339);
nand U36 (N_36,In_215,In_67);
nand U37 (N_37,In_116,In_252);
nor U38 (N_38,In_33,In_462);
nand U39 (N_39,In_181,In_285);
or U40 (N_40,In_98,In_188);
nand U41 (N_41,In_185,In_401);
or U42 (N_42,In_251,In_326);
or U43 (N_43,In_402,In_350);
and U44 (N_44,In_57,In_189);
nor U45 (N_45,In_246,In_368);
nor U46 (N_46,In_198,In_266);
nor U47 (N_47,In_296,In_4);
and U48 (N_48,In_30,In_65);
xnor U49 (N_49,In_400,In_119);
and U50 (N_50,In_60,In_499);
nor U51 (N_51,In_120,In_254);
nand U52 (N_52,N_25,In_301);
or U53 (N_53,In_124,N_38);
nand U54 (N_54,In_481,In_258);
nor U55 (N_55,In_343,In_23);
nand U56 (N_56,In_137,In_44);
nor U57 (N_57,In_480,In_443);
and U58 (N_58,In_445,In_341);
and U59 (N_59,In_321,In_323);
or U60 (N_60,In_130,In_361);
or U61 (N_61,In_456,In_428);
xor U62 (N_62,In_390,In_73);
or U63 (N_63,In_123,In_133);
nand U64 (N_64,In_267,In_93);
nand U65 (N_65,In_178,In_195);
nand U66 (N_66,In_35,In_74);
nand U67 (N_67,N_7,In_387);
or U68 (N_68,In_395,In_347);
nand U69 (N_69,In_300,In_430);
nor U70 (N_70,N_24,In_31);
or U71 (N_71,In_166,In_83);
xor U72 (N_72,In_175,In_324);
nand U73 (N_73,In_404,In_12);
nand U74 (N_74,In_384,In_230);
nand U75 (N_75,N_42,In_346);
or U76 (N_76,In_202,In_168);
nand U77 (N_77,In_210,In_442);
or U78 (N_78,In_411,In_451);
and U79 (N_79,In_255,In_39);
or U80 (N_80,In_18,In_279);
and U81 (N_81,In_491,In_261);
nand U82 (N_82,N_14,In_344);
or U83 (N_83,N_8,In_359);
and U84 (N_84,In_217,In_423);
and U85 (N_85,In_490,In_58);
nand U86 (N_86,In_433,In_221);
nand U87 (N_87,N_10,In_264);
and U88 (N_88,In_420,In_297);
and U89 (N_89,N_3,In_268);
or U90 (N_90,In_94,In_314);
and U91 (N_91,In_471,In_146);
and U92 (N_92,In_436,In_191);
nand U93 (N_93,In_394,In_291);
nand U94 (N_94,In_238,In_327);
and U95 (N_95,In_200,In_371);
or U96 (N_96,In_331,In_466);
nor U97 (N_97,N_37,N_6);
nand U98 (N_98,In_204,In_237);
nand U99 (N_99,In_357,In_257);
nor U100 (N_100,In_140,In_32);
xor U101 (N_101,In_447,In_338);
nor U102 (N_102,In_235,In_241);
nand U103 (N_103,In_378,In_482);
nor U104 (N_104,In_162,In_138);
and U105 (N_105,In_16,N_77);
or U106 (N_106,N_4,In_207);
and U107 (N_107,N_12,In_362);
nand U108 (N_108,N_41,In_169);
and U109 (N_109,In_170,In_380);
nor U110 (N_110,In_444,In_14);
or U111 (N_111,N_61,N_20);
and U112 (N_112,In_495,In_417);
nand U113 (N_113,In_472,In_459);
and U114 (N_114,N_70,In_29);
nor U115 (N_115,In_135,In_76);
nor U116 (N_116,In_440,In_25);
nor U117 (N_117,In_345,In_68);
nand U118 (N_118,N_83,In_115);
nor U119 (N_119,In_396,In_439);
nand U120 (N_120,In_11,In_22);
nand U121 (N_121,In_286,N_27);
nor U122 (N_122,In_243,In_46);
and U123 (N_123,In_372,In_488);
and U124 (N_124,In_358,In_88);
or U125 (N_125,N_29,In_302);
nand U126 (N_126,In_274,In_19);
nor U127 (N_127,N_72,N_18);
nand U128 (N_128,In_9,In_143);
nand U129 (N_129,In_1,N_21);
nand U130 (N_130,In_149,In_26);
nand U131 (N_131,N_11,N_19);
nor U132 (N_132,In_479,N_94);
and U133 (N_133,In_183,In_449);
xnor U134 (N_134,N_46,In_464);
nand U135 (N_135,N_45,In_410);
nor U136 (N_136,N_52,In_245);
nor U137 (N_137,In_218,N_75);
and U138 (N_138,In_320,In_309);
nor U139 (N_139,In_72,In_277);
or U140 (N_140,In_103,N_81);
or U141 (N_141,N_67,In_110);
or U142 (N_142,In_227,In_17);
or U143 (N_143,In_421,In_194);
nor U144 (N_144,In_64,In_414);
nor U145 (N_145,In_407,In_20);
or U146 (N_146,In_182,In_434);
nand U147 (N_147,In_250,In_377);
and U148 (N_148,In_335,In_216);
or U149 (N_149,In_275,N_48);
and U150 (N_150,N_98,N_130);
nand U151 (N_151,N_99,N_85);
nand U152 (N_152,N_114,In_81);
nand U153 (N_153,N_76,In_231);
nor U154 (N_154,N_31,N_0);
nand U155 (N_155,In_473,N_33);
nor U156 (N_156,N_131,In_317);
nor U157 (N_157,In_256,In_127);
and U158 (N_158,In_365,In_349);
nor U159 (N_159,In_452,In_403);
nand U160 (N_160,In_136,In_313);
nand U161 (N_161,In_262,N_26);
nand U162 (N_162,N_147,N_54);
or U163 (N_163,N_140,N_49);
and U164 (N_164,N_113,In_376);
and U165 (N_165,N_35,N_129);
nand U166 (N_166,N_55,N_63);
nor U167 (N_167,In_61,In_386);
or U168 (N_168,In_298,In_59);
nor U169 (N_169,N_136,In_219);
or U170 (N_170,In_355,In_408);
nor U171 (N_171,In_139,N_15);
nor U172 (N_172,In_107,In_49);
nor U173 (N_173,In_211,In_311);
nor U174 (N_174,In_333,In_485);
or U175 (N_175,In_458,N_137);
nand U176 (N_176,In_56,N_133);
or U177 (N_177,In_337,N_36);
or U178 (N_178,In_356,N_109);
nand U179 (N_179,In_496,In_330);
and U180 (N_180,In_379,In_282);
nand U181 (N_181,N_65,N_44);
nand U182 (N_182,N_106,In_315);
and U183 (N_183,In_159,In_214);
or U184 (N_184,In_228,In_51);
and U185 (N_185,In_90,In_369);
or U186 (N_186,In_155,N_139);
and U187 (N_187,In_415,In_269);
nand U188 (N_188,N_112,In_281);
and U189 (N_189,In_117,In_153);
nand U190 (N_190,N_105,In_463);
nand U191 (N_191,In_461,N_111);
nand U192 (N_192,In_310,In_36);
nand U193 (N_193,N_132,N_60);
nor U194 (N_194,N_102,N_56);
and U195 (N_195,In_299,In_265);
and U196 (N_196,In_486,In_89);
or U197 (N_197,In_190,In_244);
nor U198 (N_198,In_91,N_143);
nand U199 (N_199,In_145,In_332);
and U200 (N_200,N_2,N_53);
nand U201 (N_201,In_75,In_419);
nand U202 (N_202,In_273,N_164);
or U203 (N_203,N_116,In_69);
nor U204 (N_204,N_185,In_453);
and U205 (N_205,N_178,In_393);
nor U206 (N_206,In_259,N_127);
and U207 (N_207,In_460,In_37);
and U208 (N_208,In_307,N_160);
xor U209 (N_209,In_82,N_198);
nand U210 (N_210,In_224,In_382);
and U211 (N_211,In_114,In_164);
and U212 (N_212,N_23,In_494);
nor U213 (N_213,N_91,N_108);
nor U214 (N_214,In_352,N_122);
xor U215 (N_215,In_118,In_437);
and U216 (N_216,In_70,In_134);
nand U217 (N_217,N_159,N_190);
nand U218 (N_218,N_150,N_158);
or U219 (N_219,In_187,N_135);
nand U220 (N_220,In_441,In_288);
and U221 (N_221,N_180,N_152);
and U222 (N_222,N_172,In_426);
nand U223 (N_223,N_97,N_141);
or U224 (N_224,N_173,In_290);
and U225 (N_225,N_84,In_406);
nand U226 (N_226,N_16,N_22);
or U227 (N_227,N_151,In_469);
and U228 (N_228,N_119,N_169);
nand U229 (N_229,In_121,In_354);
and U230 (N_230,In_454,In_239);
and U231 (N_231,In_28,N_9);
nor U232 (N_232,N_191,In_38);
and U233 (N_233,N_28,N_149);
nor U234 (N_234,In_66,In_295);
nor U235 (N_235,In_87,In_381);
nor U236 (N_236,N_181,In_305);
nand U237 (N_237,In_223,In_467);
and U238 (N_238,In_289,In_8);
or U239 (N_239,N_118,In_319);
nor U240 (N_240,In_171,In_141);
and U241 (N_241,In_100,N_145);
nor U242 (N_242,In_113,N_68);
nor U243 (N_243,N_165,In_489);
or U244 (N_244,N_79,In_493);
and U245 (N_245,In_470,N_195);
nand U246 (N_246,In_48,N_40);
nor U247 (N_247,In_429,In_413);
nand U248 (N_248,In_498,N_155);
and U249 (N_249,In_5,N_101);
or U250 (N_250,N_66,In_455);
nor U251 (N_251,N_146,In_225);
and U252 (N_252,N_34,In_99);
nand U253 (N_253,In_151,In_128);
or U254 (N_254,N_232,In_40);
and U255 (N_255,N_194,N_214);
or U256 (N_256,N_204,In_363);
nand U257 (N_257,In_108,In_287);
or U258 (N_258,N_239,N_187);
and U259 (N_259,In_62,N_242);
nor U260 (N_260,In_249,In_283);
and U261 (N_261,In_111,In_477);
nand U262 (N_262,N_120,N_222);
and U263 (N_263,N_89,N_144);
nor U264 (N_264,N_215,In_383);
nand U265 (N_265,In_293,In_21);
or U266 (N_266,In_206,In_165);
and U267 (N_267,N_211,N_13);
nand U268 (N_268,N_229,N_64);
and U269 (N_269,N_92,In_342);
or U270 (N_270,N_138,N_103);
or U271 (N_271,In_316,In_222);
and U272 (N_272,In_92,In_42);
nand U273 (N_273,N_221,N_205);
nor U274 (N_274,In_270,In_483);
or U275 (N_275,In_122,In_27);
and U276 (N_276,In_179,In_147);
nor U277 (N_277,In_163,N_71);
and U278 (N_278,N_128,N_90);
nand U279 (N_279,N_58,N_104);
and U280 (N_280,N_184,N_197);
nor U281 (N_281,N_168,N_162);
nand U282 (N_282,In_177,N_47);
nor U283 (N_283,N_57,In_340);
nand U284 (N_284,In_240,N_154);
or U285 (N_285,N_212,In_272);
nand U286 (N_286,N_238,N_236);
and U287 (N_287,N_226,N_5);
xor U288 (N_288,N_225,In_465);
or U289 (N_289,In_129,N_176);
and U290 (N_290,N_100,N_174);
nand U291 (N_291,N_209,N_78);
or U292 (N_292,In_144,In_101);
nor U293 (N_293,In_260,N_74);
nand U294 (N_294,N_183,In_174);
nor U295 (N_295,N_244,In_132);
or U296 (N_296,N_30,In_276);
or U297 (N_297,In_425,N_123);
nor U298 (N_298,In_446,N_107);
nand U299 (N_299,In_97,In_52);
nor U300 (N_300,N_50,N_96);
or U301 (N_301,N_203,In_154);
or U302 (N_302,N_200,N_246);
nand U303 (N_303,N_110,N_234);
and U304 (N_304,N_230,In_34);
nor U305 (N_305,N_240,N_237);
xor U306 (N_306,N_170,N_249);
nand U307 (N_307,N_32,N_51);
and U308 (N_308,N_43,N_245);
and U309 (N_309,In_220,In_484);
xor U310 (N_310,N_235,In_53);
nor U311 (N_311,In_142,N_280);
nand U312 (N_312,N_295,N_296);
or U313 (N_313,In_448,In_336);
or U314 (N_314,N_219,N_257);
xor U315 (N_315,N_291,In_312);
xnor U316 (N_316,N_276,N_189);
and U317 (N_317,N_223,In_192);
and U318 (N_318,N_82,N_217);
or U319 (N_319,In_487,N_287);
and U320 (N_320,N_177,N_277);
nor U321 (N_321,N_278,N_115);
nand U322 (N_322,N_250,N_156);
xor U323 (N_323,N_252,N_88);
or U324 (N_324,N_282,In_150);
or U325 (N_325,N_175,In_366);
and U326 (N_326,N_210,In_374);
nand U327 (N_327,In_247,In_167);
or U328 (N_328,N_213,In_416);
nor U329 (N_329,In_388,N_17);
nor U330 (N_330,N_256,N_292);
and U331 (N_331,N_228,N_264);
nor U332 (N_332,N_216,In_306);
or U333 (N_333,In_292,N_1);
nand U334 (N_334,N_269,N_260);
nor U335 (N_335,N_124,N_186);
nand U336 (N_336,In_152,N_188);
or U337 (N_337,N_167,In_45);
and U338 (N_338,In_438,N_196);
and U339 (N_339,In_367,In_161);
nand U340 (N_340,In_409,N_293);
or U341 (N_341,N_95,In_176);
xor U342 (N_342,In_497,N_207);
or U343 (N_343,In_213,In_77);
nand U344 (N_344,N_59,In_334);
xor U345 (N_345,N_87,N_233);
and U346 (N_346,In_84,N_289);
nor U347 (N_347,In_263,N_288);
nor U348 (N_348,N_69,N_262);
nand U349 (N_349,In_102,N_62);
nand U350 (N_350,In_125,In_364);
nand U351 (N_351,In_375,N_319);
nor U352 (N_352,In_373,N_326);
nand U353 (N_353,In_450,N_182);
or U354 (N_354,N_323,N_307);
or U355 (N_355,N_259,N_268);
nor U356 (N_356,N_279,N_309);
nor U357 (N_357,N_261,In_397);
nor U358 (N_358,In_475,N_251);
and U359 (N_359,N_171,N_308);
or U360 (N_360,In_201,N_273);
and U361 (N_361,N_302,N_286);
nand U362 (N_362,N_339,In_104);
or U363 (N_363,N_39,In_212);
nand U364 (N_364,N_314,In_24);
or U365 (N_365,N_344,N_281);
and U366 (N_366,N_349,N_316);
or U367 (N_367,N_248,In_2);
and U368 (N_368,N_231,In_203);
nand U369 (N_369,N_255,N_337);
and U370 (N_370,N_247,N_335);
nand U371 (N_371,In_6,N_311);
nand U372 (N_372,N_299,In_7);
nand U373 (N_373,In_391,In_158);
nor U374 (N_374,N_317,N_313);
and U375 (N_375,N_341,N_199);
nand U376 (N_376,N_270,N_148);
and U377 (N_377,In_180,N_153);
nand U378 (N_378,N_285,N_193);
xor U379 (N_379,N_73,N_284);
nand U380 (N_380,In_196,N_202);
or U381 (N_381,N_330,N_327);
nor U382 (N_382,N_324,N_266);
and U383 (N_383,N_328,N_243);
nand U384 (N_384,In_131,N_346);
or U385 (N_385,N_320,N_322);
and U386 (N_386,N_241,N_321);
nor U387 (N_387,N_227,In_234);
or U388 (N_388,In_294,N_192);
or U389 (N_389,N_166,N_271);
nor U390 (N_390,In_193,N_294);
nand U391 (N_391,N_342,In_418);
and U392 (N_392,N_315,N_283);
nand U393 (N_393,N_121,N_300);
or U394 (N_394,N_297,In_412);
nor U395 (N_395,N_275,In_160);
nor U396 (N_396,N_258,N_345);
nor U397 (N_397,N_305,N_125);
or U398 (N_398,N_301,N_331);
or U399 (N_399,N_208,N_333);
and U400 (N_400,N_369,N_254);
xor U401 (N_401,N_338,N_303);
and U402 (N_402,N_376,In_322);
nand U403 (N_403,N_360,N_86);
nor U404 (N_404,N_389,N_380);
nand U405 (N_405,N_290,N_343);
or U406 (N_406,N_312,N_157);
or U407 (N_407,N_134,N_383);
nor U408 (N_408,N_355,N_126);
nor U409 (N_409,N_368,N_386);
nor U410 (N_410,N_201,N_272);
xnor U411 (N_411,N_347,N_265);
or U412 (N_412,N_224,N_359);
and U413 (N_413,N_253,N_267);
nor U414 (N_414,N_353,N_377);
nor U415 (N_415,N_348,N_340);
nor U416 (N_416,N_334,In_353);
nand U417 (N_417,N_336,N_354);
and U418 (N_418,N_163,N_395);
nand U419 (N_419,N_374,N_263);
nor U420 (N_420,N_364,N_385);
nand U421 (N_421,N_361,N_387);
nor U422 (N_422,N_373,N_206);
and U423 (N_423,N_142,N_332);
nand U424 (N_424,N_397,N_304);
nor U425 (N_425,In_431,In_13);
nand U426 (N_426,N_325,N_367);
nor U427 (N_427,N_366,N_384);
or U428 (N_428,N_370,N_357);
or U429 (N_429,N_356,N_310);
nand U430 (N_430,N_379,In_248);
nor U431 (N_431,N_93,N_392);
and U432 (N_432,N_274,N_329);
nand U433 (N_433,N_398,In_232);
or U434 (N_434,N_381,N_117);
or U435 (N_435,In_15,N_318);
nand U436 (N_436,N_351,N_220);
nand U437 (N_437,N_365,N_306);
nand U438 (N_438,N_80,N_371);
nand U439 (N_439,N_362,N_358);
and U440 (N_440,N_363,N_372);
and U441 (N_441,N_298,N_391);
and U442 (N_442,N_394,N_378);
nor U443 (N_443,In_199,N_350);
nor U444 (N_444,N_388,N_396);
or U445 (N_445,N_375,N_399);
nand U446 (N_446,N_161,In_10);
xnor U447 (N_447,N_218,N_179);
nand U448 (N_448,N_390,N_382);
or U449 (N_449,N_352,N_393);
and U450 (N_450,N_446,N_429);
and U451 (N_451,N_404,N_413);
and U452 (N_452,N_414,N_427);
or U453 (N_453,N_432,N_438);
nand U454 (N_454,N_422,N_442);
nand U455 (N_455,N_447,N_416);
nand U456 (N_456,N_408,N_435);
nor U457 (N_457,N_445,N_430);
and U458 (N_458,N_420,N_426);
or U459 (N_459,N_403,N_405);
nand U460 (N_460,N_440,N_407);
xnor U461 (N_461,N_433,N_406);
and U462 (N_462,N_425,N_409);
nor U463 (N_463,N_401,N_411);
nand U464 (N_464,N_423,N_428);
nand U465 (N_465,N_443,N_412);
nand U466 (N_466,N_421,N_434);
and U467 (N_467,N_448,N_400);
or U468 (N_468,N_410,N_439);
or U469 (N_469,N_415,N_444);
nor U470 (N_470,N_417,N_437);
nor U471 (N_471,N_441,N_419);
or U472 (N_472,N_418,N_449);
or U473 (N_473,N_431,N_424);
or U474 (N_474,N_402,N_436);
nor U475 (N_475,N_431,N_426);
or U476 (N_476,N_442,N_413);
and U477 (N_477,N_445,N_426);
xor U478 (N_478,N_442,N_434);
and U479 (N_479,N_439,N_423);
or U480 (N_480,N_439,N_443);
nor U481 (N_481,N_405,N_427);
and U482 (N_482,N_410,N_418);
nand U483 (N_483,N_420,N_409);
nand U484 (N_484,N_446,N_402);
and U485 (N_485,N_412,N_405);
xnor U486 (N_486,N_415,N_443);
and U487 (N_487,N_409,N_412);
nor U488 (N_488,N_425,N_416);
nor U489 (N_489,N_400,N_423);
nand U490 (N_490,N_444,N_412);
and U491 (N_491,N_411,N_447);
or U492 (N_492,N_437,N_416);
and U493 (N_493,N_425,N_417);
and U494 (N_494,N_401,N_419);
nor U495 (N_495,N_426,N_443);
xor U496 (N_496,N_405,N_436);
nand U497 (N_497,N_441,N_426);
or U498 (N_498,N_412,N_432);
nor U499 (N_499,N_408,N_440);
nor U500 (N_500,N_489,N_477);
and U501 (N_501,N_490,N_466);
nor U502 (N_502,N_491,N_474);
nor U503 (N_503,N_475,N_498);
or U504 (N_504,N_499,N_478);
or U505 (N_505,N_492,N_487);
nand U506 (N_506,N_485,N_450);
and U507 (N_507,N_476,N_462);
nand U508 (N_508,N_467,N_496);
nor U509 (N_509,N_483,N_497);
nand U510 (N_510,N_470,N_464);
and U511 (N_511,N_486,N_494);
or U512 (N_512,N_456,N_461);
nor U513 (N_513,N_482,N_452);
nand U514 (N_514,N_457,N_488);
and U515 (N_515,N_458,N_451);
nand U516 (N_516,N_493,N_481);
and U517 (N_517,N_465,N_453);
or U518 (N_518,N_471,N_459);
nand U519 (N_519,N_479,N_495);
and U520 (N_520,N_468,N_480);
or U521 (N_521,N_454,N_472);
nand U522 (N_522,N_469,N_484);
nand U523 (N_523,N_455,N_473);
nor U524 (N_524,N_463,N_460);
or U525 (N_525,N_457,N_452);
or U526 (N_526,N_477,N_479);
and U527 (N_527,N_486,N_496);
nand U528 (N_528,N_488,N_499);
nor U529 (N_529,N_461,N_455);
or U530 (N_530,N_486,N_452);
and U531 (N_531,N_479,N_468);
nor U532 (N_532,N_495,N_497);
and U533 (N_533,N_491,N_475);
nor U534 (N_534,N_484,N_476);
or U535 (N_535,N_469,N_489);
or U536 (N_536,N_491,N_485);
or U537 (N_537,N_461,N_491);
and U538 (N_538,N_485,N_474);
or U539 (N_539,N_473,N_478);
nor U540 (N_540,N_454,N_450);
or U541 (N_541,N_493,N_459);
nor U542 (N_542,N_470,N_495);
nand U543 (N_543,N_484,N_483);
nand U544 (N_544,N_472,N_459);
nand U545 (N_545,N_496,N_489);
nor U546 (N_546,N_472,N_486);
nor U547 (N_547,N_467,N_476);
nor U548 (N_548,N_490,N_463);
nor U549 (N_549,N_463,N_489);
nand U550 (N_550,N_507,N_509);
nand U551 (N_551,N_500,N_515);
nand U552 (N_552,N_529,N_541);
or U553 (N_553,N_519,N_524);
nor U554 (N_554,N_502,N_535);
or U555 (N_555,N_546,N_504);
and U556 (N_556,N_523,N_545);
and U557 (N_557,N_511,N_528);
nand U558 (N_558,N_506,N_527);
nand U559 (N_559,N_510,N_516);
nand U560 (N_560,N_548,N_531);
nand U561 (N_561,N_536,N_518);
or U562 (N_562,N_514,N_543);
nor U563 (N_563,N_540,N_533);
nand U564 (N_564,N_503,N_505);
or U565 (N_565,N_520,N_547);
nand U566 (N_566,N_513,N_522);
nor U567 (N_567,N_517,N_508);
or U568 (N_568,N_525,N_501);
nand U569 (N_569,N_544,N_542);
nor U570 (N_570,N_537,N_512);
nand U571 (N_571,N_538,N_521);
or U572 (N_572,N_539,N_534);
and U573 (N_573,N_530,N_526);
nor U574 (N_574,N_549,N_532);
nor U575 (N_575,N_533,N_513);
and U576 (N_576,N_541,N_518);
nand U577 (N_577,N_548,N_503);
xnor U578 (N_578,N_509,N_502);
nor U579 (N_579,N_508,N_539);
nand U580 (N_580,N_532,N_531);
nand U581 (N_581,N_504,N_549);
and U582 (N_582,N_536,N_532);
or U583 (N_583,N_502,N_543);
nand U584 (N_584,N_517,N_520);
nor U585 (N_585,N_534,N_530);
nand U586 (N_586,N_539,N_544);
and U587 (N_587,N_537,N_545);
nor U588 (N_588,N_526,N_520);
nand U589 (N_589,N_526,N_508);
nand U590 (N_590,N_530,N_505);
nand U591 (N_591,N_511,N_513);
and U592 (N_592,N_521,N_536);
or U593 (N_593,N_519,N_526);
and U594 (N_594,N_517,N_503);
nor U595 (N_595,N_536,N_514);
and U596 (N_596,N_518,N_512);
nand U597 (N_597,N_515,N_539);
or U598 (N_598,N_545,N_540);
and U599 (N_599,N_535,N_537);
or U600 (N_600,N_599,N_585);
and U601 (N_601,N_560,N_580);
and U602 (N_602,N_569,N_591);
and U603 (N_603,N_550,N_584);
and U604 (N_604,N_598,N_554);
nor U605 (N_605,N_581,N_568);
and U606 (N_606,N_565,N_553);
nand U607 (N_607,N_556,N_558);
and U608 (N_608,N_590,N_588);
nor U609 (N_609,N_597,N_595);
or U610 (N_610,N_579,N_557);
or U611 (N_611,N_582,N_594);
nor U612 (N_612,N_592,N_593);
nor U613 (N_613,N_596,N_576);
nand U614 (N_614,N_567,N_587);
nor U615 (N_615,N_570,N_552);
and U616 (N_616,N_559,N_573);
or U617 (N_617,N_571,N_586);
or U618 (N_618,N_555,N_561);
nor U619 (N_619,N_562,N_564);
nand U620 (N_620,N_551,N_583);
and U621 (N_621,N_574,N_589);
nor U622 (N_622,N_566,N_563);
and U623 (N_623,N_577,N_578);
or U624 (N_624,N_572,N_575);
and U625 (N_625,N_579,N_586);
nand U626 (N_626,N_585,N_561);
or U627 (N_627,N_593,N_554);
nor U628 (N_628,N_597,N_593);
or U629 (N_629,N_589,N_562);
nand U630 (N_630,N_586,N_578);
nor U631 (N_631,N_566,N_559);
nor U632 (N_632,N_585,N_581);
or U633 (N_633,N_576,N_552);
or U634 (N_634,N_588,N_589);
or U635 (N_635,N_592,N_597);
and U636 (N_636,N_568,N_594);
nor U637 (N_637,N_595,N_590);
nand U638 (N_638,N_595,N_573);
nor U639 (N_639,N_597,N_598);
nand U640 (N_640,N_581,N_567);
xnor U641 (N_641,N_582,N_586);
or U642 (N_642,N_594,N_556);
nand U643 (N_643,N_596,N_551);
or U644 (N_644,N_581,N_566);
and U645 (N_645,N_582,N_584);
nor U646 (N_646,N_574,N_588);
nand U647 (N_647,N_552,N_551);
nor U648 (N_648,N_585,N_588);
nor U649 (N_649,N_571,N_591);
or U650 (N_650,N_649,N_635);
nor U651 (N_651,N_636,N_623);
nor U652 (N_652,N_620,N_609);
and U653 (N_653,N_646,N_608);
nor U654 (N_654,N_625,N_644);
or U655 (N_655,N_622,N_614);
nand U656 (N_656,N_629,N_628);
or U657 (N_657,N_645,N_637);
nand U658 (N_658,N_616,N_648);
nor U659 (N_659,N_643,N_618);
or U660 (N_660,N_638,N_621);
and U661 (N_661,N_605,N_647);
or U662 (N_662,N_611,N_603);
nand U663 (N_663,N_601,N_633);
nand U664 (N_664,N_634,N_612);
and U665 (N_665,N_600,N_610);
and U666 (N_666,N_613,N_615);
nand U667 (N_667,N_617,N_631);
nand U668 (N_668,N_604,N_640);
xnor U669 (N_669,N_630,N_619);
and U670 (N_670,N_602,N_624);
nor U671 (N_671,N_607,N_627);
or U672 (N_672,N_606,N_626);
nor U673 (N_673,N_642,N_641);
nor U674 (N_674,N_632,N_639);
and U675 (N_675,N_617,N_611);
or U676 (N_676,N_630,N_640);
nand U677 (N_677,N_642,N_634);
nor U678 (N_678,N_628,N_633);
nand U679 (N_679,N_629,N_604);
or U680 (N_680,N_644,N_632);
or U681 (N_681,N_637,N_610);
or U682 (N_682,N_611,N_626);
nor U683 (N_683,N_638,N_631);
nand U684 (N_684,N_649,N_618);
or U685 (N_685,N_630,N_611);
nand U686 (N_686,N_626,N_609);
nor U687 (N_687,N_640,N_636);
nand U688 (N_688,N_639,N_605);
or U689 (N_689,N_623,N_640);
nor U690 (N_690,N_638,N_617);
nor U691 (N_691,N_625,N_619);
nand U692 (N_692,N_637,N_634);
nor U693 (N_693,N_603,N_639);
and U694 (N_694,N_649,N_603);
and U695 (N_695,N_636,N_607);
nor U696 (N_696,N_637,N_604);
and U697 (N_697,N_603,N_614);
and U698 (N_698,N_611,N_631);
and U699 (N_699,N_627,N_635);
and U700 (N_700,N_675,N_671);
nor U701 (N_701,N_667,N_660);
nor U702 (N_702,N_698,N_659);
nor U703 (N_703,N_669,N_690);
and U704 (N_704,N_681,N_665);
nand U705 (N_705,N_668,N_692);
and U706 (N_706,N_679,N_683);
nor U707 (N_707,N_689,N_658);
nor U708 (N_708,N_673,N_656);
nor U709 (N_709,N_677,N_680);
nand U710 (N_710,N_655,N_693);
xor U711 (N_711,N_687,N_670);
and U712 (N_712,N_653,N_685);
nand U713 (N_713,N_650,N_682);
and U714 (N_714,N_663,N_664);
nor U715 (N_715,N_686,N_661);
nand U716 (N_716,N_674,N_657);
nor U717 (N_717,N_651,N_696);
and U718 (N_718,N_678,N_684);
nand U719 (N_719,N_654,N_694);
or U720 (N_720,N_662,N_652);
and U721 (N_721,N_691,N_676);
or U722 (N_722,N_672,N_697);
or U723 (N_723,N_695,N_666);
xnor U724 (N_724,N_688,N_699);
nand U725 (N_725,N_650,N_671);
nor U726 (N_726,N_677,N_672);
nor U727 (N_727,N_672,N_684);
and U728 (N_728,N_689,N_681);
nand U729 (N_729,N_679,N_688);
nor U730 (N_730,N_678,N_659);
nand U731 (N_731,N_653,N_664);
and U732 (N_732,N_674,N_672);
nand U733 (N_733,N_689,N_673);
nand U734 (N_734,N_667,N_688);
or U735 (N_735,N_665,N_656);
xor U736 (N_736,N_691,N_697);
nand U737 (N_737,N_684,N_662);
nand U738 (N_738,N_668,N_675);
nor U739 (N_739,N_659,N_692);
nand U740 (N_740,N_670,N_680);
xor U741 (N_741,N_678,N_699);
nor U742 (N_742,N_684,N_661);
nor U743 (N_743,N_678,N_669);
and U744 (N_744,N_667,N_665);
or U745 (N_745,N_691,N_653);
xor U746 (N_746,N_689,N_686);
or U747 (N_747,N_691,N_693);
or U748 (N_748,N_681,N_691);
or U749 (N_749,N_697,N_670);
and U750 (N_750,N_749,N_704);
xor U751 (N_751,N_716,N_745);
nor U752 (N_752,N_705,N_723);
nor U753 (N_753,N_737,N_736);
nor U754 (N_754,N_739,N_708);
or U755 (N_755,N_714,N_710);
and U756 (N_756,N_724,N_709);
nor U757 (N_757,N_731,N_727);
nand U758 (N_758,N_746,N_747);
nand U759 (N_759,N_720,N_711);
nor U760 (N_760,N_701,N_721);
and U761 (N_761,N_725,N_734);
or U762 (N_762,N_740,N_728);
or U763 (N_763,N_712,N_738);
nor U764 (N_764,N_742,N_719);
and U765 (N_765,N_733,N_726);
nor U766 (N_766,N_741,N_707);
and U767 (N_767,N_744,N_706);
and U768 (N_768,N_718,N_730);
or U769 (N_769,N_722,N_732);
or U770 (N_770,N_729,N_713);
and U771 (N_771,N_715,N_703);
nand U772 (N_772,N_700,N_702);
and U773 (N_773,N_748,N_735);
nor U774 (N_774,N_717,N_743);
or U775 (N_775,N_706,N_739);
nor U776 (N_776,N_721,N_743);
nor U777 (N_777,N_732,N_733);
or U778 (N_778,N_711,N_738);
and U779 (N_779,N_744,N_749);
nor U780 (N_780,N_738,N_705);
or U781 (N_781,N_705,N_745);
nor U782 (N_782,N_731,N_716);
nor U783 (N_783,N_720,N_740);
nand U784 (N_784,N_727,N_701);
nand U785 (N_785,N_702,N_744);
nor U786 (N_786,N_700,N_743);
or U787 (N_787,N_722,N_707);
or U788 (N_788,N_717,N_710);
nor U789 (N_789,N_724,N_749);
nor U790 (N_790,N_707,N_731);
or U791 (N_791,N_704,N_722);
nor U792 (N_792,N_721,N_712);
nand U793 (N_793,N_724,N_742);
or U794 (N_794,N_725,N_744);
or U795 (N_795,N_703,N_705);
and U796 (N_796,N_704,N_700);
and U797 (N_797,N_725,N_746);
nor U798 (N_798,N_715,N_733);
or U799 (N_799,N_723,N_718);
nand U800 (N_800,N_776,N_791);
or U801 (N_801,N_790,N_797);
nor U802 (N_802,N_760,N_768);
xnor U803 (N_803,N_792,N_782);
or U804 (N_804,N_779,N_765);
nand U805 (N_805,N_795,N_784);
or U806 (N_806,N_781,N_750);
or U807 (N_807,N_794,N_761);
or U808 (N_808,N_786,N_766);
or U809 (N_809,N_775,N_751);
nand U810 (N_810,N_799,N_759);
nor U811 (N_811,N_769,N_772);
or U812 (N_812,N_764,N_787);
and U813 (N_813,N_762,N_758);
nand U814 (N_814,N_774,N_756);
nor U815 (N_815,N_789,N_777);
nand U816 (N_816,N_770,N_771);
xor U817 (N_817,N_773,N_755);
nor U818 (N_818,N_780,N_788);
nand U819 (N_819,N_752,N_754);
nor U820 (N_820,N_753,N_793);
or U821 (N_821,N_785,N_778);
nor U822 (N_822,N_798,N_783);
or U823 (N_823,N_796,N_767);
and U824 (N_824,N_757,N_763);
nand U825 (N_825,N_766,N_770);
or U826 (N_826,N_778,N_789);
and U827 (N_827,N_752,N_795);
xnor U828 (N_828,N_776,N_768);
or U829 (N_829,N_775,N_799);
and U830 (N_830,N_757,N_753);
or U831 (N_831,N_792,N_795);
or U832 (N_832,N_796,N_782);
and U833 (N_833,N_762,N_772);
and U834 (N_834,N_775,N_768);
nor U835 (N_835,N_787,N_750);
and U836 (N_836,N_768,N_789);
and U837 (N_837,N_796,N_784);
xor U838 (N_838,N_785,N_790);
nor U839 (N_839,N_767,N_764);
and U840 (N_840,N_788,N_751);
nor U841 (N_841,N_769,N_799);
or U842 (N_842,N_754,N_768);
or U843 (N_843,N_783,N_769);
or U844 (N_844,N_798,N_762);
nand U845 (N_845,N_795,N_765);
nand U846 (N_846,N_795,N_786);
and U847 (N_847,N_786,N_791);
nor U848 (N_848,N_750,N_792);
and U849 (N_849,N_789,N_783);
or U850 (N_850,N_821,N_814);
nor U851 (N_851,N_816,N_828);
or U852 (N_852,N_832,N_831);
nor U853 (N_853,N_805,N_807);
and U854 (N_854,N_836,N_819);
or U855 (N_855,N_843,N_849);
or U856 (N_856,N_837,N_842);
nor U857 (N_857,N_804,N_824);
nor U858 (N_858,N_839,N_801);
nor U859 (N_859,N_834,N_813);
nor U860 (N_860,N_833,N_827);
nand U861 (N_861,N_838,N_830);
nand U862 (N_862,N_815,N_817);
or U863 (N_863,N_847,N_820);
or U864 (N_864,N_818,N_823);
or U865 (N_865,N_825,N_803);
xnor U866 (N_866,N_800,N_810);
and U867 (N_867,N_806,N_829);
and U868 (N_868,N_848,N_808);
nor U869 (N_869,N_844,N_846);
or U870 (N_870,N_826,N_802);
and U871 (N_871,N_841,N_845);
xor U872 (N_872,N_811,N_840);
or U873 (N_873,N_822,N_835);
nand U874 (N_874,N_812,N_809);
nor U875 (N_875,N_832,N_823);
or U876 (N_876,N_820,N_812);
nand U877 (N_877,N_806,N_821);
nand U878 (N_878,N_806,N_800);
nor U879 (N_879,N_845,N_848);
or U880 (N_880,N_844,N_816);
or U881 (N_881,N_820,N_833);
or U882 (N_882,N_803,N_818);
or U883 (N_883,N_824,N_811);
nor U884 (N_884,N_823,N_842);
or U885 (N_885,N_805,N_847);
and U886 (N_886,N_800,N_808);
and U887 (N_887,N_840,N_835);
nor U888 (N_888,N_844,N_837);
nor U889 (N_889,N_817,N_840);
or U890 (N_890,N_849,N_846);
or U891 (N_891,N_825,N_821);
nor U892 (N_892,N_823,N_805);
or U893 (N_893,N_820,N_838);
and U894 (N_894,N_812,N_802);
and U895 (N_895,N_849,N_823);
and U896 (N_896,N_846,N_847);
nor U897 (N_897,N_822,N_815);
nand U898 (N_898,N_827,N_800);
or U899 (N_899,N_823,N_821);
nand U900 (N_900,N_864,N_870);
or U901 (N_901,N_899,N_882);
and U902 (N_902,N_898,N_893);
nand U903 (N_903,N_874,N_895);
xnor U904 (N_904,N_887,N_851);
nand U905 (N_905,N_894,N_873);
and U906 (N_906,N_868,N_862);
nand U907 (N_907,N_884,N_866);
nor U908 (N_908,N_890,N_863);
nand U909 (N_909,N_869,N_878);
nor U910 (N_910,N_856,N_897);
nand U911 (N_911,N_867,N_871);
nand U912 (N_912,N_880,N_859);
nor U913 (N_913,N_881,N_850);
nand U914 (N_914,N_891,N_854);
nor U915 (N_915,N_886,N_865);
or U916 (N_916,N_858,N_885);
nand U917 (N_917,N_876,N_883);
nor U918 (N_918,N_889,N_875);
nor U919 (N_919,N_860,N_853);
nand U920 (N_920,N_861,N_855);
xor U921 (N_921,N_872,N_879);
nand U922 (N_922,N_888,N_857);
nand U923 (N_923,N_896,N_877);
and U924 (N_924,N_852,N_892);
and U925 (N_925,N_897,N_881);
nand U926 (N_926,N_873,N_853);
xnor U927 (N_927,N_852,N_890);
nor U928 (N_928,N_883,N_878);
or U929 (N_929,N_875,N_888);
nor U930 (N_930,N_861,N_866);
nor U931 (N_931,N_888,N_861);
or U932 (N_932,N_861,N_897);
nor U933 (N_933,N_872,N_897);
nand U934 (N_934,N_896,N_886);
or U935 (N_935,N_860,N_865);
nand U936 (N_936,N_863,N_867);
and U937 (N_937,N_894,N_870);
nand U938 (N_938,N_854,N_890);
and U939 (N_939,N_889,N_899);
nor U940 (N_940,N_882,N_892);
nor U941 (N_941,N_860,N_893);
nor U942 (N_942,N_886,N_860);
nor U943 (N_943,N_877,N_867);
nor U944 (N_944,N_863,N_860);
and U945 (N_945,N_880,N_889);
nand U946 (N_946,N_868,N_864);
nand U947 (N_947,N_871,N_879);
or U948 (N_948,N_868,N_892);
nor U949 (N_949,N_879,N_883);
nand U950 (N_950,N_937,N_929);
xor U951 (N_951,N_903,N_941);
nand U952 (N_952,N_909,N_927);
or U953 (N_953,N_939,N_907);
and U954 (N_954,N_915,N_921);
nor U955 (N_955,N_906,N_926);
or U956 (N_956,N_935,N_946);
or U957 (N_957,N_914,N_912);
nor U958 (N_958,N_901,N_911);
xnor U959 (N_959,N_945,N_922);
nor U960 (N_960,N_923,N_934);
nand U961 (N_961,N_938,N_917);
or U962 (N_962,N_905,N_943);
or U963 (N_963,N_924,N_942);
or U964 (N_964,N_947,N_908);
nor U965 (N_965,N_913,N_933);
nor U966 (N_966,N_932,N_904);
nand U967 (N_967,N_920,N_940);
or U968 (N_968,N_931,N_944);
or U969 (N_969,N_928,N_902);
nor U970 (N_970,N_900,N_949);
nand U971 (N_971,N_948,N_919);
and U972 (N_972,N_918,N_936);
and U973 (N_973,N_910,N_916);
nor U974 (N_974,N_925,N_930);
and U975 (N_975,N_947,N_928);
nand U976 (N_976,N_941,N_901);
and U977 (N_977,N_944,N_909);
and U978 (N_978,N_936,N_901);
or U979 (N_979,N_946,N_931);
nand U980 (N_980,N_924,N_916);
nand U981 (N_981,N_942,N_905);
or U982 (N_982,N_924,N_918);
or U983 (N_983,N_907,N_922);
nand U984 (N_984,N_904,N_930);
nand U985 (N_985,N_939,N_948);
xor U986 (N_986,N_940,N_913);
or U987 (N_987,N_937,N_922);
or U988 (N_988,N_942,N_916);
xnor U989 (N_989,N_941,N_935);
nor U990 (N_990,N_936,N_907);
or U991 (N_991,N_936,N_906);
or U992 (N_992,N_912,N_904);
or U993 (N_993,N_908,N_912);
nand U994 (N_994,N_901,N_928);
nor U995 (N_995,N_908,N_931);
nor U996 (N_996,N_909,N_940);
or U997 (N_997,N_922,N_919);
nor U998 (N_998,N_938,N_918);
and U999 (N_999,N_941,N_912);
nand U1000 (N_1000,N_961,N_957);
xor U1001 (N_1001,N_994,N_950);
or U1002 (N_1002,N_956,N_993);
nor U1003 (N_1003,N_981,N_990);
or U1004 (N_1004,N_973,N_955);
nand U1005 (N_1005,N_975,N_966);
and U1006 (N_1006,N_951,N_996);
or U1007 (N_1007,N_971,N_987);
or U1008 (N_1008,N_984,N_967);
and U1009 (N_1009,N_976,N_962);
nand U1010 (N_1010,N_965,N_992);
or U1011 (N_1011,N_959,N_952);
nand U1012 (N_1012,N_997,N_977);
and U1013 (N_1013,N_974,N_983);
nand U1014 (N_1014,N_954,N_995);
or U1015 (N_1015,N_980,N_972);
nand U1016 (N_1016,N_991,N_989);
nand U1017 (N_1017,N_985,N_964);
or U1018 (N_1018,N_998,N_986);
or U1019 (N_1019,N_960,N_978);
nand U1020 (N_1020,N_953,N_982);
xor U1021 (N_1021,N_969,N_999);
and U1022 (N_1022,N_963,N_988);
nor U1023 (N_1023,N_958,N_970);
and U1024 (N_1024,N_968,N_979);
and U1025 (N_1025,N_976,N_983);
nor U1026 (N_1026,N_999,N_990);
nand U1027 (N_1027,N_977,N_990);
nor U1028 (N_1028,N_980,N_968);
nor U1029 (N_1029,N_965,N_975);
nor U1030 (N_1030,N_998,N_991);
nand U1031 (N_1031,N_978,N_966);
nand U1032 (N_1032,N_966,N_957);
nand U1033 (N_1033,N_981,N_984);
nor U1034 (N_1034,N_950,N_987);
nor U1035 (N_1035,N_956,N_994);
nor U1036 (N_1036,N_992,N_960);
nand U1037 (N_1037,N_970,N_992);
or U1038 (N_1038,N_952,N_985);
and U1039 (N_1039,N_978,N_994);
nor U1040 (N_1040,N_965,N_995);
or U1041 (N_1041,N_975,N_953);
nand U1042 (N_1042,N_951,N_973);
nand U1043 (N_1043,N_961,N_964);
nor U1044 (N_1044,N_975,N_963);
or U1045 (N_1045,N_995,N_989);
nand U1046 (N_1046,N_981,N_953);
and U1047 (N_1047,N_957,N_951);
nor U1048 (N_1048,N_991,N_961);
and U1049 (N_1049,N_951,N_972);
nand U1050 (N_1050,N_1038,N_1029);
and U1051 (N_1051,N_1031,N_1004);
xnor U1052 (N_1052,N_1009,N_1049);
nor U1053 (N_1053,N_1039,N_1028);
nand U1054 (N_1054,N_1002,N_1012);
or U1055 (N_1055,N_1006,N_1046);
or U1056 (N_1056,N_1035,N_1045);
or U1057 (N_1057,N_1020,N_1015);
or U1058 (N_1058,N_1013,N_1026);
nand U1059 (N_1059,N_1021,N_1043);
nand U1060 (N_1060,N_1023,N_1011);
and U1061 (N_1061,N_1018,N_1032);
or U1062 (N_1062,N_1007,N_1014);
nand U1063 (N_1063,N_1017,N_1033);
nand U1064 (N_1064,N_1003,N_1016);
nor U1065 (N_1065,N_1025,N_1001);
or U1066 (N_1066,N_1030,N_1044);
nand U1067 (N_1067,N_1042,N_1008);
and U1068 (N_1068,N_1024,N_1010);
nand U1069 (N_1069,N_1047,N_1022);
or U1070 (N_1070,N_1019,N_1041);
nand U1071 (N_1071,N_1036,N_1027);
or U1072 (N_1072,N_1040,N_1037);
nand U1073 (N_1073,N_1005,N_1048);
and U1074 (N_1074,N_1000,N_1034);
and U1075 (N_1075,N_1010,N_1013);
nand U1076 (N_1076,N_1038,N_1033);
nand U1077 (N_1077,N_1046,N_1030);
or U1078 (N_1078,N_1017,N_1043);
or U1079 (N_1079,N_1013,N_1011);
or U1080 (N_1080,N_1031,N_1021);
nand U1081 (N_1081,N_1003,N_1043);
nor U1082 (N_1082,N_1029,N_1034);
nand U1083 (N_1083,N_1015,N_1023);
or U1084 (N_1084,N_1031,N_1000);
nand U1085 (N_1085,N_1004,N_1019);
or U1086 (N_1086,N_1008,N_1049);
nor U1087 (N_1087,N_1035,N_1021);
nand U1088 (N_1088,N_1002,N_1023);
or U1089 (N_1089,N_1045,N_1028);
nor U1090 (N_1090,N_1013,N_1004);
or U1091 (N_1091,N_1046,N_1014);
or U1092 (N_1092,N_1003,N_1031);
and U1093 (N_1093,N_1030,N_1042);
nor U1094 (N_1094,N_1003,N_1034);
or U1095 (N_1095,N_1027,N_1035);
xor U1096 (N_1096,N_1019,N_1000);
nand U1097 (N_1097,N_1042,N_1047);
and U1098 (N_1098,N_1000,N_1015);
nand U1099 (N_1099,N_1037,N_1013);
and U1100 (N_1100,N_1088,N_1084);
nand U1101 (N_1101,N_1071,N_1051);
and U1102 (N_1102,N_1062,N_1092);
nand U1103 (N_1103,N_1067,N_1082);
nand U1104 (N_1104,N_1076,N_1056);
nand U1105 (N_1105,N_1065,N_1075);
nor U1106 (N_1106,N_1052,N_1090);
nand U1107 (N_1107,N_1083,N_1063);
nor U1108 (N_1108,N_1096,N_1070);
nand U1109 (N_1109,N_1064,N_1094);
nor U1110 (N_1110,N_1095,N_1059);
nand U1111 (N_1111,N_1089,N_1068);
nor U1112 (N_1112,N_1061,N_1085);
and U1113 (N_1113,N_1081,N_1097);
nand U1114 (N_1114,N_1054,N_1086);
nand U1115 (N_1115,N_1073,N_1069);
and U1116 (N_1116,N_1050,N_1066);
and U1117 (N_1117,N_1074,N_1080);
nand U1118 (N_1118,N_1099,N_1058);
or U1119 (N_1119,N_1091,N_1078);
nand U1120 (N_1120,N_1079,N_1053);
nor U1121 (N_1121,N_1055,N_1060);
or U1122 (N_1122,N_1077,N_1072);
or U1123 (N_1123,N_1087,N_1057);
nand U1124 (N_1124,N_1093,N_1098);
nor U1125 (N_1125,N_1052,N_1060);
or U1126 (N_1126,N_1077,N_1062);
or U1127 (N_1127,N_1057,N_1091);
or U1128 (N_1128,N_1051,N_1052);
nor U1129 (N_1129,N_1064,N_1086);
or U1130 (N_1130,N_1062,N_1091);
nand U1131 (N_1131,N_1091,N_1052);
nand U1132 (N_1132,N_1089,N_1081);
nor U1133 (N_1133,N_1065,N_1068);
nor U1134 (N_1134,N_1087,N_1091);
or U1135 (N_1135,N_1062,N_1074);
or U1136 (N_1136,N_1093,N_1064);
or U1137 (N_1137,N_1068,N_1095);
nor U1138 (N_1138,N_1097,N_1096);
and U1139 (N_1139,N_1097,N_1090);
and U1140 (N_1140,N_1061,N_1087);
and U1141 (N_1141,N_1097,N_1085);
nor U1142 (N_1142,N_1052,N_1067);
and U1143 (N_1143,N_1050,N_1074);
nor U1144 (N_1144,N_1072,N_1080);
nand U1145 (N_1145,N_1076,N_1071);
or U1146 (N_1146,N_1071,N_1081);
nor U1147 (N_1147,N_1090,N_1063);
and U1148 (N_1148,N_1073,N_1076);
nor U1149 (N_1149,N_1053,N_1097);
nor U1150 (N_1150,N_1128,N_1125);
and U1151 (N_1151,N_1126,N_1117);
or U1152 (N_1152,N_1104,N_1110);
nor U1153 (N_1153,N_1103,N_1138);
or U1154 (N_1154,N_1132,N_1129);
nor U1155 (N_1155,N_1136,N_1144);
and U1156 (N_1156,N_1147,N_1111);
nand U1157 (N_1157,N_1123,N_1127);
nor U1158 (N_1158,N_1120,N_1134);
nor U1159 (N_1159,N_1108,N_1143);
nor U1160 (N_1160,N_1140,N_1109);
nand U1161 (N_1161,N_1124,N_1114);
and U1162 (N_1162,N_1137,N_1118);
nand U1163 (N_1163,N_1133,N_1148);
and U1164 (N_1164,N_1121,N_1102);
nor U1165 (N_1165,N_1100,N_1115);
and U1166 (N_1166,N_1101,N_1141);
and U1167 (N_1167,N_1119,N_1145);
nor U1168 (N_1168,N_1139,N_1105);
and U1169 (N_1169,N_1107,N_1116);
nand U1170 (N_1170,N_1122,N_1135);
nor U1171 (N_1171,N_1113,N_1130);
or U1172 (N_1172,N_1146,N_1112);
or U1173 (N_1173,N_1106,N_1131);
and U1174 (N_1174,N_1142,N_1149);
and U1175 (N_1175,N_1113,N_1138);
nor U1176 (N_1176,N_1110,N_1140);
nand U1177 (N_1177,N_1107,N_1137);
and U1178 (N_1178,N_1113,N_1142);
and U1179 (N_1179,N_1108,N_1106);
nor U1180 (N_1180,N_1125,N_1134);
or U1181 (N_1181,N_1149,N_1134);
and U1182 (N_1182,N_1135,N_1101);
nand U1183 (N_1183,N_1138,N_1106);
and U1184 (N_1184,N_1116,N_1108);
and U1185 (N_1185,N_1131,N_1139);
nor U1186 (N_1186,N_1149,N_1105);
nand U1187 (N_1187,N_1114,N_1112);
and U1188 (N_1188,N_1108,N_1109);
xnor U1189 (N_1189,N_1104,N_1130);
nand U1190 (N_1190,N_1136,N_1126);
and U1191 (N_1191,N_1146,N_1147);
or U1192 (N_1192,N_1136,N_1142);
or U1193 (N_1193,N_1108,N_1146);
nor U1194 (N_1194,N_1103,N_1117);
nand U1195 (N_1195,N_1107,N_1136);
nand U1196 (N_1196,N_1125,N_1136);
nand U1197 (N_1197,N_1109,N_1127);
and U1198 (N_1198,N_1101,N_1129);
and U1199 (N_1199,N_1121,N_1109);
or U1200 (N_1200,N_1170,N_1157);
or U1201 (N_1201,N_1158,N_1194);
nand U1202 (N_1202,N_1187,N_1167);
nor U1203 (N_1203,N_1180,N_1179);
nand U1204 (N_1204,N_1192,N_1184);
nor U1205 (N_1205,N_1182,N_1155);
or U1206 (N_1206,N_1188,N_1195);
nor U1207 (N_1207,N_1154,N_1199);
nor U1208 (N_1208,N_1183,N_1172);
and U1209 (N_1209,N_1166,N_1159);
and U1210 (N_1210,N_1175,N_1164);
or U1211 (N_1211,N_1165,N_1153);
nand U1212 (N_1212,N_1191,N_1185);
or U1213 (N_1213,N_1150,N_1193);
and U1214 (N_1214,N_1196,N_1168);
and U1215 (N_1215,N_1177,N_1156);
and U1216 (N_1216,N_1169,N_1173);
and U1217 (N_1217,N_1198,N_1176);
nor U1218 (N_1218,N_1186,N_1174);
and U1219 (N_1219,N_1152,N_1189);
and U1220 (N_1220,N_1178,N_1161);
and U1221 (N_1221,N_1190,N_1151);
nand U1222 (N_1222,N_1171,N_1160);
nand U1223 (N_1223,N_1181,N_1162);
or U1224 (N_1224,N_1197,N_1163);
or U1225 (N_1225,N_1171,N_1158);
nor U1226 (N_1226,N_1169,N_1183);
nor U1227 (N_1227,N_1177,N_1180);
and U1228 (N_1228,N_1170,N_1181);
nand U1229 (N_1229,N_1155,N_1176);
or U1230 (N_1230,N_1163,N_1186);
nand U1231 (N_1231,N_1199,N_1194);
nor U1232 (N_1232,N_1178,N_1180);
and U1233 (N_1233,N_1160,N_1165);
nand U1234 (N_1234,N_1188,N_1164);
or U1235 (N_1235,N_1158,N_1155);
and U1236 (N_1236,N_1163,N_1179);
nand U1237 (N_1237,N_1179,N_1197);
or U1238 (N_1238,N_1173,N_1168);
or U1239 (N_1239,N_1166,N_1187);
or U1240 (N_1240,N_1189,N_1162);
and U1241 (N_1241,N_1187,N_1169);
and U1242 (N_1242,N_1170,N_1189);
and U1243 (N_1243,N_1165,N_1190);
or U1244 (N_1244,N_1160,N_1177);
or U1245 (N_1245,N_1188,N_1157);
nor U1246 (N_1246,N_1152,N_1194);
or U1247 (N_1247,N_1184,N_1166);
and U1248 (N_1248,N_1186,N_1169);
or U1249 (N_1249,N_1183,N_1165);
nor U1250 (N_1250,N_1222,N_1230);
or U1251 (N_1251,N_1236,N_1217);
nor U1252 (N_1252,N_1229,N_1232);
nand U1253 (N_1253,N_1228,N_1234);
and U1254 (N_1254,N_1247,N_1200);
xor U1255 (N_1255,N_1216,N_1227);
nor U1256 (N_1256,N_1209,N_1241);
nand U1257 (N_1257,N_1248,N_1203);
nand U1258 (N_1258,N_1243,N_1226);
nor U1259 (N_1259,N_1204,N_1244);
and U1260 (N_1260,N_1218,N_1235);
and U1261 (N_1261,N_1223,N_1212);
and U1262 (N_1262,N_1206,N_1207);
nor U1263 (N_1263,N_1239,N_1249);
nand U1264 (N_1264,N_1211,N_1221);
and U1265 (N_1265,N_1240,N_1219);
and U1266 (N_1266,N_1233,N_1242);
and U1267 (N_1267,N_1220,N_1201);
and U1268 (N_1268,N_1213,N_1210);
and U1269 (N_1269,N_1208,N_1224);
nand U1270 (N_1270,N_1205,N_1231);
nand U1271 (N_1271,N_1238,N_1245);
nand U1272 (N_1272,N_1202,N_1246);
or U1273 (N_1273,N_1237,N_1225);
nor U1274 (N_1274,N_1214,N_1215);
and U1275 (N_1275,N_1207,N_1245);
nand U1276 (N_1276,N_1228,N_1240);
or U1277 (N_1277,N_1221,N_1246);
nor U1278 (N_1278,N_1217,N_1203);
nand U1279 (N_1279,N_1213,N_1247);
or U1280 (N_1280,N_1210,N_1216);
nor U1281 (N_1281,N_1249,N_1208);
and U1282 (N_1282,N_1201,N_1239);
and U1283 (N_1283,N_1241,N_1227);
nand U1284 (N_1284,N_1237,N_1231);
xor U1285 (N_1285,N_1235,N_1212);
nand U1286 (N_1286,N_1225,N_1233);
nand U1287 (N_1287,N_1231,N_1223);
and U1288 (N_1288,N_1209,N_1206);
and U1289 (N_1289,N_1242,N_1231);
and U1290 (N_1290,N_1249,N_1241);
or U1291 (N_1291,N_1200,N_1226);
nand U1292 (N_1292,N_1235,N_1220);
and U1293 (N_1293,N_1211,N_1230);
or U1294 (N_1294,N_1231,N_1210);
or U1295 (N_1295,N_1201,N_1247);
and U1296 (N_1296,N_1222,N_1208);
nand U1297 (N_1297,N_1216,N_1201);
nor U1298 (N_1298,N_1246,N_1223);
nand U1299 (N_1299,N_1226,N_1225);
nand U1300 (N_1300,N_1279,N_1264);
nor U1301 (N_1301,N_1290,N_1295);
nor U1302 (N_1302,N_1291,N_1293);
xor U1303 (N_1303,N_1256,N_1271);
and U1304 (N_1304,N_1259,N_1278);
and U1305 (N_1305,N_1280,N_1285);
and U1306 (N_1306,N_1261,N_1266);
and U1307 (N_1307,N_1283,N_1253);
nand U1308 (N_1308,N_1287,N_1254);
and U1309 (N_1309,N_1276,N_1281);
nand U1310 (N_1310,N_1268,N_1251);
or U1311 (N_1311,N_1270,N_1255);
or U1312 (N_1312,N_1284,N_1252);
nand U1313 (N_1313,N_1298,N_1274);
or U1314 (N_1314,N_1297,N_1267);
or U1315 (N_1315,N_1260,N_1288);
or U1316 (N_1316,N_1258,N_1262);
nand U1317 (N_1317,N_1273,N_1282);
xor U1318 (N_1318,N_1286,N_1269);
nor U1319 (N_1319,N_1272,N_1289);
nand U1320 (N_1320,N_1299,N_1292);
nor U1321 (N_1321,N_1275,N_1296);
and U1322 (N_1322,N_1277,N_1257);
nor U1323 (N_1323,N_1265,N_1294);
nand U1324 (N_1324,N_1263,N_1250);
nor U1325 (N_1325,N_1279,N_1276);
nand U1326 (N_1326,N_1294,N_1297);
or U1327 (N_1327,N_1254,N_1251);
or U1328 (N_1328,N_1273,N_1274);
or U1329 (N_1329,N_1280,N_1297);
nor U1330 (N_1330,N_1271,N_1250);
nand U1331 (N_1331,N_1297,N_1291);
nand U1332 (N_1332,N_1295,N_1272);
nor U1333 (N_1333,N_1282,N_1260);
and U1334 (N_1334,N_1288,N_1285);
nand U1335 (N_1335,N_1258,N_1293);
xor U1336 (N_1336,N_1291,N_1276);
nor U1337 (N_1337,N_1257,N_1284);
nand U1338 (N_1338,N_1254,N_1282);
or U1339 (N_1339,N_1277,N_1254);
nor U1340 (N_1340,N_1273,N_1263);
or U1341 (N_1341,N_1279,N_1267);
nand U1342 (N_1342,N_1291,N_1277);
nand U1343 (N_1343,N_1291,N_1251);
nor U1344 (N_1344,N_1279,N_1258);
xor U1345 (N_1345,N_1287,N_1280);
nor U1346 (N_1346,N_1251,N_1252);
nor U1347 (N_1347,N_1252,N_1276);
nand U1348 (N_1348,N_1281,N_1280);
nand U1349 (N_1349,N_1287,N_1276);
or U1350 (N_1350,N_1312,N_1335);
nor U1351 (N_1351,N_1338,N_1347);
nor U1352 (N_1352,N_1330,N_1331);
nand U1353 (N_1353,N_1340,N_1346);
nor U1354 (N_1354,N_1305,N_1343);
and U1355 (N_1355,N_1314,N_1323);
nor U1356 (N_1356,N_1308,N_1348);
xor U1357 (N_1357,N_1344,N_1329);
and U1358 (N_1358,N_1345,N_1309);
and U1359 (N_1359,N_1306,N_1304);
and U1360 (N_1360,N_1313,N_1316);
nor U1361 (N_1361,N_1319,N_1303);
or U1362 (N_1362,N_1302,N_1349);
and U1363 (N_1363,N_1322,N_1333);
and U1364 (N_1364,N_1341,N_1337);
nor U1365 (N_1365,N_1324,N_1307);
xnor U1366 (N_1366,N_1327,N_1336);
nand U1367 (N_1367,N_1342,N_1328);
or U1368 (N_1368,N_1320,N_1310);
or U1369 (N_1369,N_1325,N_1326);
nor U1370 (N_1370,N_1321,N_1339);
and U1371 (N_1371,N_1315,N_1317);
nor U1372 (N_1372,N_1332,N_1311);
and U1373 (N_1373,N_1301,N_1300);
and U1374 (N_1374,N_1318,N_1334);
nor U1375 (N_1375,N_1346,N_1329);
and U1376 (N_1376,N_1329,N_1306);
nor U1377 (N_1377,N_1340,N_1309);
nand U1378 (N_1378,N_1327,N_1333);
xnor U1379 (N_1379,N_1338,N_1314);
nor U1380 (N_1380,N_1346,N_1315);
nor U1381 (N_1381,N_1326,N_1344);
nand U1382 (N_1382,N_1314,N_1306);
nor U1383 (N_1383,N_1311,N_1331);
nor U1384 (N_1384,N_1334,N_1336);
nor U1385 (N_1385,N_1314,N_1332);
and U1386 (N_1386,N_1345,N_1332);
nor U1387 (N_1387,N_1335,N_1323);
and U1388 (N_1388,N_1320,N_1330);
nor U1389 (N_1389,N_1300,N_1349);
nor U1390 (N_1390,N_1305,N_1334);
or U1391 (N_1391,N_1312,N_1344);
nand U1392 (N_1392,N_1305,N_1304);
nand U1393 (N_1393,N_1319,N_1344);
or U1394 (N_1394,N_1318,N_1315);
nand U1395 (N_1395,N_1327,N_1306);
nand U1396 (N_1396,N_1325,N_1322);
nand U1397 (N_1397,N_1323,N_1300);
nand U1398 (N_1398,N_1305,N_1326);
nand U1399 (N_1399,N_1324,N_1305);
nand U1400 (N_1400,N_1360,N_1393);
nand U1401 (N_1401,N_1374,N_1396);
nand U1402 (N_1402,N_1359,N_1395);
nand U1403 (N_1403,N_1363,N_1384);
nor U1404 (N_1404,N_1391,N_1368);
or U1405 (N_1405,N_1397,N_1386);
nand U1406 (N_1406,N_1380,N_1364);
and U1407 (N_1407,N_1375,N_1392);
or U1408 (N_1408,N_1352,N_1351);
and U1409 (N_1409,N_1354,N_1382);
or U1410 (N_1410,N_1353,N_1376);
and U1411 (N_1411,N_1350,N_1394);
nand U1412 (N_1412,N_1390,N_1362);
or U1413 (N_1413,N_1378,N_1366);
and U1414 (N_1414,N_1365,N_1399);
and U1415 (N_1415,N_1389,N_1398);
nor U1416 (N_1416,N_1377,N_1361);
nor U1417 (N_1417,N_1357,N_1383);
and U1418 (N_1418,N_1379,N_1367);
or U1419 (N_1419,N_1358,N_1381);
nor U1420 (N_1420,N_1388,N_1372);
and U1421 (N_1421,N_1373,N_1355);
nor U1422 (N_1422,N_1370,N_1385);
xor U1423 (N_1423,N_1371,N_1356);
nand U1424 (N_1424,N_1369,N_1387);
nor U1425 (N_1425,N_1365,N_1394);
nor U1426 (N_1426,N_1386,N_1382);
and U1427 (N_1427,N_1375,N_1385);
or U1428 (N_1428,N_1376,N_1374);
nor U1429 (N_1429,N_1369,N_1356);
or U1430 (N_1430,N_1365,N_1356);
nor U1431 (N_1431,N_1364,N_1355);
or U1432 (N_1432,N_1363,N_1397);
or U1433 (N_1433,N_1392,N_1397);
or U1434 (N_1434,N_1376,N_1399);
nor U1435 (N_1435,N_1391,N_1365);
nor U1436 (N_1436,N_1386,N_1351);
or U1437 (N_1437,N_1393,N_1383);
nand U1438 (N_1438,N_1367,N_1387);
nor U1439 (N_1439,N_1371,N_1379);
nand U1440 (N_1440,N_1380,N_1390);
nor U1441 (N_1441,N_1369,N_1371);
or U1442 (N_1442,N_1368,N_1352);
and U1443 (N_1443,N_1389,N_1382);
and U1444 (N_1444,N_1373,N_1376);
or U1445 (N_1445,N_1392,N_1388);
nand U1446 (N_1446,N_1397,N_1361);
nand U1447 (N_1447,N_1395,N_1376);
nor U1448 (N_1448,N_1380,N_1393);
xnor U1449 (N_1449,N_1355,N_1350);
or U1450 (N_1450,N_1412,N_1405);
and U1451 (N_1451,N_1448,N_1409);
or U1452 (N_1452,N_1411,N_1421);
nand U1453 (N_1453,N_1432,N_1424);
nand U1454 (N_1454,N_1431,N_1416);
nand U1455 (N_1455,N_1428,N_1437);
nor U1456 (N_1456,N_1445,N_1420);
nand U1457 (N_1457,N_1444,N_1447);
nand U1458 (N_1458,N_1400,N_1415);
and U1459 (N_1459,N_1413,N_1423);
nor U1460 (N_1460,N_1408,N_1449);
nand U1461 (N_1461,N_1414,N_1441);
nor U1462 (N_1462,N_1446,N_1443);
nor U1463 (N_1463,N_1422,N_1439);
or U1464 (N_1464,N_1417,N_1401);
nand U1465 (N_1465,N_1426,N_1404);
nor U1466 (N_1466,N_1429,N_1442);
nor U1467 (N_1467,N_1433,N_1438);
nor U1468 (N_1468,N_1410,N_1407);
nand U1469 (N_1469,N_1419,N_1418);
nand U1470 (N_1470,N_1425,N_1435);
nand U1471 (N_1471,N_1436,N_1403);
or U1472 (N_1472,N_1406,N_1427);
or U1473 (N_1473,N_1440,N_1430);
and U1474 (N_1474,N_1434,N_1402);
nand U1475 (N_1475,N_1402,N_1420);
or U1476 (N_1476,N_1409,N_1405);
nor U1477 (N_1477,N_1424,N_1408);
or U1478 (N_1478,N_1423,N_1421);
or U1479 (N_1479,N_1441,N_1402);
nor U1480 (N_1480,N_1400,N_1405);
or U1481 (N_1481,N_1420,N_1432);
nand U1482 (N_1482,N_1419,N_1441);
nand U1483 (N_1483,N_1415,N_1402);
nor U1484 (N_1484,N_1404,N_1430);
nand U1485 (N_1485,N_1449,N_1414);
or U1486 (N_1486,N_1434,N_1404);
or U1487 (N_1487,N_1432,N_1448);
or U1488 (N_1488,N_1408,N_1407);
or U1489 (N_1489,N_1432,N_1401);
nor U1490 (N_1490,N_1410,N_1425);
and U1491 (N_1491,N_1449,N_1442);
and U1492 (N_1492,N_1428,N_1434);
and U1493 (N_1493,N_1425,N_1445);
nor U1494 (N_1494,N_1427,N_1430);
and U1495 (N_1495,N_1429,N_1418);
nand U1496 (N_1496,N_1410,N_1421);
or U1497 (N_1497,N_1417,N_1449);
nand U1498 (N_1498,N_1431,N_1427);
or U1499 (N_1499,N_1423,N_1408);
or U1500 (N_1500,N_1474,N_1491);
nor U1501 (N_1501,N_1493,N_1453);
nand U1502 (N_1502,N_1488,N_1490);
and U1503 (N_1503,N_1480,N_1459);
nor U1504 (N_1504,N_1454,N_1476);
xnor U1505 (N_1505,N_1466,N_1468);
and U1506 (N_1506,N_1497,N_1487);
nor U1507 (N_1507,N_1495,N_1475);
nor U1508 (N_1508,N_1467,N_1483);
and U1509 (N_1509,N_1471,N_1499);
or U1510 (N_1510,N_1482,N_1481);
or U1511 (N_1511,N_1472,N_1492);
and U1512 (N_1512,N_1479,N_1460);
nand U1513 (N_1513,N_1478,N_1498);
and U1514 (N_1514,N_1451,N_1469);
nor U1515 (N_1515,N_1484,N_1465);
or U1516 (N_1516,N_1489,N_1464);
or U1517 (N_1517,N_1462,N_1485);
nor U1518 (N_1518,N_1461,N_1486);
and U1519 (N_1519,N_1450,N_1458);
nand U1520 (N_1520,N_1455,N_1457);
nand U1521 (N_1521,N_1496,N_1470);
nor U1522 (N_1522,N_1473,N_1456);
or U1523 (N_1523,N_1463,N_1477);
and U1524 (N_1524,N_1494,N_1452);
nor U1525 (N_1525,N_1461,N_1466);
nand U1526 (N_1526,N_1483,N_1471);
or U1527 (N_1527,N_1495,N_1496);
nor U1528 (N_1528,N_1471,N_1480);
and U1529 (N_1529,N_1459,N_1478);
nand U1530 (N_1530,N_1476,N_1480);
nand U1531 (N_1531,N_1471,N_1472);
or U1532 (N_1532,N_1462,N_1484);
nor U1533 (N_1533,N_1471,N_1492);
xor U1534 (N_1534,N_1460,N_1466);
nor U1535 (N_1535,N_1478,N_1467);
xor U1536 (N_1536,N_1496,N_1453);
and U1537 (N_1537,N_1461,N_1455);
or U1538 (N_1538,N_1477,N_1483);
and U1539 (N_1539,N_1498,N_1482);
nand U1540 (N_1540,N_1461,N_1464);
or U1541 (N_1541,N_1452,N_1482);
nand U1542 (N_1542,N_1467,N_1487);
nand U1543 (N_1543,N_1463,N_1483);
xor U1544 (N_1544,N_1484,N_1461);
nor U1545 (N_1545,N_1485,N_1499);
and U1546 (N_1546,N_1457,N_1482);
xnor U1547 (N_1547,N_1468,N_1490);
or U1548 (N_1548,N_1450,N_1497);
nor U1549 (N_1549,N_1470,N_1455);
nand U1550 (N_1550,N_1547,N_1513);
or U1551 (N_1551,N_1532,N_1536);
nor U1552 (N_1552,N_1533,N_1541);
and U1553 (N_1553,N_1539,N_1538);
or U1554 (N_1554,N_1520,N_1527);
nand U1555 (N_1555,N_1521,N_1535);
or U1556 (N_1556,N_1503,N_1504);
nand U1557 (N_1557,N_1508,N_1500);
or U1558 (N_1558,N_1502,N_1540);
or U1559 (N_1559,N_1542,N_1522);
nand U1560 (N_1560,N_1510,N_1548);
nor U1561 (N_1561,N_1516,N_1501);
or U1562 (N_1562,N_1506,N_1515);
nor U1563 (N_1563,N_1525,N_1518);
and U1564 (N_1564,N_1543,N_1537);
nand U1565 (N_1565,N_1546,N_1524);
or U1566 (N_1566,N_1511,N_1545);
nor U1567 (N_1567,N_1534,N_1530);
and U1568 (N_1568,N_1526,N_1519);
or U1569 (N_1569,N_1514,N_1523);
nor U1570 (N_1570,N_1544,N_1528);
nor U1571 (N_1571,N_1529,N_1549);
and U1572 (N_1572,N_1517,N_1509);
or U1573 (N_1573,N_1505,N_1531);
or U1574 (N_1574,N_1512,N_1507);
nor U1575 (N_1575,N_1501,N_1511);
or U1576 (N_1576,N_1540,N_1505);
nor U1577 (N_1577,N_1514,N_1535);
nor U1578 (N_1578,N_1545,N_1508);
or U1579 (N_1579,N_1507,N_1519);
nor U1580 (N_1580,N_1518,N_1545);
nand U1581 (N_1581,N_1502,N_1509);
or U1582 (N_1582,N_1501,N_1547);
nand U1583 (N_1583,N_1545,N_1519);
and U1584 (N_1584,N_1508,N_1512);
nor U1585 (N_1585,N_1524,N_1545);
and U1586 (N_1586,N_1536,N_1507);
nor U1587 (N_1587,N_1537,N_1522);
or U1588 (N_1588,N_1507,N_1537);
nand U1589 (N_1589,N_1542,N_1535);
or U1590 (N_1590,N_1546,N_1512);
nor U1591 (N_1591,N_1542,N_1549);
and U1592 (N_1592,N_1521,N_1542);
or U1593 (N_1593,N_1540,N_1528);
or U1594 (N_1594,N_1542,N_1548);
and U1595 (N_1595,N_1500,N_1529);
nand U1596 (N_1596,N_1534,N_1539);
xor U1597 (N_1597,N_1527,N_1523);
and U1598 (N_1598,N_1541,N_1531);
and U1599 (N_1599,N_1513,N_1546);
nor U1600 (N_1600,N_1550,N_1558);
or U1601 (N_1601,N_1572,N_1586);
nand U1602 (N_1602,N_1599,N_1588);
or U1603 (N_1603,N_1570,N_1577);
nand U1604 (N_1604,N_1573,N_1571);
and U1605 (N_1605,N_1567,N_1595);
and U1606 (N_1606,N_1576,N_1593);
and U1607 (N_1607,N_1590,N_1553);
nor U1608 (N_1608,N_1597,N_1575);
nand U1609 (N_1609,N_1579,N_1580);
nand U1610 (N_1610,N_1578,N_1566);
nor U1611 (N_1611,N_1592,N_1555);
nand U1612 (N_1612,N_1581,N_1563);
nand U1613 (N_1613,N_1585,N_1564);
or U1614 (N_1614,N_1591,N_1557);
and U1615 (N_1615,N_1589,N_1587);
nor U1616 (N_1616,N_1556,N_1552);
nand U1617 (N_1617,N_1551,N_1560);
nor U1618 (N_1618,N_1594,N_1574);
nand U1619 (N_1619,N_1568,N_1565);
nor U1620 (N_1620,N_1559,N_1596);
nand U1621 (N_1621,N_1562,N_1582);
nand U1622 (N_1622,N_1584,N_1569);
nor U1623 (N_1623,N_1598,N_1561);
or U1624 (N_1624,N_1554,N_1583);
or U1625 (N_1625,N_1555,N_1566);
nor U1626 (N_1626,N_1558,N_1562);
nand U1627 (N_1627,N_1550,N_1572);
xnor U1628 (N_1628,N_1596,N_1566);
or U1629 (N_1629,N_1580,N_1574);
nor U1630 (N_1630,N_1586,N_1597);
nor U1631 (N_1631,N_1553,N_1582);
or U1632 (N_1632,N_1562,N_1556);
nand U1633 (N_1633,N_1567,N_1598);
or U1634 (N_1634,N_1573,N_1580);
nor U1635 (N_1635,N_1572,N_1580);
nand U1636 (N_1636,N_1555,N_1599);
nand U1637 (N_1637,N_1592,N_1574);
and U1638 (N_1638,N_1565,N_1584);
xor U1639 (N_1639,N_1592,N_1561);
and U1640 (N_1640,N_1593,N_1564);
and U1641 (N_1641,N_1564,N_1561);
and U1642 (N_1642,N_1580,N_1585);
nand U1643 (N_1643,N_1559,N_1586);
nor U1644 (N_1644,N_1564,N_1598);
nor U1645 (N_1645,N_1581,N_1551);
or U1646 (N_1646,N_1594,N_1584);
and U1647 (N_1647,N_1589,N_1578);
or U1648 (N_1648,N_1563,N_1561);
or U1649 (N_1649,N_1561,N_1550);
nand U1650 (N_1650,N_1638,N_1632);
and U1651 (N_1651,N_1601,N_1614);
nand U1652 (N_1652,N_1622,N_1603);
nand U1653 (N_1653,N_1633,N_1647);
nand U1654 (N_1654,N_1607,N_1621);
or U1655 (N_1655,N_1635,N_1612);
nand U1656 (N_1656,N_1602,N_1628);
and U1657 (N_1657,N_1631,N_1616);
and U1658 (N_1658,N_1604,N_1613);
nand U1659 (N_1659,N_1609,N_1610);
or U1660 (N_1660,N_1637,N_1623);
and U1661 (N_1661,N_1626,N_1645);
or U1662 (N_1662,N_1643,N_1615);
and U1663 (N_1663,N_1649,N_1640);
or U1664 (N_1664,N_1620,N_1630);
or U1665 (N_1665,N_1639,N_1605);
nand U1666 (N_1666,N_1629,N_1618);
or U1667 (N_1667,N_1636,N_1646);
or U1668 (N_1668,N_1606,N_1627);
nand U1669 (N_1669,N_1624,N_1644);
and U1670 (N_1670,N_1608,N_1648);
nor U1671 (N_1671,N_1619,N_1634);
or U1672 (N_1672,N_1600,N_1641);
nand U1673 (N_1673,N_1611,N_1617);
or U1674 (N_1674,N_1642,N_1625);
nand U1675 (N_1675,N_1620,N_1641);
nand U1676 (N_1676,N_1604,N_1617);
or U1677 (N_1677,N_1622,N_1610);
or U1678 (N_1678,N_1623,N_1642);
nand U1679 (N_1679,N_1631,N_1636);
or U1680 (N_1680,N_1608,N_1637);
nor U1681 (N_1681,N_1644,N_1645);
nand U1682 (N_1682,N_1637,N_1640);
nand U1683 (N_1683,N_1636,N_1617);
nor U1684 (N_1684,N_1625,N_1614);
nor U1685 (N_1685,N_1639,N_1638);
or U1686 (N_1686,N_1629,N_1601);
or U1687 (N_1687,N_1644,N_1601);
or U1688 (N_1688,N_1627,N_1629);
nor U1689 (N_1689,N_1649,N_1642);
nand U1690 (N_1690,N_1634,N_1604);
or U1691 (N_1691,N_1604,N_1641);
or U1692 (N_1692,N_1631,N_1634);
nor U1693 (N_1693,N_1619,N_1636);
or U1694 (N_1694,N_1646,N_1617);
and U1695 (N_1695,N_1631,N_1641);
and U1696 (N_1696,N_1631,N_1603);
nor U1697 (N_1697,N_1608,N_1635);
nand U1698 (N_1698,N_1606,N_1649);
nand U1699 (N_1699,N_1645,N_1614);
nor U1700 (N_1700,N_1690,N_1685);
nand U1701 (N_1701,N_1665,N_1698);
or U1702 (N_1702,N_1651,N_1664);
nand U1703 (N_1703,N_1674,N_1696);
and U1704 (N_1704,N_1678,N_1683);
and U1705 (N_1705,N_1677,N_1662);
nor U1706 (N_1706,N_1661,N_1657);
or U1707 (N_1707,N_1682,N_1684);
nand U1708 (N_1708,N_1671,N_1652);
or U1709 (N_1709,N_1658,N_1656);
nor U1710 (N_1710,N_1666,N_1688);
or U1711 (N_1711,N_1692,N_1654);
nor U1712 (N_1712,N_1660,N_1669);
nor U1713 (N_1713,N_1686,N_1679);
nand U1714 (N_1714,N_1659,N_1694);
nor U1715 (N_1715,N_1655,N_1681);
nand U1716 (N_1716,N_1687,N_1697);
nor U1717 (N_1717,N_1695,N_1693);
xnor U1718 (N_1718,N_1650,N_1699);
and U1719 (N_1719,N_1663,N_1672);
nor U1720 (N_1720,N_1667,N_1673);
xor U1721 (N_1721,N_1689,N_1668);
nor U1722 (N_1722,N_1676,N_1653);
and U1723 (N_1723,N_1670,N_1680);
and U1724 (N_1724,N_1675,N_1691);
nor U1725 (N_1725,N_1678,N_1664);
nor U1726 (N_1726,N_1694,N_1688);
nand U1727 (N_1727,N_1672,N_1671);
nor U1728 (N_1728,N_1673,N_1678);
nor U1729 (N_1729,N_1656,N_1650);
nor U1730 (N_1730,N_1668,N_1665);
and U1731 (N_1731,N_1696,N_1684);
or U1732 (N_1732,N_1658,N_1661);
nor U1733 (N_1733,N_1666,N_1656);
nand U1734 (N_1734,N_1650,N_1675);
and U1735 (N_1735,N_1651,N_1672);
nand U1736 (N_1736,N_1685,N_1667);
or U1737 (N_1737,N_1656,N_1686);
nor U1738 (N_1738,N_1689,N_1660);
and U1739 (N_1739,N_1652,N_1691);
nand U1740 (N_1740,N_1687,N_1694);
nor U1741 (N_1741,N_1663,N_1666);
and U1742 (N_1742,N_1683,N_1698);
or U1743 (N_1743,N_1672,N_1683);
nand U1744 (N_1744,N_1672,N_1654);
nand U1745 (N_1745,N_1680,N_1656);
or U1746 (N_1746,N_1697,N_1652);
and U1747 (N_1747,N_1652,N_1667);
or U1748 (N_1748,N_1677,N_1654);
or U1749 (N_1749,N_1652,N_1669);
or U1750 (N_1750,N_1743,N_1715);
nand U1751 (N_1751,N_1742,N_1712);
nand U1752 (N_1752,N_1735,N_1721);
and U1753 (N_1753,N_1720,N_1749);
and U1754 (N_1754,N_1710,N_1744);
nand U1755 (N_1755,N_1701,N_1700);
and U1756 (N_1756,N_1724,N_1737);
and U1757 (N_1757,N_1708,N_1707);
and U1758 (N_1758,N_1727,N_1716);
and U1759 (N_1759,N_1732,N_1705);
and U1760 (N_1760,N_1746,N_1729);
nand U1761 (N_1761,N_1726,N_1706);
nand U1762 (N_1762,N_1733,N_1725);
or U1763 (N_1763,N_1734,N_1748);
nor U1764 (N_1764,N_1709,N_1745);
and U1765 (N_1765,N_1747,N_1717);
nor U1766 (N_1766,N_1719,N_1722);
nor U1767 (N_1767,N_1740,N_1730);
nor U1768 (N_1768,N_1702,N_1736);
and U1769 (N_1769,N_1738,N_1711);
or U1770 (N_1770,N_1718,N_1704);
nand U1771 (N_1771,N_1728,N_1731);
nand U1772 (N_1772,N_1713,N_1703);
nor U1773 (N_1773,N_1741,N_1739);
and U1774 (N_1774,N_1723,N_1714);
nand U1775 (N_1775,N_1745,N_1731);
or U1776 (N_1776,N_1731,N_1713);
and U1777 (N_1777,N_1738,N_1705);
and U1778 (N_1778,N_1703,N_1744);
and U1779 (N_1779,N_1700,N_1719);
and U1780 (N_1780,N_1747,N_1729);
and U1781 (N_1781,N_1742,N_1703);
nand U1782 (N_1782,N_1706,N_1710);
xnor U1783 (N_1783,N_1734,N_1725);
nand U1784 (N_1784,N_1713,N_1744);
and U1785 (N_1785,N_1731,N_1737);
or U1786 (N_1786,N_1740,N_1731);
nand U1787 (N_1787,N_1709,N_1737);
and U1788 (N_1788,N_1730,N_1728);
nand U1789 (N_1789,N_1707,N_1701);
and U1790 (N_1790,N_1743,N_1722);
nor U1791 (N_1791,N_1738,N_1714);
nand U1792 (N_1792,N_1716,N_1737);
or U1793 (N_1793,N_1711,N_1703);
nor U1794 (N_1794,N_1723,N_1718);
nand U1795 (N_1795,N_1703,N_1743);
or U1796 (N_1796,N_1739,N_1716);
and U1797 (N_1797,N_1722,N_1708);
or U1798 (N_1798,N_1727,N_1726);
nor U1799 (N_1799,N_1712,N_1700);
nand U1800 (N_1800,N_1777,N_1759);
and U1801 (N_1801,N_1766,N_1789);
or U1802 (N_1802,N_1763,N_1783);
nor U1803 (N_1803,N_1768,N_1758);
and U1804 (N_1804,N_1778,N_1774);
or U1805 (N_1805,N_1797,N_1793);
and U1806 (N_1806,N_1755,N_1761);
or U1807 (N_1807,N_1751,N_1792);
or U1808 (N_1808,N_1787,N_1773);
or U1809 (N_1809,N_1785,N_1772);
and U1810 (N_1810,N_1769,N_1786);
and U1811 (N_1811,N_1796,N_1756);
nand U1812 (N_1812,N_1760,N_1765);
nand U1813 (N_1813,N_1764,N_1770);
and U1814 (N_1814,N_1799,N_1784);
nand U1815 (N_1815,N_1798,N_1791);
or U1816 (N_1816,N_1781,N_1762);
nand U1817 (N_1817,N_1782,N_1752);
nor U1818 (N_1818,N_1750,N_1779);
and U1819 (N_1819,N_1790,N_1753);
or U1820 (N_1820,N_1794,N_1795);
nand U1821 (N_1821,N_1757,N_1775);
nand U1822 (N_1822,N_1788,N_1780);
and U1823 (N_1823,N_1767,N_1771);
or U1824 (N_1824,N_1754,N_1776);
or U1825 (N_1825,N_1798,N_1756);
or U1826 (N_1826,N_1757,N_1774);
nand U1827 (N_1827,N_1763,N_1771);
nand U1828 (N_1828,N_1750,N_1769);
nand U1829 (N_1829,N_1770,N_1775);
or U1830 (N_1830,N_1758,N_1772);
nor U1831 (N_1831,N_1790,N_1771);
nand U1832 (N_1832,N_1761,N_1758);
and U1833 (N_1833,N_1755,N_1799);
and U1834 (N_1834,N_1762,N_1760);
and U1835 (N_1835,N_1795,N_1789);
and U1836 (N_1836,N_1787,N_1764);
or U1837 (N_1837,N_1783,N_1771);
nor U1838 (N_1838,N_1797,N_1762);
nor U1839 (N_1839,N_1763,N_1758);
or U1840 (N_1840,N_1766,N_1762);
nand U1841 (N_1841,N_1752,N_1798);
nand U1842 (N_1842,N_1752,N_1791);
or U1843 (N_1843,N_1786,N_1756);
xnor U1844 (N_1844,N_1788,N_1751);
xnor U1845 (N_1845,N_1755,N_1766);
or U1846 (N_1846,N_1765,N_1774);
nor U1847 (N_1847,N_1779,N_1777);
xnor U1848 (N_1848,N_1753,N_1774);
xor U1849 (N_1849,N_1760,N_1775);
and U1850 (N_1850,N_1822,N_1838);
and U1851 (N_1851,N_1843,N_1825);
and U1852 (N_1852,N_1804,N_1845);
or U1853 (N_1853,N_1814,N_1811);
or U1854 (N_1854,N_1837,N_1803);
nor U1855 (N_1855,N_1817,N_1810);
or U1856 (N_1856,N_1808,N_1832);
and U1857 (N_1857,N_1848,N_1847);
nor U1858 (N_1858,N_1813,N_1849);
or U1859 (N_1859,N_1828,N_1835);
nand U1860 (N_1860,N_1821,N_1836);
nor U1861 (N_1861,N_1826,N_1846);
and U1862 (N_1862,N_1844,N_1841);
or U1863 (N_1863,N_1809,N_1842);
or U1864 (N_1864,N_1818,N_1816);
nand U1865 (N_1865,N_1802,N_1801);
and U1866 (N_1866,N_1829,N_1824);
or U1867 (N_1867,N_1827,N_1806);
nor U1868 (N_1868,N_1815,N_1805);
nor U1869 (N_1869,N_1820,N_1812);
nand U1870 (N_1870,N_1834,N_1800);
xor U1871 (N_1871,N_1823,N_1839);
xor U1872 (N_1872,N_1840,N_1819);
nor U1873 (N_1873,N_1830,N_1831);
and U1874 (N_1874,N_1833,N_1807);
and U1875 (N_1875,N_1800,N_1826);
or U1876 (N_1876,N_1820,N_1809);
nor U1877 (N_1877,N_1844,N_1834);
nor U1878 (N_1878,N_1826,N_1834);
nand U1879 (N_1879,N_1800,N_1819);
and U1880 (N_1880,N_1838,N_1821);
xnor U1881 (N_1881,N_1815,N_1809);
xor U1882 (N_1882,N_1832,N_1807);
and U1883 (N_1883,N_1814,N_1837);
or U1884 (N_1884,N_1835,N_1843);
and U1885 (N_1885,N_1817,N_1847);
nor U1886 (N_1886,N_1810,N_1818);
or U1887 (N_1887,N_1833,N_1803);
and U1888 (N_1888,N_1846,N_1838);
and U1889 (N_1889,N_1810,N_1805);
xnor U1890 (N_1890,N_1826,N_1835);
nor U1891 (N_1891,N_1835,N_1842);
nand U1892 (N_1892,N_1841,N_1829);
and U1893 (N_1893,N_1846,N_1832);
or U1894 (N_1894,N_1837,N_1834);
or U1895 (N_1895,N_1801,N_1809);
nand U1896 (N_1896,N_1831,N_1819);
nor U1897 (N_1897,N_1815,N_1836);
nand U1898 (N_1898,N_1829,N_1807);
and U1899 (N_1899,N_1821,N_1812);
nor U1900 (N_1900,N_1858,N_1890);
or U1901 (N_1901,N_1869,N_1862);
and U1902 (N_1902,N_1891,N_1850);
nand U1903 (N_1903,N_1893,N_1899);
nor U1904 (N_1904,N_1884,N_1879);
or U1905 (N_1905,N_1883,N_1878);
or U1906 (N_1906,N_1896,N_1894);
nand U1907 (N_1907,N_1871,N_1897);
or U1908 (N_1908,N_1885,N_1889);
nor U1909 (N_1909,N_1887,N_1873);
or U1910 (N_1910,N_1856,N_1866);
nand U1911 (N_1911,N_1854,N_1860);
nor U1912 (N_1912,N_1874,N_1892);
nand U1913 (N_1913,N_1852,N_1861);
nor U1914 (N_1914,N_1870,N_1876);
or U1915 (N_1915,N_1881,N_1875);
nor U1916 (N_1916,N_1872,N_1863);
or U1917 (N_1917,N_1882,N_1851);
or U1918 (N_1918,N_1864,N_1888);
nor U1919 (N_1919,N_1898,N_1865);
nand U1920 (N_1920,N_1857,N_1895);
nand U1921 (N_1921,N_1880,N_1877);
or U1922 (N_1922,N_1867,N_1853);
nor U1923 (N_1923,N_1868,N_1859);
nand U1924 (N_1924,N_1886,N_1855);
nor U1925 (N_1925,N_1878,N_1857);
nand U1926 (N_1926,N_1866,N_1887);
and U1927 (N_1927,N_1872,N_1858);
nor U1928 (N_1928,N_1864,N_1854);
or U1929 (N_1929,N_1879,N_1869);
nand U1930 (N_1930,N_1861,N_1856);
or U1931 (N_1931,N_1860,N_1879);
or U1932 (N_1932,N_1873,N_1899);
nor U1933 (N_1933,N_1875,N_1892);
nor U1934 (N_1934,N_1862,N_1877);
or U1935 (N_1935,N_1873,N_1868);
nor U1936 (N_1936,N_1890,N_1850);
or U1937 (N_1937,N_1862,N_1873);
nor U1938 (N_1938,N_1888,N_1894);
and U1939 (N_1939,N_1879,N_1888);
nor U1940 (N_1940,N_1868,N_1865);
nor U1941 (N_1941,N_1858,N_1880);
xor U1942 (N_1942,N_1893,N_1851);
nor U1943 (N_1943,N_1872,N_1885);
nand U1944 (N_1944,N_1871,N_1850);
and U1945 (N_1945,N_1878,N_1874);
or U1946 (N_1946,N_1873,N_1852);
or U1947 (N_1947,N_1877,N_1869);
nand U1948 (N_1948,N_1898,N_1876);
nand U1949 (N_1949,N_1886,N_1896);
xnor U1950 (N_1950,N_1919,N_1922);
and U1951 (N_1951,N_1930,N_1928);
nor U1952 (N_1952,N_1927,N_1909);
and U1953 (N_1953,N_1916,N_1942);
or U1954 (N_1954,N_1915,N_1941);
xnor U1955 (N_1955,N_1918,N_1939);
nor U1956 (N_1956,N_1949,N_1914);
or U1957 (N_1957,N_1907,N_1901);
and U1958 (N_1958,N_1905,N_1917);
nor U1959 (N_1959,N_1944,N_1912);
nand U1960 (N_1960,N_1904,N_1908);
and U1961 (N_1961,N_1929,N_1920);
nand U1962 (N_1962,N_1924,N_1902);
and U1963 (N_1963,N_1935,N_1932);
nand U1964 (N_1964,N_1910,N_1903);
or U1965 (N_1965,N_1945,N_1948);
and U1966 (N_1966,N_1937,N_1900);
nand U1967 (N_1967,N_1926,N_1947);
nor U1968 (N_1968,N_1906,N_1936);
and U1969 (N_1969,N_1938,N_1940);
nand U1970 (N_1970,N_1911,N_1934);
nor U1971 (N_1971,N_1921,N_1923);
nand U1972 (N_1972,N_1913,N_1943);
or U1973 (N_1973,N_1933,N_1925);
nor U1974 (N_1974,N_1946,N_1931);
nor U1975 (N_1975,N_1935,N_1943);
nand U1976 (N_1976,N_1934,N_1928);
or U1977 (N_1977,N_1932,N_1915);
nor U1978 (N_1978,N_1940,N_1934);
or U1979 (N_1979,N_1929,N_1933);
nor U1980 (N_1980,N_1905,N_1920);
nor U1981 (N_1981,N_1912,N_1905);
or U1982 (N_1982,N_1924,N_1922);
xor U1983 (N_1983,N_1923,N_1924);
or U1984 (N_1984,N_1935,N_1903);
nand U1985 (N_1985,N_1937,N_1908);
and U1986 (N_1986,N_1927,N_1920);
nand U1987 (N_1987,N_1915,N_1927);
nand U1988 (N_1988,N_1932,N_1946);
xor U1989 (N_1989,N_1942,N_1900);
or U1990 (N_1990,N_1900,N_1920);
and U1991 (N_1991,N_1947,N_1904);
and U1992 (N_1992,N_1934,N_1904);
and U1993 (N_1993,N_1949,N_1916);
nand U1994 (N_1994,N_1921,N_1907);
or U1995 (N_1995,N_1905,N_1901);
or U1996 (N_1996,N_1922,N_1928);
nor U1997 (N_1997,N_1909,N_1941);
nand U1998 (N_1998,N_1934,N_1925);
and U1999 (N_1999,N_1904,N_1933);
or U2000 (N_2000,N_1952,N_1983);
or U2001 (N_2001,N_1993,N_1963);
and U2002 (N_2002,N_1970,N_1954);
and U2003 (N_2003,N_1955,N_1977);
nor U2004 (N_2004,N_1960,N_1972);
and U2005 (N_2005,N_1976,N_1978);
or U2006 (N_2006,N_1981,N_1961);
and U2007 (N_2007,N_1958,N_1992);
nand U2008 (N_2008,N_1991,N_1950);
and U2009 (N_2009,N_1965,N_1956);
or U2010 (N_2010,N_1988,N_1980);
and U2011 (N_2011,N_1985,N_1964);
nand U2012 (N_2012,N_1984,N_1953);
or U2013 (N_2013,N_1966,N_1971);
and U2014 (N_2014,N_1995,N_1973);
nand U2015 (N_2015,N_1967,N_1996);
and U2016 (N_2016,N_1959,N_1999);
nor U2017 (N_2017,N_1957,N_1962);
nand U2018 (N_2018,N_1986,N_1994);
nor U2019 (N_2019,N_1989,N_1987);
nor U2020 (N_2020,N_1969,N_1975);
or U2021 (N_2021,N_1990,N_1951);
nor U2022 (N_2022,N_1998,N_1982);
or U2023 (N_2023,N_1979,N_1997);
nor U2024 (N_2024,N_1974,N_1968);
nand U2025 (N_2025,N_1988,N_1986);
nand U2026 (N_2026,N_1974,N_1998);
or U2027 (N_2027,N_1986,N_1993);
and U2028 (N_2028,N_1974,N_1986);
and U2029 (N_2029,N_1970,N_1959);
or U2030 (N_2030,N_1978,N_1986);
nor U2031 (N_2031,N_1982,N_1958);
nand U2032 (N_2032,N_1955,N_1982);
and U2033 (N_2033,N_1995,N_1985);
nand U2034 (N_2034,N_1985,N_1955);
and U2035 (N_2035,N_1996,N_1993);
nand U2036 (N_2036,N_1983,N_1958);
nand U2037 (N_2037,N_1964,N_1959);
and U2038 (N_2038,N_1960,N_1985);
and U2039 (N_2039,N_1971,N_1981);
and U2040 (N_2040,N_1995,N_1965);
or U2041 (N_2041,N_1984,N_1960);
or U2042 (N_2042,N_1989,N_1991);
nor U2043 (N_2043,N_1981,N_1970);
and U2044 (N_2044,N_1970,N_1972);
or U2045 (N_2045,N_1971,N_1967);
and U2046 (N_2046,N_1953,N_1957);
nor U2047 (N_2047,N_1975,N_1997);
and U2048 (N_2048,N_1989,N_1968);
xor U2049 (N_2049,N_1962,N_1997);
nor U2050 (N_2050,N_2040,N_2031);
nand U2051 (N_2051,N_2005,N_2024);
nand U2052 (N_2052,N_2039,N_2000);
or U2053 (N_2053,N_2018,N_2010);
nand U2054 (N_2054,N_2049,N_2032);
nand U2055 (N_2055,N_2033,N_2016);
and U2056 (N_2056,N_2046,N_2035);
or U2057 (N_2057,N_2022,N_2044);
nand U2058 (N_2058,N_2043,N_2002);
or U2059 (N_2059,N_2034,N_2023);
nor U2060 (N_2060,N_2047,N_2026);
nand U2061 (N_2061,N_2007,N_2041);
nor U2062 (N_2062,N_2036,N_2011);
or U2063 (N_2063,N_2042,N_2037);
nand U2064 (N_2064,N_2004,N_2027);
nand U2065 (N_2065,N_2030,N_2020);
or U2066 (N_2066,N_2021,N_2013);
nor U2067 (N_2067,N_2045,N_2017);
nor U2068 (N_2068,N_2006,N_2028);
or U2069 (N_2069,N_2014,N_2001);
or U2070 (N_2070,N_2008,N_2038);
nor U2071 (N_2071,N_2012,N_2003);
or U2072 (N_2072,N_2019,N_2015);
nand U2073 (N_2073,N_2048,N_2009);
and U2074 (N_2074,N_2025,N_2029);
nor U2075 (N_2075,N_2020,N_2048);
and U2076 (N_2076,N_2037,N_2001);
nand U2077 (N_2077,N_2029,N_2045);
nor U2078 (N_2078,N_2036,N_2025);
and U2079 (N_2079,N_2017,N_2028);
nor U2080 (N_2080,N_2019,N_2040);
nor U2081 (N_2081,N_2046,N_2017);
and U2082 (N_2082,N_2030,N_2036);
and U2083 (N_2083,N_2004,N_2033);
nand U2084 (N_2084,N_2041,N_2034);
nor U2085 (N_2085,N_2033,N_2009);
and U2086 (N_2086,N_2026,N_2009);
nor U2087 (N_2087,N_2009,N_2042);
or U2088 (N_2088,N_2049,N_2045);
or U2089 (N_2089,N_2027,N_2010);
nor U2090 (N_2090,N_2036,N_2018);
nor U2091 (N_2091,N_2026,N_2040);
nand U2092 (N_2092,N_2047,N_2006);
nor U2093 (N_2093,N_2029,N_2009);
and U2094 (N_2094,N_2014,N_2020);
and U2095 (N_2095,N_2048,N_2021);
xnor U2096 (N_2096,N_2030,N_2026);
nor U2097 (N_2097,N_2009,N_2004);
or U2098 (N_2098,N_2047,N_2044);
nor U2099 (N_2099,N_2020,N_2018);
or U2100 (N_2100,N_2050,N_2056);
and U2101 (N_2101,N_2053,N_2075);
and U2102 (N_2102,N_2074,N_2093);
nor U2103 (N_2103,N_2062,N_2089);
nand U2104 (N_2104,N_2069,N_2083);
nor U2105 (N_2105,N_2066,N_2095);
nor U2106 (N_2106,N_2063,N_2094);
nor U2107 (N_2107,N_2059,N_2070);
and U2108 (N_2108,N_2057,N_2051);
and U2109 (N_2109,N_2068,N_2078);
nand U2110 (N_2110,N_2076,N_2054);
xor U2111 (N_2111,N_2099,N_2092);
nand U2112 (N_2112,N_2064,N_2067);
nor U2113 (N_2113,N_2080,N_2088);
nand U2114 (N_2114,N_2097,N_2082);
xnor U2115 (N_2115,N_2090,N_2060);
nor U2116 (N_2116,N_2098,N_2079);
or U2117 (N_2117,N_2065,N_2081);
or U2118 (N_2118,N_2072,N_2085);
or U2119 (N_2119,N_2058,N_2071);
nand U2120 (N_2120,N_2096,N_2052);
nand U2121 (N_2121,N_2087,N_2055);
nor U2122 (N_2122,N_2084,N_2073);
nand U2123 (N_2123,N_2086,N_2077);
and U2124 (N_2124,N_2091,N_2061);
and U2125 (N_2125,N_2090,N_2093);
and U2126 (N_2126,N_2084,N_2080);
nand U2127 (N_2127,N_2088,N_2076);
or U2128 (N_2128,N_2053,N_2056);
nand U2129 (N_2129,N_2064,N_2069);
nor U2130 (N_2130,N_2076,N_2092);
nor U2131 (N_2131,N_2070,N_2089);
and U2132 (N_2132,N_2066,N_2055);
nand U2133 (N_2133,N_2065,N_2073);
nor U2134 (N_2134,N_2089,N_2061);
nand U2135 (N_2135,N_2096,N_2064);
or U2136 (N_2136,N_2067,N_2081);
and U2137 (N_2137,N_2084,N_2099);
and U2138 (N_2138,N_2054,N_2094);
or U2139 (N_2139,N_2076,N_2051);
nor U2140 (N_2140,N_2089,N_2055);
or U2141 (N_2141,N_2099,N_2074);
nand U2142 (N_2142,N_2072,N_2090);
and U2143 (N_2143,N_2062,N_2067);
and U2144 (N_2144,N_2092,N_2073);
and U2145 (N_2145,N_2063,N_2062);
and U2146 (N_2146,N_2076,N_2070);
nor U2147 (N_2147,N_2083,N_2099);
nand U2148 (N_2148,N_2064,N_2060);
or U2149 (N_2149,N_2051,N_2077);
and U2150 (N_2150,N_2113,N_2146);
nor U2151 (N_2151,N_2109,N_2107);
nand U2152 (N_2152,N_2123,N_2130);
and U2153 (N_2153,N_2120,N_2140);
and U2154 (N_2154,N_2148,N_2108);
nand U2155 (N_2155,N_2135,N_2106);
nor U2156 (N_2156,N_2132,N_2118);
or U2157 (N_2157,N_2134,N_2124);
or U2158 (N_2158,N_2121,N_2104);
and U2159 (N_2159,N_2102,N_2145);
nand U2160 (N_2160,N_2139,N_2126);
or U2161 (N_2161,N_2111,N_2129);
nand U2162 (N_2162,N_2138,N_2143);
or U2163 (N_2163,N_2141,N_2136);
nor U2164 (N_2164,N_2128,N_2122);
and U2165 (N_2165,N_2147,N_2127);
nand U2166 (N_2166,N_2137,N_2103);
nand U2167 (N_2167,N_2149,N_2142);
nor U2168 (N_2168,N_2133,N_2100);
and U2169 (N_2169,N_2116,N_2125);
nor U2170 (N_2170,N_2112,N_2131);
nor U2171 (N_2171,N_2114,N_2110);
nor U2172 (N_2172,N_2144,N_2101);
nor U2173 (N_2173,N_2105,N_2117);
nand U2174 (N_2174,N_2115,N_2119);
xnor U2175 (N_2175,N_2130,N_2149);
nor U2176 (N_2176,N_2137,N_2140);
and U2177 (N_2177,N_2122,N_2108);
nor U2178 (N_2178,N_2119,N_2128);
or U2179 (N_2179,N_2108,N_2123);
nand U2180 (N_2180,N_2124,N_2110);
nor U2181 (N_2181,N_2146,N_2119);
or U2182 (N_2182,N_2116,N_2121);
nor U2183 (N_2183,N_2149,N_2115);
and U2184 (N_2184,N_2103,N_2118);
nand U2185 (N_2185,N_2131,N_2106);
or U2186 (N_2186,N_2118,N_2111);
and U2187 (N_2187,N_2119,N_2147);
xor U2188 (N_2188,N_2123,N_2133);
nor U2189 (N_2189,N_2115,N_2110);
and U2190 (N_2190,N_2116,N_2128);
nand U2191 (N_2191,N_2100,N_2134);
nor U2192 (N_2192,N_2122,N_2142);
nand U2193 (N_2193,N_2113,N_2115);
or U2194 (N_2194,N_2146,N_2139);
nand U2195 (N_2195,N_2106,N_2122);
and U2196 (N_2196,N_2114,N_2120);
nand U2197 (N_2197,N_2132,N_2102);
or U2198 (N_2198,N_2146,N_2149);
nand U2199 (N_2199,N_2103,N_2129);
or U2200 (N_2200,N_2175,N_2196);
or U2201 (N_2201,N_2181,N_2179);
or U2202 (N_2202,N_2153,N_2194);
nand U2203 (N_2203,N_2193,N_2190);
or U2204 (N_2204,N_2154,N_2169);
nor U2205 (N_2205,N_2185,N_2159);
or U2206 (N_2206,N_2187,N_2168);
and U2207 (N_2207,N_2170,N_2186);
or U2208 (N_2208,N_2160,N_2177);
and U2209 (N_2209,N_2157,N_2174);
nand U2210 (N_2210,N_2198,N_2173);
nand U2211 (N_2211,N_2164,N_2167);
nor U2212 (N_2212,N_2199,N_2191);
nand U2213 (N_2213,N_2197,N_2178);
nand U2214 (N_2214,N_2182,N_2151);
nor U2215 (N_2215,N_2195,N_2189);
xor U2216 (N_2216,N_2163,N_2180);
nand U2217 (N_2217,N_2171,N_2166);
or U2218 (N_2218,N_2150,N_2176);
nor U2219 (N_2219,N_2162,N_2158);
nand U2220 (N_2220,N_2188,N_2156);
and U2221 (N_2221,N_2152,N_2192);
nand U2222 (N_2222,N_2183,N_2184);
or U2223 (N_2223,N_2172,N_2165);
nor U2224 (N_2224,N_2155,N_2161);
nor U2225 (N_2225,N_2184,N_2198);
or U2226 (N_2226,N_2189,N_2159);
and U2227 (N_2227,N_2194,N_2193);
and U2228 (N_2228,N_2168,N_2199);
nor U2229 (N_2229,N_2184,N_2153);
nor U2230 (N_2230,N_2188,N_2198);
and U2231 (N_2231,N_2199,N_2176);
nand U2232 (N_2232,N_2188,N_2170);
nor U2233 (N_2233,N_2192,N_2178);
or U2234 (N_2234,N_2194,N_2182);
nor U2235 (N_2235,N_2194,N_2166);
or U2236 (N_2236,N_2156,N_2154);
and U2237 (N_2237,N_2160,N_2178);
nor U2238 (N_2238,N_2189,N_2186);
and U2239 (N_2239,N_2192,N_2183);
or U2240 (N_2240,N_2187,N_2174);
nor U2241 (N_2241,N_2171,N_2198);
or U2242 (N_2242,N_2151,N_2181);
and U2243 (N_2243,N_2162,N_2176);
xnor U2244 (N_2244,N_2177,N_2150);
or U2245 (N_2245,N_2175,N_2168);
or U2246 (N_2246,N_2156,N_2181);
nor U2247 (N_2247,N_2175,N_2164);
nand U2248 (N_2248,N_2199,N_2172);
nand U2249 (N_2249,N_2189,N_2184);
nand U2250 (N_2250,N_2217,N_2243);
nand U2251 (N_2251,N_2244,N_2237);
or U2252 (N_2252,N_2234,N_2231);
nor U2253 (N_2253,N_2201,N_2223);
or U2254 (N_2254,N_2240,N_2228);
nand U2255 (N_2255,N_2236,N_2232);
nor U2256 (N_2256,N_2212,N_2200);
xor U2257 (N_2257,N_2226,N_2211);
nand U2258 (N_2258,N_2235,N_2218);
and U2259 (N_2259,N_2204,N_2242);
and U2260 (N_2260,N_2215,N_2220);
nand U2261 (N_2261,N_2225,N_2205);
nand U2262 (N_2262,N_2249,N_2245);
or U2263 (N_2263,N_2214,N_2239);
nand U2264 (N_2264,N_2247,N_2209);
nor U2265 (N_2265,N_2202,N_2248);
nand U2266 (N_2266,N_2222,N_2238);
nor U2267 (N_2267,N_2219,N_2216);
nand U2268 (N_2268,N_2206,N_2227);
or U2269 (N_2269,N_2224,N_2233);
or U2270 (N_2270,N_2246,N_2210);
or U2271 (N_2271,N_2230,N_2229);
nand U2272 (N_2272,N_2221,N_2203);
xor U2273 (N_2273,N_2207,N_2213);
or U2274 (N_2274,N_2241,N_2208);
and U2275 (N_2275,N_2220,N_2229);
and U2276 (N_2276,N_2230,N_2208);
or U2277 (N_2277,N_2232,N_2220);
or U2278 (N_2278,N_2209,N_2233);
nand U2279 (N_2279,N_2206,N_2224);
nor U2280 (N_2280,N_2241,N_2239);
and U2281 (N_2281,N_2234,N_2205);
and U2282 (N_2282,N_2234,N_2248);
and U2283 (N_2283,N_2209,N_2224);
nor U2284 (N_2284,N_2200,N_2235);
and U2285 (N_2285,N_2210,N_2241);
or U2286 (N_2286,N_2200,N_2233);
nand U2287 (N_2287,N_2212,N_2216);
nand U2288 (N_2288,N_2231,N_2248);
or U2289 (N_2289,N_2230,N_2202);
nor U2290 (N_2290,N_2237,N_2216);
and U2291 (N_2291,N_2245,N_2235);
nand U2292 (N_2292,N_2246,N_2241);
and U2293 (N_2293,N_2230,N_2232);
nor U2294 (N_2294,N_2234,N_2218);
and U2295 (N_2295,N_2204,N_2246);
nor U2296 (N_2296,N_2206,N_2217);
or U2297 (N_2297,N_2225,N_2230);
nor U2298 (N_2298,N_2244,N_2207);
nand U2299 (N_2299,N_2234,N_2243);
or U2300 (N_2300,N_2278,N_2292);
nor U2301 (N_2301,N_2289,N_2287);
or U2302 (N_2302,N_2299,N_2256);
nand U2303 (N_2303,N_2274,N_2284);
nor U2304 (N_2304,N_2266,N_2294);
nand U2305 (N_2305,N_2276,N_2270);
or U2306 (N_2306,N_2258,N_2252);
and U2307 (N_2307,N_2268,N_2280);
nor U2308 (N_2308,N_2275,N_2261);
and U2309 (N_2309,N_2296,N_2251);
or U2310 (N_2310,N_2282,N_2272);
and U2311 (N_2311,N_2288,N_2265);
nand U2312 (N_2312,N_2290,N_2254);
and U2313 (N_2313,N_2283,N_2259);
or U2314 (N_2314,N_2281,N_2271);
nor U2315 (N_2315,N_2273,N_2255);
or U2316 (N_2316,N_2297,N_2286);
or U2317 (N_2317,N_2260,N_2250);
and U2318 (N_2318,N_2269,N_2291);
or U2319 (N_2319,N_2253,N_2279);
or U2320 (N_2320,N_2293,N_2295);
or U2321 (N_2321,N_2257,N_2263);
nor U2322 (N_2322,N_2267,N_2277);
or U2323 (N_2323,N_2264,N_2285);
nor U2324 (N_2324,N_2298,N_2262);
nand U2325 (N_2325,N_2274,N_2271);
nor U2326 (N_2326,N_2275,N_2269);
nand U2327 (N_2327,N_2266,N_2285);
or U2328 (N_2328,N_2283,N_2275);
nor U2329 (N_2329,N_2289,N_2270);
nor U2330 (N_2330,N_2279,N_2256);
or U2331 (N_2331,N_2277,N_2276);
and U2332 (N_2332,N_2266,N_2267);
and U2333 (N_2333,N_2260,N_2291);
or U2334 (N_2334,N_2270,N_2269);
and U2335 (N_2335,N_2299,N_2290);
and U2336 (N_2336,N_2254,N_2299);
nand U2337 (N_2337,N_2250,N_2280);
nor U2338 (N_2338,N_2289,N_2273);
and U2339 (N_2339,N_2280,N_2274);
nor U2340 (N_2340,N_2270,N_2294);
or U2341 (N_2341,N_2290,N_2284);
or U2342 (N_2342,N_2290,N_2275);
and U2343 (N_2343,N_2250,N_2256);
nand U2344 (N_2344,N_2296,N_2269);
nand U2345 (N_2345,N_2296,N_2261);
or U2346 (N_2346,N_2289,N_2260);
and U2347 (N_2347,N_2298,N_2273);
nand U2348 (N_2348,N_2298,N_2290);
or U2349 (N_2349,N_2272,N_2296);
nor U2350 (N_2350,N_2323,N_2318);
and U2351 (N_2351,N_2334,N_2348);
nand U2352 (N_2352,N_2319,N_2321);
and U2353 (N_2353,N_2327,N_2346);
nor U2354 (N_2354,N_2310,N_2301);
or U2355 (N_2355,N_2331,N_2326);
nor U2356 (N_2356,N_2309,N_2329);
nor U2357 (N_2357,N_2316,N_2333);
nor U2358 (N_2358,N_2306,N_2328);
or U2359 (N_2359,N_2325,N_2338);
and U2360 (N_2360,N_2343,N_2315);
xor U2361 (N_2361,N_2347,N_2313);
nor U2362 (N_2362,N_2322,N_2304);
and U2363 (N_2363,N_2332,N_2342);
nor U2364 (N_2364,N_2349,N_2335);
and U2365 (N_2365,N_2307,N_2317);
or U2366 (N_2366,N_2311,N_2344);
nand U2367 (N_2367,N_2302,N_2336);
nor U2368 (N_2368,N_2330,N_2324);
nand U2369 (N_2369,N_2339,N_2341);
nor U2370 (N_2370,N_2314,N_2320);
nand U2371 (N_2371,N_2337,N_2305);
nand U2372 (N_2372,N_2300,N_2345);
nand U2373 (N_2373,N_2312,N_2308);
and U2374 (N_2374,N_2303,N_2340);
nand U2375 (N_2375,N_2342,N_2321);
nand U2376 (N_2376,N_2316,N_2345);
nand U2377 (N_2377,N_2338,N_2308);
nand U2378 (N_2378,N_2306,N_2339);
nand U2379 (N_2379,N_2314,N_2302);
nand U2380 (N_2380,N_2338,N_2317);
nand U2381 (N_2381,N_2312,N_2306);
and U2382 (N_2382,N_2305,N_2344);
and U2383 (N_2383,N_2327,N_2321);
nand U2384 (N_2384,N_2302,N_2325);
nor U2385 (N_2385,N_2313,N_2342);
xor U2386 (N_2386,N_2311,N_2343);
or U2387 (N_2387,N_2302,N_2303);
nor U2388 (N_2388,N_2333,N_2317);
or U2389 (N_2389,N_2315,N_2333);
nor U2390 (N_2390,N_2318,N_2305);
nor U2391 (N_2391,N_2333,N_2337);
nor U2392 (N_2392,N_2320,N_2322);
and U2393 (N_2393,N_2327,N_2333);
xnor U2394 (N_2394,N_2308,N_2329);
nand U2395 (N_2395,N_2310,N_2347);
and U2396 (N_2396,N_2316,N_2314);
xnor U2397 (N_2397,N_2304,N_2301);
or U2398 (N_2398,N_2335,N_2339);
nand U2399 (N_2399,N_2310,N_2318);
nor U2400 (N_2400,N_2353,N_2394);
or U2401 (N_2401,N_2371,N_2390);
or U2402 (N_2402,N_2396,N_2365);
or U2403 (N_2403,N_2381,N_2361);
nand U2404 (N_2404,N_2399,N_2352);
nand U2405 (N_2405,N_2372,N_2389);
nor U2406 (N_2406,N_2375,N_2391);
nor U2407 (N_2407,N_2383,N_2359);
nand U2408 (N_2408,N_2379,N_2377);
nand U2409 (N_2409,N_2366,N_2397);
and U2410 (N_2410,N_2370,N_2386);
nand U2411 (N_2411,N_2355,N_2356);
nand U2412 (N_2412,N_2395,N_2364);
nand U2413 (N_2413,N_2354,N_2384);
or U2414 (N_2414,N_2362,N_2374);
or U2415 (N_2415,N_2382,N_2385);
nand U2416 (N_2416,N_2378,N_2350);
nor U2417 (N_2417,N_2357,N_2387);
or U2418 (N_2418,N_2367,N_2360);
or U2419 (N_2419,N_2358,N_2388);
nand U2420 (N_2420,N_2380,N_2369);
or U2421 (N_2421,N_2393,N_2398);
nor U2422 (N_2422,N_2373,N_2351);
xor U2423 (N_2423,N_2363,N_2376);
or U2424 (N_2424,N_2368,N_2392);
and U2425 (N_2425,N_2387,N_2384);
and U2426 (N_2426,N_2398,N_2396);
or U2427 (N_2427,N_2358,N_2352);
nand U2428 (N_2428,N_2389,N_2379);
nand U2429 (N_2429,N_2360,N_2382);
and U2430 (N_2430,N_2396,N_2394);
nor U2431 (N_2431,N_2395,N_2392);
and U2432 (N_2432,N_2370,N_2353);
or U2433 (N_2433,N_2383,N_2362);
and U2434 (N_2434,N_2386,N_2360);
or U2435 (N_2435,N_2395,N_2376);
nand U2436 (N_2436,N_2390,N_2385);
and U2437 (N_2437,N_2377,N_2357);
and U2438 (N_2438,N_2373,N_2399);
and U2439 (N_2439,N_2354,N_2399);
or U2440 (N_2440,N_2394,N_2397);
nand U2441 (N_2441,N_2375,N_2397);
nand U2442 (N_2442,N_2385,N_2355);
or U2443 (N_2443,N_2368,N_2395);
or U2444 (N_2444,N_2383,N_2360);
nand U2445 (N_2445,N_2392,N_2354);
and U2446 (N_2446,N_2396,N_2383);
nor U2447 (N_2447,N_2372,N_2393);
and U2448 (N_2448,N_2358,N_2359);
nor U2449 (N_2449,N_2375,N_2393);
or U2450 (N_2450,N_2429,N_2424);
xnor U2451 (N_2451,N_2440,N_2409);
nor U2452 (N_2452,N_2420,N_2428);
or U2453 (N_2453,N_2406,N_2419);
nand U2454 (N_2454,N_2422,N_2405);
or U2455 (N_2455,N_2413,N_2441);
nand U2456 (N_2456,N_2418,N_2400);
nand U2457 (N_2457,N_2401,N_2410);
nand U2458 (N_2458,N_2403,N_2415);
nor U2459 (N_2459,N_2448,N_2425);
and U2460 (N_2460,N_2416,N_2433);
nand U2461 (N_2461,N_2435,N_2412);
xor U2462 (N_2462,N_2404,N_2445);
nor U2463 (N_2463,N_2437,N_2421);
or U2464 (N_2464,N_2432,N_2414);
or U2465 (N_2465,N_2439,N_2443);
nor U2466 (N_2466,N_2438,N_2436);
nand U2467 (N_2467,N_2442,N_2408);
nand U2468 (N_2468,N_2407,N_2427);
or U2469 (N_2469,N_2447,N_2449);
or U2470 (N_2470,N_2426,N_2402);
and U2471 (N_2471,N_2423,N_2430);
nand U2472 (N_2472,N_2434,N_2417);
or U2473 (N_2473,N_2444,N_2431);
nor U2474 (N_2474,N_2446,N_2411);
nand U2475 (N_2475,N_2438,N_2405);
or U2476 (N_2476,N_2400,N_2420);
nand U2477 (N_2477,N_2415,N_2414);
nand U2478 (N_2478,N_2408,N_2426);
nand U2479 (N_2479,N_2423,N_2440);
and U2480 (N_2480,N_2406,N_2400);
or U2481 (N_2481,N_2435,N_2449);
and U2482 (N_2482,N_2428,N_2435);
nor U2483 (N_2483,N_2437,N_2435);
nand U2484 (N_2484,N_2413,N_2448);
or U2485 (N_2485,N_2418,N_2404);
and U2486 (N_2486,N_2411,N_2406);
xor U2487 (N_2487,N_2443,N_2444);
or U2488 (N_2488,N_2403,N_2434);
and U2489 (N_2489,N_2444,N_2418);
nand U2490 (N_2490,N_2415,N_2442);
and U2491 (N_2491,N_2420,N_2402);
nand U2492 (N_2492,N_2427,N_2426);
nand U2493 (N_2493,N_2440,N_2402);
nand U2494 (N_2494,N_2422,N_2447);
or U2495 (N_2495,N_2439,N_2406);
nor U2496 (N_2496,N_2400,N_2436);
nand U2497 (N_2497,N_2409,N_2449);
and U2498 (N_2498,N_2436,N_2430);
and U2499 (N_2499,N_2436,N_2442);
nand U2500 (N_2500,N_2476,N_2462);
nand U2501 (N_2501,N_2474,N_2493);
and U2502 (N_2502,N_2480,N_2482);
nand U2503 (N_2503,N_2488,N_2485);
or U2504 (N_2504,N_2478,N_2469);
or U2505 (N_2505,N_2468,N_2492);
nand U2506 (N_2506,N_2477,N_2465);
or U2507 (N_2507,N_2471,N_2470);
or U2508 (N_2508,N_2481,N_2453);
or U2509 (N_2509,N_2466,N_2490);
or U2510 (N_2510,N_2461,N_2497);
nor U2511 (N_2511,N_2495,N_2450);
and U2512 (N_2512,N_2494,N_2458);
nand U2513 (N_2513,N_2459,N_2464);
and U2514 (N_2514,N_2455,N_2463);
xor U2515 (N_2515,N_2454,N_2472);
or U2516 (N_2516,N_2452,N_2479);
nand U2517 (N_2517,N_2498,N_2473);
nor U2518 (N_2518,N_2456,N_2483);
nor U2519 (N_2519,N_2475,N_2496);
and U2520 (N_2520,N_2451,N_2499);
nand U2521 (N_2521,N_2486,N_2457);
nand U2522 (N_2522,N_2487,N_2489);
nor U2523 (N_2523,N_2460,N_2484);
and U2524 (N_2524,N_2467,N_2491);
nand U2525 (N_2525,N_2475,N_2453);
nand U2526 (N_2526,N_2466,N_2452);
nor U2527 (N_2527,N_2463,N_2477);
or U2528 (N_2528,N_2456,N_2451);
nor U2529 (N_2529,N_2490,N_2474);
nor U2530 (N_2530,N_2498,N_2470);
nor U2531 (N_2531,N_2484,N_2497);
nor U2532 (N_2532,N_2468,N_2493);
nor U2533 (N_2533,N_2451,N_2465);
or U2534 (N_2534,N_2484,N_2478);
or U2535 (N_2535,N_2486,N_2467);
and U2536 (N_2536,N_2476,N_2479);
nor U2537 (N_2537,N_2465,N_2462);
or U2538 (N_2538,N_2466,N_2451);
or U2539 (N_2539,N_2482,N_2498);
or U2540 (N_2540,N_2494,N_2465);
or U2541 (N_2541,N_2466,N_2496);
and U2542 (N_2542,N_2471,N_2450);
nor U2543 (N_2543,N_2494,N_2472);
nor U2544 (N_2544,N_2454,N_2480);
and U2545 (N_2545,N_2481,N_2468);
or U2546 (N_2546,N_2468,N_2464);
nor U2547 (N_2547,N_2466,N_2472);
nand U2548 (N_2548,N_2454,N_2493);
or U2549 (N_2549,N_2496,N_2486);
or U2550 (N_2550,N_2534,N_2515);
and U2551 (N_2551,N_2514,N_2530);
and U2552 (N_2552,N_2548,N_2541);
and U2553 (N_2553,N_2533,N_2546);
and U2554 (N_2554,N_2529,N_2511);
or U2555 (N_2555,N_2531,N_2538);
nor U2556 (N_2556,N_2521,N_2524);
and U2557 (N_2557,N_2545,N_2523);
or U2558 (N_2558,N_2518,N_2509);
or U2559 (N_2559,N_2501,N_2536);
nand U2560 (N_2560,N_2526,N_2507);
nand U2561 (N_2561,N_2500,N_2543);
nor U2562 (N_2562,N_2519,N_2525);
nand U2563 (N_2563,N_2508,N_2528);
nor U2564 (N_2564,N_2506,N_2547);
nand U2565 (N_2565,N_2540,N_2539);
nand U2566 (N_2566,N_2513,N_2504);
nor U2567 (N_2567,N_2502,N_2503);
and U2568 (N_2568,N_2517,N_2505);
nor U2569 (N_2569,N_2549,N_2520);
and U2570 (N_2570,N_2542,N_2532);
and U2571 (N_2571,N_2527,N_2510);
and U2572 (N_2572,N_2537,N_2512);
and U2573 (N_2573,N_2522,N_2516);
nand U2574 (N_2574,N_2544,N_2535);
and U2575 (N_2575,N_2510,N_2521);
nor U2576 (N_2576,N_2504,N_2535);
nand U2577 (N_2577,N_2548,N_2529);
and U2578 (N_2578,N_2500,N_2540);
nand U2579 (N_2579,N_2517,N_2526);
or U2580 (N_2580,N_2514,N_2537);
nand U2581 (N_2581,N_2541,N_2519);
or U2582 (N_2582,N_2522,N_2523);
nand U2583 (N_2583,N_2537,N_2526);
and U2584 (N_2584,N_2525,N_2540);
nand U2585 (N_2585,N_2507,N_2534);
and U2586 (N_2586,N_2519,N_2531);
or U2587 (N_2587,N_2515,N_2512);
nor U2588 (N_2588,N_2545,N_2524);
nand U2589 (N_2589,N_2542,N_2540);
nand U2590 (N_2590,N_2524,N_2546);
nand U2591 (N_2591,N_2520,N_2531);
nor U2592 (N_2592,N_2516,N_2515);
or U2593 (N_2593,N_2510,N_2523);
and U2594 (N_2594,N_2535,N_2537);
nor U2595 (N_2595,N_2539,N_2533);
nor U2596 (N_2596,N_2500,N_2529);
or U2597 (N_2597,N_2500,N_2516);
nand U2598 (N_2598,N_2534,N_2531);
or U2599 (N_2599,N_2502,N_2517);
xor U2600 (N_2600,N_2594,N_2587);
and U2601 (N_2601,N_2589,N_2592);
nand U2602 (N_2602,N_2573,N_2555);
or U2603 (N_2603,N_2599,N_2577);
nand U2604 (N_2604,N_2552,N_2565);
nor U2605 (N_2605,N_2567,N_2576);
nor U2606 (N_2606,N_2572,N_2580);
or U2607 (N_2607,N_2557,N_2583);
nor U2608 (N_2608,N_2578,N_2561);
or U2609 (N_2609,N_2571,N_2553);
and U2610 (N_2610,N_2584,N_2563);
nand U2611 (N_2611,N_2570,N_2596);
nor U2612 (N_2612,N_2579,N_2593);
or U2613 (N_2613,N_2591,N_2564);
and U2614 (N_2614,N_2588,N_2569);
nor U2615 (N_2615,N_2559,N_2586);
nor U2616 (N_2616,N_2568,N_2581);
nand U2617 (N_2617,N_2560,N_2595);
nand U2618 (N_2618,N_2574,N_2585);
or U2619 (N_2619,N_2566,N_2551);
nand U2620 (N_2620,N_2550,N_2558);
or U2621 (N_2621,N_2556,N_2554);
or U2622 (N_2622,N_2582,N_2575);
or U2623 (N_2623,N_2590,N_2562);
xor U2624 (N_2624,N_2597,N_2598);
or U2625 (N_2625,N_2552,N_2588);
nor U2626 (N_2626,N_2570,N_2593);
or U2627 (N_2627,N_2578,N_2568);
or U2628 (N_2628,N_2579,N_2584);
and U2629 (N_2629,N_2582,N_2559);
and U2630 (N_2630,N_2552,N_2560);
or U2631 (N_2631,N_2550,N_2595);
or U2632 (N_2632,N_2593,N_2553);
or U2633 (N_2633,N_2573,N_2558);
or U2634 (N_2634,N_2566,N_2561);
nand U2635 (N_2635,N_2565,N_2564);
and U2636 (N_2636,N_2579,N_2594);
or U2637 (N_2637,N_2587,N_2574);
nand U2638 (N_2638,N_2553,N_2598);
xnor U2639 (N_2639,N_2551,N_2565);
xor U2640 (N_2640,N_2575,N_2579);
nor U2641 (N_2641,N_2562,N_2583);
or U2642 (N_2642,N_2560,N_2577);
and U2643 (N_2643,N_2552,N_2572);
or U2644 (N_2644,N_2595,N_2589);
or U2645 (N_2645,N_2593,N_2565);
nand U2646 (N_2646,N_2581,N_2588);
or U2647 (N_2647,N_2595,N_2563);
and U2648 (N_2648,N_2560,N_2568);
nand U2649 (N_2649,N_2574,N_2555);
and U2650 (N_2650,N_2603,N_2619);
nand U2651 (N_2651,N_2633,N_2616);
nor U2652 (N_2652,N_2629,N_2609);
nand U2653 (N_2653,N_2642,N_2648);
nor U2654 (N_2654,N_2611,N_2630);
and U2655 (N_2655,N_2618,N_2620);
or U2656 (N_2656,N_2649,N_2613);
nand U2657 (N_2657,N_2621,N_2610);
nand U2658 (N_2658,N_2625,N_2644);
nand U2659 (N_2659,N_2634,N_2624);
and U2660 (N_2660,N_2623,N_2637);
and U2661 (N_2661,N_2626,N_2636);
nand U2662 (N_2662,N_2632,N_2643);
xnor U2663 (N_2663,N_2639,N_2615);
nor U2664 (N_2664,N_2638,N_2631);
or U2665 (N_2665,N_2605,N_2617);
xor U2666 (N_2666,N_2607,N_2608);
and U2667 (N_2667,N_2604,N_2646);
or U2668 (N_2668,N_2647,N_2628);
or U2669 (N_2669,N_2614,N_2645);
or U2670 (N_2670,N_2640,N_2601);
nor U2671 (N_2671,N_2627,N_2600);
nor U2672 (N_2672,N_2641,N_2635);
and U2673 (N_2673,N_2622,N_2606);
and U2674 (N_2674,N_2602,N_2612);
or U2675 (N_2675,N_2619,N_2608);
nor U2676 (N_2676,N_2646,N_2625);
nor U2677 (N_2677,N_2606,N_2635);
nand U2678 (N_2678,N_2647,N_2610);
and U2679 (N_2679,N_2608,N_2642);
or U2680 (N_2680,N_2600,N_2633);
nor U2681 (N_2681,N_2613,N_2627);
nor U2682 (N_2682,N_2625,N_2635);
nor U2683 (N_2683,N_2624,N_2649);
and U2684 (N_2684,N_2601,N_2647);
nor U2685 (N_2685,N_2621,N_2600);
nand U2686 (N_2686,N_2633,N_2643);
or U2687 (N_2687,N_2635,N_2619);
and U2688 (N_2688,N_2636,N_2613);
nand U2689 (N_2689,N_2611,N_2644);
nor U2690 (N_2690,N_2602,N_2638);
nand U2691 (N_2691,N_2626,N_2635);
or U2692 (N_2692,N_2635,N_2634);
or U2693 (N_2693,N_2631,N_2647);
or U2694 (N_2694,N_2606,N_2646);
xnor U2695 (N_2695,N_2649,N_2631);
nor U2696 (N_2696,N_2617,N_2647);
xnor U2697 (N_2697,N_2626,N_2622);
nand U2698 (N_2698,N_2645,N_2629);
or U2699 (N_2699,N_2625,N_2643);
nor U2700 (N_2700,N_2666,N_2689);
nand U2701 (N_2701,N_2660,N_2673);
or U2702 (N_2702,N_2668,N_2677);
or U2703 (N_2703,N_2683,N_2685);
and U2704 (N_2704,N_2662,N_2652);
and U2705 (N_2705,N_2658,N_2664);
and U2706 (N_2706,N_2661,N_2656);
or U2707 (N_2707,N_2691,N_2671);
nand U2708 (N_2708,N_2669,N_2680);
nand U2709 (N_2709,N_2688,N_2699);
or U2710 (N_2710,N_2675,N_2657);
nor U2711 (N_2711,N_2687,N_2659);
and U2712 (N_2712,N_2670,N_2697);
nor U2713 (N_2713,N_2665,N_2667);
nand U2714 (N_2714,N_2692,N_2672);
nor U2715 (N_2715,N_2694,N_2650);
nor U2716 (N_2716,N_2684,N_2693);
and U2717 (N_2717,N_2681,N_2686);
nand U2718 (N_2718,N_2653,N_2676);
and U2719 (N_2719,N_2678,N_2654);
or U2720 (N_2720,N_2651,N_2679);
or U2721 (N_2721,N_2698,N_2682);
or U2722 (N_2722,N_2696,N_2674);
nor U2723 (N_2723,N_2695,N_2690);
or U2724 (N_2724,N_2655,N_2663);
and U2725 (N_2725,N_2699,N_2695);
or U2726 (N_2726,N_2656,N_2679);
nor U2727 (N_2727,N_2656,N_2682);
nor U2728 (N_2728,N_2687,N_2680);
nand U2729 (N_2729,N_2668,N_2673);
nand U2730 (N_2730,N_2699,N_2669);
and U2731 (N_2731,N_2656,N_2668);
and U2732 (N_2732,N_2681,N_2656);
nor U2733 (N_2733,N_2650,N_2688);
and U2734 (N_2734,N_2699,N_2691);
nor U2735 (N_2735,N_2677,N_2686);
nor U2736 (N_2736,N_2669,N_2684);
or U2737 (N_2737,N_2662,N_2682);
or U2738 (N_2738,N_2685,N_2652);
and U2739 (N_2739,N_2693,N_2655);
nand U2740 (N_2740,N_2661,N_2685);
or U2741 (N_2741,N_2692,N_2673);
and U2742 (N_2742,N_2691,N_2694);
nand U2743 (N_2743,N_2694,N_2666);
nor U2744 (N_2744,N_2693,N_2670);
and U2745 (N_2745,N_2679,N_2685);
nand U2746 (N_2746,N_2656,N_2653);
nor U2747 (N_2747,N_2665,N_2698);
or U2748 (N_2748,N_2678,N_2687);
nor U2749 (N_2749,N_2680,N_2672);
nand U2750 (N_2750,N_2747,N_2703);
or U2751 (N_2751,N_2723,N_2700);
and U2752 (N_2752,N_2749,N_2725);
and U2753 (N_2753,N_2708,N_2709);
nand U2754 (N_2754,N_2739,N_2716);
nand U2755 (N_2755,N_2718,N_2705);
xor U2756 (N_2756,N_2719,N_2724);
or U2757 (N_2757,N_2706,N_2711);
or U2758 (N_2758,N_2737,N_2731);
nor U2759 (N_2759,N_2745,N_2744);
and U2760 (N_2760,N_2728,N_2727);
and U2761 (N_2761,N_2712,N_2732);
or U2762 (N_2762,N_2717,N_2736);
and U2763 (N_2763,N_2710,N_2713);
nand U2764 (N_2764,N_2729,N_2740);
or U2765 (N_2765,N_2707,N_2721);
and U2766 (N_2766,N_2735,N_2720);
nor U2767 (N_2767,N_2738,N_2746);
nor U2768 (N_2768,N_2701,N_2733);
and U2769 (N_2769,N_2726,N_2734);
or U2770 (N_2770,N_2704,N_2741);
xnor U2771 (N_2771,N_2742,N_2702);
and U2772 (N_2772,N_2722,N_2743);
nand U2773 (N_2773,N_2730,N_2748);
nor U2774 (N_2774,N_2715,N_2714);
nand U2775 (N_2775,N_2708,N_2729);
nor U2776 (N_2776,N_2746,N_2739);
nor U2777 (N_2777,N_2715,N_2734);
or U2778 (N_2778,N_2710,N_2734);
and U2779 (N_2779,N_2745,N_2704);
nand U2780 (N_2780,N_2717,N_2726);
nor U2781 (N_2781,N_2715,N_2731);
nor U2782 (N_2782,N_2725,N_2743);
nor U2783 (N_2783,N_2733,N_2729);
nand U2784 (N_2784,N_2741,N_2727);
nor U2785 (N_2785,N_2744,N_2720);
nand U2786 (N_2786,N_2716,N_2718);
nor U2787 (N_2787,N_2707,N_2724);
and U2788 (N_2788,N_2703,N_2722);
nor U2789 (N_2789,N_2745,N_2734);
nor U2790 (N_2790,N_2745,N_2721);
or U2791 (N_2791,N_2746,N_2718);
nor U2792 (N_2792,N_2728,N_2709);
xnor U2793 (N_2793,N_2703,N_2738);
or U2794 (N_2794,N_2728,N_2722);
and U2795 (N_2795,N_2749,N_2733);
or U2796 (N_2796,N_2732,N_2702);
nor U2797 (N_2797,N_2746,N_2740);
and U2798 (N_2798,N_2704,N_2738);
nor U2799 (N_2799,N_2742,N_2743);
and U2800 (N_2800,N_2759,N_2750);
nor U2801 (N_2801,N_2787,N_2778);
nor U2802 (N_2802,N_2784,N_2773);
and U2803 (N_2803,N_2776,N_2790);
nand U2804 (N_2804,N_2753,N_2770);
and U2805 (N_2805,N_2795,N_2799);
or U2806 (N_2806,N_2792,N_2780);
nor U2807 (N_2807,N_2757,N_2754);
or U2808 (N_2808,N_2756,N_2766);
nor U2809 (N_2809,N_2774,N_2789);
or U2810 (N_2810,N_2760,N_2751);
nor U2811 (N_2811,N_2767,N_2793);
nor U2812 (N_2812,N_2761,N_2772);
nor U2813 (N_2813,N_2763,N_2797);
nor U2814 (N_2814,N_2755,N_2783);
or U2815 (N_2815,N_2781,N_2764);
or U2816 (N_2816,N_2752,N_2762);
or U2817 (N_2817,N_2769,N_2796);
or U2818 (N_2818,N_2782,N_2779);
or U2819 (N_2819,N_2798,N_2758);
or U2820 (N_2820,N_2765,N_2777);
nor U2821 (N_2821,N_2768,N_2771);
and U2822 (N_2822,N_2785,N_2794);
and U2823 (N_2823,N_2788,N_2791);
and U2824 (N_2824,N_2786,N_2775);
or U2825 (N_2825,N_2798,N_2793);
or U2826 (N_2826,N_2767,N_2771);
and U2827 (N_2827,N_2770,N_2778);
or U2828 (N_2828,N_2787,N_2771);
nand U2829 (N_2829,N_2755,N_2792);
or U2830 (N_2830,N_2769,N_2759);
or U2831 (N_2831,N_2793,N_2777);
or U2832 (N_2832,N_2762,N_2783);
nand U2833 (N_2833,N_2798,N_2772);
nand U2834 (N_2834,N_2763,N_2769);
or U2835 (N_2835,N_2764,N_2792);
nor U2836 (N_2836,N_2758,N_2785);
xor U2837 (N_2837,N_2773,N_2791);
nand U2838 (N_2838,N_2797,N_2786);
or U2839 (N_2839,N_2760,N_2764);
nor U2840 (N_2840,N_2796,N_2793);
nand U2841 (N_2841,N_2755,N_2778);
or U2842 (N_2842,N_2760,N_2762);
and U2843 (N_2843,N_2776,N_2799);
nand U2844 (N_2844,N_2774,N_2760);
nor U2845 (N_2845,N_2786,N_2779);
nor U2846 (N_2846,N_2770,N_2768);
and U2847 (N_2847,N_2761,N_2781);
nor U2848 (N_2848,N_2750,N_2784);
nand U2849 (N_2849,N_2757,N_2774);
nor U2850 (N_2850,N_2800,N_2841);
and U2851 (N_2851,N_2811,N_2806);
and U2852 (N_2852,N_2804,N_2831);
nand U2853 (N_2853,N_2822,N_2846);
and U2854 (N_2854,N_2801,N_2826);
or U2855 (N_2855,N_2844,N_2823);
nor U2856 (N_2856,N_2816,N_2821);
nand U2857 (N_2857,N_2833,N_2836);
and U2858 (N_2858,N_2848,N_2827);
nor U2859 (N_2859,N_2815,N_2809);
nor U2860 (N_2860,N_2832,N_2805);
nor U2861 (N_2861,N_2818,N_2819);
nor U2862 (N_2862,N_2847,N_2810);
nor U2863 (N_2863,N_2803,N_2807);
and U2864 (N_2864,N_2842,N_2825);
nor U2865 (N_2865,N_2838,N_2843);
and U2866 (N_2866,N_2814,N_2802);
nor U2867 (N_2867,N_2808,N_2824);
nor U2868 (N_2868,N_2820,N_2829);
or U2869 (N_2869,N_2839,N_2834);
nor U2870 (N_2870,N_2845,N_2828);
nand U2871 (N_2871,N_2830,N_2837);
nand U2872 (N_2872,N_2835,N_2817);
nand U2873 (N_2873,N_2840,N_2813);
nor U2874 (N_2874,N_2849,N_2812);
and U2875 (N_2875,N_2804,N_2849);
or U2876 (N_2876,N_2848,N_2823);
and U2877 (N_2877,N_2822,N_2824);
nand U2878 (N_2878,N_2842,N_2815);
and U2879 (N_2879,N_2843,N_2813);
and U2880 (N_2880,N_2806,N_2819);
and U2881 (N_2881,N_2803,N_2837);
nand U2882 (N_2882,N_2842,N_2813);
nand U2883 (N_2883,N_2837,N_2834);
xor U2884 (N_2884,N_2841,N_2836);
nor U2885 (N_2885,N_2833,N_2844);
and U2886 (N_2886,N_2823,N_2820);
nand U2887 (N_2887,N_2821,N_2801);
or U2888 (N_2888,N_2813,N_2816);
xnor U2889 (N_2889,N_2813,N_2800);
and U2890 (N_2890,N_2834,N_2821);
or U2891 (N_2891,N_2819,N_2843);
and U2892 (N_2892,N_2838,N_2848);
or U2893 (N_2893,N_2836,N_2817);
xnor U2894 (N_2894,N_2805,N_2844);
nor U2895 (N_2895,N_2808,N_2832);
nor U2896 (N_2896,N_2822,N_2810);
xor U2897 (N_2897,N_2802,N_2825);
nor U2898 (N_2898,N_2808,N_2813);
xnor U2899 (N_2899,N_2846,N_2839);
nand U2900 (N_2900,N_2861,N_2865);
and U2901 (N_2901,N_2885,N_2852);
and U2902 (N_2902,N_2871,N_2854);
nand U2903 (N_2903,N_2855,N_2876);
nor U2904 (N_2904,N_2856,N_2890);
xor U2905 (N_2905,N_2853,N_2898);
or U2906 (N_2906,N_2860,N_2892);
nand U2907 (N_2907,N_2896,N_2866);
nor U2908 (N_2908,N_2883,N_2880);
nand U2909 (N_2909,N_2882,N_2867);
nor U2910 (N_2910,N_2877,N_2864);
and U2911 (N_2911,N_2897,N_2858);
nand U2912 (N_2912,N_2850,N_2879);
nor U2913 (N_2913,N_2889,N_2899);
nor U2914 (N_2914,N_2881,N_2886);
nand U2915 (N_2915,N_2863,N_2851);
nand U2916 (N_2916,N_2857,N_2874);
and U2917 (N_2917,N_2894,N_2893);
or U2918 (N_2918,N_2884,N_2888);
and U2919 (N_2919,N_2869,N_2873);
nor U2920 (N_2920,N_2887,N_2872);
nor U2921 (N_2921,N_2868,N_2878);
or U2922 (N_2922,N_2859,N_2891);
or U2923 (N_2923,N_2870,N_2875);
or U2924 (N_2924,N_2862,N_2895);
or U2925 (N_2925,N_2858,N_2882);
or U2926 (N_2926,N_2858,N_2869);
and U2927 (N_2927,N_2891,N_2852);
and U2928 (N_2928,N_2871,N_2851);
nor U2929 (N_2929,N_2883,N_2863);
or U2930 (N_2930,N_2863,N_2869);
or U2931 (N_2931,N_2891,N_2892);
nor U2932 (N_2932,N_2885,N_2871);
nand U2933 (N_2933,N_2858,N_2895);
nand U2934 (N_2934,N_2896,N_2877);
and U2935 (N_2935,N_2871,N_2888);
or U2936 (N_2936,N_2861,N_2884);
nor U2937 (N_2937,N_2879,N_2860);
or U2938 (N_2938,N_2881,N_2853);
and U2939 (N_2939,N_2851,N_2865);
nand U2940 (N_2940,N_2853,N_2889);
nor U2941 (N_2941,N_2892,N_2867);
nand U2942 (N_2942,N_2861,N_2851);
nor U2943 (N_2943,N_2853,N_2875);
nand U2944 (N_2944,N_2859,N_2852);
or U2945 (N_2945,N_2856,N_2865);
and U2946 (N_2946,N_2896,N_2879);
and U2947 (N_2947,N_2854,N_2867);
or U2948 (N_2948,N_2860,N_2878);
nand U2949 (N_2949,N_2854,N_2870);
or U2950 (N_2950,N_2917,N_2933);
nand U2951 (N_2951,N_2931,N_2943);
and U2952 (N_2952,N_2949,N_2938);
nor U2953 (N_2953,N_2900,N_2920);
and U2954 (N_2954,N_2901,N_2903);
or U2955 (N_2955,N_2922,N_2935);
and U2956 (N_2956,N_2911,N_2937);
and U2957 (N_2957,N_2934,N_2944);
nor U2958 (N_2958,N_2914,N_2916);
nor U2959 (N_2959,N_2923,N_2940);
and U2960 (N_2960,N_2936,N_2939);
nor U2961 (N_2961,N_2905,N_2915);
and U2962 (N_2962,N_2928,N_2918);
nand U2963 (N_2963,N_2902,N_2932);
and U2964 (N_2964,N_2927,N_2948);
and U2965 (N_2965,N_2945,N_2946);
and U2966 (N_2966,N_2926,N_2942);
nand U2967 (N_2967,N_2921,N_2906);
or U2968 (N_2968,N_2947,N_2925);
or U2969 (N_2969,N_2924,N_2904);
nor U2970 (N_2970,N_2929,N_2930);
or U2971 (N_2971,N_2912,N_2941);
or U2972 (N_2972,N_2910,N_2919);
or U2973 (N_2973,N_2909,N_2908);
or U2974 (N_2974,N_2913,N_2907);
nor U2975 (N_2975,N_2945,N_2928);
nand U2976 (N_2976,N_2941,N_2908);
or U2977 (N_2977,N_2902,N_2919);
or U2978 (N_2978,N_2935,N_2924);
nor U2979 (N_2979,N_2914,N_2905);
nand U2980 (N_2980,N_2916,N_2931);
nor U2981 (N_2981,N_2902,N_2920);
and U2982 (N_2982,N_2907,N_2930);
nand U2983 (N_2983,N_2934,N_2949);
nand U2984 (N_2984,N_2936,N_2929);
nand U2985 (N_2985,N_2909,N_2932);
nand U2986 (N_2986,N_2911,N_2932);
or U2987 (N_2987,N_2918,N_2925);
or U2988 (N_2988,N_2912,N_2930);
and U2989 (N_2989,N_2930,N_2939);
nand U2990 (N_2990,N_2908,N_2925);
nor U2991 (N_2991,N_2932,N_2940);
nor U2992 (N_2992,N_2905,N_2934);
nor U2993 (N_2993,N_2904,N_2919);
nor U2994 (N_2994,N_2912,N_2905);
nor U2995 (N_2995,N_2915,N_2920);
and U2996 (N_2996,N_2921,N_2927);
nor U2997 (N_2997,N_2903,N_2919);
or U2998 (N_2998,N_2932,N_2943);
or U2999 (N_2999,N_2932,N_2917);
and UO_0 (O_0,N_2958,N_2986);
nor UO_1 (O_1,N_2959,N_2976);
nor UO_2 (O_2,N_2982,N_2991);
or UO_3 (O_3,N_2990,N_2979);
nand UO_4 (O_4,N_2984,N_2994);
nor UO_5 (O_5,N_2993,N_2997);
or UO_6 (O_6,N_2967,N_2980);
nand UO_7 (O_7,N_2987,N_2973);
nand UO_8 (O_8,N_2974,N_2965);
or UO_9 (O_9,N_2963,N_2988);
and UO_10 (O_10,N_2971,N_2953);
or UO_11 (O_11,N_2960,N_2964);
nor UO_12 (O_12,N_2962,N_2977);
or UO_13 (O_13,N_2952,N_2975);
nand UO_14 (O_14,N_2981,N_2996);
or UO_15 (O_15,N_2957,N_2978);
nand UO_16 (O_16,N_2972,N_2992);
or UO_17 (O_17,N_2956,N_2961);
nor UO_18 (O_18,N_2968,N_2966);
and UO_19 (O_19,N_2998,N_2983);
and UO_20 (O_20,N_2970,N_2951);
nor UO_21 (O_21,N_2995,N_2985);
or UO_22 (O_22,N_2955,N_2969);
nand UO_23 (O_23,N_2954,N_2999);
nor UO_24 (O_24,N_2950,N_2989);
nor UO_25 (O_25,N_2988,N_2983);
nand UO_26 (O_26,N_2977,N_2996);
nor UO_27 (O_27,N_2994,N_2953);
or UO_28 (O_28,N_2986,N_2952);
and UO_29 (O_29,N_2970,N_2983);
nor UO_30 (O_30,N_2988,N_2968);
nor UO_31 (O_31,N_2981,N_2954);
or UO_32 (O_32,N_2991,N_2980);
or UO_33 (O_33,N_2953,N_2993);
nor UO_34 (O_34,N_2971,N_2955);
and UO_35 (O_35,N_2972,N_2962);
and UO_36 (O_36,N_2971,N_2977);
and UO_37 (O_37,N_2989,N_2965);
and UO_38 (O_38,N_2983,N_2961);
nand UO_39 (O_39,N_2986,N_2995);
or UO_40 (O_40,N_2990,N_2983);
nand UO_41 (O_41,N_2991,N_2961);
or UO_42 (O_42,N_2988,N_2992);
nor UO_43 (O_43,N_2981,N_2985);
and UO_44 (O_44,N_2973,N_2950);
nand UO_45 (O_45,N_2972,N_2973);
and UO_46 (O_46,N_2974,N_2950);
nor UO_47 (O_47,N_2981,N_2971);
nor UO_48 (O_48,N_2996,N_2964);
and UO_49 (O_49,N_2985,N_2994);
nand UO_50 (O_50,N_2996,N_2967);
or UO_51 (O_51,N_2989,N_2973);
or UO_52 (O_52,N_2959,N_2999);
or UO_53 (O_53,N_2990,N_2975);
nand UO_54 (O_54,N_2983,N_2960);
nor UO_55 (O_55,N_2970,N_2986);
or UO_56 (O_56,N_2973,N_2975);
nor UO_57 (O_57,N_2971,N_2970);
nor UO_58 (O_58,N_2983,N_2974);
or UO_59 (O_59,N_2998,N_2989);
nand UO_60 (O_60,N_2963,N_2970);
and UO_61 (O_61,N_2968,N_2993);
nor UO_62 (O_62,N_2987,N_2980);
and UO_63 (O_63,N_2967,N_2965);
nand UO_64 (O_64,N_2990,N_2968);
nand UO_65 (O_65,N_2966,N_2992);
and UO_66 (O_66,N_2984,N_2993);
nor UO_67 (O_67,N_2994,N_2980);
nand UO_68 (O_68,N_2994,N_2976);
nor UO_69 (O_69,N_2953,N_2950);
nand UO_70 (O_70,N_2963,N_2967);
and UO_71 (O_71,N_2962,N_2993);
or UO_72 (O_72,N_2965,N_2950);
nand UO_73 (O_73,N_2987,N_2963);
and UO_74 (O_74,N_2970,N_2955);
and UO_75 (O_75,N_2976,N_2955);
and UO_76 (O_76,N_2968,N_2963);
nand UO_77 (O_77,N_2958,N_2993);
nor UO_78 (O_78,N_2994,N_2970);
and UO_79 (O_79,N_2956,N_2957);
or UO_80 (O_80,N_2960,N_2969);
and UO_81 (O_81,N_2984,N_2965);
nand UO_82 (O_82,N_2977,N_2981);
and UO_83 (O_83,N_2994,N_2963);
nand UO_84 (O_84,N_2952,N_2968);
or UO_85 (O_85,N_2964,N_2977);
nand UO_86 (O_86,N_2995,N_2980);
and UO_87 (O_87,N_2964,N_2981);
and UO_88 (O_88,N_2987,N_2959);
and UO_89 (O_89,N_2979,N_2963);
and UO_90 (O_90,N_2984,N_2966);
nor UO_91 (O_91,N_2982,N_2997);
nand UO_92 (O_92,N_2989,N_2951);
nand UO_93 (O_93,N_2960,N_2995);
and UO_94 (O_94,N_2962,N_2992);
nor UO_95 (O_95,N_2971,N_2993);
nor UO_96 (O_96,N_2984,N_2995);
nand UO_97 (O_97,N_2952,N_2960);
or UO_98 (O_98,N_2961,N_2960);
or UO_99 (O_99,N_2992,N_2973);
or UO_100 (O_100,N_2954,N_2998);
nand UO_101 (O_101,N_2981,N_2989);
and UO_102 (O_102,N_2975,N_2972);
or UO_103 (O_103,N_2971,N_2991);
or UO_104 (O_104,N_2966,N_2987);
and UO_105 (O_105,N_2980,N_2986);
or UO_106 (O_106,N_2975,N_2974);
nand UO_107 (O_107,N_2995,N_2970);
or UO_108 (O_108,N_2969,N_2981);
or UO_109 (O_109,N_2979,N_2994);
and UO_110 (O_110,N_2996,N_2978);
nand UO_111 (O_111,N_2989,N_2955);
and UO_112 (O_112,N_2992,N_2980);
or UO_113 (O_113,N_2954,N_2961);
and UO_114 (O_114,N_2982,N_2964);
or UO_115 (O_115,N_2992,N_2960);
and UO_116 (O_116,N_2967,N_2970);
xor UO_117 (O_117,N_2986,N_2967);
nor UO_118 (O_118,N_2985,N_2970);
and UO_119 (O_119,N_2993,N_2999);
or UO_120 (O_120,N_2974,N_2979);
and UO_121 (O_121,N_2984,N_2975);
or UO_122 (O_122,N_2987,N_2975);
and UO_123 (O_123,N_2977,N_2993);
nand UO_124 (O_124,N_2975,N_2982);
nor UO_125 (O_125,N_2968,N_2991);
nor UO_126 (O_126,N_2969,N_2980);
and UO_127 (O_127,N_2972,N_2977);
or UO_128 (O_128,N_2956,N_2973);
nor UO_129 (O_129,N_2994,N_2962);
or UO_130 (O_130,N_2954,N_2986);
nor UO_131 (O_131,N_2964,N_2990);
nand UO_132 (O_132,N_2970,N_2954);
nand UO_133 (O_133,N_2995,N_2977);
and UO_134 (O_134,N_2993,N_2995);
xor UO_135 (O_135,N_2976,N_2970);
or UO_136 (O_136,N_2975,N_2966);
and UO_137 (O_137,N_2976,N_2987);
nor UO_138 (O_138,N_2979,N_2997);
and UO_139 (O_139,N_2986,N_2972);
nand UO_140 (O_140,N_2988,N_2993);
or UO_141 (O_141,N_2970,N_2957);
nor UO_142 (O_142,N_2967,N_2968);
or UO_143 (O_143,N_2952,N_2955);
nand UO_144 (O_144,N_2997,N_2963);
and UO_145 (O_145,N_2998,N_2969);
and UO_146 (O_146,N_2951,N_2962);
and UO_147 (O_147,N_2984,N_2996);
nand UO_148 (O_148,N_2964,N_2991);
nor UO_149 (O_149,N_2970,N_2999);
nor UO_150 (O_150,N_2969,N_2950);
or UO_151 (O_151,N_2962,N_2999);
and UO_152 (O_152,N_2972,N_2955);
and UO_153 (O_153,N_2970,N_2998);
nor UO_154 (O_154,N_2956,N_2958);
nor UO_155 (O_155,N_2993,N_2994);
nand UO_156 (O_156,N_2989,N_2962);
and UO_157 (O_157,N_2975,N_2978);
nand UO_158 (O_158,N_2953,N_2951);
nand UO_159 (O_159,N_2963,N_2952);
nor UO_160 (O_160,N_2991,N_2956);
nor UO_161 (O_161,N_2973,N_2951);
nand UO_162 (O_162,N_2983,N_2992);
nor UO_163 (O_163,N_2989,N_2971);
or UO_164 (O_164,N_2970,N_2968);
nand UO_165 (O_165,N_2953,N_2968);
and UO_166 (O_166,N_2964,N_2993);
and UO_167 (O_167,N_2972,N_2982);
and UO_168 (O_168,N_2967,N_2977);
nand UO_169 (O_169,N_2974,N_2951);
and UO_170 (O_170,N_2985,N_2968);
or UO_171 (O_171,N_2992,N_2964);
or UO_172 (O_172,N_2964,N_2951);
nor UO_173 (O_173,N_2968,N_2980);
or UO_174 (O_174,N_2985,N_2963);
nor UO_175 (O_175,N_2950,N_2988);
and UO_176 (O_176,N_2963,N_2990);
nor UO_177 (O_177,N_2974,N_2980);
nor UO_178 (O_178,N_2963,N_2989);
nand UO_179 (O_179,N_2956,N_2984);
or UO_180 (O_180,N_2994,N_2997);
or UO_181 (O_181,N_2973,N_2955);
nand UO_182 (O_182,N_2965,N_2966);
nor UO_183 (O_183,N_2965,N_2963);
and UO_184 (O_184,N_2972,N_2960);
nor UO_185 (O_185,N_2992,N_2953);
and UO_186 (O_186,N_2959,N_2993);
nand UO_187 (O_187,N_2955,N_2956);
nand UO_188 (O_188,N_2956,N_2970);
or UO_189 (O_189,N_2987,N_2968);
nor UO_190 (O_190,N_2952,N_2958);
and UO_191 (O_191,N_2965,N_2980);
or UO_192 (O_192,N_2994,N_2974);
nand UO_193 (O_193,N_2968,N_2984);
nand UO_194 (O_194,N_2968,N_2955);
nor UO_195 (O_195,N_2957,N_2967);
nand UO_196 (O_196,N_2961,N_2993);
or UO_197 (O_197,N_2967,N_2951);
nor UO_198 (O_198,N_2961,N_2989);
or UO_199 (O_199,N_2989,N_2966);
nand UO_200 (O_200,N_2972,N_2978);
or UO_201 (O_201,N_2964,N_2963);
nand UO_202 (O_202,N_2962,N_2984);
or UO_203 (O_203,N_2997,N_2969);
nand UO_204 (O_204,N_2984,N_2954);
xnor UO_205 (O_205,N_2982,N_2990);
and UO_206 (O_206,N_2997,N_2958);
or UO_207 (O_207,N_2995,N_2981);
nor UO_208 (O_208,N_2994,N_2990);
or UO_209 (O_209,N_2993,N_2950);
or UO_210 (O_210,N_2986,N_2994);
nor UO_211 (O_211,N_2986,N_2968);
nor UO_212 (O_212,N_2980,N_2999);
and UO_213 (O_213,N_2971,N_2980);
or UO_214 (O_214,N_2959,N_2966);
or UO_215 (O_215,N_2957,N_2960);
and UO_216 (O_216,N_2966,N_2979);
and UO_217 (O_217,N_2962,N_2976);
and UO_218 (O_218,N_2964,N_2971);
and UO_219 (O_219,N_2965,N_2962);
or UO_220 (O_220,N_2959,N_2962);
or UO_221 (O_221,N_2982,N_2984);
nand UO_222 (O_222,N_2977,N_2988);
nor UO_223 (O_223,N_2998,N_2972);
or UO_224 (O_224,N_2981,N_2983);
nor UO_225 (O_225,N_2966,N_2983);
and UO_226 (O_226,N_2990,N_2981);
nand UO_227 (O_227,N_2965,N_2959);
nor UO_228 (O_228,N_2990,N_2986);
and UO_229 (O_229,N_2959,N_2950);
nand UO_230 (O_230,N_2990,N_2984);
or UO_231 (O_231,N_2991,N_2990);
nor UO_232 (O_232,N_2953,N_2960);
nor UO_233 (O_233,N_2974,N_2987);
nand UO_234 (O_234,N_2968,N_2992);
nor UO_235 (O_235,N_2974,N_2982);
and UO_236 (O_236,N_2956,N_2976);
nand UO_237 (O_237,N_2977,N_2990);
and UO_238 (O_238,N_2985,N_2975);
nor UO_239 (O_239,N_2993,N_2987);
nand UO_240 (O_240,N_2988,N_2959);
nand UO_241 (O_241,N_2969,N_2966);
nand UO_242 (O_242,N_2959,N_2963);
nor UO_243 (O_243,N_2972,N_2980);
nand UO_244 (O_244,N_2979,N_2978);
and UO_245 (O_245,N_2993,N_2970);
nor UO_246 (O_246,N_2958,N_2957);
nand UO_247 (O_247,N_2989,N_2960);
nand UO_248 (O_248,N_2993,N_2976);
nor UO_249 (O_249,N_2966,N_2952);
nand UO_250 (O_250,N_2969,N_2999);
nor UO_251 (O_251,N_2978,N_2986);
nand UO_252 (O_252,N_2967,N_2999);
or UO_253 (O_253,N_2969,N_2991);
and UO_254 (O_254,N_2994,N_2960);
nor UO_255 (O_255,N_2992,N_2963);
or UO_256 (O_256,N_2996,N_2971);
and UO_257 (O_257,N_2951,N_2987);
or UO_258 (O_258,N_2981,N_2959);
and UO_259 (O_259,N_2952,N_2973);
nor UO_260 (O_260,N_2962,N_2974);
nand UO_261 (O_261,N_2986,N_2966);
or UO_262 (O_262,N_2970,N_2996);
nor UO_263 (O_263,N_2955,N_2951);
and UO_264 (O_264,N_2960,N_2981);
and UO_265 (O_265,N_2967,N_2966);
and UO_266 (O_266,N_2953,N_2955);
nor UO_267 (O_267,N_2991,N_2987);
and UO_268 (O_268,N_2980,N_2996);
or UO_269 (O_269,N_2964,N_2994);
nor UO_270 (O_270,N_2952,N_2972);
nor UO_271 (O_271,N_2960,N_2979);
nand UO_272 (O_272,N_2954,N_2956);
and UO_273 (O_273,N_2982,N_2998);
or UO_274 (O_274,N_2993,N_2979);
or UO_275 (O_275,N_2953,N_2972);
and UO_276 (O_276,N_2950,N_2977);
nor UO_277 (O_277,N_2962,N_2966);
nand UO_278 (O_278,N_2986,N_2963);
or UO_279 (O_279,N_2957,N_2982);
nand UO_280 (O_280,N_2990,N_2965);
nand UO_281 (O_281,N_2962,N_2950);
or UO_282 (O_282,N_2967,N_2969);
nor UO_283 (O_283,N_2999,N_2951);
and UO_284 (O_284,N_2954,N_2960);
nand UO_285 (O_285,N_2965,N_2951);
and UO_286 (O_286,N_2994,N_2989);
or UO_287 (O_287,N_2997,N_2985);
nand UO_288 (O_288,N_2977,N_2986);
or UO_289 (O_289,N_2991,N_2957);
nand UO_290 (O_290,N_2991,N_2965);
xor UO_291 (O_291,N_2977,N_2951);
nand UO_292 (O_292,N_2985,N_2990);
nor UO_293 (O_293,N_2953,N_2977);
nand UO_294 (O_294,N_2978,N_2989);
and UO_295 (O_295,N_2957,N_2999);
and UO_296 (O_296,N_2964,N_2980);
and UO_297 (O_297,N_2975,N_2977);
or UO_298 (O_298,N_2989,N_2968);
nand UO_299 (O_299,N_2952,N_2978);
and UO_300 (O_300,N_2953,N_2995);
and UO_301 (O_301,N_2988,N_2981);
xor UO_302 (O_302,N_2995,N_2952);
nand UO_303 (O_303,N_2994,N_2967);
nand UO_304 (O_304,N_2992,N_2985);
nor UO_305 (O_305,N_2996,N_2986);
nand UO_306 (O_306,N_2981,N_2987);
nand UO_307 (O_307,N_2989,N_2982);
and UO_308 (O_308,N_2994,N_2992);
or UO_309 (O_309,N_2950,N_2967);
nor UO_310 (O_310,N_2964,N_2999);
nor UO_311 (O_311,N_2967,N_2997);
and UO_312 (O_312,N_2975,N_2951);
or UO_313 (O_313,N_2969,N_2983);
nor UO_314 (O_314,N_2954,N_2988);
or UO_315 (O_315,N_2958,N_2955);
nand UO_316 (O_316,N_2972,N_2954);
or UO_317 (O_317,N_2995,N_2969);
xnor UO_318 (O_318,N_2961,N_2955);
and UO_319 (O_319,N_2969,N_2962);
and UO_320 (O_320,N_2969,N_2954);
or UO_321 (O_321,N_2991,N_2952);
nor UO_322 (O_322,N_2978,N_2964);
or UO_323 (O_323,N_2956,N_2959);
nor UO_324 (O_324,N_2959,N_2969);
nand UO_325 (O_325,N_2969,N_2970);
or UO_326 (O_326,N_2997,N_2996);
nand UO_327 (O_327,N_2982,N_2978);
nand UO_328 (O_328,N_2999,N_2992);
nand UO_329 (O_329,N_2999,N_2987);
nor UO_330 (O_330,N_2997,N_2984);
xnor UO_331 (O_331,N_2957,N_2969);
or UO_332 (O_332,N_2958,N_2999);
nand UO_333 (O_333,N_2974,N_2986);
nand UO_334 (O_334,N_2955,N_2982);
or UO_335 (O_335,N_2985,N_2972);
nand UO_336 (O_336,N_2984,N_2992);
and UO_337 (O_337,N_2978,N_2950);
nand UO_338 (O_338,N_2991,N_2994);
nand UO_339 (O_339,N_2978,N_2959);
nor UO_340 (O_340,N_2992,N_2979);
or UO_341 (O_341,N_2990,N_2971);
and UO_342 (O_342,N_2980,N_2951);
nor UO_343 (O_343,N_2964,N_2972);
nor UO_344 (O_344,N_2972,N_2989);
nand UO_345 (O_345,N_2997,N_2975);
xnor UO_346 (O_346,N_2967,N_2952);
or UO_347 (O_347,N_2959,N_2951);
or UO_348 (O_348,N_2995,N_2988);
nor UO_349 (O_349,N_2973,N_2998);
nor UO_350 (O_350,N_2986,N_2984);
and UO_351 (O_351,N_2996,N_2992);
and UO_352 (O_352,N_2975,N_2989);
or UO_353 (O_353,N_2969,N_2979);
nand UO_354 (O_354,N_2983,N_2989);
nand UO_355 (O_355,N_2958,N_2982);
and UO_356 (O_356,N_2979,N_2954);
and UO_357 (O_357,N_2956,N_2972);
or UO_358 (O_358,N_2952,N_2976);
nand UO_359 (O_359,N_2972,N_2988);
or UO_360 (O_360,N_2974,N_2995);
nor UO_361 (O_361,N_2966,N_2980);
or UO_362 (O_362,N_2951,N_2963);
nor UO_363 (O_363,N_2970,N_2980);
and UO_364 (O_364,N_2978,N_2976);
and UO_365 (O_365,N_2990,N_2972);
or UO_366 (O_366,N_2990,N_2989);
nand UO_367 (O_367,N_2965,N_2996);
nor UO_368 (O_368,N_2952,N_2977);
or UO_369 (O_369,N_2955,N_2993);
or UO_370 (O_370,N_2954,N_2950);
or UO_371 (O_371,N_2993,N_2992);
or UO_372 (O_372,N_2977,N_2974);
or UO_373 (O_373,N_2978,N_2994);
or UO_374 (O_374,N_2979,N_2951);
nand UO_375 (O_375,N_2968,N_2951);
and UO_376 (O_376,N_2985,N_2962);
nor UO_377 (O_377,N_2994,N_2973);
nand UO_378 (O_378,N_2957,N_2959);
or UO_379 (O_379,N_2985,N_2967);
or UO_380 (O_380,N_2965,N_2975);
nor UO_381 (O_381,N_2984,N_2951);
nor UO_382 (O_382,N_2951,N_2994);
or UO_383 (O_383,N_2963,N_2955);
nor UO_384 (O_384,N_2964,N_2998);
or UO_385 (O_385,N_2988,N_2979);
or UO_386 (O_386,N_2974,N_2953);
nor UO_387 (O_387,N_2957,N_2979);
or UO_388 (O_388,N_2952,N_2962);
nor UO_389 (O_389,N_2993,N_2983);
and UO_390 (O_390,N_2982,N_2971);
and UO_391 (O_391,N_2989,N_2986);
nand UO_392 (O_392,N_2983,N_2956);
xnor UO_393 (O_393,N_2992,N_2998);
or UO_394 (O_394,N_2969,N_2951);
and UO_395 (O_395,N_2991,N_2958);
and UO_396 (O_396,N_2992,N_2970);
or UO_397 (O_397,N_2990,N_2966);
or UO_398 (O_398,N_2968,N_2977);
and UO_399 (O_399,N_2959,N_2970);
xor UO_400 (O_400,N_2980,N_2978);
nand UO_401 (O_401,N_2975,N_2962);
nand UO_402 (O_402,N_2965,N_2961);
nor UO_403 (O_403,N_2962,N_2991);
and UO_404 (O_404,N_2964,N_2952);
or UO_405 (O_405,N_2979,N_2999);
xnor UO_406 (O_406,N_2993,N_2956);
nand UO_407 (O_407,N_2977,N_2963);
nor UO_408 (O_408,N_2965,N_2955);
nand UO_409 (O_409,N_2968,N_2969);
or UO_410 (O_410,N_2954,N_2978);
and UO_411 (O_411,N_2984,N_2972);
or UO_412 (O_412,N_2980,N_2993);
or UO_413 (O_413,N_2979,N_2958);
xor UO_414 (O_414,N_2953,N_2980);
nor UO_415 (O_415,N_2986,N_2975);
or UO_416 (O_416,N_2999,N_2982);
nand UO_417 (O_417,N_2962,N_2986);
and UO_418 (O_418,N_2999,N_2955);
nand UO_419 (O_419,N_2990,N_2959);
nand UO_420 (O_420,N_2996,N_2973);
and UO_421 (O_421,N_2983,N_2991);
and UO_422 (O_422,N_2952,N_2992);
nor UO_423 (O_423,N_2957,N_2964);
nand UO_424 (O_424,N_2952,N_2994);
and UO_425 (O_425,N_2974,N_2976);
nor UO_426 (O_426,N_2961,N_2979);
nand UO_427 (O_427,N_2983,N_2972);
nand UO_428 (O_428,N_2998,N_2963);
xor UO_429 (O_429,N_2959,N_2989);
and UO_430 (O_430,N_2968,N_2978);
nand UO_431 (O_431,N_2990,N_2999);
nand UO_432 (O_432,N_2986,N_2961);
or UO_433 (O_433,N_2976,N_2983);
nand UO_434 (O_434,N_2967,N_2998);
or UO_435 (O_435,N_2990,N_2970);
nand UO_436 (O_436,N_2969,N_2978);
nor UO_437 (O_437,N_2965,N_2960);
or UO_438 (O_438,N_2968,N_2997);
nand UO_439 (O_439,N_2963,N_2973);
nand UO_440 (O_440,N_2984,N_2957);
and UO_441 (O_441,N_2981,N_2963);
nand UO_442 (O_442,N_2995,N_2971);
or UO_443 (O_443,N_2995,N_2987);
or UO_444 (O_444,N_2966,N_2956);
or UO_445 (O_445,N_2995,N_2956);
and UO_446 (O_446,N_2989,N_2984);
or UO_447 (O_447,N_2987,N_2969);
or UO_448 (O_448,N_2961,N_2987);
and UO_449 (O_449,N_2997,N_2988);
nand UO_450 (O_450,N_2968,N_2975);
or UO_451 (O_451,N_2961,N_2964);
and UO_452 (O_452,N_2964,N_2973);
nor UO_453 (O_453,N_2973,N_2999);
nor UO_454 (O_454,N_2961,N_2988);
and UO_455 (O_455,N_2976,N_2989);
nor UO_456 (O_456,N_2982,N_2966);
or UO_457 (O_457,N_2950,N_2985);
nor UO_458 (O_458,N_2956,N_2981);
nand UO_459 (O_459,N_2965,N_2976);
nor UO_460 (O_460,N_2951,N_2966);
nand UO_461 (O_461,N_2970,N_2978);
and UO_462 (O_462,N_2966,N_2958);
or UO_463 (O_463,N_2962,N_2982);
or UO_464 (O_464,N_2965,N_2979);
or UO_465 (O_465,N_2963,N_2954);
nor UO_466 (O_466,N_2977,N_2978);
or UO_467 (O_467,N_2964,N_2976);
and UO_468 (O_468,N_2984,N_2974);
nand UO_469 (O_469,N_2995,N_2978);
nor UO_470 (O_470,N_2987,N_2952);
or UO_471 (O_471,N_2971,N_2978);
and UO_472 (O_472,N_2965,N_2994);
nor UO_473 (O_473,N_2953,N_2976);
and UO_474 (O_474,N_2983,N_2977);
nor UO_475 (O_475,N_2960,N_2962);
nor UO_476 (O_476,N_2980,N_2954);
or UO_477 (O_477,N_2976,N_2973);
nor UO_478 (O_478,N_2988,N_2978);
xnor UO_479 (O_479,N_2985,N_2977);
and UO_480 (O_480,N_2984,N_2985);
nor UO_481 (O_481,N_2986,N_2976);
or UO_482 (O_482,N_2978,N_2993);
and UO_483 (O_483,N_2978,N_2955);
nor UO_484 (O_484,N_2996,N_2974);
nand UO_485 (O_485,N_2976,N_2963);
nor UO_486 (O_486,N_2986,N_2992);
nand UO_487 (O_487,N_2985,N_2982);
or UO_488 (O_488,N_2978,N_2981);
or UO_489 (O_489,N_2985,N_2959);
nor UO_490 (O_490,N_2953,N_2983);
nor UO_491 (O_491,N_2984,N_2953);
xnor UO_492 (O_492,N_2956,N_2965);
and UO_493 (O_493,N_2971,N_2984);
nor UO_494 (O_494,N_2961,N_2994);
nand UO_495 (O_495,N_2971,N_2998);
and UO_496 (O_496,N_2991,N_2975);
or UO_497 (O_497,N_2999,N_2981);
and UO_498 (O_498,N_2961,N_2966);
and UO_499 (O_499,N_2952,N_2971);
endmodule