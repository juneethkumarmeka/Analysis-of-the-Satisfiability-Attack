module basic_1000_10000_1500_2_levels_1xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5002,N_5004,N_5005,N_5007,N_5008,N_5009,N_5011,N_5012,N_5015,N_5018,N_5019,N_5020,N_5021,N_5022,N_5027,N_5028,N_5029,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5039,N_5040,N_5042,N_5043,N_5044,N_5045,N_5046,N_5048,N_5049,N_5050,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5061,N_5065,N_5066,N_5068,N_5069,N_5071,N_5072,N_5074,N_5075,N_5076,N_5077,N_5080,N_5081,N_5083,N_5084,N_5087,N_5088,N_5090,N_5091,N_5092,N_5093,N_5095,N_5098,N_5101,N_5102,N_5105,N_5107,N_5110,N_5111,N_5112,N_5113,N_5114,N_5117,N_5118,N_5122,N_5123,N_5125,N_5126,N_5127,N_5131,N_5132,N_5133,N_5134,N_5136,N_5137,N_5138,N_5139,N_5140,N_5143,N_5145,N_5147,N_5148,N_5149,N_5151,N_5152,N_5153,N_5155,N_5156,N_5157,N_5159,N_5162,N_5164,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5178,N_5179,N_5180,N_5181,N_5182,N_5184,N_5186,N_5188,N_5190,N_5192,N_5193,N_5194,N_5195,N_5196,N_5198,N_5204,N_5208,N_5209,N_5210,N_5211,N_5212,N_5214,N_5215,N_5216,N_5219,N_5220,N_5221,N_5222,N_5224,N_5227,N_5228,N_5229,N_5230,N_5231,N_5234,N_5235,N_5237,N_5238,N_5240,N_5241,N_5242,N_5245,N_5246,N_5247,N_5248,N_5251,N_5252,N_5256,N_5258,N_5260,N_5261,N_5262,N_5263,N_5264,N_5266,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5280,N_5281,N_5285,N_5286,N_5287,N_5290,N_5291,N_5293,N_5294,N_5296,N_5297,N_5299,N_5303,N_5305,N_5306,N_5309,N_5310,N_5311,N_5313,N_5314,N_5316,N_5317,N_5319,N_5320,N_5321,N_5322,N_5323,N_5325,N_5326,N_5331,N_5332,N_5334,N_5335,N_5337,N_5338,N_5339,N_5341,N_5345,N_5346,N_5347,N_5348,N_5351,N_5352,N_5353,N_5354,N_5356,N_5357,N_5358,N_5361,N_5362,N_5363,N_5364,N_5365,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5385,N_5386,N_5387,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5400,N_5401,N_5404,N_5409,N_5410,N_5412,N_5413,N_5415,N_5418,N_5419,N_5420,N_5422,N_5423,N_5424,N_5425,N_5427,N_5428,N_5429,N_5430,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5441,N_5442,N_5444,N_5446,N_5451,N_5455,N_5456,N_5458,N_5460,N_5461,N_5462,N_5465,N_5466,N_5469,N_5470,N_5472,N_5473,N_5474,N_5475,N_5477,N_5478,N_5482,N_5483,N_5487,N_5488,N_5490,N_5491,N_5495,N_5496,N_5497,N_5498,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5516,N_5517,N_5518,N_5519,N_5520,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5531,N_5532,N_5534,N_5535,N_5536,N_5540,N_5541,N_5542,N_5543,N_5545,N_5547,N_5549,N_5551,N_5552,N_5555,N_5556,N_5560,N_5561,N_5564,N_5565,N_5567,N_5568,N_5569,N_5573,N_5574,N_5575,N_5576,N_5578,N_5579,N_5581,N_5582,N_5583,N_5588,N_5589,N_5590,N_5592,N_5593,N_5594,N_5596,N_5598,N_5600,N_5602,N_5603,N_5605,N_5606,N_5607,N_5608,N_5611,N_5615,N_5616,N_5617,N_5619,N_5622,N_5624,N_5628,N_5629,N_5630,N_5631,N_5632,N_5635,N_5638,N_5640,N_5641,N_5643,N_5645,N_5646,N_5650,N_5653,N_5654,N_5655,N_5657,N_5660,N_5662,N_5663,N_5664,N_5665,N_5666,N_5668,N_5670,N_5671,N_5672,N_5674,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5684,N_5686,N_5687,N_5688,N_5689,N_5691,N_5694,N_5695,N_5696,N_5697,N_5699,N_5704,N_5706,N_5707,N_5709,N_5711,N_5713,N_5717,N_5720,N_5721,N_5724,N_5727,N_5729,N_5730,N_5732,N_5733,N_5735,N_5736,N_5742,N_5743,N_5744,N_5746,N_5748,N_5749,N_5750,N_5753,N_5756,N_5757,N_5759,N_5761,N_5763,N_5764,N_5765,N_5766,N_5768,N_5769,N_5770,N_5771,N_5773,N_5774,N_5776,N_5777,N_5778,N_5780,N_5781,N_5782,N_5783,N_5785,N_5787,N_5788,N_5789,N_5793,N_5797,N_5798,N_5800,N_5803,N_5805,N_5806,N_5807,N_5811,N_5813,N_5814,N_5817,N_5818,N_5819,N_5822,N_5823,N_5825,N_5826,N_5829,N_5831,N_5834,N_5835,N_5836,N_5837,N_5839,N_5840,N_5841,N_5843,N_5844,N_5845,N_5849,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5860,N_5863,N_5864,N_5867,N_5871,N_5873,N_5877,N_5879,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5888,N_5891,N_5892,N_5894,N_5897,N_5900,N_5902,N_5908,N_5911,N_5912,N_5914,N_5916,N_5917,N_5920,N_5921,N_5922,N_5924,N_5926,N_5930,N_5931,N_5933,N_5934,N_5936,N_5937,N_5938,N_5940,N_5942,N_5943,N_5945,N_5946,N_5947,N_5951,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5961,N_5962,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5976,N_5980,N_5981,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5993,N_5994,N_5996,N_5997,N_5998,N_6000,N_6001,N_6002,N_6004,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6015,N_6016,N_6017,N_6018,N_6020,N_6021,N_6022,N_6025,N_6026,N_6027,N_6028,N_6029,N_6031,N_6033,N_6034,N_6037,N_6040,N_6041,N_6043,N_6044,N_6045,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6056,N_6058,N_6059,N_6060,N_6065,N_6067,N_6069,N_6072,N_6073,N_6074,N_6077,N_6079,N_6080,N_6081,N_6082,N_6083,N_6086,N_6089,N_6090,N_6091,N_6092,N_6095,N_6098,N_6099,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6108,N_6109,N_6111,N_6113,N_6115,N_6117,N_6120,N_6122,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6133,N_6134,N_6136,N_6139,N_6143,N_6145,N_6146,N_6148,N_6151,N_6152,N_6154,N_6155,N_6156,N_6157,N_6158,N_6160,N_6161,N_6162,N_6163,N_6164,N_6168,N_6170,N_6171,N_6174,N_6175,N_6177,N_6178,N_6181,N_6182,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6197,N_6198,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6210,N_6212,N_6213,N_6214,N_6215,N_6217,N_6218,N_6220,N_6225,N_6227,N_6229,N_6234,N_6236,N_6238,N_6239,N_6241,N_6242,N_6243,N_6244,N_6248,N_6249,N_6250,N_6251,N_6254,N_6255,N_6256,N_6259,N_6261,N_6262,N_6263,N_6264,N_6265,N_6267,N_6269,N_6270,N_6272,N_6273,N_6276,N_6278,N_6281,N_6282,N_6284,N_6285,N_6288,N_6289,N_6290,N_6293,N_6295,N_6296,N_6297,N_6298,N_6299,N_6302,N_6303,N_6304,N_6307,N_6308,N_6310,N_6311,N_6312,N_6313,N_6319,N_6321,N_6322,N_6323,N_6324,N_6326,N_6327,N_6330,N_6331,N_6332,N_6333,N_6335,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6345,N_6346,N_6347,N_6350,N_6351,N_6353,N_6354,N_6356,N_6358,N_6359,N_6360,N_6361,N_6362,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6372,N_6373,N_6374,N_6376,N_6378,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6388,N_6389,N_6391,N_6392,N_6393,N_6394,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6404,N_6405,N_6406,N_6408,N_6410,N_6412,N_6413,N_6414,N_6415,N_6417,N_6418,N_6420,N_6421,N_6422,N_6423,N_6427,N_6428,N_6429,N_6430,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6440,N_6441,N_6442,N_6444,N_6446,N_6447,N_6448,N_6449,N_6450,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6464,N_6465,N_6466,N_6468,N_6469,N_6471,N_6473,N_6474,N_6475,N_6480,N_6482,N_6483,N_6484,N_6485,N_6487,N_6492,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6507,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6518,N_6520,N_6522,N_6523,N_6524,N_6525,N_6526,N_6529,N_6530,N_6533,N_6534,N_6536,N_6537,N_6539,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6549,N_6550,N_6552,N_6553,N_6556,N_6557,N_6558,N_6559,N_6560,N_6563,N_6564,N_6566,N_6569,N_6570,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6579,N_6580,N_6581,N_6582,N_6583,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6596,N_6597,N_6598,N_6599,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6612,N_6613,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6628,N_6630,N_6632,N_6634,N_6641,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6653,N_6655,N_6657,N_6658,N_6662,N_6663,N_6664,N_6667,N_6668,N_6669,N_6670,N_6672,N_6673,N_6676,N_6680,N_6683,N_6684,N_6688,N_6689,N_6690,N_6693,N_6696,N_6697,N_6698,N_6701,N_6702,N_6703,N_6707,N_6709,N_6711,N_6715,N_6718,N_6719,N_6721,N_6722,N_6723,N_6725,N_6727,N_6728,N_6729,N_6731,N_6734,N_6736,N_6737,N_6738,N_6741,N_6743,N_6745,N_6746,N_6747,N_6748,N_6749,N_6754,N_6757,N_6761,N_6762,N_6763,N_6764,N_6765,N_6767,N_6770,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6780,N_6782,N_6786,N_6788,N_6791,N_6793,N_6796,N_6797,N_6802,N_6805,N_6806,N_6807,N_6810,N_6811,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6824,N_6825,N_6827,N_6829,N_6830,N_6831,N_6832,N_6833,N_6835,N_6839,N_6840,N_6842,N_6843,N_6844,N_6845,N_6848,N_6852,N_6853,N_6854,N_6856,N_6857,N_6858,N_6860,N_6861,N_6862,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6873,N_6875,N_6876,N_6877,N_6881,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6897,N_6898,N_6900,N_6901,N_6904,N_6906,N_6907,N_6908,N_6911,N_6912,N_6916,N_6919,N_6921,N_6922,N_6923,N_6924,N_6926,N_6927,N_6929,N_6930,N_6933,N_6934,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6945,N_6947,N_6948,N_6949,N_6953,N_6955,N_6957,N_6959,N_6961,N_6962,N_6965,N_6966,N_6967,N_6968,N_6969,N_6971,N_6972,N_6973,N_6975,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6987,N_6988,N_6990,N_6991,N_6993,N_6994,N_6999,N_7003,N_7004,N_7008,N_7010,N_7011,N_7012,N_7013,N_7015,N_7020,N_7021,N_7023,N_7025,N_7026,N_7027,N_7029,N_7031,N_7032,N_7034,N_7035,N_7036,N_7038,N_7039,N_7041,N_7045,N_7048,N_7049,N_7050,N_7051,N_7053,N_7054,N_7055,N_7056,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7066,N_7072,N_7073,N_7074,N_7077,N_7078,N_7079,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7091,N_7093,N_7094,N_7096,N_7097,N_7099,N_7100,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7125,N_7126,N_7128,N_7130,N_7131,N_7132,N_7134,N_7136,N_7138,N_7140,N_7141,N_7142,N_7143,N_7147,N_7148,N_7149,N_7151,N_7153,N_7154,N_7155,N_7156,N_7157,N_7159,N_7160,N_7161,N_7162,N_7163,N_7166,N_7168,N_7170,N_7172,N_7174,N_7175,N_7176,N_7182,N_7183,N_7186,N_7188,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7198,N_7199,N_7201,N_7202,N_7203,N_7204,N_7205,N_7208,N_7209,N_7210,N_7211,N_7213,N_7216,N_7217,N_7218,N_7220,N_7221,N_7223,N_7224,N_7230,N_7231,N_7234,N_7235,N_7236,N_7237,N_7240,N_7241,N_7245,N_7246,N_7248,N_7249,N_7253,N_7254,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7268,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7282,N_7283,N_7284,N_7286,N_7288,N_7289,N_7294,N_7295,N_7296,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7310,N_7311,N_7312,N_7318,N_7319,N_7322,N_7323,N_7324,N_7325,N_7328,N_7329,N_7330,N_7331,N_7334,N_7338,N_7340,N_7341,N_7343,N_7345,N_7347,N_7348,N_7349,N_7350,N_7351,N_7354,N_7356,N_7358,N_7359,N_7361,N_7362,N_7363,N_7366,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7376,N_7378,N_7381,N_7384,N_7388,N_7389,N_7390,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7404,N_7405,N_7406,N_7408,N_7411,N_7412,N_7413,N_7415,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7427,N_7428,N_7431,N_7432,N_7433,N_7435,N_7436,N_7440,N_7442,N_7444,N_7445,N_7446,N_7451,N_7452,N_7453,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7462,N_7463,N_7469,N_7471,N_7473,N_7474,N_7475,N_7476,N_7479,N_7480,N_7484,N_7485,N_7486,N_7488,N_7491,N_7492,N_7493,N_7494,N_7496,N_7497,N_7499,N_7500,N_7501,N_7502,N_7504,N_7507,N_7509,N_7510,N_7512,N_7515,N_7516,N_7518,N_7520,N_7523,N_7524,N_7525,N_7526,N_7528,N_7531,N_7534,N_7535,N_7537,N_7542,N_7543,N_7545,N_7547,N_7548,N_7553,N_7556,N_7558,N_7560,N_7561,N_7563,N_7565,N_7566,N_7567,N_7570,N_7571,N_7572,N_7573,N_7574,N_7576,N_7578,N_7581,N_7583,N_7584,N_7586,N_7587,N_7588,N_7590,N_7592,N_7594,N_7596,N_7597,N_7598,N_7599,N_7604,N_7605,N_7607,N_7608,N_7610,N_7611,N_7612,N_7614,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7625,N_7626,N_7627,N_7629,N_7630,N_7633,N_7634,N_7637,N_7638,N_7639,N_7640,N_7641,N_7643,N_7644,N_7645,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7657,N_7658,N_7659,N_7661,N_7666,N_7668,N_7670,N_7673,N_7674,N_7675,N_7677,N_7681,N_7684,N_7685,N_7686,N_7689,N_7690,N_7691,N_7692,N_7694,N_7696,N_7697,N_7698,N_7699,N_7701,N_7703,N_7705,N_7706,N_7708,N_7712,N_7713,N_7714,N_7715,N_7717,N_7719,N_7720,N_7721,N_7722,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7734,N_7735,N_7737,N_7738,N_7740,N_7744,N_7745,N_7746,N_7748,N_7750,N_7753,N_7756,N_7757,N_7758,N_7760,N_7761,N_7764,N_7765,N_7766,N_7767,N_7768,N_7771,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7786,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7798,N_7799,N_7800,N_7802,N_7804,N_7805,N_7809,N_7813,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7824,N_7825,N_7827,N_7828,N_7829,N_7831,N_7833,N_7834,N_7837,N_7838,N_7839,N_7841,N_7842,N_7843,N_7844,N_7845,N_7847,N_7849,N_7852,N_7854,N_7856,N_7857,N_7858,N_7863,N_7866,N_7868,N_7869,N_7871,N_7872,N_7873,N_7874,N_7875,N_7877,N_7878,N_7882,N_7886,N_7896,N_7897,N_7898,N_7899,N_7901,N_7902,N_7903,N_7906,N_7908,N_7911,N_7914,N_7917,N_7920,N_7922,N_7923,N_7924,N_7925,N_7926,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7936,N_7938,N_7939,N_7940,N_7944,N_7945,N_7947,N_7948,N_7952,N_7954,N_7955,N_7956,N_7957,N_7959,N_7960,N_7961,N_7962,N_7964,N_7966,N_7968,N_7970,N_7971,N_7972,N_7974,N_7977,N_7978,N_7979,N_7980,N_7983,N_7985,N_7987,N_7988,N_7989,N_7990,N_7991,N_7994,N_7995,N_7996,N_7997,N_8000,N_8003,N_8005,N_8007,N_8011,N_8014,N_8015,N_8016,N_8017,N_8019,N_8022,N_8023,N_8024,N_8026,N_8027,N_8028,N_8029,N_8030,N_8038,N_8039,N_8040,N_8041,N_8043,N_8044,N_8045,N_8046,N_8047,N_8049,N_8050,N_8051,N_8053,N_8056,N_8057,N_8058,N_8060,N_8061,N_8065,N_8066,N_8067,N_8068,N_8069,N_8072,N_8073,N_8074,N_8075,N_8076,N_8078,N_8080,N_8083,N_8086,N_8087,N_8088,N_8089,N_8090,N_8092,N_8093,N_8095,N_8099,N_8100,N_8103,N_8104,N_8106,N_8108,N_8112,N_8114,N_8115,N_8117,N_8118,N_8119,N_8120,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8138,N_8139,N_8140,N_8142,N_8143,N_8146,N_8149,N_8151,N_8152,N_8154,N_8155,N_8156,N_8157,N_8158,N_8161,N_8162,N_8164,N_8165,N_8168,N_8170,N_8172,N_8175,N_8176,N_8179,N_8180,N_8181,N_8182,N_8184,N_8187,N_8188,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8200,N_8203,N_8205,N_8206,N_8209,N_8210,N_8211,N_8213,N_8214,N_8215,N_8216,N_8217,N_8219,N_8220,N_8222,N_8223,N_8225,N_8226,N_8228,N_8229,N_8232,N_8233,N_8236,N_8240,N_8241,N_8246,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8256,N_8258,N_8260,N_8261,N_8262,N_8263,N_8264,N_8266,N_8267,N_8269,N_8270,N_8271,N_8272,N_8277,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8291,N_8292,N_8294,N_8296,N_8298,N_8300,N_8301,N_8304,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8316,N_8317,N_8319,N_8320,N_8323,N_8324,N_8325,N_8327,N_8328,N_8331,N_8332,N_8334,N_8335,N_8336,N_8337,N_8338,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8349,N_8350,N_8351,N_8352,N_8355,N_8357,N_8358,N_8359,N_8360,N_8362,N_8363,N_8364,N_8365,N_8368,N_8370,N_8376,N_8377,N_8378,N_8382,N_8384,N_8385,N_8386,N_8387,N_8391,N_8392,N_8396,N_8398,N_8400,N_8401,N_8403,N_8404,N_8405,N_8408,N_8410,N_8411,N_8412,N_8413,N_8415,N_8416,N_8417,N_8419,N_8424,N_8425,N_8427,N_8428,N_8429,N_8430,N_8431,N_8433,N_8435,N_8436,N_8437,N_8438,N_8440,N_8441,N_8442,N_8447,N_8448,N_8449,N_8451,N_8453,N_8454,N_8457,N_8458,N_8459,N_8461,N_8462,N_8463,N_8467,N_8469,N_8470,N_8471,N_8473,N_8474,N_8475,N_8476,N_8479,N_8480,N_8482,N_8483,N_8486,N_8487,N_8488,N_8489,N_8490,N_8493,N_8496,N_8499,N_8500,N_8501,N_8502,N_8504,N_8506,N_8507,N_8510,N_8512,N_8514,N_8515,N_8517,N_8521,N_8522,N_8523,N_8524,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8538,N_8539,N_8541,N_8543,N_8544,N_8546,N_8547,N_8550,N_8551,N_8553,N_8557,N_8558,N_8559,N_8560,N_8564,N_8565,N_8566,N_8568,N_8569,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8580,N_8581,N_8582,N_8585,N_8589,N_8592,N_8593,N_8594,N_8595,N_8598,N_8599,N_8602,N_8603,N_8604,N_8606,N_8611,N_8613,N_8616,N_8618,N_8619,N_8620,N_8621,N_8622,N_8625,N_8627,N_8630,N_8631,N_8632,N_8634,N_8637,N_8639,N_8640,N_8641,N_8644,N_8645,N_8646,N_8648,N_8651,N_8652,N_8653,N_8655,N_8657,N_8658,N_8659,N_8663,N_8664,N_8665,N_8666,N_8667,N_8669,N_8670,N_8672,N_8673,N_8674,N_8675,N_8677,N_8680,N_8682,N_8683,N_8684,N_8686,N_8687,N_8689,N_8690,N_8691,N_8692,N_8693,N_8695,N_8698,N_8699,N_8701,N_8702,N_8704,N_8705,N_8706,N_8707,N_8709,N_8710,N_8712,N_8714,N_8715,N_8718,N_8720,N_8722,N_8723,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8735,N_8737,N_8739,N_8740,N_8742,N_8744,N_8746,N_8747,N_8750,N_8751,N_8752,N_8753,N_8754,N_8757,N_8758,N_8759,N_8761,N_8764,N_8765,N_8766,N_8768,N_8770,N_8773,N_8774,N_8776,N_8777,N_8783,N_8784,N_8786,N_8787,N_8788,N_8789,N_8792,N_8793,N_8794,N_8795,N_8797,N_8799,N_8801,N_8802,N_8804,N_8805,N_8806,N_8807,N_8808,N_8811,N_8812,N_8813,N_8817,N_8819,N_8820,N_8821,N_8822,N_8824,N_8825,N_8826,N_8828,N_8831,N_8833,N_8836,N_8837,N_8838,N_8839,N_8840,N_8842,N_8843,N_8844,N_8845,N_8847,N_8851,N_8852,N_8855,N_8856,N_8858,N_8860,N_8862,N_8864,N_8865,N_8869,N_8871,N_8872,N_8874,N_8875,N_8877,N_8879,N_8880,N_8881,N_8882,N_8886,N_8890,N_8891,N_8892,N_8895,N_8897,N_8898,N_8899,N_8900,N_8901,N_8903,N_8904,N_8905,N_8907,N_8908,N_8909,N_8911,N_8912,N_8916,N_8917,N_8919,N_8920,N_8921,N_8922,N_8923,N_8925,N_8926,N_8928,N_8930,N_8938,N_8939,N_8941,N_8943,N_8945,N_8946,N_8949,N_8951,N_8952,N_8953,N_8958,N_8959,N_8961,N_8962,N_8964,N_8965,N_8966,N_8967,N_8969,N_8970,N_8974,N_8975,N_8979,N_8985,N_8987,N_8988,N_8990,N_8991,N_8993,N_8994,N_8995,N_8998,N_8999,N_9000,N_9001,N_9003,N_9005,N_9006,N_9011,N_9013,N_9016,N_9017,N_9018,N_9019,N_9020,N_9022,N_9024,N_9025,N_9026,N_9028,N_9031,N_9033,N_9034,N_9035,N_9037,N_9038,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9050,N_9051,N_9053,N_9056,N_9057,N_9058,N_9059,N_9060,N_9062,N_9064,N_9067,N_9068,N_9070,N_9071,N_9074,N_9076,N_9078,N_9079,N_9080,N_9081,N_9083,N_9084,N_9085,N_9086,N_9089,N_9090,N_9091,N_9092,N_9093,N_9096,N_9098,N_9099,N_9102,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9112,N_9113,N_9114,N_9118,N_9120,N_9121,N_9122,N_9125,N_9126,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9138,N_9139,N_9141,N_9142,N_9143,N_9144,N_9145,N_9147,N_9148,N_9150,N_9152,N_9154,N_9155,N_9156,N_9157,N_9159,N_9160,N_9161,N_9162,N_9164,N_9165,N_9166,N_9167,N_9175,N_9176,N_9177,N_9179,N_9184,N_9185,N_9191,N_9192,N_9195,N_9198,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9211,N_9213,N_9214,N_9215,N_9216,N_9219,N_9221,N_9222,N_9223,N_9224,N_9225,N_9227,N_9229,N_9231,N_9236,N_9237,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9248,N_9249,N_9250,N_9251,N_9253,N_9254,N_9255,N_9258,N_9259,N_9263,N_9265,N_9268,N_9269,N_9270,N_9273,N_9274,N_9275,N_9276,N_9278,N_9281,N_9282,N_9283,N_9285,N_9286,N_9289,N_9290,N_9293,N_9295,N_9297,N_9300,N_9301,N_9303,N_9304,N_9307,N_9308,N_9309,N_9310,N_9312,N_9314,N_9317,N_9321,N_9324,N_9325,N_9326,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9337,N_9339,N_9340,N_9341,N_9345,N_9346,N_9349,N_9350,N_9353,N_9354,N_9355,N_9357,N_9358,N_9359,N_9360,N_9364,N_9365,N_9366,N_9370,N_9371,N_9372,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9383,N_9384,N_9385,N_9390,N_9392,N_9393,N_9397,N_9398,N_9399,N_9400,N_9401,N_9406,N_9408,N_9409,N_9411,N_9413,N_9415,N_9416,N_9417,N_9420,N_9421,N_9425,N_9427,N_9432,N_9433,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9442,N_9444,N_9445,N_9447,N_9449,N_9450,N_9453,N_9454,N_9456,N_9457,N_9459,N_9460,N_9463,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9474,N_9476,N_9480,N_9481,N_9483,N_9484,N_9485,N_9486,N_9488,N_9490,N_9493,N_9494,N_9498,N_9500,N_9501,N_9505,N_9507,N_9508,N_9512,N_9515,N_9516,N_9520,N_9523,N_9526,N_9527,N_9531,N_9533,N_9535,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9547,N_9548,N_9549,N_9550,N_9551,N_9553,N_9555,N_9556,N_9557,N_9558,N_9561,N_9562,N_9563,N_9564,N_9565,N_9567,N_9568,N_9572,N_9576,N_9578,N_9581,N_9584,N_9586,N_9587,N_9589,N_9590,N_9593,N_9599,N_9600,N_9602,N_9603,N_9606,N_9607,N_9608,N_9610,N_9611,N_9615,N_9616,N_9620,N_9621,N_9622,N_9624,N_9627,N_9628,N_9629,N_9630,N_9631,N_9638,N_9641,N_9642,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9652,N_9653,N_9656,N_9657,N_9659,N_9660,N_9661,N_9665,N_9666,N_9668,N_9670,N_9673,N_9676,N_9678,N_9680,N_9682,N_9683,N_9684,N_9685,N_9686,N_9690,N_9691,N_9692,N_9693,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9702,N_9703,N_9704,N_9709,N_9710,N_9712,N_9717,N_9718,N_9724,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9734,N_9735,N_9737,N_9738,N_9739,N_9741,N_9743,N_9745,N_9746,N_9747,N_9749,N_9751,N_9752,N_9753,N_9754,N_9758,N_9759,N_9761,N_9762,N_9764,N_9768,N_9769,N_9771,N_9776,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9787,N_9789,N_9790,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9803,N_9804,N_9805,N_9807,N_9808,N_9811,N_9813,N_9814,N_9819,N_9820,N_9821,N_9822,N_9823,N_9825,N_9827,N_9829,N_9830,N_9832,N_9833,N_9834,N_9835,N_9837,N_9840,N_9841,N_9842,N_9845,N_9846,N_9848,N_9849,N_9850,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9862,N_9864,N_9866,N_9867,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9891,N_9892,N_9897,N_9901,N_9905,N_9906,N_9907,N_9908,N_9909,N_9911,N_9916,N_9919,N_9920,N_9922,N_9923,N_9926,N_9927,N_9928,N_9929,N_9930,N_9932,N_9933,N_9935,N_9937,N_9939,N_9941,N_9942,N_9945,N_9946,N_9952,N_9953,N_9954,N_9956,N_9959,N_9962,N_9966,N_9967,N_9968,N_9969,N_9971,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9982,N_9985,N_9986,N_9988,N_9989,N_9990,N_9991,N_9993,N_9995,N_9997,N_9998,N_9999;
nor U0 (N_0,In_147,In_2);
nor U1 (N_1,In_76,In_482);
or U2 (N_2,In_185,In_276);
nand U3 (N_3,In_573,In_626);
nor U4 (N_4,In_907,In_307);
or U5 (N_5,In_43,In_240);
nor U6 (N_6,In_989,In_612);
or U7 (N_7,In_685,In_505);
or U8 (N_8,In_911,In_639);
and U9 (N_9,In_69,In_208);
nand U10 (N_10,In_705,In_228);
or U11 (N_11,In_458,In_812);
nand U12 (N_12,In_818,In_938);
or U13 (N_13,In_936,In_671);
nor U14 (N_14,In_85,In_679);
nand U15 (N_15,In_686,In_214);
or U16 (N_16,In_105,In_328);
nor U17 (N_17,In_922,In_225);
nor U18 (N_18,In_864,In_319);
nand U19 (N_19,In_39,In_150);
and U20 (N_20,In_347,In_336);
and U21 (N_21,In_879,In_599);
and U22 (N_22,In_921,In_721);
or U23 (N_23,In_764,In_650);
or U24 (N_24,In_253,In_28);
and U25 (N_25,In_373,In_83);
and U26 (N_26,In_412,In_992);
nor U27 (N_27,In_905,In_937);
nand U28 (N_28,In_116,In_115);
and U29 (N_29,In_29,In_748);
nor U30 (N_30,In_407,In_57);
nor U31 (N_31,In_746,In_363);
and U32 (N_32,In_545,In_689);
xor U33 (N_33,In_168,In_435);
or U34 (N_34,In_522,In_80);
nor U35 (N_35,In_733,In_598);
nor U36 (N_36,In_575,In_957);
nand U37 (N_37,In_148,In_813);
or U38 (N_38,In_223,In_273);
and U39 (N_39,In_314,In_695);
and U40 (N_40,In_279,In_299);
or U41 (N_41,In_187,In_403);
and U42 (N_42,In_1,In_344);
nor U43 (N_43,In_133,In_761);
and U44 (N_44,In_313,In_296);
or U45 (N_45,In_239,In_350);
and U46 (N_46,In_975,In_574);
nor U47 (N_47,In_884,In_503);
xnor U48 (N_48,In_123,In_739);
nor U49 (N_49,In_162,In_742);
nand U50 (N_50,In_471,In_124);
nand U51 (N_51,In_196,In_656);
nor U52 (N_52,In_953,In_252);
nor U53 (N_53,In_785,In_464);
and U54 (N_54,In_60,In_384);
nand U55 (N_55,In_469,In_920);
or U56 (N_56,In_21,In_615);
nand U57 (N_57,In_231,In_594);
or U58 (N_58,In_362,In_206);
or U59 (N_59,In_32,In_366);
nand U60 (N_60,In_266,In_845);
and U61 (N_61,In_811,In_275);
nand U62 (N_62,In_866,In_112);
or U63 (N_63,In_788,In_341);
or U64 (N_64,In_747,In_767);
or U65 (N_65,In_491,In_357);
nor U66 (N_66,In_199,In_261);
or U67 (N_67,In_258,In_862);
nand U68 (N_68,In_380,In_566);
nand U69 (N_69,In_146,In_91);
and U70 (N_70,In_847,In_918);
or U71 (N_71,In_257,In_932);
or U72 (N_72,In_820,In_359);
or U73 (N_73,In_236,In_106);
nor U74 (N_74,In_409,In_321);
or U75 (N_75,In_803,In_644);
and U76 (N_76,In_438,In_432);
nand U77 (N_77,In_801,In_8);
nand U78 (N_78,In_455,In_474);
nor U79 (N_79,In_323,In_465);
nor U80 (N_80,In_923,In_487);
and U81 (N_81,In_293,In_641);
nand U82 (N_82,In_578,In_821);
or U83 (N_83,In_254,In_400);
nand U84 (N_84,In_84,In_183);
nand U85 (N_85,In_556,In_593);
nand U86 (N_86,In_349,In_824);
or U87 (N_87,In_743,In_779);
nand U88 (N_88,In_842,In_625);
and U89 (N_89,In_834,In_451);
and U90 (N_90,In_128,In_353);
nand U91 (N_91,In_521,In_961);
nand U92 (N_92,In_62,In_483);
or U93 (N_93,In_145,In_394);
nand U94 (N_94,In_885,In_881);
and U95 (N_95,In_745,In_850);
and U96 (N_96,In_832,In_86);
and U97 (N_97,In_538,In_586);
nor U98 (N_98,In_81,In_662);
nor U99 (N_99,In_246,In_98);
or U100 (N_100,In_502,In_172);
nand U101 (N_101,In_161,In_496);
nor U102 (N_102,In_376,In_697);
nand U103 (N_103,In_778,In_609);
and U104 (N_104,In_737,In_655);
or U105 (N_105,In_910,In_681);
nand U106 (N_106,In_383,In_342);
nand U107 (N_107,In_659,In_237);
nand U108 (N_108,In_12,In_125);
or U109 (N_109,In_762,In_372);
nand U110 (N_110,In_719,In_295);
nor U111 (N_111,In_444,In_523);
or U112 (N_112,In_893,In_960);
xor U113 (N_113,In_683,In_647);
and U114 (N_114,In_859,In_776);
and U115 (N_115,In_397,In_54);
nor U116 (N_116,In_871,In_805);
nor U117 (N_117,In_5,In_423);
nor U118 (N_118,In_951,In_622);
or U119 (N_119,In_526,In_520);
and U120 (N_120,In_63,In_638);
nand U121 (N_121,In_354,In_170);
and U122 (N_122,In_408,In_964);
and U123 (N_123,In_554,In_138);
and U124 (N_124,In_606,In_485);
nor U125 (N_125,In_666,In_959);
nand U126 (N_126,In_463,In_867);
and U127 (N_127,In_238,In_7);
nor U128 (N_128,In_101,In_445);
and U129 (N_129,In_391,In_934);
nor U130 (N_130,In_816,In_188);
nand U131 (N_131,In_795,In_506);
or U132 (N_132,In_969,In_770);
and U133 (N_133,In_660,In_591);
and U134 (N_134,In_164,In_944);
nand U135 (N_135,In_930,In_282);
and U136 (N_136,In_153,In_744);
or U137 (N_137,In_830,In_272);
nor U138 (N_138,In_6,In_348);
nand U139 (N_139,In_840,In_883);
nor U140 (N_140,In_13,In_904);
nor U141 (N_141,In_614,In_725);
nand U142 (N_142,In_220,In_175);
nand U143 (N_143,In_571,In_548);
nor U144 (N_144,In_413,In_14);
and U145 (N_145,In_815,In_632);
nand U146 (N_146,In_939,In_966);
nand U147 (N_147,In_58,In_418);
or U148 (N_148,In_994,In_310);
nor U149 (N_149,In_66,In_304);
or U150 (N_150,In_916,In_687);
and U151 (N_151,In_972,In_207);
or U152 (N_152,In_479,In_473);
and U153 (N_153,In_322,In_20);
nand U154 (N_154,In_298,In_750);
nand U155 (N_155,In_781,In_46);
nand U156 (N_156,In_387,In_169);
and U157 (N_157,In_792,In_259);
and U158 (N_158,In_540,In_51);
nor U159 (N_159,In_552,In_915);
or U160 (N_160,In_771,In_769);
and U161 (N_161,In_967,In_588);
nand U162 (N_162,In_617,In_592);
and U163 (N_163,In_467,In_203);
nand U164 (N_164,In_814,In_962);
nand U165 (N_165,In_835,In_182);
and U166 (N_166,In_596,In_783);
nor U167 (N_167,In_708,In_416);
nor U168 (N_168,In_952,In_848);
or U169 (N_169,In_171,In_700);
nor U170 (N_170,In_600,In_649);
nor U171 (N_171,In_541,In_525);
nand U172 (N_172,In_947,In_292);
and U173 (N_173,In_255,In_470);
nand U174 (N_174,In_59,In_104);
and U175 (N_175,In_368,In_901);
and U176 (N_176,In_621,In_657);
or U177 (N_177,In_518,In_958);
nand U178 (N_178,In_831,In_836);
or U179 (N_179,In_11,In_977);
nand U180 (N_180,In_855,In_702);
xnor U181 (N_181,In_318,In_999);
and U182 (N_182,In_204,In_753);
nand U183 (N_183,In_511,In_144);
nand U184 (N_184,In_449,In_773);
and U185 (N_185,In_232,In_378);
and U186 (N_186,In_306,In_218);
or U187 (N_187,In_330,In_61);
nor U188 (N_188,In_47,In_24);
or U189 (N_189,In_942,In_131);
or U190 (N_190,In_197,In_555);
nor U191 (N_191,In_443,In_324);
or U192 (N_192,In_72,In_121);
and U193 (N_193,In_235,In_134);
nand U194 (N_194,In_544,In_210);
and U195 (N_195,In_664,In_414);
or U196 (N_196,In_417,In_120);
and U197 (N_197,In_281,In_114);
or U198 (N_198,In_287,In_283);
nor U199 (N_199,In_732,In_529);
nand U200 (N_200,In_559,In_519);
nor U201 (N_201,In_233,In_722);
nor U202 (N_202,In_530,In_741);
or U203 (N_203,In_846,In_434);
nand U204 (N_204,In_853,In_422);
or U205 (N_205,In_68,In_804);
nor U206 (N_206,In_429,In_177);
nand U207 (N_207,In_256,In_558);
or U208 (N_208,In_174,In_466);
nor U209 (N_209,In_668,In_995);
nor U210 (N_210,In_978,In_179);
or U211 (N_211,In_262,In_894);
nand U212 (N_212,In_67,In_565);
nor U213 (N_213,In_288,In_583);
nand U214 (N_214,In_335,In_286);
nor U215 (N_215,In_97,In_189);
nor U216 (N_216,In_878,In_221);
nand U217 (N_217,In_343,In_714);
nand U218 (N_218,In_504,In_532);
nand U219 (N_219,In_49,In_637);
and U220 (N_220,In_900,In_401);
or U221 (N_221,In_410,In_265);
or U222 (N_222,In_9,In_277);
nand U223 (N_223,In_452,In_667);
and U224 (N_224,In_152,In_151);
and U225 (N_225,In_488,In_178);
nand U226 (N_226,In_984,In_917);
or U227 (N_227,In_946,In_988);
nand U228 (N_228,In_379,In_680);
or U229 (N_229,In_56,In_316);
nor U230 (N_230,In_800,In_3);
and U231 (N_231,In_982,In_19);
or U232 (N_232,In_456,In_828);
nor U233 (N_233,In_833,In_186);
nand U234 (N_234,In_102,In_751);
or U235 (N_235,In_852,In_109);
and U236 (N_236,In_300,In_364);
or U237 (N_237,In_727,In_285);
nand U238 (N_238,In_774,In_809);
or U239 (N_239,In_549,In_396);
and U240 (N_240,In_513,In_297);
nor U241 (N_241,In_360,In_428);
nor U242 (N_242,In_242,In_79);
nor U243 (N_243,In_216,In_375);
or U244 (N_244,In_913,In_707);
and U245 (N_245,In_797,In_858);
nand U246 (N_246,In_440,In_584);
nand U247 (N_247,In_215,In_611);
or U248 (N_248,In_636,In_669);
or U249 (N_249,In_499,In_829);
nor U250 (N_250,In_572,In_709);
nor U251 (N_251,In_587,In_699);
nand U252 (N_252,In_241,In_30);
or U253 (N_253,In_176,In_457);
and U254 (N_254,In_624,In_926);
and U255 (N_255,In_949,In_385);
or U256 (N_256,In_654,In_437);
xor U257 (N_257,In_759,In_426);
or U258 (N_258,In_524,In_880);
nor U259 (N_259,In_280,In_462);
nor U260 (N_260,In_735,In_997);
nand U261 (N_261,In_736,In_4);
nor U262 (N_262,In_585,In_531);
or U263 (N_263,In_720,In_561);
or U264 (N_264,In_857,In_854);
nor U265 (N_265,In_912,In_516);
nand U266 (N_266,In_230,In_201);
nor U267 (N_267,In_431,In_244);
nor U268 (N_268,In_663,In_406);
nor U269 (N_269,In_251,In_874);
and U270 (N_270,In_645,In_260);
nor U271 (N_271,In_553,In_222);
nor U272 (N_272,In_477,In_983);
nand U273 (N_273,In_768,In_547);
nand U274 (N_274,In_710,In_790);
nand U275 (N_275,In_184,In_390);
or U276 (N_276,In_843,In_212);
and U277 (N_277,In_122,In_26);
nand U278 (N_278,In_369,In_90);
nor U279 (N_279,In_711,In_421);
or U280 (N_280,In_48,In_358);
nand U281 (N_281,In_264,In_892);
nor U282 (N_282,In_500,In_510);
nor U283 (N_283,In_906,In_427);
or U284 (N_284,In_37,In_929);
or U285 (N_285,In_851,In_158);
nor U286 (N_286,In_326,In_629);
nor U287 (N_287,In_154,In_633);
and U288 (N_288,In_448,In_684);
or U289 (N_289,In_974,In_726);
xnor U290 (N_290,In_193,In_17);
or U291 (N_291,In_163,In_772);
or U292 (N_292,In_924,In_602);
and U293 (N_293,In_863,In_870);
and U294 (N_294,In_963,In_317);
and U295 (N_295,In_758,In_284);
or U296 (N_296,In_908,In_712);
or U297 (N_297,In_998,In_381);
or U298 (N_298,In_113,In_673);
nand U299 (N_299,In_333,In_940);
and U300 (N_300,In_601,In_0);
nor U301 (N_301,In_579,In_291);
nor U302 (N_302,In_945,In_430);
nand U303 (N_303,In_425,In_34);
nor U304 (N_304,In_87,In_393);
nor U305 (N_305,In_875,In_620);
nand U306 (N_306,In_674,In_787);
or U307 (N_307,In_899,In_895);
or U308 (N_308,In_33,In_570);
nor U309 (N_309,In_305,In_877);
or U310 (N_310,In_569,In_143);
or U311 (N_311,In_92,In_882);
nand U312 (N_312,In_191,In_688);
and U313 (N_313,In_868,In_527);
nor U314 (N_314,In_42,In_370);
nand U315 (N_315,In_386,In_634);
nand U316 (N_316,In_919,In_311);
and U317 (N_317,In_546,In_22);
or U318 (N_318,In_607,In_166);
nor U319 (N_319,In_971,In_447);
nand U320 (N_320,In_52,In_195);
nor U321 (N_321,In_325,In_399);
or U322 (N_322,In_740,In_202);
nand U323 (N_323,In_65,In_490);
nand U324 (N_324,In_514,In_234);
nand U325 (N_325,In_970,In_653);
nand U326 (N_326,In_716,In_346);
xnor U327 (N_327,In_563,In_95);
and U328 (N_328,In_534,In_229);
and U329 (N_329,In_658,In_564);
or U330 (N_330,In_249,In_613);
and U331 (N_331,In_623,In_796);
or U332 (N_332,In_903,In_289);
nor U333 (N_333,In_642,In_860);
and U334 (N_334,In_180,In_107);
and U335 (N_335,In_312,In_701);
nor U336 (N_336,In_135,In_139);
nor U337 (N_337,In_337,In_888);
and U338 (N_338,In_137,In_44);
and U339 (N_339,In_551,In_749);
nor U340 (N_340,In_424,In_476);
and U341 (N_341,In_351,In_765);
nor U342 (N_342,In_539,In_766);
nand U343 (N_343,In_165,In_799);
nor U344 (N_344,In_340,In_806);
nor U345 (N_345,In_108,In_25);
nor U346 (N_346,In_294,In_509);
nor U347 (N_347,In_693,In_808);
nor U348 (N_348,In_315,In_398);
and U349 (N_349,In_619,In_439);
and U350 (N_350,In_590,In_224);
nand U351 (N_351,In_752,In_478);
or U352 (N_352,In_757,In_724);
nor U353 (N_353,In_392,In_149);
or U354 (N_354,In_338,In_278);
nor U355 (N_355,In_979,In_595);
or U356 (N_356,In_75,In_494);
nor U357 (N_357,In_717,In_303);
or U358 (N_358,In_713,In_651);
nand U359 (N_359,In_980,In_446);
or U360 (N_360,In_486,In_382);
nand U361 (N_361,In_802,In_301);
and U362 (N_362,In_755,In_492);
nand U363 (N_363,In_100,In_395);
nand U364 (N_364,In_205,In_226);
and U365 (N_365,In_460,In_955);
nor U366 (N_366,In_628,In_643);
nand U367 (N_367,In_608,In_672);
nor U368 (N_368,In_82,In_433);
or U369 (N_369,In_793,In_371);
nor U370 (N_370,In_71,In_64);
nor U371 (N_371,In_985,In_302);
or U372 (N_372,In_898,In_118);
nor U373 (N_373,In_675,In_27);
nand U374 (N_374,In_826,In_198);
and U375 (N_375,In_497,In_646);
or U376 (N_376,In_111,In_484);
nor U377 (N_377,In_780,In_495);
nand U378 (N_378,In_876,In_308);
nor U379 (N_379,In_18,In_55);
nand U380 (N_380,In_243,In_130);
and U381 (N_381,In_132,In_290);
and U382 (N_382,In_784,In_856);
nor U383 (N_383,In_475,In_38);
or U384 (N_384,In_692,In_227);
nor U385 (N_385,In_419,In_156);
nor U386 (N_386,In_167,In_515);
nand U387 (N_387,In_827,In_786);
and U388 (N_388,In_441,In_420);
nand U389 (N_389,In_190,In_40);
nand U390 (N_390,In_309,In_16);
and U391 (N_391,In_823,In_248);
nand U392 (N_392,In_789,In_782);
nand U393 (N_393,In_603,In_956);
nor U394 (N_394,In_209,In_537);
xnor U395 (N_395,In_192,In_247);
or U396 (N_396,In_567,In_798);
nor U397 (N_397,In_140,In_844);
nand U398 (N_398,In_610,In_332);
nor U399 (N_399,In_173,In_703);
nor U400 (N_400,In_127,In_159);
and U401 (N_401,In_734,In_715);
or U402 (N_402,In_652,In_869);
nor U403 (N_403,In_914,In_891);
nor U404 (N_404,In_691,In_41);
nand U405 (N_405,In_760,In_838);
nor U406 (N_406,In_630,In_15);
and U407 (N_407,In_542,In_841);
and U408 (N_408,In_902,In_480);
nor U409 (N_409,In_678,In_738);
nor U410 (N_410,In_694,In_690);
nand U411 (N_411,In_157,In_718);
or U412 (N_412,In_129,In_508);
nor U413 (N_413,In_987,In_777);
nand U414 (N_414,In_450,In_896);
nor U415 (N_415,In_897,In_817);
or U416 (N_416,In_461,In_459);
or U417 (N_417,In_493,In_50);
nand U418 (N_418,In_928,In_991);
nor U419 (N_419,In_402,In_489);
nor U420 (N_420,In_512,In_339);
xnor U421 (N_421,In_635,In_211);
nor U422 (N_422,In_200,In_23);
and U423 (N_423,In_365,In_976);
nand U424 (N_424,In_141,In_94);
nand U425 (N_425,In_36,In_819);
nor U426 (N_426,In_730,In_676);
nand U427 (N_427,In_909,In_731);
nand U428 (N_428,In_754,In_160);
nor U429 (N_429,In_589,In_388);
nand U430 (N_430,In_270,In_577);
and U431 (N_431,In_950,In_810);
or U432 (N_432,In_698,In_73);
nor U433 (N_433,In_45,In_973);
nor U434 (N_434,In_791,In_374);
nor U435 (N_435,In_965,In_933);
or U436 (N_436,In_861,In_93);
and U437 (N_437,In_377,In_329);
or U438 (N_438,In_88,In_728);
and U439 (N_439,In_35,In_729);
and U440 (N_440,In_155,In_581);
nand U441 (N_441,In_181,In_562);
nor U442 (N_442,In_996,In_568);
and U443 (N_443,In_775,In_361);
nand U444 (N_444,In_631,In_948);
or U445 (N_445,In_849,In_99);
nor U446 (N_446,In_763,In_943);
nand U447 (N_447,In_356,In_661);
xnor U448 (N_448,In_126,In_543);
or U449 (N_449,In_136,In_405);
and U450 (N_450,In_935,In_696);
nor U451 (N_451,In_404,In_890);
or U452 (N_452,In_550,In_822);
and U453 (N_453,In_331,In_263);
and U454 (N_454,In_825,In_528);
nor U455 (N_455,In_665,In_536);
and U456 (N_456,In_472,In_367);
nor U457 (N_457,In_453,In_271);
nor U458 (N_458,In_557,In_670);
and U459 (N_459,In_886,In_411);
and U460 (N_460,In_535,In_931);
nor U461 (N_461,In_250,In_345);
nand U462 (N_462,In_89,In_10);
or U463 (N_463,In_70,In_968);
and U464 (N_464,In_119,In_103);
nor U465 (N_465,In_219,In_267);
and U466 (N_466,In_274,In_481);
nor U467 (N_467,In_677,In_501);
or U468 (N_468,In_604,In_327);
or U469 (N_469,In_468,In_320);
nor U470 (N_470,In_269,In_723);
or U471 (N_471,In_704,In_53);
nand U472 (N_472,In_533,In_78);
and U473 (N_473,In_213,In_245);
and U474 (N_474,In_576,In_142);
nor U475 (N_475,In_442,In_807);
and U476 (N_476,In_77,In_981);
nand U477 (N_477,In_560,In_682);
nor U478 (N_478,In_597,In_865);
nand U479 (N_479,In_117,In_706);
or U480 (N_480,In_839,In_616);
nand U481 (N_481,In_986,In_648);
or U482 (N_482,In_217,In_941);
and U483 (N_483,In_640,In_74);
nor U484 (N_484,In_580,In_110);
nand U485 (N_485,In_507,In_794);
or U486 (N_486,In_355,In_872);
nand U487 (N_487,In_889,In_990);
and U488 (N_488,In_96,In_756);
and U489 (N_489,In_927,In_582);
and U490 (N_490,In_605,In_415);
or U491 (N_491,In_498,In_925);
nand U492 (N_492,In_436,In_887);
nand U493 (N_493,In_837,In_268);
and U494 (N_494,In_517,In_618);
and U495 (N_495,In_31,In_993);
or U496 (N_496,In_194,In_454);
and U497 (N_497,In_389,In_352);
nand U498 (N_498,In_873,In_334);
nand U499 (N_499,In_954,In_627);
nor U500 (N_500,In_826,In_354);
or U501 (N_501,In_935,In_384);
and U502 (N_502,In_20,In_740);
nand U503 (N_503,In_661,In_497);
or U504 (N_504,In_738,In_291);
and U505 (N_505,In_195,In_874);
nor U506 (N_506,In_221,In_988);
or U507 (N_507,In_622,In_645);
and U508 (N_508,In_193,In_240);
nor U509 (N_509,In_288,In_521);
or U510 (N_510,In_290,In_270);
and U511 (N_511,In_719,In_941);
or U512 (N_512,In_173,In_379);
nand U513 (N_513,In_392,In_418);
nor U514 (N_514,In_684,In_846);
or U515 (N_515,In_522,In_82);
nor U516 (N_516,In_389,In_535);
or U517 (N_517,In_409,In_676);
and U518 (N_518,In_826,In_884);
nor U519 (N_519,In_335,In_860);
or U520 (N_520,In_90,In_190);
nand U521 (N_521,In_920,In_957);
and U522 (N_522,In_875,In_693);
and U523 (N_523,In_654,In_158);
nand U524 (N_524,In_973,In_499);
and U525 (N_525,In_795,In_37);
nand U526 (N_526,In_955,In_790);
or U527 (N_527,In_110,In_920);
nand U528 (N_528,In_42,In_45);
and U529 (N_529,In_45,In_669);
nand U530 (N_530,In_983,In_203);
nor U531 (N_531,In_985,In_822);
and U532 (N_532,In_381,In_824);
or U533 (N_533,In_786,In_421);
or U534 (N_534,In_448,In_735);
nor U535 (N_535,In_867,In_282);
nor U536 (N_536,In_575,In_531);
nor U537 (N_537,In_487,In_791);
nand U538 (N_538,In_770,In_436);
and U539 (N_539,In_699,In_763);
nor U540 (N_540,In_909,In_639);
or U541 (N_541,In_969,In_836);
nor U542 (N_542,In_186,In_382);
and U543 (N_543,In_777,In_332);
nor U544 (N_544,In_824,In_936);
nor U545 (N_545,In_665,In_758);
nand U546 (N_546,In_964,In_618);
or U547 (N_547,In_737,In_987);
nand U548 (N_548,In_982,In_347);
or U549 (N_549,In_125,In_488);
nor U550 (N_550,In_800,In_271);
and U551 (N_551,In_953,In_115);
nor U552 (N_552,In_860,In_998);
or U553 (N_553,In_984,In_80);
nand U554 (N_554,In_190,In_694);
or U555 (N_555,In_491,In_668);
nand U556 (N_556,In_856,In_973);
and U557 (N_557,In_186,In_999);
nor U558 (N_558,In_187,In_563);
and U559 (N_559,In_69,In_570);
and U560 (N_560,In_246,In_698);
and U561 (N_561,In_726,In_301);
nor U562 (N_562,In_26,In_111);
and U563 (N_563,In_588,In_120);
and U564 (N_564,In_797,In_357);
nand U565 (N_565,In_103,In_711);
or U566 (N_566,In_455,In_791);
or U567 (N_567,In_199,In_851);
nor U568 (N_568,In_814,In_642);
and U569 (N_569,In_888,In_822);
nand U570 (N_570,In_820,In_35);
and U571 (N_571,In_408,In_813);
or U572 (N_572,In_280,In_535);
or U573 (N_573,In_609,In_844);
or U574 (N_574,In_809,In_243);
or U575 (N_575,In_930,In_47);
nand U576 (N_576,In_97,In_315);
or U577 (N_577,In_296,In_347);
or U578 (N_578,In_721,In_652);
nand U579 (N_579,In_440,In_415);
nor U580 (N_580,In_327,In_32);
and U581 (N_581,In_143,In_246);
or U582 (N_582,In_587,In_363);
nor U583 (N_583,In_44,In_767);
nor U584 (N_584,In_330,In_59);
or U585 (N_585,In_760,In_165);
and U586 (N_586,In_905,In_430);
and U587 (N_587,In_534,In_736);
and U588 (N_588,In_340,In_538);
and U589 (N_589,In_654,In_542);
or U590 (N_590,In_277,In_695);
or U591 (N_591,In_723,In_897);
nor U592 (N_592,In_158,In_161);
nand U593 (N_593,In_841,In_822);
nand U594 (N_594,In_500,In_472);
or U595 (N_595,In_853,In_284);
nor U596 (N_596,In_62,In_818);
or U597 (N_597,In_844,In_658);
nand U598 (N_598,In_725,In_236);
and U599 (N_599,In_676,In_826);
nor U600 (N_600,In_570,In_186);
nor U601 (N_601,In_86,In_841);
nor U602 (N_602,In_836,In_714);
nand U603 (N_603,In_721,In_583);
nand U604 (N_604,In_509,In_965);
nand U605 (N_605,In_523,In_209);
nand U606 (N_606,In_317,In_818);
nand U607 (N_607,In_618,In_703);
nand U608 (N_608,In_106,In_668);
nand U609 (N_609,In_690,In_351);
nand U610 (N_610,In_512,In_508);
or U611 (N_611,In_396,In_759);
nand U612 (N_612,In_459,In_978);
nand U613 (N_613,In_239,In_551);
and U614 (N_614,In_383,In_850);
nor U615 (N_615,In_632,In_227);
and U616 (N_616,In_647,In_456);
nand U617 (N_617,In_371,In_885);
or U618 (N_618,In_515,In_821);
or U619 (N_619,In_625,In_650);
or U620 (N_620,In_575,In_996);
nand U621 (N_621,In_832,In_744);
nand U622 (N_622,In_347,In_949);
nor U623 (N_623,In_669,In_872);
nor U624 (N_624,In_193,In_251);
or U625 (N_625,In_398,In_343);
nand U626 (N_626,In_695,In_683);
and U627 (N_627,In_748,In_643);
nand U628 (N_628,In_238,In_78);
nor U629 (N_629,In_549,In_407);
or U630 (N_630,In_991,In_271);
and U631 (N_631,In_108,In_402);
and U632 (N_632,In_286,In_430);
and U633 (N_633,In_247,In_625);
nor U634 (N_634,In_113,In_442);
nand U635 (N_635,In_782,In_641);
xor U636 (N_636,In_646,In_537);
xnor U637 (N_637,In_484,In_766);
and U638 (N_638,In_224,In_912);
and U639 (N_639,In_891,In_924);
and U640 (N_640,In_574,In_473);
or U641 (N_641,In_827,In_346);
or U642 (N_642,In_327,In_962);
nor U643 (N_643,In_86,In_155);
or U644 (N_644,In_910,In_398);
or U645 (N_645,In_706,In_124);
or U646 (N_646,In_533,In_531);
and U647 (N_647,In_962,In_245);
and U648 (N_648,In_223,In_330);
nand U649 (N_649,In_258,In_683);
and U650 (N_650,In_589,In_551);
nand U651 (N_651,In_253,In_291);
nand U652 (N_652,In_657,In_167);
nand U653 (N_653,In_142,In_958);
or U654 (N_654,In_20,In_844);
nand U655 (N_655,In_630,In_874);
or U656 (N_656,In_469,In_162);
and U657 (N_657,In_925,In_24);
nand U658 (N_658,In_769,In_532);
nor U659 (N_659,In_364,In_4);
nand U660 (N_660,In_897,In_656);
and U661 (N_661,In_796,In_41);
nor U662 (N_662,In_612,In_665);
nand U663 (N_663,In_742,In_557);
nand U664 (N_664,In_989,In_182);
nor U665 (N_665,In_714,In_477);
and U666 (N_666,In_988,In_793);
nor U667 (N_667,In_788,In_755);
and U668 (N_668,In_444,In_795);
or U669 (N_669,In_892,In_471);
or U670 (N_670,In_983,In_842);
or U671 (N_671,In_388,In_745);
nor U672 (N_672,In_683,In_903);
and U673 (N_673,In_625,In_187);
or U674 (N_674,In_19,In_913);
and U675 (N_675,In_163,In_825);
and U676 (N_676,In_173,In_935);
nand U677 (N_677,In_107,In_330);
or U678 (N_678,In_580,In_991);
and U679 (N_679,In_274,In_198);
nor U680 (N_680,In_620,In_178);
or U681 (N_681,In_846,In_204);
nand U682 (N_682,In_993,In_210);
nor U683 (N_683,In_362,In_448);
or U684 (N_684,In_133,In_171);
or U685 (N_685,In_369,In_301);
or U686 (N_686,In_958,In_526);
and U687 (N_687,In_554,In_149);
and U688 (N_688,In_642,In_291);
and U689 (N_689,In_969,In_806);
nor U690 (N_690,In_758,In_873);
nand U691 (N_691,In_852,In_314);
and U692 (N_692,In_220,In_783);
or U693 (N_693,In_904,In_10);
nand U694 (N_694,In_470,In_848);
nand U695 (N_695,In_311,In_200);
nor U696 (N_696,In_379,In_977);
nand U697 (N_697,In_246,In_838);
nor U698 (N_698,In_286,In_884);
or U699 (N_699,In_409,In_520);
or U700 (N_700,In_577,In_321);
nor U701 (N_701,In_720,In_810);
nand U702 (N_702,In_582,In_531);
nor U703 (N_703,In_775,In_127);
or U704 (N_704,In_360,In_344);
nand U705 (N_705,In_615,In_692);
or U706 (N_706,In_65,In_103);
nand U707 (N_707,In_566,In_332);
and U708 (N_708,In_199,In_752);
and U709 (N_709,In_259,In_892);
nand U710 (N_710,In_286,In_199);
and U711 (N_711,In_946,In_547);
nor U712 (N_712,In_118,In_749);
and U713 (N_713,In_436,In_993);
nand U714 (N_714,In_144,In_266);
and U715 (N_715,In_738,In_578);
nand U716 (N_716,In_576,In_795);
or U717 (N_717,In_50,In_177);
and U718 (N_718,In_130,In_588);
nor U719 (N_719,In_253,In_894);
nand U720 (N_720,In_163,In_200);
xor U721 (N_721,In_18,In_962);
or U722 (N_722,In_448,In_810);
or U723 (N_723,In_615,In_386);
and U724 (N_724,In_659,In_558);
nand U725 (N_725,In_59,In_907);
nand U726 (N_726,In_13,In_470);
nor U727 (N_727,In_887,In_36);
and U728 (N_728,In_997,In_357);
nor U729 (N_729,In_199,In_929);
or U730 (N_730,In_702,In_689);
nand U731 (N_731,In_375,In_51);
nand U732 (N_732,In_949,In_988);
or U733 (N_733,In_415,In_999);
nand U734 (N_734,In_129,In_266);
and U735 (N_735,In_888,In_932);
and U736 (N_736,In_602,In_8);
nand U737 (N_737,In_96,In_495);
nand U738 (N_738,In_840,In_133);
and U739 (N_739,In_964,In_299);
or U740 (N_740,In_833,In_785);
or U741 (N_741,In_509,In_314);
or U742 (N_742,In_337,In_71);
nand U743 (N_743,In_921,In_890);
or U744 (N_744,In_66,In_64);
nand U745 (N_745,In_212,In_750);
nor U746 (N_746,In_623,In_766);
or U747 (N_747,In_248,In_406);
and U748 (N_748,In_722,In_806);
nand U749 (N_749,In_370,In_451);
xor U750 (N_750,In_676,In_375);
and U751 (N_751,In_525,In_990);
nand U752 (N_752,In_682,In_820);
or U753 (N_753,In_847,In_772);
or U754 (N_754,In_96,In_473);
nand U755 (N_755,In_446,In_234);
or U756 (N_756,In_207,In_25);
nand U757 (N_757,In_898,In_901);
or U758 (N_758,In_647,In_511);
and U759 (N_759,In_693,In_698);
and U760 (N_760,In_706,In_381);
and U761 (N_761,In_211,In_289);
or U762 (N_762,In_716,In_862);
and U763 (N_763,In_732,In_763);
and U764 (N_764,In_328,In_39);
nor U765 (N_765,In_378,In_594);
or U766 (N_766,In_270,In_984);
nand U767 (N_767,In_131,In_204);
nand U768 (N_768,In_921,In_627);
and U769 (N_769,In_126,In_673);
nand U770 (N_770,In_514,In_941);
nor U771 (N_771,In_603,In_413);
and U772 (N_772,In_613,In_371);
nor U773 (N_773,In_307,In_462);
and U774 (N_774,In_684,In_649);
or U775 (N_775,In_662,In_350);
and U776 (N_776,In_331,In_87);
or U777 (N_777,In_355,In_768);
nor U778 (N_778,In_767,In_709);
nand U779 (N_779,In_792,In_955);
and U780 (N_780,In_941,In_439);
or U781 (N_781,In_36,In_528);
or U782 (N_782,In_865,In_885);
nor U783 (N_783,In_758,In_191);
and U784 (N_784,In_848,In_123);
or U785 (N_785,In_181,In_48);
nand U786 (N_786,In_732,In_38);
and U787 (N_787,In_203,In_721);
and U788 (N_788,In_869,In_882);
nand U789 (N_789,In_744,In_423);
or U790 (N_790,In_608,In_320);
nand U791 (N_791,In_642,In_297);
nand U792 (N_792,In_455,In_465);
and U793 (N_793,In_519,In_18);
or U794 (N_794,In_831,In_611);
or U795 (N_795,In_484,In_50);
and U796 (N_796,In_875,In_942);
nand U797 (N_797,In_615,In_214);
and U798 (N_798,In_820,In_301);
and U799 (N_799,In_418,In_676);
and U800 (N_800,In_215,In_468);
or U801 (N_801,In_799,In_465);
or U802 (N_802,In_747,In_885);
nand U803 (N_803,In_498,In_832);
nand U804 (N_804,In_171,In_140);
and U805 (N_805,In_916,In_764);
nand U806 (N_806,In_518,In_502);
or U807 (N_807,In_721,In_595);
or U808 (N_808,In_62,In_526);
or U809 (N_809,In_467,In_700);
nand U810 (N_810,In_305,In_278);
nor U811 (N_811,In_702,In_839);
and U812 (N_812,In_160,In_520);
and U813 (N_813,In_243,In_708);
and U814 (N_814,In_704,In_305);
nor U815 (N_815,In_938,In_452);
or U816 (N_816,In_34,In_311);
nand U817 (N_817,In_208,In_599);
nand U818 (N_818,In_287,In_686);
nor U819 (N_819,In_45,In_633);
or U820 (N_820,In_250,In_915);
nand U821 (N_821,In_691,In_34);
nor U822 (N_822,In_183,In_872);
nand U823 (N_823,In_236,In_686);
or U824 (N_824,In_185,In_614);
nand U825 (N_825,In_931,In_360);
and U826 (N_826,In_389,In_321);
and U827 (N_827,In_485,In_675);
nand U828 (N_828,In_792,In_140);
or U829 (N_829,In_543,In_398);
or U830 (N_830,In_129,In_295);
and U831 (N_831,In_847,In_285);
and U832 (N_832,In_620,In_531);
or U833 (N_833,In_399,In_355);
and U834 (N_834,In_808,In_50);
nor U835 (N_835,In_663,In_201);
or U836 (N_836,In_671,In_847);
nor U837 (N_837,In_710,In_233);
or U838 (N_838,In_14,In_603);
or U839 (N_839,In_961,In_325);
nand U840 (N_840,In_505,In_719);
nor U841 (N_841,In_302,In_239);
nand U842 (N_842,In_708,In_57);
nand U843 (N_843,In_388,In_733);
or U844 (N_844,In_129,In_261);
and U845 (N_845,In_173,In_88);
or U846 (N_846,In_330,In_615);
nand U847 (N_847,In_470,In_88);
nand U848 (N_848,In_259,In_812);
or U849 (N_849,In_988,In_7);
or U850 (N_850,In_317,In_98);
and U851 (N_851,In_527,In_99);
and U852 (N_852,In_219,In_519);
or U853 (N_853,In_187,In_979);
or U854 (N_854,In_185,In_750);
or U855 (N_855,In_941,In_548);
nand U856 (N_856,In_541,In_852);
and U857 (N_857,In_747,In_821);
or U858 (N_858,In_650,In_790);
and U859 (N_859,In_349,In_974);
nand U860 (N_860,In_737,In_60);
and U861 (N_861,In_659,In_474);
nor U862 (N_862,In_8,In_627);
and U863 (N_863,In_253,In_40);
nor U864 (N_864,In_122,In_292);
nor U865 (N_865,In_507,In_231);
nor U866 (N_866,In_923,In_826);
or U867 (N_867,In_185,In_855);
nand U868 (N_868,In_909,In_417);
nor U869 (N_869,In_902,In_767);
and U870 (N_870,In_579,In_650);
nor U871 (N_871,In_839,In_928);
or U872 (N_872,In_915,In_854);
nor U873 (N_873,In_28,In_855);
and U874 (N_874,In_434,In_866);
nor U875 (N_875,In_934,In_535);
or U876 (N_876,In_892,In_222);
or U877 (N_877,In_674,In_383);
nor U878 (N_878,In_669,In_227);
nor U879 (N_879,In_951,In_991);
nand U880 (N_880,In_240,In_987);
and U881 (N_881,In_635,In_33);
or U882 (N_882,In_718,In_974);
or U883 (N_883,In_450,In_731);
and U884 (N_884,In_182,In_72);
and U885 (N_885,In_565,In_805);
xor U886 (N_886,In_216,In_263);
and U887 (N_887,In_492,In_13);
nor U888 (N_888,In_9,In_743);
and U889 (N_889,In_728,In_349);
or U890 (N_890,In_145,In_474);
and U891 (N_891,In_339,In_299);
or U892 (N_892,In_848,In_95);
or U893 (N_893,In_96,In_255);
nand U894 (N_894,In_737,In_172);
nor U895 (N_895,In_174,In_726);
or U896 (N_896,In_834,In_933);
or U897 (N_897,In_448,In_329);
nor U898 (N_898,In_36,In_125);
or U899 (N_899,In_12,In_559);
or U900 (N_900,In_745,In_959);
or U901 (N_901,In_337,In_498);
and U902 (N_902,In_429,In_604);
and U903 (N_903,In_979,In_866);
nor U904 (N_904,In_674,In_40);
and U905 (N_905,In_76,In_586);
and U906 (N_906,In_976,In_261);
nand U907 (N_907,In_329,In_646);
nand U908 (N_908,In_963,In_942);
and U909 (N_909,In_165,In_223);
nand U910 (N_910,In_393,In_53);
or U911 (N_911,In_147,In_744);
nand U912 (N_912,In_946,In_363);
nor U913 (N_913,In_232,In_565);
nand U914 (N_914,In_624,In_855);
xnor U915 (N_915,In_989,In_652);
nor U916 (N_916,In_959,In_243);
and U917 (N_917,In_37,In_967);
nor U918 (N_918,In_975,In_588);
nor U919 (N_919,In_632,In_849);
or U920 (N_920,In_677,In_10);
or U921 (N_921,In_83,In_375);
nand U922 (N_922,In_200,In_454);
and U923 (N_923,In_79,In_864);
nand U924 (N_924,In_560,In_928);
or U925 (N_925,In_761,In_810);
and U926 (N_926,In_987,In_358);
and U927 (N_927,In_274,In_736);
and U928 (N_928,In_211,In_343);
nand U929 (N_929,In_746,In_3);
nand U930 (N_930,In_71,In_265);
nand U931 (N_931,In_900,In_468);
nand U932 (N_932,In_688,In_661);
nand U933 (N_933,In_628,In_538);
and U934 (N_934,In_693,In_379);
or U935 (N_935,In_155,In_140);
nor U936 (N_936,In_453,In_174);
and U937 (N_937,In_395,In_864);
or U938 (N_938,In_220,In_487);
nand U939 (N_939,In_107,In_699);
nor U940 (N_940,In_124,In_163);
nor U941 (N_941,In_190,In_675);
nor U942 (N_942,In_59,In_297);
nor U943 (N_943,In_927,In_388);
or U944 (N_944,In_382,In_322);
nand U945 (N_945,In_946,In_240);
nor U946 (N_946,In_10,In_445);
or U947 (N_947,In_192,In_89);
nor U948 (N_948,In_861,In_477);
and U949 (N_949,In_296,In_333);
nand U950 (N_950,In_561,In_249);
nor U951 (N_951,In_101,In_894);
and U952 (N_952,In_785,In_885);
nor U953 (N_953,In_890,In_419);
nor U954 (N_954,In_575,In_483);
nand U955 (N_955,In_817,In_149);
nor U956 (N_956,In_594,In_72);
or U957 (N_957,In_856,In_574);
nor U958 (N_958,In_632,In_171);
nand U959 (N_959,In_854,In_285);
or U960 (N_960,In_578,In_348);
nor U961 (N_961,In_282,In_411);
nand U962 (N_962,In_749,In_738);
nor U963 (N_963,In_36,In_490);
or U964 (N_964,In_83,In_46);
and U965 (N_965,In_357,In_178);
or U966 (N_966,In_450,In_45);
nand U967 (N_967,In_928,In_847);
or U968 (N_968,In_312,In_677);
and U969 (N_969,In_259,In_406);
or U970 (N_970,In_570,In_610);
nor U971 (N_971,In_768,In_504);
nand U972 (N_972,In_87,In_801);
nand U973 (N_973,In_631,In_396);
nand U974 (N_974,In_856,In_552);
nor U975 (N_975,In_878,In_546);
and U976 (N_976,In_939,In_876);
and U977 (N_977,In_59,In_236);
nor U978 (N_978,In_925,In_503);
nand U979 (N_979,In_769,In_785);
nor U980 (N_980,In_896,In_458);
or U981 (N_981,In_190,In_253);
or U982 (N_982,In_524,In_16);
or U983 (N_983,In_488,In_617);
nor U984 (N_984,In_605,In_632);
or U985 (N_985,In_616,In_674);
nand U986 (N_986,In_541,In_334);
nand U987 (N_987,In_293,In_733);
nand U988 (N_988,In_205,In_867);
nor U989 (N_989,In_172,In_320);
nor U990 (N_990,In_589,In_233);
nand U991 (N_991,In_663,In_258);
or U992 (N_992,In_473,In_331);
nor U993 (N_993,In_585,In_95);
and U994 (N_994,In_329,In_349);
nor U995 (N_995,In_51,In_962);
or U996 (N_996,In_400,In_966);
and U997 (N_997,In_499,In_953);
nand U998 (N_998,In_745,In_728);
nor U999 (N_999,In_655,In_279);
and U1000 (N_1000,In_100,In_795);
and U1001 (N_1001,In_713,In_313);
and U1002 (N_1002,In_230,In_53);
xor U1003 (N_1003,In_398,In_410);
nor U1004 (N_1004,In_201,In_520);
or U1005 (N_1005,In_584,In_619);
or U1006 (N_1006,In_391,In_311);
nor U1007 (N_1007,In_525,In_132);
nor U1008 (N_1008,In_755,In_352);
nand U1009 (N_1009,In_853,In_711);
nand U1010 (N_1010,In_334,In_859);
or U1011 (N_1011,In_685,In_209);
nor U1012 (N_1012,In_653,In_537);
and U1013 (N_1013,In_439,In_358);
nor U1014 (N_1014,In_481,In_897);
nor U1015 (N_1015,In_700,In_333);
nand U1016 (N_1016,In_136,In_978);
and U1017 (N_1017,In_180,In_279);
nor U1018 (N_1018,In_767,In_246);
or U1019 (N_1019,In_265,In_603);
and U1020 (N_1020,In_955,In_70);
nor U1021 (N_1021,In_537,In_997);
and U1022 (N_1022,In_189,In_978);
nand U1023 (N_1023,In_279,In_625);
nand U1024 (N_1024,In_203,In_764);
and U1025 (N_1025,In_299,In_437);
nand U1026 (N_1026,In_865,In_253);
or U1027 (N_1027,In_842,In_613);
nand U1028 (N_1028,In_395,In_729);
or U1029 (N_1029,In_612,In_360);
or U1030 (N_1030,In_703,In_434);
nand U1031 (N_1031,In_914,In_976);
nand U1032 (N_1032,In_496,In_582);
nand U1033 (N_1033,In_961,In_655);
nand U1034 (N_1034,In_27,In_171);
nor U1035 (N_1035,In_236,In_173);
nand U1036 (N_1036,In_920,In_763);
and U1037 (N_1037,In_455,In_996);
and U1038 (N_1038,In_365,In_848);
or U1039 (N_1039,In_44,In_606);
nand U1040 (N_1040,In_260,In_808);
nor U1041 (N_1041,In_330,In_540);
nand U1042 (N_1042,In_147,In_768);
and U1043 (N_1043,In_656,In_333);
nand U1044 (N_1044,In_270,In_60);
and U1045 (N_1045,In_940,In_306);
or U1046 (N_1046,In_189,In_498);
or U1047 (N_1047,In_518,In_827);
nand U1048 (N_1048,In_24,In_952);
nor U1049 (N_1049,In_555,In_191);
or U1050 (N_1050,In_209,In_495);
and U1051 (N_1051,In_758,In_489);
and U1052 (N_1052,In_655,In_623);
and U1053 (N_1053,In_907,In_30);
or U1054 (N_1054,In_337,In_214);
or U1055 (N_1055,In_331,In_401);
and U1056 (N_1056,In_846,In_20);
nor U1057 (N_1057,In_107,In_517);
and U1058 (N_1058,In_81,In_340);
or U1059 (N_1059,In_789,In_351);
and U1060 (N_1060,In_194,In_92);
nor U1061 (N_1061,In_710,In_153);
nor U1062 (N_1062,In_534,In_38);
and U1063 (N_1063,In_511,In_712);
or U1064 (N_1064,In_392,In_579);
or U1065 (N_1065,In_886,In_79);
and U1066 (N_1066,In_390,In_541);
or U1067 (N_1067,In_661,In_89);
or U1068 (N_1068,In_880,In_563);
nand U1069 (N_1069,In_930,In_776);
nand U1070 (N_1070,In_65,In_113);
nor U1071 (N_1071,In_962,In_156);
nor U1072 (N_1072,In_513,In_322);
nand U1073 (N_1073,In_913,In_74);
or U1074 (N_1074,In_678,In_770);
or U1075 (N_1075,In_539,In_33);
nor U1076 (N_1076,In_275,In_853);
and U1077 (N_1077,In_26,In_140);
nor U1078 (N_1078,In_451,In_155);
or U1079 (N_1079,In_400,In_349);
or U1080 (N_1080,In_272,In_475);
or U1081 (N_1081,In_753,In_769);
nand U1082 (N_1082,In_72,In_354);
and U1083 (N_1083,In_845,In_241);
and U1084 (N_1084,In_204,In_526);
nor U1085 (N_1085,In_977,In_330);
nand U1086 (N_1086,In_126,In_452);
nand U1087 (N_1087,In_63,In_959);
and U1088 (N_1088,In_865,In_549);
nor U1089 (N_1089,In_83,In_8);
or U1090 (N_1090,In_281,In_798);
or U1091 (N_1091,In_308,In_688);
or U1092 (N_1092,In_197,In_420);
or U1093 (N_1093,In_488,In_669);
nor U1094 (N_1094,In_593,In_327);
nor U1095 (N_1095,In_39,In_975);
nand U1096 (N_1096,In_63,In_805);
or U1097 (N_1097,In_18,In_964);
nand U1098 (N_1098,In_674,In_842);
and U1099 (N_1099,In_128,In_516);
nor U1100 (N_1100,In_395,In_941);
nand U1101 (N_1101,In_169,In_674);
nand U1102 (N_1102,In_646,In_147);
nor U1103 (N_1103,In_705,In_328);
xnor U1104 (N_1104,In_438,In_788);
nor U1105 (N_1105,In_272,In_181);
or U1106 (N_1106,In_418,In_929);
nor U1107 (N_1107,In_383,In_454);
nor U1108 (N_1108,In_501,In_783);
nand U1109 (N_1109,In_89,In_623);
and U1110 (N_1110,In_308,In_541);
nand U1111 (N_1111,In_170,In_621);
or U1112 (N_1112,In_313,In_72);
nand U1113 (N_1113,In_945,In_397);
nor U1114 (N_1114,In_40,In_728);
nand U1115 (N_1115,In_487,In_520);
nor U1116 (N_1116,In_404,In_643);
nand U1117 (N_1117,In_83,In_388);
nor U1118 (N_1118,In_630,In_389);
nor U1119 (N_1119,In_87,In_421);
or U1120 (N_1120,In_828,In_173);
nor U1121 (N_1121,In_287,In_603);
and U1122 (N_1122,In_535,In_103);
nor U1123 (N_1123,In_568,In_108);
or U1124 (N_1124,In_962,In_731);
nand U1125 (N_1125,In_177,In_713);
nand U1126 (N_1126,In_498,In_730);
nand U1127 (N_1127,In_567,In_728);
and U1128 (N_1128,In_154,In_366);
and U1129 (N_1129,In_299,In_123);
nor U1130 (N_1130,In_574,In_878);
and U1131 (N_1131,In_163,In_819);
or U1132 (N_1132,In_386,In_885);
and U1133 (N_1133,In_134,In_507);
nand U1134 (N_1134,In_63,In_411);
nand U1135 (N_1135,In_409,In_697);
and U1136 (N_1136,In_52,In_275);
or U1137 (N_1137,In_801,In_908);
and U1138 (N_1138,In_892,In_938);
or U1139 (N_1139,In_93,In_316);
nor U1140 (N_1140,In_517,In_532);
nor U1141 (N_1141,In_28,In_23);
nor U1142 (N_1142,In_374,In_840);
nand U1143 (N_1143,In_274,In_802);
nand U1144 (N_1144,In_10,In_724);
or U1145 (N_1145,In_520,In_957);
nor U1146 (N_1146,In_451,In_945);
nor U1147 (N_1147,In_359,In_464);
and U1148 (N_1148,In_466,In_502);
nand U1149 (N_1149,In_470,In_948);
nand U1150 (N_1150,In_290,In_859);
and U1151 (N_1151,In_902,In_518);
nor U1152 (N_1152,In_38,In_71);
nor U1153 (N_1153,In_214,In_592);
nand U1154 (N_1154,In_229,In_289);
xnor U1155 (N_1155,In_246,In_811);
or U1156 (N_1156,In_664,In_883);
or U1157 (N_1157,In_362,In_361);
or U1158 (N_1158,In_929,In_974);
nand U1159 (N_1159,In_275,In_865);
nand U1160 (N_1160,In_39,In_71);
or U1161 (N_1161,In_662,In_833);
nand U1162 (N_1162,In_872,In_751);
nand U1163 (N_1163,In_426,In_672);
and U1164 (N_1164,In_556,In_951);
and U1165 (N_1165,In_820,In_135);
nor U1166 (N_1166,In_200,In_665);
or U1167 (N_1167,In_268,In_158);
and U1168 (N_1168,In_347,In_100);
and U1169 (N_1169,In_856,In_643);
xor U1170 (N_1170,In_942,In_429);
or U1171 (N_1171,In_636,In_138);
nand U1172 (N_1172,In_150,In_898);
nand U1173 (N_1173,In_665,In_113);
or U1174 (N_1174,In_522,In_703);
or U1175 (N_1175,In_707,In_167);
nand U1176 (N_1176,In_675,In_88);
and U1177 (N_1177,In_271,In_533);
and U1178 (N_1178,In_749,In_109);
or U1179 (N_1179,In_77,In_219);
nor U1180 (N_1180,In_843,In_383);
nand U1181 (N_1181,In_628,In_921);
nor U1182 (N_1182,In_117,In_91);
nand U1183 (N_1183,In_549,In_630);
and U1184 (N_1184,In_707,In_727);
nor U1185 (N_1185,In_942,In_694);
or U1186 (N_1186,In_382,In_568);
or U1187 (N_1187,In_633,In_580);
or U1188 (N_1188,In_944,In_194);
or U1189 (N_1189,In_622,In_730);
and U1190 (N_1190,In_247,In_146);
nor U1191 (N_1191,In_47,In_778);
nand U1192 (N_1192,In_5,In_226);
nor U1193 (N_1193,In_489,In_679);
or U1194 (N_1194,In_685,In_519);
and U1195 (N_1195,In_824,In_674);
or U1196 (N_1196,In_452,In_569);
and U1197 (N_1197,In_450,In_812);
or U1198 (N_1198,In_653,In_194);
nand U1199 (N_1199,In_836,In_849);
nand U1200 (N_1200,In_49,In_819);
nor U1201 (N_1201,In_528,In_998);
and U1202 (N_1202,In_736,In_541);
nor U1203 (N_1203,In_592,In_215);
and U1204 (N_1204,In_538,In_877);
nor U1205 (N_1205,In_572,In_359);
or U1206 (N_1206,In_824,In_603);
nor U1207 (N_1207,In_331,In_40);
nand U1208 (N_1208,In_420,In_239);
nor U1209 (N_1209,In_371,In_261);
nor U1210 (N_1210,In_475,In_382);
or U1211 (N_1211,In_786,In_112);
or U1212 (N_1212,In_933,In_239);
and U1213 (N_1213,In_293,In_852);
nand U1214 (N_1214,In_761,In_479);
and U1215 (N_1215,In_602,In_278);
nand U1216 (N_1216,In_952,In_984);
or U1217 (N_1217,In_664,In_292);
or U1218 (N_1218,In_22,In_54);
or U1219 (N_1219,In_991,In_93);
or U1220 (N_1220,In_13,In_56);
and U1221 (N_1221,In_6,In_253);
nand U1222 (N_1222,In_898,In_35);
or U1223 (N_1223,In_799,In_291);
nand U1224 (N_1224,In_680,In_895);
and U1225 (N_1225,In_699,In_322);
and U1226 (N_1226,In_74,In_467);
and U1227 (N_1227,In_610,In_520);
or U1228 (N_1228,In_857,In_595);
or U1229 (N_1229,In_220,In_198);
or U1230 (N_1230,In_652,In_512);
or U1231 (N_1231,In_137,In_110);
or U1232 (N_1232,In_726,In_124);
nor U1233 (N_1233,In_671,In_704);
nand U1234 (N_1234,In_212,In_217);
or U1235 (N_1235,In_768,In_449);
or U1236 (N_1236,In_252,In_602);
and U1237 (N_1237,In_552,In_907);
or U1238 (N_1238,In_167,In_839);
or U1239 (N_1239,In_410,In_963);
nand U1240 (N_1240,In_168,In_778);
nand U1241 (N_1241,In_935,In_52);
or U1242 (N_1242,In_223,In_243);
nand U1243 (N_1243,In_43,In_371);
xnor U1244 (N_1244,In_728,In_422);
and U1245 (N_1245,In_220,In_68);
nand U1246 (N_1246,In_74,In_906);
or U1247 (N_1247,In_362,In_172);
nand U1248 (N_1248,In_210,In_376);
or U1249 (N_1249,In_974,In_815);
nor U1250 (N_1250,In_463,In_576);
nor U1251 (N_1251,In_974,In_669);
nand U1252 (N_1252,In_73,In_553);
nor U1253 (N_1253,In_826,In_296);
and U1254 (N_1254,In_684,In_280);
nor U1255 (N_1255,In_224,In_349);
nand U1256 (N_1256,In_550,In_36);
and U1257 (N_1257,In_295,In_487);
and U1258 (N_1258,In_711,In_192);
and U1259 (N_1259,In_345,In_71);
or U1260 (N_1260,In_953,In_162);
or U1261 (N_1261,In_151,In_283);
nand U1262 (N_1262,In_54,In_861);
nand U1263 (N_1263,In_476,In_123);
and U1264 (N_1264,In_90,In_873);
nand U1265 (N_1265,In_593,In_449);
or U1266 (N_1266,In_170,In_387);
nand U1267 (N_1267,In_393,In_517);
nand U1268 (N_1268,In_999,In_896);
or U1269 (N_1269,In_674,In_965);
and U1270 (N_1270,In_960,In_484);
and U1271 (N_1271,In_559,In_187);
nand U1272 (N_1272,In_363,In_325);
and U1273 (N_1273,In_72,In_589);
nor U1274 (N_1274,In_403,In_988);
nand U1275 (N_1275,In_561,In_243);
nand U1276 (N_1276,In_987,In_380);
and U1277 (N_1277,In_887,In_185);
nor U1278 (N_1278,In_450,In_220);
or U1279 (N_1279,In_936,In_445);
nand U1280 (N_1280,In_289,In_772);
and U1281 (N_1281,In_393,In_898);
and U1282 (N_1282,In_863,In_11);
and U1283 (N_1283,In_436,In_976);
or U1284 (N_1284,In_797,In_549);
nor U1285 (N_1285,In_432,In_552);
nor U1286 (N_1286,In_563,In_59);
nand U1287 (N_1287,In_524,In_853);
and U1288 (N_1288,In_104,In_52);
nor U1289 (N_1289,In_983,In_154);
or U1290 (N_1290,In_449,In_222);
nor U1291 (N_1291,In_864,In_827);
nand U1292 (N_1292,In_908,In_760);
nor U1293 (N_1293,In_223,In_39);
and U1294 (N_1294,In_911,In_592);
or U1295 (N_1295,In_978,In_916);
nor U1296 (N_1296,In_636,In_742);
or U1297 (N_1297,In_810,In_566);
nor U1298 (N_1298,In_395,In_663);
nand U1299 (N_1299,In_535,In_451);
nand U1300 (N_1300,In_13,In_162);
or U1301 (N_1301,In_840,In_500);
nand U1302 (N_1302,In_855,In_148);
nand U1303 (N_1303,In_575,In_682);
nor U1304 (N_1304,In_574,In_648);
nand U1305 (N_1305,In_988,In_309);
nand U1306 (N_1306,In_663,In_714);
nand U1307 (N_1307,In_295,In_195);
and U1308 (N_1308,In_550,In_597);
and U1309 (N_1309,In_902,In_507);
and U1310 (N_1310,In_488,In_683);
and U1311 (N_1311,In_293,In_16);
or U1312 (N_1312,In_67,In_936);
and U1313 (N_1313,In_700,In_485);
nand U1314 (N_1314,In_344,In_75);
nor U1315 (N_1315,In_902,In_487);
nand U1316 (N_1316,In_194,In_33);
and U1317 (N_1317,In_331,In_559);
or U1318 (N_1318,In_651,In_405);
nand U1319 (N_1319,In_998,In_842);
or U1320 (N_1320,In_480,In_651);
or U1321 (N_1321,In_486,In_639);
and U1322 (N_1322,In_977,In_684);
nor U1323 (N_1323,In_393,In_65);
xnor U1324 (N_1324,In_603,In_437);
and U1325 (N_1325,In_905,In_465);
or U1326 (N_1326,In_760,In_741);
nand U1327 (N_1327,In_792,In_709);
or U1328 (N_1328,In_249,In_533);
nor U1329 (N_1329,In_480,In_418);
and U1330 (N_1330,In_640,In_791);
nand U1331 (N_1331,In_174,In_397);
nand U1332 (N_1332,In_308,In_154);
nand U1333 (N_1333,In_545,In_325);
and U1334 (N_1334,In_981,In_512);
and U1335 (N_1335,In_734,In_937);
nand U1336 (N_1336,In_863,In_861);
and U1337 (N_1337,In_292,In_566);
and U1338 (N_1338,In_385,In_35);
and U1339 (N_1339,In_316,In_97);
and U1340 (N_1340,In_975,In_345);
nor U1341 (N_1341,In_167,In_628);
and U1342 (N_1342,In_236,In_253);
nand U1343 (N_1343,In_381,In_921);
nand U1344 (N_1344,In_203,In_544);
nor U1345 (N_1345,In_912,In_842);
and U1346 (N_1346,In_871,In_33);
nand U1347 (N_1347,In_303,In_282);
nand U1348 (N_1348,In_305,In_220);
nor U1349 (N_1349,In_660,In_338);
and U1350 (N_1350,In_283,In_257);
nand U1351 (N_1351,In_593,In_29);
or U1352 (N_1352,In_978,In_724);
and U1353 (N_1353,In_383,In_329);
and U1354 (N_1354,In_375,In_135);
and U1355 (N_1355,In_444,In_789);
nor U1356 (N_1356,In_236,In_938);
nand U1357 (N_1357,In_734,In_100);
and U1358 (N_1358,In_102,In_984);
and U1359 (N_1359,In_530,In_307);
nor U1360 (N_1360,In_529,In_224);
nor U1361 (N_1361,In_267,In_700);
and U1362 (N_1362,In_430,In_358);
or U1363 (N_1363,In_350,In_434);
and U1364 (N_1364,In_899,In_524);
and U1365 (N_1365,In_797,In_785);
nor U1366 (N_1366,In_999,In_589);
or U1367 (N_1367,In_836,In_755);
and U1368 (N_1368,In_576,In_998);
nor U1369 (N_1369,In_112,In_336);
nand U1370 (N_1370,In_258,In_954);
nor U1371 (N_1371,In_972,In_320);
or U1372 (N_1372,In_964,In_861);
and U1373 (N_1373,In_185,In_38);
and U1374 (N_1374,In_167,In_188);
or U1375 (N_1375,In_339,In_669);
or U1376 (N_1376,In_326,In_589);
and U1377 (N_1377,In_636,In_473);
or U1378 (N_1378,In_607,In_134);
and U1379 (N_1379,In_973,In_181);
nor U1380 (N_1380,In_168,In_364);
nand U1381 (N_1381,In_803,In_450);
nor U1382 (N_1382,In_653,In_120);
nand U1383 (N_1383,In_731,In_267);
and U1384 (N_1384,In_682,In_724);
nand U1385 (N_1385,In_481,In_413);
nand U1386 (N_1386,In_460,In_810);
nand U1387 (N_1387,In_624,In_1);
nor U1388 (N_1388,In_431,In_797);
nor U1389 (N_1389,In_607,In_817);
nand U1390 (N_1390,In_853,In_806);
nor U1391 (N_1391,In_514,In_472);
nand U1392 (N_1392,In_199,In_633);
and U1393 (N_1393,In_296,In_637);
nor U1394 (N_1394,In_222,In_848);
or U1395 (N_1395,In_145,In_433);
nor U1396 (N_1396,In_454,In_148);
or U1397 (N_1397,In_741,In_257);
nand U1398 (N_1398,In_667,In_823);
or U1399 (N_1399,In_951,In_412);
nor U1400 (N_1400,In_628,In_332);
nor U1401 (N_1401,In_255,In_859);
nor U1402 (N_1402,In_565,In_332);
nand U1403 (N_1403,In_680,In_604);
nand U1404 (N_1404,In_854,In_841);
nand U1405 (N_1405,In_568,In_415);
or U1406 (N_1406,In_619,In_49);
nor U1407 (N_1407,In_13,In_181);
nand U1408 (N_1408,In_651,In_525);
nand U1409 (N_1409,In_963,In_183);
or U1410 (N_1410,In_624,In_994);
or U1411 (N_1411,In_303,In_153);
nand U1412 (N_1412,In_79,In_973);
nand U1413 (N_1413,In_903,In_176);
or U1414 (N_1414,In_876,In_198);
and U1415 (N_1415,In_39,In_698);
or U1416 (N_1416,In_647,In_454);
nor U1417 (N_1417,In_759,In_620);
or U1418 (N_1418,In_52,In_534);
nand U1419 (N_1419,In_182,In_681);
nand U1420 (N_1420,In_733,In_15);
or U1421 (N_1421,In_645,In_530);
nand U1422 (N_1422,In_14,In_786);
nand U1423 (N_1423,In_657,In_162);
and U1424 (N_1424,In_134,In_253);
nand U1425 (N_1425,In_374,In_660);
or U1426 (N_1426,In_284,In_803);
nor U1427 (N_1427,In_959,In_965);
nand U1428 (N_1428,In_271,In_21);
or U1429 (N_1429,In_608,In_921);
nand U1430 (N_1430,In_305,In_756);
xnor U1431 (N_1431,In_115,In_565);
and U1432 (N_1432,In_818,In_100);
nor U1433 (N_1433,In_92,In_950);
or U1434 (N_1434,In_54,In_160);
nor U1435 (N_1435,In_113,In_283);
or U1436 (N_1436,In_371,In_937);
nor U1437 (N_1437,In_396,In_359);
or U1438 (N_1438,In_44,In_774);
nand U1439 (N_1439,In_356,In_602);
nor U1440 (N_1440,In_66,In_863);
nor U1441 (N_1441,In_487,In_570);
or U1442 (N_1442,In_338,In_405);
nor U1443 (N_1443,In_338,In_858);
nand U1444 (N_1444,In_766,In_213);
nor U1445 (N_1445,In_749,In_504);
or U1446 (N_1446,In_825,In_328);
nor U1447 (N_1447,In_207,In_33);
and U1448 (N_1448,In_732,In_455);
xnor U1449 (N_1449,In_641,In_44);
nor U1450 (N_1450,In_917,In_944);
nand U1451 (N_1451,In_965,In_979);
or U1452 (N_1452,In_414,In_975);
nor U1453 (N_1453,In_644,In_613);
and U1454 (N_1454,In_371,In_7);
nor U1455 (N_1455,In_608,In_765);
or U1456 (N_1456,In_850,In_548);
and U1457 (N_1457,In_780,In_385);
xor U1458 (N_1458,In_744,In_706);
or U1459 (N_1459,In_280,In_834);
nor U1460 (N_1460,In_23,In_849);
or U1461 (N_1461,In_440,In_750);
or U1462 (N_1462,In_368,In_78);
and U1463 (N_1463,In_901,In_71);
and U1464 (N_1464,In_319,In_61);
and U1465 (N_1465,In_181,In_249);
nor U1466 (N_1466,In_402,In_589);
nor U1467 (N_1467,In_710,In_632);
or U1468 (N_1468,In_282,In_406);
nand U1469 (N_1469,In_705,In_845);
and U1470 (N_1470,In_473,In_834);
nor U1471 (N_1471,In_150,In_522);
and U1472 (N_1472,In_109,In_715);
nand U1473 (N_1473,In_653,In_445);
or U1474 (N_1474,In_791,In_686);
and U1475 (N_1475,In_964,In_730);
nor U1476 (N_1476,In_288,In_562);
nand U1477 (N_1477,In_326,In_981);
or U1478 (N_1478,In_207,In_999);
nor U1479 (N_1479,In_650,In_200);
and U1480 (N_1480,In_732,In_650);
and U1481 (N_1481,In_327,In_555);
or U1482 (N_1482,In_931,In_724);
nand U1483 (N_1483,In_852,In_382);
nand U1484 (N_1484,In_848,In_547);
or U1485 (N_1485,In_813,In_684);
nand U1486 (N_1486,In_132,In_237);
nor U1487 (N_1487,In_529,In_547);
and U1488 (N_1488,In_709,In_46);
nand U1489 (N_1489,In_704,In_616);
or U1490 (N_1490,In_146,In_775);
nand U1491 (N_1491,In_791,In_351);
or U1492 (N_1492,In_514,In_626);
or U1493 (N_1493,In_203,In_148);
nor U1494 (N_1494,In_894,In_442);
and U1495 (N_1495,In_750,In_506);
nor U1496 (N_1496,In_30,In_904);
and U1497 (N_1497,In_904,In_106);
and U1498 (N_1498,In_541,In_321);
nor U1499 (N_1499,In_731,In_573);
nand U1500 (N_1500,In_720,In_931);
nor U1501 (N_1501,In_513,In_567);
nand U1502 (N_1502,In_753,In_94);
nand U1503 (N_1503,In_139,In_381);
nand U1504 (N_1504,In_992,In_699);
nor U1505 (N_1505,In_214,In_566);
or U1506 (N_1506,In_958,In_307);
or U1507 (N_1507,In_802,In_798);
and U1508 (N_1508,In_419,In_796);
nand U1509 (N_1509,In_687,In_150);
or U1510 (N_1510,In_582,In_588);
and U1511 (N_1511,In_469,In_81);
nor U1512 (N_1512,In_158,In_523);
and U1513 (N_1513,In_178,In_525);
nor U1514 (N_1514,In_757,In_354);
or U1515 (N_1515,In_76,In_827);
or U1516 (N_1516,In_642,In_952);
and U1517 (N_1517,In_144,In_466);
or U1518 (N_1518,In_693,In_612);
nor U1519 (N_1519,In_44,In_272);
nand U1520 (N_1520,In_635,In_223);
and U1521 (N_1521,In_885,In_440);
nor U1522 (N_1522,In_583,In_395);
or U1523 (N_1523,In_861,In_235);
or U1524 (N_1524,In_52,In_192);
nand U1525 (N_1525,In_59,In_408);
or U1526 (N_1526,In_380,In_105);
or U1527 (N_1527,In_407,In_940);
nor U1528 (N_1528,In_698,In_793);
and U1529 (N_1529,In_591,In_858);
nand U1530 (N_1530,In_262,In_54);
or U1531 (N_1531,In_52,In_923);
nand U1532 (N_1532,In_806,In_768);
and U1533 (N_1533,In_491,In_711);
or U1534 (N_1534,In_453,In_651);
nor U1535 (N_1535,In_822,In_251);
and U1536 (N_1536,In_998,In_668);
nor U1537 (N_1537,In_460,In_545);
and U1538 (N_1538,In_793,In_118);
or U1539 (N_1539,In_782,In_43);
or U1540 (N_1540,In_613,In_761);
nor U1541 (N_1541,In_257,In_61);
and U1542 (N_1542,In_530,In_971);
and U1543 (N_1543,In_146,In_259);
and U1544 (N_1544,In_301,In_828);
nand U1545 (N_1545,In_753,In_969);
or U1546 (N_1546,In_37,In_369);
nor U1547 (N_1547,In_20,In_967);
nand U1548 (N_1548,In_47,In_562);
nand U1549 (N_1549,In_435,In_293);
or U1550 (N_1550,In_903,In_153);
nor U1551 (N_1551,In_836,In_466);
nor U1552 (N_1552,In_111,In_911);
or U1553 (N_1553,In_419,In_484);
nor U1554 (N_1554,In_772,In_737);
nor U1555 (N_1555,In_361,In_199);
nand U1556 (N_1556,In_120,In_708);
or U1557 (N_1557,In_333,In_737);
and U1558 (N_1558,In_42,In_187);
nand U1559 (N_1559,In_311,In_459);
nor U1560 (N_1560,In_598,In_659);
and U1561 (N_1561,In_934,In_307);
or U1562 (N_1562,In_586,In_481);
or U1563 (N_1563,In_542,In_662);
or U1564 (N_1564,In_586,In_531);
and U1565 (N_1565,In_928,In_595);
nand U1566 (N_1566,In_898,In_244);
and U1567 (N_1567,In_86,In_459);
or U1568 (N_1568,In_97,In_27);
and U1569 (N_1569,In_845,In_756);
nor U1570 (N_1570,In_459,In_221);
and U1571 (N_1571,In_821,In_770);
or U1572 (N_1572,In_22,In_17);
nand U1573 (N_1573,In_110,In_391);
nor U1574 (N_1574,In_246,In_181);
nor U1575 (N_1575,In_51,In_36);
nand U1576 (N_1576,In_600,In_663);
or U1577 (N_1577,In_739,In_764);
or U1578 (N_1578,In_927,In_589);
and U1579 (N_1579,In_581,In_337);
and U1580 (N_1580,In_161,In_891);
nor U1581 (N_1581,In_458,In_106);
or U1582 (N_1582,In_385,In_563);
or U1583 (N_1583,In_964,In_578);
nor U1584 (N_1584,In_755,In_49);
or U1585 (N_1585,In_18,In_483);
nand U1586 (N_1586,In_363,In_824);
or U1587 (N_1587,In_123,In_5);
nand U1588 (N_1588,In_473,In_94);
nand U1589 (N_1589,In_188,In_429);
or U1590 (N_1590,In_909,In_855);
and U1591 (N_1591,In_192,In_60);
nand U1592 (N_1592,In_609,In_727);
or U1593 (N_1593,In_46,In_447);
or U1594 (N_1594,In_838,In_584);
nand U1595 (N_1595,In_740,In_92);
nor U1596 (N_1596,In_184,In_741);
or U1597 (N_1597,In_124,In_859);
and U1598 (N_1598,In_216,In_940);
nand U1599 (N_1599,In_555,In_875);
nand U1600 (N_1600,In_853,In_78);
nand U1601 (N_1601,In_88,In_798);
nor U1602 (N_1602,In_124,In_492);
and U1603 (N_1603,In_68,In_728);
and U1604 (N_1604,In_44,In_301);
or U1605 (N_1605,In_171,In_426);
or U1606 (N_1606,In_778,In_863);
and U1607 (N_1607,In_996,In_836);
nor U1608 (N_1608,In_575,In_958);
nor U1609 (N_1609,In_34,In_142);
nand U1610 (N_1610,In_588,In_256);
or U1611 (N_1611,In_72,In_650);
and U1612 (N_1612,In_369,In_627);
nor U1613 (N_1613,In_491,In_978);
and U1614 (N_1614,In_231,In_93);
or U1615 (N_1615,In_116,In_916);
and U1616 (N_1616,In_501,In_52);
nand U1617 (N_1617,In_492,In_980);
and U1618 (N_1618,In_443,In_175);
and U1619 (N_1619,In_381,In_510);
nand U1620 (N_1620,In_488,In_518);
and U1621 (N_1621,In_173,In_153);
and U1622 (N_1622,In_485,In_713);
and U1623 (N_1623,In_249,In_347);
nand U1624 (N_1624,In_735,In_710);
and U1625 (N_1625,In_248,In_780);
nor U1626 (N_1626,In_447,In_242);
or U1627 (N_1627,In_697,In_767);
nor U1628 (N_1628,In_42,In_5);
nand U1629 (N_1629,In_269,In_419);
or U1630 (N_1630,In_9,In_168);
or U1631 (N_1631,In_825,In_956);
nor U1632 (N_1632,In_875,In_827);
nor U1633 (N_1633,In_104,In_856);
nand U1634 (N_1634,In_408,In_346);
and U1635 (N_1635,In_130,In_68);
or U1636 (N_1636,In_27,In_446);
and U1637 (N_1637,In_673,In_698);
or U1638 (N_1638,In_273,In_831);
nor U1639 (N_1639,In_194,In_482);
nor U1640 (N_1640,In_179,In_24);
or U1641 (N_1641,In_550,In_86);
and U1642 (N_1642,In_679,In_664);
nor U1643 (N_1643,In_296,In_507);
xor U1644 (N_1644,In_633,In_725);
nor U1645 (N_1645,In_517,In_716);
and U1646 (N_1646,In_851,In_676);
nand U1647 (N_1647,In_506,In_125);
nor U1648 (N_1648,In_364,In_631);
nand U1649 (N_1649,In_770,In_478);
and U1650 (N_1650,In_635,In_800);
xnor U1651 (N_1651,In_831,In_18);
nor U1652 (N_1652,In_347,In_165);
nand U1653 (N_1653,In_615,In_852);
nand U1654 (N_1654,In_623,In_275);
nand U1655 (N_1655,In_773,In_494);
nand U1656 (N_1656,In_11,In_55);
nor U1657 (N_1657,In_595,In_441);
nor U1658 (N_1658,In_996,In_596);
nor U1659 (N_1659,In_224,In_193);
and U1660 (N_1660,In_254,In_88);
nand U1661 (N_1661,In_286,In_607);
nor U1662 (N_1662,In_364,In_320);
or U1663 (N_1663,In_402,In_759);
nor U1664 (N_1664,In_115,In_712);
nand U1665 (N_1665,In_465,In_776);
nor U1666 (N_1666,In_482,In_595);
and U1667 (N_1667,In_714,In_830);
or U1668 (N_1668,In_30,In_294);
nor U1669 (N_1669,In_828,In_421);
nand U1670 (N_1670,In_790,In_112);
or U1671 (N_1671,In_615,In_47);
nand U1672 (N_1672,In_174,In_686);
nor U1673 (N_1673,In_454,In_545);
nor U1674 (N_1674,In_652,In_927);
nor U1675 (N_1675,In_134,In_559);
or U1676 (N_1676,In_804,In_79);
nor U1677 (N_1677,In_400,In_525);
and U1678 (N_1678,In_972,In_501);
nand U1679 (N_1679,In_441,In_119);
nor U1680 (N_1680,In_490,In_180);
or U1681 (N_1681,In_801,In_946);
nand U1682 (N_1682,In_93,In_272);
or U1683 (N_1683,In_439,In_65);
nand U1684 (N_1684,In_314,In_228);
or U1685 (N_1685,In_123,In_697);
nor U1686 (N_1686,In_521,In_752);
and U1687 (N_1687,In_941,In_545);
nand U1688 (N_1688,In_501,In_281);
and U1689 (N_1689,In_56,In_361);
and U1690 (N_1690,In_172,In_1);
and U1691 (N_1691,In_756,In_742);
and U1692 (N_1692,In_970,In_260);
or U1693 (N_1693,In_746,In_927);
and U1694 (N_1694,In_866,In_637);
nand U1695 (N_1695,In_132,In_6);
and U1696 (N_1696,In_750,In_83);
nor U1697 (N_1697,In_162,In_955);
and U1698 (N_1698,In_631,In_885);
nor U1699 (N_1699,In_943,In_448);
nor U1700 (N_1700,In_430,In_139);
nor U1701 (N_1701,In_374,In_591);
xor U1702 (N_1702,In_284,In_246);
nor U1703 (N_1703,In_663,In_611);
nor U1704 (N_1704,In_428,In_157);
and U1705 (N_1705,In_971,In_569);
or U1706 (N_1706,In_145,In_812);
or U1707 (N_1707,In_997,In_345);
and U1708 (N_1708,In_75,In_880);
nor U1709 (N_1709,In_136,In_918);
and U1710 (N_1710,In_231,In_482);
and U1711 (N_1711,In_811,In_270);
and U1712 (N_1712,In_232,In_903);
and U1713 (N_1713,In_689,In_682);
nand U1714 (N_1714,In_302,In_733);
and U1715 (N_1715,In_229,In_703);
and U1716 (N_1716,In_268,In_217);
or U1717 (N_1717,In_704,In_840);
nand U1718 (N_1718,In_18,In_528);
or U1719 (N_1719,In_394,In_23);
nand U1720 (N_1720,In_61,In_32);
or U1721 (N_1721,In_972,In_879);
and U1722 (N_1722,In_560,In_552);
nor U1723 (N_1723,In_123,In_738);
nand U1724 (N_1724,In_680,In_573);
nor U1725 (N_1725,In_773,In_838);
nand U1726 (N_1726,In_470,In_778);
or U1727 (N_1727,In_607,In_739);
nor U1728 (N_1728,In_801,In_268);
nor U1729 (N_1729,In_13,In_245);
or U1730 (N_1730,In_866,In_171);
and U1731 (N_1731,In_874,In_789);
nand U1732 (N_1732,In_960,In_635);
and U1733 (N_1733,In_896,In_279);
nand U1734 (N_1734,In_236,In_546);
nor U1735 (N_1735,In_384,In_277);
and U1736 (N_1736,In_822,In_30);
or U1737 (N_1737,In_109,In_307);
and U1738 (N_1738,In_596,In_763);
nor U1739 (N_1739,In_228,In_275);
or U1740 (N_1740,In_182,In_66);
or U1741 (N_1741,In_253,In_648);
and U1742 (N_1742,In_749,In_788);
and U1743 (N_1743,In_802,In_441);
nand U1744 (N_1744,In_485,In_806);
and U1745 (N_1745,In_272,In_256);
or U1746 (N_1746,In_455,In_163);
nand U1747 (N_1747,In_174,In_725);
nand U1748 (N_1748,In_509,In_365);
and U1749 (N_1749,In_537,In_739);
nand U1750 (N_1750,In_408,In_283);
nor U1751 (N_1751,In_212,In_171);
nand U1752 (N_1752,In_124,In_531);
and U1753 (N_1753,In_933,In_906);
or U1754 (N_1754,In_890,In_89);
nor U1755 (N_1755,In_7,In_536);
nor U1756 (N_1756,In_674,In_490);
nand U1757 (N_1757,In_716,In_977);
and U1758 (N_1758,In_634,In_826);
or U1759 (N_1759,In_763,In_445);
nand U1760 (N_1760,In_720,In_485);
nor U1761 (N_1761,In_263,In_550);
nand U1762 (N_1762,In_880,In_681);
and U1763 (N_1763,In_13,In_678);
nand U1764 (N_1764,In_975,In_139);
or U1765 (N_1765,In_429,In_222);
nand U1766 (N_1766,In_346,In_405);
nand U1767 (N_1767,In_743,In_730);
nand U1768 (N_1768,In_786,In_290);
xnor U1769 (N_1769,In_581,In_748);
nand U1770 (N_1770,In_264,In_66);
xor U1771 (N_1771,In_709,In_992);
nor U1772 (N_1772,In_406,In_155);
nor U1773 (N_1773,In_713,In_629);
or U1774 (N_1774,In_280,In_822);
or U1775 (N_1775,In_324,In_430);
and U1776 (N_1776,In_261,In_217);
nor U1777 (N_1777,In_464,In_115);
or U1778 (N_1778,In_21,In_397);
or U1779 (N_1779,In_881,In_554);
or U1780 (N_1780,In_871,In_737);
or U1781 (N_1781,In_331,In_164);
and U1782 (N_1782,In_931,In_815);
nor U1783 (N_1783,In_656,In_700);
and U1784 (N_1784,In_996,In_955);
nand U1785 (N_1785,In_832,In_989);
or U1786 (N_1786,In_125,In_884);
nand U1787 (N_1787,In_837,In_677);
nor U1788 (N_1788,In_110,In_50);
and U1789 (N_1789,In_213,In_637);
xnor U1790 (N_1790,In_915,In_528);
nor U1791 (N_1791,In_672,In_20);
nor U1792 (N_1792,In_836,In_769);
or U1793 (N_1793,In_509,In_919);
nand U1794 (N_1794,In_803,In_748);
nand U1795 (N_1795,In_11,In_722);
or U1796 (N_1796,In_93,In_123);
or U1797 (N_1797,In_589,In_980);
or U1798 (N_1798,In_592,In_653);
and U1799 (N_1799,In_686,In_719);
and U1800 (N_1800,In_847,In_221);
nor U1801 (N_1801,In_724,In_853);
nor U1802 (N_1802,In_701,In_304);
nor U1803 (N_1803,In_977,In_535);
and U1804 (N_1804,In_937,In_879);
nand U1805 (N_1805,In_390,In_262);
and U1806 (N_1806,In_499,In_408);
or U1807 (N_1807,In_393,In_743);
or U1808 (N_1808,In_76,In_41);
or U1809 (N_1809,In_708,In_774);
or U1810 (N_1810,In_818,In_798);
nor U1811 (N_1811,In_999,In_904);
and U1812 (N_1812,In_563,In_372);
nor U1813 (N_1813,In_884,In_565);
nand U1814 (N_1814,In_846,In_451);
and U1815 (N_1815,In_612,In_400);
and U1816 (N_1816,In_149,In_386);
nor U1817 (N_1817,In_828,In_694);
or U1818 (N_1818,In_114,In_499);
nor U1819 (N_1819,In_778,In_344);
or U1820 (N_1820,In_171,In_654);
nor U1821 (N_1821,In_260,In_683);
nand U1822 (N_1822,In_356,In_934);
nand U1823 (N_1823,In_561,In_733);
nor U1824 (N_1824,In_799,In_483);
nor U1825 (N_1825,In_236,In_734);
nand U1826 (N_1826,In_219,In_13);
nand U1827 (N_1827,In_361,In_28);
nand U1828 (N_1828,In_311,In_899);
nand U1829 (N_1829,In_376,In_589);
nand U1830 (N_1830,In_258,In_158);
nand U1831 (N_1831,In_3,In_889);
nand U1832 (N_1832,In_541,In_83);
nand U1833 (N_1833,In_273,In_121);
or U1834 (N_1834,In_988,In_935);
and U1835 (N_1835,In_83,In_228);
nor U1836 (N_1836,In_312,In_173);
or U1837 (N_1837,In_298,In_56);
nor U1838 (N_1838,In_184,In_882);
and U1839 (N_1839,In_921,In_709);
or U1840 (N_1840,In_367,In_359);
or U1841 (N_1841,In_617,In_194);
nand U1842 (N_1842,In_23,In_864);
and U1843 (N_1843,In_822,In_405);
and U1844 (N_1844,In_573,In_20);
and U1845 (N_1845,In_152,In_446);
or U1846 (N_1846,In_8,In_743);
or U1847 (N_1847,In_923,In_806);
or U1848 (N_1848,In_379,In_938);
or U1849 (N_1849,In_543,In_766);
and U1850 (N_1850,In_207,In_110);
nor U1851 (N_1851,In_117,In_582);
nor U1852 (N_1852,In_630,In_791);
nand U1853 (N_1853,In_674,In_461);
nand U1854 (N_1854,In_600,In_766);
and U1855 (N_1855,In_72,In_995);
and U1856 (N_1856,In_240,In_925);
nor U1857 (N_1857,In_609,In_694);
or U1858 (N_1858,In_893,In_228);
and U1859 (N_1859,In_357,In_137);
nor U1860 (N_1860,In_310,In_766);
and U1861 (N_1861,In_854,In_141);
nand U1862 (N_1862,In_471,In_345);
nand U1863 (N_1863,In_422,In_197);
nor U1864 (N_1864,In_840,In_751);
nor U1865 (N_1865,In_396,In_516);
nand U1866 (N_1866,In_563,In_754);
nor U1867 (N_1867,In_160,In_172);
or U1868 (N_1868,In_290,In_756);
nor U1869 (N_1869,In_168,In_183);
nand U1870 (N_1870,In_964,In_51);
or U1871 (N_1871,In_174,In_180);
nor U1872 (N_1872,In_449,In_353);
and U1873 (N_1873,In_670,In_641);
or U1874 (N_1874,In_371,In_365);
and U1875 (N_1875,In_374,In_955);
and U1876 (N_1876,In_604,In_990);
or U1877 (N_1877,In_319,In_619);
nand U1878 (N_1878,In_96,In_721);
nor U1879 (N_1879,In_969,In_70);
and U1880 (N_1880,In_731,In_747);
and U1881 (N_1881,In_658,In_731);
nand U1882 (N_1882,In_281,In_892);
and U1883 (N_1883,In_855,In_792);
nor U1884 (N_1884,In_99,In_19);
or U1885 (N_1885,In_742,In_892);
and U1886 (N_1886,In_539,In_900);
and U1887 (N_1887,In_944,In_588);
nand U1888 (N_1888,In_985,In_818);
and U1889 (N_1889,In_693,In_861);
and U1890 (N_1890,In_704,In_64);
and U1891 (N_1891,In_734,In_903);
nor U1892 (N_1892,In_405,In_143);
nand U1893 (N_1893,In_850,In_702);
nand U1894 (N_1894,In_666,In_264);
nand U1895 (N_1895,In_805,In_816);
and U1896 (N_1896,In_228,In_261);
or U1897 (N_1897,In_607,In_790);
and U1898 (N_1898,In_976,In_666);
nor U1899 (N_1899,In_712,In_321);
nand U1900 (N_1900,In_558,In_342);
nand U1901 (N_1901,In_52,In_616);
nor U1902 (N_1902,In_350,In_899);
nor U1903 (N_1903,In_646,In_907);
and U1904 (N_1904,In_668,In_566);
nor U1905 (N_1905,In_262,In_555);
nor U1906 (N_1906,In_0,In_748);
or U1907 (N_1907,In_127,In_544);
and U1908 (N_1908,In_109,In_261);
and U1909 (N_1909,In_71,In_792);
nor U1910 (N_1910,In_472,In_256);
nor U1911 (N_1911,In_227,In_849);
nand U1912 (N_1912,In_994,In_936);
or U1913 (N_1913,In_475,In_781);
and U1914 (N_1914,In_663,In_936);
nand U1915 (N_1915,In_135,In_955);
and U1916 (N_1916,In_764,In_855);
nand U1917 (N_1917,In_560,In_352);
or U1918 (N_1918,In_308,In_819);
xor U1919 (N_1919,In_664,In_52);
nand U1920 (N_1920,In_776,In_401);
or U1921 (N_1921,In_429,In_908);
and U1922 (N_1922,In_762,In_800);
nand U1923 (N_1923,In_256,In_226);
nor U1924 (N_1924,In_194,In_517);
nand U1925 (N_1925,In_363,In_690);
or U1926 (N_1926,In_275,In_779);
nand U1927 (N_1927,In_3,In_0);
or U1928 (N_1928,In_598,In_133);
nand U1929 (N_1929,In_388,In_986);
or U1930 (N_1930,In_96,In_257);
nor U1931 (N_1931,In_430,In_45);
nand U1932 (N_1932,In_802,In_59);
nor U1933 (N_1933,In_932,In_363);
nand U1934 (N_1934,In_983,In_988);
or U1935 (N_1935,In_11,In_470);
nor U1936 (N_1936,In_925,In_916);
nor U1937 (N_1937,In_651,In_153);
nand U1938 (N_1938,In_401,In_980);
nand U1939 (N_1939,In_620,In_652);
and U1940 (N_1940,In_420,In_616);
nor U1941 (N_1941,In_222,In_470);
nand U1942 (N_1942,In_386,In_749);
and U1943 (N_1943,In_286,In_587);
and U1944 (N_1944,In_480,In_586);
xnor U1945 (N_1945,In_14,In_931);
or U1946 (N_1946,In_645,In_869);
nand U1947 (N_1947,In_915,In_287);
or U1948 (N_1948,In_523,In_864);
nor U1949 (N_1949,In_967,In_993);
and U1950 (N_1950,In_404,In_299);
and U1951 (N_1951,In_499,In_376);
and U1952 (N_1952,In_859,In_288);
or U1953 (N_1953,In_104,In_365);
nand U1954 (N_1954,In_378,In_766);
nand U1955 (N_1955,In_6,In_144);
or U1956 (N_1956,In_355,In_774);
and U1957 (N_1957,In_788,In_952);
or U1958 (N_1958,In_734,In_702);
and U1959 (N_1959,In_354,In_781);
and U1960 (N_1960,In_995,In_552);
or U1961 (N_1961,In_42,In_961);
nor U1962 (N_1962,In_13,In_573);
nand U1963 (N_1963,In_33,In_658);
or U1964 (N_1964,In_747,In_491);
or U1965 (N_1965,In_374,In_141);
and U1966 (N_1966,In_32,In_156);
and U1967 (N_1967,In_646,In_12);
or U1968 (N_1968,In_942,In_862);
or U1969 (N_1969,In_999,In_128);
and U1970 (N_1970,In_847,In_514);
or U1971 (N_1971,In_232,In_363);
and U1972 (N_1972,In_418,In_324);
and U1973 (N_1973,In_326,In_397);
and U1974 (N_1974,In_72,In_478);
nor U1975 (N_1975,In_664,In_131);
nand U1976 (N_1976,In_548,In_986);
nand U1977 (N_1977,In_949,In_26);
or U1978 (N_1978,In_15,In_323);
nor U1979 (N_1979,In_607,In_369);
and U1980 (N_1980,In_637,In_422);
and U1981 (N_1981,In_681,In_506);
nand U1982 (N_1982,In_223,In_830);
nand U1983 (N_1983,In_291,In_30);
nor U1984 (N_1984,In_687,In_600);
nor U1985 (N_1985,In_940,In_571);
nand U1986 (N_1986,In_886,In_929);
nand U1987 (N_1987,In_310,In_442);
nor U1988 (N_1988,In_845,In_483);
or U1989 (N_1989,In_981,In_686);
and U1990 (N_1990,In_999,In_922);
nor U1991 (N_1991,In_80,In_902);
and U1992 (N_1992,In_89,In_345);
or U1993 (N_1993,In_729,In_319);
nand U1994 (N_1994,In_0,In_704);
or U1995 (N_1995,In_541,In_530);
nor U1996 (N_1996,In_127,In_276);
nand U1997 (N_1997,In_61,In_233);
nor U1998 (N_1998,In_642,In_46);
nor U1999 (N_1999,In_878,In_975);
nor U2000 (N_2000,In_796,In_10);
nor U2001 (N_2001,In_821,In_287);
nor U2002 (N_2002,In_407,In_197);
or U2003 (N_2003,In_911,In_824);
nor U2004 (N_2004,In_822,In_596);
nand U2005 (N_2005,In_269,In_167);
or U2006 (N_2006,In_147,In_516);
and U2007 (N_2007,In_611,In_496);
or U2008 (N_2008,In_322,In_677);
or U2009 (N_2009,In_356,In_873);
nor U2010 (N_2010,In_457,In_772);
nand U2011 (N_2011,In_326,In_482);
nand U2012 (N_2012,In_915,In_452);
nand U2013 (N_2013,In_849,In_384);
nor U2014 (N_2014,In_103,In_79);
and U2015 (N_2015,In_562,In_739);
nand U2016 (N_2016,In_442,In_728);
or U2017 (N_2017,In_447,In_290);
nand U2018 (N_2018,In_309,In_996);
nor U2019 (N_2019,In_263,In_523);
and U2020 (N_2020,In_403,In_230);
nand U2021 (N_2021,In_614,In_252);
and U2022 (N_2022,In_779,In_345);
nor U2023 (N_2023,In_465,In_104);
or U2024 (N_2024,In_418,In_777);
nand U2025 (N_2025,In_574,In_544);
or U2026 (N_2026,In_487,In_933);
and U2027 (N_2027,In_63,In_461);
or U2028 (N_2028,In_301,In_214);
and U2029 (N_2029,In_113,In_996);
or U2030 (N_2030,In_828,In_463);
or U2031 (N_2031,In_324,In_440);
nand U2032 (N_2032,In_878,In_52);
nor U2033 (N_2033,In_697,In_336);
nor U2034 (N_2034,In_631,In_21);
and U2035 (N_2035,In_236,In_972);
nor U2036 (N_2036,In_392,In_445);
and U2037 (N_2037,In_545,In_44);
or U2038 (N_2038,In_425,In_342);
or U2039 (N_2039,In_529,In_680);
nand U2040 (N_2040,In_949,In_53);
nor U2041 (N_2041,In_364,In_672);
or U2042 (N_2042,In_8,In_121);
and U2043 (N_2043,In_214,In_186);
or U2044 (N_2044,In_935,In_514);
nand U2045 (N_2045,In_601,In_401);
nand U2046 (N_2046,In_502,In_850);
nor U2047 (N_2047,In_598,In_712);
nor U2048 (N_2048,In_535,In_745);
nor U2049 (N_2049,In_347,In_101);
nand U2050 (N_2050,In_703,In_950);
or U2051 (N_2051,In_403,In_253);
nand U2052 (N_2052,In_837,In_599);
nor U2053 (N_2053,In_350,In_9);
or U2054 (N_2054,In_395,In_236);
nand U2055 (N_2055,In_846,In_734);
or U2056 (N_2056,In_106,In_395);
and U2057 (N_2057,In_550,In_843);
or U2058 (N_2058,In_972,In_51);
or U2059 (N_2059,In_929,In_139);
and U2060 (N_2060,In_975,In_624);
nand U2061 (N_2061,In_783,In_116);
nand U2062 (N_2062,In_998,In_763);
and U2063 (N_2063,In_286,In_343);
or U2064 (N_2064,In_967,In_411);
or U2065 (N_2065,In_734,In_139);
nor U2066 (N_2066,In_879,In_609);
nor U2067 (N_2067,In_352,In_562);
nand U2068 (N_2068,In_797,In_193);
nand U2069 (N_2069,In_103,In_782);
nand U2070 (N_2070,In_843,In_992);
or U2071 (N_2071,In_836,In_973);
or U2072 (N_2072,In_185,In_513);
nand U2073 (N_2073,In_761,In_252);
and U2074 (N_2074,In_388,In_677);
or U2075 (N_2075,In_130,In_853);
nand U2076 (N_2076,In_813,In_858);
nand U2077 (N_2077,In_514,In_249);
nor U2078 (N_2078,In_360,In_136);
nor U2079 (N_2079,In_581,In_749);
nand U2080 (N_2080,In_376,In_103);
nand U2081 (N_2081,In_619,In_206);
nand U2082 (N_2082,In_702,In_912);
nor U2083 (N_2083,In_858,In_662);
or U2084 (N_2084,In_75,In_532);
nor U2085 (N_2085,In_672,In_67);
or U2086 (N_2086,In_280,In_605);
and U2087 (N_2087,In_910,In_477);
nor U2088 (N_2088,In_212,In_719);
and U2089 (N_2089,In_906,In_629);
nand U2090 (N_2090,In_170,In_81);
or U2091 (N_2091,In_565,In_455);
nand U2092 (N_2092,In_230,In_978);
and U2093 (N_2093,In_276,In_123);
nand U2094 (N_2094,In_281,In_595);
and U2095 (N_2095,In_395,In_397);
nor U2096 (N_2096,In_208,In_441);
nand U2097 (N_2097,In_475,In_958);
nand U2098 (N_2098,In_611,In_917);
and U2099 (N_2099,In_948,In_351);
and U2100 (N_2100,In_178,In_588);
nor U2101 (N_2101,In_948,In_707);
nand U2102 (N_2102,In_916,In_503);
and U2103 (N_2103,In_283,In_832);
and U2104 (N_2104,In_962,In_993);
xor U2105 (N_2105,In_101,In_946);
and U2106 (N_2106,In_543,In_262);
nand U2107 (N_2107,In_797,In_994);
nor U2108 (N_2108,In_13,In_604);
nand U2109 (N_2109,In_16,In_749);
or U2110 (N_2110,In_391,In_834);
and U2111 (N_2111,In_305,In_468);
nand U2112 (N_2112,In_751,In_788);
or U2113 (N_2113,In_578,In_139);
nand U2114 (N_2114,In_625,In_731);
and U2115 (N_2115,In_708,In_943);
and U2116 (N_2116,In_818,In_459);
nor U2117 (N_2117,In_541,In_149);
or U2118 (N_2118,In_467,In_826);
nor U2119 (N_2119,In_963,In_19);
and U2120 (N_2120,In_229,In_590);
or U2121 (N_2121,In_349,In_694);
or U2122 (N_2122,In_776,In_761);
or U2123 (N_2123,In_630,In_881);
nor U2124 (N_2124,In_159,In_899);
and U2125 (N_2125,In_269,In_407);
nor U2126 (N_2126,In_695,In_647);
nand U2127 (N_2127,In_884,In_920);
nand U2128 (N_2128,In_640,In_86);
nand U2129 (N_2129,In_276,In_62);
or U2130 (N_2130,In_819,In_104);
or U2131 (N_2131,In_903,In_469);
or U2132 (N_2132,In_796,In_854);
and U2133 (N_2133,In_571,In_589);
and U2134 (N_2134,In_693,In_558);
nand U2135 (N_2135,In_393,In_490);
and U2136 (N_2136,In_214,In_419);
nor U2137 (N_2137,In_784,In_339);
nand U2138 (N_2138,In_195,In_505);
and U2139 (N_2139,In_912,In_496);
nand U2140 (N_2140,In_60,In_656);
nor U2141 (N_2141,In_353,In_857);
nand U2142 (N_2142,In_659,In_444);
or U2143 (N_2143,In_983,In_638);
nand U2144 (N_2144,In_416,In_3);
nor U2145 (N_2145,In_151,In_774);
or U2146 (N_2146,In_589,In_997);
or U2147 (N_2147,In_347,In_570);
nor U2148 (N_2148,In_474,In_457);
and U2149 (N_2149,In_165,In_153);
or U2150 (N_2150,In_947,In_829);
or U2151 (N_2151,In_389,In_989);
and U2152 (N_2152,In_38,In_560);
or U2153 (N_2153,In_962,In_557);
and U2154 (N_2154,In_20,In_693);
or U2155 (N_2155,In_953,In_236);
nand U2156 (N_2156,In_57,In_301);
and U2157 (N_2157,In_886,In_128);
nor U2158 (N_2158,In_659,In_214);
and U2159 (N_2159,In_270,In_492);
or U2160 (N_2160,In_82,In_711);
or U2161 (N_2161,In_380,In_635);
xor U2162 (N_2162,In_236,In_723);
and U2163 (N_2163,In_102,In_887);
and U2164 (N_2164,In_55,In_801);
nand U2165 (N_2165,In_76,In_707);
nor U2166 (N_2166,In_284,In_505);
nor U2167 (N_2167,In_558,In_233);
nor U2168 (N_2168,In_976,In_583);
nand U2169 (N_2169,In_500,In_863);
and U2170 (N_2170,In_772,In_782);
and U2171 (N_2171,In_159,In_495);
nand U2172 (N_2172,In_19,In_536);
or U2173 (N_2173,In_113,In_985);
or U2174 (N_2174,In_938,In_880);
nor U2175 (N_2175,In_376,In_234);
nor U2176 (N_2176,In_428,In_442);
or U2177 (N_2177,In_855,In_820);
or U2178 (N_2178,In_274,In_24);
nor U2179 (N_2179,In_530,In_995);
and U2180 (N_2180,In_323,In_277);
nand U2181 (N_2181,In_57,In_406);
nor U2182 (N_2182,In_246,In_833);
and U2183 (N_2183,In_745,In_670);
or U2184 (N_2184,In_285,In_403);
and U2185 (N_2185,In_487,In_125);
or U2186 (N_2186,In_847,In_888);
xnor U2187 (N_2187,In_920,In_660);
or U2188 (N_2188,In_942,In_606);
or U2189 (N_2189,In_680,In_43);
and U2190 (N_2190,In_92,In_885);
nand U2191 (N_2191,In_267,In_119);
nor U2192 (N_2192,In_441,In_919);
nor U2193 (N_2193,In_414,In_329);
and U2194 (N_2194,In_483,In_153);
or U2195 (N_2195,In_816,In_247);
or U2196 (N_2196,In_309,In_394);
and U2197 (N_2197,In_18,In_900);
xor U2198 (N_2198,In_248,In_554);
or U2199 (N_2199,In_701,In_806);
or U2200 (N_2200,In_187,In_5);
nor U2201 (N_2201,In_528,In_95);
and U2202 (N_2202,In_429,In_952);
or U2203 (N_2203,In_819,In_251);
or U2204 (N_2204,In_974,In_761);
nand U2205 (N_2205,In_327,In_350);
nand U2206 (N_2206,In_198,In_845);
and U2207 (N_2207,In_618,In_351);
nor U2208 (N_2208,In_203,In_12);
nor U2209 (N_2209,In_95,In_967);
or U2210 (N_2210,In_342,In_626);
or U2211 (N_2211,In_289,In_639);
and U2212 (N_2212,In_805,In_801);
or U2213 (N_2213,In_133,In_71);
nor U2214 (N_2214,In_416,In_718);
nand U2215 (N_2215,In_341,In_592);
nor U2216 (N_2216,In_638,In_53);
or U2217 (N_2217,In_824,In_469);
nand U2218 (N_2218,In_431,In_124);
and U2219 (N_2219,In_202,In_438);
or U2220 (N_2220,In_613,In_148);
or U2221 (N_2221,In_556,In_398);
nor U2222 (N_2222,In_809,In_127);
xnor U2223 (N_2223,In_562,In_610);
nand U2224 (N_2224,In_90,In_592);
nor U2225 (N_2225,In_517,In_940);
nor U2226 (N_2226,In_991,In_359);
nor U2227 (N_2227,In_203,In_825);
nor U2228 (N_2228,In_538,In_988);
or U2229 (N_2229,In_190,In_981);
nor U2230 (N_2230,In_769,In_834);
nand U2231 (N_2231,In_194,In_296);
and U2232 (N_2232,In_240,In_871);
nor U2233 (N_2233,In_349,In_992);
nor U2234 (N_2234,In_314,In_828);
nor U2235 (N_2235,In_835,In_347);
nand U2236 (N_2236,In_172,In_436);
nor U2237 (N_2237,In_344,In_914);
or U2238 (N_2238,In_377,In_151);
or U2239 (N_2239,In_589,In_479);
nand U2240 (N_2240,In_597,In_224);
nor U2241 (N_2241,In_806,In_748);
nand U2242 (N_2242,In_525,In_953);
and U2243 (N_2243,In_40,In_108);
and U2244 (N_2244,In_426,In_702);
or U2245 (N_2245,In_156,In_611);
nor U2246 (N_2246,In_160,In_342);
nor U2247 (N_2247,In_37,In_485);
and U2248 (N_2248,In_243,In_453);
xnor U2249 (N_2249,In_952,In_101);
and U2250 (N_2250,In_179,In_115);
nand U2251 (N_2251,In_508,In_954);
nor U2252 (N_2252,In_427,In_775);
or U2253 (N_2253,In_928,In_672);
and U2254 (N_2254,In_33,In_910);
nand U2255 (N_2255,In_754,In_136);
xnor U2256 (N_2256,In_547,In_187);
and U2257 (N_2257,In_531,In_516);
and U2258 (N_2258,In_174,In_148);
nand U2259 (N_2259,In_469,In_936);
nand U2260 (N_2260,In_265,In_984);
nor U2261 (N_2261,In_749,In_102);
nand U2262 (N_2262,In_804,In_516);
or U2263 (N_2263,In_809,In_201);
or U2264 (N_2264,In_411,In_336);
and U2265 (N_2265,In_747,In_640);
and U2266 (N_2266,In_837,In_418);
nor U2267 (N_2267,In_429,In_564);
and U2268 (N_2268,In_393,In_255);
nand U2269 (N_2269,In_849,In_394);
or U2270 (N_2270,In_612,In_875);
and U2271 (N_2271,In_303,In_64);
nand U2272 (N_2272,In_79,In_949);
or U2273 (N_2273,In_45,In_387);
nor U2274 (N_2274,In_658,In_84);
nand U2275 (N_2275,In_7,In_512);
and U2276 (N_2276,In_736,In_374);
and U2277 (N_2277,In_113,In_890);
nand U2278 (N_2278,In_876,In_222);
and U2279 (N_2279,In_84,In_698);
and U2280 (N_2280,In_555,In_455);
and U2281 (N_2281,In_16,In_761);
xnor U2282 (N_2282,In_865,In_490);
and U2283 (N_2283,In_53,In_261);
nor U2284 (N_2284,In_599,In_471);
and U2285 (N_2285,In_491,In_328);
and U2286 (N_2286,In_611,In_965);
or U2287 (N_2287,In_69,In_268);
and U2288 (N_2288,In_685,In_231);
nor U2289 (N_2289,In_151,In_839);
and U2290 (N_2290,In_244,In_902);
nor U2291 (N_2291,In_640,In_572);
nor U2292 (N_2292,In_458,In_955);
or U2293 (N_2293,In_729,In_251);
nor U2294 (N_2294,In_693,In_106);
nor U2295 (N_2295,In_355,In_590);
nand U2296 (N_2296,In_629,In_129);
or U2297 (N_2297,In_142,In_532);
or U2298 (N_2298,In_409,In_911);
nor U2299 (N_2299,In_242,In_399);
nor U2300 (N_2300,In_563,In_254);
and U2301 (N_2301,In_572,In_969);
nand U2302 (N_2302,In_187,In_903);
and U2303 (N_2303,In_986,In_937);
nor U2304 (N_2304,In_347,In_753);
nand U2305 (N_2305,In_459,In_929);
nand U2306 (N_2306,In_429,In_586);
and U2307 (N_2307,In_704,In_983);
nand U2308 (N_2308,In_462,In_929);
or U2309 (N_2309,In_838,In_459);
or U2310 (N_2310,In_796,In_1);
and U2311 (N_2311,In_674,In_940);
and U2312 (N_2312,In_185,In_845);
or U2313 (N_2313,In_767,In_997);
or U2314 (N_2314,In_266,In_546);
or U2315 (N_2315,In_698,In_873);
nor U2316 (N_2316,In_521,In_600);
nor U2317 (N_2317,In_607,In_457);
and U2318 (N_2318,In_396,In_817);
or U2319 (N_2319,In_849,In_454);
and U2320 (N_2320,In_36,In_870);
nand U2321 (N_2321,In_342,In_405);
nor U2322 (N_2322,In_42,In_900);
or U2323 (N_2323,In_600,In_760);
nand U2324 (N_2324,In_205,In_797);
nand U2325 (N_2325,In_59,In_430);
and U2326 (N_2326,In_466,In_769);
nor U2327 (N_2327,In_488,In_144);
and U2328 (N_2328,In_890,In_429);
or U2329 (N_2329,In_387,In_19);
nand U2330 (N_2330,In_842,In_932);
or U2331 (N_2331,In_39,In_17);
nor U2332 (N_2332,In_585,In_440);
nor U2333 (N_2333,In_974,In_559);
or U2334 (N_2334,In_845,In_591);
nor U2335 (N_2335,In_62,In_426);
nor U2336 (N_2336,In_388,In_202);
and U2337 (N_2337,In_510,In_864);
or U2338 (N_2338,In_585,In_608);
or U2339 (N_2339,In_770,In_919);
or U2340 (N_2340,In_568,In_888);
nand U2341 (N_2341,In_299,In_607);
nand U2342 (N_2342,In_24,In_428);
nand U2343 (N_2343,In_90,In_729);
and U2344 (N_2344,In_24,In_446);
nand U2345 (N_2345,In_980,In_722);
nand U2346 (N_2346,In_69,In_696);
nor U2347 (N_2347,In_483,In_641);
nor U2348 (N_2348,In_232,In_140);
nand U2349 (N_2349,In_929,In_316);
and U2350 (N_2350,In_100,In_634);
nor U2351 (N_2351,In_897,In_556);
and U2352 (N_2352,In_415,In_913);
nor U2353 (N_2353,In_407,In_85);
nor U2354 (N_2354,In_535,In_486);
and U2355 (N_2355,In_345,In_794);
nand U2356 (N_2356,In_455,In_832);
or U2357 (N_2357,In_157,In_485);
nor U2358 (N_2358,In_678,In_86);
and U2359 (N_2359,In_743,In_583);
nand U2360 (N_2360,In_769,In_641);
and U2361 (N_2361,In_257,In_821);
or U2362 (N_2362,In_401,In_201);
or U2363 (N_2363,In_487,In_90);
nor U2364 (N_2364,In_533,In_847);
nand U2365 (N_2365,In_88,In_789);
nand U2366 (N_2366,In_332,In_755);
or U2367 (N_2367,In_168,In_601);
nor U2368 (N_2368,In_524,In_561);
nor U2369 (N_2369,In_806,In_128);
and U2370 (N_2370,In_397,In_82);
or U2371 (N_2371,In_59,In_300);
nor U2372 (N_2372,In_549,In_446);
or U2373 (N_2373,In_829,In_596);
and U2374 (N_2374,In_844,In_815);
or U2375 (N_2375,In_860,In_890);
nand U2376 (N_2376,In_12,In_250);
nor U2377 (N_2377,In_272,In_100);
nor U2378 (N_2378,In_225,In_880);
or U2379 (N_2379,In_961,In_488);
nand U2380 (N_2380,In_431,In_913);
nor U2381 (N_2381,In_113,In_35);
nand U2382 (N_2382,In_606,In_973);
nand U2383 (N_2383,In_181,In_934);
or U2384 (N_2384,In_787,In_737);
nor U2385 (N_2385,In_757,In_421);
or U2386 (N_2386,In_132,In_931);
nor U2387 (N_2387,In_577,In_134);
nand U2388 (N_2388,In_946,In_978);
nor U2389 (N_2389,In_251,In_228);
nor U2390 (N_2390,In_582,In_485);
nand U2391 (N_2391,In_713,In_803);
nand U2392 (N_2392,In_849,In_375);
or U2393 (N_2393,In_605,In_507);
or U2394 (N_2394,In_481,In_84);
nand U2395 (N_2395,In_236,In_108);
and U2396 (N_2396,In_201,In_786);
nand U2397 (N_2397,In_750,In_135);
nand U2398 (N_2398,In_364,In_596);
nand U2399 (N_2399,In_285,In_46);
and U2400 (N_2400,In_768,In_129);
and U2401 (N_2401,In_439,In_557);
and U2402 (N_2402,In_663,In_796);
and U2403 (N_2403,In_850,In_952);
or U2404 (N_2404,In_147,In_671);
and U2405 (N_2405,In_493,In_922);
or U2406 (N_2406,In_855,In_922);
or U2407 (N_2407,In_200,In_67);
nand U2408 (N_2408,In_250,In_353);
and U2409 (N_2409,In_877,In_61);
or U2410 (N_2410,In_655,In_113);
nand U2411 (N_2411,In_156,In_445);
nor U2412 (N_2412,In_490,In_554);
nand U2413 (N_2413,In_814,In_284);
nand U2414 (N_2414,In_135,In_499);
nor U2415 (N_2415,In_738,In_919);
nor U2416 (N_2416,In_348,In_739);
or U2417 (N_2417,In_929,In_489);
or U2418 (N_2418,In_54,In_336);
nand U2419 (N_2419,In_466,In_455);
and U2420 (N_2420,In_908,In_984);
and U2421 (N_2421,In_655,In_484);
or U2422 (N_2422,In_838,In_312);
and U2423 (N_2423,In_397,In_928);
nor U2424 (N_2424,In_154,In_270);
or U2425 (N_2425,In_788,In_338);
and U2426 (N_2426,In_638,In_230);
and U2427 (N_2427,In_59,In_825);
and U2428 (N_2428,In_539,In_708);
nor U2429 (N_2429,In_354,In_922);
nor U2430 (N_2430,In_9,In_812);
or U2431 (N_2431,In_434,In_933);
or U2432 (N_2432,In_753,In_162);
and U2433 (N_2433,In_9,In_822);
and U2434 (N_2434,In_886,In_853);
nand U2435 (N_2435,In_552,In_922);
and U2436 (N_2436,In_631,In_630);
or U2437 (N_2437,In_632,In_993);
nand U2438 (N_2438,In_59,In_728);
nand U2439 (N_2439,In_493,In_476);
or U2440 (N_2440,In_128,In_589);
and U2441 (N_2441,In_831,In_796);
and U2442 (N_2442,In_600,In_232);
or U2443 (N_2443,In_542,In_125);
and U2444 (N_2444,In_677,In_285);
or U2445 (N_2445,In_82,In_639);
or U2446 (N_2446,In_663,In_900);
nor U2447 (N_2447,In_301,In_140);
and U2448 (N_2448,In_637,In_594);
or U2449 (N_2449,In_257,In_22);
nor U2450 (N_2450,In_411,In_809);
nand U2451 (N_2451,In_516,In_337);
nor U2452 (N_2452,In_323,In_536);
and U2453 (N_2453,In_444,In_173);
or U2454 (N_2454,In_15,In_473);
nand U2455 (N_2455,In_772,In_800);
nand U2456 (N_2456,In_90,In_477);
nor U2457 (N_2457,In_298,In_874);
nand U2458 (N_2458,In_724,In_290);
and U2459 (N_2459,In_464,In_168);
nand U2460 (N_2460,In_389,In_99);
nand U2461 (N_2461,In_855,In_962);
nand U2462 (N_2462,In_846,In_402);
nor U2463 (N_2463,In_627,In_865);
or U2464 (N_2464,In_599,In_228);
nand U2465 (N_2465,In_384,In_217);
nor U2466 (N_2466,In_756,In_810);
and U2467 (N_2467,In_41,In_857);
and U2468 (N_2468,In_575,In_368);
or U2469 (N_2469,In_941,In_919);
and U2470 (N_2470,In_298,In_869);
nand U2471 (N_2471,In_588,In_999);
nor U2472 (N_2472,In_832,In_4);
nor U2473 (N_2473,In_2,In_806);
nand U2474 (N_2474,In_198,In_696);
or U2475 (N_2475,In_845,In_230);
nor U2476 (N_2476,In_243,In_156);
nand U2477 (N_2477,In_638,In_514);
nand U2478 (N_2478,In_748,In_727);
nand U2479 (N_2479,In_982,In_153);
and U2480 (N_2480,In_331,In_430);
or U2481 (N_2481,In_73,In_292);
or U2482 (N_2482,In_425,In_390);
nand U2483 (N_2483,In_601,In_913);
or U2484 (N_2484,In_829,In_720);
nand U2485 (N_2485,In_273,In_872);
and U2486 (N_2486,In_57,In_997);
and U2487 (N_2487,In_168,In_677);
nand U2488 (N_2488,In_991,In_458);
xnor U2489 (N_2489,In_418,In_333);
or U2490 (N_2490,In_534,In_283);
nand U2491 (N_2491,In_882,In_594);
and U2492 (N_2492,In_186,In_653);
nor U2493 (N_2493,In_0,In_77);
nor U2494 (N_2494,In_196,In_840);
or U2495 (N_2495,In_119,In_625);
nor U2496 (N_2496,In_690,In_225);
nor U2497 (N_2497,In_378,In_251);
and U2498 (N_2498,In_767,In_613);
nand U2499 (N_2499,In_929,In_192);
nor U2500 (N_2500,In_475,In_868);
and U2501 (N_2501,In_82,In_39);
nand U2502 (N_2502,In_614,In_386);
nor U2503 (N_2503,In_360,In_393);
nor U2504 (N_2504,In_252,In_577);
nor U2505 (N_2505,In_721,In_826);
and U2506 (N_2506,In_350,In_34);
nand U2507 (N_2507,In_107,In_704);
nand U2508 (N_2508,In_831,In_602);
nor U2509 (N_2509,In_666,In_826);
and U2510 (N_2510,In_288,In_460);
nor U2511 (N_2511,In_469,In_522);
nor U2512 (N_2512,In_258,In_44);
nor U2513 (N_2513,In_961,In_616);
nand U2514 (N_2514,In_14,In_269);
nor U2515 (N_2515,In_688,In_210);
nor U2516 (N_2516,In_289,In_898);
nand U2517 (N_2517,In_721,In_694);
nand U2518 (N_2518,In_834,In_363);
and U2519 (N_2519,In_585,In_642);
or U2520 (N_2520,In_493,In_414);
and U2521 (N_2521,In_939,In_244);
nand U2522 (N_2522,In_346,In_79);
or U2523 (N_2523,In_740,In_482);
nand U2524 (N_2524,In_107,In_455);
nor U2525 (N_2525,In_486,In_357);
or U2526 (N_2526,In_336,In_447);
and U2527 (N_2527,In_696,In_99);
nand U2528 (N_2528,In_891,In_871);
nor U2529 (N_2529,In_274,In_562);
and U2530 (N_2530,In_16,In_502);
and U2531 (N_2531,In_473,In_184);
and U2532 (N_2532,In_125,In_17);
and U2533 (N_2533,In_112,In_316);
nand U2534 (N_2534,In_598,In_219);
nor U2535 (N_2535,In_268,In_966);
nand U2536 (N_2536,In_511,In_44);
nor U2537 (N_2537,In_413,In_28);
and U2538 (N_2538,In_871,In_595);
nand U2539 (N_2539,In_274,In_103);
or U2540 (N_2540,In_829,In_41);
and U2541 (N_2541,In_57,In_526);
nor U2542 (N_2542,In_861,In_661);
and U2543 (N_2543,In_400,In_47);
nor U2544 (N_2544,In_193,In_771);
nand U2545 (N_2545,In_107,In_821);
or U2546 (N_2546,In_715,In_171);
nor U2547 (N_2547,In_145,In_816);
or U2548 (N_2548,In_539,In_112);
or U2549 (N_2549,In_971,In_606);
nor U2550 (N_2550,In_275,In_730);
or U2551 (N_2551,In_486,In_105);
nor U2552 (N_2552,In_170,In_31);
nor U2553 (N_2553,In_226,In_490);
or U2554 (N_2554,In_174,In_859);
and U2555 (N_2555,In_508,In_352);
nor U2556 (N_2556,In_445,In_747);
nand U2557 (N_2557,In_338,In_438);
and U2558 (N_2558,In_238,In_741);
and U2559 (N_2559,In_208,In_46);
or U2560 (N_2560,In_351,In_640);
and U2561 (N_2561,In_380,In_709);
or U2562 (N_2562,In_7,In_246);
and U2563 (N_2563,In_58,In_205);
or U2564 (N_2564,In_358,In_799);
nand U2565 (N_2565,In_168,In_371);
nand U2566 (N_2566,In_926,In_37);
nand U2567 (N_2567,In_856,In_660);
or U2568 (N_2568,In_439,In_748);
or U2569 (N_2569,In_925,In_779);
nor U2570 (N_2570,In_696,In_136);
nor U2571 (N_2571,In_181,In_317);
or U2572 (N_2572,In_15,In_822);
nor U2573 (N_2573,In_627,In_277);
or U2574 (N_2574,In_987,In_471);
and U2575 (N_2575,In_714,In_416);
or U2576 (N_2576,In_111,In_190);
nand U2577 (N_2577,In_421,In_615);
and U2578 (N_2578,In_260,In_325);
nand U2579 (N_2579,In_359,In_461);
nand U2580 (N_2580,In_391,In_232);
and U2581 (N_2581,In_937,In_300);
and U2582 (N_2582,In_645,In_563);
xor U2583 (N_2583,In_772,In_688);
nand U2584 (N_2584,In_930,In_890);
nand U2585 (N_2585,In_484,In_679);
and U2586 (N_2586,In_260,In_430);
nand U2587 (N_2587,In_202,In_336);
nand U2588 (N_2588,In_573,In_327);
nor U2589 (N_2589,In_15,In_795);
or U2590 (N_2590,In_291,In_247);
and U2591 (N_2591,In_644,In_388);
or U2592 (N_2592,In_296,In_570);
nor U2593 (N_2593,In_72,In_250);
nor U2594 (N_2594,In_912,In_780);
nand U2595 (N_2595,In_48,In_598);
nand U2596 (N_2596,In_278,In_494);
and U2597 (N_2597,In_396,In_918);
nand U2598 (N_2598,In_706,In_426);
and U2599 (N_2599,In_404,In_112);
or U2600 (N_2600,In_869,In_669);
and U2601 (N_2601,In_464,In_67);
nor U2602 (N_2602,In_956,In_346);
nor U2603 (N_2603,In_280,In_811);
or U2604 (N_2604,In_729,In_436);
nor U2605 (N_2605,In_751,In_168);
nor U2606 (N_2606,In_536,In_432);
or U2607 (N_2607,In_581,In_879);
and U2608 (N_2608,In_770,In_330);
nand U2609 (N_2609,In_662,In_663);
nor U2610 (N_2610,In_26,In_987);
nor U2611 (N_2611,In_570,In_622);
and U2612 (N_2612,In_157,In_441);
or U2613 (N_2613,In_450,In_25);
or U2614 (N_2614,In_358,In_349);
nor U2615 (N_2615,In_608,In_316);
and U2616 (N_2616,In_740,In_9);
nand U2617 (N_2617,In_775,In_597);
or U2618 (N_2618,In_674,In_14);
nor U2619 (N_2619,In_659,In_371);
or U2620 (N_2620,In_467,In_675);
and U2621 (N_2621,In_511,In_80);
nand U2622 (N_2622,In_401,In_890);
or U2623 (N_2623,In_678,In_814);
and U2624 (N_2624,In_867,In_561);
nor U2625 (N_2625,In_195,In_233);
and U2626 (N_2626,In_778,In_893);
and U2627 (N_2627,In_512,In_394);
or U2628 (N_2628,In_169,In_39);
and U2629 (N_2629,In_391,In_150);
or U2630 (N_2630,In_854,In_864);
and U2631 (N_2631,In_585,In_413);
and U2632 (N_2632,In_335,In_57);
nor U2633 (N_2633,In_450,In_91);
nor U2634 (N_2634,In_589,In_517);
nor U2635 (N_2635,In_85,In_284);
nand U2636 (N_2636,In_716,In_586);
or U2637 (N_2637,In_811,In_300);
nor U2638 (N_2638,In_321,In_523);
or U2639 (N_2639,In_489,In_775);
and U2640 (N_2640,In_446,In_472);
and U2641 (N_2641,In_47,In_355);
nand U2642 (N_2642,In_708,In_356);
or U2643 (N_2643,In_136,In_227);
nor U2644 (N_2644,In_855,In_363);
xnor U2645 (N_2645,In_430,In_201);
and U2646 (N_2646,In_76,In_344);
and U2647 (N_2647,In_835,In_474);
or U2648 (N_2648,In_219,In_131);
and U2649 (N_2649,In_842,In_20);
nor U2650 (N_2650,In_720,In_142);
and U2651 (N_2651,In_931,In_949);
and U2652 (N_2652,In_744,In_541);
or U2653 (N_2653,In_500,In_536);
nand U2654 (N_2654,In_242,In_339);
xnor U2655 (N_2655,In_576,In_682);
and U2656 (N_2656,In_937,In_485);
and U2657 (N_2657,In_138,In_184);
nand U2658 (N_2658,In_888,In_987);
nand U2659 (N_2659,In_523,In_902);
nor U2660 (N_2660,In_139,In_138);
and U2661 (N_2661,In_392,In_789);
and U2662 (N_2662,In_347,In_102);
or U2663 (N_2663,In_766,In_693);
nor U2664 (N_2664,In_334,In_429);
or U2665 (N_2665,In_52,In_326);
or U2666 (N_2666,In_291,In_713);
or U2667 (N_2667,In_630,In_136);
nand U2668 (N_2668,In_723,In_250);
nor U2669 (N_2669,In_780,In_443);
nand U2670 (N_2670,In_226,In_951);
xor U2671 (N_2671,In_310,In_334);
nand U2672 (N_2672,In_804,In_394);
nand U2673 (N_2673,In_97,In_36);
nand U2674 (N_2674,In_722,In_308);
and U2675 (N_2675,In_580,In_185);
nor U2676 (N_2676,In_73,In_298);
nor U2677 (N_2677,In_552,In_38);
and U2678 (N_2678,In_335,In_825);
nor U2679 (N_2679,In_457,In_556);
and U2680 (N_2680,In_884,In_508);
and U2681 (N_2681,In_588,In_492);
and U2682 (N_2682,In_166,In_229);
and U2683 (N_2683,In_905,In_466);
nand U2684 (N_2684,In_39,In_938);
or U2685 (N_2685,In_174,In_830);
nand U2686 (N_2686,In_622,In_178);
and U2687 (N_2687,In_262,In_865);
or U2688 (N_2688,In_974,In_748);
or U2689 (N_2689,In_781,In_103);
nor U2690 (N_2690,In_876,In_237);
nor U2691 (N_2691,In_639,In_415);
or U2692 (N_2692,In_829,In_614);
or U2693 (N_2693,In_305,In_26);
or U2694 (N_2694,In_61,In_802);
nor U2695 (N_2695,In_323,In_236);
nor U2696 (N_2696,In_841,In_898);
nand U2697 (N_2697,In_435,In_259);
or U2698 (N_2698,In_480,In_172);
nor U2699 (N_2699,In_142,In_561);
nand U2700 (N_2700,In_700,In_854);
and U2701 (N_2701,In_427,In_813);
and U2702 (N_2702,In_789,In_10);
nor U2703 (N_2703,In_332,In_868);
nand U2704 (N_2704,In_348,In_559);
nand U2705 (N_2705,In_955,In_313);
or U2706 (N_2706,In_287,In_891);
nand U2707 (N_2707,In_104,In_463);
nand U2708 (N_2708,In_737,In_522);
or U2709 (N_2709,In_446,In_613);
nand U2710 (N_2710,In_174,In_899);
and U2711 (N_2711,In_691,In_661);
nor U2712 (N_2712,In_592,In_850);
nand U2713 (N_2713,In_914,In_808);
and U2714 (N_2714,In_272,In_814);
or U2715 (N_2715,In_750,In_131);
or U2716 (N_2716,In_985,In_778);
or U2717 (N_2717,In_281,In_15);
and U2718 (N_2718,In_709,In_387);
or U2719 (N_2719,In_125,In_515);
nor U2720 (N_2720,In_655,In_522);
or U2721 (N_2721,In_517,In_438);
nor U2722 (N_2722,In_108,In_482);
xor U2723 (N_2723,In_179,In_509);
and U2724 (N_2724,In_389,In_342);
nor U2725 (N_2725,In_312,In_12);
nand U2726 (N_2726,In_549,In_452);
or U2727 (N_2727,In_137,In_944);
nand U2728 (N_2728,In_356,In_235);
nor U2729 (N_2729,In_457,In_281);
nor U2730 (N_2730,In_631,In_457);
nand U2731 (N_2731,In_338,In_412);
or U2732 (N_2732,In_912,In_514);
nor U2733 (N_2733,In_23,In_317);
nor U2734 (N_2734,In_931,In_589);
or U2735 (N_2735,In_218,In_149);
or U2736 (N_2736,In_345,In_40);
nand U2737 (N_2737,In_567,In_889);
nand U2738 (N_2738,In_999,In_95);
nor U2739 (N_2739,In_40,In_348);
or U2740 (N_2740,In_932,In_192);
or U2741 (N_2741,In_616,In_252);
and U2742 (N_2742,In_360,In_99);
nor U2743 (N_2743,In_160,In_227);
and U2744 (N_2744,In_555,In_416);
or U2745 (N_2745,In_647,In_334);
or U2746 (N_2746,In_982,In_298);
or U2747 (N_2747,In_707,In_480);
and U2748 (N_2748,In_6,In_238);
nand U2749 (N_2749,In_934,In_566);
or U2750 (N_2750,In_450,In_986);
and U2751 (N_2751,In_0,In_59);
and U2752 (N_2752,In_401,In_58);
or U2753 (N_2753,In_248,In_685);
nand U2754 (N_2754,In_433,In_875);
and U2755 (N_2755,In_241,In_855);
nor U2756 (N_2756,In_2,In_413);
nor U2757 (N_2757,In_885,In_683);
and U2758 (N_2758,In_65,In_933);
nand U2759 (N_2759,In_176,In_821);
nor U2760 (N_2760,In_797,In_905);
nand U2761 (N_2761,In_811,In_900);
nand U2762 (N_2762,In_200,In_16);
nand U2763 (N_2763,In_868,In_681);
nor U2764 (N_2764,In_215,In_383);
xor U2765 (N_2765,In_672,In_103);
and U2766 (N_2766,In_111,In_988);
nand U2767 (N_2767,In_503,In_730);
or U2768 (N_2768,In_442,In_83);
or U2769 (N_2769,In_132,In_245);
or U2770 (N_2770,In_835,In_908);
nor U2771 (N_2771,In_506,In_672);
or U2772 (N_2772,In_460,In_133);
nor U2773 (N_2773,In_658,In_587);
xor U2774 (N_2774,In_329,In_720);
nand U2775 (N_2775,In_255,In_541);
nor U2776 (N_2776,In_258,In_977);
nor U2777 (N_2777,In_996,In_218);
and U2778 (N_2778,In_206,In_674);
and U2779 (N_2779,In_620,In_684);
and U2780 (N_2780,In_325,In_864);
nor U2781 (N_2781,In_838,In_378);
nor U2782 (N_2782,In_944,In_274);
nor U2783 (N_2783,In_49,In_290);
and U2784 (N_2784,In_304,In_964);
nor U2785 (N_2785,In_788,In_322);
xnor U2786 (N_2786,In_199,In_844);
and U2787 (N_2787,In_485,In_602);
or U2788 (N_2788,In_703,In_67);
or U2789 (N_2789,In_525,In_481);
nand U2790 (N_2790,In_266,In_311);
nor U2791 (N_2791,In_663,In_724);
or U2792 (N_2792,In_575,In_941);
or U2793 (N_2793,In_703,In_452);
and U2794 (N_2794,In_585,In_625);
nor U2795 (N_2795,In_148,In_269);
nor U2796 (N_2796,In_177,In_797);
nor U2797 (N_2797,In_312,In_940);
and U2798 (N_2798,In_493,In_735);
nand U2799 (N_2799,In_66,In_259);
nand U2800 (N_2800,In_297,In_152);
or U2801 (N_2801,In_46,In_903);
and U2802 (N_2802,In_409,In_259);
and U2803 (N_2803,In_303,In_198);
nor U2804 (N_2804,In_100,In_987);
nor U2805 (N_2805,In_903,In_145);
and U2806 (N_2806,In_169,In_943);
nor U2807 (N_2807,In_678,In_29);
nand U2808 (N_2808,In_467,In_161);
and U2809 (N_2809,In_431,In_809);
nor U2810 (N_2810,In_841,In_676);
nand U2811 (N_2811,In_86,In_48);
nor U2812 (N_2812,In_13,In_770);
and U2813 (N_2813,In_958,In_986);
nor U2814 (N_2814,In_570,In_76);
or U2815 (N_2815,In_62,In_625);
and U2816 (N_2816,In_398,In_370);
or U2817 (N_2817,In_781,In_836);
or U2818 (N_2818,In_215,In_387);
and U2819 (N_2819,In_87,In_224);
nor U2820 (N_2820,In_605,In_923);
or U2821 (N_2821,In_783,In_323);
or U2822 (N_2822,In_371,In_59);
nand U2823 (N_2823,In_88,In_383);
nand U2824 (N_2824,In_296,In_724);
and U2825 (N_2825,In_682,In_18);
nand U2826 (N_2826,In_301,In_8);
or U2827 (N_2827,In_574,In_863);
nor U2828 (N_2828,In_888,In_119);
and U2829 (N_2829,In_138,In_549);
nor U2830 (N_2830,In_186,In_405);
xor U2831 (N_2831,In_995,In_498);
or U2832 (N_2832,In_6,In_718);
or U2833 (N_2833,In_167,In_483);
nand U2834 (N_2834,In_769,In_359);
or U2835 (N_2835,In_63,In_177);
and U2836 (N_2836,In_696,In_520);
and U2837 (N_2837,In_993,In_787);
and U2838 (N_2838,In_748,In_650);
nand U2839 (N_2839,In_170,In_886);
nand U2840 (N_2840,In_188,In_588);
nand U2841 (N_2841,In_855,In_973);
and U2842 (N_2842,In_161,In_576);
or U2843 (N_2843,In_864,In_368);
nand U2844 (N_2844,In_812,In_592);
or U2845 (N_2845,In_497,In_156);
nand U2846 (N_2846,In_569,In_416);
or U2847 (N_2847,In_93,In_105);
nand U2848 (N_2848,In_122,In_55);
or U2849 (N_2849,In_30,In_78);
or U2850 (N_2850,In_766,In_376);
or U2851 (N_2851,In_967,In_210);
nor U2852 (N_2852,In_423,In_10);
and U2853 (N_2853,In_163,In_21);
nand U2854 (N_2854,In_528,In_270);
and U2855 (N_2855,In_72,In_507);
and U2856 (N_2856,In_116,In_514);
and U2857 (N_2857,In_110,In_615);
nor U2858 (N_2858,In_600,In_164);
nor U2859 (N_2859,In_822,In_636);
nand U2860 (N_2860,In_713,In_807);
and U2861 (N_2861,In_355,In_967);
xnor U2862 (N_2862,In_218,In_723);
nand U2863 (N_2863,In_121,In_781);
and U2864 (N_2864,In_714,In_223);
or U2865 (N_2865,In_194,In_325);
or U2866 (N_2866,In_836,In_708);
and U2867 (N_2867,In_54,In_516);
nand U2868 (N_2868,In_96,In_903);
or U2869 (N_2869,In_704,In_154);
and U2870 (N_2870,In_685,In_380);
nor U2871 (N_2871,In_832,In_104);
and U2872 (N_2872,In_899,In_956);
and U2873 (N_2873,In_715,In_500);
nor U2874 (N_2874,In_492,In_241);
nand U2875 (N_2875,In_418,In_692);
nand U2876 (N_2876,In_992,In_136);
and U2877 (N_2877,In_572,In_85);
or U2878 (N_2878,In_38,In_938);
nand U2879 (N_2879,In_230,In_812);
nand U2880 (N_2880,In_119,In_95);
or U2881 (N_2881,In_516,In_298);
nor U2882 (N_2882,In_618,In_414);
and U2883 (N_2883,In_370,In_768);
nand U2884 (N_2884,In_929,In_129);
or U2885 (N_2885,In_812,In_697);
or U2886 (N_2886,In_575,In_582);
nor U2887 (N_2887,In_707,In_597);
and U2888 (N_2888,In_811,In_141);
or U2889 (N_2889,In_877,In_805);
or U2890 (N_2890,In_432,In_15);
or U2891 (N_2891,In_339,In_409);
nand U2892 (N_2892,In_582,In_860);
and U2893 (N_2893,In_951,In_360);
xor U2894 (N_2894,In_400,In_252);
and U2895 (N_2895,In_896,In_25);
nand U2896 (N_2896,In_804,In_268);
or U2897 (N_2897,In_477,In_669);
nand U2898 (N_2898,In_916,In_750);
nand U2899 (N_2899,In_311,In_236);
nor U2900 (N_2900,In_71,In_684);
nand U2901 (N_2901,In_476,In_486);
and U2902 (N_2902,In_560,In_435);
nand U2903 (N_2903,In_152,In_789);
nor U2904 (N_2904,In_435,In_692);
nand U2905 (N_2905,In_257,In_569);
or U2906 (N_2906,In_143,In_133);
nor U2907 (N_2907,In_867,In_324);
or U2908 (N_2908,In_984,In_43);
or U2909 (N_2909,In_200,In_882);
nand U2910 (N_2910,In_241,In_675);
nor U2911 (N_2911,In_115,In_63);
nand U2912 (N_2912,In_889,In_539);
nor U2913 (N_2913,In_481,In_997);
nand U2914 (N_2914,In_175,In_274);
nand U2915 (N_2915,In_894,In_300);
nand U2916 (N_2916,In_478,In_79);
nand U2917 (N_2917,In_699,In_68);
or U2918 (N_2918,In_340,In_581);
and U2919 (N_2919,In_919,In_477);
or U2920 (N_2920,In_530,In_977);
and U2921 (N_2921,In_66,In_634);
nand U2922 (N_2922,In_62,In_32);
and U2923 (N_2923,In_797,In_608);
nor U2924 (N_2924,In_505,In_296);
nand U2925 (N_2925,In_861,In_437);
and U2926 (N_2926,In_934,In_404);
or U2927 (N_2927,In_608,In_198);
nor U2928 (N_2928,In_710,In_100);
nor U2929 (N_2929,In_560,In_122);
and U2930 (N_2930,In_596,In_64);
and U2931 (N_2931,In_159,In_78);
nand U2932 (N_2932,In_991,In_15);
or U2933 (N_2933,In_199,In_757);
nand U2934 (N_2934,In_743,In_64);
or U2935 (N_2935,In_199,In_913);
nand U2936 (N_2936,In_489,In_719);
and U2937 (N_2937,In_844,In_379);
and U2938 (N_2938,In_982,In_288);
and U2939 (N_2939,In_613,In_57);
nand U2940 (N_2940,In_871,In_501);
nor U2941 (N_2941,In_225,In_577);
or U2942 (N_2942,In_459,In_623);
and U2943 (N_2943,In_786,In_27);
and U2944 (N_2944,In_496,In_690);
nor U2945 (N_2945,In_386,In_181);
and U2946 (N_2946,In_383,In_908);
and U2947 (N_2947,In_903,In_966);
and U2948 (N_2948,In_883,In_250);
and U2949 (N_2949,In_513,In_548);
nor U2950 (N_2950,In_356,In_276);
nand U2951 (N_2951,In_18,In_441);
or U2952 (N_2952,In_325,In_585);
nand U2953 (N_2953,In_298,In_697);
nor U2954 (N_2954,In_593,In_15);
nor U2955 (N_2955,In_31,In_465);
nor U2956 (N_2956,In_612,In_984);
or U2957 (N_2957,In_453,In_870);
nor U2958 (N_2958,In_918,In_365);
or U2959 (N_2959,In_162,In_157);
or U2960 (N_2960,In_758,In_776);
nand U2961 (N_2961,In_457,In_318);
and U2962 (N_2962,In_109,In_492);
nor U2963 (N_2963,In_394,In_401);
nor U2964 (N_2964,In_803,In_330);
and U2965 (N_2965,In_595,In_831);
and U2966 (N_2966,In_408,In_812);
or U2967 (N_2967,In_894,In_937);
xnor U2968 (N_2968,In_848,In_778);
nand U2969 (N_2969,In_588,In_642);
and U2970 (N_2970,In_476,In_807);
nand U2971 (N_2971,In_102,In_169);
and U2972 (N_2972,In_317,In_318);
and U2973 (N_2973,In_15,In_510);
or U2974 (N_2974,In_639,In_776);
nand U2975 (N_2975,In_49,In_813);
nand U2976 (N_2976,In_19,In_346);
and U2977 (N_2977,In_717,In_21);
nand U2978 (N_2978,In_845,In_175);
or U2979 (N_2979,In_571,In_233);
nor U2980 (N_2980,In_429,In_957);
or U2981 (N_2981,In_569,In_336);
and U2982 (N_2982,In_378,In_678);
nand U2983 (N_2983,In_396,In_753);
and U2984 (N_2984,In_382,In_196);
nand U2985 (N_2985,In_46,In_515);
or U2986 (N_2986,In_27,In_453);
nand U2987 (N_2987,In_724,In_411);
nor U2988 (N_2988,In_823,In_36);
or U2989 (N_2989,In_59,In_913);
or U2990 (N_2990,In_961,In_933);
nor U2991 (N_2991,In_662,In_546);
and U2992 (N_2992,In_571,In_705);
and U2993 (N_2993,In_419,In_765);
nor U2994 (N_2994,In_703,In_20);
or U2995 (N_2995,In_468,In_867);
or U2996 (N_2996,In_354,In_321);
or U2997 (N_2997,In_588,In_451);
or U2998 (N_2998,In_196,In_135);
nor U2999 (N_2999,In_26,In_340);
or U3000 (N_3000,In_694,In_657);
and U3001 (N_3001,In_479,In_453);
and U3002 (N_3002,In_611,In_870);
nand U3003 (N_3003,In_40,In_657);
nand U3004 (N_3004,In_809,In_980);
and U3005 (N_3005,In_546,In_241);
and U3006 (N_3006,In_270,In_688);
nor U3007 (N_3007,In_658,In_684);
and U3008 (N_3008,In_874,In_748);
or U3009 (N_3009,In_315,In_189);
and U3010 (N_3010,In_237,In_63);
nand U3011 (N_3011,In_639,In_37);
or U3012 (N_3012,In_421,In_463);
and U3013 (N_3013,In_907,In_638);
and U3014 (N_3014,In_230,In_619);
nand U3015 (N_3015,In_207,In_391);
nand U3016 (N_3016,In_899,In_776);
nor U3017 (N_3017,In_182,In_139);
or U3018 (N_3018,In_436,In_563);
nand U3019 (N_3019,In_185,In_472);
or U3020 (N_3020,In_433,In_415);
xor U3021 (N_3021,In_640,In_403);
nor U3022 (N_3022,In_715,In_440);
nand U3023 (N_3023,In_990,In_317);
nand U3024 (N_3024,In_377,In_478);
nor U3025 (N_3025,In_575,In_919);
or U3026 (N_3026,In_845,In_504);
and U3027 (N_3027,In_63,In_34);
nand U3028 (N_3028,In_685,In_53);
nor U3029 (N_3029,In_615,In_357);
and U3030 (N_3030,In_770,In_889);
or U3031 (N_3031,In_705,In_66);
and U3032 (N_3032,In_352,In_264);
and U3033 (N_3033,In_95,In_228);
and U3034 (N_3034,In_170,In_233);
and U3035 (N_3035,In_743,In_938);
and U3036 (N_3036,In_779,In_752);
or U3037 (N_3037,In_323,In_764);
or U3038 (N_3038,In_79,In_358);
and U3039 (N_3039,In_621,In_19);
and U3040 (N_3040,In_708,In_142);
or U3041 (N_3041,In_713,In_268);
nor U3042 (N_3042,In_824,In_724);
or U3043 (N_3043,In_401,In_138);
or U3044 (N_3044,In_21,In_875);
nor U3045 (N_3045,In_351,In_636);
and U3046 (N_3046,In_404,In_698);
nor U3047 (N_3047,In_476,In_212);
and U3048 (N_3048,In_792,In_500);
or U3049 (N_3049,In_458,In_388);
or U3050 (N_3050,In_664,In_703);
nor U3051 (N_3051,In_919,In_744);
or U3052 (N_3052,In_514,In_307);
and U3053 (N_3053,In_938,In_198);
or U3054 (N_3054,In_650,In_621);
nand U3055 (N_3055,In_816,In_578);
or U3056 (N_3056,In_755,In_153);
and U3057 (N_3057,In_417,In_990);
and U3058 (N_3058,In_45,In_358);
nor U3059 (N_3059,In_767,In_483);
nand U3060 (N_3060,In_205,In_595);
and U3061 (N_3061,In_713,In_696);
xor U3062 (N_3062,In_312,In_400);
nand U3063 (N_3063,In_612,In_57);
nand U3064 (N_3064,In_584,In_637);
or U3065 (N_3065,In_80,In_886);
nand U3066 (N_3066,In_163,In_603);
nand U3067 (N_3067,In_581,In_545);
and U3068 (N_3068,In_553,In_168);
or U3069 (N_3069,In_478,In_116);
nand U3070 (N_3070,In_426,In_399);
and U3071 (N_3071,In_689,In_471);
and U3072 (N_3072,In_639,In_884);
or U3073 (N_3073,In_717,In_647);
and U3074 (N_3074,In_561,In_717);
nand U3075 (N_3075,In_918,In_812);
or U3076 (N_3076,In_207,In_249);
nand U3077 (N_3077,In_909,In_847);
nand U3078 (N_3078,In_242,In_133);
nor U3079 (N_3079,In_103,In_34);
nand U3080 (N_3080,In_939,In_282);
nor U3081 (N_3081,In_77,In_662);
or U3082 (N_3082,In_393,In_940);
or U3083 (N_3083,In_821,In_591);
nand U3084 (N_3084,In_414,In_319);
and U3085 (N_3085,In_84,In_925);
nand U3086 (N_3086,In_447,In_91);
nand U3087 (N_3087,In_927,In_809);
and U3088 (N_3088,In_334,In_185);
or U3089 (N_3089,In_176,In_779);
or U3090 (N_3090,In_12,In_564);
nor U3091 (N_3091,In_894,In_845);
and U3092 (N_3092,In_550,In_407);
nand U3093 (N_3093,In_490,In_945);
or U3094 (N_3094,In_921,In_806);
nand U3095 (N_3095,In_879,In_574);
nand U3096 (N_3096,In_300,In_303);
nand U3097 (N_3097,In_158,In_555);
or U3098 (N_3098,In_416,In_700);
nand U3099 (N_3099,In_739,In_690);
or U3100 (N_3100,In_129,In_584);
and U3101 (N_3101,In_682,In_242);
and U3102 (N_3102,In_19,In_134);
xor U3103 (N_3103,In_64,In_299);
nand U3104 (N_3104,In_367,In_982);
and U3105 (N_3105,In_110,In_725);
xnor U3106 (N_3106,In_689,In_200);
and U3107 (N_3107,In_927,In_301);
nand U3108 (N_3108,In_948,In_578);
and U3109 (N_3109,In_445,In_387);
nor U3110 (N_3110,In_521,In_767);
nor U3111 (N_3111,In_860,In_767);
nor U3112 (N_3112,In_660,In_411);
or U3113 (N_3113,In_498,In_48);
nand U3114 (N_3114,In_865,In_524);
nand U3115 (N_3115,In_578,In_380);
nand U3116 (N_3116,In_680,In_136);
or U3117 (N_3117,In_690,In_426);
xor U3118 (N_3118,In_578,In_131);
nor U3119 (N_3119,In_470,In_152);
nor U3120 (N_3120,In_433,In_41);
or U3121 (N_3121,In_67,In_48);
nor U3122 (N_3122,In_135,In_980);
and U3123 (N_3123,In_83,In_437);
and U3124 (N_3124,In_623,In_522);
and U3125 (N_3125,In_631,In_73);
nor U3126 (N_3126,In_213,In_46);
and U3127 (N_3127,In_802,In_178);
nand U3128 (N_3128,In_776,In_319);
xor U3129 (N_3129,In_503,In_561);
nor U3130 (N_3130,In_765,In_377);
nand U3131 (N_3131,In_741,In_547);
and U3132 (N_3132,In_753,In_337);
nand U3133 (N_3133,In_353,In_987);
nor U3134 (N_3134,In_349,In_705);
nor U3135 (N_3135,In_881,In_449);
nand U3136 (N_3136,In_199,In_313);
or U3137 (N_3137,In_631,In_162);
and U3138 (N_3138,In_393,In_734);
nand U3139 (N_3139,In_99,In_48);
and U3140 (N_3140,In_228,In_912);
nor U3141 (N_3141,In_749,In_477);
nand U3142 (N_3142,In_972,In_239);
nor U3143 (N_3143,In_129,In_842);
or U3144 (N_3144,In_226,In_760);
and U3145 (N_3145,In_620,In_836);
and U3146 (N_3146,In_849,In_730);
or U3147 (N_3147,In_142,In_102);
and U3148 (N_3148,In_311,In_195);
nor U3149 (N_3149,In_736,In_731);
and U3150 (N_3150,In_754,In_405);
and U3151 (N_3151,In_766,In_560);
and U3152 (N_3152,In_66,In_288);
nor U3153 (N_3153,In_128,In_575);
nand U3154 (N_3154,In_666,In_282);
and U3155 (N_3155,In_251,In_398);
xnor U3156 (N_3156,In_863,In_206);
nand U3157 (N_3157,In_170,In_610);
nor U3158 (N_3158,In_837,In_421);
nand U3159 (N_3159,In_426,In_157);
nor U3160 (N_3160,In_905,In_970);
and U3161 (N_3161,In_67,In_44);
or U3162 (N_3162,In_888,In_842);
nand U3163 (N_3163,In_564,In_590);
nand U3164 (N_3164,In_758,In_671);
nand U3165 (N_3165,In_704,In_32);
nand U3166 (N_3166,In_765,In_319);
and U3167 (N_3167,In_823,In_482);
or U3168 (N_3168,In_974,In_311);
or U3169 (N_3169,In_284,In_198);
nand U3170 (N_3170,In_785,In_722);
nand U3171 (N_3171,In_662,In_528);
nor U3172 (N_3172,In_408,In_451);
nor U3173 (N_3173,In_965,In_400);
or U3174 (N_3174,In_168,In_692);
nand U3175 (N_3175,In_358,In_119);
and U3176 (N_3176,In_790,In_361);
nor U3177 (N_3177,In_266,In_948);
or U3178 (N_3178,In_850,In_514);
nor U3179 (N_3179,In_882,In_99);
or U3180 (N_3180,In_286,In_675);
nor U3181 (N_3181,In_519,In_417);
nand U3182 (N_3182,In_486,In_9);
nand U3183 (N_3183,In_864,In_915);
and U3184 (N_3184,In_446,In_830);
nor U3185 (N_3185,In_805,In_626);
nand U3186 (N_3186,In_307,In_836);
or U3187 (N_3187,In_286,In_163);
and U3188 (N_3188,In_241,In_586);
nor U3189 (N_3189,In_733,In_25);
nand U3190 (N_3190,In_599,In_548);
nand U3191 (N_3191,In_617,In_996);
and U3192 (N_3192,In_471,In_203);
and U3193 (N_3193,In_415,In_64);
nor U3194 (N_3194,In_44,In_570);
and U3195 (N_3195,In_623,In_963);
or U3196 (N_3196,In_259,In_486);
or U3197 (N_3197,In_787,In_762);
or U3198 (N_3198,In_871,In_990);
nor U3199 (N_3199,In_873,In_651);
nand U3200 (N_3200,In_279,In_448);
xor U3201 (N_3201,In_862,In_698);
nor U3202 (N_3202,In_423,In_734);
and U3203 (N_3203,In_543,In_550);
nand U3204 (N_3204,In_623,In_759);
or U3205 (N_3205,In_373,In_777);
and U3206 (N_3206,In_20,In_52);
and U3207 (N_3207,In_279,In_369);
nor U3208 (N_3208,In_828,In_759);
xnor U3209 (N_3209,In_933,In_198);
and U3210 (N_3210,In_218,In_675);
nand U3211 (N_3211,In_370,In_503);
or U3212 (N_3212,In_246,In_795);
nand U3213 (N_3213,In_206,In_939);
or U3214 (N_3214,In_520,In_302);
nand U3215 (N_3215,In_299,In_838);
and U3216 (N_3216,In_266,In_630);
and U3217 (N_3217,In_538,In_126);
and U3218 (N_3218,In_23,In_353);
nand U3219 (N_3219,In_843,In_998);
nand U3220 (N_3220,In_776,In_602);
nand U3221 (N_3221,In_234,In_549);
nor U3222 (N_3222,In_161,In_536);
nor U3223 (N_3223,In_309,In_307);
and U3224 (N_3224,In_595,In_830);
nor U3225 (N_3225,In_925,In_412);
nor U3226 (N_3226,In_482,In_208);
and U3227 (N_3227,In_288,In_670);
nand U3228 (N_3228,In_886,In_549);
nand U3229 (N_3229,In_398,In_876);
nand U3230 (N_3230,In_918,In_216);
nand U3231 (N_3231,In_966,In_601);
nand U3232 (N_3232,In_494,In_116);
nand U3233 (N_3233,In_80,In_535);
and U3234 (N_3234,In_846,In_559);
nor U3235 (N_3235,In_127,In_693);
or U3236 (N_3236,In_570,In_456);
nand U3237 (N_3237,In_452,In_864);
nand U3238 (N_3238,In_608,In_863);
nand U3239 (N_3239,In_351,In_877);
or U3240 (N_3240,In_784,In_42);
and U3241 (N_3241,In_634,In_30);
nor U3242 (N_3242,In_419,In_112);
or U3243 (N_3243,In_45,In_500);
nand U3244 (N_3244,In_103,In_874);
nand U3245 (N_3245,In_591,In_134);
nor U3246 (N_3246,In_104,In_243);
or U3247 (N_3247,In_361,In_885);
nand U3248 (N_3248,In_555,In_595);
nand U3249 (N_3249,In_363,In_724);
or U3250 (N_3250,In_569,In_651);
nand U3251 (N_3251,In_53,In_602);
nand U3252 (N_3252,In_539,In_689);
or U3253 (N_3253,In_624,In_676);
nor U3254 (N_3254,In_48,In_264);
and U3255 (N_3255,In_815,In_843);
nor U3256 (N_3256,In_387,In_482);
nor U3257 (N_3257,In_270,In_362);
xnor U3258 (N_3258,In_425,In_87);
or U3259 (N_3259,In_285,In_933);
nor U3260 (N_3260,In_139,In_876);
and U3261 (N_3261,In_289,In_869);
nand U3262 (N_3262,In_415,In_427);
nand U3263 (N_3263,In_994,In_481);
or U3264 (N_3264,In_925,In_404);
nor U3265 (N_3265,In_381,In_272);
nand U3266 (N_3266,In_500,In_497);
nand U3267 (N_3267,In_572,In_318);
or U3268 (N_3268,In_206,In_33);
nor U3269 (N_3269,In_146,In_544);
and U3270 (N_3270,In_802,In_324);
nor U3271 (N_3271,In_959,In_747);
nor U3272 (N_3272,In_136,In_262);
and U3273 (N_3273,In_560,In_315);
or U3274 (N_3274,In_977,In_674);
xnor U3275 (N_3275,In_974,In_680);
or U3276 (N_3276,In_216,In_163);
nor U3277 (N_3277,In_879,In_147);
or U3278 (N_3278,In_899,In_370);
nor U3279 (N_3279,In_89,In_995);
or U3280 (N_3280,In_720,In_278);
or U3281 (N_3281,In_604,In_485);
nor U3282 (N_3282,In_165,In_455);
nor U3283 (N_3283,In_930,In_321);
nor U3284 (N_3284,In_911,In_976);
and U3285 (N_3285,In_521,In_942);
nor U3286 (N_3286,In_464,In_151);
and U3287 (N_3287,In_422,In_515);
nand U3288 (N_3288,In_363,In_667);
nand U3289 (N_3289,In_508,In_892);
nor U3290 (N_3290,In_722,In_698);
nand U3291 (N_3291,In_242,In_475);
nor U3292 (N_3292,In_17,In_511);
and U3293 (N_3293,In_783,In_860);
and U3294 (N_3294,In_517,In_177);
and U3295 (N_3295,In_76,In_743);
nor U3296 (N_3296,In_435,In_596);
nor U3297 (N_3297,In_563,In_6);
and U3298 (N_3298,In_353,In_227);
or U3299 (N_3299,In_961,In_138);
or U3300 (N_3300,In_766,In_645);
or U3301 (N_3301,In_516,In_467);
nor U3302 (N_3302,In_886,In_65);
and U3303 (N_3303,In_178,In_266);
or U3304 (N_3304,In_120,In_923);
nand U3305 (N_3305,In_822,In_206);
nor U3306 (N_3306,In_580,In_201);
nor U3307 (N_3307,In_221,In_981);
nor U3308 (N_3308,In_372,In_225);
nand U3309 (N_3309,In_39,In_6);
or U3310 (N_3310,In_755,In_223);
nor U3311 (N_3311,In_775,In_609);
or U3312 (N_3312,In_435,In_554);
nand U3313 (N_3313,In_67,In_312);
nor U3314 (N_3314,In_414,In_186);
nand U3315 (N_3315,In_822,In_921);
and U3316 (N_3316,In_596,In_238);
nor U3317 (N_3317,In_739,In_591);
and U3318 (N_3318,In_463,In_870);
or U3319 (N_3319,In_835,In_503);
nor U3320 (N_3320,In_818,In_85);
nor U3321 (N_3321,In_801,In_804);
nor U3322 (N_3322,In_825,In_211);
nand U3323 (N_3323,In_137,In_67);
and U3324 (N_3324,In_788,In_317);
xor U3325 (N_3325,In_852,In_608);
nand U3326 (N_3326,In_867,In_235);
nand U3327 (N_3327,In_140,In_598);
nor U3328 (N_3328,In_176,In_678);
or U3329 (N_3329,In_192,In_663);
nor U3330 (N_3330,In_411,In_635);
and U3331 (N_3331,In_847,In_101);
nor U3332 (N_3332,In_408,In_808);
and U3333 (N_3333,In_829,In_19);
and U3334 (N_3334,In_650,In_159);
or U3335 (N_3335,In_136,In_766);
nand U3336 (N_3336,In_951,In_191);
or U3337 (N_3337,In_94,In_822);
and U3338 (N_3338,In_949,In_454);
nand U3339 (N_3339,In_445,In_989);
and U3340 (N_3340,In_212,In_200);
nand U3341 (N_3341,In_991,In_890);
or U3342 (N_3342,In_387,In_332);
nand U3343 (N_3343,In_149,In_550);
nor U3344 (N_3344,In_826,In_14);
nand U3345 (N_3345,In_86,In_136);
xnor U3346 (N_3346,In_481,In_580);
nor U3347 (N_3347,In_805,In_528);
or U3348 (N_3348,In_232,In_863);
or U3349 (N_3349,In_583,In_983);
or U3350 (N_3350,In_928,In_883);
nor U3351 (N_3351,In_551,In_854);
nor U3352 (N_3352,In_513,In_216);
or U3353 (N_3353,In_338,In_174);
nand U3354 (N_3354,In_615,In_246);
or U3355 (N_3355,In_397,In_664);
nor U3356 (N_3356,In_740,In_970);
or U3357 (N_3357,In_616,In_285);
nor U3358 (N_3358,In_797,In_187);
or U3359 (N_3359,In_376,In_702);
nor U3360 (N_3360,In_65,In_502);
or U3361 (N_3361,In_311,In_818);
or U3362 (N_3362,In_65,In_697);
nand U3363 (N_3363,In_433,In_332);
and U3364 (N_3364,In_130,In_244);
and U3365 (N_3365,In_168,In_559);
and U3366 (N_3366,In_708,In_295);
or U3367 (N_3367,In_468,In_221);
nand U3368 (N_3368,In_313,In_100);
or U3369 (N_3369,In_218,In_704);
and U3370 (N_3370,In_589,In_170);
and U3371 (N_3371,In_691,In_805);
nor U3372 (N_3372,In_66,In_783);
nand U3373 (N_3373,In_446,In_730);
nand U3374 (N_3374,In_448,In_805);
or U3375 (N_3375,In_507,In_550);
nand U3376 (N_3376,In_371,In_572);
or U3377 (N_3377,In_155,In_731);
and U3378 (N_3378,In_151,In_926);
nand U3379 (N_3379,In_251,In_763);
or U3380 (N_3380,In_91,In_659);
nor U3381 (N_3381,In_947,In_573);
nand U3382 (N_3382,In_85,In_0);
nor U3383 (N_3383,In_968,In_155);
nor U3384 (N_3384,In_589,In_37);
and U3385 (N_3385,In_817,In_776);
and U3386 (N_3386,In_501,In_331);
nor U3387 (N_3387,In_900,In_709);
and U3388 (N_3388,In_740,In_415);
and U3389 (N_3389,In_189,In_609);
nand U3390 (N_3390,In_510,In_988);
nor U3391 (N_3391,In_912,In_219);
nand U3392 (N_3392,In_461,In_478);
nor U3393 (N_3393,In_1,In_905);
nor U3394 (N_3394,In_934,In_227);
or U3395 (N_3395,In_656,In_98);
and U3396 (N_3396,In_529,In_83);
and U3397 (N_3397,In_551,In_271);
nor U3398 (N_3398,In_123,In_572);
nand U3399 (N_3399,In_119,In_904);
and U3400 (N_3400,In_281,In_475);
nor U3401 (N_3401,In_309,In_593);
or U3402 (N_3402,In_225,In_424);
and U3403 (N_3403,In_186,In_864);
nand U3404 (N_3404,In_697,In_600);
nand U3405 (N_3405,In_789,In_551);
nand U3406 (N_3406,In_642,In_410);
nand U3407 (N_3407,In_929,In_812);
nor U3408 (N_3408,In_185,In_687);
and U3409 (N_3409,In_798,In_772);
nor U3410 (N_3410,In_7,In_437);
nor U3411 (N_3411,In_258,In_583);
and U3412 (N_3412,In_359,In_815);
and U3413 (N_3413,In_889,In_32);
nand U3414 (N_3414,In_52,In_457);
and U3415 (N_3415,In_773,In_584);
nand U3416 (N_3416,In_768,In_153);
and U3417 (N_3417,In_316,In_3);
and U3418 (N_3418,In_356,In_850);
nor U3419 (N_3419,In_149,In_403);
or U3420 (N_3420,In_665,In_68);
nand U3421 (N_3421,In_313,In_45);
or U3422 (N_3422,In_561,In_935);
and U3423 (N_3423,In_20,In_433);
nand U3424 (N_3424,In_287,In_670);
nand U3425 (N_3425,In_716,In_671);
or U3426 (N_3426,In_78,In_984);
and U3427 (N_3427,In_263,In_851);
nor U3428 (N_3428,In_366,In_980);
nand U3429 (N_3429,In_296,In_740);
and U3430 (N_3430,In_23,In_280);
and U3431 (N_3431,In_829,In_863);
and U3432 (N_3432,In_443,In_18);
nand U3433 (N_3433,In_481,In_734);
or U3434 (N_3434,In_790,In_427);
and U3435 (N_3435,In_390,In_697);
nor U3436 (N_3436,In_793,In_5);
and U3437 (N_3437,In_786,In_359);
nor U3438 (N_3438,In_197,In_904);
nand U3439 (N_3439,In_263,In_125);
xnor U3440 (N_3440,In_660,In_853);
nand U3441 (N_3441,In_871,In_38);
nand U3442 (N_3442,In_36,In_669);
nor U3443 (N_3443,In_37,In_539);
and U3444 (N_3444,In_417,In_450);
nand U3445 (N_3445,In_870,In_84);
nand U3446 (N_3446,In_52,In_222);
nand U3447 (N_3447,In_296,In_986);
and U3448 (N_3448,In_878,In_501);
nor U3449 (N_3449,In_121,In_785);
and U3450 (N_3450,In_577,In_716);
nand U3451 (N_3451,In_939,In_799);
nor U3452 (N_3452,In_442,In_731);
and U3453 (N_3453,In_918,In_871);
or U3454 (N_3454,In_21,In_314);
nor U3455 (N_3455,In_504,In_935);
and U3456 (N_3456,In_769,In_721);
nor U3457 (N_3457,In_165,In_726);
or U3458 (N_3458,In_44,In_762);
nand U3459 (N_3459,In_337,In_801);
and U3460 (N_3460,In_733,In_470);
nor U3461 (N_3461,In_163,In_612);
nand U3462 (N_3462,In_927,In_164);
and U3463 (N_3463,In_345,In_447);
nor U3464 (N_3464,In_92,In_549);
and U3465 (N_3465,In_122,In_54);
and U3466 (N_3466,In_559,In_268);
nor U3467 (N_3467,In_444,In_266);
nand U3468 (N_3468,In_836,In_96);
xor U3469 (N_3469,In_384,In_473);
or U3470 (N_3470,In_25,In_291);
nor U3471 (N_3471,In_870,In_874);
nand U3472 (N_3472,In_614,In_275);
nand U3473 (N_3473,In_51,In_836);
or U3474 (N_3474,In_117,In_581);
nand U3475 (N_3475,In_236,In_679);
or U3476 (N_3476,In_543,In_964);
nor U3477 (N_3477,In_123,In_953);
or U3478 (N_3478,In_876,In_734);
nand U3479 (N_3479,In_860,In_558);
or U3480 (N_3480,In_676,In_348);
and U3481 (N_3481,In_144,In_233);
and U3482 (N_3482,In_257,In_3);
nor U3483 (N_3483,In_906,In_595);
nand U3484 (N_3484,In_438,In_525);
and U3485 (N_3485,In_932,In_931);
and U3486 (N_3486,In_744,In_372);
and U3487 (N_3487,In_939,In_751);
and U3488 (N_3488,In_139,In_249);
nand U3489 (N_3489,In_193,In_851);
or U3490 (N_3490,In_611,In_546);
or U3491 (N_3491,In_967,In_568);
nand U3492 (N_3492,In_559,In_662);
nor U3493 (N_3493,In_815,In_535);
and U3494 (N_3494,In_437,In_482);
nor U3495 (N_3495,In_285,In_21);
nand U3496 (N_3496,In_231,In_405);
nor U3497 (N_3497,In_384,In_397);
or U3498 (N_3498,In_871,In_846);
and U3499 (N_3499,In_389,In_494);
nor U3500 (N_3500,In_257,In_836);
nand U3501 (N_3501,In_904,In_420);
nand U3502 (N_3502,In_497,In_128);
and U3503 (N_3503,In_736,In_15);
and U3504 (N_3504,In_682,In_504);
nor U3505 (N_3505,In_289,In_972);
and U3506 (N_3506,In_180,In_368);
nand U3507 (N_3507,In_738,In_312);
nand U3508 (N_3508,In_792,In_869);
or U3509 (N_3509,In_588,In_329);
nand U3510 (N_3510,In_797,In_530);
nand U3511 (N_3511,In_415,In_558);
nand U3512 (N_3512,In_762,In_853);
or U3513 (N_3513,In_205,In_357);
nand U3514 (N_3514,In_114,In_342);
nor U3515 (N_3515,In_529,In_412);
or U3516 (N_3516,In_753,In_734);
nand U3517 (N_3517,In_905,In_671);
nand U3518 (N_3518,In_787,In_530);
or U3519 (N_3519,In_990,In_817);
and U3520 (N_3520,In_770,In_942);
xnor U3521 (N_3521,In_833,In_824);
nand U3522 (N_3522,In_432,In_278);
nand U3523 (N_3523,In_558,In_5);
nor U3524 (N_3524,In_851,In_56);
nor U3525 (N_3525,In_840,In_887);
or U3526 (N_3526,In_969,In_647);
and U3527 (N_3527,In_3,In_763);
or U3528 (N_3528,In_679,In_432);
nor U3529 (N_3529,In_526,In_46);
or U3530 (N_3530,In_134,In_203);
nor U3531 (N_3531,In_97,In_385);
nand U3532 (N_3532,In_656,In_19);
nand U3533 (N_3533,In_781,In_513);
xor U3534 (N_3534,In_31,In_133);
nand U3535 (N_3535,In_436,In_635);
nor U3536 (N_3536,In_881,In_686);
nor U3537 (N_3537,In_813,In_905);
and U3538 (N_3538,In_629,In_651);
and U3539 (N_3539,In_667,In_130);
or U3540 (N_3540,In_388,In_467);
nor U3541 (N_3541,In_201,In_284);
and U3542 (N_3542,In_87,In_17);
nand U3543 (N_3543,In_764,In_917);
or U3544 (N_3544,In_652,In_8);
or U3545 (N_3545,In_701,In_256);
and U3546 (N_3546,In_467,In_609);
nor U3547 (N_3547,In_635,In_748);
or U3548 (N_3548,In_264,In_569);
nand U3549 (N_3549,In_574,In_899);
or U3550 (N_3550,In_621,In_886);
or U3551 (N_3551,In_171,In_142);
or U3552 (N_3552,In_675,In_784);
nand U3553 (N_3553,In_433,In_985);
and U3554 (N_3554,In_887,In_742);
nand U3555 (N_3555,In_704,In_780);
or U3556 (N_3556,In_275,In_537);
or U3557 (N_3557,In_491,In_589);
nor U3558 (N_3558,In_930,In_750);
nor U3559 (N_3559,In_168,In_118);
and U3560 (N_3560,In_676,In_926);
nand U3561 (N_3561,In_238,In_480);
nor U3562 (N_3562,In_339,In_333);
and U3563 (N_3563,In_731,In_251);
nand U3564 (N_3564,In_927,In_752);
nor U3565 (N_3565,In_617,In_222);
or U3566 (N_3566,In_740,In_161);
nand U3567 (N_3567,In_91,In_49);
nor U3568 (N_3568,In_82,In_550);
nor U3569 (N_3569,In_887,In_796);
and U3570 (N_3570,In_477,In_299);
nand U3571 (N_3571,In_701,In_234);
or U3572 (N_3572,In_453,In_538);
nand U3573 (N_3573,In_759,In_932);
nand U3574 (N_3574,In_266,In_529);
or U3575 (N_3575,In_344,In_240);
nand U3576 (N_3576,In_526,In_109);
nor U3577 (N_3577,In_82,In_882);
or U3578 (N_3578,In_755,In_990);
nand U3579 (N_3579,In_998,In_965);
nor U3580 (N_3580,In_542,In_576);
nand U3581 (N_3581,In_466,In_925);
nor U3582 (N_3582,In_68,In_92);
and U3583 (N_3583,In_148,In_753);
nand U3584 (N_3584,In_573,In_715);
or U3585 (N_3585,In_55,In_591);
or U3586 (N_3586,In_301,In_338);
and U3587 (N_3587,In_360,In_132);
or U3588 (N_3588,In_334,In_162);
nor U3589 (N_3589,In_85,In_138);
or U3590 (N_3590,In_844,In_965);
or U3591 (N_3591,In_390,In_695);
nand U3592 (N_3592,In_73,In_656);
nor U3593 (N_3593,In_213,In_65);
nor U3594 (N_3594,In_570,In_123);
nor U3595 (N_3595,In_848,In_565);
nor U3596 (N_3596,In_901,In_177);
or U3597 (N_3597,In_375,In_828);
nand U3598 (N_3598,In_437,In_652);
and U3599 (N_3599,In_282,In_152);
and U3600 (N_3600,In_800,In_813);
or U3601 (N_3601,In_74,In_889);
nor U3602 (N_3602,In_37,In_285);
or U3603 (N_3603,In_441,In_124);
nor U3604 (N_3604,In_541,In_365);
or U3605 (N_3605,In_846,In_594);
or U3606 (N_3606,In_786,In_788);
nand U3607 (N_3607,In_568,In_17);
nor U3608 (N_3608,In_846,In_808);
nand U3609 (N_3609,In_38,In_296);
and U3610 (N_3610,In_152,In_605);
nor U3611 (N_3611,In_670,In_264);
nor U3612 (N_3612,In_123,In_213);
nand U3613 (N_3613,In_159,In_92);
nand U3614 (N_3614,In_807,In_436);
nand U3615 (N_3615,In_928,In_338);
and U3616 (N_3616,In_10,In_435);
and U3617 (N_3617,In_154,In_959);
and U3618 (N_3618,In_292,In_121);
or U3619 (N_3619,In_384,In_396);
or U3620 (N_3620,In_354,In_366);
nand U3621 (N_3621,In_753,In_237);
nand U3622 (N_3622,In_923,In_917);
nand U3623 (N_3623,In_301,In_122);
or U3624 (N_3624,In_654,In_931);
or U3625 (N_3625,In_424,In_195);
and U3626 (N_3626,In_24,In_501);
nor U3627 (N_3627,In_890,In_808);
or U3628 (N_3628,In_858,In_724);
nor U3629 (N_3629,In_457,In_552);
or U3630 (N_3630,In_886,In_433);
nand U3631 (N_3631,In_885,In_484);
nor U3632 (N_3632,In_719,In_237);
or U3633 (N_3633,In_284,In_437);
nor U3634 (N_3634,In_441,In_567);
or U3635 (N_3635,In_355,In_188);
and U3636 (N_3636,In_618,In_393);
nor U3637 (N_3637,In_413,In_221);
or U3638 (N_3638,In_974,In_503);
and U3639 (N_3639,In_323,In_166);
and U3640 (N_3640,In_312,In_10);
nand U3641 (N_3641,In_76,In_560);
nand U3642 (N_3642,In_734,In_925);
nor U3643 (N_3643,In_312,In_861);
nand U3644 (N_3644,In_178,In_249);
nand U3645 (N_3645,In_841,In_229);
nand U3646 (N_3646,In_914,In_746);
nand U3647 (N_3647,In_717,In_232);
and U3648 (N_3648,In_469,In_253);
nor U3649 (N_3649,In_779,In_73);
or U3650 (N_3650,In_101,In_707);
nand U3651 (N_3651,In_85,In_342);
or U3652 (N_3652,In_340,In_150);
and U3653 (N_3653,In_354,In_873);
and U3654 (N_3654,In_939,In_431);
nor U3655 (N_3655,In_44,In_362);
and U3656 (N_3656,In_105,In_523);
or U3657 (N_3657,In_427,In_300);
nor U3658 (N_3658,In_277,In_833);
and U3659 (N_3659,In_112,In_382);
and U3660 (N_3660,In_216,In_47);
and U3661 (N_3661,In_650,In_292);
or U3662 (N_3662,In_474,In_136);
nand U3663 (N_3663,In_939,In_678);
and U3664 (N_3664,In_688,In_455);
and U3665 (N_3665,In_645,In_117);
nand U3666 (N_3666,In_305,In_615);
or U3667 (N_3667,In_39,In_198);
or U3668 (N_3668,In_792,In_50);
nand U3669 (N_3669,In_756,In_175);
or U3670 (N_3670,In_715,In_152);
nand U3671 (N_3671,In_357,In_142);
nor U3672 (N_3672,In_193,In_847);
nand U3673 (N_3673,In_514,In_546);
or U3674 (N_3674,In_193,In_361);
or U3675 (N_3675,In_129,In_91);
or U3676 (N_3676,In_168,In_159);
nand U3677 (N_3677,In_518,In_510);
and U3678 (N_3678,In_525,In_976);
nor U3679 (N_3679,In_543,In_566);
nand U3680 (N_3680,In_887,In_326);
nand U3681 (N_3681,In_289,In_344);
nand U3682 (N_3682,In_963,In_145);
nor U3683 (N_3683,In_700,In_325);
or U3684 (N_3684,In_818,In_246);
or U3685 (N_3685,In_5,In_332);
or U3686 (N_3686,In_126,In_80);
nor U3687 (N_3687,In_391,In_909);
and U3688 (N_3688,In_211,In_294);
nor U3689 (N_3689,In_924,In_475);
and U3690 (N_3690,In_218,In_569);
nand U3691 (N_3691,In_680,In_50);
or U3692 (N_3692,In_275,In_106);
and U3693 (N_3693,In_506,In_543);
nand U3694 (N_3694,In_888,In_801);
or U3695 (N_3695,In_920,In_811);
nor U3696 (N_3696,In_180,In_128);
nor U3697 (N_3697,In_562,In_10);
and U3698 (N_3698,In_44,In_326);
or U3699 (N_3699,In_257,In_382);
or U3700 (N_3700,In_757,In_255);
and U3701 (N_3701,In_839,In_367);
and U3702 (N_3702,In_457,In_217);
or U3703 (N_3703,In_640,In_849);
or U3704 (N_3704,In_868,In_652);
and U3705 (N_3705,In_534,In_919);
nor U3706 (N_3706,In_793,In_934);
and U3707 (N_3707,In_20,In_449);
and U3708 (N_3708,In_512,In_287);
nand U3709 (N_3709,In_36,In_733);
and U3710 (N_3710,In_249,In_321);
nand U3711 (N_3711,In_58,In_979);
nand U3712 (N_3712,In_712,In_135);
or U3713 (N_3713,In_239,In_236);
nor U3714 (N_3714,In_411,In_149);
nor U3715 (N_3715,In_148,In_153);
and U3716 (N_3716,In_25,In_681);
nor U3717 (N_3717,In_658,In_883);
nand U3718 (N_3718,In_173,In_919);
or U3719 (N_3719,In_924,In_562);
nand U3720 (N_3720,In_962,In_976);
or U3721 (N_3721,In_787,In_392);
nand U3722 (N_3722,In_605,In_23);
or U3723 (N_3723,In_969,In_68);
or U3724 (N_3724,In_120,In_539);
nor U3725 (N_3725,In_25,In_194);
nand U3726 (N_3726,In_418,In_543);
or U3727 (N_3727,In_453,In_245);
nand U3728 (N_3728,In_498,In_853);
nand U3729 (N_3729,In_460,In_113);
nand U3730 (N_3730,In_332,In_528);
nand U3731 (N_3731,In_602,In_947);
nand U3732 (N_3732,In_482,In_617);
nor U3733 (N_3733,In_564,In_537);
nand U3734 (N_3734,In_299,In_259);
nand U3735 (N_3735,In_245,In_445);
or U3736 (N_3736,In_362,In_665);
nand U3737 (N_3737,In_634,In_909);
and U3738 (N_3738,In_271,In_593);
nor U3739 (N_3739,In_156,In_257);
and U3740 (N_3740,In_780,In_461);
and U3741 (N_3741,In_244,In_634);
or U3742 (N_3742,In_618,In_861);
or U3743 (N_3743,In_618,In_295);
and U3744 (N_3744,In_92,In_355);
and U3745 (N_3745,In_182,In_393);
and U3746 (N_3746,In_865,In_79);
nand U3747 (N_3747,In_821,In_598);
or U3748 (N_3748,In_227,In_953);
and U3749 (N_3749,In_881,In_340);
nand U3750 (N_3750,In_162,In_258);
or U3751 (N_3751,In_120,In_451);
and U3752 (N_3752,In_243,In_339);
and U3753 (N_3753,In_178,In_749);
nor U3754 (N_3754,In_824,In_786);
or U3755 (N_3755,In_590,In_10);
nand U3756 (N_3756,In_892,In_611);
or U3757 (N_3757,In_402,In_293);
nand U3758 (N_3758,In_825,In_237);
and U3759 (N_3759,In_876,In_49);
or U3760 (N_3760,In_30,In_300);
nor U3761 (N_3761,In_41,In_782);
or U3762 (N_3762,In_287,In_942);
or U3763 (N_3763,In_597,In_645);
nand U3764 (N_3764,In_163,In_478);
nor U3765 (N_3765,In_988,In_572);
nand U3766 (N_3766,In_350,In_843);
and U3767 (N_3767,In_141,In_787);
nand U3768 (N_3768,In_171,In_351);
nor U3769 (N_3769,In_867,In_970);
or U3770 (N_3770,In_506,In_556);
nand U3771 (N_3771,In_186,In_523);
or U3772 (N_3772,In_9,In_364);
nand U3773 (N_3773,In_279,In_882);
and U3774 (N_3774,In_292,In_583);
or U3775 (N_3775,In_202,In_42);
nand U3776 (N_3776,In_8,In_821);
and U3777 (N_3777,In_739,In_330);
or U3778 (N_3778,In_406,In_910);
or U3779 (N_3779,In_988,In_531);
or U3780 (N_3780,In_167,In_740);
or U3781 (N_3781,In_283,In_266);
and U3782 (N_3782,In_33,In_1);
and U3783 (N_3783,In_745,In_232);
or U3784 (N_3784,In_68,In_539);
and U3785 (N_3785,In_882,In_316);
nor U3786 (N_3786,In_809,In_962);
or U3787 (N_3787,In_395,In_447);
or U3788 (N_3788,In_921,In_956);
nand U3789 (N_3789,In_612,In_145);
nand U3790 (N_3790,In_95,In_6);
nor U3791 (N_3791,In_971,In_202);
nor U3792 (N_3792,In_37,In_800);
and U3793 (N_3793,In_856,In_635);
nand U3794 (N_3794,In_379,In_278);
and U3795 (N_3795,In_140,In_592);
or U3796 (N_3796,In_229,In_902);
or U3797 (N_3797,In_604,In_611);
nand U3798 (N_3798,In_86,In_941);
nor U3799 (N_3799,In_109,In_138);
nor U3800 (N_3800,In_833,In_637);
or U3801 (N_3801,In_310,In_424);
nor U3802 (N_3802,In_567,In_151);
nand U3803 (N_3803,In_199,In_624);
nor U3804 (N_3804,In_429,In_205);
or U3805 (N_3805,In_541,In_13);
nand U3806 (N_3806,In_288,In_848);
and U3807 (N_3807,In_301,In_106);
nor U3808 (N_3808,In_886,In_353);
or U3809 (N_3809,In_602,In_366);
and U3810 (N_3810,In_867,In_877);
and U3811 (N_3811,In_962,In_533);
xnor U3812 (N_3812,In_769,In_513);
and U3813 (N_3813,In_694,In_511);
and U3814 (N_3814,In_882,In_613);
or U3815 (N_3815,In_990,In_963);
nor U3816 (N_3816,In_592,In_966);
nand U3817 (N_3817,In_958,In_781);
and U3818 (N_3818,In_37,In_758);
or U3819 (N_3819,In_862,In_342);
nand U3820 (N_3820,In_882,In_871);
and U3821 (N_3821,In_246,In_151);
nor U3822 (N_3822,In_652,In_728);
or U3823 (N_3823,In_86,In_823);
and U3824 (N_3824,In_402,In_86);
nor U3825 (N_3825,In_307,In_45);
nand U3826 (N_3826,In_63,In_640);
or U3827 (N_3827,In_732,In_726);
nor U3828 (N_3828,In_414,In_51);
nand U3829 (N_3829,In_323,In_452);
or U3830 (N_3830,In_445,In_297);
nor U3831 (N_3831,In_822,In_996);
or U3832 (N_3832,In_651,In_795);
and U3833 (N_3833,In_404,In_695);
nand U3834 (N_3834,In_238,In_201);
and U3835 (N_3835,In_613,In_624);
and U3836 (N_3836,In_696,In_775);
nor U3837 (N_3837,In_978,In_597);
or U3838 (N_3838,In_961,In_228);
or U3839 (N_3839,In_379,In_794);
and U3840 (N_3840,In_172,In_601);
nand U3841 (N_3841,In_675,In_103);
nor U3842 (N_3842,In_117,In_87);
nor U3843 (N_3843,In_807,In_866);
or U3844 (N_3844,In_272,In_74);
and U3845 (N_3845,In_425,In_815);
and U3846 (N_3846,In_200,In_294);
and U3847 (N_3847,In_318,In_214);
or U3848 (N_3848,In_276,In_752);
and U3849 (N_3849,In_825,In_841);
nor U3850 (N_3850,In_80,In_751);
or U3851 (N_3851,In_235,In_163);
and U3852 (N_3852,In_94,In_280);
and U3853 (N_3853,In_81,In_1);
and U3854 (N_3854,In_742,In_930);
and U3855 (N_3855,In_58,In_529);
nand U3856 (N_3856,In_657,In_368);
and U3857 (N_3857,In_70,In_714);
nand U3858 (N_3858,In_499,In_414);
nor U3859 (N_3859,In_126,In_196);
nand U3860 (N_3860,In_689,In_778);
and U3861 (N_3861,In_383,In_837);
nand U3862 (N_3862,In_451,In_594);
nand U3863 (N_3863,In_488,In_716);
and U3864 (N_3864,In_666,In_532);
nand U3865 (N_3865,In_411,In_661);
nor U3866 (N_3866,In_868,In_504);
nand U3867 (N_3867,In_146,In_437);
or U3868 (N_3868,In_752,In_67);
nand U3869 (N_3869,In_739,In_749);
xor U3870 (N_3870,In_451,In_500);
or U3871 (N_3871,In_696,In_81);
nor U3872 (N_3872,In_232,In_121);
nor U3873 (N_3873,In_664,In_874);
and U3874 (N_3874,In_831,In_259);
or U3875 (N_3875,In_827,In_531);
or U3876 (N_3876,In_211,In_77);
or U3877 (N_3877,In_634,In_55);
nor U3878 (N_3878,In_728,In_325);
and U3879 (N_3879,In_727,In_100);
xor U3880 (N_3880,In_653,In_801);
nand U3881 (N_3881,In_459,In_335);
and U3882 (N_3882,In_143,In_391);
or U3883 (N_3883,In_511,In_874);
nor U3884 (N_3884,In_382,In_56);
and U3885 (N_3885,In_749,In_203);
nor U3886 (N_3886,In_960,In_185);
or U3887 (N_3887,In_775,In_979);
and U3888 (N_3888,In_94,In_824);
and U3889 (N_3889,In_947,In_918);
nand U3890 (N_3890,In_222,In_624);
nand U3891 (N_3891,In_861,In_743);
nand U3892 (N_3892,In_90,In_697);
xor U3893 (N_3893,In_381,In_41);
nand U3894 (N_3894,In_289,In_259);
or U3895 (N_3895,In_43,In_845);
nand U3896 (N_3896,In_6,In_4);
nand U3897 (N_3897,In_753,In_638);
nor U3898 (N_3898,In_160,In_747);
nor U3899 (N_3899,In_119,In_870);
nand U3900 (N_3900,In_576,In_252);
and U3901 (N_3901,In_363,In_644);
nor U3902 (N_3902,In_640,In_799);
or U3903 (N_3903,In_68,In_564);
xnor U3904 (N_3904,In_281,In_936);
nand U3905 (N_3905,In_169,In_107);
and U3906 (N_3906,In_739,In_213);
or U3907 (N_3907,In_305,In_403);
nor U3908 (N_3908,In_67,In_347);
nand U3909 (N_3909,In_964,In_457);
nand U3910 (N_3910,In_558,In_644);
nand U3911 (N_3911,In_959,In_740);
or U3912 (N_3912,In_215,In_161);
nand U3913 (N_3913,In_209,In_351);
nor U3914 (N_3914,In_585,In_60);
or U3915 (N_3915,In_685,In_69);
or U3916 (N_3916,In_256,In_753);
nand U3917 (N_3917,In_452,In_201);
or U3918 (N_3918,In_355,In_17);
nand U3919 (N_3919,In_501,In_922);
or U3920 (N_3920,In_398,In_934);
nand U3921 (N_3921,In_106,In_58);
and U3922 (N_3922,In_17,In_124);
nand U3923 (N_3923,In_214,In_690);
nor U3924 (N_3924,In_702,In_34);
or U3925 (N_3925,In_138,In_675);
and U3926 (N_3926,In_954,In_99);
nand U3927 (N_3927,In_154,In_59);
and U3928 (N_3928,In_208,In_939);
and U3929 (N_3929,In_207,In_462);
or U3930 (N_3930,In_169,In_520);
nor U3931 (N_3931,In_478,In_634);
and U3932 (N_3932,In_633,In_973);
or U3933 (N_3933,In_970,In_109);
and U3934 (N_3934,In_331,In_74);
nand U3935 (N_3935,In_448,In_393);
nand U3936 (N_3936,In_626,In_950);
nor U3937 (N_3937,In_514,In_149);
nand U3938 (N_3938,In_313,In_949);
nor U3939 (N_3939,In_985,In_982);
nor U3940 (N_3940,In_352,In_758);
or U3941 (N_3941,In_450,In_56);
or U3942 (N_3942,In_463,In_432);
nor U3943 (N_3943,In_253,In_72);
and U3944 (N_3944,In_133,In_507);
or U3945 (N_3945,In_120,In_101);
nand U3946 (N_3946,In_51,In_794);
nand U3947 (N_3947,In_861,In_837);
and U3948 (N_3948,In_12,In_949);
nor U3949 (N_3949,In_473,In_31);
nand U3950 (N_3950,In_19,In_192);
and U3951 (N_3951,In_585,In_607);
nor U3952 (N_3952,In_629,In_926);
and U3953 (N_3953,In_120,In_254);
or U3954 (N_3954,In_139,In_873);
or U3955 (N_3955,In_879,In_946);
nand U3956 (N_3956,In_897,In_303);
nor U3957 (N_3957,In_691,In_642);
nand U3958 (N_3958,In_107,In_615);
nand U3959 (N_3959,In_857,In_216);
nor U3960 (N_3960,In_447,In_508);
and U3961 (N_3961,In_128,In_252);
nand U3962 (N_3962,In_690,In_253);
or U3963 (N_3963,In_939,In_946);
nor U3964 (N_3964,In_576,In_336);
and U3965 (N_3965,In_432,In_89);
nor U3966 (N_3966,In_938,In_130);
or U3967 (N_3967,In_397,In_45);
or U3968 (N_3968,In_304,In_289);
or U3969 (N_3969,In_396,In_142);
nand U3970 (N_3970,In_929,In_504);
and U3971 (N_3971,In_561,In_482);
nand U3972 (N_3972,In_560,In_790);
nor U3973 (N_3973,In_950,In_192);
nor U3974 (N_3974,In_671,In_130);
and U3975 (N_3975,In_335,In_994);
nand U3976 (N_3976,In_566,In_352);
nand U3977 (N_3977,In_910,In_476);
nor U3978 (N_3978,In_106,In_387);
nand U3979 (N_3979,In_89,In_877);
or U3980 (N_3980,In_546,In_254);
nor U3981 (N_3981,In_992,In_711);
nand U3982 (N_3982,In_464,In_738);
and U3983 (N_3983,In_291,In_40);
and U3984 (N_3984,In_397,In_931);
and U3985 (N_3985,In_28,In_371);
and U3986 (N_3986,In_584,In_813);
nor U3987 (N_3987,In_565,In_154);
and U3988 (N_3988,In_179,In_829);
nor U3989 (N_3989,In_480,In_555);
nor U3990 (N_3990,In_66,In_914);
nand U3991 (N_3991,In_260,In_865);
nand U3992 (N_3992,In_847,In_362);
nor U3993 (N_3993,In_764,In_702);
nand U3994 (N_3994,In_122,In_659);
and U3995 (N_3995,In_543,In_611);
nand U3996 (N_3996,In_603,In_958);
nor U3997 (N_3997,In_795,In_599);
and U3998 (N_3998,In_237,In_312);
and U3999 (N_3999,In_149,In_607);
or U4000 (N_4000,In_450,In_622);
nor U4001 (N_4001,In_118,In_61);
and U4002 (N_4002,In_785,In_762);
nor U4003 (N_4003,In_360,In_543);
nand U4004 (N_4004,In_290,In_83);
and U4005 (N_4005,In_119,In_774);
or U4006 (N_4006,In_558,In_880);
and U4007 (N_4007,In_172,In_681);
or U4008 (N_4008,In_753,In_884);
nor U4009 (N_4009,In_937,In_643);
or U4010 (N_4010,In_616,In_745);
nand U4011 (N_4011,In_369,In_489);
nand U4012 (N_4012,In_320,In_904);
or U4013 (N_4013,In_799,In_228);
nand U4014 (N_4014,In_936,In_666);
or U4015 (N_4015,In_884,In_401);
nor U4016 (N_4016,In_275,In_321);
nand U4017 (N_4017,In_413,In_984);
nand U4018 (N_4018,In_64,In_258);
xnor U4019 (N_4019,In_755,In_997);
or U4020 (N_4020,In_879,In_297);
nor U4021 (N_4021,In_898,In_571);
nand U4022 (N_4022,In_298,In_746);
nand U4023 (N_4023,In_219,In_559);
nand U4024 (N_4024,In_826,In_814);
nor U4025 (N_4025,In_73,In_872);
nand U4026 (N_4026,In_322,In_987);
or U4027 (N_4027,In_997,In_108);
and U4028 (N_4028,In_993,In_529);
nor U4029 (N_4029,In_906,In_514);
or U4030 (N_4030,In_181,In_835);
nand U4031 (N_4031,In_688,In_675);
or U4032 (N_4032,In_194,In_750);
or U4033 (N_4033,In_50,In_346);
xnor U4034 (N_4034,In_642,In_998);
and U4035 (N_4035,In_628,In_258);
and U4036 (N_4036,In_53,In_723);
nand U4037 (N_4037,In_301,In_25);
and U4038 (N_4038,In_919,In_309);
nor U4039 (N_4039,In_902,In_728);
nand U4040 (N_4040,In_724,In_701);
and U4041 (N_4041,In_845,In_597);
nor U4042 (N_4042,In_711,In_628);
nand U4043 (N_4043,In_690,In_8);
or U4044 (N_4044,In_127,In_385);
and U4045 (N_4045,In_878,In_14);
nand U4046 (N_4046,In_243,In_930);
nor U4047 (N_4047,In_627,In_276);
nand U4048 (N_4048,In_1,In_943);
and U4049 (N_4049,In_83,In_124);
nor U4050 (N_4050,In_472,In_687);
and U4051 (N_4051,In_490,In_353);
and U4052 (N_4052,In_721,In_244);
nand U4053 (N_4053,In_26,In_665);
nand U4054 (N_4054,In_3,In_692);
nor U4055 (N_4055,In_805,In_620);
nor U4056 (N_4056,In_959,In_651);
or U4057 (N_4057,In_27,In_858);
or U4058 (N_4058,In_619,In_112);
nor U4059 (N_4059,In_821,In_516);
or U4060 (N_4060,In_363,In_848);
nand U4061 (N_4061,In_142,In_950);
nor U4062 (N_4062,In_836,In_214);
and U4063 (N_4063,In_595,In_894);
nor U4064 (N_4064,In_731,In_402);
nor U4065 (N_4065,In_137,In_739);
nand U4066 (N_4066,In_374,In_762);
nand U4067 (N_4067,In_940,In_624);
and U4068 (N_4068,In_868,In_679);
and U4069 (N_4069,In_119,In_792);
and U4070 (N_4070,In_895,In_795);
nor U4071 (N_4071,In_232,In_698);
and U4072 (N_4072,In_368,In_722);
and U4073 (N_4073,In_507,In_328);
nor U4074 (N_4074,In_694,In_900);
nand U4075 (N_4075,In_196,In_92);
or U4076 (N_4076,In_93,In_590);
or U4077 (N_4077,In_910,In_682);
nor U4078 (N_4078,In_470,In_191);
and U4079 (N_4079,In_799,In_301);
nand U4080 (N_4080,In_990,In_944);
nand U4081 (N_4081,In_165,In_666);
and U4082 (N_4082,In_960,In_831);
and U4083 (N_4083,In_674,In_526);
nand U4084 (N_4084,In_210,In_428);
nor U4085 (N_4085,In_727,In_518);
nor U4086 (N_4086,In_577,In_354);
nand U4087 (N_4087,In_364,In_876);
or U4088 (N_4088,In_246,In_227);
and U4089 (N_4089,In_548,In_305);
nand U4090 (N_4090,In_981,In_83);
or U4091 (N_4091,In_275,In_722);
nand U4092 (N_4092,In_747,In_644);
nor U4093 (N_4093,In_119,In_191);
nand U4094 (N_4094,In_920,In_772);
or U4095 (N_4095,In_141,In_425);
or U4096 (N_4096,In_589,In_225);
or U4097 (N_4097,In_340,In_668);
nand U4098 (N_4098,In_784,In_802);
or U4099 (N_4099,In_865,In_722);
or U4100 (N_4100,In_866,In_751);
or U4101 (N_4101,In_560,In_360);
nor U4102 (N_4102,In_12,In_425);
nand U4103 (N_4103,In_597,In_401);
nand U4104 (N_4104,In_759,In_316);
nand U4105 (N_4105,In_683,In_514);
or U4106 (N_4106,In_530,In_918);
and U4107 (N_4107,In_688,In_553);
nor U4108 (N_4108,In_408,In_794);
or U4109 (N_4109,In_807,In_46);
nor U4110 (N_4110,In_723,In_777);
nand U4111 (N_4111,In_817,In_407);
or U4112 (N_4112,In_687,In_727);
nand U4113 (N_4113,In_107,In_159);
nand U4114 (N_4114,In_846,In_426);
nand U4115 (N_4115,In_43,In_292);
and U4116 (N_4116,In_169,In_593);
nand U4117 (N_4117,In_722,In_903);
nand U4118 (N_4118,In_231,In_500);
nor U4119 (N_4119,In_823,In_15);
and U4120 (N_4120,In_342,In_576);
nor U4121 (N_4121,In_78,In_806);
or U4122 (N_4122,In_725,In_467);
nor U4123 (N_4123,In_403,In_537);
and U4124 (N_4124,In_352,In_298);
and U4125 (N_4125,In_812,In_336);
nand U4126 (N_4126,In_680,In_865);
nand U4127 (N_4127,In_683,In_745);
and U4128 (N_4128,In_727,In_242);
or U4129 (N_4129,In_966,In_203);
and U4130 (N_4130,In_882,In_559);
or U4131 (N_4131,In_505,In_254);
or U4132 (N_4132,In_790,In_544);
nor U4133 (N_4133,In_40,In_559);
nand U4134 (N_4134,In_925,In_357);
or U4135 (N_4135,In_438,In_989);
nor U4136 (N_4136,In_901,In_128);
and U4137 (N_4137,In_873,In_10);
or U4138 (N_4138,In_494,In_364);
nor U4139 (N_4139,In_862,In_635);
or U4140 (N_4140,In_738,In_527);
nor U4141 (N_4141,In_272,In_923);
or U4142 (N_4142,In_556,In_207);
or U4143 (N_4143,In_370,In_817);
nor U4144 (N_4144,In_698,In_718);
nand U4145 (N_4145,In_507,In_55);
nand U4146 (N_4146,In_927,In_110);
nand U4147 (N_4147,In_533,In_747);
nand U4148 (N_4148,In_598,In_181);
and U4149 (N_4149,In_82,In_723);
and U4150 (N_4150,In_914,In_979);
and U4151 (N_4151,In_458,In_727);
nand U4152 (N_4152,In_767,In_133);
and U4153 (N_4153,In_956,In_726);
and U4154 (N_4154,In_427,In_465);
and U4155 (N_4155,In_989,In_43);
nand U4156 (N_4156,In_344,In_662);
nor U4157 (N_4157,In_146,In_89);
xnor U4158 (N_4158,In_579,In_585);
and U4159 (N_4159,In_283,In_478);
nand U4160 (N_4160,In_283,In_658);
nand U4161 (N_4161,In_901,In_690);
nand U4162 (N_4162,In_200,In_369);
nand U4163 (N_4163,In_540,In_328);
or U4164 (N_4164,In_361,In_216);
or U4165 (N_4165,In_75,In_664);
or U4166 (N_4166,In_241,In_565);
or U4167 (N_4167,In_966,In_404);
nand U4168 (N_4168,In_501,In_549);
nand U4169 (N_4169,In_922,In_231);
nor U4170 (N_4170,In_112,In_683);
or U4171 (N_4171,In_917,In_224);
and U4172 (N_4172,In_667,In_600);
nor U4173 (N_4173,In_692,In_583);
nand U4174 (N_4174,In_941,In_349);
nor U4175 (N_4175,In_896,In_830);
nand U4176 (N_4176,In_959,In_415);
and U4177 (N_4177,In_418,In_68);
nand U4178 (N_4178,In_608,In_2);
or U4179 (N_4179,In_18,In_912);
or U4180 (N_4180,In_855,In_863);
nand U4181 (N_4181,In_602,In_909);
nand U4182 (N_4182,In_45,In_330);
nand U4183 (N_4183,In_546,In_711);
and U4184 (N_4184,In_507,In_342);
nor U4185 (N_4185,In_475,In_24);
nand U4186 (N_4186,In_29,In_843);
nor U4187 (N_4187,In_179,In_75);
or U4188 (N_4188,In_816,In_534);
nor U4189 (N_4189,In_115,In_34);
or U4190 (N_4190,In_77,In_960);
nor U4191 (N_4191,In_279,In_521);
nor U4192 (N_4192,In_373,In_579);
nor U4193 (N_4193,In_966,In_220);
nor U4194 (N_4194,In_34,In_844);
or U4195 (N_4195,In_936,In_476);
nor U4196 (N_4196,In_284,In_900);
or U4197 (N_4197,In_615,In_225);
nor U4198 (N_4198,In_328,In_769);
or U4199 (N_4199,In_542,In_591);
nor U4200 (N_4200,In_928,In_509);
or U4201 (N_4201,In_268,In_9);
nor U4202 (N_4202,In_633,In_276);
nor U4203 (N_4203,In_447,In_989);
nor U4204 (N_4204,In_929,In_166);
nand U4205 (N_4205,In_129,In_407);
nor U4206 (N_4206,In_416,In_862);
or U4207 (N_4207,In_851,In_332);
and U4208 (N_4208,In_609,In_41);
nor U4209 (N_4209,In_116,In_975);
nand U4210 (N_4210,In_395,In_808);
nand U4211 (N_4211,In_328,In_7);
nor U4212 (N_4212,In_788,In_196);
nor U4213 (N_4213,In_408,In_100);
or U4214 (N_4214,In_28,In_103);
or U4215 (N_4215,In_154,In_278);
or U4216 (N_4216,In_607,In_455);
or U4217 (N_4217,In_500,In_331);
and U4218 (N_4218,In_190,In_965);
nor U4219 (N_4219,In_393,In_253);
nand U4220 (N_4220,In_598,In_147);
or U4221 (N_4221,In_969,In_432);
nor U4222 (N_4222,In_871,In_79);
nand U4223 (N_4223,In_827,In_808);
nor U4224 (N_4224,In_300,In_356);
nand U4225 (N_4225,In_815,In_469);
and U4226 (N_4226,In_11,In_341);
nor U4227 (N_4227,In_193,In_340);
or U4228 (N_4228,In_388,In_362);
nand U4229 (N_4229,In_35,In_879);
or U4230 (N_4230,In_858,In_279);
nand U4231 (N_4231,In_883,In_370);
and U4232 (N_4232,In_119,In_818);
nor U4233 (N_4233,In_728,In_205);
or U4234 (N_4234,In_741,In_280);
nand U4235 (N_4235,In_611,In_688);
nand U4236 (N_4236,In_526,In_438);
nor U4237 (N_4237,In_667,In_728);
xor U4238 (N_4238,In_154,In_147);
or U4239 (N_4239,In_14,In_935);
nand U4240 (N_4240,In_766,In_347);
nor U4241 (N_4241,In_901,In_160);
nand U4242 (N_4242,In_95,In_566);
nor U4243 (N_4243,In_991,In_352);
or U4244 (N_4244,In_977,In_849);
and U4245 (N_4245,In_720,In_733);
or U4246 (N_4246,In_718,In_915);
and U4247 (N_4247,In_465,In_385);
nand U4248 (N_4248,In_892,In_645);
nand U4249 (N_4249,In_106,In_738);
nor U4250 (N_4250,In_37,In_634);
nor U4251 (N_4251,In_846,In_673);
nand U4252 (N_4252,In_583,In_968);
and U4253 (N_4253,In_16,In_40);
nand U4254 (N_4254,In_88,In_228);
and U4255 (N_4255,In_488,In_154);
or U4256 (N_4256,In_514,In_251);
nand U4257 (N_4257,In_357,In_535);
or U4258 (N_4258,In_787,In_542);
or U4259 (N_4259,In_96,In_659);
or U4260 (N_4260,In_239,In_850);
nor U4261 (N_4261,In_835,In_882);
and U4262 (N_4262,In_910,In_320);
and U4263 (N_4263,In_355,In_313);
nor U4264 (N_4264,In_219,In_90);
or U4265 (N_4265,In_332,In_629);
nand U4266 (N_4266,In_294,In_675);
nand U4267 (N_4267,In_554,In_641);
and U4268 (N_4268,In_745,In_618);
and U4269 (N_4269,In_785,In_955);
and U4270 (N_4270,In_26,In_841);
nor U4271 (N_4271,In_874,In_439);
and U4272 (N_4272,In_860,In_934);
or U4273 (N_4273,In_31,In_972);
nor U4274 (N_4274,In_358,In_428);
nor U4275 (N_4275,In_858,In_320);
and U4276 (N_4276,In_833,In_53);
nand U4277 (N_4277,In_126,In_300);
nand U4278 (N_4278,In_594,In_944);
nand U4279 (N_4279,In_84,In_979);
nand U4280 (N_4280,In_105,In_243);
and U4281 (N_4281,In_674,In_45);
nand U4282 (N_4282,In_656,In_884);
nand U4283 (N_4283,In_35,In_11);
and U4284 (N_4284,In_544,In_746);
and U4285 (N_4285,In_92,In_36);
nand U4286 (N_4286,In_108,In_180);
or U4287 (N_4287,In_839,In_102);
or U4288 (N_4288,In_931,In_58);
and U4289 (N_4289,In_392,In_672);
or U4290 (N_4290,In_604,In_535);
nand U4291 (N_4291,In_818,In_843);
and U4292 (N_4292,In_228,In_693);
nor U4293 (N_4293,In_948,In_273);
nor U4294 (N_4294,In_128,In_45);
or U4295 (N_4295,In_327,In_578);
nand U4296 (N_4296,In_583,In_925);
nor U4297 (N_4297,In_242,In_540);
nor U4298 (N_4298,In_422,In_89);
nor U4299 (N_4299,In_469,In_947);
nand U4300 (N_4300,In_394,In_991);
nand U4301 (N_4301,In_939,In_264);
nor U4302 (N_4302,In_306,In_39);
nand U4303 (N_4303,In_350,In_781);
or U4304 (N_4304,In_190,In_205);
nor U4305 (N_4305,In_296,In_749);
and U4306 (N_4306,In_688,In_150);
nor U4307 (N_4307,In_140,In_530);
nand U4308 (N_4308,In_52,In_119);
nor U4309 (N_4309,In_967,In_54);
and U4310 (N_4310,In_789,In_941);
nor U4311 (N_4311,In_898,In_818);
nand U4312 (N_4312,In_152,In_862);
and U4313 (N_4313,In_120,In_67);
nand U4314 (N_4314,In_206,In_51);
nand U4315 (N_4315,In_858,In_893);
nor U4316 (N_4316,In_107,In_366);
nand U4317 (N_4317,In_564,In_128);
or U4318 (N_4318,In_436,In_386);
and U4319 (N_4319,In_525,In_865);
nand U4320 (N_4320,In_34,In_870);
and U4321 (N_4321,In_951,In_292);
nor U4322 (N_4322,In_451,In_912);
nand U4323 (N_4323,In_511,In_643);
or U4324 (N_4324,In_101,In_683);
nor U4325 (N_4325,In_291,In_45);
and U4326 (N_4326,In_392,In_751);
nand U4327 (N_4327,In_463,In_983);
nand U4328 (N_4328,In_801,In_597);
or U4329 (N_4329,In_592,In_451);
nor U4330 (N_4330,In_523,In_834);
nor U4331 (N_4331,In_957,In_736);
nor U4332 (N_4332,In_211,In_194);
nand U4333 (N_4333,In_311,In_478);
and U4334 (N_4334,In_336,In_390);
nand U4335 (N_4335,In_822,In_279);
nor U4336 (N_4336,In_402,In_350);
or U4337 (N_4337,In_348,In_675);
or U4338 (N_4338,In_549,In_880);
nand U4339 (N_4339,In_573,In_407);
nor U4340 (N_4340,In_970,In_926);
nor U4341 (N_4341,In_488,In_500);
or U4342 (N_4342,In_78,In_255);
or U4343 (N_4343,In_829,In_221);
nor U4344 (N_4344,In_734,In_43);
and U4345 (N_4345,In_297,In_26);
or U4346 (N_4346,In_627,In_686);
nand U4347 (N_4347,In_2,In_630);
nor U4348 (N_4348,In_878,In_947);
nor U4349 (N_4349,In_229,In_983);
nor U4350 (N_4350,In_996,In_0);
or U4351 (N_4351,In_663,In_162);
and U4352 (N_4352,In_993,In_680);
or U4353 (N_4353,In_248,In_856);
and U4354 (N_4354,In_990,In_254);
nor U4355 (N_4355,In_888,In_32);
and U4356 (N_4356,In_847,In_490);
and U4357 (N_4357,In_570,In_394);
and U4358 (N_4358,In_724,In_131);
and U4359 (N_4359,In_625,In_926);
nor U4360 (N_4360,In_246,In_908);
nand U4361 (N_4361,In_362,In_516);
or U4362 (N_4362,In_407,In_632);
nand U4363 (N_4363,In_752,In_655);
nand U4364 (N_4364,In_86,In_986);
nand U4365 (N_4365,In_256,In_139);
or U4366 (N_4366,In_604,In_360);
nor U4367 (N_4367,In_553,In_978);
and U4368 (N_4368,In_242,In_84);
nand U4369 (N_4369,In_509,In_63);
nor U4370 (N_4370,In_110,In_192);
nand U4371 (N_4371,In_655,In_564);
nand U4372 (N_4372,In_342,In_361);
nor U4373 (N_4373,In_668,In_542);
or U4374 (N_4374,In_389,In_167);
nor U4375 (N_4375,In_76,In_909);
nand U4376 (N_4376,In_999,In_461);
and U4377 (N_4377,In_732,In_720);
or U4378 (N_4378,In_474,In_391);
nor U4379 (N_4379,In_94,In_539);
nand U4380 (N_4380,In_643,In_131);
or U4381 (N_4381,In_581,In_911);
nand U4382 (N_4382,In_256,In_771);
and U4383 (N_4383,In_961,In_597);
nor U4384 (N_4384,In_845,In_790);
and U4385 (N_4385,In_859,In_402);
and U4386 (N_4386,In_161,In_806);
and U4387 (N_4387,In_152,In_761);
nand U4388 (N_4388,In_135,In_748);
nand U4389 (N_4389,In_655,In_950);
nand U4390 (N_4390,In_329,In_278);
and U4391 (N_4391,In_182,In_487);
or U4392 (N_4392,In_959,In_807);
and U4393 (N_4393,In_686,In_234);
or U4394 (N_4394,In_181,In_511);
nor U4395 (N_4395,In_236,In_607);
and U4396 (N_4396,In_745,In_853);
nor U4397 (N_4397,In_381,In_783);
and U4398 (N_4398,In_378,In_245);
and U4399 (N_4399,In_140,In_671);
nor U4400 (N_4400,In_94,In_525);
nor U4401 (N_4401,In_225,In_976);
and U4402 (N_4402,In_651,In_412);
nand U4403 (N_4403,In_984,In_382);
nor U4404 (N_4404,In_555,In_550);
and U4405 (N_4405,In_264,In_823);
nor U4406 (N_4406,In_626,In_82);
or U4407 (N_4407,In_48,In_808);
nor U4408 (N_4408,In_850,In_19);
or U4409 (N_4409,In_470,In_558);
and U4410 (N_4410,In_388,In_973);
nor U4411 (N_4411,In_236,In_174);
nand U4412 (N_4412,In_560,In_161);
nand U4413 (N_4413,In_781,In_984);
and U4414 (N_4414,In_558,In_30);
nand U4415 (N_4415,In_74,In_572);
or U4416 (N_4416,In_155,In_884);
nand U4417 (N_4417,In_240,In_647);
or U4418 (N_4418,In_535,In_514);
or U4419 (N_4419,In_833,In_555);
nor U4420 (N_4420,In_766,In_120);
nor U4421 (N_4421,In_943,In_604);
and U4422 (N_4422,In_325,In_789);
nand U4423 (N_4423,In_235,In_956);
or U4424 (N_4424,In_558,In_21);
or U4425 (N_4425,In_367,In_280);
or U4426 (N_4426,In_567,In_865);
or U4427 (N_4427,In_525,In_756);
or U4428 (N_4428,In_718,In_10);
or U4429 (N_4429,In_356,In_381);
or U4430 (N_4430,In_58,In_472);
nand U4431 (N_4431,In_177,In_759);
and U4432 (N_4432,In_340,In_277);
or U4433 (N_4433,In_214,In_538);
nand U4434 (N_4434,In_397,In_874);
nor U4435 (N_4435,In_899,In_721);
or U4436 (N_4436,In_92,In_986);
and U4437 (N_4437,In_333,In_455);
nor U4438 (N_4438,In_305,In_34);
and U4439 (N_4439,In_807,In_1);
and U4440 (N_4440,In_500,In_223);
and U4441 (N_4441,In_202,In_186);
and U4442 (N_4442,In_37,In_193);
and U4443 (N_4443,In_688,In_71);
or U4444 (N_4444,In_20,In_60);
and U4445 (N_4445,In_449,In_670);
nand U4446 (N_4446,In_84,In_207);
and U4447 (N_4447,In_611,In_937);
or U4448 (N_4448,In_975,In_655);
nand U4449 (N_4449,In_330,In_421);
and U4450 (N_4450,In_909,In_823);
nand U4451 (N_4451,In_196,In_351);
nor U4452 (N_4452,In_784,In_741);
nand U4453 (N_4453,In_242,In_252);
and U4454 (N_4454,In_495,In_103);
nor U4455 (N_4455,In_458,In_271);
and U4456 (N_4456,In_337,In_175);
nand U4457 (N_4457,In_265,In_967);
nand U4458 (N_4458,In_842,In_715);
and U4459 (N_4459,In_790,In_289);
or U4460 (N_4460,In_536,In_322);
and U4461 (N_4461,In_544,In_705);
nor U4462 (N_4462,In_591,In_109);
or U4463 (N_4463,In_470,In_902);
nand U4464 (N_4464,In_678,In_631);
or U4465 (N_4465,In_195,In_332);
nor U4466 (N_4466,In_294,In_623);
and U4467 (N_4467,In_212,In_711);
or U4468 (N_4468,In_14,In_521);
or U4469 (N_4469,In_616,In_714);
nor U4470 (N_4470,In_325,In_261);
nand U4471 (N_4471,In_649,In_144);
nor U4472 (N_4472,In_131,In_125);
nor U4473 (N_4473,In_869,In_544);
or U4474 (N_4474,In_209,In_382);
nor U4475 (N_4475,In_323,In_878);
or U4476 (N_4476,In_611,In_63);
or U4477 (N_4477,In_106,In_19);
nand U4478 (N_4478,In_848,In_353);
or U4479 (N_4479,In_911,In_115);
and U4480 (N_4480,In_591,In_722);
nand U4481 (N_4481,In_235,In_647);
nor U4482 (N_4482,In_484,In_904);
and U4483 (N_4483,In_299,In_91);
nor U4484 (N_4484,In_733,In_860);
or U4485 (N_4485,In_543,In_623);
and U4486 (N_4486,In_469,In_212);
and U4487 (N_4487,In_400,In_502);
or U4488 (N_4488,In_659,In_674);
and U4489 (N_4489,In_596,In_184);
nand U4490 (N_4490,In_542,In_178);
nand U4491 (N_4491,In_283,In_754);
or U4492 (N_4492,In_342,In_753);
xor U4493 (N_4493,In_81,In_819);
nor U4494 (N_4494,In_615,In_808);
or U4495 (N_4495,In_132,In_145);
and U4496 (N_4496,In_160,In_968);
nor U4497 (N_4497,In_161,In_752);
and U4498 (N_4498,In_158,In_391);
or U4499 (N_4499,In_625,In_323);
or U4500 (N_4500,In_586,In_954);
and U4501 (N_4501,In_852,In_773);
and U4502 (N_4502,In_909,In_805);
nor U4503 (N_4503,In_595,In_874);
and U4504 (N_4504,In_357,In_155);
or U4505 (N_4505,In_257,In_278);
or U4506 (N_4506,In_215,In_534);
or U4507 (N_4507,In_287,In_302);
and U4508 (N_4508,In_410,In_300);
or U4509 (N_4509,In_348,In_100);
and U4510 (N_4510,In_168,In_515);
nand U4511 (N_4511,In_76,In_341);
nor U4512 (N_4512,In_992,In_405);
and U4513 (N_4513,In_276,In_292);
or U4514 (N_4514,In_72,In_782);
nor U4515 (N_4515,In_930,In_460);
nand U4516 (N_4516,In_206,In_183);
or U4517 (N_4517,In_532,In_412);
and U4518 (N_4518,In_948,In_435);
nand U4519 (N_4519,In_562,In_745);
nor U4520 (N_4520,In_490,In_797);
nand U4521 (N_4521,In_404,In_125);
nor U4522 (N_4522,In_249,In_334);
and U4523 (N_4523,In_898,In_10);
nand U4524 (N_4524,In_952,In_914);
nand U4525 (N_4525,In_478,In_592);
nor U4526 (N_4526,In_165,In_304);
or U4527 (N_4527,In_116,In_281);
and U4528 (N_4528,In_943,In_401);
and U4529 (N_4529,In_967,In_490);
or U4530 (N_4530,In_52,In_397);
nand U4531 (N_4531,In_908,In_257);
and U4532 (N_4532,In_515,In_241);
nor U4533 (N_4533,In_486,In_815);
nor U4534 (N_4534,In_429,In_640);
or U4535 (N_4535,In_114,In_497);
and U4536 (N_4536,In_392,In_308);
nor U4537 (N_4537,In_997,In_515);
nor U4538 (N_4538,In_523,In_386);
nor U4539 (N_4539,In_784,In_125);
nand U4540 (N_4540,In_995,In_651);
or U4541 (N_4541,In_650,In_466);
nor U4542 (N_4542,In_747,In_867);
and U4543 (N_4543,In_501,In_86);
and U4544 (N_4544,In_853,In_675);
nand U4545 (N_4545,In_226,In_475);
or U4546 (N_4546,In_995,In_869);
or U4547 (N_4547,In_519,In_181);
nand U4548 (N_4548,In_863,In_796);
nor U4549 (N_4549,In_939,In_299);
nand U4550 (N_4550,In_416,In_158);
nor U4551 (N_4551,In_810,In_294);
and U4552 (N_4552,In_733,In_248);
and U4553 (N_4553,In_645,In_593);
nor U4554 (N_4554,In_644,In_271);
and U4555 (N_4555,In_576,In_394);
or U4556 (N_4556,In_398,In_636);
nand U4557 (N_4557,In_928,In_264);
or U4558 (N_4558,In_730,In_475);
and U4559 (N_4559,In_361,In_710);
nor U4560 (N_4560,In_605,In_508);
or U4561 (N_4561,In_109,In_910);
nand U4562 (N_4562,In_784,In_637);
and U4563 (N_4563,In_721,In_229);
and U4564 (N_4564,In_990,In_955);
or U4565 (N_4565,In_872,In_742);
or U4566 (N_4566,In_224,In_942);
nand U4567 (N_4567,In_175,In_556);
nor U4568 (N_4568,In_84,In_888);
nand U4569 (N_4569,In_86,In_872);
nand U4570 (N_4570,In_968,In_299);
nor U4571 (N_4571,In_911,In_297);
or U4572 (N_4572,In_580,In_233);
or U4573 (N_4573,In_631,In_332);
nor U4574 (N_4574,In_990,In_711);
nand U4575 (N_4575,In_350,In_922);
or U4576 (N_4576,In_490,In_10);
and U4577 (N_4577,In_427,In_352);
nor U4578 (N_4578,In_313,In_66);
nor U4579 (N_4579,In_497,In_263);
or U4580 (N_4580,In_497,In_291);
or U4581 (N_4581,In_0,In_886);
nand U4582 (N_4582,In_281,In_700);
nand U4583 (N_4583,In_84,In_198);
and U4584 (N_4584,In_905,In_533);
and U4585 (N_4585,In_905,In_529);
nor U4586 (N_4586,In_93,In_220);
nand U4587 (N_4587,In_140,In_518);
or U4588 (N_4588,In_416,In_464);
nor U4589 (N_4589,In_589,In_351);
nor U4590 (N_4590,In_157,In_952);
xor U4591 (N_4591,In_248,In_879);
nor U4592 (N_4592,In_85,In_695);
nand U4593 (N_4593,In_641,In_491);
nand U4594 (N_4594,In_96,In_188);
nand U4595 (N_4595,In_409,In_646);
or U4596 (N_4596,In_544,In_200);
nand U4597 (N_4597,In_600,In_440);
and U4598 (N_4598,In_835,In_720);
nor U4599 (N_4599,In_478,In_541);
nor U4600 (N_4600,In_847,In_648);
nand U4601 (N_4601,In_67,In_24);
nand U4602 (N_4602,In_830,In_171);
and U4603 (N_4603,In_77,In_582);
nor U4604 (N_4604,In_474,In_404);
nand U4605 (N_4605,In_22,In_969);
and U4606 (N_4606,In_928,In_687);
and U4607 (N_4607,In_180,In_248);
xnor U4608 (N_4608,In_504,In_233);
nand U4609 (N_4609,In_217,In_831);
nand U4610 (N_4610,In_65,In_407);
and U4611 (N_4611,In_78,In_960);
or U4612 (N_4612,In_173,In_819);
nor U4613 (N_4613,In_871,In_106);
nand U4614 (N_4614,In_260,In_795);
or U4615 (N_4615,In_960,In_165);
nor U4616 (N_4616,In_65,In_668);
or U4617 (N_4617,In_756,In_342);
and U4618 (N_4618,In_107,In_779);
and U4619 (N_4619,In_312,In_272);
nand U4620 (N_4620,In_764,In_729);
nand U4621 (N_4621,In_435,In_735);
nor U4622 (N_4622,In_716,In_450);
nor U4623 (N_4623,In_111,In_540);
nor U4624 (N_4624,In_822,In_76);
or U4625 (N_4625,In_86,In_408);
and U4626 (N_4626,In_642,In_469);
or U4627 (N_4627,In_641,In_117);
or U4628 (N_4628,In_35,In_285);
and U4629 (N_4629,In_257,In_420);
or U4630 (N_4630,In_135,In_743);
and U4631 (N_4631,In_564,In_785);
nor U4632 (N_4632,In_461,In_611);
or U4633 (N_4633,In_663,In_573);
and U4634 (N_4634,In_231,In_341);
nor U4635 (N_4635,In_961,In_686);
nor U4636 (N_4636,In_867,In_281);
nand U4637 (N_4637,In_179,In_814);
nand U4638 (N_4638,In_544,In_390);
nand U4639 (N_4639,In_373,In_883);
and U4640 (N_4640,In_857,In_195);
nand U4641 (N_4641,In_956,In_246);
or U4642 (N_4642,In_982,In_820);
and U4643 (N_4643,In_657,In_791);
nand U4644 (N_4644,In_985,In_966);
nand U4645 (N_4645,In_409,In_310);
or U4646 (N_4646,In_506,In_120);
nor U4647 (N_4647,In_519,In_745);
or U4648 (N_4648,In_416,In_829);
nor U4649 (N_4649,In_48,In_540);
nor U4650 (N_4650,In_635,In_716);
nand U4651 (N_4651,In_751,In_181);
nand U4652 (N_4652,In_512,In_700);
nor U4653 (N_4653,In_753,In_465);
nand U4654 (N_4654,In_192,In_734);
or U4655 (N_4655,In_104,In_954);
or U4656 (N_4656,In_393,In_469);
and U4657 (N_4657,In_902,In_347);
and U4658 (N_4658,In_645,In_223);
nand U4659 (N_4659,In_208,In_884);
and U4660 (N_4660,In_877,In_470);
nand U4661 (N_4661,In_462,In_903);
nor U4662 (N_4662,In_420,In_90);
and U4663 (N_4663,In_138,In_233);
nand U4664 (N_4664,In_80,In_384);
and U4665 (N_4665,In_20,In_391);
nor U4666 (N_4666,In_1,In_559);
xor U4667 (N_4667,In_252,In_454);
nand U4668 (N_4668,In_513,In_344);
nand U4669 (N_4669,In_961,In_848);
xnor U4670 (N_4670,In_739,In_153);
or U4671 (N_4671,In_211,In_529);
and U4672 (N_4672,In_627,In_720);
nand U4673 (N_4673,In_779,In_768);
and U4674 (N_4674,In_680,In_588);
nor U4675 (N_4675,In_827,In_404);
and U4676 (N_4676,In_941,In_11);
nor U4677 (N_4677,In_908,In_593);
and U4678 (N_4678,In_566,In_459);
nor U4679 (N_4679,In_520,In_80);
nand U4680 (N_4680,In_226,In_616);
or U4681 (N_4681,In_577,In_606);
or U4682 (N_4682,In_151,In_595);
nand U4683 (N_4683,In_88,In_48);
nand U4684 (N_4684,In_395,In_360);
nand U4685 (N_4685,In_585,In_336);
nand U4686 (N_4686,In_575,In_635);
and U4687 (N_4687,In_963,In_947);
nor U4688 (N_4688,In_221,In_803);
nor U4689 (N_4689,In_116,In_787);
nand U4690 (N_4690,In_307,In_83);
nor U4691 (N_4691,In_575,In_578);
or U4692 (N_4692,In_885,In_124);
or U4693 (N_4693,In_592,In_164);
nor U4694 (N_4694,In_590,In_169);
nand U4695 (N_4695,In_37,In_373);
or U4696 (N_4696,In_396,In_72);
and U4697 (N_4697,In_261,In_407);
and U4698 (N_4698,In_410,In_853);
nor U4699 (N_4699,In_744,In_443);
nor U4700 (N_4700,In_390,In_93);
nand U4701 (N_4701,In_495,In_805);
nor U4702 (N_4702,In_946,In_274);
nor U4703 (N_4703,In_870,In_377);
nand U4704 (N_4704,In_622,In_700);
nand U4705 (N_4705,In_280,In_274);
and U4706 (N_4706,In_913,In_411);
nand U4707 (N_4707,In_351,In_903);
nor U4708 (N_4708,In_365,In_974);
or U4709 (N_4709,In_479,In_870);
nor U4710 (N_4710,In_970,In_382);
nor U4711 (N_4711,In_586,In_543);
and U4712 (N_4712,In_891,In_507);
nand U4713 (N_4713,In_295,In_994);
and U4714 (N_4714,In_207,In_629);
or U4715 (N_4715,In_375,In_538);
nor U4716 (N_4716,In_707,In_692);
nor U4717 (N_4717,In_22,In_315);
and U4718 (N_4718,In_152,In_878);
and U4719 (N_4719,In_3,In_78);
nand U4720 (N_4720,In_612,In_659);
and U4721 (N_4721,In_925,In_350);
nor U4722 (N_4722,In_736,In_322);
nand U4723 (N_4723,In_36,In_740);
or U4724 (N_4724,In_39,In_748);
nor U4725 (N_4725,In_733,In_308);
nand U4726 (N_4726,In_527,In_115);
and U4727 (N_4727,In_1,In_204);
nor U4728 (N_4728,In_783,In_337);
nand U4729 (N_4729,In_147,In_115);
or U4730 (N_4730,In_157,In_166);
and U4731 (N_4731,In_424,In_237);
nand U4732 (N_4732,In_308,In_896);
nor U4733 (N_4733,In_992,In_622);
and U4734 (N_4734,In_675,In_284);
nor U4735 (N_4735,In_887,In_825);
nor U4736 (N_4736,In_122,In_546);
and U4737 (N_4737,In_160,In_480);
or U4738 (N_4738,In_463,In_424);
and U4739 (N_4739,In_663,In_133);
xor U4740 (N_4740,In_435,In_459);
nand U4741 (N_4741,In_226,In_130);
nor U4742 (N_4742,In_564,In_300);
or U4743 (N_4743,In_276,In_535);
and U4744 (N_4744,In_408,In_24);
nor U4745 (N_4745,In_330,In_720);
nor U4746 (N_4746,In_795,In_187);
nand U4747 (N_4747,In_641,In_826);
or U4748 (N_4748,In_748,In_422);
nand U4749 (N_4749,In_436,In_740);
nor U4750 (N_4750,In_43,In_573);
or U4751 (N_4751,In_169,In_697);
nor U4752 (N_4752,In_515,In_648);
nand U4753 (N_4753,In_967,In_553);
nand U4754 (N_4754,In_762,In_981);
nor U4755 (N_4755,In_992,In_149);
and U4756 (N_4756,In_521,In_83);
nor U4757 (N_4757,In_62,In_195);
or U4758 (N_4758,In_375,In_740);
nor U4759 (N_4759,In_557,In_584);
and U4760 (N_4760,In_492,In_790);
nand U4761 (N_4761,In_898,In_269);
or U4762 (N_4762,In_817,In_514);
nand U4763 (N_4763,In_468,In_68);
or U4764 (N_4764,In_923,In_751);
and U4765 (N_4765,In_947,In_268);
and U4766 (N_4766,In_87,In_784);
and U4767 (N_4767,In_143,In_742);
nor U4768 (N_4768,In_510,In_781);
and U4769 (N_4769,In_748,In_957);
nor U4770 (N_4770,In_28,In_796);
nor U4771 (N_4771,In_996,In_13);
nand U4772 (N_4772,In_758,In_833);
nand U4773 (N_4773,In_105,In_132);
nand U4774 (N_4774,In_345,In_833);
and U4775 (N_4775,In_919,In_191);
nand U4776 (N_4776,In_270,In_140);
or U4777 (N_4777,In_371,In_727);
and U4778 (N_4778,In_296,In_893);
nor U4779 (N_4779,In_718,In_325);
and U4780 (N_4780,In_639,In_796);
and U4781 (N_4781,In_492,In_143);
or U4782 (N_4782,In_902,In_406);
or U4783 (N_4783,In_694,In_992);
nor U4784 (N_4784,In_974,In_494);
xnor U4785 (N_4785,In_455,In_728);
nor U4786 (N_4786,In_735,In_676);
nand U4787 (N_4787,In_233,In_586);
nand U4788 (N_4788,In_569,In_629);
and U4789 (N_4789,In_36,In_428);
nand U4790 (N_4790,In_687,In_806);
or U4791 (N_4791,In_287,In_626);
xor U4792 (N_4792,In_464,In_84);
or U4793 (N_4793,In_397,In_519);
nand U4794 (N_4794,In_853,In_183);
nand U4795 (N_4795,In_545,In_74);
nand U4796 (N_4796,In_709,In_902);
nor U4797 (N_4797,In_654,In_12);
and U4798 (N_4798,In_79,In_598);
nand U4799 (N_4799,In_642,In_989);
nor U4800 (N_4800,In_754,In_362);
or U4801 (N_4801,In_877,In_909);
or U4802 (N_4802,In_861,In_278);
nor U4803 (N_4803,In_334,In_105);
or U4804 (N_4804,In_180,In_666);
and U4805 (N_4805,In_369,In_975);
nor U4806 (N_4806,In_443,In_963);
nand U4807 (N_4807,In_9,In_823);
nor U4808 (N_4808,In_833,In_43);
and U4809 (N_4809,In_819,In_312);
nor U4810 (N_4810,In_500,In_504);
and U4811 (N_4811,In_670,In_182);
or U4812 (N_4812,In_988,In_901);
nor U4813 (N_4813,In_330,In_925);
nor U4814 (N_4814,In_8,In_171);
nand U4815 (N_4815,In_9,In_100);
and U4816 (N_4816,In_164,In_79);
nor U4817 (N_4817,In_280,In_579);
or U4818 (N_4818,In_655,In_230);
and U4819 (N_4819,In_73,In_363);
or U4820 (N_4820,In_150,In_792);
nor U4821 (N_4821,In_480,In_791);
or U4822 (N_4822,In_284,In_130);
and U4823 (N_4823,In_454,In_742);
nand U4824 (N_4824,In_412,In_919);
nand U4825 (N_4825,In_164,In_366);
or U4826 (N_4826,In_887,In_568);
and U4827 (N_4827,In_964,In_520);
nand U4828 (N_4828,In_542,In_76);
or U4829 (N_4829,In_326,In_605);
and U4830 (N_4830,In_834,In_568);
and U4831 (N_4831,In_148,In_156);
nand U4832 (N_4832,In_530,In_655);
nor U4833 (N_4833,In_214,In_71);
nand U4834 (N_4834,In_125,In_260);
or U4835 (N_4835,In_611,In_227);
nor U4836 (N_4836,In_671,In_480);
nor U4837 (N_4837,In_770,In_849);
and U4838 (N_4838,In_368,In_110);
nand U4839 (N_4839,In_499,In_476);
xor U4840 (N_4840,In_199,In_279);
nand U4841 (N_4841,In_887,In_830);
nand U4842 (N_4842,In_971,In_170);
and U4843 (N_4843,In_507,In_44);
nand U4844 (N_4844,In_337,In_335);
and U4845 (N_4845,In_5,In_504);
and U4846 (N_4846,In_346,In_732);
or U4847 (N_4847,In_548,In_139);
and U4848 (N_4848,In_572,In_901);
nor U4849 (N_4849,In_590,In_503);
nor U4850 (N_4850,In_914,In_88);
nor U4851 (N_4851,In_771,In_519);
or U4852 (N_4852,In_524,In_93);
xnor U4853 (N_4853,In_231,In_534);
nor U4854 (N_4854,In_197,In_975);
nor U4855 (N_4855,In_928,In_309);
and U4856 (N_4856,In_48,In_553);
nor U4857 (N_4857,In_602,In_151);
or U4858 (N_4858,In_829,In_150);
nand U4859 (N_4859,In_16,In_332);
nand U4860 (N_4860,In_74,In_47);
nand U4861 (N_4861,In_778,In_190);
and U4862 (N_4862,In_857,In_725);
or U4863 (N_4863,In_128,In_9);
nor U4864 (N_4864,In_566,In_992);
nor U4865 (N_4865,In_934,In_997);
nor U4866 (N_4866,In_629,In_525);
nand U4867 (N_4867,In_241,In_939);
and U4868 (N_4868,In_400,In_986);
nand U4869 (N_4869,In_226,In_993);
nor U4870 (N_4870,In_890,In_276);
nor U4871 (N_4871,In_532,In_739);
nand U4872 (N_4872,In_224,In_442);
nand U4873 (N_4873,In_809,In_88);
nor U4874 (N_4874,In_501,In_430);
xnor U4875 (N_4875,In_342,In_310);
nand U4876 (N_4876,In_470,In_603);
and U4877 (N_4877,In_950,In_889);
nand U4878 (N_4878,In_514,In_167);
or U4879 (N_4879,In_683,In_128);
or U4880 (N_4880,In_505,In_54);
nand U4881 (N_4881,In_859,In_37);
nor U4882 (N_4882,In_377,In_12);
and U4883 (N_4883,In_535,In_130);
nor U4884 (N_4884,In_650,In_646);
nor U4885 (N_4885,In_466,In_250);
or U4886 (N_4886,In_315,In_506);
nor U4887 (N_4887,In_385,In_877);
or U4888 (N_4888,In_532,In_346);
or U4889 (N_4889,In_269,In_914);
xor U4890 (N_4890,In_521,In_550);
nor U4891 (N_4891,In_840,In_854);
nor U4892 (N_4892,In_908,In_836);
nand U4893 (N_4893,In_447,In_613);
or U4894 (N_4894,In_457,In_155);
nand U4895 (N_4895,In_262,In_814);
nor U4896 (N_4896,In_920,In_950);
nand U4897 (N_4897,In_380,In_981);
nor U4898 (N_4898,In_773,In_305);
and U4899 (N_4899,In_713,In_494);
or U4900 (N_4900,In_830,In_112);
nand U4901 (N_4901,In_579,In_742);
nor U4902 (N_4902,In_376,In_979);
nor U4903 (N_4903,In_288,In_165);
and U4904 (N_4904,In_589,In_988);
and U4905 (N_4905,In_383,In_829);
or U4906 (N_4906,In_416,In_354);
nor U4907 (N_4907,In_923,In_666);
and U4908 (N_4908,In_567,In_462);
nand U4909 (N_4909,In_352,In_749);
and U4910 (N_4910,In_592,In_254);
and U4911 (N_4911,In_122,In_373);
or U4912 (N_4912,In_84,In_573);
nor U4913 (N_4913,In_397,In_989);
or U4914 (N_4914,In_155,In_172);
nand U4915 (N_4915,In_305,In_30);
or U4916 (N_4916,In_250,In_811);
and U4917 (N_4917,In_174,In_808);
and U4918 (N_4918,In_931,In_742);
or U4919 (N_4919,In_608,In_603);
and U4920 (N_4920,In_896,In_442);
or U4921 (N_4921,In_891,In_786);
and U4922 (N_4922,In_752,In_257);
nand U4923 (N_4923,In_730,In_483);
and U4924 (N_4924,In_141,In_339);
or U4925 (N_4925,In_530,In_702);
or U4926 (N_4926,In_469,In_198);
and U4927 (N_4927,In_755,In_573);
nor U4928 (N_4928,In_703,In_221);
nor U4929 (N_4929,In_950,In_293);
nor U4930 (N_4930,In_681,In_509);
and U4931 (N_4931,In_323,In_369);
nor U4932 (N_4932,In_299,In_795);
nor U4933 (N_4933,In_649,In_419);
xnor U4934 (N_4934,In_752,In_390);
or U4935 (N_4935,In_327,In_967);
or U4936 (N_4936,In_125,In_185);
nand U4937 (N_4937,In_124,In_190);
xor U4938 (N_4938,In_330,In_445);
nor U4939 (N_4939,In_386,In_362);
and U4940 (N_4940,In_740,In_882);
and U4941 (N_4941,In_785,In_854);
and U4942 (N_4942,In_98,In_571);
nand U4943 (N_4943,In_107,In_468);
nor U4944 (N_4944,In_51,In_311);
and U4945 (N_4945,In_893,In_762);
nor U4946 (N_4946,In_839,In_343);
or U4947 (N_4947,In_837,In_33);
nor U4948 (N_4948,In_405,In_169);
nor U4949 (N_4949,In_845,In_346);
and U4950 (N_4950,In_509,In_530);
and U4951 (N_4951,In_87,In_499);
and U4952 (N_4952,In_221,In_421);
or U4953 (N_4953,In_377,In_700);
nand U4954 (N_4954,In_208,In_555);
and U4955 (N_4955,In_755,In_887);
and U4956 (N_4956,In_335,In_568);
nor U4957 (N_4957,In_519,In_212);
and U4958 (N_4958,In_227,In_550);
or U4959 (N_4959,In_976,In_83);
and U4960 (N_4960,In_567,In_819);
nand U4961 (N_4961,In_626,In_172);
nand U4962 (N_4962,In_671,In_866);
nor U4963 (N_4963,In_350,In_291);
nor U4964 (N_4964,In_182,In_109);
nand U4965 (N_4965,In_96,In_683);
and U4966 (N_4966,In_918,In_418);
and U4967 (N_4967,In_49,In_817);
or U4968 (N_4968,In_466,In_648);
or U4969 (N_4969,In_405,In_307);
and U4970 (N_4970,In_312,In_126);
nor U4971 (N_4971,In_369,In_187);
nor U4972 (N_4972,In_734,In_673);
nand U4973 (N_4973,In_201,In_428);
nor U4974 (N_4974,In_555,In_702);
and U4975 (N_4975,In_653,In_154);
nand U4976 (N_4976,In_733,In_937);
nand U4977 (N_4977,In_865,In_755);
or U4978 (N_4978,In_414,In_193);
nand U4979 (N_4979,In_583,In_390);
nor U4980 (N_4980,In_653,In_451);
nand U4981 (N_4981,In_889,In_688);
and U4982 (N_4982,In_278,In_389);
nor U4983 (N_4983,In_342,In_621);
nand U4984 (N_4984,In_191,In_477);
and U4985 (N_4985,In_996,In_541);
nor U4986 (N_4986,In_529,In_377);
nor U4987 (N_4987,In_955,In_326);
and U4988 (N_4988,In_59,In_82);
or U4989 (N_4989,In_946,In_768);
nand U4990 (N_4990,In_553,In_709);
nor U4991 (N_4991,In_307,In_100);
nand U4992 (N_4992,In_723,In_921);
and U4993 (N_4993,In_205,In_696);
or U4994 (N_4994,In_900,In_60);
nor U4995 (N_4995,In_632,In_483);
nand U4996 (N_4996,In_684,In_781);
or U4997 (N_4997,In_979,In_712);
and U4998 (N_4998,In_648,In_338);
and U4999 (N_4999,In_565,In_859);
nand U5000 (N_5000,N_444,N_1117);
nor U5001 (N_5001,N_372,N_1192);
and U5002 (N_5002,N_4054,N_4492);
or U5003 (N_5003,N_4770,N_3186);
and U5004 (N_5004,N_3163,N_1486);
and U5005 (N_5005,N_1844,N_151);
and U5006 (N_5006,N_2263,N_2524);
nand U5007 (N_5007,N_1735,N_1739);
nor U5008 (N_5008,N_982,N_3395);
and U5009 (N_5009,N_4013,N_1618);
nand U5010 (N_5010,N_3685,N_2493);
nand U5011 (N_5011,N_2227,N_899);
or U5012 (N_5012,N_2710,N_3076);
nor U5013 (N_5013,N_2570,N_2839);
or U5014 (N_5014,N_2682,N_2612);
nand U5015 (N_5015,N_3023,N_4474);
nor U5016 (N_5016,N_686,N_1639);
or U5017 (N_5017,N_506,N_4023);
nand U5018 (N_5018,N_2985,N_1129);
nand U5019 (N_5019,N_486,N_36);
nor U5020 (N_5020,N_4070,N_4445);
and U5021 (N_5021,N_1080,N_4015);
nand U5022 (N_5022,N_4508,N_4617);
nand U5023 (N_5023,N_3248,N_1855);
or U5024 (N_5024,N_3993,N_2108);
and U5025 (N_5025,N_1598,N_1343);
or U5026 (N_5026,N_605,N_1632);
and U5027 (N_5027,N_503,N_4484);
and U5028 (N_5028,N_1877,N_3058);
nand U5029 (N_5029,N_4560,N_4343);
or U5030 (N_5030,N_4181,N_3630);
nand U5031 (N_5031,N_2064,N_139);
nor U5032 (N_5032,N_3373,N_4465);
nor U5033 (N_5033,N_1969,N_1744);
nor U5034 (N_5034,N_3224,N_1407);
nand U5035 (N_5035,N_2453,N_3897);
or U5036 (N_5036,N_2684,N_642);
nand U5037 (N_5037,N_1549,N_1303);
or U5038 (N_5038,N_2473,N_3736);
nor U5039 (N_5039,N_2865,N_1966);
nor U5040 (N_5040,N_821,N_1714);
or U5041 (N_5041,N_4435,N_534);
nand U5042 (N_5042,N_3497,N_2260);
or U5043 (N_5043,N_1792,N_3220);
nor U5044 (N_5044,N_4548,N_4965);
or U5045 (N_5045,N_1937,N_2954);
nor U5046 (N_5046,N_790,N_2430);
and U5047 (N_5047,N_3940,N_857);
or U5048 (N_5048,N_2491,N_970);
nand U5049 (N_5049,N_1317,N_2097);
or U5050 (N_5050,N_3892,N_1910);
and U5051 (N_5051,N_4934,N_634);
or U5052 (N_5052,N_2550,N_4165);
nand U5053 (N_5053,N_255,N_4220);
and U5054 (N_5054,N_2480,N_1124);
and U5055 (N_5055,N_4340,N_907);
nand U5056 (N_5056,N_3251,N_1933);
nand U5057 (N_5057,N_1110,N_3860);
nand U5058 (N_5058,N_3250,N_4736);
and U5059 (N_5059,N_4229,N_3692);
nand U5060 (N_5060,N_657,N_2349);
and U5061 (N_5061,N_3672,N_2271);
nand U5062 (N_5062,N_1690,N_2777);
nor U5063 (N_5063,N_3558,N_2114);
nor U5064 (N_5064,N_4392,N_4576);
nor U5065 (N_5065,N_3164,N_3124);
nand U5066 (N_5066,N_1372,N_2992);
and U5067 (N_5067,N_4931,N_904);
nor U5068 (N_5068,N_505,N_4602);
nor U5069 (N_5069,N_636,N_3763);
nor U5070 (N_5070,N_1912,N_3934);
and U5071 (N_5071,N_2462,N_1298);
or U5072 (N_5072,N_1740,N_2551);
nand U5073 (N_5073,N_2672,N_524);
and U5074 (N_5074,N_1016,N_4946);
and U5075 (N_5075,N_2334,N_1929);
nor U5076 (N_5076,N_720,N_3286);
or U5077 (N_5077,N_2737,N_2871);
and U5078 (N_5078,N_2003,N_2258);
or U5079 (N_5079,N_4802,N_4101);
and U5080 (N_5080,N_2369,N_4851);
nor U5081 (N_5081,N_4417,N_2747);
nor U5082 (N_5082,N_2160,N_1069);
nor U5083 (N_5083,N_3389,N_3211);
and U5084 (N_5084,N_1767,N_2885);
nor U5085 (N_5085,N_1351,N_3204);
or U5086 (N_5086,N_2537,N_4914);
nand U5087 (N_5087,N_3208,N_173);
or U5088 (N_5088,N_1798,N_1000);
or U5089 (N_5089,N_3380,N_23);
or U5090 (N_5090,N_3840,N_253);
and U5091 (N_5091,N_1199,N_3863);
or U5092 (N_5092,N_4145,N_2866);
nand U5093 (N_5093,N_2047,N_203);
nor U5094 (N_5094,N_4859,N_4519);
or U5095 (N_5095,N_4098,N_4144);
and U5096 (N_5096,N_3241,N_575);
or U5097 (N_5097,N_1946,N_752);
or U5098 (N_5098,N_2891,N_4709);
nand U5099 (N_5099,N_4655,N_1224);
or U5100 (N_5100,N_206,N_1930);
nand U5101 (N_5101,N_3138,N_1770);
or U5102 (N_5102,N_4948,N_3219);
nor U5103 (N_5103,N_3240,N_1120);
and U5104 (N_5104,N_83,N_263);
or U5105 (N_5105,N_1736,N_3107);
or U5106 (N_5106,N_383,N_4459);
or U5107 (N_5107,N_3571,N_2649);
nand U5108 (N_5108,N_2020,N_1516);
and U5109 (N_5109,N_4500,N_822);
nor U5110 (N_5110,N_861,N_2039);
nor U5111 (N_5111,N_3661,N_727);
and U5112 (N_5112,N_4955,N_525);
nor U5113 (N_5113,N_1007,N_4318);
nor U5114 (N_5114,N_1834,N_1132);
nor U5115 (N_5115,N_1480,N_4885);
and U5116 (N_5116,N_4678,N_4276);
nor U5117 (N_5117,N_3991,N_682);
or U5118 (N_5118,N_2997,N_3668);
nor U5119 (N_5119,N_146,N_14);
nand U5120 (N_5120,N_4926,N_239);
nor U5121 (N_5121,N_1524,N_1887);
and U5122 (N_5122,N_3605,N_1630);
and U5123 (N_5123,N_377,N_1608);
nor U5124 (N_5124,N_4712,N_1920);
nor U5125 (N_5125,N_449,N_554);
and U5126 (N_5126,N_4158,N_1315);
nand U5127 (N_5127,N_1496,N_2613);
and U5128 (N_5128,N_2446,N_2341);
and U5129 (N_5129,N_660,N_4745);
nor U5130 (N_5130,N_4415,N_1021);
nor U5131 (N_5131,N_2938,N_1779);
nand U5132 (N_5132,N_4938,N_4426);
or U5133 (N_5133,N_334,N_1533);
nand U5134 (N_5134,N_2956,N_2439);
xnor U5135 (N_5135,N_4669,N_4811);
nor U5136 (N_5136,N_1745,N_4947);
xnor U5137 (N_5137,N_3575,N_4640);
and U5138 (N_5138,N_2784,N_1253);
or U5139 (N_5139,N_679,N_1698);
or U5140 (N_5140,N_1200,N_322);
nand U5141 (N_5141,N_2195,N_2496);
nand U5142 (N_5142,N_3399,N_853);
and U5143 (N_5143,N_4383,N_1824);
or U5144 (N_5144,N_1170,N_1577);
or U5145 (N_5145,N_1626,N_2045);
and U5146 (N_5146,N_1164,N_1741);
or U5147 (N_5147,N_467,N_2397);
nor U5148 (N_5148,N_90,N_1126);
nor U5149 (N_5149,N_2536,N_1391);
nand U5150 (N_5150,N_3742,N_2478);
nand U5151 (N_5151,N_2847,N_2266);
nor U5152 (N_5152,N_2224,N_1842);
nand U5153 (N_5153,N_3818,N_3213);
nand U5154 (N_5154,N_4431,N_4992);
or U5155 (N_5155,N_4226,N_91);
and U5156 (N_5156,N_72,N_20);
and U5157 (N_5157,N_3748,N_3858);
nor U5158 (N_5158,N_1028,N_2025);
or U5159 (N_5159,N_4516,N_1430);
nand U5160 (N_5160,N_885,N_1364);
or U5161 (N_5161,N_3889,N_3313);
or U5162 (N_5162,N_1325,N_748);
and U5163 (N_5163,N_1288,N_60);
nand U5164 (N_5164,N_3063,N_2301);
nor U5165 (N_5165,N_665,N_3724);
or U5166 (N_5166,N_1870,N_1456);
nand U5167 (N_5167,N_4333,N_4803);
nand U5168 (N_5168,N_2075,N_2786);
and U5169 (N_5169,N_4214,N_2983);
nand U5170 (N_5170,N_4533,N_2772);
nor U5171 (N_5171,N_4607,N_2256);
nor U5172 (N_5172,N_456,N_1528);
and U5173 (N_5173,N_3882,N_3546);
or U5174 (N_5174,N_4530,N_1014);
nand U5175 (N_5175,N_2245,N_3223);
nor U5176 (N_5176,N_3830,N_4471);
nor U5177 (N_5177,N_3712,N_1167);
nand U5178 (N_5178,N_2925,N_2782);
or U5179 (N_5179,N_788,N_3236);
and U5180 (N_5180,N_1070,N_569);
and U5181 (N_5181,N_1783,N_2624);
nor U5182 (N_5182,N_2166,N_939);
nor U5183 (N_5183,N_1894,N_1888);
and U5184 (N_5184,N_1086,N_2506);
nand U5185 (N_5185,N_1241,N_145);
or U5186 (N_5186,N_71,N_520);
nand U5187 (N_5187,N_4048,N_2987);
nor U5188 (N_5188,N_3357,N_722);
and U5189 (N_5189,N_3841,N_4767);
or U5190 (N_5190,N_4882,N_3664);
or U5191 (N_5191,N_1780,N_823);
nand U5192 (N_5192,N_2519,N_883);
or U5193 (N_5193,N_4105,N_2094);
nand U5194 (N_5194,N_4238,N_2947);
nor U5195 (N_5195,N_3310,N_1475);
nor U5196 (N_5196,N_4826,N_3682);
and U5197 (N_5197,N_1096,N_4843);
nand U5198 (N_5198,N_4986,N_556);
nor U5199 (N_5199,N_1296,N_4470);
or U5200 (N_5200,N_3962,N_3606);
and U5201 (N_5201,N_2741,N_2633);
nand U5202 (N_5202,N_2530,N_990);
and U5203 (N_5203,N_3235,N_1039);
and U5204 (N_5204,N_1077,N_3658);
or U5205 (N_5205,N_1062,N_840);
and U5206 (N_5206,N_1902,N_188);
nor U5207 (N_5207,N_479,N_726);
and U5208 (N_5208,N_3548,N_3227);
and U5209 (N_5209,N_2518,N_931);
or U5210 (N_5210,N_1708,N_4361);
or U5211 (N_5211,N_4962,N_851);
and U5212 (N_5212,N_2356,N_3083);
nand U5213 (N_5213,N_4246,N_1355);
and U5214 (N_5214,N_3465,N_3690);
nor U5215 (N_5215,N_379,N_2126);
nand U5216 (N_5216,N_1316,N_3677);
nor U5217 (N_5217,N_954,N_2474);
nand U5218 (N_5218,N_4805,N_1468);
nor U5219 (N_5219,N_4132,N_3563);
or U5220 (N_5220,N_2599,N_1172);
nand U5221 (N_5221,N_2238,N_4814);
nand U5222 (N_5222,N_412,N_1071);
nor U5223 (N_5223,N_3833,N_4266);
or U5224 (N_5224,N_542,N_1243);
xnor U5225 (N_5225,N_2667,N_1018);
or U5226 (N_5226,N_4960,N_2350);
or U5227 (N_5227,N_599,N_3469);
nand U5228 (N_5228,N_3887,N_419);
and U5229 (N_5229,N_2348,N_4375);
and U5230 (N_5230,N_3280,N_3092);
and U5231 (N_5231,N_314,N_46);
and U5232 (N_5232,N_149,N_2372);
nand U5233 (N_5233,N_3955,N_442);
or U5234 (N_5234,N_4171,N_528);
nand U5235 (N_5235,N_1293,N_409);
or U5236 (N_5236,N_956,N_2509);
or U5237 (N_5237,N_4020,N_1793);
or U5238 (N_5238,N_4439,N_4644);
nor U5239 (N_5239,N_2981,N_3266);
and U5240 (N_5240,N_2713,N_154);
nor U5241 (N_5241,N_889,N_3614);
or U5242 (N_5242,N_342,N_4487);
and U5243 (N_5243,N_3303,N_652);
nand U5244 (N_5244,N_4553,N_1410);
nor U5245 (N_5245,N_714,N_877);
nand U5246 (N_5246,N_2444,N_3354);
or U5247 (N_5247,N_610,N_737);
and U5248 (N_5248,N_4968,N_4604);
nand U5249 (N_5249,N_3120,N_2610);
and U5250 (N_5250,N_4209,N_4497);
nand U5251 (N_5251,N_1811,N_4094);
or U5252 (N_5252,N_356,N_1350);
nor U5253 (N_5253,N_1665,N_2054);
nor U5254 (N_5254,N_3191,N_3845);
or U5255 (N_5255,N_2803,N_296);
and U5256 (N_5256,N_4033,N_3823);
or U5257 (N_5257,N_2225,N_1279);
or U5258 (N_5258,N_3147,N_1890);
nand U5259 (N_5259,N_3511,N_4215);
or U5260 (N_5260,N_220,N_1619);
or U5261 (N_5261,N_4577,N_3330);
and U5262 (N_5262,N_3988,N_1271);
or U5263 (N_5263,N_4322,N_277);
or U5264 (N_5264,N_3564,N_4893);
nand U5265 (N_5265,N_2948,N_2659);
nor U5266 (N_5266,N_1839,N_2124);
or U5267 (N_5267,N_186,N_3372);
and U5268 (N_5268,N_3527,N_4026);
nand U5269 (N_5269,N_275,N_219);
and U5270 (N_5270,N_3306,N_4664);
nand U5271 (N_5271,N_2823,N_3838);
and U5272 (N_5272,N_4073,N_300);
and U5273 (N_5273,N_3526,N_1130);
nor U5274 (N_5274,N_517,N_2587);
or U5275 (N_5275,N_4772,N_4583);
nand U5276 (N_5276,N_4835,N_2525);
and U5277 (N_5277,N_3435,N_3275);
xor U5278 (N_5278,N_3181,N_4526);
or U5279 (N_5279,N_3461,N_3206);
xor U5280 (N_5280,N_4536,N_308);
nand U5281 (N_5281,N_2147,N_629);
nor U5282 (N_5282,N_1936,N_4909);
nand U5283 (N_5283,N_3479,N_3944);
nand U5284 (N_5284,N_1586,N_2130);
xnor U5285 (N_5285,N_457,N_4385);
or U5286 (N_5286,N_2877,N_4099);
or U5287 (N_5287,N_4989,N_1712);
or U5288 (N_5288,N_204,N_4100);
nand U5289 (N_5289,N_2693,N_3570);
nor U5290 (N_5290,N_4278,N_2297);
nor U5291 (N_5291,N_2377,N_2978);
and U5292 (N_5292,N_1076,N_4956);
and U5293 (N_5293,N_349,N_3488);
nor U5294 (N_5294,N_2156,N_2151);
nor U5295 (N_5295,N_2016,N_1587);
nand U5296 (N_5296,N_1155,N_3801);
or U5297 (N_5297,N_150,N_3369);
nand U5298 (N_5298,N_4045,N_2230);
and U5299 (N_5299,N_2766,N_2416);
nor U5300 (N_5300,N_1173,N_2785);
nor U5301 (N_5301,N_2799,N_62);
and U5302 (N_5302,N_288,N_2109);
and U5303 (N_5303,N_1585,N_2205);
and U5304 (N_5304,N_3390,N_3103);
and U5305 (N_5305,N_4812,N_3339);
nand U5306 (N_5306,N_1319,N_2869);
or U5307 (N_5307,N_75,N_3169);
and U5308 (N_5308,N_4705,N_2084);
nor U5309 (N_5309,N_3591,N_1385);
and U5310 (N_5310,N_4394,N_411);
nand U5311 (N_5311,N_4999,N_633);
nor U5312 (N_5312,N_2457,N_656);
and U5313 (N_5313,N_1038,N_3981);
nand U5314 (N_5314,N_4566,N_1747);
nor U5315 (N_5315,N_3604,N_4346);
or U5316 (N_5316,N_4206,N_704);
nor U5317 (N_5317,N_2485,N_2870);
or U5318 (N_5318,N_18,N_465);
nand U5319 (N_5319,N_2332,N_1924);
or U5320 (N_5320,N_654,N_1852);
and U5321 (N_5321,N_1334,N_3466);
and U5322 (N_5322,N_4550,N_2744);
nand U5323 (N_5323,N_998,N_3464);
or U5324 (N_5324,N_1254,N_1345);
and U5325 (N_5325,N_2723,N_3542);
nor U5326 (N_5326,N_3550,N_933);
or U5327 (N_5327,N_3289,N_2059);
nor U5328 (N_5328,N_3761,N_3803);
nand U5329 (N_5329,N_1008,N_4258);
and U5330 (N_5330,N_557,N_3589);
and U5331 (N_5331,N_261,N_4155);
nand U5332 (N_5332,N_4510,N_1653);
nand U5333 (N_5333,N_4028,N_1649);
or U5334 (N_5334,N_2021,N_3738);
or U5335 (N_5335,N_155,N_1127);
and U5336 (N_5336,N_1651,N_2361);
nand U5337 (N_5337,N_974,N_4599);
and U5338 (N_5338,N_3540,N_2759);
or U5339 (N_5339,N_2597,N_3336);
nand U5340 (N_5340,N_1928,N_3855);
nor U5341 (N_5341,N_107,N_1221);
and U5342 (N_5342,N_4320,N_3709);
nand U5343 (N_5343,N_2774,N_2176);
or U5344 (N_5344,N_713,N_3018);
nor U5345 (N_5345,N_3210,N_600);
nor U5346 (N_5346,N_2223,N_3068);
or U5347 (N_5347,N_1664,N_1203);
nand U5348 (N_5348,N_4696,N_214);
or U5349 (N_5349,N_3997,N_319);
or U5350 (N_5350,N_2635,N_655);
nand U5351 (N_5351,N_1274,N_271);
or U5352 (N_5352,N_3077,N_3758);
or U5353 (N_5353,N_2917,N_1416);
nand U5354 (N_5354,N_2831,N_371);
and U5355 (N_5355,N_1571,N_4614);
or U5356 (N_5356,N_1359,N_2492);
nor U5357 (N_5357,N_1846,N_1948);
nand U5358 (N_5358,N_2449,N_2140);
nand U5359 (N_5359,N_4891,N_3381);
or U5360 (N_5360,N_4674,N_984);
or U5361 (N_5361,N_1988,N_496);
nor U5362 (N_5362,N_4954,N_2152);
nor U5363 (N_5363,N_3295,N_1575);
nor U5364 (N_5364,N_133,N_2378);
and U5365 (N_5365,N_2296,N_2555);
and U5366 (N_5366,N_1283,N_3481);
or U5367 (N_5367,N_800,N_3839);
or U5368 (N_5368,N_2526,N_4286);
and U5369 (N_5369,N_4725,N_3300);
and U5370 (N_5370,N_473,N_3975);
nand U5371 (N_5371,N_3704,N_4507);
nor U5372 (N_5372,N_1300,N_2508);
nor U5373 (N_5373,N_290,N_1118);
nand U5374 (N_5374,N_2190,N_4555);
and U5375 (N_5375,N_3999,N_3462);
or U5376 (N_5376,N_3960,N_1799);
nand U5377 (N_5377,N_2502,N_1593);
xnor U5378 (N_5378,N_4032,N_1573);
and U5379 (N_5379,N_41,N_4252);
nor U5380 (N_5380,N_1926,N_847);
nand U5381 (N_5381,N_2005,N_1160);
or U5382 (N_5382,N_3739,N_2820);
or U5383 (N_5383,N_1449,N_160);
nand U5384 (N_5384,N_3653,N_17);
and U5385 (N_5385,N_1092,N_3291);
nand U5386 (N_5386,N_4239,N_2058);
and U5387 (N_5387,N_4866,N_3276);
or U5388 (N_5388,N_2791,N_4869);
and U5389 (N_5389,N_795,N_1610);
nor U5390 (N_5390,N_2712,N_3420);
and U5391 (N_5391,N_3128,N_462);
nor U5392 (N_5392,N_819,N_1204);
or U5393 (N_5393,N_3190,N_3544);
nor U5394 (N_5394,N_3750,N_4865);
or U5395 (N_5395,N_4088,N_2619);
or U5396 (N_5396,N_1976,N_1764);
or U5397 (N_5397,N_2796,N_2608);
nor U5398 (N_5398,N_67,N_2117);
or U5399 (N_5399,N_59,N_2155);
nor U5400 (N_5400,N_2862,N_241);
nand U5401 (N_5401,N_4633,N_1578);
or U5402 (N_5402,N_3859,N_3322);
nand U5403 (N_5403,N_3700,N_3885);
or U5404 (N_5404,N_4029,N_4845);
nand U5405 (N_5405,N_3894,N_3360);
or U5406 (N_5406,N_744,N_4634);
and U5407 (N_5407,N_421,N_1089);
and U5408 (N_5408,N_1668,N_381);
nand U5409 (N_5409,N_4842,N_2330);
nor U5410 (N_5410,N_389,N_3207);
or U5411 (N_5411,N_3167,N_2445);
nand U5412 (N_5412,N_4227,N_4213);
or U5413 (N_5413,N_208,N_2584);
nor U5414 (N_5414,N_135,N_3556);
and U5415 (N_5415,N_981,N_3710);
nand U5416 (N_5416,N_4858,N_2211);
or U5417 (N_5417,N_3057,N_3132);
nor U5418 (N_5418,N_724,N_4959);
or U5419 (N_5419,N_3467,N_594);
nand U5420 (N_5420,N_985,N_690);
nand U5421 (N_5421,N_3886,N_212);
and U5422 (N_5422,N_967,N_2670);
or U5423 (N_5423,N_3601,N_3829);
nand U5424 (N_5424,N_1542,N_1817);
nor U5425 (N_5425,N_1900,N_1399);
nor U5426 (N_5426,N_3269,N_2000);
and U5427 (N_5427,N_3099,N_2314);
and U5428 (N_5428,N_2251,N_4328);
or U5429 (N_5429,N_3890,N_519);
nand U5430 (N_5430,N_3939,N_305);
or U5431 (N_5431,N_2973,N_4060);
nor U5432 (N_5432,N_4037,N_10);
nand U5433 (N_5433,N_4034,N_649);
and U5434 (N_5434,N_695,N_390);
or U5435 (N_5435,N_2364,N_3054);
and U5436 (N_5436,N_4224,N_4436);
nand U5437 (N_5437,N_687,N_3179);
nor U5438 (N_5438,N_2407,N_875);
and U5439 (N_5439,N_4850,N_838);
nand U5440 (N_5440,N_1037,N_2320);
or U5441 (N_5441,N_4222,N_639);
and U5442 (N_5442,N_3945,N_490);
or U5443 (N_5443,N_1795,N_4758);
or U5444 (N_5444,N_1252,N_454);
nor U5445 (N_5445,N_2215,N_1153);
or U5446 (N_5446,N_3875,N_3490);
or U5447 (N_5447,N_363,N_3644);
nand U5448 (N_5448,N_1255,N_1382);
and U5449 (N_5449,N_2734,N_1590);
nor U5450 (N_5450,N_1017,N_4190);
or U5451 (N_5451,N_2110,N_1574);
nand U5452 (N_5452,N_427,N_3493);
nand U5453 (N_5453,N_2809,N_3331);
and U5454 (N_5454,N_2007,N_3559);
nor U5455 (N_5455,N_4639,N_3194);
or U5456 (N_5456,N_2770,N_2437);
or U5457 (N_5457,N_4801,N_4317);
or U5458 (N_5458,N_958,N_4513);
nand U5459 (N_5459,N_750,N_2062);
nor U5460 (N_5460,N_404,N_4069);
nand U5461 (N_5461,N_3162,N_3309);
and U5462 (N_5462,N_258,N_2669);
nor U5463 (N_5463,N_925,N_4661);
nand U5464 (N_5464,N_1613,N_105);
or U5465 (N_5465,N_1511,N_3543);
nor U5466 (N_5466,N_38,N_2347);
or U5467 (N_5467,N_307,N_3880);
nor U5468 (N_5468,N_1581,N_1065);
and U5469 (N_5469,N_1318,N_3611);
and U5470 (N_5470,N_611,N_969);
or U5471 (N_5471,N_3701,N_2235);
and U5472 (N_5472,N_3359,N_297);
nand U5473 (N_5473,N_3911,N_3495);
and U5474 (N_5474,N_2136,N_3424);
nand U5475 (N_5475,N_2685,N_3429);
nand U5476 (N_5476,N_3531,N_1907);
and U5477 (N_5477,N_3032,N_2467);
nand U5478 (N_5478,N_3024,N_2528);
nor U5479 (N_5479,N_4730,N_2312);
or U5480 (N_5480,N_191,N_4575);
nor U5481 (N_5481,N_347,N_1191);
nand U5482 (N_5482,N_3470,N_4864);
nor U5483 (N_5483,N_2501,N_3102);
and U5484 (N_5484,N_92,N_3595);
nor U5485 (N_5485,N_4440,N_2585);
and U5486 (N_5486,N_1050,N_927);
and U5487 (N_5487,N_3626,N_2452);
and U5488 (N_5488,N_3528,N_812);
and U5489 (N_5489,N_4387,N_1436);
and U5490 (N_5490,N_1683,N_4977);
nor U5491 (N_5491,N_3505,N_286);
nand U5492 (N_5492,N_645,N_3974);
nor U5493 (N_5493,N_710,N_1195);
and U5494 (N_5494,N_4641,N_4489);
or U5495 (N_5495,N_2466,N_4189);
nor U5496 (N_5496,N_1339,N_1519);
and U5497 (N_5497,N_4254,N_4442);
and U5498 (N_5498,N_2929,N_493);
nor U5499 (N_5499,N_1370,N_1344);
nor U5500 (N_5500,N_549,N_4460);
and U5501 (N_5501,N_337,N_3699);
and U5502 (N_5502,N_4559,N_4515);
nand U5503 (N_5503,N_1433,N_3687);
and U5504 (N_5504,N_2505,N_489);
nand U5505 (N_5505,N_986,N_328);
and U5506 (N_5506,N_612,N_3349);
nor U5507 (N_5507,N_382,N_3480);
or U5508 (N_5508,N_1211,N_2776);
nand U5509 (N_5509,N_2639,N_2708);
nor U5510 (N_5510,N_3854,N_2658);
or U5511 (N_5511,N_1876,N_1663);
or U5512 (N_5512,N_2958,N_2887);
nand U5513 (N_5513,N_1403,N_2834);
nand U5514 (N_5514,N_1384,N_576);
nand U5515 (N_5515,N_230,N_3176);
and U5516 (N_5516,N_1368,N_1159);
and U5517 (N_5517,N_4787,N_3089);
nor U5518 (N_5518,N_2923,N_2798);
and U5519 (N_5519,N_622,N_3686);
nand U5520 (N_5520,N_2515,N_3284);
nor U5521 (N_5521,N_1506,N_201);
nor U5522 (N_5522,N_908,N_3517);
and U5523 (N_5523,N_1108,N_4355);
nor U5524 (N_5524,N_4233,N_4594);
nor U5525 (N_5525,N_589,N_1045);
or U5526 (N_5526,N_2135,N_3101);
nand U5527 (N_5527,N_2222,N_1242);
or U5528 (N_5528,N_515,N_581);
nand U5529 (N_5529,N_4126,N_4403);
nor U5530 (N_5530,N_1095,N_4827);
nand U5531 (N_5531,N_3499,N_4702);
nor U5532 (N_5532,N_1617,N_86);
and U5533 (N_5533,N_2792,N_1457);
or U5534 (N_5534,N_910,N_4870);
nor U5535 (N_5535,N_4081,N_1908);
nor U5536 (N_5536,N_3452,N_1947);
nand U5537 (N_5537,N_3351,N_1987);
or U5538 (N_5538,N_4592,N_4097);
and U5539 (N_5539,N_4211,N_1205);
nor U5540 (N_5540,N_2797,N_3971);
nand U5541 (N_5541,N_1941,N_1927);
nor U5542 (N_5542,N_4315,N_2636);
and U5543 (N_5543,N_1588,N_3016);
and U5544 (N_5544,N_3009,N_1371);
and U5545 (N_5545,N_1423,N_4244);
and U5546 (N_5546,N_4953,N_2647);
or U5547 (N_5547,N_4283,N_4253);
and U5548 (N_5548,N_207,N_1748);
nand U5549 (N_5549,N_2728,N_2512);
and U5550 (N_5550,N_539,N_1526);
and U5551 (N_5551,N_1105,N_2595);
nor U5552 (N_5552,N_4593,N_1361);
nand U5553 (N_5553,N_4425,N_966);
nand U5554 (N_5554,N_1951,N_1629);
or U5555 (N_5555,N_3192,N_164);
nor U5556 (N_5556,N_3258,N_4648);
nor U5557 (N_5557,N_4228,N_429);
nand U5558 (N_5558,N_4062,N_2050);
or U5559 (N_5559,N_85,N_1463);
and U5560 (N_5560,N_2226,N_2720);
and U5561 (N_5561,N_4464,N_4567);
nand U5562 (N_5562,N_2254,N_3702);
nor U5563 (N_5563,N_760,N_3970);
and U5564 (N_5564,N_791,N_2856);
nor U5565 (N_5565,N_616,N_3426);
or U5566 (N_5566,N_134,N_1067);
and U5567 (N_5567,N_794,N_1725);
and U5568 (N_5568,N_4950,N_769);
and U5569 (N_5569,N_1671,N_1097);
and U5570 (N_5570,N_1494,N_1087);
or U5571 (N_5571,N_4963,N_2666);
xnor U5572 (N_5572,N_4907,N_623);
nor U5573 (N_5573,N_1843,N_384);
nor U5574 (N_5574,N_2873,N_4653);
nand U5575 (N_5575,N_232,N_3486);
nand U5576 (N_5576,N_4915,N_1025);
and U5577 (N_5577,N_1544,N_352);
and U5578 (N_5578,N_181,N_2221);
and U5579 (N_5579,N_2032,N_4540);
nor U5580 (N_5580,N_1450,N_4535);
xnor U5581 (N_5581,N_4797,N_3274);
or U5582 (N_5582,N_1766,N_2030);
nand U5583 (N_5583,N_2168,N_3002);
and U5584 (N_5584,N_614,N_4349);
or U5585 (N_5585,N_2122,N_3247);
or U5586 (N_5586,N_1721,N_310);
and U5587 (N_5587,N_4297,N_2511);
nor U5588 (N_5588,N_285,N_138);
nand U5589 (N_5589,N_2357,N_4719);
or U5590 (N_5590,N_2589,N_3904);
nand U5591 (N_5591,N_2403,N_2008);
nor U5592 (N_5592,N_2678,N_1352);
nand U5593 (N_5593,N_4872,N_335);
or U5594 (N_5594,N_3098,N_3121);
nand U5595 (N_5595,N_193,N_4857);
or U5596 (N_5596,N_4332,N_4076);
or U5597 (N_5597,N_61,N_4585);
and U5598 (N_5598,N_132,N_3364);
nand U5599 (N_5599,N_4491,N_1709);
or U5600 (N_5600,N_2717,N_3114);
or U5601 (N_5601,N_1667,N_1994);
and U5602 (N_5602,N_3583,N_706);
or U5603 (N_5603,N_3329,N_2464);
or U5604 (N_5604,N_451,N_3916);
and U5605 (N_5605,N_804,N_4262);
and U5606 (N_5606,N_3387,N_2620);
nor U5607 (N_5607,N_4057,N_1232);
nand U5608 (N_5608,N_3652,N_4486);
and U5609 (N_5609,N_4223,N_3819);
or U5610 (N_5610,N_4973,N_354);
and U5611 (N_5611,N_1658,N_3406);
nor U5612 (N_5612,N_2494,N_2427);
nor U5613 (N_5613,N_1104,N_3643);
nand U5614 (N_5614,N_2232,N_3954);
and U5615 (N_5615,N_1848,N_601);
nand U5616 (N_5616,N_4853,N_1309);
nor U5617 (N_5617,N_688,N_3573);
nor U5618 (N_5618,N_3625,N_30);
xor U5619 (N_5619,N_292,N_2295);
or U5620 (N_5620,N_2704,N_4849);
and U5621 (N_5621,N_4140,N_1723);
nor U5622 (N_5622,N_360,N_2541);
nor U5623 (N_5623,N_1459,N_1705);
nor U5624 (N_5624,N_4469,N_1801);
or U5625 (N_5625,N_735,N_3534);
or U5626 (N_5626,N_474,N_4518);
nand U5627 (N_5627,N_2841,N_4207);
nand U5628 (N_5628,N_1791,N_2617);
or U5629 (N_5629,N_625,N_619);
nand U5630 (N_5630,N_3134,N_1061);
nand U5631 (N_5631,N_4447,N_2857);
or U5632 (N_5632,N_2889,N_2687);
and U5633 (N_5633,N_2788,N_1850);
or U5634 (N_5634,N_1538,N_77);
and U5635 (N_5635,N_1595,N_2413);
and U5636 (N_5636,N_2127,N_4879);
nor U5637 (N_5637,N_3202,N_237);
nor U5638 (N_5638,N_84,N_365);
nor U5639 (N_5639,N_2833,N_698);
and U5640 (N_5640,N_890,N_119);
or U5641 (N_5641,N_2252,N_4546);
and U5642 (N_5642,N_793,N_1991);
or U5643 (N_5643,N_751,N_3753);
nor U5644 (N_5644,N_2346,N_1443);
nand U5645 (N_5645,N_2034,N_2998);
or U5646 (N_5646,N_2688,N_1942);
and U5647 (N_5647,N_414,N_957);
nand U5648 (N_5648,N_2479,N_596);
and U5649 (N_5649,N_1330,N_2686);
or U5650 (N_5650,N_3834,N_3290);
or U5651 (N_5651,N_4305,N_1289);
or U5652 (N_5652,N_4776,N_716);
nor U5653 (N_5653,N_3731,N_1760);
nor U5654 (N_5654,N_2606,N_568);
nand U5655 (N_5655,N_2024,N_2583);
xor U5656 (N_5656,N_4410,N_729);
nand U5657 (N_5657,N_4765,N_2547);
and U5658 (N_5658,N_4428,N_1609);
nor U5659 (N_5659,N_1185,N_667);
nor U5660 (N_5660,N_3483,N_4605);
nand U5661 (N_5661,N_4477,N_3669);
and U5662 (N_5662,N_2764,N_3003);
nand U5663 (N_5663,N_3927,N_2644);
nand U5664 (N_5664,N_4943,N_1980);
or U5665 (N_5665,N_2510,N_3283);
nor U5666 (N_5666,N_3572,N_3510);
and U5667 (N_5667,N_4658,N_37);
nand U5668 (N_5668,N_3396,N_3341);
and U5669 (N_5669,N_4167,N_2354);
nand U5670 (N_5670,N_248,N_1281);
nor U5671 (N_5671,N_3929,N_1622);
nand U5672 (N_5672,N_1788,N_21);
and U5673 (N_5673,N_4756,N_3715);
or U5674 (N_5674,N_4568,N_1762);
and U5675 (N_5675,N_2868,N_2216);
and U5676 (N_5676,N_3228,N_2414);
nand U5677 (N_5677,N_4116,N_118);
or U5678 (N_5678,N_4393,N_2590);
nor U5679 (N_5679,N_1049,N_2272);
nor U5680 (N_5680,N_3515,N_3442);
nor U5681 (N_5681,N_3909,N_4509);
or U5682 (N_5682,N_4025,N_1732);
nand U5683 (N_5683,N_685,N_3772);
nor U5684 (N_5684,N_872,N_3512);
nand U5685 (N_5685,N_2181,N_4232);
nand U5686 (N_5686,N_2447,N_2813);
and U5687 (N_5687,N_3811,N_2768);
nand U5688 (N_5688,N_1420,N_2375);
and U5689 (N_5689,N_4616,N_1597);
nand U5690 (N_5690,N_1970,N_4642);
nor U5691 (N_5691,N_4446,N_1212);
nor U5692 (N_5692,N_2640,N_4717);
nor U5693 (N_5693,N_1218,N_3050);
nor U5694 (N_5694,N_1131,N_1209);
nor U5695 (N_5695,N_4921,N_778);
nand U5696 (N_5696,N_2592,N_3814);
and U5697 (N_5697,N_4847,N_4250);
nor U5698 (N_5698,N_949,N_4312);
nor U5699 (N_5699,N_4044,N_3607);
nor U5700 (N_5700,N_4216,N_2757);
or U5701 (N_5701,N_1426,N_231);
nor U5702 (N_5702,N_1560,N_2072);
and U5703 (N_5703,N_521,N_1227);
nor U5704 (N_5704,N_1697,N_4074);
nor U5705 (N_5705,N_1903,N_2656);
and U5706 (N_5706,N_579,N_2352);
nor U5707 (N_5707,N_732,N_1260);
nor U5708 (N_5708,N_3302,N_900);
nand U5709 (N_5709,N_743,N_4296);
nor U5710 (N_5710,N_3376,N_309);
or U5711 (N_5711,N_1180,N_4688);
and U5712 (N_5712,N_2240,N_367);
nand U5713 (N_5713,N_4339,N_2787);
nor U5714 (N_5714,N_1645,N_1679);
or U5715 (N_5715,N_2498,N_694);
or U5716 (N_5716,N_723,N_641);
nand U5717 (N_5717,N_3525,N_4125);
nor U5718 (N_5718,N_3638,N_1369);
and U5719 (N_5719,N_1270,N_2533);
nand U5720 (N_5720,N_4659,N_4557);
or U5721 (N_5721,N_4817,N_2692);
nor U5722 (N_5722,N_4396,N_501);
or U5723 (N_5723,N_3616,N_408);
or U5724 (N_5724,N_1865,N_4752);
and U5725 (N_5725,N_4897,N_3600);
or U5726 (N_5726,N_1471,N_2443);
nand U5727 (N_5727,N_1802,N_4130);
nand U5728 (N_5728,N_2182,N_1757);
nor U5729 (N_5729,N_3825,N_2634);
and U5730 (N_5730,N_1648,N_4041);
and U5731 (N_5731,N_2779,N_1965);
or U5732 (N_5732,N_1383,N_3632);
or U5733 (N_5733,N_210,N_321);
nand U5734 (N_5734,N_4645,N_2701);
or U5735 (N_5735,N_2175,N_4981);
or U5736 (N_5736,N_4668,N_225);
nor U5737 (N_5737,N_4056,N_1438);
nor U5738 (N_5738,N_2844,N_2459);
nand U5739 (N_5739,N_4078,N_3287);
nand U5740 (N_5740,N_4341,N_4114);
or U5741 (N_5741,N_3716,N_4038);
and U5742 (N_5742,N_1123,N_903);
and U5743 (N_5743,N_2031,N_2288);
or U5744 (N_5744,N_1011,N_148);
nor U5745 (N_5745,N_268,N_259);
nor U5746 (N_5746,N_3808,N_540);
and U5747 (N_5747,N_3468,N_3173);
and U5748 (N_5748,N_3130,N_1313);
and U5749 (N_5749,N_1042,N_2046);
or U5750 (N_5750,N_1308,N_3535);
nand U5751 (N_5751,N_2689,N_228);
or U5752 (N_5752,N_378,N_3001);
nand U5753 (N_5753,N_1427,N_2690);
nor U5754 (N_5754,N_3888,N_1179);
and U5755 (N_5755,N_4504,N_3157);
nor U5756 (N_5756,N_507,N_4432);
nor U5757 (N_5757,N_3737,N_3297);
or U5758 (N_5758,N_1728,N_4148);
or U5759 (N_5759,N_3145,N_792);
nand U5760 (N_5760,N_3131,N_432);
nand U5761 (N_5761,N_452,N_4374);
or U5762 (N_5762,N_1056,N_2521);
nor U5763 (N_5763,N_1365,N_418);
or U5764 (N_5764,N_4080,N_4338);
and U5765 (N_5765,N_826,N_4306);
nand U5766 (N_5766,N_971,N_508);
nor U5767 (N_5767,N_3707,N_4755);
nand U5768 (N_5768,N_2373,N_1547);
or U5769 (N_5769,N_2129,N_1673);
nand U5770 (N_5770,N_1950,N_2044);
nand U5771 (N_5771,N_2469,N_1557);
or U5772 (N_5772,N_891,N_2851);
and U5773 (N_5773,N_3273,N_3949);
and U5774 (N_5774,N_200,N_3007);
nand U5775 (N_5775,N_373,N_1996);
nor U5776 (N_5776,N_2629,N_1958);
and U5777 (N_5777,N_830,N_2431);
nand U5778 (N_5778,N_4092,N_756);
nand U5779 (N_5779,N_2277,N_2854);
nand U5780 (N_5780,N_4763,N_1414);
and U5781 (N_5781,N_3586,N_4578);
or U5782 (N_5782,N_4743,N_829);
nor U5783 (N_5783,N_874,N_3416);
or U5784 (N_5784,N_3150,N_753);
or U5785 (N_5785,N_591,N_157);
xor U5786 (N_5786,N_4839,N_2470);
nor U5787 (N_5787,N_1604,N_1895);
or U5788 (N_5788,N_4543,N_147);
or U5789 (N_5789,N_2163,N_4694);
nand U5790 (N_5790,N_3928,N_817);
or U5791 (N_5791,N_495,N_190);
and U5792 (N_5792,N_1580,N_684);
nor U5793 (N_5793,N_304,N_1302);
or U5794 (N_5794,N_4195,N_2607);
and U5795 (N_5795,N_1481,N_3603);
and U5796 (N_5796,N_3484,N_2729);
or U5797 (N_5797,N_4704,N_2898);
and U5798 (N_5798,N_362,N_4146);
nor U5799 (N_5799,N_2864,N_1431);
and U5800 (N_5800,N_4632,N_1662);
and U5801 (N_5801,N_4043,N_25);
and U5802 (N_5802,N_4483,N_2926);
and U5803 (N_5803,N_3567,N_3122);
or U5804 (N_5804,N_4796,N_192);
nor U5805 (N_5805,N_3805,N_1797);
nor U5806 (N_5806,N_4660,N_1024);
nor U5807 (N_5807,N_1661,N_1845);
and U5808 (N_5808,N_4539,N_962);
nor U5809 (N_5809,N_3218,N_1554);
nand U5810 (N_5810,N_628,N_2388);
and U5811 (N_5811,N_4360,N_740);
or U5812 (N_5812,N_543,N_1719);
nand U5813 (N_5813,N_2646,N_3239);
and U5814 (N_5814,N_1052,N_3506);
and U5815 (N_5815,N_287,N_2208);
and U5816 (N_5816,N_3978,N_1445);
and U5817 (N_5817,N_4287,N_4370);
or U5818 (N_5818,N_3612,N_3837);
nand U5819 (N_5819,N_4579,N_3910);
nor U5820 (N_5820,N_834,N_1919);
or U5821 (N_5821,N_1794,N_3895);
nand U5822 (N_5822,N_3019,N_712);
or U5823 (N_5823,N_2317,N_3870);
and U5824 (N_5824,N_1418,N_3768);
and U5825 (N_5825,N_1893,N_1367);
or U5826 (N_5826,N_997,N_3337);
or U5827 (N_5827,N_2705,N_3402);
nor U5828 (N_5828,N_2626,N_317);
nand U5829 (N_5829,N_1790,N_3878);
or U5830 (N_5830,N_2726,N_2250);
or U5831 (N_5831,N_928,N_1536);
or U5832 (N_5832,N_1680,N_3537);
and U5833 (N_5833,N_127,N_1320);
nor U5834 (N_5834,N_3698,N_3800);
and U5835 (N_5835,N_1592,N_4121);
nand U5836 (N_5836,N_2150,N_1152);
and U5837 (N_5837,N_4707,N_2806);
and U5838 (N_5838,N_4376,N_702);
and U5839 (N_5839,N_54,N_249);
and U5840 (N_5840,N_358,N_1559);
nand U5841 (N_5841,N_1029,N_2894);
and U5842 (N_5842,N_511,N_843);
and U5843 (N_5843,N_3217,N_4691);
nor U5844 (N_5844,N_536,N_1914);
or U5845 (N_5845,N_2273,N_3513);
and U5846 (N_5846,N_806,N_4277);
xor U5847 (N_5847,N_2384,N_4768);
and U5848 (N_5848,N_4110,N_662);
or U5849 (N_5849,N_4422,N_1548);
nand U5850 (N_5850,N_182,N_1441);
and U5851 (N_5851,N_2832,N_736);
xor U5852 (N_5852,N_852,N_1491);
and U5853 (N_5853,N_2391,N_4647);
nand U5854 (N_5854,N_4761,N_2477);
nor U5855 (N_5855,N_3021,N_4871);
and U5856 (N_5856,N_2386,N_3618);
nand U5857 (N_5857,N_1823,N_1157);
nor U5858 (N_5858,N_1186,N_3096);
nor U5859 (N_5859,N_3340,N_571);
or U5860 (N_5860,N_3957,N_593);
nor U5861 (N_5861,N_4525,N_3914);
or U5862 (N_5862,N_4203,N_912);
nand U5863 (N_5863,N_497,N_413);
or U5864 (N_5864,N_16,N_2203);
nand U5865 (N_5865,N_4502,N_2167);
or U5866 (N_5866,N_4654,N_97);
and U5867 (N_5867,N_2842,N_2490);
nor U5868 (N_5868,N_3667,N_4363);
nand U5869 (N_5869,N_537,N_1612);
nand U5870 (N_5870,N_130,N_425);
nor U5871 (N_5871,N_1116,N_2400);
and U5872 (N_5872,N_1,N_2960);
nor U5873 (N_5873,N_2192,N_3861);
nand U5874 (N_5874,N_2229,N_1499);
nand U5875 (N_5875,N_3388,N_728);
nand U5876 (N_5876,N_2310,N_2291);
nand U5877 (N_5877,N_116,N_859);
nor U5878 (N_5878,N_2243,N_4050);
and U5879 (N_5879,N_2542,N_2293);
or U5880 (N_5880,N_1231,N_2006);
and U5881 (N_5881,N_1717,N_3177);
nand U5882 (N_5882,N_1267,N_3455);
nor U5883 (N_5883,N_3129,N_1217);
nor U5884 (N_5884,N_4429,N_2318);
and U5885 (N_5885,N_1073,N_2331);
nor U5886 (N_5886,N_1981,N_1148);
nand U5887 (N_5887,N_19,N_4294);
nand U5888 (N_5888,N_2753,N_4923);
and U5889 (N_5889,N_2828,N_2179);
or U5890 (N_5890,N_2071,N_1005);
or U5891 (N_5891,N_125,N_4913);
nor U5892 (N_5892,N_2628,N_4493);
and U5893 (N_5893,N_940,N_3590);
and U5894 (N_5894,N_1269,N_1133);
or U5895 (N_5895,N_3696,N_1301);
and U5896 (N_5896,N_3675,N_2435);
or U5897 (N_5897,N_4586,N_320);
or U5898 (N_5898,N_3872,N_278);
nand U5899 (N_5899,N_2995,N_898);
and U5900 (N_5900,N_4786,N_3585);
or U5901 (N_5901,N_345,N_2063);
nand U5902 (N_5902,N_3857,N_256);
and U5903 (N_5903,N_3326,N_3972);
or U5904 (N_5904,N_4988,N_3793);
nor U5905 (N_5905,N_3796,N_1558);
nor U5906 (N_5906,N_4760,N_624);
nand U5907 (N_5907,N_4301,N_4626);
nand U5908 (N_5908,N_3417,N_1248);
and U5909 (N_5909,N_3529,N_2499);
and U5910 (N_5910,N_4359,N_3320);
nor U5911 (N_5911,N_2991,N_1473);
nor U5912 (N_5912,N_2976,N_1729);
nand U5913 (N_5913,N_763,N_3478);
and U5914 (N_5914,N_4362,N_538);
nor U5915 (N_5915,N_2458,N_3361);
or U5916 (N_5916,N_4903,N_1957);
or U5917 (N_5917,N_953,N_1809);
or U5918 (N_5918,N_1949,N_2967);
and U5919 (N_5919,N_2763,N_993);
and U5920 (N_5920,N_4329,N_2316);
nor U5921 (N_5921,N_818,N_1755);
nand U5922 (N_5922,N_2497,N_3816);
or U5923 (N_5923,N_1746,N_3333);
nor U5924 (N_5924,N_1607,N_1053);
nand U5925 (N_5925,N_4917,N_2548);
nor U5926 (N_5926,N_3325,N_260);
or U5927 (N_5927,N_162,N_4856);
or U5928 (N_5928,N_3229,N_1238);
and U5929 (N_5929,N_884,N_1774);
or U5930 (N_5930,N_3245,N_3789);
and U5931 (N_5931,N_1967,N_2681);
nand U5932 (N_5932,N_2233,N_4156);
nand U5933 (N_5933,N_250,N_4371);
and U5934 (N_5934,N_1857,N_1229);
nand U5935 (N_5935,N_44,N_4878);
nand U5936 (N_5936,N_4325,N_3463);
or U5937 (N_5937,N_2103,N_3041);
nor U5938 (N_5938,N_4138,N_1759);
nor U5939 (N_5939,N_4993,N_4202);
and U5940 (N_5940,N_3125,N_3596);
nand U5941 (N_5941,N_3231,N_4064);
nor U5942 (N_5942,N_1081,N_3706);
and U5943 (N_5943,N_1168,N_2598);
nor U5944 (N_5944,N_2475,N_4932);
or U5945 (N_5945,N_1295,N_916);
nand U5946 (N_5946,N_4547,N_968);
and U5947 (N_5947,N_4580,N_3597);
nor U5948 (N_5948,N_2267,N_3718);
nand U5949 (N_5949,N_994,N_640);
and U5950 (N_5950,N_582,N_3081);
and U5951 (N_5951,N_1726,N_3335);
and U5952 (N_5952,N_3649,N_2662);
and U5953 (N_5953,N_2800,N_4612);
nand U5954 (N_5954,N_2552,N_2428);
nor U5955 (N_5955,N_4275,N_1393);
and U5956 (N_5956,N_2100,N_244);
and U5957 (N_5957,N_4829,N_717);
nor U5958 (N_5958,N_265,N_3343);
or U5959 (N_5959,N_4180,N_4747);
and U5960 (N_5960,N_2043,N_2116);
or U5961 (N_5961,N_703,N_4908);
nand U5962 (N_5962,N_4479,N_2471);
or U5963 (N_5963,N_2440,N_4002);
and U5964 (N_5964,N_3458,N_70);
and U5965 (N_5965,N_136,N_252);
nand U5966 (N_5966,N_4741,N_651);
nor U5967 (N_5967,N_2460,N_3029);
nand U5968 (N_5968,N_3293,N_2187);
nand U5969 (N_5969,N_386,N_4461);
or U5970 (N_5970,N_3726,N_2483);
or U5971 (N_5971,N_1055,N_4692);
nand U5972 (N_5972,N_2749,N_2605);
nor U5973 (N_5973,N_2507,N_4310);
or U5974 (N_5974,N_692,N_3973);
nor U5975 (N_5975,N_2945,N_4900);
or U5976 (N_5976,N_2614,N_169);
and U5977 (N_5977,N_4259,N_4672);
or U5978 (N_5978,N_3398,N_370);
nor U5979 (N_5979,N_2172,N_1503);
or U5980 (N_5980,N_1136,N_2429);
nand U5981 (N_5981,N_2170,N_2132);
or U5982 (N_5982,N_1688,N_1660);
and U5983 (N_5983,N_4083,N_2559);
xor U5984 (N_5984,N_1068,N_4976);
nor U5985 (N_5985,N_799,N_948);
or U5986 (N_5986,N_1066,N_1060);
or U5987 (N_5987,N_3411,N_4367);
nand U5988 (N_5988,N_3990,N_3319);
or U5989 (N_5989,N_3541,N_8);
and U5990 (N_5990,N_1830,N_2213);
or U5991 (N_5991,N_2657,N_1638);
and U5992 (N_5992,N_3781,N_745);
or U5993 (N_5993,N_531,N_2422);
or U5994 (N_5994,N_35,N_1812);
or U5995 (N_5995,N_2580,N_4545);
and U5996 (N_5996,N_3368,N_4350);
nand U5997 (N_5997,N_3933,N_2370);
nor U5998 (N_5998,N_3085,N_4584);
and U5999 (N_5999,N_1019,N_4901);
nand U6000 (N_6000,N_4676,N_1576);
or U6001 (N_6001,N_3580,N_3299);
nand U6002 (N_6002,N_2653,N_1512);
and U6003 (N_6003,N_4087,N_2683);
or U6004 (N_6004,N_2093,N_242);
or U6005 (N_6005,N_613,N_2884);
xor U6006 (N_6006,N_3317,N_1337);
and U6007 (N_6007,N_3986,N_1488);
and U6008 (N_6008,N_2158,N_1868);
and U6009 (N_6009,N_4405,N_541);
nor U6010 (N_6010,N_869,N_522);
and U6011 (N_6011,N_4035,N_1210);
xnor U6012 (N_6012,N_4303,N_1827);
nor U6013 (N_6013,N_3899,N_1861);
nand U6014 (N_6014,N_2159,N_4534);
nor U6015 (N_6015,N_2199,N_1244);
nand U6016 (N_6016,N_80,N_2804);
and U6017 (N_6017,N_1743,N_2625);
or U6018 (N_6018,N_238,N_4384);
and U6019 (N_6019,N_4314,N_3384);
and U6020 (N_6020,N_109,N_1026);
nor U6021 (N_6021,N_2735,N_2722);
and U6022 (N_6022,N_1415,N_2557);
or U6023 (N_6023,N_1631,N_4728);
or U6024 (N_6024,N_1700,N_2643);
and U6025 (N_6025,N_3437,N_2148);
and U6026 (N_6026,N_1883,N_1819);
nand U6027 (N_6027,N_3233,N_2137);
or U6028 (N_6028,N_1310,N_2781);
or U6029 (N_6029,N_2922,N_2914);
nor U6030 (N_6030,N_1703,N_747);
or U6031 (N_6031,N_272,N_4815);
nand U6032 (N_6032,N_3998,N_2835);
or U6033 (N_6033,N_423,N_3105);
nor U6034 (N_6034,N_4537,N_3762);
and U6035 (N_6035,N_2304,N_3729);
and U6036 (N_6036,N_450,N_815);
or U6037 (N_6037,N_3214,N_2421);
or U6038 (N_6038,N_2715,N_4818);
and U6039 (N_6039,N_3166,N_89);
nand U6040 (N_6040,N_635,N_398);
or U6041 (N_6041,N_4982,N_1341);
nand U6042 (N_6042,N_707,N_3594);
or U6043 (N_6043,N_2994,N_3253);
and U6044 (N_6044,N_4153,N_3485);
and U6045 (N_6045,N_1047,N_3244);
and U6046 (N_6046,N_1402,N_1467);
or U6047 (N_6047,N_4448,N_1400);
or U6048 (N_6048,N_2123,N_709);
and U6049 (N_6049,N_3025,N_4424);
and U6050 (N_6050,N_1921,N_4139);
or U6051 (N_6051,N_1814,N_1111);
and U6052 (N_6052,N_2042,N_2966);
nor U6053 (N_6053,N_2420,N_2908);
nand U6054 (N_6054,N_2918,N_2270);
or U6055 (N_6055,N_42,N_3868);
and U6056 (N_6056,N_1984,N_3433);
nor U6057 (N_6057,N_2184,N_833);
and U6058 (N_6058,N_4588,N_3810);
or U6059 (N_6059,N_2183,N_2696);
or U6060 (N_6060,N_3508,N_3946);
and U6061 (N_6061,N_3598,N_2913);
and U6062 (N_6062,N_3602,N_4754);
nor U6063 (N_6063,N_94,N_977);
and U6064 (N_6064,N_3256,N_3923);
and U6065 (N_6065,N_3873,N_2338);
nand U6066 (N_6066,N_3056,N_3111);
nor U6067 (N_6067,N_1093,N_3170);
nand U6068 (N_6068,N_2988,N_2088);
nor U6069 (N_6069,N_3415,N_518);
nor U6070 (N_6070,N_1633,N_4187);
and U6071 (N_6071,N_4862,N_391);
and U6072 (N_6072,N_2013,N_2204);
and U6073 (N_6073,N_4358,N_1702);
or U6074 (N_6074,N_1754,N_1875);
nor U6075 (N_6075,N_4521,N_1041);
nor U6076 (N_6076,N_3200,N_3547);
nor U6077 (N_6077,N_3011,N_1220);
and U6078 (N_6078,N_2014,N_2661);
nor U6079 (N_6079,N_4066,N_3579);
nor U6080 (N_6080,N_1768,N_814);
nand U6081 (N_6081,N_2801,N_2952);
or U6082 (N_6082,N_3272,N_4103);
nor U6083 (N_6083,N_960,N_3959);
and U6084 (N_6084,N_766,N_439);
nand U6085 (N_6085,N_1911,N_3370);
nand U6086 (N_6086,N_240,N_2099);
xor U6087 (N_6087,N_3237,N_1678);
nor U6088 (N_6088,N_1711,N_3171);
xor U6089 (N_6089,N_311,N_2858);
nand U6090 (N_6090,N_4419,N_1880);
nand U6091 (N_6091,N_1147,N_1562);
or U6092 (N_6092,N_4894,N_2795);
and U6093 (N_6093,N_3645,N_2324);
or U6094 (N_6094,N_550,N_2055);
nor U6095 (N_6095,N_2695,N_4106);
or U6096 (N_6096,N_3198,N_4774);
nand U6097 (N_6097,N_2398,N_4051);
or U6098 (N_6098,N_3044,N_1259);
nand U6099 (N_6099,N_3792,N_681);
and U6100 (N_6100,N_159,N_4382);
or U6101 (N_6101,N_4495,N_2326);
and U6102 (N_6102,N_631,N_560);
nand U6103 (N_6103,N_4001,N_1765);
and U6104 (N_6104,N_2214,N_816);
nand U6105 (N_6105,N_2287,N_929);
and U6106 (N_6106,N_4663,N_455);
or U6107 (N_6107,N_1654,N_3430);
nand U6108 (N_6108,N_4319,N_2322);
nand U6109 (N_6109,N_3629,N_463);
nor U6110 (N_6110,N_331,N_1643);
nand U6111 (N_6111,N_1826,N_2944);
nand U6112 (N_6112,N_2450,N_2185);
and U6113 (N_6113,N_3574,N_2932);
and U6114 (N_6114,N_4208,N_1388);
nand U6115 (N_6115,N_1256,N_1072);
and U6116 (N_6116,N_2694,N_3065);
nand U6117 (N_6117,N_2073,N_4629);
nand U6118 (N_6118,N_4031,N_1621);
and U6119 (N_6119,N_3062,N_4698);
and U6120 (N_6120,N_1258,N_2102);
nand U6121 (N_6121,N_3087,N_1346);
or U6122 (N_6122,N_2961,N_1057);
nand U6123 (N_6123,N_3334,N_4961);
and U6124 (N_6124,N_3942,N_4898);
or U6125 (N_6125,N_1197,N_1146);
nand U6126 (N_6126,N_4183,N_4618);
nor U6127 (N_6127,N_4005,N_3881);
nor U6128 (N_6128,N_4284,N_4129);
nor U6129 (N_6129,N_4398,N_65);
or U6130 (N_6130,N_2486,N_3386);
nand U6131 (N_6131,N_512,N_4010);
nor U6132 (N_6132,N_2284,N_435);
nand U6133 (N_6133,N_3160,N_1773);
nor U6134 (N_6134,N_870,N_879);
and U6135 (N_6135,N_1193,N_825);
or U6136 (N_6136,N_2594,N_2335);
and U6137 (N_6137,N_4944,N_2989);
nor U6138 (N_6138,N_2415,N_4172);
nor U6139 (N_6139,N_4104,N_1482);
and U6140 (N_6140,N_1064,N_1644);
nor U6141 (N_6141,N_4119,N_3725);
and U6142 (N_6142,N_2972,N_944);
and U6143 (N_6143,N_1939,N_2652);
or U6144 (N_6144,N_4689,N_4368);
and U6145 (N_6145,N_1553,N_786);
or U6146 (N_6146,N_1046,N_4437);
or U6147 (N_6147,N_4455,N_773);
and U6148 (N_6148,N_1923,N_3394);
and U6149 (N_6149,N_4159,N_4149);
nor U6150 (N_6150,N_2249,N_782);
or U6151 (N_6151,N_1145,N_2807);
and U6152 (N_6152,N_2783,N_3159);
or U6153 (N_6153,N_3045,N_1545);
and U6154 (N_6154,N_1462,N_376);
nand U6155 (N_6155,N_4910,N_669);
nand U6156 (N_6156,N_2860,N_1478);
xor U6157 (N_6157,N_341,N_4863);
nor U6158 (N_6158,N_1389,N_291);
and U6159 (N_6159,N_3771,N_3952);
and U6160 (N_6160,N_544,N_2970);
or U6161 (N_6161,N_3199,N_4241);
or U6162 (N_6162,N_1314,N_3958);
nor U6163 (N_6163,N_4194,N_2850);
or U6164 (N_6164,N_3538,N_1171);
and U6165 (N_6165,N_3148,N_2274);
or U6166 (N_6166,N_4527,N_1102);
nand U6167 (N_6167,N_3817,N_1447);
nor U6168 (N_6168,N_394,N_3995);
and U6169 (N_6169,N_3673,N_4684);
and U6170 (N_6170,N_3900,N_1685);
and U6171 (N_6171,N_1245,N_693);
or U6172 (N_6172,N_3844,N_4690);
or U6173 (N_6173,N_523,N_123);
nand U6174 (N_6174,N_1841,N_4677);
nor U6175 (N_6175,N_2441,N_3977);
nor U6176 (N_6176,N_1202,N_936);
and U6177 (N_6177,N_4794,N_1464);
and U6178 (N_6178,N_2366,N_516);
nand U6179 (N_6179,N_3185,N_4998);
and U6180 (N_6180,N_730,N_262);
nand U6181 (N_6181,N_2755,N_1395);
nand U6182 (N_6182,N_2406,N_3938);
nand U6183 (N_6183,N_1079,N_3504);
and U6184 (N_6184,N_731,N_3786);
or U6185 (N_6185,N_4846,N_4942);
and U6186 (N_6186,N_475,N_4700);
or U6187 (N_6187,N_2802,N_1963);
and U6188 (N_6188,N_4930,N_4089);
nor U6189 (N_6189,N_513,N_2209);
and U6190 (N_6190,N_2572,N_416);
and U6191 (N_6191,N_802,N_1932);
and U6192 (N_6192,N_783,N_2959);
and U6193 (N_6193,N_4166,N_4458);
nor U6194 (N_6194,N_4657,N_4452);
and U6195 (N_6195,N_3004,N_3449);
nand U6196 (N_6196,N_243,N_1692);
and U6197 (N_6197,N_4280,N_1432);
nor U6198 (N_6198,N_4844,N_4600);
and U6199 (N_6199,N_1292,N_1234);
nor U6200 (N_6200,N_2950,N_4683);
nor U6201 (N_6201,N_2927,N_3551);
nand U6202 (N_6202,N_315,N_762);
nor U6203 (N_6203,N_2825,N_4506);
nand U6204 (N_6204,N_2402,N_1362);
nand U6205 (N_6205,N_1878,N_1641);
and U6206 (N_6206,N_1670,N_995);
and U6207 (N_6207,N_3292,N_643);
xnor U6208 (N_6208,N_3849,N_1034);
and U6209 (N_6209,N_4257,N_2067);
or U6210 (N_6210,N_725,N_2817);
nand U6211 (N_6211,N_1501,N_1831);
or U6212 (N_6212,N_4751,N_0);
and U6213 (N_6213,N_1530,N_3651);
xor U6214 (N_6214,N_2035,N_172);
nor U6215 (N_6215,N_4715,N_4798);
or U6216 (N_6216,N_3822,N_1002);
or U6217 (N_6217,N_3755,N_1531);
and U6218 (N_6218,N_1959,N_66);
and U6219 (N_6219,N_3730,N_4449);
nor U6220 (N_6220,N_1184,N_2977);
nand U6221 (N_6221,N_1527,N_4945);
nor U6222 (N_6222,N_3740,N_2228);
nor U6223 (N_6223,N_4248,N_983);
and U6224 (N_6224,N_1579,N_2104);
nor U6225 (N_6225,N_2196,N_461);
and U6226 (N_6226,N_1084,N_120);
nor U6227 (N_6227,N_4940,N_4373);
or U6228 (N_6228,N_3015,N_1239);
nand U6229 (N_6229,N_1465,N_585);
or U6230 (N_6230,N_4188,N_3042);
xnor U6231 (N_6231,N_221,N_4150);
and U6232 (N_6232,N_4196,N_1401);
nand U6233 (N_6233,N_4749,N_1206);
nand U6234 (N_6234,N_168,N_27);
or U6235 (N_6235,N_832,N_53);
nor U6236 (N_6236,N_2463,N_672);
nand U6237 (N_6237,N_1357,N_1128);
or U6238 (N_6238,N_3503,N_739);
or U6239 (N_6239,N_1198,N_2886);
or U6240 (N_6240,N_708,N_1119);
nor U6241 (N_6241,N_2345,N_4175);
nor U6242 (N_6242,N_3249,N_4807);
and U6243 (N_6243,N_947,N_2826);
nor U6244 (N_6244,N_3094,N_4631);
nor U6245 (N_6245,N_4523,N_2083);
nor U6246 (N_6246,N_2808,N_2294);
and U6247 (N_6247,N_2461,N_4710);
nor U6248 (N_6248,N_1742,N_4236);
nor U6249 (N_6249,N_332,N_3262);
nor U6250 (N_6250,N_2278,N_3752);
or U6251 (N_6251,N_1106,N_24);
nand U6252 (N_6252,N_3338,N_3943);
nor U6253 (N_6253,N_2193,N_3473);
nor U6254 (N_6254,N_4840,N_923);
nand U6255 (N_6255,N_2746,N_3347);
and U6256 (N_6256,N_3061,N_1777);
nor U6257 (N_6257,N_4615,N_2876);
nor U6258 (N_6258,N_876,N_410);
or U6259 (N_6259,N_2756,N_3037);
or U6260 (N_6260,N_1505,N_4059);
nand U6261 (N_6261,N_3271,N_4895);
and U6262 (N_6262,N_4096,N_4769);
or U6263 (N_6263,N_798,N_1181);
nor U6264 (N_6264,N_211,N_4200);
and U6265 (N_6265,N_3757,N_216);
or U6266 (N_6266,N_2543,N_282);
nor U6267 (N_6267,N_4263,N_2725);
or U6268 (N_6268,N_2142,N_2360);
and U6269 (N_6269,N_4979,N_2139);
and U6270 (N_6270,N_3362,N_1230);
nand U6271 (N_6271,N_4162,N_4619);
nor U6272 (N_6272,N_680,N_3767);
or U6273 (N_6273,N_1509,N_1614);
or U6274 (N_6274,N_4957,N_670);
nor U6275 (N_6275,N_3379,N_4737);
nor U6276 (N_6276,N_4681,N_781);
nand U6277 (N_6277,N_4983,N_2911);
nor U6278 (N_6278,N_4697,N_2553);
and U6279 (N_6279,N_3397,N_2417);
and U6280 (N_6280,N_1985,N_4964);
and U6281 (N_6281,N_3296,N_1635);
and U6282 (N_6282,N_2247,N_4995);
nor U6283 (N_6283,N_4498,N_1158);
and U6284 (N_6284,N_1853,N_4806);
nand U6285 (N_6285,N_1837,N_301);
or U6286 (N_6286,N_3864,N_1636);
xor U6287 (N_6287,N_4939,N_4952);
and U6288 (N_6288,N_3010,N_2307);
nor U6289 (N_6289,N_3135,N_3842);
nor U6290 (N_6290,N_2732,N_2392);
nor U6291 (N_6291,N_1497,N_850);
or U6292 (N_6292,N_1867,N_2675);
and U6293 (N_6293,N_4264,N_4381);
and U6294 (N_6294,N_3891,N_4418);
nor U6295 (N_6295,N_1390,N_3311);
and U6296 (N_6296,N_1338,N_1546);
nor U6297 (N_6297,N_4409,N_3414);
nand U6298 (N_6298,N_1990,N_4656);
nand U6299 (N_6299,N_4978,N_3963);
and U6300 (N_6300,N_2082,N_2115);
and U6301 (N_6301,N_2068,N_3671);
nand U6302 (N_6302,N_570,N_4433);
and U6303 (N_6303,N_3298,N_4799);
nand U6304 (N_6304,N_2091,N_3133);
nand U6305 (N_6305,N_2201,N_3070);
or U6306 (N_6306,N_1627,N_4364);
nor U6307 (N_6307,N_4186,N_2882);
nand U6308 (N_6308,N_808,N_2716);
or U6309 (N_6309,N_4721,N_3806);
nor U6310 (N_6310,N_4191,N_115);
nor U6311 (N_6311,N_3382,N_4789);
or U6312 (N_6312,N_865,N_2872);
nand U6313 (N_6313,N_4750,N_4379);
nand U6314 (N_6314,N_1477,N_368);
or U6315 (N_6315,N_4609,N_2999);
or U6316 (N_6316,N_3104,N_4201);
nand U6317 (N_6317,N_2535,N_4994);
or U6318 (N_6318,N_1606,N_2219);
or U6319 (N_6319,N_955,N_2979);
and U6320 (N_6320,N_4503,N_178);
xor U6321 (N_6321,N_56,N_401);
nand U6322 (N_6322,N_4052,N_1208);
or U6323 (N_6323,N_4311,N_658);
nor U6324 (N_6324,N_2265,N_2516);
nand U6325 (N_6325,N_4018,N_2112);
and U6326 (N_6326,N_3703,N_1602);
nand U6327 (N_6327,N_4178,N_478);
nor U6328 (N_6328,N_780,N_3523);
nand U6329 (N_6329,N_1863,N_4075);
and U6330 (N_6330,N_3097,N_3695);
nand U6331 (N_6331,N_82,N_4260);
and U6332 (N_6332,N_254,N_2276);
nand U6333 (N_6333,N_338,N_4544);
nand U6334 (N_6334,N_4434,N_1568);
and U6335 (N_6335,N_1822,N_2611);
or U6336 (N_6336,N_2651,N_2596);
or U6337 (N_6337,N_303,N_856);
nor U6338 (N_6338,N_4225,N_759);
or U6339 (N_6339,N_4966,N_1525);
nor U6340 (N_6340,N_494,N_4169);
and U6341 (N_6341,N_4300,N_565);
nand U6342 (N_6342,N_2282,N_2733);
nand U6343 (N_6343,N_2775,N_2438);
or U6344 (N_6344,N_1262,N_3717);
and U6345 (N_6345,N_163,N_3948);
and U6346 (N_6346,N_1796,N_68);
nand U6347 (N_6347,N_4899,N_2867);
or U6348 (N_6348,N_312,N_1469);
nand U6349 (N_6349,N_3683,N_1716);
or U6350 (N_6350,N_3866,N_504);
and U6351 (N_6351,N_592,N_2412);
nor U6352 (N_6352,N_2793,N_420);
nor U6353 (N_6353,N_3277,N_4335);
nor U6354 (N_6354,N_1847,N_197);
nor U6355 (N_6355,N_4643,N_1889);
nand U6356 (N_6356,N_3434,N_1782);
nor U6357 (N_6357,N_3530,N_4746);
nor U6358 (N_6358,N_3749,N_1675);
and U6359 (N_6359,N_273,N_2309);
nand U6360 (N_6360,N_4764,N_4077);
or U6361 (N_6361,N_213,N_2144);
or U6362 (N_6362,N_3263,N_3100);
nor U6363 (N_6363,N_2040,N_2336);
or U6364 (N_6364,N_4680,N_4569);
and U6365 (N_6365,N_1485,N_721);
nor U6366 (N_6366,N_2141,N_4984);
or U6367 (N_6367,N_3113,N_2600);
and U6368 (N_6368,N_572,N_3518);
and U6369 (N_6369,N_627,N_2546);
or U6370 (N_6370,N_805,N_187);
or U6371 (N_6371,N_3846,N_4997);
nor U6372 (N_6372,N_4467,N_3059);
or U6373 (N_6373,N_4193,N_4549);
or U6374 (N_6374,N_1196,N_774);
nand U6375 (N_6375,N_878,N_3828);
and U6376 (N_6376,N_4791,N_1650);
nor U6377 (N_6377,N_1312,N_2709);
or U6378 (N_6378,N_4974,N_587);
nor U6379 (N_6379,N_3654,N_4601);
or U6380 (N_6380,N_4941,N_4404);
nand U6381 (N_6381,N_1815,N_402);
nand U6382 (N_6382,N_2878,N_668);
or U6383 (N_6383,N_2077,N_4777);
nor U6384 (N_6384,N_3066,N_1724);
nor U6385 (N_6385,N_1813,N_1411);
nor U6386 (N_6386,N_989,N_3438);
nand U6387 (N_6387,N_3046,N_3693);
or U6388 (N_6388,N_4430,N_4833);
or U6389 (N_6389,N_1689,N_2076);
nand U6390 (N_6390,N_4969,N_4450);
nor U6391 (N_6391,N_1307,N_4058);
nor U6392 (N_6392,N_895,N_2514);
or U6393 (N_6393,N_548,N_2579);
or U6394 (N_6394,N_1975,N_355);
or U6395 (N_6395,N_4703,N_3489);
or U6396 (N_6396,N_3621,N_2);
nand U6397 (N_6397,N_224,N_1710);
and U6398 (N_6398,N_2118,N_2532);
or U6399 (N_6399,N_3474,N_3967);
nor U6400 (N_6400,N_4877,N_559);
and U6401 (N_6401,N_3144,N_4141);
nand U6402 (N_6402,N_3216,N_2677);
nor U6403 (N_6403,N_2487,N_4808);
and U6404 (N_6404,N_603,N_1183);
and U6405 (N_6405,N_1997,N_1860);
or U6406 (N_6406,N_1647,N_3521);
and U6407 (N_6407,N_4996,N_1236);
and U6408 (N_6408,N_887,N_1187);
or U6409 (N_6409,N_3869,N_1514);
nand U6410 (N_6410,N_1446,N_4753);
nor U6411 (N_6411,N_742,N_3705);
or U6412 (N_6412,N_1634,N_218);
or U6413 (N_6413,N_1961,N_3920);
nor U6414 (N_6414,N_2111,N_4855);
or U6415 (N_6415,N_3172,N_3454);
or U6416 (N_6416,N_2264,N_4511);
and U6417 (N_6417,N_1901,N_2880);
and U6418 (N_6418,N_4365,N_2963);
or U6419 (N_6419,N_3728,N_4008);
nand U6420 (N_6420,N_2405,N_4249);
xor U6421 (N_6421,N_2206,N_1493);
nand U6422 (N_6422,N_2750,N_3175);
and U6423 (N_6423,N_1101,N_598);
or U6424 (N_6424,N_1734,N_1322);
or U6425 (N_6425,N_897,N_3554);
or U6426 (N_6426,N_659,N_4473);
nor U6427 (N_6427,N_586,N_1324);
nor U6428 (N_6428,N_399,N_3392);
nor U6429 (N_6429,N_313,N_4413);
and U6430 (N_6430,N_4011,N_1333);
or U6431 (N_6431,N_2838,N_1048);
nand U6432 (N_6432,N_863,N_3365);
nor U6433 (N_6433,N_1327,N_3264);
nand U6434 (N_6434,N_4219,N_426);
or U6435 (N_6435,N_4135,N_2074);
and U6436 (N_6436,N_959,N_4454);
nand U6437 (N_6437,N_3353,N_2098);
or U6438 (N_6438,N_2303,N_1974);
nand U6439 (N_6439,N_2837,N_1141);
or U6440 (N_6440,N_98,N_3374);
or U6441 (N_6441,N_2342,N_2962);
and U6442 (N_6442,N_453,N_3371);
nor U6443 (N_6443,N_784,N_3327);
nand U6444 (N_6444,N_3565,N_2389);
nor U6445 (N_6445,N_1656,N_2571);
and U6446 (N_6446,N_1178,N_1772);
nand U6447 (N_6447,N_3647,N_4124);
nand U6448 (N_6448,N_5,N_330);
and U6449 (N_6449,N_1377,N_583);
and U6450 (N_6450,N_4625,N_3913);
nor U6451 (N_6451,N_2125,N_3152);
or U6452 (N_6452,N_653,N_4610);
nand U6453 (N_6453,N_1366,N_3270);
or U6454 (N_6454,N_1810,N_1044);
or U6455 (N_6455,N_2337,N_99);
or U6456 (N_6456,N_215,N_3267);
and U6457 (N_6457,N_1532,N_2563);
nand U6458 (N_6458,N_3108,N_2949);
or U6459 (N_6459,N_2975,N_827);
xnor U6460 (N_6460,N_281,N_3584);
nand U6461 (N_6461,N_836,N_3031);
and U6462 (N_6462,N_4781,N_4792);
and U6463 (N_6463,N_143,N_196);
nand U6464 (N_6464,N_359,N_2289);
and U6465 (N_6465,N_2387,N_3610);
nand U6466 (N_6466,N_3500,N_837);
and U6467 (N_6467,N_1872,N_3569);
or U6468 (N_6468,N_388,N_3344);
or U6469 (N_6469,N_3146,N_380);
nor U6470 (N_6470,N_4572,N_403);
and U6471 (N_6471,N_2641,N_1169);
nor U6472 (N_6472,N_466,N_2748);
nor U6473 (N_6473,N_4261,N_942);
nand U6474 (N_6474,N_3196,N_1871);
nand U6475 (N_6475,N_2121,N_3000);
nand U6476 (N_6476,N_3678,N_964);
or U6477 (N_6477,N_1374,N_117);
nor U6478 (N_6478,N_533,N_1348);
and U6479 (N_6479,N_3142,N_2904);
and U6480 (N_6480,N_1882,N_3783);
nand U6481 (N_6481,N_3637,N_4288);
and U6482 (N_6482,N_3622,N_3633);
nand U6483 (N_6483,N_2482,N_3836);
nor U6484 (N_6484,N_2292,N_1107);
or U6485 (N_6485,N_3912,N_2631);
and U6486 (N_6486,N_4904,N_393);
nor U6487 (N_6487,N_4552,N_348);
xor U6488 (N_6488,N_3127,N_532);
and U6489 (N_6489,N_2554,N_325);
nor U6490 (N_6490,N_4488,N_1424);
and U6491 (N_6491,N_106,N_1027);
or U6492 (N_6492,N_1235,N_3441);
nand U6493 (N_6493,N_4268,N_4174);
nor U6494 (N_6494,N_3745,N_3791);
nor U6495 (N_6495,N_2197,N_1832);
and U6496 (N_6496,N_1955,N_4117);
nor U6497 (N_6497,N_326,N_3655);
nand U6498 (N_6498,N_2248,N_3735);
or U6499 (N_6499,N_4102,N_4667);
or U6500 (N_6500,N_1862,N_174);
nand U6501 (N_6501,N_3378,N_4326);
and U6502 (N_6502,N_2968,N_4285);
and U6503 (N_6503,N_1284,N_2544);
nand U6504 (N_6504,N_3403,N_3440);
nand U6505 (N_6505,N_4016,N_2311);
and U6506 (N_6506,N_683,N_1539);
and U6507 (N_6507,N_1751,N_1640);
nor U6508 (N_6508,N_3785,N_2815);
nor U6509 (N_6509,N_4255,N_4086);
nor U6510 (N_6510,N_3187,N_3953);
or U6511 (N_6511,N_2762,N_1451);
and U6512 (N_6512,N_1349,N_2401);
nor U6513 (N_6513,N_3936,N_1358);
nand U6514 (N_6514,N_183,N_464);
nor U6515 (N_6515,N_3049,N_546);
nor U6516 (N_6516,N_3321,N_3400);
or U6517 (N_6517,N_855,N_2026);
nor U6518 (N_6518,N_2242,N_295);
nor U6519 (N_6519,N_4063,N_607);
nor U6520 (N_6520,N_2426,N_3226);
and U6521 (N_6521,N_3301,N_2080);
nand U6522 (N_6522,N_4047,N_4421);
nand U6523 (N_6523,N_1803,N_1666);
and U6524 (N_6524,N_3324,N_882);
nand U6525 (N_6525,N_1115,N_1360);
nor U6526 (N_6526,N_4883,N_3456);
or U6527 (N_6527,N_2946,N_3876);
and U6528 (N_6528,N_1913,N_2410);
nor U6529 (N_6529,N_2719,N_4151);
nand U6530 (N_6530,N_3316,N_1720);
nor U6531 (N_6531,N_4675,N_2863);
nand U6532 (N_6532,N_3754,N_789);
nand U6533 (N_6533,N_4331,N_1535);
and U6534 (N_6534,N_1250,N_677);
or U6535 (N_6535,N_4686,N_2106);
and U6536 (N_6536,N_2742,N_1594);
nand U6537 (N_6537,N_1686,N_2721);
nand U6538 (N_6538,N_4478,N_3459);
nand U6539 (N_6539,N_438,N_1182);
or U6540 (N_6540,N_3561,N_3674);
and U6541 (N_6541,N_749,N_4788);
or U6542 (N_6542,N_2070,N_2582);
nor U6543 (N_6543,N_3812,N_4245);
and U6544 (N_6544,N_2765,N_1059);
nand U6545 (N_6545,N_3348,N_3901);
and U6546 (N_6546,N_4824,N_1215);
nor U6547 (N_6547,N_4936,N_2874);
nand U6548 (N_6548,N_2556,N_161);
or U6549 (N_6549,N_4337,N_3918);
and U6550 (N_6550,N_1453,N_1551);
and U6551 (N_6551,N_3619,N_2162);
nor U6552 (N_6552,N_3071,N_3930);
and U6553 (N_6553,N_2668,N_2424);
and U6554 (N_6554,N_279,N_2161);
or U6555 (N_6555,N_26,N_3209);
nor U6556 (N_6556,N_3095,N_3879);
nor U6557 (N_6557,N_1458,N_4496);
or U6558 (N_6558,N_2339,N_2385);
nand U6559 (N_6559,N_1082,N_2846);
or U6560 (N_6560,N_4251,N_620);
and U6561 (N_6561,N_476,N_1363);
or U6562 (N_6562,N_3795,N_4739);
or U6563 (N_6563,N_1897,N_502);
and U6564 (N_6564,N_1684,N_2738);
nand U6565 (N_6565,N_4021,N_758);
or U6566 (N_6566,N_93,N_104);
nor U6567 (N_6567,N_1529,N_3221);
or U6568 (N_6568,N_3576,N_3775);
xnor U6569 (N_6569,N_2409,N_1962);
and U6570 (N_6570,N_1655,N_848);
or U6571 (N_6571,N_227,N_3498);
and U6572 (N_6572,N_4348,N_644);
or U6573 (N_6573,N_1603,N_2089);
nor U6574 (N_6574,N_700,N_2812);
or U6575 (N_6575,N_886,N_801);
or U6576 (N_6576,N_3636,N_3802);
xor U6577 (N_6577,N_1510,N_922);
nand U6578 (N_6578,N_229,N_1408);
or U6579 (N_6579,N_3961,N_820);
and U6580 (N_6580,N_165,N_919);
nand U6581 (N_6581,N_1429,N_3980);
nand U6582 (N_6582,N_3174,N_1421);
or U6583 (N_6583,N_921,N_3119);
and U6584 (N_6584,N_2731,N_3922);
and U6585 (N_6585,N_711,N_4274);
and U6586 (N_6586,N_3421,N_1489);
or U6587 (N_6587,N_2220,N_1161);
nor U6588 (N_6588,N_3947,N_3475);
and U6589 (N_6589,N_1623,N_1682);
or U6590 (N_6590,N_2638,N_3994);
nand U6591 (N_6591,N_2411,N_4980);
nor U6592 (N_6592,N_2890,N_2261);
nor U6593 (N_6593,N_2165,N_4695);
nand U6594 (N_6594,N_2171,N_1495);
or U6595 (N_6595,N_2906,N_4514);
nor U6596 (N_6596,N_4134,N_1422);
nor U6597 (N_6597,N_4868,N_1100);
or U6598 (N_6598,N_4608,N_555);
or U6599 (N_6599,N_3203,N_854);
nand U6600 (N_6600,N_4221,N_3197);
nand U6601 (N_6601,N_1556,N_1858);
and U6602 (N_6602,N_991,N_4007);
nor U6603 (N_6603,N_558,N_4810);
and U6604 (N_6604,N_1490,N_4046);
nand U6605 (N_6605,N_2673,N_100);
nand U6606 (N_6606,N_630,N_4395);
nand U6607 (N_6607,N_1659,N_1098);
nor U6608 (N_6608,N_1859,N_1265);
nand U6609 (N_6609,N_2355,N_4876);
nor U6610 (N_6610,N_4345,N_1375);
nor U6611 (N_6611,N_2231,N_978);
nor U6612 (N_6612,N_1696,N_4852);
nor U6613 (N_6613,N_911,N_3539);
nand U6614 (N_6614,N_397,N_514);
or U6615 (N_6615,N_980,N_4985);
nand U6616 (N_6616,N_3670,N_3903);
nor U6617 (N_6617,N_3487,N_2727);
nor U6618 (N_6618,N_39,N_4757);
nand U6619 (N_6619,N_719,N_4780);
or U6620 (N_6620,N_2174,N_1781);
nor U6621 (N_6621,N_2645,N_2943);
nand U6622 (N_6622,N_3780,N_2910);
and U6623 (N_6623,N_999,N_483);
nand U6624 (N_6624,N_839,N_4273);
nor U6625 (N_6625,N_2164,N_4218);
nand U6626 (N_6626,N_3074,N_22);
nor U6627 (N_6627,N_4595,N_3158);
or U6628 (N_6628,N_1276,N_3966);
nand U6629 (N_6629,N_1691,N_3545);
or U6630 (N_6630,N_3898,N_2935);
nand U6631 (N_6631,N_2761,N_3189);
nor U6632 (N_6632,N_1417,N_1342);
nor U6633 (N_6633,N_2758,N_3615);
nor U6634 (N_6634,N_245,N_1584);
nand U6635 (N_6635,N_2399,N_2145);
or U6636 (N_6636,N_3222,N_3022);
nand U6637 (N_6637,N_1332,N_2969);
nand U6638 (N_6638,N_1233,N_1022);
or U6639 (N_6639,N_2942,N_433);
or U6640 (N_6640,N_1789,N_1964);
and U6641 (N_6641,N_597,N_4342);
nor U6642 (N_6642,N_3557,N_3697);
nor U6643 (N_6643,N_1282,N_351);
nand U6644 (N_6644,N_2359,N_3477);
and U6645 (N_6645,N_4916,N_4443);
and U6646 (N_6646,N_1572,N_4079);
or U6647 (N_6647,N_387,N_1379);
or U6648 (N_6648,N_2455,N_2351);
nand U6649 (N_6649,N_3017,N_4874);
and U6650 (N_6650,N_3281,N_1681);
or U6651 (N_6651,N_1785,N_1952);
nand U6652 (N_6652,N_417,N_618);
nor U6653 (N_6653,N_1993,N_4210);
and U6654 (N_6654,N_718,N_3482);
and U6655 (N_6655,N_318,N_1012);
xnor U6656 (N_6656,N_4627,N_4055);
or U6657 (N_6657,N_2433,N_1808);
nor U6658 (N_6658,N_4987,N_4157);
nor U6659 (N_6659,N_4407,N_3969);
nand U6660 (N_6660,N_166,N_366);
nand U6661 (N_6661,N_2500,N_4480);
nand U6662 (N_6662,N_1820,N_274);
nand U6663 (N_6663,N_4036,N_2191);
or U6664 (N_6664,N_1460,N_2616);
and U6665 (N_6665,N_460,N_1909);
nand U6666 (N_6666,N_4009,N_1727);
and U6667 (N_6667,N_4173,N_58);
or U6668 (N_6668,N_2268,N_2895);
nand U6669 (N_6669,N_3385,N_3079);
nor U6670 (N_6670,N_4290,N_3363);
nor U6671 (N_6671,N_4881,N_1905);
nor U6672 (N_6672,N_1078,N_236);
or U6673 (N_6673,N_4650,N_3708);
xnor U6674 (N_6674,N_950,N_3278);
nand U6675 (N_6675,N_2280,N_1404);
nor U6676 (N_6676,N_2937,N_3109);
nor U6677 (N_6677,N_1109,N_2065);
and U6678 (N_6678,N_1149,N_551);
or U6679 (N_6679,N_764,N_1904);
nor U6680 (N_6680,N_1713,N_3778);
and U6681 (N_6681,N_445,N_4620);
and U6682 (N_6682,N_137,N_588);
or U6683 (N_6683,N_918,N_1771);
nand U6684 (N_6684,N_3318,N_2134);
and U6685 (N_6685,N_179,N_3149);
and U6686 (N_6686,N_3514,N_3536);
nand U6687 (N_6687,N_3212,N_4184);
nand U6688 (N_6688,N_4004,N_4289);
nand U6689 (N_6689,N_73,N_1896);
and U6690 (N_6690,N_176,N_2697);
nand U6691 (N_6691,N_195,N_2434);
nor U6692 (N_6692,N_1381,N_3156);
or U6693 (N_6693,N_302,N_2321);
nand U6694 (N_6694,N_3680,N_4528);
and U6695 (N_6695,N_3450,N_1419);
nor U6696 (N_6696,N_3684,N_3161);
nand U6697 (N_6697,N_2086,N_1151);
nand U6698 (N_6698,N_1934,N_2495);
or U6699 (N_6699,N_3798,N_2488);
or U6700 (N_6700,N_2630,N_2706);
nand U6701 (N_6701,N_3116,N_3404);
or U6702 (N_6702,N_509,N_57);
or U6703 (N_6703,N_715,N_2984);
and U6704 (N_6704,N_3764,N_1704);
nor U6705 (N_6705,N_902,N_1004);
nor U6706 (N_6706,N_1470,N_3088);
or U6707 (N_6707,N_4638,N_4713);
nor U6708 (N_6708,N_4293,N_2371);
nand U6709 (N_6709,N_2931,N_1999);
or U6710 (N_6710,N_4646,N_2009);
or U6711 (N_6711,N_3826,N_1437);
nand U6712 (N_6712,N_3137,N_1020);
xnor U6713 (N_6713,N_3243,N_4369);
nor U6714 (N_6714,N_4291,N_563);
nand U6715 (N_6715,N_3178,N_2830);
nand U6716 (N_6716,N_754,N_2367);
nand U6717 (N_6717,N_4581,N_2237);
nand U6718 (N_6718,N_2365,N_2395);
or U6719 (N_6719,N_2604,N_4416);
or U6720 (N_6720,N_3719,N_3827);
and U6721 (N_6721,N_2940,N_4327);
and U6722 (N_6722,N_4012,N_4951);
or U6723 (N_6723,N_2269,N_757);
nor U6724 (N_6724,N_2095,N_3225);
nor U6725 (N_6725,N_2707,N_1968);
nor U6726 (N_6726,N_553,N_498);
nor U6727 (N_6727,N_1504,N_492);
nor U6728 (N_6728,N_4611,N_2011);
nand U6729 (N_6729,N_2061,N_4597);
and U6730 (N_6730,N_1982,N_1885);
and U6731 (N_6731,N_3168,N_4281);
nor U6732 (N_6732,N_674,N_2676);
nand U6733 (N_6733,N_2540,N_1669);
or U6734 (N_6734,N_866,N_4727);
nand U6735 (N_6735,N_4170,N_329);
and U6736 (N_6736,N_1922,N_841);
or U6737 (N_6737,N_4867,N_609);
and U6738 (N_6738,N_4321,N_2306);
nor U6739 (N_6739,N_626,N_2368);
nor U6740 (N_6740,N_2818,N_3877);
and U6741 (N_6741,N_1237,N_1699);
nor U6742 (N_6742,N_327,N_447);
nand U6743 (N_6743,N_3951,N_1869);
and U6744 (N_6744,N_3623,N_3907);
nor U6745 (N_6745,N_3642,N_574);
nand U6746 (N_6746,N_4836,N_1805);
nor U6747 (N_6747,N_1971,N_4880);
nor U6748 (N_6748,N_3305,N_3255);
and U6749 (N_6749,N_1866,N_4687);
and U6750 (N_6750,N_122,N_4481);
nand U6751 (N_6751,N_264,N_2845);
nor U6752 (N_6752,N_3871,N_2648);
and U6753 (N_6753,N_1479,N_1412);
nor U6754 (N_6754,N_941,N_4462);
or U6755 (N_6755,N_470,N_2051);
and U6756 (N_6756,N_3136,N_76);
nor U6757 (N_6757,N_2476,N_1285);
nand U6758 (N_6758,N_1166,N_3252);
or U6759 (N_6759,N_3408,N_1207);
or U6760 (N_6760,N_3195,N_2642);
and U6761 (N_6761,N_2374,N_4603);
or U6762 (N_6762,N_4971,N_3985);
nand U6763 (N_6763,N_336,N_3723);
or U6764 (N_6764,N_1321,N_1566);
or U6765 (N_6765,N_4828,N_3774);
and U6766 (N_6766,N_4635,N_1806);
and U6767 (N_6767,N_3115,N_1818);
or U6768 (N_6768,N_4270,N_357);
and U6769 (N_6769,N_2778,N_3375);
or U6770 (N_6770,N_79,N_2919);
or U6771 (N_6771,N_4179,N_1474);
nand U6772 (N_6772,N_1201,N_4651);
and U6773 (N_6773,N_1620,N_2575);
nor U6774 (N_6774,N_4017,N_1394);
or U6775 (N_6775,N_2974,N_2394);
and U6776 (N_6776,N_3507,N_4485);
or U6777 (N_6777,N_615,N_3713);
and U6778 (N_6778,N_2451,N_845);
and U6779 (N_6779,N_2881,N_4556);
or U6780 (N_6780,N_3592,N_3581);
or U6781 (N_6781,N_1425,N_1010);
or U6782 (N_6782,N_4400,N_32);
nand U6783 (N_6783,N_1935,N_2993);
and U6784 (N_6784,N_3756,N_2513);
nor U6785 (N_6785,N_1642,N_4494);
or U6786 (N_6786,N_1775,N_881);
nor U6787 (N_6787,N_428,N_4472);
and U6788 (N_6788,N_2383,N_2836);
and U6789 (N_6789,N_4505,N_545);
nor U6790 (N_6790,N_1175,N_1083);
nor U6791 (N_6791,N_3356,N_52);
and U6792 (N_6792,N_1816,N_1054);
nor U6793 (N_6793,N_3624,N_487);
nand U6794 (N_6794,N_2591,N_1616);
and U6795 (N_6795,N_3568,N_3867);
and U6796 (N_6796,N_3688,N_2902);
nand U6797 (N_6797,N_4093,N_499);
nand U6798 (N_6798,N_1088,N_4168);
nor U6799 (N_6799,N_3391,N_1015);
nand U6800 (N_6800,N_4888,N_3082);
nor U6801 (N_6801,N_3139,N_4860);
or U6802 (N_6802,N_298,N_1264);
and U6803 (N_6803,N_1763,N_4854);
nor U6804 (N_6804,N_1272,N_2234);
or U6805 (N_6805,N_2905,N_1601);
and U6806 (N_6806,N_4120,N_3126);
and U6807 (N_6807,N_4019,N_2539);
and U6808 (N_6808,N_3036,N_1249);
and U6809 (N_6809,N_1956,N_1354);
or U6810 (N_6810,N_3491,N_415);
nor U6811 (N_6811,N_2113,N_4356);
or U6812 (N_6812,N_4271,N_4427);
nand U6813 (N_6813,N_1787,N_530);
or U6814 (N_6814,N_1983,N_2568);
or U6815 (N_6815,N_4107,N_2012);
or U6816 (N_6816,N_144,N_1944);
or U6817 (N_6817,N_2028,N_3323);
nand U6818 (N_6818,N_4154,N_4905);
or U6819 (N_6819,N_4723,N_2090);
nand U6820 (N_6820,N_3533,N_4889);
and U6821 (N_6821,N_1513,N_1439);
nor U6822 (N_6822,N_481,N_2957);
or U6823 (N_6823,N_4775,N_3847);
or U6824 (N_6824,N_3850,N_1113);
nor U6825 (N_6825,N_2578,N_4726);
or U6826 (N_6826,N_1892,N_3051);
nor U6827 (N_6827,N_2143,N_1323);
nor U6828 (N_6828,N_2425,N_1188);
xor U6829 (N_6829,N_3874,N_3084);
and U6830 (N_6830,N_1677,N_4068);
and U6831 (N_6831,N_768,N_2085);
nor U6832 (N_6832,N_1849,N_2131);
nand U6833 (N_6833,N_1063,N_1125);
or U6834 (N_6834,N_1144,N_257);
nand U6835 (N_6835,N_2593,N_4053);
or U6836 (N_6836,N_976,N_103);
and U6837 (N_6837,N_2390,N_1013);
nand U6838 (N_6838,N_2038,N_3711);
nand U6839 (N_6839,N_1646,N_4820);
nand U6840 (N_6840,N_2718,N_2920);
nor U6841 (N_6841,N_3784,N_2419);
or U6842 (N_6842,N_2255,N_1340);
and U6843 (N_6843,N_3427,N_316);
or U6844 (N_6844,N_2200,N_51);
and U6845 (N_6845,N_350,N_1838);
and U6846 (N_6846,N_233,N_29);
or U6847 (N_6847,N_3932,N_199);
nand U6848 (N_6848,N_2699,N_1409);
or U6849 (N_6849,N_738,N_3522);
nor U6850 (N_6850,N_4551,N_364);
and U6851 (N_6851,N_590,N_223);
nor U6852 (N_6852,N_3853,N_2448);
or U6853 (N_6853,N_3635,N_3201);
nor U6854 (N_6854,N_3639,N_4401);
or U6855 (N_6855,N_293,N_2194);
nor U6856 (N_6856,N_2456,N_765);
and U6857 (N_6857,N_1864,N_4309);
nand U6858 (N_6858,N_3106,N_3193);
or U6859 (N_6859,N_4109,N_1305);
nand U6860 (N_6860,N_1596,N_198);
nor U6861 (N_6861,N_3232,N_3496);
nor U6862 (N_6862,N_1694,N_1628);
and U6863 (N_6863,N_1840,N_580);
nand U6864 (N_6864,N_2036,N_1454);
nor U6865 (N_6865,N_267,N_2861);
or U6866 (N_6866,N_4622,N_1534);
or U6867 (N_6867,N_3052,N_4920);
nand U6868 (N_6868,N_1515,N_4071);
nand U6869 (N_6869,N_1150,N_2101);
and U6870 (N_6870,N_142,N_3294);
nand U6871 (N_6871,N_621,N_3034);
nand U6872 (N_6872,N_3242,N_930);
nor U6873 (N_6873,N_4571,N_3941);
nand U6874 (N_6874,N_4919,N_824);
nor U6875 (N_6875,N_4061,N_3720);
and U6876 (N_6876,N_385,N_1738);
or U6877 (N_6877,N_167,N_2576);
nand U6878 (N_6878,N_2029,N_1452);
nor U6879 (N_6879,N_3444,N_344);
nand U6880 (N_6880,N_1251,N_131);
nor U6881 (N_6881,N_2454,N_3968);
or U6882 (N_6882,N_1979,N_1989);
and U6883 (N_6883,N_1753,N_3153);
nor U6884 (N_6884,N_1226,N_3694);
and U6885 (N_6885,N_124,N_2069);
nor U6886 (N_6886,N_4128,N_1541);
nor U6887 (N_6887,N_2010,N_3282);
and U6888 (N_6888,N_4706,N_4482);
nor U6889 (N_6889,N_1434,N_2829);
and U6890 (N_6890,N_1033,N_4198);
nand U6891 (N_6891,N_2207,N_3917);
or U6892 (N_6892,N_3609,N_374);
nor U6893 (N_6893,N_47,N_4466);
nor U6894 (N_6894,N_4444,N_2558);
or U6895 (N_6895,N_1397,N_4324);
or U6896 (N_6896,N_485,N_1737);
nand U6897 (N_6897,N_1565,N_4975);
and U6898 (N_6898,N_2004,N_3315);
nor U6899 (N_6899,N_2298,N_1378);
nor U6900 (N_6900,N_431,N_2745);
nor U6901 (N_6901,N_2897,N_905);
or U6902 (N_6902,N_4861,N_2665);
or U6903 (N_6903,N_2805,N_1583);
and U6904 (N_6904,N_2472,N_1290);
nor U6905 (N_6905,N_527,N_4000);
or U6906 (N_6906,N_4800,N_1103);
or U6907 (N_6907,N_3457,N_3154);
nor U6908 (N_6908,N_3552,N_2015);
and U6909 (N_6909,N_2315,N_4234);
or U6910 (N_6910,N_2138,N_1750);
and U6911 (N_6911,N_3992,N_2564);
nand U6912 (N_6912,N_4299,N_1032);
nand U6913 (N_6913,N_1995,N_2915);
nand U6914 (N_6914,N_4391,N_4918);
and U6915 (N_6915,N_4282,N_892);
nor U6916 (N_6916,N_2353,N_4176);
nor U6917 (N_6917,N_369,N_3776);
nand U6918 (N_6918,N_965,N_4779);
nand U6919 (N_6919,N_3555,N_1291);
nor U6920 (N_6920,N_171,N_4804);
and U6921 (N_6921,N_2824,N_797);
and U6922 (N_6922,N_2586,N_4468);
nor U6923 (N_6923,N_3577,N_2262);
and U6924 (N_6924,N_4670,N_3982);
or U6925 (N_6925,N_741,N_2621);
nand U6926 (N_6926,N_2468,N_3666);
nand U6927 (N_6927,N_526,N_4970);
and U6928 (N_6928,N_2323,N_2092);
nand U6929 (N_6929,N_3520,N_1387);
nor U6930 (N_6930,N_2951,N_2714);
nand U6931 (N_6931,N_3090,N_4990);
and U6932 (N_6932,N_1143,N_4790);
or U6933 (N_6933,N_987,N_3908);
or U6934 (N_6934,N_4848,N_3787);
and U6935 (N_6935,N_2381,N_1329);
nand U6936 (N_6936,N_1373,N_4711);
nand U6937 (N_6937,N_1931,N_1715);
nor U6938 (N_6938,N_459,N_1406);
nand U6939 (N_6939,N_2404,N_3436);
and U6940 (N_6940,N_3641,N_2022);
or U6941 (N_6941,N_2380,N_2739);
nand U6942 (N_6942,N_4247,N_2052);
nand U6943 (N_6943,N_566,N_3734);
and U6944 (N_6944,N_3285,N_776);
nand U6945 (N_6945,N_996,N_4738);
or U6946 (N_6946,N_4554,N_1693);
and U6947 (N_6947,N_4887,N_3314);
nand U6948 (N_6948,N_2023,N_126);
nor U6949 (N_6949,N_2325,N_422);
nand U6950 (N_6950,N_4377,N_2567);
and U6951 (N_6951,N_1800,N_4929);
or U6952 (N_6952,N_4030,N_353);
nor U6953 (N_6953,N_909,N_2305);
nand U6954 (N_6954,N_3013,N_1615);
nor U6955 (N_6955,N_4735,N_2924);
or U6956 (N_6956,N_434,N_3345);
nand U6957 (N_6957,N_2754,N_3979);
nor U6958 (N_6958,N_1507,N_153);
and U6959 (N_6959,N_194,N_2241);
nand U6960 (N_6960,N_1943,N_3428);
nor U6961 (N_6961,N_915,N_705);
and U6962 (N_6962,N_3807,N_4771);
nand U6963 (N_6963,N_4830,N_1986);
or U6964 (N_6964,N_284,N_156);
nor U6965 (N_6965,N_3883,N_650);
nand U6966 (N_6966,N_4490,N_4679);
or U6967 (N_6967,N_246,N_2538);
nor U6968 (N_6968,N_4778,N_2153);
and U6969 (N_6969,N_2615,N_2907);
nand U6970 (N_6970,N_6,N_3799);
xor U6971 (N_6971,N_1138,N_184);
or U6972 (N_6972,N_1835,N_3355);
nor U6973 (N_6973,N_2107,N_578);
nand U6974 (N_6974,N_4733,N_3741);
nor U6975 (N_6975,N_3984,N_1733);
and U6976 (N_6976,N_4067,N_4564);
or U6977 (N_6977,N_1442,N_3234);
nand U6978 (N_6978,N_2980,N_772);
or U6979 (N_6979,N_2408,N_3304);
nor U6980 (N_6980,N_400,N_2936);
or U6981 (N_6981,N_2393,N_480);
nand U6982 (N_6982,N_1625,N_2852);
or U6983 (N_6983,N_4623,N_4708);
and U6984 (N_6984,N_2740,N_2990);
nor U6985 (N_6985,N_4351,N_3851);
nor U6986 (N_6986,N_2810,N_3425);
nor U6987 (N_6987,N_2308,N_811);
nand U6988 (N_6988,N_3744,N_2177);
nor U6989 (N_6989,N_1487,N_3358);
nor U6990 (N_6990,N_2259,N_2909);
nor U6991 (N_6991,N_4177,N_4541);
and U6992 (N_6992,N_4729,N_2154);
nor U6993 (N_6993,N_4873,N_4890);
nand U6994 (N_6994,N_1992,N_678);
nand U6995 (N_6995,N_3476,N_3759);
nand U6996 (N_6996,N_4352,N_3377);
nor U6997 (N_6997,N_1392,N_2078);
and U6998 (N_6998,N_4082,N_4624);
nor U6999 (N_6999,N_4137,N_3078);
nand U7000 (N_7000,N_1821,N_3328);
xor U7001 (N_7001,N_1009,N_2504);
nor U7002 (N_7002,N_4279,N_4912);
nand U7003 (N_7003,N_4517,N_4822);
nand U7004 (N_7004,N_2048,N_1978);
and U7005 (N_7005,N_938,N_3043);
or U7006 (N_7006,N_2875,N_4111);
nand U7007 (N_7007,N_3721,N_4441);
nand U7008 (N_7008,N_3312,N_846);
or U7009 (N_7009,N_1006,N_4722);
and U7010 (N_7010,N_1036,N_3012);
nor U7011 (N_7011,N_4357,N_3183);
or U7012 (N_7012,N_4685,N_3471);
nor U7013 (N_7013,N_604,N_1953);
nand U7014 (N_7014,N_2239,N_3794);
or U7015 (N_7015,N_4532,N_1520);
nor U7016 (N_7016,N_111,N_2319);
and U7017 (N_7017,N_4832,N_1550);
or U7018 (N_7018,N_1891,N_4131);
nand U7019 (N_7019,N_2079,N_4133);
and U7020 (N_7020,N_1099,N_2057);
nand U7021 (N_7021,N_4590,N_1287);
nor U7022 (N_7022,N_4773,N_4242);
nor U7023 (N_7023,N_4896,N_1954);
or U7024 (N_7024,N_323,N_1730);
or U7025 (N_7025,N_3925,N_4389);
and U7026 (N_7026,N_3921,N_3852);
nand U7027 (N_7027,N_1328,N_4967);
and U7028 (N_7028,N_3732,N_3451);
or U7029 (N_7029,N_3915,N_430);
or U7030 (N_7030,N_849,N_4267);
nor U7031 (N_7031,N_2588,N_4699);
or U7032 (N_7032,N_2120,N_2210);
or U7033 (N_7033,N_1701,N_3410);
nand U7034 (N_7034,N_3352,N_4673);
and U7035 (N_7035,N_1833,N_2327);
nand U7036 (N_7036,N_3005,N_2534);
or U7037 (N_7037,N_1518,N_4922);
and U7038 (N_7038,N_4024,N_1672);
nand U7039 (N_7039,N_1874,N_392);
nor U7040 (N_7040,N_4003,N_4693);
nor U7041 (N_7041,N_917,N_831);
nor U7042 (N_7042,N_1440,N_217);
or U7043 (N_7043,N_3439,N_1918);
and U7044 (N_7044,N_914,N_3069);
nand U7045 (N_7045,N_632,N_4152);
nor U7046 (N_7046,N_129,N_3727);
or U7047 (N_7047,N_573,N_4716);
nor U7048 (N_7048,N_446,N_2442);
and U7049 (N_7049,N_595,N_1873);
nand U7050 (N_7050,N_1035,N_3342);
and U7051 (N_7051,N_4972,N_2671);
nor U7052 (N_7052,N_482,N_491);
nor U7053 (N_7053,N_3519,N_2146);
nor U7054 (N_7054,N_4744,N_1294);
or U7055 (N_7055,N_3620,N_3743);
and U7056 (N_7056,N_2149,N_2105);
and U7057 (N_7057,N_3665,N_1915);
or U7058 (N_7058,N_675,N_2933);
and U7059 (N_7059,N_1135,N_3627);
nand U7060 (N_7060,N_3040,N_4884);
nor U7061 (N_7061,N_696,N_2066);
nor U7062 (N_7062,N_1396,N_4272);
or U7063 (N_7063,N_606,N_3401);
or U7064 (N_7064,N_266,N_3048);
and U7065 (N_7065,N_4875,N_1804);
nor U7066 (N_7066,N_2982,N_4354);
nor U7067 (N_7067,N_2883,N_1280);
and U7068 (N_7068,N_2049,N_1413);
and U7069 (N_7069,N_1040,N_4542);
and U7070 (N_7070,N_1240,N_4606);
and U7071 (N_7071,N_1213,N_3566);
nor U7072 (N_7072,N_3650,N_2561);
nor U7073 (N_7073,N_2002,N_202);
or U7074 (N_7074,N_552,N_1706);
or U7075 (N_7075,N_4958,N_896);
nor U7076 (N_7076,N_1074,N_3412);
nand U7077 (N_7077,N_3902,N_4906);
and U7078 (N_7078,N_3419,N_2650);
or U7079 (N_7079,N_1023,N_3184);
and U7080 (N_7080,N_3080,N_4192);
nand U7081 (N_7081,N_1275,N_4816);
nand U7082 (N_7082,N_1001,N_1134);
nor U7083 (N_7083,N_1674,N_3020);
nand U7084 (N_7084,N_2893,N_4886);
or U7085 (N_7085,N_1266,N_1916);
or U7086 (N_7086,N_175,N_2033);
or U7087 (N_7087,N_701,N_3502);
nand U7088 (N_7088,N_2679,N_4524);
nor U7089 (N_7089,N_1973,N_4714);
nand U7090 (N_7090,N_2771,N_2680);
nor U7091 (N_7091,N_3259,N_1543);
nand U7092 (N_7092,N_2941,N_648);
and U7093 (N_7093,N_1190,N_4636);
and U7094 (N_7094,N_935,N_3151);
nor U7095 (N_7095,N_4399,N_2892);
nand U7096 (N_7096,N_771,N_3835);
and U7097 (N_7097,N_4841,N_1257);
nor U7098 (N_7098,N_1326,N_3028);
nand U7099 (N_7099,N_2743,N_3460);
nor U7100 (N_7100,N_3747,N_2627);
nand U7101 (N_7101,N_4420,N_4783);
and U7102 (N_7102,N_1552,N_4423);
and U7103 (N_7103,N_1297,N_4621);
nor U7104 (N_7104,N_1154,N_3659);
and U7105 (N_7105,N_3788,N_407);
and U7106 (N_7106,N_1695,N_4666);
or U7107 (N_7107,N_3516,N_4671);
or U7108 (N_7108,N_1521,N_3773);
or U7109 (N_7109,N_1561,N_3617);
or U7110 (N_7110,N_2244,N_2711);
nand U7111 (N_7111,N_1945,N_4295);
nor U7112 (N_7112,N_661,N_4565);
nand U7113 (N_7113,N_2423,N_1879);
and U7114 (N_7114,N_3582,N_4463);
or U7115 (N_7115,N_1228,N_562);
and U7116 (N_7116,N_3956,N_2133);
and U7117 (N_7117,N_4531,N_251);
nor U7118 (N_7118,N_906,N_1657);
and U7119 (N_7119,N_2996,N_1537);
nand U7120 (N_7120,N_4039,N_1189);
and U7121 (N_7121,N_1807,N_785);
nand U7122 (N_7122,N_4925,N_4748);
xnor U7123 (N_7123,N_676,N_1466);
nor U7124 (N_7124,N_4123,N_1500);
nor U7125 (N_7125,N_1749,N_1508);
and U7126 (N_7126,N_1247,N_2816);
nand U7127 (N_7127,N_226,N_867);
or U7128 (N_7128,N_1051,N_2724);
nor U7129 (N_7129,N_3813,N_4453);
and U7130 (N_7130,N_2790,N_2814);
or U7131 (N_7131,N_2018,N_396);
nand U7132 (N_7132,N_170,N_699);
nand U7133 (N_7133,N_1306,N_3215);
or U7134 (N_7134,N_1261,N_4821);
and U7135 (N_7135,N_951,N_269);
nand U7136 (N_7136,N_1492,N_49);
or U7137 (N_7137,N_4217,N_4118);
nand U7138 (N_7138,N_500,N_2253);
nor U7139 (N_7139,N_1502,N_3790);
and U7140 (N_7140,N_477,N_2246);
and U7141 (N_7141,N_3691,N_2751);
and U7142 (N_7142,N_1075,N_1299);
nor U7143 (N_7143,N_128,N_3560);
or U7144 (N_7144,N_2279,N_2358);
xor U7145 (N_7145,N_4512,N_972);
or U7146 (N_7146,N_4795,N_2577);
nand U7147 (N_7147,N_2283,N_2855);
nor U7148 (N_7148,N_2418,N_3553);
or U7149 (N_7149,N_4085,N_2562);
or U7150 (N_7150,N_2637,N_3924);
or U7151 (N_7151,N_2545,N_3926);
and U7152 (N_7152,N_2290,N_4587);
nor U7153 (N_7153,N_2618,N_4014);
and U7154 (N_7154,N_3038,N_1222);
or U7155 (N_7155,N_3856,N_4538);
and U7156 (N_7156,N_4813,N_4204);
nand U7157 (N_7157,N_1960,N_2363);
or U7158 (N_7158,N_7,N_4927);
nor U7159 (N_7159,N_4662,N_2853);
nor U7160 (N_7160,N_469,N_34);
and U7161 (N_7161,N_1214,N_920);
or U7162 (N_7162,N_1444,N_2928);
nor U7163 (N_7163,N_4378,N_3765);
and U7164 (N_7164,N_913,N_3053);
and U7165 (N_7165,N_3447,N_437);
xnor U7166 (N_7166,N_3722,N_283);
or U7167 (N_7167,N_1398,N_3809);
or U7168 (N_7168,N_934,N_1386);
or U7169 (N_7169,N_443,N_280);
or U7170 (N_7170,N_4323,N_2840);
or U7171 (N_7171,N_3662,N_4366);
nand U7172 (N_7172,N_937,N_3188);
nand U7173 (N_7173,N_2663,N_2517);
nand U7174 (N_7174,N_1121,N_1177);
xnor U7175 (N_7175,N_3072,N_2691);
nand U7176 (N_7176,N_3308,N_4637);
and U7177 (N_7177,N_3008,N_2912);
nor U7178 (N_7178,N_1043,N_2037);
and U7179 (N_7179,N_4949,N_1652);
or U7180 (N_7180,N_4499,N_1784);
nand U7181 (N_7181,N_2674,N_924);
or U7182 (N_7182,N_666,N_3407);
nor U7183 (N_7183,N_4006,N_3608);
nand U7184 (N_7184,N_4933,N_9);
and U7185 (N_7185,N_4562,N_2060);
and U7186 (N_7186,N_1854,N_4561);
and U7187 (N_7187,N_1884,N_4718);
and U7188 (N_7188,N_2827,N_3448);
nand U7189 (N_7189,N_2560,N_2859);
and U7190 (N_7190,N_4230,N_4185);
nand U7191 (N_7191,N_862,N_488);
and U7192 (N_7192,N_3593,N_3634);
or U7193 (N_7193,N_1600,N_28);
and U7194 (N_7194,N_3422,N_2794);
nor U7195 (N_7195,N_4935,N_2752);
nand U7196 (N_7196,N_1162,N_1769);
or U7197 (N_7197,N_4924,N_1564);
or U7198 (N_7198,N_2622,N_4022);
xor U7199 (N_7199,N_2087,N_3628);
or U7200 (N_7200,N_2660,N_4834);
nand U7201 (N_7201,N_3782,N_2180);
nor U7202 (N_7202,N_1611,N_2664);
and U7203 (N_7203,N_2396,N_3613);
and U7204 (N_7204,N_113,N_4302);
nor U7205 (N_7205,N_1718,N_4682);
and U7206 (N_7206,N_4762,N_779);
and U7207 (N_7207,N_3648,N_4902);
and U7208 (N_7208,N_2901,N_992);
nand U7209 (N_7209,N_1605,N_2178);
and U7210 (N_7210,N_102,N_561);
or U7211 (N_7211,N_3893,N_4784);
and U7212 (N_7212,N_3770,N_3182);
nand U7213 (N_7213,N_4147,N_1498);
or U7214 (N_7214,N_842,N_646);
or U7215 (N_7215,N_2173,N_1707);
nor U7216 (N_7216,N_3599,N_3086);
nand U7217 (N_7217,N_108,N_1435);
and U7218 (N_7218,N_3047,N_96);
nor U7219 (N_7219,N_1731,N_3896);
nand U7220 (N_7220,N_4652,N_484);
and U7221 (N_7221,N_3769,N_177);
nor U7222 (N_7222,N_4402,N_3155);
and U7223 (N_7223,N_343,N_1091);
or U7224 (N_7224,N_3820,N_3472);
and U7225 (N_7225,N_3640,N_3679);
nand U7226 (N_7226,N_926,N_1277);
nand U7227 (N_7227,N_1925,N_1555);
nor U7228 (N_7228,N_1523,N_2769);
nor U7229 (N_7229,N_3862,N_4197);
and U7230 (N_7230,N_3367,N_4732);
and U7231 (N_7231,N_4438,N_1336);
and U7232 (N_7232,N_796,N_1219);
or U7233 (N_7233,N_3562,N_1448);
and U7234 (N_7234,N_436,N_270);
and U7235 (N_7235,N_4372,N_1761);
nand U7236 (N_7236,N_4928,N_2432);
or U7237 (N_7237,N_2654,N_3035);
or U7238 (N_7238,N_3443,N_4837);
and U7239 (N_7239,N_1472,N_121);
and U7240 (N_7240,N_2340,N_3843);
or U7241 (N_7241,N_112,N_1031);
nor U7242 (N_7242,N_2843,N_4334);
and U7243 (N_7243,N_3027,N_2362);
nor U7244 (N_7244,N_4386,N_2821);
or U7245 (N_7245,N_1752,N_4785);
and U7246 (N_7246,N_1347,N_95);
nand U7247 (N_7247,N_617,N_4256);
nand U7248 (N_7248,N_4766,N_1676);
nor U7249 (N_7249,N_1263,N_3393);
nor U7250 (N_7250,N_4347,N_1225);
nand U7251 (N_7251,N_961,N_975);
nor U7252 (N_7252,N_2609,N_247);
nand U7253 (N_7253,N_734,N_4613);
and U7254 (N_7254,N_1223,N_3409);
and U7255 (N_7255,N_1331,N_873);
nand U7256 (N_7256,N_3268,N_3663);
or U7257 (N_7257,N_2603,N_4809);
or U7258 (N_7258,N_2703,N_276);
nand U7259 (N_7259,N_2212,N_4269);
nor U7260 (N_7260,N_807,N_74);
and U7261 (N_7261,N_4240,N_1881);
and U7262 (N_7262,N_3423,N_3824);
nand U7263 (N_7263,N_4164,N_2903);
or U7264 (N_7264,N_2217,N_3091);
and U7265 (N_7265,N_3656,N_2819);
and U7266 (N_7266,N_2285,N_602);
nor U7267 (N_7267,N_3815,N_3532);
nand U7268 (N_7268,N_4163,N_1484);
and U7269 (N_7269,N_1405,N_1758);
nand U7270 (N_7270,N_3073,N_3307);
nor U7271 (N_7271,N_4072,N_2299);
or U7272 (N_7272,N_3112,N_577);
nor U7273 (N_7273,N_2549,N_3996);
and U7274 (N_7274,N_2921,N_664);
or U7275 (N_7275,N_222,N_2623);
nand U7276 (N_7276,N_4724,N_4143);
nand U7277 (N_7277,N_3779,N_12);
nor U7278 (N_7278,N_234,N_2302);
nor U7279 (N_7279,N_3006,N_346);
nor U7280 (N_7280,N_3987,N_3205);
nand U7281 (N_7281,N_673,N_2188);
and U7282 (N_7282,N_3033,N_4313);
or U7283 (N_7283,N_3905,N_2189);
and U7284 (N_7284,N_2027,N_2888);
or U7285 (N_7285,N_69,N_1156);
and U7286 (N_7286,N_1194,N_4501);
nand U7287 (N_7287,N_1722,N_3919);
xnor U7288 (N_7288,N_3165,N_1756);
or U7289 (N_7289,N_1058,N_2019);
and U7290 (N_7290,N_2344,N_2700);
or U7291 (N_7291,N_2169,N_2379);
and U7292 (N_7292,N_4084,N_4108);
and U7293 (N_7293,N_4456,N_1268);
nand U7294 (N_7294,N_3588,N_2789);
nand U7295 (N_7295,N_4598,N_1938);
nor U7296 (N_7296,N_3265,N_3413);
nor U7297 (N_7297,N_152,N_2198);
nor U7298 (N_7298,N_1569,N_767);
and U7299 (N_7299,N_1335,N_1163);
and U7300 (N_7300,N_871,N_4243);
nor U7301 (N_7301,N_2581,N_663);
nand U7302 (N_7302,N_4336,N_777);
and U7303 (N_7303,N_1380,N_547);
or U7304 (N_7304,N_471,N_4406);
nor U7305 (N_7305,N_3760,N_3093);
or U7306 (N_7306,N_3123,N_1476);
or U7307 (N_7307,N_1522,N_4911);
nor U7308 (N_7308,N_1778,N_3);
and U7309 (N_7309,N_2934,N_88);
or U7310 (N_7310,N_48,N_4161);
or U7311 (N_7311,N_2573,N_2569);
or U7312 (N_7312,N_1825,N_3865);
or U7313 (N_7313,N_1886,N_4412);
or U7314 (N_7314,N_205,N_4390);
and U7315 (N_7315,N_1906,N_4573);
and U7316 (N_7316,N_4734,N_3831);
and U7317 (N_7317,N_2128,N_2056);
and U7318 (N_7318,N_3681,N_2566);
nor U7319 (N_7319,N_2930,N_1977);
and U7320 (N_7320,N_2481,N_50);
and U7321 (N_7321,N_1570,N_40);
nor U7322 (N_7322,N_4231,N_180);
nor U7323 (N_7323,N_1090,N_2955);
nor U7324 (N_7324,N_3260,N_4353);
nand U7325 (N_7325,N_4160,N_3906);
and U7326 (N_7326,N_2281,N_3964);
or U7327 (N_7327,N_787,N_4665);
nand U7328 (N_7328,N_4065,N_4027);
and U7329 (N_7329,N_770,N_2300);
nand U7330 (N_7330,N_3453,N_3797);
and U7331 (N_7331,N_1094,N_140);
or U7332 (N_7332,N_2899,N_4591);
and U7333 (N_7333,N_3383,N_637);
or U7334 (N_7334,N_2574,N_4040);
or U7335 (N_7335,N_440,N_1828);
nor U7336 (N_7336,N_3445,N_4205);
and U7337 (N_7337,N_952,N_647);
or U7338 (N_7338,N_3230,N_3405);
nor U7339 (N_7339,N_1899,N_3676);
and U7340 (N_7340,N_1687,N_567);
and U7341 (N_7341,N_3660,N_4476);
and U7342 (N_7342,N_2520,N_3350);
and U7343 (N_7343,N_2503,N_3117);
nand U7344 (N_7344,N_4740,N_761);
or U7345 (N_7345,N_4042,N_4520);
and U7346 (N_7346,N_2484,N_3884);
nor U7347 (N_7347,N_4411,N_4049);
nand U7348 (N_7348,N_4991,N_2698);
or U7349 (N_7349,N_4558,N_2329);
xor U7350 (N_7350,N_2730,N_1304);
nand U7351 (N_7351,N_3931,N_2236);
or U7352 (N_7352,N_3832,N_4630);
or U7353 (N_7353,N_4112,N_2848);
nor U7354 (N_7354,N_4819,N_4720);
nor U7355 (N_7355,N_2523,N_4782);
and U7356 (N_7356,N_81,N_33);
nand U7357 (N_7357,N_4457,N_2436);
xnor U7358 (N_7358,N_988,N_2343);
and U7359 (N_7359,N_395,N_1851);
nand U7360 (N_7360,N_405,N_2900);
nand U7361 (N_7361,N_3055,N_2953);
or U7362 (N_7362,N_1122,N_2376);
or U7363 (N_7363,N_3746,N_3821);
or U7364 (N_7364,N_3935,N_1286);
nor U7365 (N_7365,N_4825,N_608);
and U7366 (N_7366,N_510,N_4212);
nand U7367 (N_7367,N_3509,N_235);
and U7368 (N_7368,N_4199,N_3631);
nand U7369 (N_7369,N_2939,N_3067);
nor U7370 (N_7370,N_2971,N_864);
or U7371 (N_7371,N_1517,N_468);
or U7372 (N_7372,N_3075,N_2333);
nor U7373 (N_7373,N_324,N_472);
nand U7374 (N_7374,N_4380,N_1624);
nand U7375 (N_7375,N_1142,N_3804);
or U7376 (N_7376,N_2257,N_4759);
and U7377 (N_7377,N_1483,N_844);
and U7378 (N_7378,N_4292,N_1836);
or U7379 (N_7379,N_3431,N_1829);
or U7380 (N_7380,N_4182,N_2529);
nor U7381 (N_7381,N_114,N_3140);
nand U7382 (N_7382,N_101,N_333);
nand U7383 (N_7383,N_1582,N_185);
and U7384 (N_7384,N_13,N_1003);
nand U7385 (N_7385,N_4330,N_4823);
nand U7386 (N_7386,N_4388,N_2760);
and U7387 (N_7387,N_3039,N_535);
and U7388 (N_7388,N_4113,N_1940);
xnor U7389 (N_7389,N_448,N_458);
nand U7390 (N_7390,N_2186,N_2986);
and U7391 (N_7391,N_1917,N_3110);
nand U7392 (N_7392,N_45,N_3288);
or U7393 (N_7393,N_880,N_2736);
nor U7394 (N_7394,N_4582,N_4475);
nor U7395 (N_7395,N_3257,N_3494);
nand U7396 (N_7396,N_4091,N_4095);
nor U7397 (N_7397,N_4316,N_1540);
and U7398 (N_7398,N_2822,N_858);
xor U7399 (N_7399,N_1856,N_3014);
nand U7400 (N_7400,N_691,N_2767);
or U7401 (N_7401,N_3657,N_3937);
nand U7402 (N_7402,N_564,N_2964);
nor U7403 (N_7403,N_2465,N_746);
nand U7404 (N_7404,N_2041,N_3492);
or U7405 (N_7405,N_4408,N_2773);
nand U7406 (N_7406,N_4304,N_4451);
and U7407 (N_7407,N_1353,N_901);
nor U7408 (N_7408,N_1085,N_894);
nor U7409 (N_7409,N_1165,N_3965);
or U7410 (N_7410,N_1599,N_1776);
nor U7411 (N_7411,N_4529,N_4235);
nor U7412 (N_7412,N_4838,N_2286);
xnor U7413 (N_7413,N_3254,N_1273);
and U7414 (N_7414,N_809,N_638);
and U7415 (N_7415,N_3950,N_3587);
or U7416 (N_7416,N_2879,N_2602);
nor U7417 (N_7417,N_1139,N_43);
and U7418 (N_7418,N_4649,N_868);
nand U7419 (N_7419,N_4793,N_64);
nand U7420 (N_7420,N_1376,N_4127);
nand U7421 (N_7421,N_1311,N_2328);
and U7422 (N_7422,N_2053,N_1972);
or U7423 (N_7423,N_2916,N_4136);
nand U7424 (N_7424,N_2565,N_2157);
nand U7425 (N_7425,N_3366,N_1112);
and U7426 (N_7426,N_3118,N_3549);
xnor U7427 (N_7427,N_3261,N_813);
nand U7428 (N_7428,N_4628,N_3989);
or U7429 (N_7429,N_3848,N_828);
nand U7430 (N_7430,N_4122,N_943);
nand U7431 (N_7431,N_3524,N_2218);
and U7432 (N_7432,N_294,N_1176);
nor U7433 (N_7433,N_1637,N_1589);
or U7434 (N_7434,N_375,N_4892);
or U7435 (N_7435,N_2313,N_3689);
nor U7436 (N_7436,N_4237,N_1140);
xor U7437 (N_7437,N_4265,N_979);
nand U7438 (N_7438,N_4397,N_2527);
and U7439 (N_7439,N_63,N_1567);
nor U7440 (N_7440,N_2780,N_2632);
and U7441 (N_7441,N_4596,N_299);
nor U7442 (N_7442,N_1137,N_4307);
nor U7443 (N_7443,N_945,N_2275);
nand U7444 (N_7444,N_2522,N_4522);
or U7445 (N_7445,N_4589,N_2811);
and U7446 (N_7446,N_55,N_406);
nor U7447 (N_7447,N_4563,N_932);
and U7448 (N_7448,N_2081,N_340);
and U7449 (N_7449,N_2531,N_810);
nor U7450 (N_7450,N_4,N_3714);
and U7451 (N_7451,N_1278,N_3030);
nand U7452 (N_7452,N_4742,N_2896);
and U7453 (N_7453,N_209,N_3141);
and U7454 (N_7454,N_424,N_1998);
and U7455 (N_7455,N_4414,N_3733);
nor U7456 (N_7456,N_1216,N_4937);
or U7457 (N_7457,N_4831,N_1246);
or U7458 (N_7458,N_4090,N_3766);
nand U7459 (N_7459,N_860,N_3976);
nand U7460 (N_7460,N_189,N_3180);
nor U7461 (N_7461,N_671,N_697);
nand U7462 (N_7462,N_2849,N_803);
nand U7463 (N_7463,N_2601,N_755);
nand U7464 (N_7464,N_2702,N_3578);
or U7465 (N_7465,N_1030,N_1461);
or U7466 (N_7466,N_31,N_2001);
and U7467 (N_7467,N_441,N_946);
and U7468 (N_7468,N_3026,N_963);
nand U7469 (N_7469,N_3346,N_1428);
nor U7470 (N_7470,N_3279,N_775);
nand U7471 (N_7471,N_584,N_2119);
or U7472 (N_7472,N_689,N_15);
or U7473 (N_7473,N_4344,N_4308);
nand U7474 (N_7474,N_289,N_11);
nand U7475 (N_7475,N_4142,N_2489);
and U7476 (N_7476,N_893,N_2202);
nor U7477 (N_7477,N_3143,N_3777);
nand U7478 (N_7478,N_3060,N_3332);
nor U7479 (N_7479,N_1174,N_141);
and U7480 (N_7480,N_110,N_2965);
or U7481 (N_7481,N_4701,N_1455);
or U7482 (N_7482,N_1563,N_339);
and U7483 (N_7483,N_3751,N_1591);
nor U7484 (N_7484,N_2017,N_361);
or U7485 (N_7485,N_4115,N_1898);
nor U7486 (N_7486,N_3246,N_1114);
or U7487 (N_7487,N_78,N_87);
and U7488 (N_7488,N_3446,N_2655);
or U7489 (N_7489,N_835,N_529);
nor U7490 (N_7490,N_3501,N_888);
and U7491 (N_7491,N_3983,N_3064);
nand U7492 (N_7492,N_4570,N_158);
nand U7493 (N_7493,N_1786,N_4731);
and U7494 (N_7494,N_306,N_3646);
nor U7495 (N_7495,N_733,N_3418);
nor U7496 (N_7496,N_2096,N_4574);
nor U7497 (N_7497,N_3238,N_3432);
nand U7498 (N_7498,N_4298,N_1356);
or U7499 (N_7499,N_973,N_2382);
and U7500 (N_7500,N_1082,N_4691);
or U7501 (N_7501,N_4633,N_1631);
nand U7502 (N_7502,N_949,N_1286);
nand U7503 (N_7503,N_3669,N_2220);
nor U7504 (N_7504,N_1408,N_4067);
and U7505 (N_7505,N_2143,N_21);
or U7506 (N_7506,N_2347,N_2854);
nand U7507 (N_7507,N_4983,N_4054);
nand U7508 (N_7508,N_1782,N_3258);
and U7509 (N_7509,N_4616,N_499);
nor U7510 (N_7510,N_2366,N_2018);
nor U7511 (N_7511,N_1367,N_1314);
nand U7512 (N_7512,N_4612,N_4833);
and U7513 (N_7513,N_660,N_2778);
nand U7514 (N_7514,N_1686,N_4010);
or U7515 (N_7515,N_2538,N_1752);
nor U7516 (N_7516,N_2642,N_4382);
nand U7517 (N_7517,N_4362,N_4408);
and U7518 (N_7518,N_3255,N_4985);
and U7519 (N_7519,N_4779,N_2871);
nor U7520 (N_7520,N_1239,N_4622);
or U7521 (N_7521,N_2318,N_975);
nand U7522 (N_7522,N_27,N_3898);
nor U7523 (N_7523,N_678,N_3870);
and U7524 (N_7524,N_3114,N_4439);
or U7525 (N_7525,N_2018,N_3824);
nor U7526 (N_7526,N_4598,N_4707);
or U7527 (N_7527,N_3624,N_2888);
or U7528 (N_7528,N_471,N_3690);
nand U7529 (N_7529,N_3413,N_791);
and U7530 (N_7530,N_3757,N_685);
nor U7531 (N_7531,N_3912,N_4614);
nor U7532 (N_7532,N_314,N_2031);
nand U7533 (N_7533,N_422,N_914);
or U7534 (N_7534,N_1671,N_4930);
nand U7535 (N_7535,N_4325,N_3536);
or U7536 (N_7536,N_2300,N_3092);
nand U7537 (N_7537,N_3479,N_3663);
nor U7538 (N_7538,N_2732,N_2823);
nor U7539 (N_7539,N_1266,N_4249);
nand U7540 (N_7540,N_815,N_1142);
and U7541 (N_7541,N_1544,N_4440);
or U7542 (N_7542,N_1905,N_517);
nor U7543 (N_7543,N_2233,N_4568);
nand U7544 (N_7544,N_503,N_2146);
or U7545 (N_7545,N_2594,N_3000);
and U7546 (N_7546,N_1172,N_4868);
nor U7547 (N_7547,N_2890,N_183);
and U7548 (N_7548,N_594,N_1534);
and U7549 (N_7549,N_736,N_3182);
nand U7550 (N_7550,N_1297,N_1606);
nand U7551 (N_7551,N_1033,N_2573);
nor U7552 (N_7552,N_4740,N_3916);
or U7553 (N_7553,N_790,N_2984);
and U7554 (N_7554,N_4903,N_2919);
nor U7555 (N_7555,N_4476,N_292);
and U7556 (N_7556,N_2650,N_1876);
or U7557 (N_7557,N_1097,N_4243);
or U7558 (N_7558,N_4439,N_4661);
and U7559 (N_7559,N_54,N_2131);
nor U7560 (N_7560,N_329,N_2529);
nor U7561 (N_7561,N_4008,N_1303);
xnor U7562 (N_7562,N_3526,N_4127);
nor U7563 (N_7563,N_833,N_3162);
nand U7564 (N_7564,N_2114,N_4757);
nor U7565 (N_7565,N_3746,N_3787);
nor U7566 (N_7566,N_2838,N_4323);
and U7567 (N_7567,N_2304,N_1678);
or U7568 (N_7568,N_1896,N_2748);
nand U7569 (N_7569,N_2570,N_4303);
and U7570 (N_7570,N_963,N_3679);
or U7571 (N_7571,N_1563,N_3175);
and U7572 (N_7572,N_2687,N_939);
or U7573 (N_7573,N_2897,N_1959);
nor U7574 (N_7574,N_1530,N_2489);
nor U7575 (N_7575,N_4927,N_3388);
or U7576 (N_7576,N_1901,N_2988);
nand U7577 (N_7577,N_853,N_1223);
or U7578 (N_7578,N_4112,N_3172);
and U7579 (N_7579,N_3877,N_3669);
and U7580 (N_7580,N_479,N_1388);
or U7581 (N_7581,N_3209,N_1490);
nor U7582 (N_7582,N_861,N_1271);
nor U7583 (N_7583,N_2735,N_3170);
or U7584 (N_7584,N_16,N_187);
or U7585 (N_7585,N_65,N_4474);
or U7586 (N_7586,N_4568,N_3386);
nor U7587 (N_7587,N_1206,N_1746);
nand U7588 (N_7588,N_40,N_1738);
or U7589 (N_7589,N_3238,N_3989);
or U7590 (N_7590,N_3034,N_4287);
and U7591 (N_7591,N_540,N_141);
nor U7592 (N_7592,N_489,N_3850);
or U7593 (N_7593,N_3661,N_1391);
nor U7594 (N_7594,N_530,N_4053);
nor U7595 (N_7595,N_2289,N_890);
nor U7596 (N_7596,N_4587,N_1440);
nand U7597 (N_7597,N_2948,N_1512);
nor U7598 (N_7598,N_1273,N_3145);
nor U7599 (N_7599,N_30,N_3638);
and U7600 (N_7600,N_2543,N_3576);
and U7601 (N_7601,N_4906,N_3541);
nand U7602 (N_7602,N_1505,N_4043);
nand U7603 (N_7603,N_3328,N_2935);
and U7604 (N_7604,N_2614,N_1234);
and U7605 (N_7605,N_1335,N_1341);
nand U7606 (N_7606,N_1360,N_4810);
nand U7607 (N_7607,N_2454,N_2681);
or U7608 (N_7608,N_4981,N_2076);
nand U7609 (N_7609,N_1519,N_1278);
nor U7610 (N_7610,N_2261,N_29);
and U7611 (N_7611,N_2852,N_2114);
or U7612 (N_7612,N_210,N_1134);
and U7613 (N_7613,N_3610,N_2177);
nand U7614 (N_7614,N_1881,N_1703);
or U7615 (N_7615,N_3559,N_1243);
nand U7616 (N_7616,N_4760,N_2253);
nor U7617 (N_7617,N_3553,N_4968);
and U7618 (N_7618,N_2660,N_2896);
xnor U7619 (N_7619,N_2568,N_2695);
and U7620 (N_7620,N_488,N_88);
nor U7621 (N_7621,N_3246,N_3576);
nand U7622 (N_7622,N_4979,N_1163);
and U7623 (N_7623,N_2991,N_4160);
or U7624 (N_7624,N_3421,N_3491);
and U7625 (N_7625,N_1152,N_3812);
nand U7626 (N_7626,N_151,N_2351);
nand U7627 (N_7627,N_2427,N_2677);
nand U7628 (N_7628,N_407,N_3758);
nand U7629 (N_7629,N_4452,N_2814);
nor U7630 (N_7630,N_1576,N_1091);
nand U7631 (N_7631,N_2421,N_2265);
or U7632 (N_7632,N_2468,N_1902);
or U7633 (N_7633,N_1500,N_4880);
nor U7634 (N_7634,N_2114,N_4120);
nand U7635 (N_7635,N_4330,N_422);
or U7636 (N_7636,N_2803,N_2633);
xor U7637 (N_7637,N_4917,N_2284);
nor U7638 (N_7638,N_1480,N_4481);
and U7639 (N_7639,N_2100,N_3936);
and U7640 (N_7640,N_3835,N_1842);
nand U7641 (N_7641,N_561,N_2052);
and U7642 (N_7642,N_1639,N_4042);
nor U7643 (N_7643,N_41,N_702);
or U7644 (N_7644,N_3914,N_1036);
or U7645 (N_7645,N_2097,N_4792);
or U7646 (N_7646,N_1060,N_3125);
and U7647 (N_7647,N_2418,N_2127);
and U7648 (N_7648,N_4673,N_4791);
nor U7649 (N_7649,N_2803,N_1234);
or U7650 (N_7650,N_437,N_3316);
nand U7651 (N_7651,N_2661,N_4900);
or U7652 (N_7652,N_4253,N_3073);
nand U7653 (N_7653,N_765,N_941);
nand U7654 (N_7654,N_4224,N_4475);
nand U7655 (N_7655,N_3768,N_320);
or U7656 (N_7656,N_3980,N_3043);
nor U7657 (N_7657,N_2048,N_4436);
nor U7658 (N_7658,N_1869,N_3181);
or U7659 (N_7659,N_1698,N_2644);
nor U7660 (N_7660,N_1840,N_893);
or U7661 (N_7661,N_475,N_4383);
nor U7662 (N_7662,N_2677,N_843);
nand U7663 (N_7663,N_2320,N_3836);
and U7664 (N_7664,N_4882,N_4991);
nor U7665 (N_7665,N_1239,N_4883);
nand U7666 (N_7666,N_2004,N_2392);
nand U7667 (N_7667,N_3013,N_4184);
nand U7668 (N_7668,N_2956,N_4247);
and U7669 (N_7669,N_2954,N_2309);
or U7670 (N_7670,N_2707,N_4387);
nand U7671 (N_7671,N_2512,N_1034);
nand U7672 (N_7672,N_3527,N_1582);
nand U7673 (N_7673,N_2406,N_663);
and U7674 (N_7674,N_3779,N_3660);
nor U7675 (N_7675,N_4834,N_4712);
or U7676 (N_7676,N_772,N_1788);
or U7677 (N_7677,N_2800,N_202);
nor U7678 (N_7678,N_1403,N_2694);
nand U7679 (N_7679,N_693,N_2543);
or U7680 (N_7680,N_722,N_3996);
xor U7681 (N_7681,N_1862,N_655);
nor U7682 (N_7682,N_3619,N_4337);
and U7683 (N_7683,N_2294,N_595);
and U7684 (N_7684,N_4279,N_1772);
nand U7685 (N_7685,N_289,N_1812);
nand U7686 (N_7686,N_4434,N_1090);
nor U7687 (N_7687,N_1326,N_2206);
and U7688 (N_7688,N_895,N_232);
or U7689 (N_7689,N_3565,N_1549);
or U7690 (N_7690,N_1057,N_2275);
or U7691 (N_7691,N_2598,N_2116);
and U7692 (N_7692,N_4159,N_127);
or U7693 (N_7693,N_4860,N_4254);
nand U7694 (N_7694,N_660,N_2585);
or U7695 (N_7695,N_1172,N_431);
nand U7696 (N_7696,N_763,N_75);
or U7697 (N_7697,N_4184,N_952);
or U7698 (N_7698,N_3467,N_57);
and U7699 (N_7699,N_771,N_2661);
nand U7700 (N_7700,N_2760,N_299);
nor U7701 (N_7701,N_2365,N_3143);
and U7702 (N_7702,N_2793,N_4087);
nor U7703 (N_7703,N_1229,N_498);
nand U7704 (N_7704,N_4407,N_980);
and U7705 (N_7705,N_1581,N_4515);
nand U7706 (N_7706,N_4835,N_1858);
or U7707 (N_7707,N_227,N_4647);
and U7708 (N_7708,N_3612,N_374);
and U7709 (N_7709,N_2647,N_2539);
xor U7710 (N_7710,N_4176,N_2672);
nand U7711 (N_7711,N_4838,N_1734);
nor U7712 (N_7712,N_2160,N_1470);
nor U7713 (N_7713,N_2887,N_877);
or U7714 (N_7714,N_3145,N_2394);
nand U7715 (N_7715,N_3540,N_2229);
nand U7716 (N_7716,N_3400,N_541);
nor U7717 (N_7717,N_4608,N_4227);
and U7718 (N_7718,N_4943,N_1273);
or U7719 (N_7719,N_3257,N_4176);
or U7720 (N_7720,N_4882,N_2579);
nor U7721 (N_7721,N_597,N_3141);
or U7722 (N_7722,N_1096,N_3359);
nand U7723 (N_7723,N_2326,N_3664);
and U7724 (N_7724,N_2288,N_3891);
or U7725 (N_7725,N_3002,N_2953);
and U7726 (N_7726,N_2559,N_4501);
or U7727 (N_7727,N_1221,N_3062);
and U7728 (N_7728,N_2924,N_1772);
nor U7729 (N_7729,N_864,N_2985);
nand U7730 (N_7730,N_4942,N_4301);
nor U7731 (N_7731,N_181,N_3440);
nand U7732 (N_7732,N_2155,N_1529);
nor U7733 (N_7733,N_4987,N_350);
or U7734 (N_7734,N_520,N_2406);
nor U7735 (N_7735,N_1482,N_3765);
nand U7736 (N_7736,N_29,N_1834);
and U7737 (N_7737,N_654,N_12);
or U7738 (N_7738,N_4242,N_2013);
and U7739 (N_7739,N_1308,N_39);
and U7740 (N_7740,N_3160,N_2937);
or U7741 (N_7741,N_1016,N_2750);
nor U7742 (N_7742,N_4985,N_186);
or U7743 (N_7743,N_4315,N_1003);
nand U7744 (N_7744,N_3094,N_88);
nand U7745 (N_7745,N_4769,N_2654);
and U7746 (N_7746,N_1906,N_4745);
nand U7747 (N_7747,N_2311,N_4358);
or U7748 (N_7748,N_4074,N_4856);
and U7749 (N_7749,N_3662,N_647);
or U7750 (N_7750,N_27,N_2631);
and U7751 (N_7751,N_433,N_3069);
nor U7752 (N_7752,N_2306,N_524);
and U7753 (N_7753,N_3944,N_4117);
and U7754 (N_7754,N_1133,N_4023);
or U7755 (N_7755,N_1677,N_4943);
nor U7756 (N_7756,N_4153,N_186);
or U7757 (N_7757,N_943,N_1538);
nand U7758 (N_7758,N_2893,N_3522);
or U7759 (N_7759,N_3842,N_604);
and U7760 (N_7760,N_3591,N_1205);
nand U7761 (N_7761,N_1058,N_956);
nand U7762 (N_7762,N_2727,N_4067);
nand U7763 (N_7763,N_600,N_2344);
nand U7764 (N_7764,N_2177,N_666);
or U7765 (N_7765,N_55,N_3282);
nor U7766 (N_7766,N_908,N_1456);
and U7767 (N_7767,N_3252,N_1038);
nor U7768 (N_7768,N_3467,N_2894);
nand U7769 (N_7769,N_3631,N_4939);
and U7770 (N_7770,N_3607,N_2910);
and U7771 (N_7771,N_4293,N_2662);
nor U7772 (N_7772,N_3693,N_3164);
nand U7773 (N_7773,N_21,N_2996);
or U7774 (N_7774,N_3894,N_232);
nor U7775 (N_7775,N_1374,N_2746);
or U7776 (N_7776,N_4463,N_2549);
nor U7777 (N_7777,N_1383,N_1913);
and U7778 (N_7778,N_3619,N_4445);
nor U7779 (N_7779,N_2934,N_4187);
nor U7780 (N_7780,N_1393,N_2700);
nand U7781 (N_7781,N_470,N_3963);
and U7782 (N_7782,N_2502,N_3741);
nand U7783 (N_7783,N_3511,N_4562);
or U7784 (N_7784,N_684,N_562);
or U7785 (N_7785,N_1654,N_4405);
and U7786 (N_7786,N_3080,N_3730);
nor U7787 (N_7787,N_4576,N_3485);
nand U7788 (N_7788,N_6,N_4235);
nor U7789 (N_7789,N_4430,N_2034);
or U7790 (N_7790,N_4997,N_489);
and U7791 (N_7791,N_4470,N_1093);
or U7792 (N_7792,N_2705,N_2065);
nor U7793 (N_7793,N_3622,N_3696);
and U7794 (N_7794,N_952,N_3724);
nand U7795 (N_7795,N_2336,N_1221);
nor U7796 (N_7796,N_1219,N_3305);
and U7797 (N_7797,N_3898,N_3381);
nor U7798 (N_7798,N_3644,N_4933);
nand U7799 (N_7799,N_2333,N_2565);
nor U7800 (N_7800,N_809,N_1903);
or U7801 (N_7801,N_486,N_4371);
or U7802 (N_7802,N_3362,N_529);
or U7803 (N_7803,N_2270,N_4935);
and U7804 (N_7804,N_1556,N_3836);
nor U7805 (N_7805,N_48,N_3522);
and U7806 (N_7806,N_359,N_1690);
nand U7807 (N_7807,N_4025,N_2988);
and U7808 (N_7808,N_4363,N_1322);
nand U7809 (N_7809,N_4243,N_3446);
nand U7810 (N_7810,N_479,N_855);
nand U7811 (N_7811,N_2548,N_128);
nor U7812 (N_7812,N_1502,N_2326);
or U7813 (N_7813,N_1,N_2223);
nor U7814 (N_7814,N_41,N_2972);
nor U7815 (N_7815,N_3746,N_2008);
nand U7816 (N_7816,N_787,N_2164);
or U7817 (N_7817,N_4508,N_2151);
and U7818 (N_7818,N_1993,N_2386);
nor U7819 (N_7819,N_3015,N_1495);
nand U7820 (N_7820,N_2446,N_2007);
or U7821 (N_7821,N_3613,N_3905);
nand U7822 (N_7822,N_115,N_4591);
and U7823 (N_7823,N_4432,N_4611);
nand U7824 (N_7824,N_781,N_3746);
or U7825 (N_7825,N_520,N_2642);
or U7826 (N_7826,N_4178,N_1329);
nor U7827 (N_7827,N_4005,N_499);
or U7828 (N_7828,N_4043,N_4288);
nand U7829 (N_7829,N_4228,N_1000);
nand U7830 (N_7830,N_3957,N_2326);
or U7831 (N_7831,N_3693,N_2504);
nand U7832 (N_7832,N_3649,N_3536);
nand U7833 (N_7833,N_3122,N_1537);
nand U7834 (N_7834,N_566,N_811);
nand U7835 (N_7835,N_2087,N_3035);
nand U7836 (N_7836,N_945,N_51);
nand U7837 (N_7837,N_73,N_844);
nand U7838 (N_7838,N_2515,N_3660);
nor U7839 (N_7839,N_4542,N_1902);
nor U7840 (N_7840,N_2104,N_4412);
and U7841 (N_7841,N_827,N_2623);
and U7842 (N_7842,N_11,N_3229);
nand U7843 (N_7843,N_617,N_371);
or U7844 (N_7844,N_2664,N_1052);
or U7845 (N_7845,N_4973,N_3266);
or U7846 (N_7846,N_1196,N_2805);
nand U7847 (N_7847,N_3828,N_4088);
nand U7848 (N_7848,N_1404,N_755);
and U7849 (N_7849,N_3794,N_1959);
nor U7850 (N_7850,N_2154,N_99);
or U7851 (N_7851,N_2456,N_1201);
or U7852 (N_7852,N_3877,N_1383);
nand U7853 (N_7853,N_1986,N_1777);
and U7854 (N_7854,N_1619,N_1514);
nor U7855 (N_7855,N_252,N_3340);
nand U7856 (N_7856,N_3313,N_3053);
nor U7857 (N_7857,N_437,N_945);
and U7858 (N_7858,N_351,N_4892);
or U7859 (N_7859,N_1255,N_1648);
nor U7860 (N_7860,N_1620,N_565);
or U7861 (N_7861,N_3856,N_1334);
and U7862 (N_7862,N_3037,N_2292);
and U7863 (N_7863,N_4980,N_4186);
nor U7864 (N_7864,N_2635,N_4234);
nand U7865 (N_7865,N_4236,N_4354);
and U7866 (N_7866,N_415,N_4814);
or U7867 (N_7867,N_2118,N_1101);
nand U7868 (N_7868,N_2441,N_3217);
or U7869 (N_7869,N_1502,N_3428);
xor U7870 (N_7870,N_255,N_340);
nand U7871 (N_7871,N_4451,N_152);
or U7872 (N_7872,N_3226,N_787);
nand U7873 (N_7873,N_3147,N_3037);
or U7874 (N_7874,N_4170,N_3134);
and U7875 (N_7875,N_2915,N_1695);
nand U7876 (N_7876,N_730,N_873);
nor U7877 (N_7877,N_127,N_1580);
nor U7878 (N_7878,N_4574,N_113);
and U7879 (N_7879,N_3329,N_928);
or U7880 (N_7880,N_2183,N_1639);
xor U7881 (N_7881,N_4684,N_1140);
and U7882 (N_7882,N_276,N_2645);
and U7883 (N_7883,N_2949,N_2072);
nand U7884 (N_7884,N_3918,N_1198);
or U7885 (N_7885,N_326,N_2897);
nor U7886 (N_7886,N_1513,N_2620);
and U7887 (N_7887,N_241,N_3805);
nor U7888 (N_7888,N_2781,N_3380);
nand U7889 (N_7889,N_3576,N_3541);
nand U7890 (N_7890,N_3985,N_3406);
xnor U7891 (N_7891,N_3314,N_3726);
and U7892 (N_7892,N_1754,N_4029);
or U7893 (N_7893,N_4547,N_4817);
and U7894 (N_7894,N_585,N_3990);
nor U7895 (N_7895,N_1498,N_2009);
and U7896 (N_7896,N_132,N_1275);
and U7897 (N_7897,N_3555,N_1402);
and U7898 (N_7898,N_779,N_1902);
and U7899 (N_7899,N_4139,N_2864);
or U7900 (N_7900,N_2314,N_2328);
or U7901 (N_7901,N_150,N_2316);
and U7902 (N_7902,N_1008,N_3288);
or U7903 (N_7903,N_2400,N_4588);
nand U7904 (N_7904,N_679,N_4565);
nand U7905 (N_7905,N_4634,N_3817);
and U7906 (N_7906,N_474,N_4218);
nor U7907 (N_7907,N_826,N_3171);
nor U7908 (N_7908,N_3634,N_4651);
and U7909 (N_7909,N_453,N_2129);
and U7910 (N_7910,N_4136,N_540);
and U7911 (N_7911,N_3796,N_4456);
nor U7912 (N_7912,N_1632,N_1493);
nor U7913 (N_7913,N_1483,N_1266);
nand U7914 (N_7914,N_3970,N_3290);
nor U7915 (N_7915,N_2192,N_3275);
or U7916 (N_7916,N_1445,N_3705);
and U7917 (N_7917,N_112,N_2978);
and U7918 (N_7918,N_1586,N_2263);
and U7919 (N_7919,N_210,N_2626);
nand U7920 (N_7920,N_257,N_3575);
or U7921 (N_7921,N_4011,N_536);
nand U7922 (N_7922,N_3886,N_1332);
or U7923 (N_7923,N_4950,N_1755);
nand U7924 (N_7924,N_1683,N_1730);
or U7925 (N_7925,N_4350,N_830);
or U7926 (N_7926,N_2196,N_4766);
nand U7927 (N_7927,N_2844,N_2316);
or U7928 (N_7928,N_1076,N_744);
nor U7929 (N_7929,N_2579,N_662);
nand U7930 (N_7930,N_3556,N_4400);
and U7931 (N_7931,N_3116,N_4590);
and U7932 (N_7932,N_4916,N_4544);
nor U7933 (N_7933,N_403,N_52);
and U7934 (N_7934,N_781,N_4600);
or U7935 (N_7935,N_2737,N_3820);
nor U7936 (N_7936,N_179,N_215);
nor U7937 (N_7937,N_2015,N_3851);
nor U7938 (N_7938,N_4849,N_2076);
or U7939 (N_7939,N_1250,N_3686);
and U7940 (N_7940,N_1218,N_115);
nand U7941 (N_7941,N_3811,N_2746);
nor U7942 (N_7942,N_3707,N_4300);
nand U7943 (N_7943,N_601,N_3400);
or U7944 (N_7944,N_785,N_3368);
nand U7945 (N_7945,N_2600,N_881);
nor U7946 (N_7946,N_4178,N_180);
nor U7947 (N_7947,N_2118,N_4546);
nor U7948 (N_7948,N_1307,N_4082);
nor U7949 (N_7949,N_814,N_1287);
or U7950 (N_7950,N_2507,N_4377);
nor U7951 (N_7951,N_2879,N_268);
nand U7952 (N_7952,N_855,N_3275);
nand U7953 (N_7953,N_4401,N_4894);
nor U7954 (N_7954,N_109,N_964);
nor U7955 (N_7955,N_4574,N_1659);
and U7956 (N_7956,N_1742,N_195);
and U7957 (N_7957,N_53,N_313);
and U7958 (N_7958,N_4780,N_747);
or U7959 (N_7959,N_3106,N_674);
nand U7960 (N_7960,N_4607,N_3762);
and U7961 (N_7961,N_3190,N_3957);
and U7962 (N_7962,N_2211,N_2123);
and U7963 (N_7963,N_750,N_2486);
nand U7964 (N_7964,N_333,N_4037);
nand U7965 (N_7965,N_219,N_4195);
and U7966 (N_7966,N_1924,N_3803);
nand U7967 (N_7967,N_685,N_4892);
nand U7968 (N_7968,N_4908,N_366);
nand U7969 (N_7969,N_4347,N_2689);
nor U7970 (N_7970,N_2134,N_829);
nand U7971 (N_7971,N_3647,N_623);
and U7972 (N_7972,N_3534,N_51);
or U7973 (N_7973,N_1135,N_3215);
or U7974 (N_7974,N_1123,N_781);
nor U7975 (N_7975,N_4382,N_2365);
or U7976 (N_7976,N_3126,N_3204);
nor U7977 (N_7977,N_4402,N_1501);
and U7978 (N_7978,N_4688,N_4515);
nand U7979 (N_7979,N_4262,N_4793);
or U7980 (N_7980,N_3069,N_4264);
or U7981 (N_7981,N_154,N_3927);
nor U7982 (N_7982,N_1813,N_2263);
and U7983 (N_7983,N_4332,N_178);
and U7984 (N_7984,N_1631,N_2715);
nor U7985 (N_7985,N_3648,N_2303);
and U7986 (N_7986,N_4529,N_3330);
and U7987 (N_7987,N_217,N_923);
nor U7988 (N_7988,N_4853,N_659);
nor U7989 (N_7989,N_4264,N_4061);
nor U7990 (N_7990,N_3437,N_4379);
nor U7991 (N_7991,N_4672,N_3096);
nand U7992 (N_7992,N_1188,N_3412);
and U7993 (N_7993,N_4601,N_2572);
nor U7994 (N_7994,N_211,N_3548);
nor U7995 (N_7995,N_3428,N_2867);
nor U7996 (N_7996,N_3861,N_3668);
nand U7997 (N_7997,N_4209,N_1781);
and U7998 (N_7998,N_1545,N_3286);
and U7999 (N_7999,N_1951,N_4244);
or U8000 (N_8000,N_2050,N_2476);
nand U8001 (N_8001,N_532,N_3117);
or U8002 (N_8002,N_2265,N_618);
and U8003 (N_8003,N_4018,N_1292);
or U8004 (N_8004,N_2039,N_985);
and U8005 (N_8005,N_2185,N_4364);
nand U8006 (N_8006,N_230,N_4704);
nor U8007 (N_8007,N_2103,N_1254);
nor U8008 (N_8008,N_4770,N_2266);
or U8009 (N_8009,N_4184,N_1044);
xor U8010 (N_8010,N_4618,N_3370);
xnor U8011 (N_8011,N_3239,N_2808);
and U8012 (N_8012,N_1907,N_3180);
nor U8013 (N_8013,N_4483,N_2038);
or U8014 (N_8014,N_1228,N_1610);
and U8015 (N_8015,N_4307,N_2296);
and U8016 (N_8016,N_1789,N_3486);
nand U8017 (N_8017,N_2414,N_111);
and U8018 (N_8018,N_4386,N_1905);
nand U8019 (N_8019,N_3802,N_2777);
nand U8020 (N_8020,N_2440,N_1234);
or U8021 (N_8021,N_2407,N_2898);
nor U8022 (N_8022,N_1790,N_3597);
and U8023 (N_8023,N_4377,N_1539);
and U8024 (N_8024,N_2492,N_2162);
or U8025 (N_8025,N_1561,N_3609);
nand U8026 (N_8026,N_3529,N_1278);
nor U8027 (N_8027,N_2268,N_263);
and U8028 (N_8028,N_2487,N_2162);
nor U8029 (N_8029,N_1064,N_4773);
nor U8030 (N_8030,N_3049,N_3151);
and U8031 (N_8031,N_4695,N_461);
nand U8032 (N_8032,N_237,N_2483);
or U8033 (N_8033,N_1619,N_39);
and U8034 (N_8034,N_926,N_4119);
nor U8035 (N_8035,N_3774,N_1311);
or U8036 (N_8036,N_316,N_4600);
and U8037 (N_8037,N_3150,N_2099);
xor U8038 (N_8038,N_4336,N_2715);
xnor U8039 (N_8039,N_4018,N_4147);
and U8040 (N_8040,N_3407,N_3618);
xnor U8041 (N_8041,N_4307,N_764);
or U8042 (N_8042,N_1280,N_783);
and U8043 (N_8043,N_1886,N_1909);
nand U8044 (N_8044,N_515,N_2835);
nand U8045 (N_8045,N_291,N_822);
and U8046 (N_8046,N_4091,N_3950);
or U8047 (N_8047,N_1025,N_3332);
xnor U8048 (N_8048,N_1485,N_2448);
nand U8049 (N_8049,N_3253,N_1574);
and U8050 (N_8050,N_2503,N_221);
nand U8051 (N_8051,N_4669,N_447);
and U8052 (N_8052,N_2264,N_1583);
or U8053 (N_8053,N_4217,N_526);
nor U8054 (N_8054,N_1399,N_2580);
nand U8055 (N_8055,N_2033,N_4324);
or U8056 (N_8056,N_2997,N_2001);
nand U8057 (N_8057,N_3814,N_4597);
or U8058 (N_8058,N_350,N_1192);
or U8059 (N_8059,N_295,N_745);
nor U8060 (N_8060,N_3628,N_3318);
or U8061 (N_8061,N_4131,N_4965);
and U8062 (N_8062,N_4540,N_732);
nor U8063 (N_8063,N_3230,N_1910);
and U8064 (N_8064,N_1807,N_556);
and U8065 (N_8065,N_4025,N_3675);
nand U8066 (N_8066,N_697,N_1441);
nor U8067 (N_8067,N_1922,N_4150);
nand U8068 (N_8068,N_1249,N_310);
and U8069 (N_8069,N_534,N_405);
and U8070 (N_8070,N_605,N_1010);
nand U8071 (N_8071,N_4997,N_2747);
nor U8072 (N_8072,N_479,N_4787);
or U8073 (N_8073,N_4897,N_4036);
or U8074 (N_8074,N_1882,N_409);
nor U8075 (N_8075,N_4698,N_4608);
and U8076 (N_8076,N_4968,N_4755);
nand U8077 (N_8077,N_3902,N_4540);
or U8078 (N_8078,N_125,N_3517);
nor U8079 (N_8079,N_212,N_4238);
nor U8080 (N_8080,N_2867,N_1932);
or U8081 (N_8081,N_616,N_487);
or U8082 (N_8082,N_2193,N_4738);
or U8083 (N_8083,N_4328,N_1072);
or U8084 (N_8084,N_2613,N_2529);
or U8085 (N_8085,N_2929,N_3999);
and U8086 (N_8086,N_1960,N_236);
and U8087 (N_8087,N_1283,N_1684);
nor U8088 (N_8088,N_2776,N_4770);
and U8089 (N_8089,N_1574,N_637);
and U8090 (N_8090,N_947,N_2674);
nor U8091 (N_8091,N_2256,N_4040);
nor U8092 (N_8092,N_1450,N_386);
nand U8093 (N_8093,N_4023,N_1809);
nor U8094 (N_8094,N_4432,N_4486);
nand U8095 (N_8095,N_2577,N_321);
and U8096 (N_8096,N_3400,N_4107);
nand U8097 (N_8097,N_4860,N_4227);
or U8098 (N_8098,N_3429,N_3247);
nand U8099 (N_8099,N_2128,N_2785);
or U8100 (N_8100,N_3129,N_2695);
nand U8101 (N_8101,N_1244,N_3038);
and U8102 (N_8102,N_512,N_3895);
or U8103 (N_8103,N_2206,N_3048);
or U8104 (N_8104,N_711,N_3446);
nand U8105 (N_8105,N_993,N_729);
and U8106 (N_8106,N_998,N_3064);
nand U8107 (N_8107,N_937,N_915);
nand U8108 (N_8108,N_2096,N_2928);
nor U8109 (N_8109,N_4344,N_1084);
and U8110 (N_8110,N_3483,N_1661);
and U8111 (N_8111,N_794,N_1190);
nand U8112 (N_8112,N_2701,N_2014);
and U8113 (N_8113,N_2886,N_4044);
and U8114 (N_8114,N_4935,N_1284);
and U8115 (N_8115,N_2710,N_1004);
nor U8116 (N_8116,N_694,N_496);
or U8117 (N_8117,N_2148,N_902);
nand U8118 (N_8118,N_23,N_3787);
nand U8119 (N_8119,N_3037,N_438);
or U8120 (N_8120,N_670,N_2369);
nor U8121 (N_8121,N_2711,N_790);
or U8122 (N_8122,N_2348,N_1701);
or U8123 (N_8123,N_4277,N_1874);
or U8124 (N_8124,N_4946,N_935);
nand U8125 (N_8125,N_1541,N_2512);
and U8126 (N_8126,N_2020,N_1535);
and U8127 (N_8127,N_34,N_804);
nand U8128 (N_8128,N_1630,N_4681);
or U8129 (N_8129,N_4298,N_206);
nor U8130 (N_8130,N_4510,N_4152);
or U8131 (N_8131,N_690,N_1146);
or U8132 (N_8132,N_4014,N_201);
and U8133 (N_8133,N_2135,N_2465);
nor U8134 (N_8134,N_593,N_1575);
or U8135 (N_8135,N_2248,N_647);
and U8136 (N_8136,N_2614,N_557);
or U8137 (N_8137,N_4641,N_3604);
nor U8138 (N_8138,N_1358,N_1463);
or U8139 (N_8139,N_2438,N_646);
nand U8140 (N_8140,N_109,N_2407);
nor U8141 (N_8141,N_449,N_1938);
nor U8142 (N_8142,N_1000,N_3993);
and U8143 (N_8143,N_1580,N_1477);
or U8144 (N_8144,N_4198,N_1997);
or U8145 (N_8145,N_2596,N_1337);
and U8146 (N_8146,N_1611,N_4599);
nand U8147 (N_8147,N_4027,N_963);
or U8148 (N_8148,N_2571,N_545);
or U8149 (N_8149,N_4797,N_1506);
and U8150 (N_8150,N_3449,N_1409);
or U8151 (N_8151,N_225,N_3637);
or U8152 (N_8152,N_3865,N_3174);
or U8153 (N_8153,N_2235,N_4473);
nand U8154 (N_8154,N_54,N_1090);
and U8155 (N_8155,N_97,N_3238);
nand U8156 (N_8156,N_2558,N_386);
and U8157 (N_8157,N_2599,N_480);
nor U8158 (N_8158,N_681,N_2700);
nor U8159 (N_8159,N_3870,N_286);
or U8160 (N_8160,N_3774,N_2664);
nand U8161 (N_8161,N_2470,N_3901);
or U8162 (N_8162,N_4642,N_3904);
nor U8163 (N_8163,N_2353,N_3979);
and U8164 (N_8164,N_810,N_1552);
and U8165 (N_8165,N_3343,N_759);
nand U8166 (N_8166,N_188,N_1641);
and U8167 (N_8167,N_1726,N_3713);
xor U8168 (N_8168,N_721,N_2438);
or U8169 (N_8169,N_3673,N_1821);
nor U8170 (N_8170,N_665,N_2640);
nor U8171 (N_8171,N_2853,N_4398);
and U8172 (N_8172,N_3457,N_2307);
and U8173 (N_8173,N_431,N_1615);
and U8174 (N_8174,N_228,N_4615);
and U8175 (N_8175,N_4838,N_2504);
nand U8176 (N_8176,N_549,N_2152);
nor U8177 (N_8177,N_4647,N_1223);
nand U8178 (N_8178,N_2137,N_4908);
nor U8179 (N_8179,N_566,N_1666);
and U8180 (N_8180,N_3157,N_3335);
and U8181 (N_8181,N_2115,N_1074);
nand U8182 (N_8182,N_1534,N_2487);
or U8183 (N_8183,N_890,N_1899);
and U8184 (N_8184,N_779,N_9);
or U8185 (N_8185,N_2504,N_4231);
nor U8186 (N_8186,N_4358,N_2303);
and U8187 (N_8187,N_1323,N_4948);
or U8188 (N_8188,N_1762,N_2599);
and U8189 (N_8189,N_291,N_2947);
or U8190 (N_8190,N_2038,N_1170);
nand U8191 (N_8191,N_2020,N_1211);
or U8192 (N_8192,N_4186,N_4393);
nand U8193 (N_8193,N_2170,N_1051);
or U8194 (N_8194,N_4393,N_3515);
and U8195 (N_8195,N_1453,N_1740);
nand U8196 (N_8196,N_2528,N_2304);
nor U8197 (N_8197,N_934,N_1351);
nand U8198 (N_8198,N_243,N_2498);
or U8199 (N_8199,N_2490,N_2210);
nand U8200 (N_8200,N_4273,N_3477);
nor U8201 (N_8201,N_3126,N_1347);
or U8202 (N_8202,N_4049,N_4182);
or U8203 (N_8203,N_2464,N_2546);
nor U8204 (N_8204,N_4529,N_1996);
and U8205 (N_8205,N_3708,N_3551);
nor U8206 (N_8206,N_989,N_3786);
nand U8207 (N_8207,N_86,N_1475);
or U8208 (N_8208,N_1426,N_302);
or U8209 (N_8209,N_1324,N_3774);
and U8210 (N_8210,N_2410,N_292);
or U8211 (N_8211,N_3189,N_638);
and U8212 (N_8212,N_1703,N_3785);
and U8213 (N_8213,N_1110,N_4106);
nand U8214 (N_8214,N_2748,N_1522);
nor U8215 (N_8215,N_4388,N_3495);
nand U8216 (N_8216,N_4667,N_1001);
nand U8217 (N_8217,N_1842,N_3853);
nand U8218 (N_8218,N_581,N_2311);
nor U8219 (N_8219,N_4140,N_1855);
or U8220 (N_8220,N_2397,N_4112);
and U8221 (N_8221,N_84,N_10);
nand U8222 (N_8222,N_3168,N_900);
and U8223 (N_8223,N_1102,N_1894);
xnor U8224 (N_8224,N_2860,N_1679);
nor U8225 (N_8225,N_4424,N_1573);
or U8226 (N_8226,N_4533,N_1080);
and U8227 (N_8227,N_4042,N_4394);
and U8228 (N_8228,N_4654,N_2457);
nand U8229 (N_8229,N_2732,N_2237);
nand U8230 (N_8230,N_1793,N_3259);
and U8231 (N_8231,N_1955,N_2690);
nor U8232 (N_8232,N_4824,N_4330);
nand U8233 (N_8233,N_2408,N_1777);
or U8234 (N_8234,N_3060,N_3335);
nor U8235 (N_8235,N_4689,N_2353);
nand U8236 (N_8236,N_2631,N_3483);
nand U8237 (N_8237,N_2569,N_3410);
nand U8238 (N_8238,N_2183,N_1103);
nand U8239 (N_8239,N_1406,N_1941);
nand U8240 (N_8240,N_2550,N_316);
nor U8241 (N_8241,N_350,N_3766);
and U8242 (N_8242,N_4212,N_4126);
or U8243 (N_8243,N_2074,N_4283);
nand U8244 (N_8244,N_3792,N_4821);
or U8245 (N_8245,N_1454,N_4016);
and U8246 (N_8246,N_4446,N_756);
and U8247 (N_8247,N_3069,N_721);
or U8248 (N_8248,N_3147,N_2724);
or U8249 (N_8249,N_3074,N_1446);
nor U8250 (N_8250,N_2743,N_4580);
and U8251 (N_8251,N_1270,N_2176);
or U8252 (N_8252,N_2608,N_2234);
nand U8253 (N_8253,N_813,N_2225);
nand U8254 (N_8254,N_4893,N_2646);
xnor U8255 (N_8255,N_2756,N_1827);
nor U8256 (N_8256,N_4678,N_3267);
nand U8257 (N_8257,N_1573,N_1571);
and U8258 (N_8258,N_3347,N_4546);
and U8259 (N_8259,N_1488,N_1437);
or U8260 (N_8260,N_4246,N_2684);
and U8261 (N_8261,N_263,N_1279);
nand U8262 (N_8262,N_4977,N_2059);
nor U8263 (N_8263,N_2714,N_3309);
nor U8264 (N_8264,N_3692,N_1767);
nand U8265 (N_8265,N_2438,N_4850);
nor U8266 (N_8266,N_3498,N_112);
and U8267 (N_8267,N_3233,N_3138);
nor U8268 (N_8268,N_4425,N_4543);
nor U8269 (N_8269,N_50,N_3486);
nor U8270 (N_8270,N_2485,N_1701);
or U8271 (N_8271,N_3148,N_604);
nand U8272 (N_8272,N_2243,N_2407);
and U8273 (N_8273,N_4413,N_3368);
nand U8274 (N_8274,N_2032,N_4459);
nor U8275 (N_8275,N_3583,N_871);
and U8276 (N_8276,N_1276,N_877);
nand U8277 (N_8277,N_2442,N_1571);
or U8278 (N_8278,N_1151,N_4069);
nor U8279 (N_8279,N_4275,N_1449);
nand U8280 (N_8280,N_3810,N_4864);
nor U8281 (N_8281,N_1231,N_511);
or U8282 (N_8282,N_3723,N_4310);
nand U8283 (N_8283,N_4853,N_367);
nand U8284 (N_8284,N_1737,N_2135);
or U8285 (N_8285,N_1297,N_2047);
or U8286 (N_8286,N_4408,N_2827);
or U8287 (N_8287,N_3079,N_3721);
or U8288 (N_8288,N_4562,N_2824);
nor U8289 (N_8289,N_2796,N_2609);
nand U8290 (N_8290,N_372,N_4542);
and U8291 (N_8291,N_4870,N_359);
nand U8292 (N_8292,N_616,N_1624);
nor U8293 (N_8293,N_2177,N_3760);
or U8294 (N_8294,N_2757,N_414);
and U8295 (N_8295,N_3917,N_496);
or U8296 (N_8296,N_563,N_971);
nor U8297 (N_8297,N_926,N_1344);
nor U8298 (N_8298,N_4667,N_1257);
nor U8299 (N_8299,N_851,N_4720);
nor U8300 (N_8300,N_1580,N_3946);
and U8301 (N_8301,N_4252,N_1381);
and U8302 (N_8302,N_206,N_4319);
or U8303 (N_8303,N_752,N_3439);
or U8304 (N_8304,N_2135,N_3729);
nand U8305 (N_8305,N_80,N_4828);
nand U8306 (N_8306,N_3764,N_2144);
and U8307 (N_8307,N_1341,N_4623);
nor U8308 (N_8308,N_757,N_4403);
nand U8309 (N_8309,N_3452,N_1770);
or U8310 (N_8310,N_214,N_4365);
nand U8311 (N_8311,N_2301,N_2034);
or U8312 (N_8312,N_4557,N_31);
or U8313 (N_8313,N_1568,N_2655);
nor U8314 (N_8314,N_1496,N_3318);
nand U8315 (N_8315,N_2230,N_486);
or U8316 (N_8316,N_4134,N_3521);
or U8317 (N_8317,N_22,N_2542);
nor U8318 (N_8318,N_4800,N_2724);
nor U8319 (N_8319,N_3844,N_892);
and U8320 (N_8320,N_3158,N_3892);
nor U8321 (N_8321,N_2647,N_4240);
nand U8322 (N_8322,N_4661,N_3781);
or U8323 (N_8323,N_4575,N_2014);
nand U8324 (N_8324,N_4295,N_4329);
or U8325 (N_8325,N_677,N_1692);
or U8326 (N_8326,N_1817,N_1580);
and U8327 (N_8327,N_771,N_2202);
nor U8328 (N_8328,N_2182,N_1788);
nand U8329 (N_8329,N_3430,N_2158);
and U8330 (N_8330,N_2536,N_3024);
nor U8331 (N_8331,N_536,N_2280);
and U8332 (N_8332,N_551,N_673);
nor U8333 (N_8333,N_2627,N_3829);
and U8334 (N_8334,N_968,N_2808);
nand U8335 (N_8335,N_4305,N_1397);
or U8336 (N_8336,N_1753,N_3071);
nor U8337 (N_8337,N_3777,N_3452);
or U8338 (N_8338,N_1019,N_3050);
and U8339 (N_8339,N_1379,N_4862);
and U8340 (N_8340,N_572,N_3396);
nor U8341 (N_8341,N_2280,N_280);
nor U8342 (N_8342,N_3218,N_4675);
nand U8343 (N_8343,N_4649,N_3437);
nand U8344 (N_8344,N_2393,N_4401);
nor U8345 (N_8345,N_2252,N_4658);
or U8346 (N_8346,N_415,N_4322);
and U8347 (N_8347,N_3897,N_844);
or U8348 (N_8348,N_2420,N_3536);
or U8349 (N_8349,N_3356,N_2240);
nand U8350 (N_8350,N_1329,N_1303);
nand U8351 (N_8351,N_1887,N_1172);
and U8352 (N_8352,N_4631,N_4641);
and U8353 (N_8353,N_2996,N_1679);
nand U8354 (N_8354,N_3192,N_1429);
nor U8355 (N_8355,N_4405,N_4534);
and U8356 (N_8356,N_4666,N_2074);
and U8357 (N_8357,N_3253,N_2507);
nand U8358 (N_8358,N_4376,N_4489);
or U8359 (N_8359,N_2415,N_4052);
and U8360 (N_8360,N_1238,N_2307);
and U8361 (N_8361,N_4727,N_2660);
and U8362 (N_8362,N_1239,N_343);
and U8363 (N_8363,N_3170,N_2860);
and U8364 (N_8364,N_4830,N_47);
or U8365 (N_8365,N_1421,N_4118);
and U8366 (N_8366,N_1854,N_2509);
or U8367 (N_8367,N_2896,N_4070);
and U8368 (N_8368,N_1692,N_1406);
or U8369 (N_8369,N_2054,N_3069);
nor U8370 (N_8370,N_2754,N_3865);
or U8371 (N_8371,N_573,N_1729);
or U8372 (N_8372,N_3915,N_2639);
or U8373 (N_8373,N_1097,N_4402);
or U8374 (N_8374,N_4522,N_688);
or U8375 (N_8375,N_4501,N_1187);
nor U8376 (N_8376,N_1535,N_3149);
or U8377 (N_8377,N_222,N_2768);
nor U8378 (N_8378,N_2508,N_46);
or U8379 (N_8379,N_1308,N_1983);
and U8380 (N_8380,N_4665,N_4764);
nor U8381 (N_8381,N_3567,N_3864);
nand U8382 (N_8382,N_116,N_4087);
or U8383 (N_8383,N_4347,N_3774);
or U8384 (N_8384,N_342,N_2244);
or U8385 (N_8385,N_2808,N_713);
nor U8386 (N_8386,N_4405,N_3981);
or U8387 (N_8387,N_3906,N_4268);
nand U8388 (N_8388,N_29,N_3790);
nor U8389 (N_8389,N_4474,N_125);
or U8390 (N_8390,N_2513,N_1612);
and U8391 (N_8391,N_3532,N_2354);
and U8392 (N_8392,N_4746,N_3800);
or U8393 (N_8393,N_4056,N_231);
nor U8394 (N_8394,N_3821,N_577);
nor U8395 (N_8395,N_4845,N_3353);
and U8396 (N_8396,N_943,N_1645);
or U8397 (N_8397,N_3720,N_1600);
nand U8398 (N_8398,N_1643,N_548);
or U8399 (N_8399,N_105,N_4073);
nor U8400 (N_8400,N_1536,N_1999);
and U8401 (N_8401,N_3779,N_4145);
nand U8402 (N_8402,N_3653,N_3554);
nor U8403 (N_8403,N_3664,N_2971);
nor U8404 (N_8404,N_4227,N_2591);
and U8405 (N_8405,N_1713,N_2500);
and U8406 (N_8406,N_1660,N_1176);
nand U8407 (N_8407,N_4392,N_222);
or U8408 (N_8408,N_2180,N_4576);
nor U8409 (N_8409,N_1787,N_3549);
nor U8410 (N_8410,N_4582,N_4155);
nand U8411 (N_8411,N_416,N_4738);
nor U8412 (N_8412,N_1943,N_3216);
nor U8413 (N_8413,N_2672,N_4385);
nand U8414 (N_8414,N_1523,N_3325);
or U8415 (N_8415,N_2577,N_1431);
nand U8416 (N_8416,N_2726,N_4738);
and U8417 (N_8417,N_4242,N_4600);
nor U8418 (N_8418,N_2194,N_1850);
nand U8419 (N_8419,N_3656,N_2714);
and U8420 (N_8420,N_3852,N_1445);
nor U8421 (N_8421,N_2552,N_35);
or U8422 (N_8422,N_4586,N_2867);
and U8423 (N_8423,N_339,N_987);
or U8424 (N_8424,N_1730,N_4137);
xor U8425 (N_8425,N_2617,N_365);
nand U8426 (N_8426,N_4794,N_2379);
and U8427 (N_8427,N_3082,N_3689);
or U8428 (N_8428,N_3835,N_1257);
nor U8429 (N_8429,N_2573,N_4169);
nor U8430 (N_8430,N_624,N_308);
nand U8431 (N_8431,N_2334,N_2991);
or U8432 (N_8432,N_4753,N_215);
and U8433 (N_8433,N_3378,N_669);
or U8434 (N_8434,N_4256,N_3147);
and U8435 (N_8435,N_4102,N_1176);
nor U8436 (N_8436,N_3745,N_1705);
nor U8437 (N_8437,N_4296,N_1547);
nand U8438 (N_8438,N_4060,N_3363);
and U8439 (N_8439,N_291,N_4276);
or U8440 (N_8440,N_2077,N_1431);
and U8441 (N_8441,N_2489,N_1686);
or U8442 (N_8442,N_2507,N_927);
nand U8443 (N_8443,N_3407,N_3771);
or U8444 (N_8444,N_168,N_3517);
or U8445 (N_8445,N_8,N_4611);
nand U8446 (N_8446,N_1497,N_4332);
or U8447 (N_8447,N_1959,N_3633);
and U8448 (N_8448,N_4481,N_3626);
and U8449 (N_8449,N_434,N_4633);
or U8450 (N_8450,N_1257,N_2565);
xor U8451 (N_8451,N_2993,N_2123);
nor U8452 (N_8452,N_1732,N_4766);
or U8453 (N_8453,N_344,N_3778);
nor U8454 (N_8454,N_3824,N_4535);
nor U8455 (N_8455,N_3791,N_3836);
or U8456 (N_8456,N_1564,N_2169);
or U8457 (N_8457,N_3510,N_2953);
nor U8458 (N_8458,N_3324,N_1708);
or U8459 (N_8459,N_934,N_3939);
or U8460 (N_8460,N_480,N_4810);
nand U8461 (N_8461,N_441,N_1791);
nor U8462 (N_8462,N_3919,N_2890);
nor U8463 (N_8463,N_3075,N_3730);
nand U8464 (N_8464,N_4158,N_2372);
and U8465 (N_8465,N_1815,N_2030);
nor U8466 (N_8466,N_4889,N_257);
and U8467 (N_8467,N_3269,N_1089);
or U8468 (N_8468,N_3631,N_844);
nand U8469 (N_8469,N_1687,N_4197);
nor U8470 (N_8470,N_3723,N_4878);
nor U8471 (N_8471,N_121,N_4838);
nand U8472 (N_8472,N_2035,N_2790);
or U8473 (N_8473,N_334,N_3991);
or U8474 (N_8474,N_3075,N_1642);
and U8475 (N_8475,N_667,N_3010);
nand U8476 (N_8476,N_3183,N_269);
nand U8477 (N_8477,N_2583,N_3807);
and U8478 (N_8478,N_703,N_1093);
nand U8479 (N_8479,N_896,N_511);
or U8480 (N_8480,N_359,N_3992);
nand U8481 (N_8481,N_2955,N_1546);
and U8482 (N_8482,N_4963,N_465);
and U8483 (N_8483,N_1240,N_3586);
and U8484 (N_8484,N_4191,N_4306);
nor U8485 (N_8485,N_4555,N_312);
nand U8486 (N_8486,N_2704,N_2903);
and U8487 (N_8487,N_2329,N_662);
and U8488 (N_8488,N_2968,N_2158);
nor U8489 (N_8489,N_4357,N_2080);
nor U8490 (N_8490,N_4078,N_2466);
or U8491 (N_8491,N_717,N_3392);
xnor U8492 (N_8492,N_4271,N_3674);
nand U8493 (N_8493,N_3284,N_1485);
nand U8494 (N_8494,N_3354,N_4013);
nand U8495 (N_8495,N_757,N_454);
and U8496 (N_8496,N_2897,N_2423);
or U8497 (N_8497,N_2877,N_2621);
nand U8498 (N_8498,N_4680,N_3655);
nor U8499 (N_8499,N_3889,N_3170);
nor U8500 (N_8500,N_3863,N_3714);
nor U8501 (N_8501,N_4519,N_4058);
nand U8502 (N_8502,N_2822,N_2017);
nand U8503 (N_8503,N_1224,N_1800);
and U8504 (N_8504,N_1140,N_3286);
or U8505 (N_8505,N_2876,N_452);
nor U8506 (N_8506,N_3954,N_122);
nand U8507 (N_8507,N_456,N_2048);
and U8508 (N_8508,N_2924,N_1366);
or U8509 (N_8509,N_913,N_2768);
and U8510 (N_8510,N_4581,N_3437);
or U8511 (N_8511,N_2730,N_4060);
and U8512 (N_8512,N_3650,N_4469);
and U8513 (N_8513,N_3784,N_1049);
nor U8514 (N_8514,N_1107,N_2216);
or U8515 (N_8515,N_311,N_1563);
nand U8516 (N_8516,N_243,N_106);
nor U8517 (N_8517,N_2486,N_3134);
or U8518 (N_8518,N_2447,N_172);
nand U8519 (N_8519,N_335,N_122);
and U8520 (N_8520,N_2272,N_441);
or U8521 (N_8521,N_518,N_315);
and U8522 (N_8522,N_2726,N_115);
nor U8523 (N_8523,N_812,N_2120);
nor U8524 (N_8524,N_3858,N_2801);
or U8525 (N_8525,N_4594,N_1494);
and U8526 (N_8526,N_4331,N_1127);
or U8527 (N_8527,N_133,N_4571);
nor U8528 (N_8528,N_4921,N_3240);
nand U8529 (N_8529,N_4337,N_3476);
nand U8530 (N_8530,N_1534,N_4144);
or U8531 (N_8531,N_66,N_3924);
nand U8532 (N_8532,N_4775,N_4397);
nor U8533 (N_8533,N_1604,N_2770);
nand U8534 (N_8534,N_327,N_4459);
and U8535 (N_8535,N_4413,N_16);
and U8536 (N_8536,N_924,N_2068);
nor U8537 (N_8537,N_377,N_749);
and U8538 (N_8538,N_1252,N_1425);
nor U8539 (N_8539,N_4425,N_3932);
nand U8540 (N_8540,N_3486,N_1463);
or U8541 (N_8541,N_2545,N_4132);
xor U8542 (N_8542,N_3483,N_220);
nand U8543 (N_8543,N_4431,N_3216);
and U8544 (N_8544,N_1433,N_4137);
xnor U8545 (N_8545,N_634,N_4208);
and U8546 (N_8546,N_143,N_250);
and U8547 (N_8547,N_1143,N_2554);
or U8548 (N_8548,N_1182,N_3995);
nor U8549 (N_8549,N_3845,N_1554);
or U8550 (N_8550,N_2093,N_2208);
nand U8551 (N_8551,N_4476,N_1337);
nor U8552 (N_8552,N_3680,N_1336);
or U8553 (N_8553,N_3456,N_1693);
or U8554 (N_8554,N_2366,N_428);
nor U8555 (N_8555,N_4824,N_4347);
and U8556 (N_8556,N_1262,N_3952);
or U8557 (N_8557,N_1144,N_109);
or U8558 (N_8558,N_3519,N_2745);
nor U8559 (N_8559,N_1248,N_1339);
nand U8560 (N_8560,N_2885,N_245);
nand U8561 (N_8561,N_2884,N_2090);
nand U8562 (N_8562,N_1675,N_268);
or U8563 (N_8563,N_1001,N_2600);
or U8564 (N_8564,N_303,N_1278);
nor U8565 (N_8565,N_2265,N_2490);
or U8566 (N_8566,N_4046,N_4080);
and U8567 (N_8567,N_1044,N_1540);
and U8568 (N_8568,N_4485,N_3758);
nor U8569 (N_8569,N_2039,N_3438);
nand U8570 (N_8570,N_3055,N_287);
nand U8571 (N_8571,N_3030,N_1931);
nor U8572 (N_8572,N_75,N_4996);
or U8573 (N_8573,N_344,N_880);
nand U8574 (N_8574,N_2169,N_2054);
nand U8575 (N_8575,N_585,N_4701);
nor U8576 (N_8576,N_3843,N_4228);
nor U8577 (N_8577,N_582,N_4538);
nand U8578 (N_8578,N_3234,N_1477);
or U8579 (N_8579,N_4880,N_1645);
or U8580 (N_8580,N_1365,N_1797);
or U8581 (N_8581,N_1452,N_269);
or U8582 (N_8582,N_3018,N_2461);
or U8583 (N_8583,N_4767,N_4675);
nor U8584 (N_8584,N_565,N_1927);
or U8585 (N_8585,N_4468,N_1722);
nand U8586 (N_8586,N_2272,N_4732);
or U8587 (N_8587,N_1719,N_208);
or U8588 (N_8588,N_2858,N_3858);
and U8589 (N_8589,N_2530,N_2337);
and U8590 (N_8590,N_1094,N_4301);
and U8591 (N_8591,N_3642,N_498);
nand U8592 (N_8592,N_3532,N_1316);
and U8593 (N_8593,N_3321,N_1211);
nor U8594 (N_8594,N_2574,N_3001);
nand U8595 (N_8595,N_3961,N_2254);
nand U8596 (N_8596,N_2998,N_4216);
and U8597 (N_8597,N_1488,N_1124);
nor U8598 (N_8598,N_3788,N_4065);
nand U8599 (N_8599,N_246,N_154);
nor U8600 (N_8600,N_2376,N_3179);
nor U8601 (N_8601,N_3293,N_3757);
or U8602 (N_8602,N_3803,N_1848);
or U8603 (N_8603,N_3241,N_2956);
nand U8604 (N_8604,N_3645,N_109);
or U8605 (N_8605,N_4457,N_4909);
xor U8606 (N_8606,N_1597,N_2058);
nor U8607 (N_8607,N_3598,N_2981);
nand U8608 (N_8608,N_4987,N_564);
and U8609 (N_8609,N_557,N_3302);
or U8610 (N_8610,N_2652,N_121);
nand U8611 (N_8611,N_1679,N_3241);
or U8612 (N_8612,N_1529,N_2640);
nand U8613 (N_8613,N_2216,N_846);
or U8614 (N_8614,N_4860,N_1080);
nor U8615 (N_8615,N_4821,N_4924);
nor U8616 (N_8616,N_1050,N_4223);
nor U8617 (N_8617,N_2393,N_707);
and U8618 (N_8618,N_4893,N_641);
or U8619 (N_8619,N_4205,N_1581);
nor U8620 (N_8620,N_3073,N_1729);
nor U8621 (N_8621,N_1288,N_304);
xor U8622 (N_8622,N_2330,N_2709);
nand U8623 (N_8623,N_54,N_3734);
and U8624 (N_8624,N_693,N_2855);
and U8625 (N_8625,N_3949,N_1735);
nor U8626 (N_8626,N_1979,N_4020);
and U8627 (N_8627,N_339,N_4652);
and U8628 (N_8628,N_2597,N_2771);
or U8629 (N_8629,N_2770,N_3714);
and U8630 (N_8630,N_4288,N_704);
nand U8631 (N_8631,N_3429,N_1048);
or U8632 (N_8632,N_312,N_1613);
and U8633 (N_8633,N_4845,N_2689);
and U8634 (N_8634,N_2789,N_3333);
and U8635 (N_8635,N_4229,N_2429);
and U8636 (N_8636,N_3580,N_3196);
nor U8637 (N_8637,N_439,N_3641);
nand U8638 (N_8638,N_1153,N_3743);
nor U8639 (N_8639,N_441,N_2864);
and U8640 (N_8640,N_2710,N_3237);
nor U8641 (N_8641,N_1233,N_3849);
nand U8642 (N_8642,N_3781,N_1626);
nand U8643 (N_8643,N_1358,N_2981);
or U8644 (N_8644,N_3575,N_877);
nand U8645 (N_8645,N_4173,N_1024);
and U8646 (N_8646,N_4876,N_4623);
nor U8647 (N_8647,N_2052,N_2665);
nor U8648 (N_8648,N_2115,N_2190);
nor U8649 (N_8649,N_2204,N_1938);
and U8650 (N_8650,N_4112,N_4382);
nor U8651 (N_8651,N_1105,N_136);
nand U8652 (N_8652,N_1864,N_3012);
nand U8653 (N_8653,N_4543,N_918);
nand U8654 (N_8654,N_2989,N_357);
xor U8655 (N_8655,N_3179,N_4850);
nand U8656 (N_8656,N_1709,N_4526);
and U8657 (N_8657,N_954,N_1);
nand U8658 (N_8658,N_2957,N_298);
nor U8659 (N_8659,N_693,N_2714);
and U8660 (N_8660,N_3450,N_2348);
or U8661 (N_8661,N_1938,N_3221);
nand U8662 (N_8662,N_2117,N_4708);
nand U8663 (N_8663,N_62,N_3669);
and U8664 (N_8664,N_2412,N_3420);
nor U8665 (N_8665,N_2287,N_3517);
and U8666 (N_8666,N_4772,N_4070);
and U8667 (N_8667,N_290,N_543);
or U8668 (N_8668,N_1961,N_4965);
or U8669 (N_8669,N_888,N_2145);
nand U8670 (N_8670,N_4176,N_3062);
nor U8671 (N_8671,N_1710,N_1803);
nand U8672 (N_8672,N_3184,N_657);
nor U8673 (N_8673,N_231,N_2866);
nor U8674 (N_8674,N_1257,N_913);
nand U8675 (N_8675,N_2269,N_889);
nand U8676 (N_8676,N_343,N_4251);
and U8677 (N_8677,N_349,N_4937);
nor U8678 (N_8678,N_3093,N_3240);
and U8679 (N_8679,N_382,N_3615);
and U8680 (N_8680,N_2694,N_1962);
nor U8681 (N_8681,N_2611,N_221);
and U8682 (N_8682,N_4967,N_3135);
or U8683 (N_8683,N_2438,N_965);
nand U8684 (N_8684,N_2829,N_3797);
nand U8685 (N_8685,N_4289,N_894);
or U8686 (N_8686,N_569,N_1996);
nor U8687 (N_8687,N_4616,N_42);
nand U8688 (N_8688,N_4242,N_3434);
nand U8689 (N_8689,N_3084,N_1124);
and U8690 (N_8690,N_2569,N_3167);
nor U8691 (N_8691,N_264,N_765);
nor U8692 (N_8692,N_259,N_1122);
nor U8693 (N_8693,N_3865,N_3857);
or U8694 (N_8694,N_2858,N_571);
nand U8695 (N_8695,N_1380,N_4035);
nor U8696 (N_8696,N_3934,N_2290);
nand U8697 (N_8697,N_2314,N_3201);
and U8698 (N_8698,N_4126,N_657);
nor U8699 (N_8699,N_399,N_3925);
nand U8700 (N_8700,N_1890,N_3790);
nand U8701 (N_8701,N_2720,N_1648);
and U8702 (N_8702,N_4580,N_1648);
nand U8703 (N_8703,N_3264,N_3687);
and U8704 (N_8704,N_224,N_2098);
and U8705 (N_8705,N_4348,N_4092);
and U8706 (N_8706,N_1192,N_752);
and U8707 (N_8707,N_3221,N_555);
and U8708 (N_8708,N_2236,N_1420);
or U8709 (N_8709,N_2578,N_2241);
nor U8710 (N_8710,N_2059,N_1207);
nor U8711 (N_8711,N_3,N_1085);
nand U8712 (N_8712,N_551,N_2446);
or U8713 (N_8713,N_338,N_3549);
nor U8714 (N_8714,N_1755,N_4435);
nor U8715 (N_8715,N_4910,N_4550);
xnor U8716 (N_8716,N_1782,N_641);
nand U8717 (N_8717,N_2899,N_2060);
nor U8718 (N_8718,N_600,N_1382);
nand U8719 (N_8719,N_109,N_607);
and U8720 (N_8720,N_1757,N_2149);
nand U8721 (N_8721,N_3253,N_4896);
or U8722 (N_8722,N_1071,N_4863);
and U8723 (N_8723,N_4752,N_4045);
nor U8724 (N_8724,N_945,N_4009);
nand U8725 (N_8725,N_2432,N_3483);
and U8726 (N_8726,N_585,N_3890);
or U8727 (N_8727,N_852,N_1739);
nand U8728 (N_8728,N_775,N_3973);
xnor U8729 (N_8729,N_4727,N_1676);
nand U8730 (N_8730,N_2245,N_878);
and U8731 (N_8731,N_3419,N_4483);
or U8732 (N_8732,N_227,N_1936);
or U8733 (N_8733,N_4534,N_4962);
and U8734 (N_8734,N_520,N_1169);
and U8735 (N_8735,N_3145,N_632);
and U8736 (N_8736,N_130,N_2158);
nand U8737 (N_8737,N_87,N_3605);
and U8738 (N_8738,N_3176,N_134);
and U8739 (N_8739,N_1614,N_3591);
nand U8740 (N_8740,N_3937,N_2684);
and U8741 (N_8741,N_3473,N_1833);
nor U8742 (N_8742,N_966,N_544);
and U8743 (N_8743,N_3516,N_581);
or U8744 (N_8744,N_3191,N_294);
nand U8745 (N_8745,N_4040,N_1641);
nor U8746 (N_8746,N_4700,N_3522);
or U8747 (N_8747,N_2978,N_3379);
xnor U8748 (N_8748,N_2565,N_4768);
nand U8749 (N_8749,N_136,N_3602);
nor U8750 (N_8750,N_2768,N_2171);
nor U8751 (N_8751,N_1503,N_4832);
nand U8752 (N_8752,N_4119,N_3642);
xor U8753 (N_8753,N_2083,N_2428);
or U8754 (N_8754,N_675,N_4176);
nor U8755 (N_8755,N_3276,N_3256);
and U8756 (N_8756,N_3603,N_3137);
or U8757 (N_8757,N_574,N_2825);
or U8758 (N_8758,N_1685,N_3436);
and U8759 (N_8759,N_552,N_4630);
and U8760 (N_8760,N_4051,N_2251);
nor U8761 (N_8761,N_4526,N_201);
nor U8762 (N_8762,N_1851,N_128);
and U8763 (N_8763,N_3529,N_1944);
nand U8764 (N_8764,N_2970,N_462);
or U8765 (N_8765,N_2905,N_19);
nor U8766 (N_8766,N_4200,N_3492);
and U8767 (N_8767,N_1832,N_1703);
and U8768 (N_8768,N_2918,N_2986);
nand U8769 (N_8769,N_3169,N_3955);
and U8770 (N_8770,N_514,N_1115);
or U8771 (N_8771,N_3388,N_2216);
and U8772 (N_8772,N_584,N_4625);
nand U8773 (N_8773,N_659,N_3005);
nor U8774 (N_8774,N_3452,N_1309);
nand U8775 (N_8775,N_958,N_1701);
nor U8776 (N_8776,N_359,N_2900);
nor U8777 (N_8777,N_3775,N_720);
and U8778 (N_8778,N_1305,N_1552);
or U8779 (N_8779,N_3142,N_141);
and U8780 (N_8780,N_222,N_4475);
nand U8781 (N_8781,N_2138,N_520);
nor U8782 (N_8782,N_2375,N_3893);
and U8783 (N_8783,N_1893,N_1013);
nor U8784 (N_8784,N_4629,N_3811);
nand U8785 (N_8785,N_4446,N_2694);
and U8786 (N_8786,N_1549,N_2755);
or U8787 (N_8787,N_4655,N_53);
nor U8788 (N_8788,N_2330,N_2967);
or U8789 (N_8789,N_732,N_2640);
and U8790 (N_8790,N_973,N_4585);
and U8791 (N_8791,N_3654,N_1351);
nand U8792 (N_8792,N_49,N_593);
and U8793 (N_8793,N_1180,N_3482);
nand U8794 (N_8794,N_4922,N_4809);
nand U8795 (N_8795,N_3699,N_3312);
or U8796 (N_8796,N_3499,N_3667);
or U8797 (N_8797,N_3748,N_1962);
and U8798 (N_8798,N_4116,N_1269);
and U8799 (N_8799,N_2494,N_547);
nor U8800 (N_8800,N_2999,N_1393);
nand U8801 (N_8801,N_4895,N_3764);
or U8802 (N_8802,N_1059,N_2544);
nor U8803 (N_8803,N_4550,N_1692);
or U8804 (N_8804,N_296,N_429);
or U8805 (N_8805,N_4068,N_3587);
nand U8806 (N_8806,N_3976,N_1642);
nor U8807 (N_8807,N_2042,N_4759);
nor U8808 (N_8808,N_1400,N_4111);
nand U8809 (N_8809,N_3188,N_2919);
nand U8810 (N_8810,N_3093,N_1157);
and U8811 (N_8811,N_402,N_257);
or U8812 (N_8812,N_663,N_1479);
nor U8813 (N_8813,N_945,N_1590);
nand U8814 (N_8814,N_88,N_2221);
and U8815 (N_8815,N_435,N_1648);
nand U8816 (N_8816,N_4304,N_2215);
or U8817 (N_8817,N_3505,N_3066);
or U8818 (N_8818,N_3560,N_3446);
nand U8819 (N_8819,N_1203,N_4499);
and U8820 (N_8820,N_1580,N_1869);
nand U8821 (N_8821,N_3901,N_2830);
nor U8822 (N_8822,N_1607,N_1723);
and U8823 (N_8823,N_3226,N_234);
and U8824 (N_8824,N_559,N_137);
and U8825 (N_8825,N_2496,N_2242);
nand U8826 (N_8826,N_3504,N_1866);
nor U8827 (N_8827,N_3284,N_1043);
or U8828 (N_8828,N_4403,N_1034);
and U8829 (N_8829,N_108,N_1207);
and U8830 (N_8830,N_2784,N_4284);
or U8831 (N_8831,N_1992,N_2895);
and U8832 (N_8832,N_219,N_514);
nand U8833 (N_8833,N_1628,N_2925);
nand U8834 (N_8834,N_4154,N_997);
nor U8835 (N_8835,N_43,N_1711);
or U8836 (N_8836,N_4634,N_1779);
nor U8837 (N_8837,N_1635,N_2019);
nor U8838 (N_8838,N_817,N_953);
and U8839 (N_8839,N_769,N_898);
and U8840 (N_8840,N_1554,N_3069);
and U8841 (N_8841,N_3340,N_4622);
nand U8842 (N_8842,N_1100,N_3933);
nand U8843 (N_8843,N_1945,N_1634);
nand U8844 (N_8844,N_4992,N_920);
nand U8845 (N_8845,N_2984,N_3027);
nand U8846 (N_8846,N_1071,N_810);
nor U8847 (N_8847,N_1255,N_1471);
or U8848 (N_8848,N_3772,N_4520);
or U8849 (N_8849,N_4164,N_3135);
and U8850 (N_8850,N_4685,N_3344);
nor U8851 (N_8851,N_4128,N_3979);
and U8852 (N_8852,N_364,N_317);
and U8853 (N_8853,N_4287,N_239);
nor U8854 (N_8854,N_998,N_4245);
and U8855 (N_8855,N_2066,N_1591);
or U8856 (N_8856,N_2730,N_3246);
or U8857 (N_8857,N_3817,N_4366);
and U8858 (N_8858,N_4996,N_2057);
and U8859 (N_8859,N_4290,N_552);
nand U8860 (N_8860,N_3901,N_2489);
and U8861 (N_8861,N_2458,N_612);
nor U8862 (N_8862,N_4477,N_3778);
and U8863 (N_8863,N_1277,N_818);
and U8864 (N_8864,N_4246,N_1413);
nand U8865 (N_8865,N_2755,N_4663);
or U8866 (N_8866,N_4723,N_708);
and U8867 (N_8867,N_3159,N_3955);
nor U8868 (N_8868,N_4820,N_3003);
or U8869 (N_8869,N_978,N_2470);
and U8870 (N_8870,N_2178,N_2411);
nor U8871 (N_8871,N_2423,N_3442);
and U8872 (N_8872,N_4200,N_2388);
nand U8873 (N_8873,N_237,N_2681);
nor U8874 (N_8874,N_54,N_3718);
nand U8875 (N_8875,N_2266,N_4258);
nand U8876 (N_8876,N_2645,N_1737);
nand U8877 (N_8877,N_2344,N_2943);
and U8878 (N_8878,N_2072,N_3139);
and U8879 (N_8879,N_2922,N_860);
or U8880 (N_8880,N_2471,N_2056);
and U8881 (N_8881,N_4138,N_4695);
nand U8882 (N_8882,N_1509,N_3132);
and U8883 (N_8883,N_4342,N_2341);
or U8884 (N_8884,N_401,N_1059);
and U8885 (N_8885,N_1369,N_3375);
and U8886 (N_8886,N_2984,N_2170);
nand U8887 (N_8887,N_4916,N_4840);
nand U8888 (N_8888,N_1954,N_2328);
or U8889 (N_8889,N_401,N_3571);
or U8890 (N_8890,N_1534,N_2943);
or U8891 (N_8891,N_4813,N_2048);
nand U8892 (N_8892,N_2816,N_3739);
xor U8893 (N_8893,N_4062,N_4021);
or U8894 (N_8894,N_4720,N_931);
nand U8895 (N_8895,N_3487,N_1480);
nor U8896 (N_8896,N_1359,N_1915);
nor U8897 (N_8897,N_480,N_4444);
nand U8898 (N_8898,N_1548,N_1181);
or U8899 (N_8899,N_2748,N_4768);
or U8900 (N_8900,N_3506,N_590);
nand U8901 (N_8901,N_1947,N_3513);
nor U8902 (N_8902,N_1130,N_3549);
and U8903 (N_8903,N_2491,N_931);
or U8904 (N_8904,N_596,N_2903);
nand U8905 (N_8905,N_4783,N_1255);
and U8906 (N_8906,N_3743,N_927);
and U8907 (N_8907,N_2367,N_399);
nor U8908 (N_8908,N_480,N_2);
nor U8909 (N_8909,N_4990,N_3085);
nand U8910 (N_8910,N_951,N_1198);
and U8911 (N_8911,N_1509,N_463);
or U8912 (N_8912,N_3143,N_3625);
nor U8913 (N_8913,N_3740,N_3641);
and U8914 (N_8914,N_2604,N_3557);
and U8915 (N_8915,N_4820,N_2059);
nor U8916 (N_8916,N_3019,N_4532);
nor U8917 (N_8917,N_102,N_4726);
nand U8918 (N_8918,N_4812,N_2099);
nand U8919 (N_8919,N_4720,N_3308);
nor U8920 (N_8920,N_4927,N_3889);
or U8921 (N_8921,N_1222,N_3745);
or U8922 (N_8922,N_145,N_3315);
nor U8923 (N_8923,N_4879,N_3628);
and U8924 (N_8924,N_26,N_3537);
nand U8925 (N_8925,N_4526,N_2394);
or U8926 (N_8926,N_4416,N_1428);
nand U8927 (N_8927,N_4696,N_4452);
or U8928 (N_8928,N_4586,N_1785);
nand U8929 (N_8929,N_3372,N_1033);
and U8930 (N_8930,N_4007,N_2814);
nand U8931 (N_8931,N_3927,N_1636);
and U8932 (N_8932,N_741,N_2422);
and U8933 (N_8933,N_4432,N_3660);
xnor U8934 (N_8934,N_4202,N_1144);
nor U8935 (N_8935,N_2259,N_2367);
xor U8936 (N_8936,N_1055,N_3129);
and U8937 (N_8937,N_2395,N_2087);
or U8938 (N_8938,N_3215,N_296);
or U8939 (N_8939,N_4108,N_502);
or U8940 (N_8940,N_4029,N_3362);
or U8941 (N_8941,N_4973,N_2628);
nand U8942 (N_8942,N_4434,N_3303);
or U8943 (N_8943,N_856,N_3356);
and U8944 (N_8944,N_3938,N_2730);
and U8945 (N_8945,N_3267,N_1984);
nor U8946 (N_8946,N_1233,N_1619);
nor U8947 (N_8947,N_3308,N_285);
and U8948 (N_8948,N_976,N_3745);
nand U8949 (N_8949,N_40,N_4162);
or U8950 (N_8950,N_3478,N_4008);
nand U8951 (N_8951,N_1695,N_320);
nand U8952 (N_8952,N_2516,N_4428);
or U8953 (N_8953,N_2405,N_1402);
nand U8954 (N_8954,N_3963,N_365);
nor U8955 (N_8955,N_757,N_4349);
nand U8956 (N_8956,N_2387,N_1713);
and U8957 (N_8957,N_4610,N_3325);
nand U8958 (N_8958,N_2777,N_4626);
nand U8959 (N_8959,N_2929,N_1080);
nor U8960 (N_8960,N_4437,N_1398);
and U8961 (N_8961,N_2924,N_3);
and U8962 (N_8962,N_2589,N_1188);
nor U8963 (N_8963,N_3589,N_4006);
nor U8964 (N_8964,N_1970,N_4536);
nor U8965 (N_8965,N_1234,N_4485);
nand U8966 (N_8966,N_1306,N_2057);
or U8967 (N_8967,N_112,N_3314);
or U8968 (N_8968,N_2656,N_1970);
or U8969 (N_8969,N_156,N_961);
or U8970 (N_8970,N_3394,N_4220);
xor U8971 (N_8971,N_2601,N_2115);
nand U8972 (N_8972,N_4696,N_77);
or U8973 (N_8973,N_1648,N_1365);
or U8974 (N_8974,N_1186,N_3859);
or U8975 (N_8975,N_2655,N_3804);
or U8976 (N_8976,N_1759,N_1020);
or U8977 (N_8977,N_4448,N_686);
nand U8978 (N_8978,N_579,N_4689);
or U8979 (N_8979,N_4423,N_703);
and U8980 (N_8980,N_305,N_3404);
or U8981 (N_8981,N_2762,N_4208);
and U8982 (N_8982,N_2262,N_3943);
nand U8983 (N_8983,N_1298,N_4104);
and U8984 (N_8984,N_2328,N_2246);
and U8985 (N_8985,N_881,N_3348);
nor U8986 (N_8986,N_1604,N_3710);
and U8987 (N_8987,N_73,N_2342);
and U8988 (N_8988,N_3754,N_1966);
or U8989 (N_8989,N_2040,N_4046);
nand U8990 (N_8990,N_2488,N_3054);
or U8991 (N_8991,N_4226,N_1045);
and U8992 (N_8992,N_4135,N_2903);
and U8993 (N_8993,N_4399,N_167);
and U8994 (N_8994,N_1833,N_1831);
nand U8995 (N_8995,N_1340,N_1359);
or U8996 (N_8996,N_1183,N_997);
and U8997 (N_8997,N_489,N_3215);
or U8998 (N_8998,N_1517,N_3158);
xor U8999 (N_8999,N_584,N_3091);
nor U9000 (N_9000,N_4474,N_3579);
nand U9001 (N_9001,N_66,N_2790);
and U9002 (N_9002,N_2364,N_4621);
and U9003 (N_9003,N_2762,N_4368);
nand U9004 (N_9004,N_3691,N_2797);
nand U9005 (N_9005,N_3439,N_3302);
and U9006 (N_9006,N_2275,N_1999);
and U9007 (N_9007,N_136,N_1393);
nor U9008 (N_9008,N_4075,N_2729);
and U9009 (N_9009,N_4005,N_1307);
and U9010 (N_9010,N_965,N_318);
and U9011 (N_9011,N_3203,N_1990);
nor U9012 (N_9012,N_3995,N_4535);
or U9013 (N_9013,N_3946,N_3723);
nor U9014 (N_9014,N_4976,N_1010);
or U9015 (N_9015,N_2410,N_4663);
nor U9016 (N_9016,N_3686,N_1832);
and U9017 (N_9017,N_2925,N_1510);
nand U9018 (N_9018,N_2072,N_2335);
or U9019 (N_9019,N_3514,N_2304);
nor U9020 (N_9020,N_2733,N_3941);
and U9021 (N_9021,N_821,N_2451);
nor U9022 (N_9022,N_4237,N_542);
nand U9023 (N_9023,N_2707,N_4931);
or U9024 (N_9024,N_121,N_961);
nor U9025 (N_9025,N_861,N_36);
or U9026 (N_9026,N_1105,N_2735);
and U9027 (N_9027,N_3728,N_1155);
nor U9028 (N_9028,N_3955,N_3334);
nor U9029 (N_9029,N_4876,N_875);
nor U9030 (N_9030,N_3508,N_715);
and U9031 (N_9031,N_3250,N_4276);
and U9032 (N_9032,N_89,N_4556);
and U9033 (N_9033,N_4223,N_1695);
and U9034 (N_9034,N_2977,N_2928);
nor U9035 (N_9035,N_651,N_1060);
nand U9036 (N_9036,N_593,N_599);
and U9037 (N_9037,N_1079,N_1400);
nor U9038 (N_9038,N_947,N_4687);
nor U9039 (N_9039,N_2757,N_2108);
or U9040 (N_9040,N_2077,N_2913);
nand U9041 (N_9041,N_310,N_583);
nor U9042 (N_9042,N_4935,N_1909);
nand U9043 (N_9043,N_1403,N_1487);
or U9044 (N_9044,N_1917,N_1254);
nor U9045 (N_9045,N_3059,N_799);
nand U9046 (N_9046,N_585,N_1493);
and U9047 (N_9047,N_711,N_3090);
nor U9048 (N_9048,N_2432,N_3907);
or U9049 (N_9049,N_1016,N_4570);
or U9050 (N_9050,N_4321,N_2962);
nand U9051 (N_9051,N_3909,N_777);
or U9052 (N_9052,N_4592,N_3495);
or U9053 (N_9053,N_4177,N_3731);
nand U9054 (N_9054,N_3756,N_578);
nor U9055 (N_9055,N_1421,N_2767);
or U9056 (N_9056,N_330,N_3380);
or U9057 (N_9057,N_4961,N_2227);
xor U9058 (N_9058,N_3240,N_4124);
nand U9059 (N_9059,N_4706,N_581);
or U9060 (N_9060,N_3781,N_4530);
and U9061 (N_9061,N_2582,N_3669);
nor U9062 (N_9062,N_676,N_1070);
nand U9063 (N_9063,N_651,N_2798);
nand U9064 (N_9064,N_853,N_2025);
and U9065 (N_9065,N_4886,N_1570);
nor U9066 (N_9066,N_1322,N_3855);
nand U9067 (N_9067,N_2671,N_4212);
nor U9068 (N_9068,N_3314,N_2217);
and U9069 (N_9069,N_3492,N_2665);
and U9070 (N_9070,N_1132,N_2749);
nor U9071 (N_9071,N_3516,N_2215);
nand U9072 (N_9072,N_1153,N_4148);
nor U9073 (N_9073,N_1212,N_57);
nor U9074 (N_9074,N_4856,N_3819);
or U9075 (N_9075,N_3525,N_2661);
and U9076 (N_9076,N_2252,N_1289);
nor U9077 (N_9077,N_3733,N_766);
nand U9078 (N_9078,N_2707,N_4227);
nor U9079 (N_9079,N_2101,N_4765);
or U9080 (N_9080,N_4015,N_1610);
nand U9081 (N_9081,N_4705,N_2388);
and U9082 (N_9082,N_463,N_4254);
nand U9083 (N_9083,N_1857,N_1772);
and U9084 (N_9084,N_3076,N_3347);
nor U9085 (N_9085,N_2988,N_1117);
nor U9086 (N_9086,N_1519,N_957);
or U9087 (N_9087,N_4023,N_3534);
or U9088 (N_9088,N_651,N_918);
or U9089 (N_9089,N_607,N_3540);
nor U9090 (N_9090,N_3766,N_1489);
and U9091 (N_9091,N_1847,N_1440);
or U9092 (N_9092,N_744,N_147);
nand U9093 (N_9093,N_223,N_3961);
nor U9094 (N_9094,N_3389,N_295);
nand U9095 (N_9095,N_2193,N_1357);
nand U9096 (N_9096,N_1490,N_1143);
nand U9097 (N_9097,N_2409,N_2368);
or U9098 (N_9098,N_979,N_4718);
nor U9099 (N_9099,N_886,N_290);
or U9100 (N_9100,N_1339,N_1288);
nor U9101 (N_9101,N_3445,N_969);
nor U9102 (N_9102,N_2661,N_3096);
or U9103 (N_9103,N_2382,N_203);
nor U9104 (N_9104,N_3779,N_3713);
or U9105 (N_9105,N_830,N_3270);
and U9106 (N_9106,N_161,N_3084);
and U9107 (N_9107,N_3209,N_2773);
or U9108 (N_9108,N_4989,N_1375);
or U9109 (N_9109,N_432,N_2527);
or U9110 (N_9110,N_1480,N_3484);
nand U9111 (N_9111,N_2190,N_3178);
or U9112 (N_9112,N_1811,N_3130);
nand U9113 (N_9113,N_288,N_1830);
nor U9114 (N_9114,N_804,N_2538);
nor U9115 (N_9115,N_4555,N_4782);
nand U9116 (N_9116,N_2706,N_4361);
nor U9117 (N_9117,N_3019,N_401);
and U9118 (N_9118,N_843,N_3631);
or U9119 (N_9119,N_3970,N_2179);
nor U9120 (N_9120,N_4209,N_4967);
nor U9121 (N_9121,N_3439,N_1178);
nor U9122 (N_9122,N_943,N_3846);
nor U9123 (N_9123,N_1774,N_4161);
or U9124 (N_9124,N_4436,N_1772);
or U9125 (N_9125,N_1030,N_3044);
or U9126 (N_9126,N_2211,N_4540);
nor U9127 (N_9127,N_2562,N_64);
nor U9128 (N_9128,N_903,N_3447);
nor U9129 (N_9129,N_3454,N_4089);
and U9130 (N_9130,N_263,N_3153);
nand U9131 (N_9131,N_3404,N_276);
nor U9132 (N_9132,N_47,N_1525);
nor U9133 (N_9133,N_1420,N_1910);
nor U9134 (N_9134,N_2987,N_3431);
nand U9135 (N_9135,N_978,N_3698);
and U9136 (N_9136,N_2671,N_4089);
or U9137 (N_9137,N_4813,N_2426);
nor U9138 (N_9138,N_1593,N_3906);
nand U9139 (N_9139,N_989,N_4646);
or U9140 (N_9140,N_3182,N_249);
nor U9141 (N_9141,N_4800,N_2525);
or U9142 (N_9142,N_2057,N_3439);
nor U9143 (N_9143,N_2452,N_1447);
and U9144 (N_9144,N_2407,N_1086);
nand U9145 (N_9145,N_604,N_4493);
nor U9146 (N_9146,N_2413,N_772);
and U9147 (N_9147,N_2159,N_1821);
nor U9148 (N_9148,N_2436,N_4454);
and U9149 (N_9149,N_1492,N_4385);
and U9150 (N_9150,N_4839,N_1935);
nor U9151 (N_9151,N_4415,N_2184);
nand U9152 (N_9152,N_936,N_875);
and U9153 (N_9153,N_397,N_1109);
or U9154 (N_9154,N_1134,N_1972);
nor U9155 (N_9155,N_1625,N_3796);
and U9156 (N_9156,N_2291,N_2063);
or U9157 (N_9157,N_2630,N_2870);
nor U9158 (N_9158,N_1047,N_4218);
and U9159 (N_9159,N_2173,N_3243);
and U9160 (N_9160,N_508,N_1619);
or U9161 (N_9161,N_4570,N_1656);
nor U9162 (N_9162,N_3496,N_2134);
nand U9163 (N_9163,N_4413,N_2730);
and U9164 (N_9164,N_3054,N_2803);
nand U9165 (N_9165,N_2474,N_2918);
or U9166 (N_9166,N_3323,N_1950);
or U9167 (N_9167,N_4621,N_4728);
nand U9168 (N_9168,N_2966,N_4554);
and U9169 (N_9169,N_2693,N_4127);
and U9170 (N_9170,N_4615,N_1848);
or U9171 (N_9171,N_4008,N_333);
or U9172 (N_9172,N_3940,N_3143);
nand U9173 (N_9173,N_3991,N_482);
nor U9174 (N_9174,N_581,N_3689);
and U9175 (N_9175,N_4650,N_812);
or U9176 (N_9176,N_3468,N_941);
or U9177 (N_9177,N_1861,N_1991);
nor U9178 (N_9178,N_1587,N_4223);
or U9179 (N_9179,N_4979,N_2992);
and U9180 (N_9180,N_4562,N_2339);
xor U9181 (N_9181,N_3939,N_3316);
or U9182 (N_9182,N_2058,N_3336);
and U9183 (N_9183,N_2911,N_1781);
and U9184 (N_9184,N_2608,N_2894);
nor U9185 (N_9185,N_1112,N_4950);
nor U9186 (N_9186,N_3891,N_1521);
and U9187 (N_9187,N_2146,N_1116);
nand U9188 (N_9188,N_1464,N_292);
or U9189 (N_9189,N_1708,N_2705);
nand U9190 (N_9190,N_2671,N_3089);
nor U9191 (N_9191,N_1641,N_4802);
and U9192 (N_9192,N_1256,N_1493);
and U9193 (N_9193,N_4954,N_1303);
nor U9194 (N_9194,N_3302,N_4182);
or U9195 (N_9195,N_2484,N_1021);
nor U9196 (N_9196,N_2136,N_4679);
nand U9197 (N_9197,N_285,N_1433);
or U9198 (N_9198,N_442,N_2957);
or U9199 (N_9199,N_2252,N_3068);
nor U9200 (N_9200,N_3714,N_4569);
and U9201 (N_9201,N_2901,N_4970);
and U9202 (N_9202,N_2628,N_2716);
and U9203 (N_9203,N_338,N_4705);
nor U9204 (N_9204,N_4414,N_3509);
and U9205 (N_9205,N_2468,N_1696);
or U9206 (N_9206,N_3958,N_448);
nand U9207 (N_9207,N_3356,N_2926);
and U9208 (N_9208,N_4870,N_546);
nor U9209 (N_9209,N_2380,N_3265);
nor U9210 (N_9210,N_4977,N_4819);
nand U9211 (N_9211,N_4627,N_274);
or U9212 (N_9212,N_4344,N_376);
nand U9213 (N_9213,N_3777,N_4469);
and U9214 (N_9214,N_3057,N_2260);
nand U9215 (N_9215,N_2245,N_228);
and U9216 (N_9216,N_2185,N_2455);
nor U9217 (N_9217,N_3608,N_1410);
and U9218 (N_9218,N_515,N_4337);
or U9219 (N_9219,N_3674,N_2739);
nor U9220 (N_9220,N_1069,N_3213);
or U9221 (N_9221,N_16,N_1581);
or U9222 (N_9222,N_753,N_204);
or U9223 (N_9223,N_3863,N_1876);
nor U9224 (N_9224,N_3561,N_460);
nand U9225 (N_9225,N_1805,N_3293);
and U9226 (N_9226,N_1430,N_3259);
and U9227 (N_9227,N_2538,N_4726);
or U9228 (N_9228,N_3990,N_4743);
nor U9229 (N_9229,N_737,N_4610);
or U9230 (N_9230,N_4573,N_2949);
and U9231 (N_9231,N_1935,N_3359);
nor U9232 (N_9232,N_1049,N_4642);
nor U9233 (N_9233,N_2166,N_2079);
or U9234 (N_9234,N_874,N_3371);
and U9235 (N_9235,N_418,N_4798);
nand U9236 (N_9236,N_4125,N_4907);
or U9237 (N_9237,N_89,N_4907);
or U9238 (N_9238,N_4998,N_4064);
nand U9239 (N_9239,N_1584,N_4315);
nor U9240 (N_9240,N_4175,N_2690);
and U9241 (N_9241,N_3650,N_1969);
nand U9242 (N_9242,N_3056,N_489);
and U9243 (N_9243,N_3517,N_3055);
nand U9244 (N_9244,N_4374,N_477);
or U9245 (N_9245,N_5,N_1245);
or U9246 (N_9246,N_2392,N_2829);
or U9247 (N_9247,N_2204,N_1106);
nor U9248 (N_9248,N_3864,N_10);
nand U9249 (N_9249,N_1271,N_4631);
nor U9250 (N_9250,N_1050,N_4229);
nor U9251 (N_9251,N_3382,N_2095);
nor U9252 (N_9252,N_2702,N_1032);
or U9253 (N_9253,N_3052,N_3434);
and U9254 (N_9254,N_1454,N_1103);
or U9255 (N_9255,N_4310,N_1468);
nor U9256 (N_9256,N_720,N_4693);
nand U9257 (N_9257,N_516,N_3695);
nor U9258 (N_9258,N_2417,N_1469);
nand U9259 (N_9259,N_4072,N_1837);
and U9260 (N_9260,N_1207,N_2704);
nor U9261 (N_9261,N_2854,N_2239);
or U9262 (N_9262,N_4823,N_2887);
nor U9263 (N_9263,N_4793,N_754);
or U9264 (N_9264,N_4571,N_928);
and U9265 (N_9265,N_2376,N_3819);
or U9266 (N_9266,N_1264,N_4478);
nand U9267 (N_9267,N_4003,N_811);
nor U9268 (N_9268,N_3518,N_1025);
nand U9269 (N_9269,N_4209,N_1516);
and U9270 (N_9270,N_3646,N_1567);
nand U9271 (N_9271,N_1980,N_4663);
and U9272 (N_9272,N_111,N_1999);
or U9273 (N_9273,N_487,N_2131);
and U9274 (N_9274,N_3101,N_2038);
or U9275 (N_9275,N_1660,N_3861);
and U9276 (N_9276,N_1415,N_2758);
and U9277 (N_9277,N_236,N_2463);
and U9278 (N_9278,N_405,N_1972);
or U9279 (N_9279,N_2169,N_3524);
nor U9280 (N_9280,N_851,N_2711);
nor U9281 (N_9281,N_3991,N_2895);
nor U9282 (N_9282,N_3093,N_3859);
nor U9283 (N_9283,N_556,N_4638);
nor U9284 (N_9284,N_1727,N_1196);
nor U9285 (N_9285,N_3947,N_2768);
and U9286 (N_9286,N_4867,N_350);
and U9287 (N_9287,N_487,N_3336);
nand U9288 (N_9288,N_1672,N_4908);
or U9289 (N_9289,N_4415,N_3008);
nand U9290 (N_9290,N_921,N_1257);
nand U9291 (N_9291,N_3557,N_4682);
or U9292 (N_9292,N_4185,N_2404);
or U9293 (N_9293,N_3666,N_4942);
nor U9294 (N_9294,N_4959,N_1305);
and U9295 (N_9295,N_2783,N_824);
nand U9296 (N_9296,N_3347,N_1050);
nor U9297 (N_9297,N_4631,N_2382);
nand U9298 (N_9298,N_4179,N_1050);
xnor U9299 (N_9299,N_3626,N_711);
and U9300 (N_9300,N_403,N_1639);
and U9301 (N_9301,N_1213,N_4549);
or U9302 (N_9302,N_3656,N_2981);
or U9303 (N_9303,N_4412,N_2986);
nand U9304 (N_9304,N_4873,N_1478);
or U9305 (N_9305,N_153,N_2678);
nor U9306 (N_9306,N_464,N_4531);
xor U9307 (N_9307,N_1730,N_4866);
and U9308 (N_9308,N_4656,N_2020);
nor U9309 (N_9309,N_802,N_4937);
and U9310 (N_9310,N_3187,N_2273);
xor U9311 (N_9311,N_213,N_2338);
xnor U9312 (N_9312,N_1797,N_4983);
nand U9313 (N_9313,N_3083,N_2486);
and U9314 (N_9314,N_2481,N_1702);
and U9315 (N_9315,N_1534,N_3831);
or U9316 (N_9316,N_3753,N_1737);
nor U9317 (N_9317,N_2765,N_4171);
and U9318 (N_9318,N_4305,N_3667);
and U9319 (N_9319,N_3761,N_1574);
nor U9320 (N_9320,N_4086,N_703);
nand U9321 (N_9321,N_438,N_2331);
xnor U9322 (N_9322,N_1457,N_2692);
nand U9323 (N_9323,N_2527,N_3759);
or U9324 (N_9324,N_73,N_4921);
or U9325 (N_9325,N_3835,N_868);
nor U9326 (N_9326,N_4903,N_1335);
and U9327 (N_9327,N_611,N_1948);
nand U9328 (N_9328,N_3812,N_3146);
or U9329 (N_9329,N_1238,N_3429);
nor U9330 (N_9330,N_4004,N_4259);
nand U9331 (N_9331,N_1300,N_135);
and U9332 (N_9332,N_2547,N_897);
and U9333 (N_9333,N_3117,N_538);
and U9334 (N_9334,N_2874,N_439);
nand U9335 (N_9335,N_2677,N_3996);
and U9336 (N_9336,N_223,N_3719);
nand U9337 (N_9337,N_3630,N_3373);
nor U9338 (N_9338,N_3513,N_2533);
nand U9339 (N_9339,N_2918,N_1148);
or U9340 (N_9340,N_3131,N_1535);
nor U9341 (N_9341,N_3659,N_2013);
nand U9342 (N_9342,N_246,N_521);
nand U9343 (N_9343,N_1020,N_1106);
and U9344 (N_9344,N_831,N_3131);
or U9345 (N_9345,N_3570,N_2760);
and U9346 (N_9346,N_2886,N_1912);
nand U9347 (N_9347,N_4740,N_2725);
or U9348 (N_9348,N_2823,N_291);
nor U9349 (N_9349,N_4780,N_735);
or U9350 (N_9350,N_1527,N_2196);
and U9351 (N_9351,N_1161,N_1151);
nand U9352 (N_9352,N_4794,N_1297);
nand U9353 (N_9353,N_4465,N_229);
or U9354 (N_9354,N_3621,N_2449);
and U9355 (N_9355,N_2491,N_3901);
and U9356 (N_9356,N_3117,N_4959);
and U9357 (N_9357,N_1024,N_2695);
or U9358 (N_9358,N_1408,N_2670);
nor U9359 (N_9359,N_412,N_754);
and U9360 (N_9360,N_731,N_1961);
nor U9361 (N_9361,N_3232,N_304);
nor U9362 (N_9362,N_664,N_1054);
nor U9363 (N_9363,N_3118,N_3677);
nand U9364 (N_9364,N_1448,N_4770);
nor U9365 (N_9365,N_3402,N_3934);
or U9366 (N_9366,N_4922,N_3708);
nor U9367 (N_9367,N_785,N_3809);
nor U9368 (N_9368,N_3429,N_3956);
and U9369 (N_9369,N_460,N_2456);
nand U9370 (N_9370,N_3613,N_66);
and U9371 (N_9371,N_2885,N_4292);
nor U9372 (N_9372,N_4842,N_4065);
nor U9373 (N_9373,N_2278,N_2202);
and U9374 (N_9374,N_750,N_2803);
or U9375 (N_9375,N_44,N_420);
nor U9376 (N_9376,N_4062,N_4813);
nor U9377 (N_9377,N_1692,N_4899);
nor U9378 (N_9378,N_4053,N_2103);
nand U9379 (N_9379,N_292,N_327);
or U9380 (N_9380,N_2853,N_970);
nand U9381 (N_9381,N_2531,N_3001);
nand U9382 (N_9382,N_3239,N_3271);
and U9383 (N_9383,N_4318,N_135);
and U9384 (N_9384,N_4319,N_343);
and U9385 (N_9385,N_1369,N_22);
or U9386 (N_9386,N_222,N_3366);
nor U9387 (N_9387,N_1906,N_2042);
nand U9388 (N_9388,N_3485,N_2030);
nand U9389 (N_9389,N_1500,N_3152);
or U9390 (N_9390,N_1498,N_854);
or U9391 (N_9391,N_3912,N_795);
nor U9392 (N_9392,N_4172,N_1988);
nor U9393 (N_9393,N_2384,N_2927);
nand U9394 (N_9394,N_43,N_4223);
nand U9395 (N_9395,N_4507,N_3411);
nor U9396 (N_9396,N_2280,N_4702);
nor U9397 (N_9397,N_3025,N_3475);
nand U9398 (N_9398,N_150,N_515);
or U9399 (N_9399,N_1794,N_2931);
nor U9400 (N_9400,N_1451,N_1222);
nor U9401 (N_9401,N_4170,N_4032);
nand U9402 (N_9402,N_2371,N_4134);
nand U9403 (N_9403,N_62,N_3482);
nor U9404 (N_9404,N_4009,N_912);
and U9405 (N_9405,N_2827,N_4367);
nor U9406 (N_9406,N_2477,N_2979);
or U9407 (N_9407,N_2979,N_1336);
and U9408 (N_9408,N_357,N_2465);
nand U9409 (N_9409,N_1305,N_1506);
nor U9410 (N_9410,N_2739,N_4424);
or U9411 (N_9411,N_49,N_4093);
xor U9412 (N_9412,N_4870,N_1272);
nand U9413 (N_9413,N_297,N_4342);
nand U9414 (N_9414,N_2886,N_4892);
nor U9415 (N_9415,N_4615,N_514);
or U9416 (N_9416,N_3808,N_4067);
nand U9417 (N_9417,N_2823,N_1310);
nand U9418 (N_9418,N_2470,N_267);
nor U9419 (N_9419,N_1533,N_1436);
or U9420 (N_9420,N_424,N_2920);
and U9421 (N_9421,N_153,N_1560);
or U9422 (N_9422,N_3730,N_3069);
nand U9423 (N_9423,N_2954,N_3556);
or U9424 (N_9424,N_1435,N_1169);
nand U9425 (N_9425,N_4076,N_1055);
nor U9426 (N_9426,N_4304,N_2012);
nor U9427 (N_9427,N_2570,N_3616);
and U9428 (N_9428,N_671,N_2838);
nand U9429 (N_9429,N_3400,N_1831);
or U9430 (N_9430,N_3396,N_652);
nor U9431 (N_9431,N_4898,N_3974);
or U9432 (N_9432,N_449,N_1776);
or U9433 (N_9433,N_2269,N_1447);
or U9434 (N_9434,N_4662,N_4471);
nor U9435 (N_9435,N_3459,N_1625);
nand U9436 (N_9436,N_3195,N_3635);
and U9437 (N_9437,N_3257,N_797);
and U9438 (N_9438,N_1251,N_1188);
and U9439 (N_9439,N_1510,N_1689);
or U9440 (N_9440,N_4505,N_2558);
or U9441 (N_9441,N_4486,N_3056);
and U9442 (N_9442,N_4436,N_4466);
and U9443 (N_9443,N_3055,N_2924);
xnor U9444 (N_9444,N_4175,N_3975);
nand U9445 (N_9445,N_3305,N_3922);
and U9446 (N_9446,N_1228,N_4455);
and U9447 (N_9447,N_478,N_403);
nand U9448 (N_9448,N_1750,N_781);
nor U9449 (N_9449,N_1201,N_3455);
and U9450 (N_9450,N_799,N_1459);
or U9451 (N_9451,N_1557,N_4384);
and U9452 (N_9452,N_4627,N_888);
nand U9453 (N_9453,N_3898,N_4388);
nor U9454 (N_9454,N_1344,N_4289);
nor U9455 (N_9455,N_341,N_1709);
or U9456 (N_9456,N_3032,N_3423);
nor U9457 (N_9457,N_3006,N_3609);
and U9458 (N_9458,N_3336,N_1242);
and U9459 (N_9459,N_1779,N_3776);
xor U9460 (N_9460,N_520,N_4009);
nand U9461 (N_9461,N_3724,N_672);
or U9462 (N_9462,N_1113,N_2359);
nor U9463 (N_9463,N_680,N_3418);
or U9464 (N_9464,N_1541,N_4647);
and U9465 (N_9465,N_2835,N_558);
nand U9466 (N_9466,N_1744,N_391);
nor U9467 (N_9467,N_3352,N_2019);
and U9468 (N_9468,N_893,N_804);
or U9469 (N_9469,N_749,N_122);
nor U9470 (N_9470,N_1677,N_4289);
or U9471 (N_9471,N_4696,N_1265);
and U9472 (N_9472,N_4578,N_4345);
nand U9473 (N_9473,N_1491,N_3107);
nand U9474 (N_9474,N_2664,N_3820);
nand U9475 (N_9475,N_834,N_248);
or U9476 (N_9476,N_1322,N_4095);
and U9477 (N_9477,N_1686,N_4367);
and U9478 (N_9478,N_2919,N_4556);
and U9479 (N_9479,N_3359,N_4203);
nand U9480 (N_9480,N_2828,N_875);
and U9481 (N_9481,N_2365,N_3347);
nor U9482 (N_9482,N_2093,N_1893);
or U9483 (N_9483,N_2181,N_1231);
nand U9484 (N_9484,N_1196,N_151);
and U9485 (N_9485,N_4444,N_4739);
and U9486 (N_9486,N_4046,N_903);
or U9487 (N_9487,N_4703,N_2862);
nand U9488 (N_9488,N_3702,N_315);
or U9489 (N_9489,N_1991,N_919);
nand U9490 (N_9490,N_202,N_4210);
and U9491 (N_9491,N_1207,N_1817);
nor U9492 (N_9492,N_4786,N_403);
and U9493 (N_9493,N_2126,N_3133);
nor U9494 (N_9494,N_4945,N_436);
nand U9495 (N_9495,N_2476,N_1573);
and U9496 (N_9496,N_1634,N_3594);
nand U9497 (N_9497,N_2985,N_685);
nor U9498 (N_9498,N_2046,N_3225);
nand U9499 (N_9499,N_1957,N_4202);
nand U9500 (N_9500,N_4580,N_3807);
nand U9501 (N_9501,N_455,N_4022);
nor U9502 (N_9502,N_891,N_4763);
or U9503 (N_9503,N_4949,N_3855);
nor U9504 (N_9504,N_3568,N_2115);
or U9505 (N_9505,N_2689,N_3253);
or U9506 (N_9506,N_436,N_290);
and U9507 (N_9507,N_1453,N_3756);
or U9508 (N_9508,N_1728,N_2818);
nor U9509 (N_9509,N_3556,N_3143);
or U9510 (N_9510,N_577,N_1910);
and U9511 (N_9511,N_249,N_4052);
or U9512 (N_9512,N_1422,N_1778);
nand U9513 (N_9513,N_1149,N_3240);
nor U9514 (N_9514,N_4080,N_4540);
nor U9515 (N_9515,N_3709,N_3796);
nor U9516 (N_9516,N_3553,N_4387);
nor U9517 (N_9517,N_1345,N_4251);
nor U9518 (N_9518,N_1683,N_2858);
and U9519 (N_9519,N_3260,N_2968);
or U9520 (N_9520,N_3710,N_2868);
nor U9521 (N_9521,N_3500,N_4285);
nand U9522 (N_9522,N_552,N_1456);
nand U9523 (N_9523,N_2690,N_4575);
nand U9524 (N_9524,N_432,N_2716);
and U9525 (N_9525,N_4070,N_1355);
nor U9526 (N_9526,N_134,N_2538);
nor U9527 (N_9527,N_1808,N_4673);
or U9528 (N_9528,N_3849,N_2622);
and U9529 (N_9529,N_1742,N_4822);
nor U9530 (N_9530,N_3578,N_1424);
and U9531 (N_9531,N_3245,N_2776);
or U9532 (N_9532,N_4740,N_801);
nand U9533 (N_9533,N_2231,N_1978);
nand U9534 (N_9534,N_4320,N_3306);
nand U9535 (N_9535,N_1575,N_449);
nand U9536 (N_9536,N_4991,N_1737);
nor U9537 (N_9537,N_3252,N_4819);
and U9538 (N_9538,N_1391,N_1656);
or U9539 (N_9539,N_193,N_2134);
nor U9540 (N_9540,N_1704,N_3403);
nand U9541 (N_9541,N_4052,N_3015);
nor U9542 (N_9542,N_2139,N_9);
nor U9543 (N_9543,N_296,N_3452);
or U9544 (N_9544,N_3730,N_944);
or U9545 (N_9545,N_1523,N_4084);
or U9546 (N_9546,N_3033,N_4931);
or U9547 (N_9547,N_3519,N_4233);
nand U9548 (N_9548,N_2332,N_2219);
and U9549 (N_9549,N_415,N_2185);
and U9550 (N_9550,N_3476,N_223);
and U9551 (N_9551,N_4858,N_2496);
nor U9552 (N_9552,N_2472,N_2789);
and U9553 (N_9553,N_2213,N_2086);
and U9554 (N_9554,N_24,N_3630);
nor U9555 (N_9555,N_2846,N_420);
or U9556 (N_9556,N_4759,N_2454);
or U9557 (N_9557,N_4122,N_441);
or U9558 (N_9558,N_2167,N_123);
and U9559 (N_9559,N_3793,N_4282);
or U9560 (N_9560,N_3498,N_3195);
or U9561 (N_9561,N_329,N_4274);
nor U9562 (N_9562,N_1761,N_3134);
nand U9563 (N_9563,N_1064,N_3539);
nand U9564 (N_9564,N_1185,N_244);
and U9565 (N_9565,N_1508,N_1207);
nor U9566 (N_9566,N_710,N_4168);
nand U9567 (N_9567,N_406,N_214);
nand U9568 (N_9568,N_4307,N_3089);
and U9569 (N_9569,N_45,N_3634);
or U9570 (N_9570,N_3745,N_902);
and U9571 (N_9571,N_613,N_2753);
and U9572 (N_9572,N_1129,N_66);
nand U9573 (N_9573,N_4665,N_3995);
nor U9574 (N_9574,N_1708,N_4386);
and U9575 (N_9575,N_4574,N_3641);
and U9576 (N_9576,N_1769,N_3422);
nor U9577 (N_9577,N_1054,N_3518);
or U9578 (N_9578,N_1834,N_4549);
nor U9579 (N_9579,N_2103,N_2948);
or U9580 (N_9580,N_3301,N_2977);
nand U9581 (N_9581,N_769,N_1858);
or U9582 (N_9582,N_4282,N_64);
nor U9583 (N_9583,N_2951,N_1199);
nand U9584 (N_9584,N_2046,N_3558);
and U9585 (N_9585,N_2996,N_3468);
xor U9586 (N_9586,N_1940,N_3050);
or U9587 (N_9587,N_4374,N_443);
or U9588 (N_9588,N_4024,N_4860);
or U9589 (N_9589,N_3908,N_756);
or U9590 (N_9590,N_4796,N_2997);
nor U9591 (N_9591,N_2121,N_1609);
and U9592 (N_9592,N_1679,N_2456);
nand U9593 (N_9593,N_2165,N_4261);
nand U9594 (N_9594,N_4977,N_499);
and U9595 (N_9595,N_2165,N_1349);
and U9596 (N_9596,N_3882,N_3382);
and U9597 (N_9597,N_1999,N_2709);
and U9598 (N_9598,N_499,N_2383);
or U9599 (N_9599,N_1657,N_4511);
and U9600 (N_9600,N_4449,N_4986);
nor U9601 (N_9601,N_1537,N_2425);
nor U9602 (N_9602,N_4808,N_1570);
nand U9603 (N_9603,N_1075,N_3914);
or U9604 (N_9604,N_3862,N_4819);
nor U9605 (N_9605,N_3881,N_2601);
nor U9606 (N_9606,N_3159,N_4865);
or U9607 (N_9607,N_4391,N_551);
nand U9608 (N_9608,N_1970,N_1250);
nand U9609 (N_9609,N_3403,N_3497);
and U9610 (N_9610,N_2455,N_1233);
and U9611 (N_9611,N_3181,N_2075);
or U9612 (N_9612,N_1685,N_34);
nor U9613 (N_9613,N_2919,N_4349);
or U9614 (N_9614,N_2776,N_3149);
nor U9615 (N_9615,N_4087,N_1580);
and U9616 (N_9616,N_4682,N_1074);
nor U9617 (N_9617,N_1880,N_2565);
nor U9618 (N_9618,N_4330,N_4754);
or U9619 (N_9619,N_4999,N_2534);
nand U9620 (N_9620,N_1456,N_4217);
nor U9621 (N_9621,N_3001,N_4296);
or U9622 (N_9622,N_3953,N_3304);
nor U9623 (N_9623,N_880,N_4803);
or U9624 (N_9624,N_3430,N_3067);
or U9625 (N_9625,N_3691,N_3758);
and U9626 (N_9626,N_4560,N_1422);
nor U9627 (N_9627,N_3574,N_3167);
or U9628 (N_9628,N_332,N_1436);
nor U9629 (N_9629,N_1970,N_1624);
or U9630 (N_9630,N_3037,N_4081);
or U9631 (N_9631,N_1097,N_2628);
nor U9632 (N_9632,N_75,N_3147);
or U9633 (N_9633,N_1040,N_1849);
or U9634 (N_9634,N_2275,N_3775);
nand U9635 (N_9635,N_1412,N_1642);
xnor U9636 (N_9636,N_4078,N_3412);
and U9637 (N_9637,N_2055,N_2127);
nor U9638 (N_9638,N_4698,N_4330);
nor U9639 (N_9639,N_1710,N_4678);
nand U9640 (N_9640,N_2741,N_3624);
or U9641 (N_9641,N_2879,N_709);
nand U9642 (N_9642,N_4364,N_1992);
xor U9643 (N_9643,N_3862,N_3512);
or U9644 (N_9644,N_937,N_84);
and U9645 (N_9645,N_4617,N_1039);
nand U9646 (N_9646,N_1715,N_3964);
and U9647 (N_9647,N_369,N_2345);
nor U9648 (N_9648,N_4313,N_2073);
nor U9649 (N_9649,N_2899,N_3758);
or U9650 (N_9650,N_1268,N_844);
nor U9651 (N_9651,N_3870,N_3325);
and U9652 (N_9652,N_2306,N_1255);
nand U9653 (N_9653,N_1834,N_3917);
and U9654 (N_9654,N_138,N_2032);
nor U9655 (N_9655,N_385,N_3644);
nor U9656 (N_9656,N_4672,N_4597);
nand U9657 (N_9657,N_1166,N_709);
or U9658 (N_9658,N_575,N_1043);
nand U9659 (N_9659,N_1984,N_3332);
nand U9660 (N_9660,N_2470,N_2972);
and U9661 (N_9661,N_119,N_2917);
nor U9662 (N_9662,N_1476,N_3265);
and U9663 (N_9663,N_661,N_1161);
nand U9664 (N_9664,N_187,N_3061);
or U9665 (N_9665,N_911,N_1988);
or U9666 (N_9666,N_4712,N_1110);
or U9667 (N_9667,N_327,N_2011);
nand U9668 (N_9668,N_4246,N_4394);
nand U9669 (N_9669,N_3107,N_1668);
nand U9670 (N_9670,N_3282,N_32);
or U9671 (N_9671,N_2588,N_1365);
and U9672 (N_9672,N_1591,N_1702);
or U9673 (N_9673,N_1821,N_2484);
nor U9674 (N_9674,N_875,N_4772);
or U9675 (N_9675,N_2663,N_159);
nand U9676 (N_9676,N_3978,N_3394);
nor U9677 (N_9677,N_3099,N_4494);
nor U9678 (N_9678,N_315,N_2498);
nor U9679 (N_9679,N_1526,N_3466);
nor U9680 (N_9680,N_914,N_1379);
nor U9681 (N_9681,N_608,N_4022);
or U9682 (N_9682,N_3403,N_1470);
or U9683 (N_9683,N_2339,N_2677);
nand U9684 (N_9684,N_105,N_3487);
nand U9685 (N_9685,N_219,N_4106);
or U9686 (N_9686,N_2562,N_4577);
or U9687 (N_9687,N_3565,N_2225);
nor U9688 (N_9688,N_1466,N_1147);
nand U9689 (N_9689,N_414,N_521);
nand U9690 (N_9690,N_29,N_2306);
nor U9691 (N_9691,N_2601,N_286);
and U9692 (N_9692,N_366,N_3372);
nor U9693 (N_9693,N_329,N_1849);
and U9694 (N_9694,N_2067,N_1931);
nand U9695 (N_9695,N_1090,N_1376);
nand U9696 (N_9696,N_2930,N_3091);
nand U9697 (N_9697,N_4534,N_3095);
and U9698 (N_9698,N_1284,N_4877);
or U9699 (N_9699,N_2769,N_1890);
or U9700 (N_9700,N_1293,N_4153);
nand U9701 (N_9701,N_4744,N_465);
or U9702 (N_9702,N_2388,N_2511);
nand U9703 (N_9703,N_4333,N_2244);
nand U9704 (N_9704,N_2940,N_4347);
nor U9705 (N_9705,N_3247,N_3490);
or U9706 (N_9706,N_4553,N_945);
nor U9707 (N_9707,N_2344,N_3156);
nand U9708 (N_9708,N_1809,N_1525);
nand U9709 (N_9709,N_2912,N_1227);
nand U9710 (N_9710,N_1509,N_2912);
nand U9711 (N_9711,N_1597,N_4832);
nand U9712 (N_9712,N_2416,N_1359);
nand U9713 (N_9713,N_4304,N_1108);
nand U9714 (N_9714,N_4545,N_2369);
or U9715 (N_9715,N_1650,N_1902);
nand U9716 (N_9716,N_2287,N_2117);
nor U9717 (N_9717,N_3444,N_3490);
or U9718 (N_9718,N_306,N_719);
or U9719 (N_9719,N_1790,N_337);
and U9720 (N_9720,N_3725,N_2736);
nor U9721 (N_9721,N_2688,N_1279);
and U9722 (N_9722,N_595,N_818);
nand U9723 (N_9723,N_569,N_2963);
nor U9724 (N_9724,N_4012,N_4603);
or U9725 (N_9725,N_1486,N_2148);
and U9726 (N_9726,N_4677,N_804);
nor U9727 (N_9727,N_1875,N_976);
and U9728 (N_9728,N_4262,N_3285);
nand U9729 (N_9729,N_1804,N_4285);
nor U9730 (N_9730,N_1118,N_4327);
xnor U9731 (N_9731,N_1896,N_1108);
and U9732 (N_9732,N_250,N_3703);
and U9733 (N_9733,N_4909,N_1718);
nand U9734 (N_9734,N_2724,N_1690);
and U9735 (N_9735,N_2415,N_3478);
and U9736 (N_9736,N_919,N_1891);
nand U9737 (N_9737,N_2090,N_843);
nor U9738 (N_9738,N_4582,N_2098);
and U9739 (N_9739,N_3327,N_1489);
nor U9740 (N_9740,N_492,N_4009);
nor U9741 (N_9741,N_2866,N_4983);
xnor U9742 (N_9742,N_2098,N_2412);
nand U9743 (N_9743,N_4188,N_325);
and U9744 (N_9744,N_2131,N_327);
nand U9745 (N_9745,N_969,N_794);
nand U9746 (N_9746,N_788,N_2689);
or U9747 (N_9747,N_4525,N_2279);
nand U9748 (N_9748,N_4077,N_3314);
nor U9749 (N_9749,N_2222,N_2785);
nor U9750 (N_9750,N_3985,N_2060);
nand U9751 (N_9751,N_3999,N_1487);
nor U9752 (N_9752,N_3954,N_3283);
nand U9753 (N_9753,N_4285,N_914);
or U9754 (N_9754,N_406,N_2893);
nor U9755 (N_9755,N_1627,N_442);
nand U9756 (N_9756,N_1689,N_4435);
nand U9757 (N_9757,N_4464,N_3461);
nand U9758 (N_9758,N_1415,N_3229);
nor U9759 (N_9759,N_4566,N_1483);
and U9760 (N_9760,N_2457,N_4627);
nand U9761 (N_9761,N_1708,N_1219);
nor U9762 (N_9762,N_4338,N_2415);
nor U9763 (N_9763,N_4098,N_4497);
or U9764 (N_9764,N_2803,N_844);
nor U9765 (N_9765,N_4020,N_3045);
or U9766 (N_9766,N_4512,N_1951);
nand U9767 (N_9767,N_4436,N_1064);
nand U9768 (N_9768,N_1484,N_3140);
nor U9769 (N_9769,N_2036,N_4792);
and U9770 (N_9770,N_1587,N_2530);
nor U9771 (N_9771,N_1567,N_1762);
nand U9772 (N_9772,N_569,N_2022);
nor U9773 (N_9773,N_4760,N_4190);
nand U9774 (N_9774,N_1957,N_1904);
or U9775 (N_9775,N_2031,N_2672);
nor U9776 (N_9776,N_841,N_1171);
nand U9777 (N_9777,N_2910,N_4719);
nor U9778 (N_9778,N_860,N_1864);
nand U9779 (N_9779,N_3493,N_2892);
nor U9780 (N_9780,N_4258,N_1763);
or U9781 (N_9781,N_3802,N_251);
or U9782 (N_9782,N_4121,N_4428);
or U9783 (N_9783,N_3877,N_1988);
and U9784 (N_9784,N_2820,N_3132);
nand U9785 (N_9785,N_4726,N_2971);
and U9786 (N_9786,N_3528,N_357);
nor U9787 (N_9787,N_3248,N_3336);
nand U9788 (N_9788,N_4432,N_655);
nand U9789 (N_9789,N_1763,N_1653);
nor U9790 (N_9790,N_3363,N_477);
nand U9791 (N_9791,N_887,N_3454);
nand U9792 (N_9792,N_4922,N_4133);
or U9793 (N_9793,N_538,N_2390);
or U9794 (N_9794,N_1611,N_3725);
nor U9795 (N_9795,N_278,N_1490);
and U9796 (N_9796,N_4708,N_4843);
nand U9797 (N_9797,N_1878,N_2532);
or U9798 (N_9798,N_1220,N_4154);
or U9799 (N_9799,N_55,N_4494);
nand U9800 (N_9800,N_612,N_2070);
nand U9801 (N_9801,N_4065,N_1885);
and U9802 (N_9802,N_4921,N_152);
nor U9803 (N_9803,N_2859,N_3547);
nand U9804 (N_9804,N_3103,N_2624);
xor U9805 (N_9805,N_1869,N_4843);
nand U9806 (N_9806,N_2513,N_4582);
or U9807 (N_9807,N_3445,N_1651);
nor U9808 (N_9808,N_4912,N_2134);
nand U9809 (N_9809,N_4859,N_3056);
nor U9810 (N_9810,N_740,N_619);
nor U9811 (N_9811,N_871,N_1482);
and U9812 (N_9812,N_1709,N_2882);
nand U9813 (N_9813,N_1769,N_4066);
nor U9814 (N_9814,N_1219,N_338);
and U9815 (N_9815,N_3256,N_987);
and U9816 (N_9816,N_4886,N_3071);
or U9817 (N_9817,N_2660,N_1696);
nand U9818 (N_9818,N_3203,N_2216);
nand U9819 (N_9819,N_3224,N_1691);
and U9820 (N_9820,N_4850,N_4529);
nand U9821 (N_9821,N_4173,N_1065);
and U9822 (N_9822,N_179,N_309);
and U9823 (N_9823,N_2512,N_2520);
or U9824 (N_9824,N_771,N_4394);
nand U9825 (N_9825,N_4520,N_2978);
and U9826 (N_9826,N_2164,N_4975);
nor U9827 (N_9827,N_4455,N_4071);
nor U9828 (N_9828,N_2214,N_929);
and U9829 (N_9829,N_447,N_775);
or U9830 (N_9830,N_1748,N_4977);
nor U9831 (N_9831,N_717,N_2627);
nor U9832 (N_9832,N_3305,N_1196);
nor U9833 (N_9833,N_3784,N_4962);
and U9834 (N_9834,N_4818,N_1319);
or U9835 (N_9835,N_678,N_4525);
nor U9836 (N_9836,N_1056,N_4430);
nand U9837 (N_9837,N_2191,N_1000);
nand U9838 (N_9838,N_2389,N_1354);
nor U9839 (N_9839,N_860,N_2483);
and U9840 (N_9840,N_3101,N_1934);
and U9841 (N_9841,N_4879,N_3886);
nor U9842 (N_9842,N_765,N_2149);
and U9843 (N_9843,N_3234,N_3203);
and U9844 (N_9844,N_2989,N_324);
nand U9845 (N_9845,N_1298,N_4787);
and U9846 (N_9846,N_1866,N_2784);
nand U9847 (N_9847,N_3813,N_4204);
and U9848 (N_9848,N_2624,N_4025);
or U9849 (N_9849,N_1936,N_3290);
nor U9850 (N_9850,N_1501,N_2435);
and U9851 (N_9851,N_1412,N_738);
nor U9852 (N_9852,N_3514,N_3691);
nand U9853 (N_9853,N_352,N_938);
nand U9854 (N_9854,N_727,N_4566);
xnor U9855 (N_9855,N_4758,N_4026);
nor U9856 (N_9856,N_621,N_1500);
or U9857 (N_9857,N_4055,N_4368);
nor U9858 (N_9858,N_1414,N_546);
and U9859 (N_9859,N_3985,N_4463);
or U9860 (N_9860,N_3479,N_3141);
and U9861 (N_9861,N_1362,N_2182);
nand U9862 (N_9862,N_4654,N_4841);
or U9863 (N_9863,N_4400,N_885);
or U9864 (N_9864,N_4480,N_4054);
and U9865 (N_9865,N_2748,N_2101);
and U9866 (N_9866,N_3113,N_2105);
or U9867 (N_9867,N_3573,N_178);
nand U9868 (N_9868,N_1082,N_2917);
nand U9869 (N_9869,N_627,N_2694);
nor U9870 (N_9870,N_2371,N_2803);
nor U9871 (N_9871,N_4152,N_3672);
nand U9872 (N_9872,N_866,N_4140);
and U9873 (N_9873,N_2938,N_17);
nand U9874 (N_9874,N_3343,N_3420);
nor U9875 (N_9875,N_1095,N_3988);
nor U9876 (N_9876,N_3774,N_4151);
nand U9877 (N_9877,N_3772,N_1471);
and U9878 (N_9878,N_1931,N_2454);
nand U9879 (N_9879,N_232,N_344);
nand U9880 (N_9880,N_979,N_1311);
or U9881 (N_9881,N_2728,N_4389);
and U9882 (N_9882,N_4270,N_4486);
nor U9883 (N_9883,N_2993,N_1753);
or U9884 (N_9884,N_4727,N_4855);
or U9885 (N_9885,N_391,N_2408);
and U9886 (N_9886,N_4115,N_3897);
nor U9887 (N_9887,N_2625,N_3527);
nand U9888 (N_9888,N_4244,N_844);
nand U9889 (N_9889,N_2218,N_15);
nand U9890 (N_9890,N_3846,N_1492);
or U9891 (N_9891,N_2691,N_1559);
xnor U9892 (N_9892,N_1142,N_4703);
nand U9893 (N_9893,N_102,N_845);
nor U9894 (N_9894,N_2320,N_2551);
nand U9895 (N_9895,N_1493,N_4782);
nand U9896 (N_9896,N_2840,N_888);
and U9897 (N_9897,N_192,N_4275);
or U9898 (N_9898,N_1933,N_1464);
and U9899 (N_9899,N_2794,N_1299);
nand U9900 (N_9900,N_1087,N_3341);
and U9901 (N_9901,N_143,N_4942);
nor U9902 (N_9902,N_1615,N_2687);
nand U9903 (N_9903,N_1270,N_570);
or U9904 (N_9904,N_43,N_2933);
nand U9905 (N_9905,N_3854,N_1915);
nand U9906 (N_9906,N_555,N_330);
nand U9907 (N_9907,N_2089,N_2351);
and U9908 (N_9908,N_583,N_3400);
nor U9909 (N_9909,N_2182,N_2319);
and U9910 (N_9910,N_4556,N_2509);
or U9911 (N_9911,N_2161,N_965);
nand U9912 (N_9912,N_747,N_722);
nor U9913 (N_9913,N_2903,N_508);
nor U9914 (N_9914,N_2783,N_1392);
nor U9915 (N_9915,N_2784,N_4148);
nor U9916 (N_9916,N_443,N_1675);
and U9917 (N_9917,N_1024,N_4989);
xnor U9918 (N_9918,N_2339,N_3066);
nand U9919 (N_9919,N_1339,N_1109);
nand U9920 (N_9920,N_296,N_2437);
nor U9921 (N_9921,N_2454,N_1830);
or U9922 (N_9922,N_3884,N_4789);
nand U9923 (N_9923,N_2382,N_1019);
nand U9924 (N_9924,N_4626,N_1661);
xor U9925 (N_9925,N_571,N_519);
or U9926 (N_9926,N_1839,N_337);
nand U9927 (N_9927,N_4672,N_4001);
and U9928 (N_9928,N_1122,N_2396);
nand U9929 (N_9929,N_3232,N_1392);
nor U9930 (N_9930,N_3568,N_4725);
nor U9931 (N_9931,N_2582,N_4325);
and U9932 (N_9932,N_2408,N_4300);
nor U9933 (N_9933,N_2648,N_645);
nor U9934 (N_9934,N_407,N_2201);
nand U9935 (N_9935,N_4335,N_109);
or U9936 (N_9936,N_1485,N_4934);
nor U9937 (N_9937,N_405,N_349);
nor U9938 (N_9938,N_1778,N_3050);
or U9939 (N_9939,N_2751,N_46);
nand U9940 (N_9940,N_3299,N_1963);
nor U9941 (N_9941,N_3532,N_4292);
and U9942 (N_9942,N_1364,N_101);
nand U9943 (N_9943,N_1167,N_4993);
and U9944 (N_9944,N_4668,N_4153);
nor U9945 (N_9945,N_3855,N_1749);
nand U9946 (N_9946,N_740,N_4375);
nand U9947 (N_9947,N_4720,N_3362);
nor U9948 (N_9948,N_2312,N_841);
or U9949 (N_9949,N_4681,N_1751);
and U9950 (N_9950,N_303,N_496);
nand U9951 (N_9951,N_2440,N_280);
and U9952 (N_9952,N_1368,N_3694);
or U9953 (N_9953,N_2873,N_1307);
and U9954 (N_9954,N_4128,N_4593);
nor U9955 (N_9955,N_1221,N_4595);
or U9956 (N_9956,N_2926,N_1170);
nand U9957 (N_9957,N_3435,N_4816);
or U9958 (N_9958,N_4237,N_3599);
or U9959 (N_9959,N_3783,N_150);
xnor U9960 (N_9960,N_784,N_1939);
nand U9961 (N_9961,N_1708,N_3755);
or U9962 (N_9962,N_4566,N_22);
nand U9963 (N_9963,N_4186,N_4982);
and U9964 (N_9964,N_1691,N_2672);
xnor U9965 (N_9965,N_2957,N_415);
or U9966 (N_9966,N_4923,N_4731);
and U9967 (N_9967,N_3407,N_948);
nand U9968 (N_9968,N_1792,N_911);
or U9969 (N_9969,N_4732,N_4318);
and U9970 (N_9970,N_4551,N_4453);
and U9971 (N_9971,N_2883,N_3658);
and U9972 (N_9972,N_1381,N_2705);
or U9973 (N_9973,N_752,N_1510);
nor U9974 (N_9974,N_1087,N_1505);
and U9975 (N_9975,N_61,N_738);
nor U9976 (N_9976,N_586,N_249);
nor U9977 (N_9977,N_3754,N_3497);
nor U9978 (N_9978,N_972,N_4121);
or U9979 (N_9979,N_3182,N_2373);
and U9980 (N_9980,N_1129,N_2033);
nand U9981 (N_9981,N_2114,N_2733);
nor U9982 (N_9982,N_3170,N_277);
nor U9983 (N_9983,N_1628,N_4210);
and U9984 (N_9984,N_3704,N_1947);
nand U9985 (N_9985,N_1537,N_4493);
nor U9986 (N_9986,N_659,N_3787);
nand U9987 (N_9987,N_2374,N_809);
and U9988 (N_9988,N_3568,N_647);
or U9989 (N_9989,N_1438,N_4353);
or U9990 (N_9990,N_907,N_3250);
or U9991 (N_9991,N_3687,N_2526);
or U9992 (N_9992,N_2192,N_2661);
nand U9993 (N_9993,N_376,N_4442);
nand U9994 (N_9994,N_887,N_191);
nor U9995 (N_9995,N_801,N_943);
nand U9996 (N_9996,N_3855,N_387);
nor U9997 (N_9997,N_4144,N_3041);
nor U9998 (N_9998,N_269,N_235);
and U9999 (N_9999,N_2297,N_1192);
or UO_0 (O_0,N_9565,N_8277);
or UO_1 (O_1,N_6497,N_7780);
or UO_2 (O_2,N_9501,N_7445);
nor UO_3 (O_3,N_8702,N_9653);
nor UO_4 (O_4,N_7789,N_8016);
or UO_5 (O_5,N_7661,N_8467);
nor UO_6 (O_6,N_7768,N_9035);
nand UO_7 (O_7,N_8325,N_6265);
nor UO_8 (O_8,N_6973,N_9526);
nand UO_9 (O_9,N_6041,N_9231);
and UO_10 (O_10,N_6353,N_5579);
nand UO_11 (O_11,N_5826,N_6929);
nor UO_12 (O_12,N_6256,N_5555);
nand UO_13 (O_13,N_6090,N_7138);
and UO_14 (O_14,N_7418,N_7172);
nand UO_15 (O_15,N_5084,N_9885);
nor UO_16 (O_16,N_6570,N_7765);
nor UO_17 (O_17,N_6168,N_8351);
or UO_18 (O_18,N_8926,N_7130);
nor UO_19 (O_19,N_8808,N_7817);
nor UO_20 (O_20,N_5483,N_5576);
or UO_21 (O_21,N_8726,N_9728);
nor UO_22 (O_22,N_6761,N_6083);
or UO_23 (O_23,N_7776,N_5527);
or UO_24 (O_24,N_9754,N_6930);
and UO_25 (O_25,N_6775,N_9650);
nor UO_26 (O_26,N_9743,N_8104);
nor UO_27 (O_27,N_6597,N_9620);
nor UO_28 (O_28,N_8990,N_6658);
and UO_29 (O_29,N_7305,N_6916);
and UO_30 (O_30,N_5776,N_6229);
or UO_31 (O_31,N_5886,N_9398);
nand UO_32 (O_32,N_9084,N_7819);
and UO_33 (O_33,N_5662,N_8120);
nand UO_34 (O_34,N_6510,N_5691);
nor UO_35 (O_35,N_6261,N_9202);
nor UO_36 (O_36,N_9114,N_7358);
nand UO_37 (O_37,N_7647,N_5849);
or UO_38 (O_38,N_8634,N_6622);
nor UO_39 (O_39,N_8308,N_8572);
nor UO_40 (O_40,N_8844,N_5594);
nor UO_41 (O_41,N_7204,N_9110);
nand UO_42 (O_42,N_7694,N_5733);
or UO_43 (O_43,N_7845,N_7983);
nand UO_44 (O_44,N_6648,N_8998);
or UO_45 (O_45,N_5689,N_9474);
nand UO_46 (O_46,N_5957,N_5945);
nand UO_47 (O_47,N_8665,N_6184);
or UO_48 (O_48,N_7436,N_6028);
and UO_49 (O_49,N_7899,N_9380);
nand UO_50 (O_50,N_6464,N_6027);
and UO_51 (O_51,N_6405,N_7485);
nor UO_52 (O_52,N_6402,N_6558);
nor UO_53 (O_53,N_9985,N_9814);
or UO_54 (O_54,N_9490,N_9131);
nor UO_55 (O_55,N_7898,N_7581);
and UO_56 (O_56,N_9966,N_6904);
nand UO_57 (O_57,N_7792,N_6840);
and UO_58 (O_58,N_7523,N_8802);
and UO_59 (O_59,N_6102,N_5181);
nand UO_60 (O_60,N_5520,N_6845);
or UO_61 (O_61,N_5348,N_7035);
nor UO_62 (O_62,N_8312,N_7246);
nand UO_63 (O_63,N_7334,N_5684);
and UO_64 (O_64,N_7011,N_9255);
or UO_65 (O_65,N_8704,N_8919);
and UO_66 (O_66,N_5029,N_5008);
nand UO_67 (O_67,N_7945,N_6644);
nand UO_68 (O_68,N_5033,N_6077);
nand UO_69 (O_69,N_9249,N_8574);
nand UO_70 (O_70,N_6128,N_8469);
or UO_71 (O_71,N_5434,N_6447);
or UO_72 (O_72,N_6213,N_6018);
or UO_73 (O_73,N_9784,N_7411);
nand UO_74 (O_74,N_5857,N_7262);
or UO_75 (O_75,N_9841,N_6457);
and UO_76 (O_76,N_7796,N_7573);
or UO_77 (O_77,N_6186,N_6824);
and UO_78 (O_78,N_6959,N_8411);
and UO_79 (O_79,N_9211,N_6312);
or UO_80 (O_80,N_9349,N_6867);
or UO_81 (O_81,N_9121,N_9044);
and UO_82 (O_82,N_8701,N_7300);
and UO_83 (O_83,N_8564,N_5156);
and UO_84 (O_84,N_8507,N_8440);
nand UO_85 (O_85,N_5306,N_8811);
and UO_86 (O_86,N_5672,N_7926);
and UO_87 (O_87,N_9769,N_5472);
or UO_88 (O_88,N_9606,N_5071);
or UO_89 (O_89,N_6626,N_7931);
nand UO_90 (O_90,N_7558,N_6881);
and UO_91 (O_91,N_8715,N_8412);
nor UO_92 (O_92,N_9629,N_5814);
nor UO_93 (O_93,N_7306,N_8892);
nand UO_94 (O_94,N_7493,N_8528);
or UO_95 (O_95,N_8995,N_7354);
nor UO_96 (O_96,N_9953,N_5296);
nor UO_97 (O_97,N_6238,N_5940);
and UO_98 (O_98,N_9543,N_8331);
and UO_99 (O_99,N_8938,N_7616);
or UO_100 (O_100,N_7308,N_8751);
or UO_101 (O_101,N_7872,N_8731);
and UO_102 (O_102,N_5275,N_5879);
or UO_103 (O_103,N_5560,N_9329);
nor UO_104 (O_104,N_7930,N_6907);
nand UO_105 (O_105,N_6065,N_6552);
and UO_106 (O_106,N_9920,N_5778);
or UO_107 (O_107,N_9333,N_8551);
nand UO_108 (O_108,N_9549,N_7302);
nor UO_109 (O_109,N_5611,N_6106);
and UO_110 (O_110,N_6815,N_5028);
and UO_111 (O_111,N_6778,N_6208);
xnor UO_112 (O_112,N_8864,N_7392);
or UO_113 (O_113,N_6308,N_7492);
or UO_114 (O_114,N_9089,N_6234);
or UO_115 (O_115,N_6026,N_5507);
or UO_116 (O_116,N_9248,N_7987);
nand UO_117 (O_117,N_7507,N_9118);
and UO_118 (O_118,N_7446,N_8536);
and UO_119 (O_119,N_5229,N_7638);
and UO_120 (O_120,N_9709,N_7054);
or UO_121 (O_121,N_7218,N_9811);
and UO_122 (O_122,N_5377,N_8039);
nor UO_123 (O_123,N_9945,N_5294);
nand UO_124 (O_124,N_5860,N_7841);
nand UO_125 (O_125,N_8154,N_8557);
nand UO_126 (O_126,N_7294,N_6888);
or UO_127 (O_127,N_8216,N_7038);
nand UO_128 (O_128,N_7729,N_5011);
xor UO_129 (O_129,N_7644,N_6487);
nor UO_130 (O_130,N_5711,N_6045);
nand UO_131 (O_131,N_7003,N_7061);
and UO_132 (O_132,N_8017,N_9244);
nand UO_133 (O_133,N_7119,N_6007);
nand UO_134 (O_134,N_5451,N_5174);
and UO_135 (O_135,N_5319,N_5400);
nand UO_136 (O_136,N_9092,N_7740);
or UO_137 (O_137,N_6204,N_9154);
nand UO_138 (O_138,N_9330,N_6456);
or UO_139 (O_139,N_6366,N_6545);
or UO_140 (O_140,N_7698,N_5192);
or UO_141 (O_141,N_8683,N_9162);
and UO_142 (O_142,N_8284,N_6523);
nand UO_143 (O_143,N_9738,N_5065);
and UO_144 (O_144,N_6515,N_8705);
nor UO_145 (O_145,N_6645,N_7767);
nor UO_146 (O_146,N_8014,N_7100);
xnor UO_147 (O_147,N_6542,N_5272);
nor UO_148 (O_148,N_8228,N_7376);
or UO_149 (O_149,N_5873,N_5167);
nand UO_150 (O_150,N_9139,N_5098);
or UO_151 (O_151,N_7619,N_6466);
or UO_152 (O_152,N_6725,N_8280);
or UO_153 (O_153,N_7726,N_6748);
or UO_154 (O_154,N_8754,N_7191);
or UO_155 (O_155,N_9533,N_8196);
nor UO_156 (O_156,N_9827,N_8714);
nor UO_157 (O_157,N_5756,N_8740);
and UO_158 (O_158,N_6857,N_7399);
and UO_159 (O_159,N_6302,N_8925);
nor UO_160 (O_160,N_5729,N_9253);
nor UO_161 (O_161,N_8246,N_5112);
nor UO_162 (O_162,N_6937,N_5000);
nor UO_163 (O_163,N_5526,N_9638);
or UO_164 (O_164,N_8943,N_5774);
and UO_165 (O_165,N_5470,N_5713);
nor UO_166 (O_166,N_8880,N_5931);
nor UO_167 (O_167,N_5699,N_7932);
nand UO_168 (O_168,N_9933,N_6105);
and UO_169 (O_169,N_7705,N_7500);
nand UO_170 (O_170,N_9589,N_8253);
nand UO_171 (O_171,N_5654,N_5184);
nand UO_172 (O_172,N_6438,N_9020);
nand UO_173 (O_173,N_6860,N_5456);
nand UO_174 (O_174,N_6843,N_5717);
or UO_175 (O_175,N_9693,N_9331);
nand UO_176 (O_176,N_7990,N_5966);
and UO_177 (O_177,N_5050,N_8900);
and UO_178 (O_178,N_5993,N_5766);
or UO_179 (O_179,N_6702,N_5305);
nand UO_180 (O_180,N_5194,N_9982);
or UO_181 (O_181,N_8223,N_5678);
nand UO_182 (O_182,N_7962,N_9401);
nor UO_183 (O_183,N_9547,N_7649);
nand UO_184 (O_184,N_9768,N_7330);
or UO_185 (O_185,N_8069,N_6617);
and UO_186 (O_186,N_8382,N_5198);
nor UO_187 (O_187,N_7906,N_5660);
and UO_188 (O_188,N_8965,N_8625);
nand UO_189 (O_189,N_6465,N_8355);
or UO_190 (O_190,N_5469,N_5436);
and UO_191 (O_191,N_8640,N_6122);
nor UO_192 (O_192,N_5974,N_9167);
and UO_193 (O_193,N_9215,N_8083);
nand UO_194 (O_194,N_5532,N_8512);
nor UO_195 (O_195,N_8594,N_5429);
and UO_196 (O_196,N_5285,N_9630);
nand UO_197 (O_197,N_7547,N_7920);
nor UO_198 (O_198,N_7713,N_5235);
nor UO_199 (O_199,N_6670,N_7988);
or UO_200 (O_200,N_8499,N_7802);
or UO_201 (O_201,N_6796,N_8664);
nor UO_202 (O_202,N_8514,N_5425);
xor UO_203 (O_203,N_7093,N_8236);
nor UO_204 (O_204,N_7587,N_8459);
or UO_205 (O_205,N_5894,N_8813);
and UO_206 (O_206,N_5753,N_7839);
nand UO_207 (O_207,N_9498,N_5567);
nor UO_208 (O_208,N_5724,N_5536);
or UO_209 (O_209,N_8795,N_5022);
or UO_210 (O_210,N_7208,N_8645);
nand UO_211 (O_211,N_9834,N_9042);
nor UO_212 (O_212,N_9542,N_5102);
or UO_213 (O_213,N_6672,N_5787);
nand UO_214 (O_214,N_8146,N_8152);
or UO_215 (O_215,N_9564,N_9051);
or UO_216 (O_216,N_7148,N_5034);
or UO_217 (O_217,N_7048,N_8471);
or UO_218 (O_218,N_6429,N_8099);
nor UO_219 (O_219,N_6254,N_9782);
nand UO_220 (O_220,N_6338,N_8581);
nand UO_221 (O_221,N_9752,N_7614);
or UO_222 (O_222,N_7451,N_8378);
and UO_223 (O_223,N_5475,N_9038);
nand UO_224 (O_224,N_6311,N_5606);
nand UO_225 (O_225,N_6536,N_8593);
or UO_226 (O_226,N_7805,N_9047);
and UO_227 (O_227,N_5379,N_5009);
or UO_228 (O_228,N_5837,N_8262);
and UO_229 (O_229,N_8209,N_7914);
nor UO_230 (O_230,N_9041,N_8391);
nand UO_231 (O_231,N_6590,N_9067);
nand UO_232 (O_232,N_6616,N_5346);
nand UO_233 (O_233,N_5921,N_9122);
or UO_234 (O_234,N_6818,N_7372);
and UO_235 (O_235,N_9698,N_9454);
nand UO_236 (O_236,N_9976,N_6673);
nor UO_237 (O_237,N_9377,N_5277);
and UO_238 (O_238,N_8323,N_8487);
or UO_239 (O_239,N_9697,N_5196);
and UO_240 (O_240,N_6875,N_7758);
nor UO_241 (O_241,N_9731,N_8291);
or UO_242 (O_242,N_5506,N_9584);
and UO_243 (O_243,N_8263,N_8476);
or UO_244 (O_244,N_7720,N_8428);
nand UO_245 (O_245,N_5676,N_9074);
nand UO_246 (O_246,N_9710,N_8267);
nand UO_247 (O_247,N_6632,N_7186);
nor UO_248 (O_248,N_7798,N_6663);
nor UO_249 (O_249,N_7640,N_7452);
and UO_250 (O_250,N_5985,N_8332);
nor UO_251 (O_251,N_5303,N_8786);
and UO_252 (O_252,N_6942,N_9132);
or UO_253 (O_253,N_6754,N_5031);
or UO_254 (O_254,N_7924,N_5228);
or UO_255 (O_255,N_6154,N_6323);
or UO_256 (O_256,N_8447,N_6773);
nor UO_257 (O_257,N_9751,N_5955);
and UO_258 (O_258,N_7113,N_5005);
or UO_259 (O_259,N_9006,N_9537);
or UO_260 (O_260,N_7820,N_6389);
or UO_261 (O_261,N_8050,N_6495);
or UO_262 (O_262,N_5933,N_7625);
or UO_263 (O_263,N_6412,N_6155);
and UO_264 (O_264,N_7674,N_9459);
and UO_265 (O_265,N_7670,N_8618);
xor UO_266 (O_266,N_7420,N_9076);
or UO_267 (O_267,N_8611,N_8657);
nand UO_268 (O_268,N_9201,N_7922);
and UO_269 (O_269,N_5058,N_8766);
nand UO_270 (O_270,N_6385,N_9057);
nand UO_271 (O_271,N_8044,N_8698);
or UO_272 (O_272,N_5214,N_7370);
nand UO_273 (O_273,N_9937,N_8674);
and UO_274 (O_274,N_8073,N_6440);
and UO_275 (O_275,N_6270,N_8003);
nor UO_276 (O_276,N_8663,N_6241);
nor UO_277 (O_277,N_9129,N_9572);
nand UO_278 (O_278,N_5858,N_8838);
or UO_279 (O_279,N_8531,N_7944);
or UO_280 (O_280,N_6471,N_7537);
or UO_281 (O_281,N_8794,N_9759);
nand UO_282 (O_282,N_9274,N_8882);
nor UO_283 (O_283,N_7627,N_5424);
nor UO_284 (O_284,N_5101,N_9214);
nor UO_285 (O_285,N_5727,N_5845);
nor UO_286 (O_286,N_7630,N_7717);
and UO_287 (O_287,N_8028,N_7668);
nand UO_288 (O_288,N_7021,N_8747);
or UO_289 (O_289,N_6999,N_6468);
nand UO_290 (O_290,N_5066,N_5641);
or UO_291 (O_291,N_6350,N_5973);
and UO_292 (O_292,N_9929,N_6346);
or UO_293 (O_293,N_9928,N_7423);
or UO_294 (O_294,N_8252,N_9718);
nor UO_295 (O_295,N_5679,N_6599);
and UO_296 (O_296,N_8828,N_7096);
nor UO_297 (O_297,N_9793,N_9494);
and UO_298 (O_298,N_6029,N_9222);
or UO_299 (O_299,N_7097,N_8905);
nand UO_300 (O_300,N_5309,N_8086);
or UO_301 (O_301,N_7050,N_5004);
and UO_302 (O_302,N_6289,N_7610);
nand UO_303 (O_303,N_5090,N_6319);
and UO_304 (O_304,N_6170,N_6747);
nand UO_305 (O_305,N_9645,N_7147);
nor UO_306 (O_306,N_5788,N_9717);
nor UO_307 (O_307,N_6475,N_9691);
nand UO_308 (O_308,N_5885,N_6908);
nor UO_309 (O_309,N_8396,N_9460);
or UO_310 (O_310,N_9390,N_8436);
nor UO_311 (O_311,N_6858,N_5956);
or UO_312 (O_312,N_7176,N_5339);
or UO_313 (O_313,N_6335,N_7417);
nand UO_314 (O_314,N_7548,N_9666);
nor UO_315 (O_315,N_7731,N_9746);
nand UO_316 (O_316,N_7282,N_9840);
nand UO_317 (O_317,N_7997,N_9993);
or UO_318 (O_318,N_8577,N_8693);
or UO_319 (O_319,N_5143,N_7192);
nor UO_320 (O_320,N_5854,N_6709);
nand UO_321 (O_321,N_5430,N_5007);
nor UO_322 (O_322,N_5516,N_7105);
and UO_323 (O_323,N_8820,N_7324);
nor UO_324 (O_324,N_5643,N_5441);
nand UO_325 (O_325,N_8311,N_9466);
nor UO_326 (O_326,N_6248,N_5299);
and UO_327 (O_327,N_7373,N_6214);
and UO_328 (O_328,N_9734,N_8317);
or UO_329 (O_329,N_8639,N_6285);
nand UO_330 (O_330,N_5474,N_6499);
nor UO_331 (O_331,N_5575,N_6647);
or UO_332 (O_332,N_8761,N_7756);
and UO_333 (O_333,N_9463,N_8404);
and UO_334 (O_334,N_9310,N_6485);
nor UO_335 (O_335,N_9562,N_5646);
and UO_336 (O_336,N_6130,N_8364);
nor UO_337 (O_337,N_9145,N_5959);
nand UO_338 (O_338,N_7809,N_9581);
or UO_339 (O_339,N_5534,N_7463);
or UO_340 (O_340,N_5138,N_7957);
nor UO_341 (O_341,N_6354,N_7590);
and UO_342 (O_342,N_5640,N_9821);
or UO_343 (O_343,N_7696,N_6033);
and UO_344 (O_344,N_5806,N_5159);
or UO_345 (O_345,N_5969,N_6895);
or UO_346 (O_346,N_7182,N_8417);
nor UO_347 (O_347,N_7259,N_8759);
or UO_348 (O_348,N_5680,N_6537);
nor UO_349 (O_349,N_7174,N_5444);
nand UO_350 (O_350,N_7570,N_8226);
nor UO_351 (O_351,N_6189,N_9803);
and UO_352 (O_352,N_6953,N_6134);
or UO_353 (O_353,N_5498,N_7804);
or UO_354 (O_354,N_9409,N_7525);
and UO_355 (O_355,N_8424,N_8045);
or UO_356 (O_356,N_5883,N_6981);
and UO_357 (O_357,N_7131,N_7666);
and UO_358 (O_358,N_9147,N_6002);
nor UO_359 (O_359,N_9480,N_8865);
nor UO_360 (O_360,N_5877,N_9128);
nand UO_361 (O_361,N_8316,N_6178);
and UO_362 (O_362,N_9776,N_8558);
or UO_363 (O_363,N_5764,N_6887);
and UO_364 (O_364,N_5122,N_9016);
nand UO_365 (O_365,N_5171,N_9143);
or UO_366 (O_366,N_6788,N_6524);
nor UO_367 (O_367,N_6127,N_9258);
and UO_368 (O_368,N_9236,N_6182);
nor UO_369 (O_369,N_5908,N_7116);
or UO_370 (O_370,N_7939,N_5263);
and UO_371 (O_371,N_8659,N_7654);
and UO_372 (O_372,N_7854,N_5074);
nor UO_373 (O_373,N_9830,N_6574);
nor UO_374 (O_374,N_6423,N_8057);
and UO_375 (O_375,N_6947,N_5687);
or UO_376 (O_376,N_9135,N_9393);
or UO_377 (O_377,N_7473,N_5088);
or UO_378 (O_378,N_8283,N_8530);
nor UO_379 (O_379,N_6994,N_9785);
or UO_380 (O_380,N_7261,N_6975);
and UO_381 (O_381,N_8742,N_9680);
and UO_382 (O_382,N_8320,N_7108);
or UO_383 (O_383,N_7388,N_5290);
or UO_384 (O_384,N_5674,N_6202);
nand UO_385 (O_385,N_5628,N_7427);
nor UO_386 (O_386,N_7078,N_9438);
nor UO_387 (O_387,N_8845,N_7824);
xnor UO_388 (O_388,N_6827,N_6586);
nand UO_389 (O_389,N_7084,N_7224);
nor UO_390 (O_390,N_6688,N_5404);
or UO_391 (O_391,N_9068,N_6054);
or UO_392 (O_392,N_7323,N_5310);
nand UO_393 (O_393,N_5971,N_8140);
nor UO_394 (O_394,N_8580,N_7994);
xor UO_395 (O_395,N_6630,N_7059);
nand UO_396 (O_396,N_7877,N_7827);
and UO_397 (O_397,N_9512,N_6201);
and UO_398 (O_398,N_8737,N_5736);
nand UO_399 (O_399,N_8161,N_5216);
nand UO_400 (O_400,N_5266,N_5123);
nand UO_401 (O_401,N_6581,N_5423);
and UO_402 (O_402,N_9340,N_5357);
or UO_403 (O_403,N_9712,N_8264);
nor UO_404 (O_404,N_9354,N_7822);
and UO_405 (O_405,N_9155,N_6120);
nand UO_406 (O_406,N_5313,N_8879);
xor UO_407 (O_407,N_7203,N_5892);
or UO_408 (O_408,N_8739,N_7066);
xnor UO_409 (O_409,N_5619,N_5367);
and UO_410 (O_410,N_5665,N_7361);
nor UO_411 (O_411,N_9799,N_7911);
nand UO_412 (O_412,N_8812,N_7209);
nand UO_413 (O_413,N_7236,N_5352);
nand UO_414 (O_414,N_5721,N_9133);
and UO_415 (O_415,N_6434,N_9859);
nand UO_416 (O_416,N_6983,N_7978);
or UO_417 (O_417,N_8899,N_6770);
nor UO_418 (O_418,N_8897,N_6933);
nand UO_419 (O_419,N_7928,N_9807);
and UO_420 (O_420,N_7618,N_9647);
nor UO_421 (O_421,N_5706,N_6313);
xor UO_422 (O_422,N_9005,N_8442);
and UO_423 (O_423,N_9682,N_9602);
nand UO_424 (O_424,N_6901,N_8123);
xnor UO_425 (O_425,N_7120,N_9798);
nor UO_426 (O_426,N_8765,N_9209);
or UO_427 (O_427,N_8517,N_7746);
nor UO_428 (O_428,N_7193,N_6386);
nand UO_429 (O_429,N_9822,N_6868);
nor UO_430 (O_430,N_5241,N_6250);
and UO_431 (O_431,N_8271,N_6474);
or UO_432 (O_432,N_6446,N_8604);
and UO_433 (O_433,N_8709,N_8807);
nor UO_434 (O_434,N_6351,N_8473);
nor UO_435 (O_435,N_6494,N_7213);
nor UO_436 (O_436,N_8961,N_8232);
and UO_437 (O_437,N_5134,N_7198);
and UO_438 (O_438,N_5942,N_7813);
and UO_439 (O_439,N_8589,N_6806);
nor UO_440 (O_440,N_6356,N_9973);
or UO_441 (O_441,N_6793,N_6711);
or UO_442 (O_442,N_6444,N_7799);
and UO_443 (O_443,N_6948,N_9399);
and UO_444 (O_444,N_8483,N_8215);
nor UO_445 (O_445,N_5358,N_8907);
nor UO_446 (O_446,N_7359,N_8124);
nand UO_447 (O_447,N_9837,N_6145);
and UO_448 (O_448,N_7008,N_5338);
nor UO_449 (O_449,N_8930,N_9050);
and UO_450 (O_450,N_5781,N_7849);
or UO_451 (O_451,N_7727,N_5321);
nand UO_452 (O_452,N_7041,N_6417);
nand UO_453 (O_453,N_6462,N_9037);
nand UO_454 (O_454,N_5968,N_9156);
and UO_455 (O_455,N_8569,N_7112);
nand UO_456 (O_456,N_6825,N_5600);
nor UO_457 (O_457,N_9846,N_9090);
or UO_458 (O_458,N_9700,N_7117);
nand UO_459 (O_459,N_5157,N_6556);
nand UO_460 (O_460,N_8718,N_8210);
and UO_461 (O_461,N_7276,N_8344);
and UO_462 (O_462,N_9371,N_8279);
nor UO_463 (O_463,N_9269,N_6866);
nor UO_464 (O_464,N_7413,N_5497);
nand UO_465 (O_465,N_5482,N_7903);
or UO_466 (O_466,N_5032,N_8205);
nor UO_467 (O_467,N_9062,N_7161);
or UO_468 (O_468,N_6303,N_5524);
and UO_469 (O_469,N_8005,N_5926);
and UO_470 (O_470,N_8842,N_5856);
nor UO_471 (O_471,N_6618,N_8448);
or UO_472 (O_472,N_7757,N_7788);
nor UO_473 (O_473,N_8368,N_9954);
nor UO_474 (O_474,N_8689,N_5884);
or UO_475 (O_475,N_9916,N_6900);
nand UO_476 (O_476,N_9729,N_7099);
and UO_477 (O_477,N_6098,N_6982);
or UO_478 (O_478,N_6060,N_5193);
nor UO_479 (O_479,N_7241,N_6980);
or UO_480 (O_480,N_7444,N_6264);
or UO_481 (O_481,N_7390,N_5048);
and UO_482 (O_482,N_6441,N_6040);
nand UO_483 (O_483,N_8117,N_8792);
nor UO_484 (O_484,N_7341,N_8539);
or UO_485 (O_485,N_8427,N_7412);
or UO_486 (O_486,N_8735,N_7303);
nor UO_487 (O_487,N_6206,N_6433);
nand UO_488 (O_488,N_6288,N_7556);
nand UO_489 (O_489,N_5248,N_9141);
and UO_490 (O_490,N_6690,N_7086);
nor UO_491 (O_491,N_5761,N_7908);
nand UO_492 (O_492,N_5394,N_9550);
nand UO_493 (O_493,N_8324,N_7509);
and UO_494 (O_494,N_8712,N_8058);
or UO_495 (O_495,N_6372,N_6381);
or UO_496 (O_496,N_8723,N_5190);
nor UO_497 (O_497,N_8869,N_6940);
or UO_498 (O_498,N_8939,N_9539);
and UO_499 (O_499,N_5547,N_7620);
and UO_500 (O_500,N_6021,N_7036);
nor UO_501 (O_501,N_5936,N_6020);
and UO_502 (O_502,N_5677,N_7432);
nand UO_503 (O_503,N_7153,N_7524);
and UO_504 (O_504,N_9229,N_5720);
nor UO_505 (O_505,N_9254,N_6185);
nand UO_506 (O_506,N_6560,N_6669);
and UO_507 (O_507,N_6625,N_5222);
and UO_508 (O_508,N_9086,N_6197);
nor UO_509 (O_509,N_5768,N_8720);
nor UO_510 (O_510,N_6897,N_5462);
nand UO_511 (O_511,N_7502,N_5386);
nand UO_512 (O_512,N_9286,N_5561);
nand UO_513 (O_513,N_6587,N_9078);
and UO_514 (O_514,N_5629,N_5287);
nand UO_515 (O_515,N_9120,N_7659);
and UO_516 (O_516,N_6181,N_7501);
and UO_517 (O_517,N_6151,N_8622);
xnor UO_518 (O_518,N_5984,N_5920);
and UO_519 (O_519,N_8860,N_5882);
or UO_520 (O_520,N_9484,N_5271);
or UO_521 (O_521,N_7760,N_7761);
nand UO_522 (O_522,N_5958,N_8486);
nand UO_523 (O_523,N_6539,N_6922);
nand UO_524 (O_524,N_6591,N_9355);
and UO_525 (O_525,N_8451,N_9312);
and UO_526 (O_526,N_8988,N_7952);
nor UO_527 (O_527,N_9184,N_6492);
nor UO_528 (O_528,N_5316,N_6174);
and UO_529 (O_529,N_9381,N_6817);
nand UO_530 (O_530,N_7869,N_9600);
nor UO_531 (O_531,N_8170,N_7560);
and UO_532 (O_532,N_6163,N_8118);
nand UO_533 (O_533,N_5797,N_5260);
or UO_534 (O_534,N_7738,N_7956);
and UO_535 (O_535,N_5543,N_9857);
nor UO_536 (O_536,N_8156,N_9932);
or UO_537 (O_537,N_5083,N_6220);
and UO_538 (O_538,N_5261,N_5021);
nor UO_539 (O_539,N_5364,N_7543);
nor UO_540 (O_540,N_7381,N_8134);
or UO_541 (O_541,N_9417,N_9488);
nand UO_542 (O_542,N_6715,N_7322);
nand UO_543 (O_543,N_5525,N_9590);
nand UO_544 (O_544,N_6919,N_9018);
or UO_545 (O_545,N_7234,N_7968);
nand UO_546 (O_546,N_9096,N_6522);
nand UO_547 (O_547,N_6101,N_8585);
or UO_548 (O_548,N_6430,N_6576);
nor UO_549 (O_549,N_7394,N_8165);
and UO_550 (O_550,N_8632,N_9668);
or UO_551 (O_551,N_5215,N_9028);
or UO_552 (O_552,N_8655,N_7288);
nand UO_553 (O_553,N_6534,N_5871);
or UO_554 (O_554,N_5983,N_9360);
nor UO_555 (O_555,N_6215,N_7980);
and UO_556 (O_556,N_7143,N_6580);
nor UO_557 (O_557,N_5596,N_8334);
and UO_558 (O_558,N_5855,N_5565);
and UO_559 (O_559,N_5529,N_5531);
nand UO_560 (O_560,N_5938,N_6657);
nor UO_561 (O_561,N_9440,N_7977);
or UO_562 (O_562,N_6734,N_5518);
nand UO_563 (O_563,N_7421,N_8490);
nand UO_564 (O_564,N_8258,N_5822);
and UO_565 (O_565,N_5270,N_8621);
or UO_566 (O_566,N_9977,N_5631);
or UO_567 (O_567,N_7563,N_6501);
and UO_568 (O_568,N_6016,N_8967);
nand UO_569 (O_569,N_5042,N_6749);
or UO_570 (O_570,N_7553,N_7708);
or UO_571 (O_571,N_9243,N_5655);
and UO_572 (O_572,N_5383,N_6892);
nand UO_573 (O_573,N_9825,N_8125);
nor UO_574 (O_574,N_6782,N_8192);
or UO_575 (O_575,N_6513,N_6161);
and UO_576 (O_576,N_5002,N_7039);
nand UO_577 (O_577,N_5508,N_7235);
and UO_578 (O_578,N_8576,N_5954);
and UO_579 (O_579,N_6428,N_5039);
nor UO_580 (O_580,N_8128,N_6437);
nand UO_581 (O_581,N_9823,N_9085);
or UO_582 (O_582,N_6707,N_8921);
nor UO_583 (O_583,N_5455,N_7366);
nor UO_584 (O_584,N_8400,N_5117);
nand UO_585 (O_585,N_7800,N_7419);
nand UO_586 (O_586,N_8504,N_7484);
nand UO_587 (O_587,N_5179,N_8901);
nor UO_588 (O_588,N_5273,N_8162);
or UO_589 (O_589,N_6362,N_8858);
nand UO_590 (O_590,N_9483,N_7284);
nand UO_591 (O_591,N_6743,N_9481);
nand UO_592 (O_592,N_9080,N_9995);
and UO_593 (O_593,N_7966,N_6593);
and UO_594 (O_594,N_7764,N_8619);
or UO_595 (O_595,N_6853,N_8862);
and UO_596 (O_596,N_5744,N_5994);
or UO_597 (O_597,N_9045,N_7136);
and UO_598 (O_598,N_9771,N_6299);
and UO_599 (O_599,N_8462,N_9192);
and UO_600 (O_600,N_9308,N_9242);
nor UO_601 (O_601,N_6157,N_5049);
and UO_602 (O_602,N_6146,N_7440);
and UO_603 (O_603,N_7462,N_6962);
nor UO_604 (O_604,N_6526,N_8015);
nor UO_605 (O_605,N_8788,N_9761);
or UO_606 (O_606,N_5512,N_9990);
nor UO_607 (O_607,N_9906,N_7025);
and UO_608 (O_608,N_7374,N_5541);
and UO_609 (O_609,N_8360,N_7240);
or UO_610 (O_610,N_7023,N_9801);
and UO_611 (O_611,N_8752,N_9026);
nor UO_612 (O_612,N_8546,N_6044);
and UO_613 (O_613,N_8653,N_8023);
or UO_614 (O_614,N_7405,N_6619);
or UO_615 (O_615,N_8524,N_5598);
nor UO_616 (O_616,N_7825,N_7750);
or UO_617 (O_617,N_5396,N_6623);
or UO_618 (O_618,N_7734,N_9856);
or UO_619 (O_619,N_7897,N_8651);
nand UO_620 (O_620,N_5162,N_8175);
or UO_621 (O_621,N_6547,N_7858);
xor UO_622 (O_622,N_6746,N_5237);
nor UO_623 (O_623,N_9033,N_9219);
and UO_624 (O_624,N_9406,N_5742);
and UO_625 (O_625,N_8510,N_5897);
and UO_626 (O_626,N_8658,N_6243);
or UO_627 (O_627,N_9628,N_6239);
nor UO_628 (O_628,N_6765,N_6073);
or UO_629 (O_629,N_5556,N_9011);
or UO_630 (O_630,N_8251,N_9659);
or UO_631 (O_631,N_9241,N_7947);
nor UO_632 (O_632,N_6304,N_9621);
nor UO_633 (O_633,N_7954,N_9523);
or UO_634 (O_634,N_7199,N_8928);
xnor UO_635 (O_635,N_6791,N_7605);
and UO_636 (O_636,N_6877,N_9328);
or UO_637 (O_637,N_6034,N_7031);
nand UO_638 (O_638,N_6807,N_7154);
or UO_639 (O_639,N_6615,N_9297);
and UO_640 (O_640,N_6927,N_9216);
nand UO_641 (O_641,N_7058,N_5365);
and UO_642 (O_642,N_6559,N_5356);
nand UO_643 (O_643,N_6516,N_7815);
or UO_644 (O_644,N_7453,N_5262);
and UO_645 (O_645,N_8875,N_9191);
and UO_646 (O_646,N_9792,N_6541);
nand UO_647 (O_647,N_9282,N_8620);
or UO_648 (O_648,N_6689,N_8730);
and UO_649 (O_649,N_8923,N_9307);
and UO_650 (O_650,N_7831,N_6207);
nand UO_651 (O_651,N_8272,N_6589);
or UO_652 (O_652,N_8214,N_9515);
nand UO_653 (O_653,N_6820,N_5170);
and UO_654 (O_654,N_7901,N_9553);
nand UO_655 (O_655,N_7081,N_7312);
nor UO_656 (O_656,N_6662,N_5180);
and UO_657 (O_657,N_6610,N_6588);
nand UO_658 (O_658,N_8912,N_6442);
or UO_659 (O_659,N_6525,N_5211);
or UO_660 (O_660,N_7594,N_7126);
nand UO_661 (O_661,N_9239,N_8310);
nand UO_662 (O_662,N_5616,N_6017);
and UO_663 (O_663,N_6938,N_6307);
or UO_664 (O_664,N_6074,N_6400);
or UO_665 (O_665,N_7648,N_7852);
nor UO_666 (O_666,N_9905,N_5036);
or UO_667 (O_667,N_9795,N_7094);
nor UO_668 (O_668,N_9545,N_5251);
nand UO_669 (O_669,N_7703,N_6814);
nand UO_670 (O_670,N_5240,N_6129);
or UO_671 (O_671,N_6924,N_7565);
nand UO_672 (O_672,N_9656,N_7163);
nand UO_673 (O_673,N_8392,N_8571);
and UO_674 (O_674,N_7721,N_6819);
and UO_675 (O_675,N_5369,N_7395);
nor UO_676 (O_676,N_8595,N_6418);
or UO_677 (O_677,N_6965,N_8991);
and UO_678 (O_678,N_7843,N_9031);
nor UO_679 (O_679,N_8164,N_7996);
and UO_680 (O_680,N_6869,N_9858);
and UO_681 (O_681,N_6731,N_5593);
nand UO_682 (O_682,N_9855,N_9684);
and UO_683 (O_683,N_5757,N_8670);
nand UO_684 (O_684,N_7778,N_5763);
nor UO_685 (O_685,N_6200,N_5139);
nand UO_686 (O_686,N_5989,N_8479);
and UO_687 (O_687,N_8061,N_6861);
or UO_688 (O_688,N_6693,N_5686);
and UO_689 (O_689,N_8119,N_7149);
and UO_690 (O_690,N_6053,N_7249);
and UO_691 (O_691,N_9213,N_5247);
nand UO_692 (O_692,N_7064,N_6741);
nand UO_693 (O_693,N_5293,N_5332);
nor UO_694 (O_694,N_8309,N_7621);
or UO_695 (O_695,N_9185,N_9225);
or UO_696 (O_696,N_8408,N_9860);
or UO_697 (O_697,N_5477,N_5077);
and UO_698 (O_698,N_5818,N_7286);
nand UO_699 (O_699,N_5953,N_7190);
and UO_700 (O_700,N_8966,N_9678);
xor UO_701 (O_701,N_9608,N_8667);
nand UO_702 (O_702,N_6529,N_6051);
or UO_703 (O_703,N_7083,N_9842);
and UO_704 (O_704,N_8774,N_7258);
nand UO_705 (O_705,N_6620,N_8352);
nand UO_706 (O_706,N_8725,N_5519);
nor UO_707 (O_707,N_9098,N_6031);
and UO_708 (O_708,N_8502,N_8401);
or UO_709 (O_709,N_8041,N_6608);
nand UO_710 (O_710,N_6511,N_7566);
and UO_711 (O_711,N_9376,N_7307);
or UO_712 (O_712,N_5069,N_9295);
and UO_713 (O_713,N_6388,N_6324);
or UO_714 (O_714,N_8095,N_6297);
and UO_715 (O_715,N_5473,N_6359);
nand UO_716 (O_716,N_8470,N_9888);
nor UO_717 (O_717,N_8184,N_8544);
xor UO_718 (O_718,N_5765,N_6729);
nand UO_719 (O_719,N_8904,N_9469);
nand UO_720 (O_720,N_7125,N_7599);
nand UO_721 (O_721,N_7109,N_9908);
nand UO_722 (O_722,N_5354,N_9790);
xnor UO_723 (O_723,N_6802,N_6310);
nand UO_724 (O_724,N_9025,N_7263);
nand UO_725 (O_725,N_7626,N_6008);
or UO_726 (O_726,N_6432,N_7029);
and UO_727 (O_727,N_9959,N_9359);
and UO_728 (O_728,N_9470,N_9648);
and UO_729 (O_729,N_7604,N_9508);
nor UO_730 (O_730,N_5943,N_9540);
nor UO_731 (O_731,N_8075,N_6500);
or UO_732 (O_732,N_6126,N_6049);
or UO_733 (O_733,N_6585,N_5823);
and UO_734 (O_734,N_9043,N_9695);
or UO_735 (O_735,N_7273,N_8506);
and UO_736 (O_736,N_5362,N_5592);
or UO_737 (O_737,N_8535,N_7055);
and UO_738 (O_738,N_6399,N_7004);
and UO_739 (O_739,N_9911,N_9370);
or UO_740 (O_740,N_8241,N_8523);
nand UO_741 (O_741,N_8217,N_8449);
nor UO_742 (O_742,N_8030,N_5045);
nor UO_743 (O_743,N_7677,N_5650);
nand UO_744 (O_744,N_9820,N_9164);
nor UO_745 (O_745,N_5478,N_6282);
nor UO_746 (O_746,N_8206,N_7496);
or UO_747 (O_747,N_8822,N_7087);
or UO_748 (O_748,N_7929,N_5785);
nand UO_749 (O_749,N_9273,N_7140);
nor UO_750 (O_750,N_7985,N_9385);
nand UO_751 (O_751,N_7406,N_5027);
nand UO_752 (O_752,N_5238,N_9281);
or UO_753 (O_753,N_8941,N_5834);
or UO_754 (O_754,N_9436,N_6607);
or UO_755 (O_755,N_6006,N_8550);
or UO_756 (O_756,N_5043,N_6380);
nand UO_757 (O_757,N_8644,N_6624);
nor UO_758 (O_758,N_9346,N_6367);
nand UO_759 (O_759,N_7194,N_9300);
nand UO_760 (O_760,N_5393,N_7790);
or UO_761 (O_761,N_8722,N_8343);
nor UO_762 (O_762,N_8489,N_7027);
and UO_763 (O_763,N_5351,N_6566);
or UO_764 (O_764,N_7612,N_8475);
and UO_765 (O_765,N_8342,N_9134);
nand UO_766 (O_766,N_9975,N_6553);
and UO_767 (O_767,N_5087,N_6427);
and UO_768 (O_768,N_5793,N_5132);
nand UO_769 (O_769,N_8783,N_6043);
nor UO_770 (O_770,N_8847,N_8327);
and UO_771 (O_771,N_8060,N_9365);
or UO_772 (O_772,N_7408,N_6218);
and UO_773 (O_773,N_6327,N_6281);
xor UO_774 (O_774,N_8855,N_7486);
or UO_775 (O_775,N_8029,N_8637);
nor UO_776 (O_776,N_9083,N_5168);
or UO_777 (O_777,N_6148,N_5569);
nand UO_778 (O_778,N_7400,N_8958);
or UO_779 (O_779,N_8306,N_5427);
nand UO_780 (O_780,N_7972,N_8296);
and UO_781 (O_781,N_9064,N_8891);
nand UO_782 (O_782,N_7195,N_9887);
and UO_783 (O_783,N_9278,N_9942);
xnor UO_784 (O_784,N_9978,N_5951);
nor UO_785 (O_785,N_7415,N_7431);
nor UO_786 (O_786,N_7202,N_9702);
nor UO_787 (O_787,N_5368,N_7995);
nor UO_788 (O_788,N_9449,N_5924);
and UO_789 (O_789,N_6968,N_7774);
nor UO_790 (O_790,N_6512,N_5057);
and UO_791 (O_791,N_5617,N_6000);
nor UO_792 (O_792,N_9160,N_8349);
and UO_793 (O_793,N_5113,N_7979);
nand UO_794 (O_794,N_8203,N_8179);
nand UO_795 (O_795,N_6115,N_5863);
or UO_796 (O_796,N_6175,N_5671);
nand UO_797 (O_797,N_7794,N_8691);
or UO_798 (O_798,N_9467,N_9555);
and UO_799 (O_799,N_6010,N_6745);
nor UO_800 (O_800,N_8746,N_5264);
or UO_801 (O_801,N_6136,N_9157);
nor UO_802 (O_802,N_8687,N_9631);
and UO_803 (O_803,N_7793,N_7991);
and UO_804 (O_804,N_9276,N_8482);
and UO_805 (O_805,N_7829,N_7690);
nand UO_806 (O_806,N_9692,N_7645);
or UO_807 (O_807,N_5624,N_6091);
nand UO_808 (O_808,N_5552,N_6376);
nor UO_809 (O_809,N_5278,N_8269);
nor UO_810 (O_810,N_5770,N_5242);
or UO_811 (O_811,N_8022,N_8051);
nor UO_812 (O_812,N_6949,N_8078);
nor UO_813 (O_813,N_8911,N_7175);
nand UO_814 (O_814,N_6579,N_5325);
nor UO_815 (O_815,N_9576,N_6436);
and UO_816 (O_816,N_9251,N_8784);
nand UO_817 (O_817,N_9764,N_8727);
nor UO_818 (O_818,N_9935,N_5509);
nor UO_819 (O_819,N_9535,N_8805);
nand UO_820 (O_820,N_7404,N_6358);
or UO_821 (O_821,N_8613,N_6081);
nand UO_822 (O_822,N_6251,N_7970);
nand UO_823 (O_823,N_6719,N_9400);
nand UO_824 (O_824,N_9897,N_6269);
or UO_825 (O_825,N_9126,N_6926);
or UO_826 (O_826,N_9781,N_9177);
or UO_827 (O_827,N_7925,N_8158);
and UO_828 (O_828,N_8288,N_9797);
or UO_829 (O_829,N_9974,N_8677);
or UO_830 (O_830,N_9450,N_8521);
or UO_831 (O_831,N_9485,N_9476);
nor UO_832 (O_832,N_5081,N_6906);
or UO_833 (O_833,N_5843,N_8744);
nand UO_834 (O_834,N_9250,N_8260);
and UO_835 (O_835,N_7168,N_5317);
nand UO_836 (O_836,N_5391,N_6596);
nand UO_837 (O_837,N_9364,N_9159);
nor UO_838 (O_838,N_6333,N_8975);
or UO_839 (O_839,N_8248,N_5867);
nand UO_840 (O_840,N_5274,N_5495);
and UO_841 (O_841,N_7455,N_6780);
nor UO_842 (O_842,N_7216,N_9848);
or UO_843 (O_843,N_7526,N_6205);
or UO_844 (O_844,N_5208,N_9586);
or UO_845 (O_845,N_6273,N_5782);
and UO_846 (O_846,N_6227,N_5297);
nand UO_847 (O_847,N_8157,N_7961);
and UO_848 (O_848,N_6832,N_8831);
and UO_849 (O_849,N_8839,N_8559);
or UO_850 (O_850,N_8405,N_7528);
nor UO_851 (O_851,N_5412,N_7494);
and UO_852 (O_852,N_7049,N_8946);
nand UO_853 (O_853,N_8648,N_7456);
and UO_854 (O_854,N_7157,N_9646);
nand UO_855 (O_855,N_7211,N_8000);
nor UO_856 (O_856,N_6171,N_5376);
nand UO_857 (O_857,N_8026,N_8692);
and UO_858 (O_858,N_5990,N_6331);
nor UO_859 (O_859,N_9427,N_7728);
or UO_860 (O_860,N_5438,N_9568);
nand UO_861 (O_861,N_5347,N_9144);
nand UO_862 (O_862,N_5496,N_6450);
nor UO_863 (O_863,N_9875,N_8358);
nor UO_864 (O_864,N_8541,N_5510);
and UO_865 (O_865,N_9421,N_8319);
nor UO_866 (O_866,N_5126,N_9690);
nand UO_867 (O_867,N_9112,N_6776);
and UO_868 (O_868,N_7684,N_7542);
or UO_869 (O_869,N_7574,N_9046);
nor UO_870 (O_870,N_9871,N_9195);
and UO_871 (O_871,N_9453,N_9337);
nor UO_872 (O_872,N_7289,N_7356);
nor UO_873 (O_873,N_7866,N_7205);
nor UO_874 (O_874,N_5707,N_6025);
or UO_875 (O_875,N_6050,N_6830);
nor UO_876 (O_876,N_6961,N_9091);
or UO_877 (O_877,N_7056,N_9221);
nor UO_878 (O_878,N_8292,N_7971);
nand UO_879 (O_879,N_9941,N_9876);
nor UO_880 (O_880,N_8294,N_7051);
and UO_881 (O_881,N_6701,N_8833);
nand UO_882 (O_882,N_7115,N_6079);
nor UO_883 (O_883,N_6703,N_8836);
nor UO_884 (O_884,N_9339,N_9735);
nor UO_885 (O_885,N_5020,N_7034);
or UO_886 (O_886,N_8213,N_5111);
nand UO_887 (O_887,N_6891,N_6727);
and UO_888 (O_888,N_8877,N_6979);
or UO_889 (O_889,N_8690,N_7657);
or UO_890 (O_890,N_7340,N_5053);
nor UO_891 (O_891,N_9341,N_7476);
and UO_892 (O_892,N_5670,N_7118);
and UO_893 (O_893,N_5528,N_8289);
or UO_894 (O_894,N_6737,N_7706);
nand UO_895 (O_895,N_5917,N_7608);
xnor UO_896 (O_896,N_6449,N_7010);
or UO_897 (O_897,N_5771,N_6244);
nand UO_898 (O_898,N_6583,N_7617);
nor UO_899 (O_899,N_7886,N_6721);
or UO_900 (O_900,N_9800,N_7210);
nand UO_901 (O_901,N_9081,N_8211);
nor UO_902 (O_902,N_5709,N_5568);
and UO_903 (O_903,N_5746,N_7685);
and UO_904 (O_904,N_8764,N_5059);
nor UO_905 (O_905,N_7576,N_8429);
or UO_906 (O_906,N_7121,N_5811);
or UO_907 (O_907,N_5182,N_7301);
nand UO_908 (O_908,N_7782,N_6398);
nor UO_909 (O_909,N_9558,N_6022);
and UO_910 (O_910,N_6015,N_5513);
nand UO_911 (O_911,N_9758,N_6164);
or UO_912 (O_912,N_9332,N_7350);
nor UO_913 (O_913,N_8249,N_5545);
nand UO_914 (O_914,N_8532,N_8200);
or UO_915 (O_915,N_9285,N_7821);
nand UO_916 (O_916,N_8093,N_9099);
or UO_917 (O_917,N_9607,N_7896);
nor UO_918 (O_918,N_6210,N_8067);
or UO_919 (O_919,N_5125,N_7633);
and UO_920 (O_920,N_5997,N_7107);
or UO_921 (O_921,N_8088,N_5900);
and UO_922 (O_922,N_6345,N_8821);
nand UO_923 (O_923,N_9416,N_6460);
nand UO_924 (O_924,N_6987,N_5988);
nand UO_925 (O_925,N_9324,N_6598);
and UO_926 (O_926,N_6736,N_8133);
xnor UO_927 (O_927,N_5209,N_8143);
and UO_928 (O_928,N_7643,N_8533);
or UO_929 (O_929,N_7959,N_5361);
or UO_930 (O_930,N_9125,N_7856);
nand UO_931 (O_931,N_7857,N_5380);
nand UO_932 (O_932,N_8496,N_7629);
nand UO_933 (O_933,N_9593,N_7510);
nand UO_934 (O_934,N_9787,N_7786);
or UO_935 (O_935,N_6392,N_9657);
nor UO_936 (O_936,N_9309,N_9854);
or UO_937 (O_937,N_8895,N_8281);
nor UO_938 (O_938,N_9383,N_6482);
or UO_939 (O_939,N_7691,N_8874);
nand UO_940 (O_940,N_8130,N_8386);
nand UO_941 (O_941,N_7020,N_5730);
nand UO_942 (O_942,N_5551,N_9093);
nand UO_943 (O_943,N_8970,N_8176);
and UO_944 (O_944,N_6592,N_7428);
and UO_945 (O_945,N_7201,N_6133);
nand UO_946 (O_946,N_8824,N_6396);
or UO_947 (O_947,N_9794,N_6448);
nor UO_948 (O_948,N_7159,N_5638);
or UO_949 (O_949,N_5916,N_9578);
nand UO_950 (O_950,N_8750,N_8074);
or UO_951 (O_951,N_6461,N_7378);
and UO_952 (O_952,N_9275,N_9660);
nor UO_953 (O_953,N_8350,N_8602);
and UO_954 (O_954,N_5805,N_6898);
nand UO_955 (O_955,N_7837,N_6284);
or UO_956 (O_956,N_7974,N_7545);
or UO_957 (O_957,N_9198,N_6086);
nor UO_958 (O_958,N_5769,N_5428);
nand UO_959 (O_959,N_8155,N_5664);
and UO_960 (O_960,N_9437,N_7650);
and UO_961 (O_961,N_7572,N_8187);
nor UO_962 (O_962,N_6544,N_8488);
nor UO_963 (O_963,N_5972,N_5976);
nand UO_964 (O_964,N_7271,N_6414);
nand UO_965 (O_965,N_7863,N_7142);
nand UO_966 (O_966,N_8463,N_9408);
and UO_967 (O_967,N_7274,N_8347);
and UO_968 (O_968,N_8728,N_7231);
nor UO_969 (O_969,N_5373,N_6921);
nand UO_970 (O_970,N_6242,N_6212);
or UO_971 (O_971,N_8384,N_6876);
or UO_972 (O_972,N_9661,N_5276);
nor UO_973 (O_973,N_6606,N_8416);
nor UO_974 (O_974,N_8419,N_7310);
nor UO_975 (O_975,N_8871,N_7592);
nand UO_976 (O_976,N_9747,N_5341);
or UO_977 (O_977,N_6263,N_9317);
nor UO_978 (O_978,N_6111,N_8500);
nor UO_979 (O_979,N_9130,N_7714);
nor UO_980 (O_980,N_6059,N_7457);
nor UO_981 (O_981,N_8652,N_5245);
nand UO_982 (O_982,N_8641,N_8987);
nor UO_983 (O_983,N_9998,N_7272);
or UO_984 (O_984,N_8920,N_9946);
and UO_985 (O_985,N_9892,N_8132);
or UO_986 (O_986,N_7278,N_8188);
nor UO_987 (O_987,N_6058,N_8753);
or UO_988 (O_988,N_6339,N_5853);
or UO_989 (O_989,N_8338,N_5844);
nand UO_990 (O_990,N_9290,N_6509);
or UO_991 (O_991,N_9372,N_5987);
nor UO_992 (O_992,N_9796,N_8695);
or UO_993 (O_993,N_9927,N_5881);
nor UO_994 (O_994,N_6698,N_5934);
or UO_995 (O_995,N_7319,N_7474);
or UO_996 (O_996,N_5922,N_9683);
and UO_997 (O_997,N_8979,N_8922);
nand UO_998 (O_998,N_9034,N_5748);
or UO_999 (O_999,N_5280,N_7166);
nor UO_1000 (O_1000,N_5040,N_6728);
or UO_1001 (O_1001,N_5409,N_9353);
or UO_1002 (O_1002,N_7515,N_6894);
nand UO_1003 (O_1003,N_9161,N_8112);
and UO_1004 (O_1004,N_7026,N_5735);
nor UO_1005 (O_1005,N_9040,N_6293);
and UO_1006 (O_1006,N_6103,N_7401);
or UO_1007 (O_1007,N_8346,N_6676);
xor UO_1008 (O_1008,N_9447,N_5093);
and UO_1009 (O_1009,N_8599,N_6520);
and UO_1010 (O_1010,N_7458,N_6109);
nand UO_1011 (O_1011,N_6911,N_6082);
nor UO_1012 (O_1012,N_7162,N_9907);
or UO_1013 (O_1013,N_8362,N_5967);
and UO_1014 (O_1014,N_6966,N_7598);
nor UO_1015 (O_1015,N_8114,N_6259);
and UO_1016 (O_1016,N_9366,N_9493);
and UO_1017 (O_1017,N_7103,N_7237);
and UO_1018 (O_1018,N_5466,N_8024);
or UO_1019 (O_1019,N_8220,N_5107);
nor UO_1020 (O_1020,N_9869,N_6757);
or UO_1021 (O_1021,N_8363,N_9148);
or UO_1022 (O_1022,N_9017,N_6422);
nand UO_1023 (O_1023,N_7771,N_9808);
nor UO_1024 (O_1024,N_9345,N_5410);
and UO_1025 (O_1025,N_9022,N_5054);
and UO_1026 (O_1026,N_7063,N_8195);
and UO_1027 (O_1027,N_8040,N_6549);
nand UO_1028 (O_1028,N_9411,N_8286);
or UO_1029 (O_1029,N_8916,N_7155);
nor UO_1030 (O_1030,N_8801,N_7697);
and UO_1031 (O_1031,N_7230,N_9870);
or UO_1032 (O_1032,N_5615,N_6236);
nor UO_1033 (O_1033,N_5668,N_9849);
and UO_1034 (O_1034,N_5397,N_6971);
and UO_1035 (O_1035,N_9433,N_8952);
nand UO_1036 (O_1036,N_9556,N_8680);
nor UO_1037 (O_1037,N_9326,N_5511);
and UO_1038 (O_1038,N_7833,N_6718);
nand UO_1039 (O_1039,N_6255,N_7077);
and UO_1040 (O_1040,N_7085,N_8410);
nand UO_1041 (O_1041,N_5981,N_7504);
or UO_1042 (O_1042,N_5549,N_6393);
nand UO_1043 (O_1043,N_6383,N_6198);
or UO_1044 (O_1044,N_8672,N_6458);
nor UO_1045 (O_1045,N_8675,N_7398);
nor UO_1046 (O_1046,N_8631,N_7073);
or UO_1047 (O_1047,N_5195,N_5018);
and UO_1048 (O_1048,N_9561,N_5420);
and UO_1049 (O_1049,N_8129,N_7777);
nand UO_1050 (O_1050,N_5800,N_9413);
and UO_1051 (O_1051,N_5131,N_7275);
or UO_1052 (O_1052,N_7329,N_8969);
or UO_1053 (O_1053,N_8430,N_5581);
and UO_1054 (O_1054,N_8566,N_7220);
nand UO_1055 (O_1055,N_7871,N_8345);
nand UO_1056 (O_1056,N_8222,N_5080);
nand UO_1057 (O_1057,N_7686,N_7842);
and UO_1058 (O_1058,N_6347,N_9176);
or UO_1059 (O_1059,N_7844,N_8282);
and UO_1060 (O_1060,N_5535,N_6374);
or UO_1061 (O_1061,N_9304,N_7104);
or UO_1062 (O_1062,N_9864,N_7753);
or UO_1063 (O_1063,N_6993,N_7134);
nand UO_1064 (O_1064,N_7766,N_7471);
and UO_1065 (O_1065,N_9832,N_5220);
nand UO_1066 (O_1066,N_9867,N_8837);
or UO_1067 (O_1067,N_6854,N_8377);
or UO_1068 (O_1068,N_8729,N_5657);
or UO_1069 (O_1069,N_8172,N_6634);
nand UO_1070 (O_1070,N_9270,N_8856);
and UO_1071 (O_1071,N_5789,N_9060);
and UO_1072 (O_1072,N_8945,N_8527);
or UO_1073 (O_1073,N_8131,N_5582);
or UO_1074 (O_1074,N_6048,N_9301);
nand UO_1075 (O_1075,N_5442,N_6330);
nand UO_1076 (O_1076,N_8666,N_9435);
and UO_1077 (O_1077,N_5256,N_5437);
and UO_1078 (O_1078,N_9872,N_9724);
or UO_1079 (O_1079,N_9704,N_5749);
and UO_1080 (O_1080,N_8287,N_8458);
nor UO_1081 (O_1081,N_5666,N_8872);
nand UO_1082 (O_1082,N_9420,N_5415);
nand UO_1083 (O_1083,N_6988,N_9056);
nand UO_1084 (O_1084,N_6408,N_7389);
nor UO_1085 (O_1085,N_6125,N_8307);
and UO_1086 (O_1086,N_5841,N_8843);
nand UO_1087 (O_1087,N_5219,N_6483);
and UO_1088 (O_1088,N_8139,N_8890);
and UO_1089 (O_1089,N_8529,N_5052);
nand UO_1090 (O_1090,N_9703,N_8673);
and UO_1091 (O_1091,N_8038,N_5681);
nand UO_1092 (O_1092,N_6762,N_8630);
or UO_1093 (O_1093,N_7277,N_7088);
and UO_1094 (O_1094,N_5169,N_6572);
or UO_1095 (O_1095,N_8768,N_8341);
and UO_1096 (O_1096,N_7878,N_5465);
nor UO_1097 (O_1097,N_7156,N_5422);
nor UO_1098 (O_1098,N_6543,N_9969);
nand UO_1099 (O_1099,N_9375,N_5092);
nand UO_1100 (O_1100,N_7597,N_7013);
nand UO_1101 (O_1101,N_7847,N_8457);
or UO_1102 (O_1102,N_8582,N_7318);
nand UO_1103 (O_1103,N_7480,N_8538);
and UO_1104 (O_1104,N_9432,N_8072);
nand UO_1105 (O_1105,N_6459,N_8522);
or UO_1106 (O_1106,N_5374,N_8047);
nand UO_1107 (O_1107,N_7745,N_5204);
and UO_1108 (O_1108,N_7296,N_9439);
or UO_1109 (O_1109,N_6394,N_7396);
nor UO_1110 (O_1110,N_5221,N_6369);
nor UO_1111 (O_1111,N_9829,N_7868);
nor UO_1112 (O_1112,N_8669,N_5732);
or UO_1113 (O_1113,N_5061,N_9616);
nor UO_1114 (O_1114,N_9627,N_7936);
nor UO_1115 (O_1115,N_6667,N_7460);
or UO_1116 (O_1116,N_9150,N_7254);
nand UO_1117 (O_1117,N_8197,N_8076);
nand UO_1118 (O_1118,N_6191,N_7653);
nand UO_1119 (O_1119,N_9862,N_6507);
and UO_1120 (O_1120,N_6738,N_9001);
or UO_1121 (O_1121,N_9673,N_8193);
nand UO_1122 (O_1122,N_7459,N_9109);
or UO_1123 (O_1123,N_9587,N_7349);
nor UO_1124 (O_1124,N_9780,N_8027);
nand UO_1125 (O_1125,N_9538,N_6177);
nor UO_1126 (O_1126,N_9445,N_6835);
or UO_1127 (O_1127,N_6605,N_7875);
nor UO_1128 (O_1128,N_9325,N_8758);
nor UO_1129 (O_1129,N_5835,N_5813);
nor UO_1130 (O_1130,N_8415,N_6546);
nor UO_1131 (O_1131,N_7114,N_8903);
nand UO_1132 (O_1132,N_8534,N_5608);
or UO_1133 (O_1133,N_7934,N_7874);
and UO_1134 (O_1134,N_5645,N_5603);
and UO_1135 (O_1135,N_7955,N_8106);
nand UO_1136 (O_1136,N_9665,N_6435);
or UO_1137 (O_1137,N_6108,N_5962);
nor UO_1138 (O_1138,N_5133,N_9468);
nor UO_1139 (O_1139,N_7673,N_8825);
or UO_1140 (O_1140,N_7012,N_8336);
or UO_1141 (O_1141,N_8092,N_6575);
nand UO_1142 (O_1142,N_9321,N_9874);
nor UO_1143 (O_1143,N_5118,N_6052);
or UO_1144 (O_1144,N_9922,N_6609);
nor UO_1145 (O_1145,N_5798,N_6870);
nand UO_1146 (O_1146,N_5578,N_5704);
nand UO_1147 (O_1147,N_9152,N_8543);
nor UO_1148 (O_1148,N_7828,N_8817);
and UO_1149 (O_1149,N_7060,N_7719);
nor UO_1150 (O_1150,N_6533,N_7938);
and UO_1151 (O_1151,N_8435,N_6811);
nor UO_1152 (O_1152,N_7960,N_7141);
nor UO_1153 (O_1153,N_8699,N_6092);
nor UO_1154 (O_1154,N_6095,N_6004);
nor UO_1155 (O_1155,N_5210,N_6113);
nand UO_1156 (O_1156,N_8732,N_5395);
nand UO_1157 (O_1157,N_6628,N_8250);
and UO_1158 (O_1158,N_6332,N_9884);
nor UO_1159 (O_1159,N_9486,N_6643);
and UO_1160 (O_1160,N_7637,N_9283);
or UO_1161 (O_1161,N_7917,N_9753);
nor UO_1162 (O_1162,N_9175,N_5314);
nand UO_1163 (O_1163,N_5419,N_6945);
nand UO_1164 (O_1164,N_6368,N_9206);
or UO_1165 (O_1165,N_8826,N_8301);
nand UO_1166 (O_1166,N_5258,N_9507);
nor UO_1167 (O_1167,N_5019,N_9379);
or UO_1168 (O_1168,N_5750,N_5780);
nand UO_1169 (O_1169,N_6829,N_8474);
nand UO_1170 (O_1170,N_6011,N_8881);
and UO_1171 (O_1171,N_6117,N_6613);
nor UO_1172 (O_1172,N_5829,N_5127);
and UO_1173 (O_1173,N_8480,N_5291);
nand UO_1174 (O_1174,N_8066,N_5970);
and UO_1175 (O_1175,N_6473,N_5435);
and UO_1176 (O_1176,N_5803,N_6886);
nand UO_1177 (O_1177,N_6786,N_8068);
nor UO_1178 (O_1178,N_6871,N_9789);
nor UO_1179 (O_1179,N_7948,N_8553);
or UO_1180 (O_1180,N_6156,N_9108);
xnor UO_1181 (O_1181,N_8592,N_5996);
nand UO_1182 (O_1182,N_9259,N_7658);
or UO_1183 (O_1183,N_8501,N_6099);
nor UO_1184 (O_1184,N_5231,N_6577);
or UO_1185 (O_1185,N_7795,N_8799);
and UO_1186 (O_1186,N_8298,N_7132);
nor UO_1187 (O_1187,N_5378,N_8181);
and UO_1188 (O_1188,N_8359,N_8056);
and UO_1189 (O_1189,N_6298,N_8616);
or UO_1190 (O_1190,N_8127,N_8398);
or UO_1191 (O_1191,N_9397,N_5653);
nor UO_1192 (O_1192,N_5148,N_8335);
or UO_1193 (O_1193,N_7584,N_6262);
and UO_1194 (O_1194,N_9615,N_6160);
and UO_1195 (O_1195,N_5055,N_9456);
or UO_1196 (O_1196,N_5783,N_5075);
and UO_1197 (O_1197,N_7074,N_6267);
nor UO_1198 (O_1198,N_9106,N_8547);
nand UO_1199 (O_1199,N_8949,N_7433);
nand UO_1200 (O_1200,N_7748,N_5914);
and UO_1201 (O_1201,N_9567,N_7362);
nor UO_1202 (O_1202,N_6496,N_5072);
nand UO_1203 (O_1203,N_7106,N_6203);
nand UO_1204 (O_1204,N_8493,N_8065);
nor UO_1205 (O_1205,N_8219,N_9053);
nor UO_1206 (O_1206,N_5175,N_7873);
nor UO_1207 (O_1207,N_7393,N_6406);
nor UO_1208 (O_1208,N_6943,N_6831);
nand UO_1209 (O_1209,N_6680,N_8819);
and UO_1210 (O_1210,N_8710,N_9465);
or UO_1211 (O_1211,N_5487,N_9739);
nor UO_1212 (O_1212,N_8575,N_9334);
or UO_1213 (O_1213,N_9237,N_6664);
nor UO_1214 (O_1214,N_7053,N_8770);
or UO_1215 (O_1215,N_5212,N_7475);
nor UO_1216 (O_1216,N_5961,N_9224);
and UO_1217 (O_1217,N_5392,N_5076);
nand UO_1218 (O_1218,N_8852,N_9415);
nor UO_1219 (O_1219,N_9741,N_8138);
nor UO_1220 (O_1220,N_6668,N_6139);
nor UO_1221 (O_1221,N_8149,N_6453);
and UO_1222 (O_1222,N_7331,N_9000);
or UO_1223 (O_1223,N_9991,N_5540);
or UO_1224 (O_1224,N_9610,N_9557);
and UO_1225 (O_1225,N_5147,N_9374);
or UO_1226 (O_1226,N_9670,N_6188);
and UO_1227 (O_1227,N_5839,N_6420);
and UO_1228 (O_1228,N_6391,N_7520);
or UO_1229 (O_1229,N_5433,N_9268);
and UO_1230 (O_1230,N_8646,N_9003);
or UO_1231 (O_1231,N_6573,N_7571);
nand UO_1232 (O_1232,N_5140,N_9901);
nor UO_1233 (O_1233,N_8385,N_5326);
and UO_1234 (O_1234,N_8365,N_9071);
or UO_1235 (O_1235,N_9611,N_5286);
and UO_1236 (O_1236,N_7641,N_8043);
and UO_1237 (O_1237,N_7735,N_5864);
nand UO_1238 (O_1238,N_5697,N_8080);
nor UO_1239 (O_1239,N_8797,N_5178);
and UO_1240 (O_1240,N_5382,N_9930);
and UO_1241 (O_1241,N_6646,N_6767);
or UO_1242 (O_1242,N_8103,N_5345);
nor UO_1243 (O_1243,N_7160,N_5446);
and UO_1244 (O_1244,N_6844,N_6360);
nor UO_1245 (O_1245,N_8441,N_7607);
nand UO_1246 (O_1246,N_8959,N_7692);
nand UO_1247 (O_1247,N_6697,N_9745);
xnor UO_1248 (O_1248,N_9686,N_5695);
and UO_1249 (O_1249,N_5607,N_8168);
and UO_1250 (O_1250,N_6278,N_9070);
nor UO_1251 (O_1251,N_6421,N_8313);
or UO_1252 (O_1252,N_5035,N_7675);
nand UO_1253 (O_1253,N_6991,N_9891);
and UO_1254 (O_1254,N_8953,N_8682);
and UO_1255 (O_1255,N_5385,N_5491);
and UO_1256 (O_1256,N_5590,N_6582);
nor UO_1257 (O_1257,N_9923,N_6249);
or UO_1258 (O_1258,N_9378,N_8707);
nand UO_1259 (O_1259,N_7062,N_5947);
or UO_1260 (O_1260,N_5991,N_5153);
or UO_1261 (O_1261,N_7170,N_8437);
and UO_1262 (O_1262,N_5234,N_6839);
nand UO_1263 (O_1263,N_7744,N_9883);
nand UO_1264 (O_1264,N_6890,N_8686);
nand UO_1265 (O_1265,N_7422,N_7311);
nor UO_1266 (O_1266,N_9649,N_9866);
nand UO_1267 (O_1267,N_8777,N_9358);
nor UO_1268 (O_1268,N_8994,N_6683);
nand UO_1269 (O_1269,N_5230,N_6550);
or UO_1270 (O_1270,N_7779,N_8886);
xnor UO_1271 (O_1271,N_5246,N_5188);
nor UO_1272 (O_1272,N_7535,N_7183);
and UO_1273 (O_1273,N_7567,N_8962);
nor UO_1274 (O_1274,N_8431,N_9303);
nand UO_1275 (O_1275,N_7518,N_6484);
or UO_1276 (O_1276,N_8370,N_8256);
nor UO_1277 (O_1277,N_9749,N_9726);
nor UO_1278 (O_1278,N_9142,N_6941);
nand UO_1279 (O_1279,N_5252,N_8304);
or UO_1280 (O_1280,N_6990,N_6384);
and UO_1281 (O_1281,N_6873,N_7499);
and UO_1282 (O_1282,N_8453,N_8974);
or UO_1283 (O_1283,N_6187,N_5056);
nor UO_1284 (O_1284,N_8515,N_8985);
and UO_1285 (O_1285,N_9203,N_9204);
nor UO_1286 (O_1286,N_9263,N_7348);
nand UO_1287 (O_1287,N_9644,N_9762);
nor UO_1288 (O_1288,N_9079,N_9058);
nor UO_1289 (O_1289,N_6969,N_7304);
nor UO_1290 (O_1290,N_5911,N_9138);
nor UO_1291 (O_1291,N_6364,N_9652);
or UO_1292 (O_1292,N_7838,N_8376);
nand UO_1293 (O_1293,N_5777,N_9986);
and UO_1294 (O_1294,N_6276,N_9819);
nand UO_1295 (O_1295,N_6480,N_8603);
or UO_1296 (O_1296,N_9227,N_5136);
nor UO_1297 (O_1297,N_7253,N_9223);
or UO_1298 (O_1298,N_8773,N_6272);
or UO_1299 (O_1299,N_8229,N_8328);
and UO_1300 (O_1300,N_6365,N_9293);
nor UO_1301 (O_1301,N_8999,N_9444);
nor UO_1302 (O_1302,N_5149,N_7737);
and UO_1303 (O_1303,N_7561,N_6225);
and UO_1304 (O_1304,N_6889,N_7681);
nand UO_1305 (O_1305,N_5759,N_5353);
nand UO_1306 (O_1306,N_5110,N_9997);
or UO_1307 (O_1307,N_5574,N_7082);
nor UO_1308 (O_1308,N_8413,N_5588);
nand UO_1309 (O_1309,N_9727,N_7435);
nand UO_1310 (O_1310,N_9425,N_8007);
or UO_1311 (O_1311,N_8804,N_7248);
nand UO_1312 (O_1312,N_5564,N_9926);
nand UO_1313 (O_1313,N_6143,N_9919);
and UO_1314 (O_1314,N_7295,N_9527);
xnor UO_1315 (O_1315,N_9166,N_5334);
xnor UO_1316 (O_1316,N_8122,N_6413);
or UO_1317 (O_1317,N_5413,N_8300);
nor UO_1318 (O_1318,N_8090,N_9500);
nor UO_1319 (O_1319,N_5688,N_7791);
nand UO_1320 (O_1320,N_7345,N_8233);
or UO_1321 (O_1321,N_7338,N_6080);
nor UO_1322 (O_1322,N_6722,N_8240);
nand UO_1323 (O_1323,N_7369,N_5137);
xor UO_1324 (O_1324,N_7730,N_7923);
nand UO_1325 (O_1325,N_7223,N_6833);
nor UO_1326 (O_1326,N_7045,N_6404);
nand UO_1327 (O_1327,N_7015,N_8908);
and UO_1328 (O_1328,N_5370,N_7283);
or UO_1329 (O_1329,N_8270,N_9551);
nand UO_1330 (O_1330,N_7816,N_7531);
and UO_1331 (O_1331,N_6939,N_9737);
nand UO_1332 (O_1332,N_6816,N_9548);
or UO_1333 (O_1333,N_5517,N_6296);
and UO_1334 (O_1334,N_6514,N_9599);
or UO_1335 (O_1335,N_6684,N_8425);
or UO_1336 (O_1336,N_8573,N_9952);
nor UO_1337 (O_1337,N_5281,N_5401);
and UO_1338 (O_1338,N_7221,N_9505);
or UO_1339 (O_1339,N_5888,N_7634);
and UO_1340 (O_1340,N_5375,N_9208);
nor UO_1341 (O_1341,N_7715,N_7722);
nand UO_1342 (O_1342,N_5573,N_8909);
or UO_1343 (O_1343,N_5311,N_9805);
nand UO_1344 (O_1344,N_5387,N_9988);
nand UO_1345 (O_1345,N_9442,N_8964);
or UO_1346 (O_1346,N_5320,N_5418);
nor UO_1347 (O_1347,N_7260,N_9024);
nor UO_1348 (O_1348,N_5946,N_6955);
nand UO_1349 (O_1349,N_6382,N_8337);
or UO_1350 (O_1350,N_6893,N_7151);
or UO_1351 (O_1351,N_5151,N_9730);
nor UO_1352 (O_1352,N_5095,N_5068);
and UO_1353 (O_1353,N_9384,N_5105);
and UO_1354 (O_1354,N_7325,N_9968);
nor UO_1355 (O_1355,N_5930,N_6340);
and UO_1356 (O_1356,N_8787,N_9531);
nor UO_1357 (O_1357,N_8840,N_6852);
or UO_1358 (O_1358,N_7072,N_5630);
nor UO_1359 (O_1359,N_5166,N_6290);
and UO_1360 (O_1360,N_8142,N_7773);
and UO_1361 (O_1361,N_8089,N_7689);
nand UO_1362 (O_1362,N_5980,N_7834);
or UO_1363 (O_1363,N_9392,N_6361);
and UO_1364 (O_1364,N_9350,N_7512);
nand UO_1365 (O_1365,N_7371,N_9850);
and UO_1366 (O_1366,N_5114,N_6885);
nor UO_1367 (O_1367,N_7265,N_7245);
nor UO_1368 (O_1368,N_7343,N_8285);
nor UO_1369 (O_1369,N_5335,N_5632);
or UO_1370 (O_1370,N_6454,N_9909);
nor UO_1371 (O_1371,N_8115,N_8135);
and UO_1372 (O_1372,N_9783,N_5164);
and UO_1373 (O_1373,N_6009,N_8433);
nor UO_1374 (O_1374,N_9179,N_9622);
nand UO_1375 (O_1375,N_6810,N_8180);
nand UO_1376 (O_1376,N_9113,N_5046);
nand UO_1377 (O_1377,N_8951,N_5965);
nand UO_1378 (O_1378,N_6774,N_8049);
or UO_1379 (O_1379,N_6342,N_5152);
and UO_1380 (O_1380,N_6498,N_6037);
or UO_1381 (O_1381,N_8387,N_7775);
nor UO_1382 (O_1382,N_7940,N_8757);
or UO_1383 (O_1383,N_5173,N_6056);
and UO_1384 (O_1384,N_5891,N_7497);
nor UO_1385 (O_1385,N_8182,N_8194);
nor UO_1386 (O_1386,N_5505,N_6069);
nor UO_1387 (O_1387,N_5589,N_5663);
or UO_1388 (O_1388,N_5542,N_6152);
and UO_1389 (O_1389,N_9541,N_6337);
and UO_1390 (O_1390,N_6848,N_5840);
xor UO_1391 (O_1391,N_9107,N_5224);
nor UO_1392 (O_1392,N_6518,N_5807);
nand UO_1393 (O_1393,N_7128,N_7268);
nor UO_1394 (O_1394,N_8917,N_8851);
or UO_1395 (O_1395,N_6777,N_6862);
nor UO_1396 (O_1396,N_6569,N_8225);
or UO_1397 (O_1397,N_8793,N_8011);
or UO_1398 (O_1398,N_9956,N_9205);
or UO_1399 (O_1399,N_5044,N_9516);
nand UO_1400 (O_1400,N_5998,N_8403);
xnor UO_1401 (O_1401,N_6295,N_7781);
nor UO_1402 (O_1402,N_9877,N_9059);
or UO_1403 (O_1403,N_7902,N_5825);
nand UO_1404 (O_1404,N_5490,N_5227);
nand UO_1405 (O_1405,N_7583,N_9105);
or UO_1406 (O_1406,N_6912,N_7491);
and UO_1407 (O_1407,N_7347,N_9696);
nand UO_1408 (O_1408,N_9873,N_9967);
nand UO_1409 (O_1409,N_6649,N_9676);
or UO_1410 (O_1410,N_7264,N_6089);
nor UO_1411 (O_1411,N_9699,N_8898);
nand UO_1412 (O_1412,N_5694,N_8806);
or UO_1413 (O_1413,N_9979,N_6856);
nor UO_1414 (O_1414,N_6978,N_9019);
or UO_1415 (O_1415,N_7651,N_6158);
nor UO_1416 (O_1416,N_5458,N_5155);
nand UO_1417 (O_1417,N_7079,N_5015);
or UO_1418 (O_1418,N_9642,N_5488);
nand UO_1419 (O_1419,N_5372,N_9624);
nand UO_1420 (O_1420,N_5912,N_6373);
and UO_1421 (O_1421,N_5363,N_8100);
nand UO_1422 (O_1422,N_9641,N_5322);
nor UO_1423 (O_1423,N_7596,N_8357);
xnor UO_1424 (O_1424,N_6410,N_9886);
and UO_1425 (O_1425,N_7639,N_7534);
nor UO_1426 (O_1426,N_8706,N_6653);
or UO_1427 (O_1427,N_6322,N_8261);
nor UO_1428 (O_1428,N_8461,N_8438);
xnor UO_1429 (O_1429,N_8568,N_9813);
nor UO_1430 (O_1430,N_5371,N_6934);
nor UO_1431 (O_1431,N_7933,N_8598);
and UO_1432 (O_1432,N_6805,N_6217);
nand UO_1433 (O_1433,N_6655,N_6797);
nand UO_1434 (O_1434,N_8776,N_5902);
nand UO_1435 (O_1435,N_6557,N_7424);
nand UO_1436 (O_1436,N_7442,N_9804);
and UO_1437 (O_1437,N_6401,N_6341);
and UO_1438 (O_1438,N_6923,N_5831);
and UO_1439 (O_1439,N_7611,N_5817);
and UO_1440 (O_1440,N_7578,N_8191);
nor UO_1441 (O_1441,N_8684,N_5432);
and UO_1442 (O_1442,N_9240,N_5461);
nor UO_1443 (O_1443,N_7964,N_5186);
and UO_1444 (O_1444,N_6397,N_7588);
nand UO_1445 (O_1445,N_9357,N_7328);
or UO_1446 (O_1446,N_9104,N_8454);
and UO_1447 (O_1447,N_7032,N_7397);
xor UO_1448 (O_1448,N_6563,N_6763);
and UO_1449 (O_1449,N_8266,N_8151);
and UO_1450 (O_1450,N_8126,N_9962);
and UO_1451 (O_1451,N_8254,N_6621);
and UO_1452 (O_1452,N_8053,N_9544);
or UO_1453 (O_1453,N_5172,N_5986);
nor UO_1454 (O_1454,N_5331,N_8606);
and UO_1455 (O_1455,N_9013,N_9563);
nor UO_1456 (O_1456,N_5696,N_9165);
and UO_1457 (O_1457,N_8560,N_5091);
or UO_1458 (O_1458,N_6321,N_9520);
nand UO_1459 (O_1459,N_8019,N_7469);
or UO_1460 (O_1460,N_8993,N_6967);
nand UO_1461 (O_1461,N_7351,N_9265);
nand UO_1462 (O_1462,N_6641,N_7479);
nor UO_1463 (O_1463,N_9207,N_6104);
nand UO_1464 (O_1464,N_5602,N_6162);
xor UO_1465 (O_1465,N_5937,N_9457);
nor UO_1466 (O_1466,N_9845,N_7699);
nand UO_1467 (O_1467,N_5819,N_6190);
or UO_1468 (O_1468,N_7882,N_7818);
nand UO_1469 (O_1469,N_7488,N_9102);
nand UO_1470 (O_1470,N_5583,N_6072);
nand UO_1471 (O_1471,N_9289,N_6001);
nand UO_1472 (O_1472,N_6326,N_9833);
and UO_1473 (O_1473,N_6455,N_7188);
nor UO_1474 (O_1474,N_6564,N_6842);
nand UO_1475 (O_1475,N_6469,N_5605);
nand UO_1476 (O_1476,N_8108,N_6957);
or UO_1477 (O_1477,N_6067,N_6612);
nor UO_1478 (O_1478,N_5836,N_9999);
nor UO_1479 (O_1479,N_7701,N_5635);
and UO_1480 (O_1480,N_8087,N_7586);
nor UO_1481 (O_1481,N_9971,N_5743);
nor UO_1482 (O_1482,N_9314,N_8565);
nor UO_1483 (O_1483,N_8046,N_6972);
and UO_1484 (O_1484,N_7516,N_5012);
and UO_1485 (O_1485,N_6764,N_9835);
nor UO_1486 (O_1486,N_9939,N_7217);
or UO_1487 (O_1487,N_8789,N_5337);
or UO_1488 (O_1488,N_5460,N_7712);
or UO_1489 (O_1489,N_8627,N_5390);
and UO_1490 (O_1490,N_7384,N_6984);
nand UO_1491 (O_1491,N_5381,N_6696);
and UO_1492 (O_1492,N_9685,N_5622);
and UO_1493 (O_1493,N_7091,N_5773);
nand UO_1494 (O_1494,N_7989,N_6378);
and UO_1495 (O_1495,N_7652,N_5323);
nor UO_1496 (O_1496,N_5145,N_7363);
nor UO_1497 (O_1497,N_9989,N_6415);
nand UO_1498 (O_1498,N_9603,N_9048);
xor UO_1499 (O_1499,N_6723,N_6530);
endmodule