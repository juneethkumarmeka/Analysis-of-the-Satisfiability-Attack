module basic_2000_20000_2500_20_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_871,In_1152);
xnor U1 (N_1,In_337,In_1122);
nor U2 (N_2,In_720,In_1178);
or U3 (N_3,In_1984,In_1309);
nor U4 (N_4,In_1431,In_1357);
nand U5 (N_5,In_339,In_783);
nand U6 (N_6,In_1366,In_960);
nand U7 (N_7,In_121,In_130);
or U8 (N_8,In_1823,In_886);
or U9 (N_9,In_425,In_921);
and U10 (N_10,In_110,In_1145);
or U11 (N_11,In_380,In_142);
and U12 (N_12,In_1260,In_1627);
xnor U13 (N_13,In_598,In_421);
nand U14 (N_14,In_325,In_1662);
or U15 (N_15,In_997,In_646);
or U16 (N_16,In_296,In_771);
nor U17 (N_17,In_1926,In_969);
xor U18 (N_18,In_1384,In_965);
nor U19 (N_19,In_1598,In_503);
and U20 (N_20,In_1115,In_1861);
or U21 (N_21,In_1890,In_1103);
and U22 (N_22,In_1585,In_849);
or U23 (N_23,In_111,In_90);
nand U24 (N_24,In_256,In_97);
and U25 (N_25,In_186,In_1077);
and U26 (N_26,In_957,In_76);
xor U27 (N_27,In_232,In_281);
nor U28 (N_28,In_1482,In_1395);
nand U29 (N_29,In_429,In_1347);
or U30 (N_30,In_1193,In_1614);
xnor U31 (N_31,In_1076,In_1953);
and U32 (N_32,In_485,In_1821);
and U33 (N_33,In_1459,In_1110);
or U34 (N_34,In_373,In_239);
nor U35 (N_35,In_363,In_1072);
xor U36 (N_36,In_740,In_1487);
nor U37 (N_37,In_623,In_192);
nand U38 (N_38,In_948,In_1742);
nor U39 (N_39,In_1223,In_1949);
xor U40 (N_40,In_1078,In_439);
and U41 (N_41,In_496,In_619);
nor U42 (N_42,In_57,In_1736);
nor U43 (N_43,In_1827,In_1690);
nor U44 (N_44,In_1005,In_126);
or U45 (N_45,In_1430,In_565);
or U46 (N_46,In_1967,In_1399);
nand U47 (N_47,In_1945,In_1878);
xor U48 (N_48,In_357,In_741);
and U49 (N_49,In_1262,In_932);
xnor U50 (N_50,In_787,In_92);
nand U51 (N_51,In_1432,In_758);
xnor U52 (N_52,In_1571,In_1270);
or U53 (N_53,In_1128,In_884);
xnor U54 (N_54,In_1481,In_198);
nand U55 (N_55,In_1304,In_665);
or U56 (N_56,In_647,In_1906);
or U57 (N_57,In_149,In_340);
or U58 (N_58,In_288,In_78);
xor U59 (N_59,In_345,In_1768);
and U60 (N_60,In_1891,In_1386);
xor U61 (N_61,In_958,In_467);
nor U62 (N_62,In_1909,In_904);
nand U63 (N_63,In_74,In_591);
xnor U64 (N_64,In_738,In_1718);
nand U65 (N_65,In_1401,In_508);
and U66 (N_66,In_768,In_1424);
nor U67 (N_67,In_767,In_581);
xnor U68 (N_68,In_1328,In_1126);
nand U69 (N_69,In_99,In_453);
nor U70 (N_70,In_642,In_1669);
and U71 (N_71,In_1325,In_1066);
and U72 (N_72,In_786,In_653);
nor U73 (N_73,In_1879,In_988);
and U74 (N_74,In_1605,In_1123);
nor U75 (N_75,In_1899,In_54);
or U76 (N_76,In_1000,In_926);
and U77 (N_77,In_788,In_689);
xnor U78 (N_78,In_67,In_1830);
nand U79 (N_79,In_11,In_1781);
nand U80 (N_80,In_1526,In_1215);
nand U81 (N_81,In_1296,In_1188);
xnor U82 (N_82,In_796,In_329);
and U83 (N_83,In_354,In_971);
nand U84 (N_84,In_275,In_1352);
nand U85 (N_85,In_167,In_637);
and U86 (N_86,In_301,In_427);
or U87 (N_87,In_1261,In_802);
nand U88 (N_88,In_1974,In_1786);
or U89 (N_89,In_136,In_91);
and U90 (N_90,In_1514,In_1449);
nor U91 (N_91,In_567,In_1273);
xnor U92 (N_92,In_657,In_199);
xnor U93 (N_93,In_1250,In_1803);
xnor U94 (N_94,In_1338,In_319);
or U95 (N_95,In_1914,In_1872);
nor U96 (N_96,In_1554,In_434);
nor U97 (N_97,In_1367,In_1682);
xnor U98 (N_98,In_910,In_853);
or U99 (N_99,In_1111,In_326);
and U100 (N_100,In_1628,In_1124);
xor U101 (N_101,In_708,In_1621);
nor U102 (N_102,In_322,In_152);
nand U103 (N_103,In_205,In_974);
or U104 (N_104,In_1797,In_596);
xor U105 (N_105,In_1944,In_519);
nand U106 (N_106,In_1980,In_473);
and U107 (N_107,In_701,In_1715);
or U108 (N_108,In_1054,In_1794);
nand U109 (N_109,In_1871,In_518);
nor U110 (N_110,In_710,In_1420);
nand U111 (N_111,In_170,In_1219);
xor U112 (N_112,In_45,In_1254);
and U113 (N_113,In_277,In_324);
nor U114 (N_114,In_38,In_1991);
or U115 (N_115,In_1600,In_1784);
or U116 (N_116,In_1677,In_1711);
nor U117 (N_117,In_1074,In_29);
nand U118 (N_118,In_552,In_1168);
xnor U119 (N_119,In_542,In_430);
or U120 (N_120,In_832,In_1575);
or U121 (N_121,In_1772,In_548);
nand U122 (N_122,In_407,In_562);
and U123 (N_123,In_108,In_1770);
and U124 (N_124,In_1735,In_1440);
and U125 (N_125,In_1313,In_1038);
or U126 (N_126,In_1229,In_1957);
and U127 (N_127,In_493,In_1622);
or U128 (N_128,In_1032,In_1593);
nand U129 (N_129,In_1933,In_1720);
and U130 (N_130,In_487,In_331);
and U131 (N_131,In_1160,In_1969);
nand U132 (N_132,In_176,In_1568);
and U133 (N_133,In_475,In_208);
nand U134 (N_134,In_1486,In_763);
nand U135 (N_135,In_1192,In_1195);
nand U136 (N_136,In_160,In_469);
nor U137 (N_137,In_987,In_1064);
or U138 (N_138,In_1322,In_1277);
and U139 (N_139,In_3,In_94);
nor U140 (N_140,In_481,In_1492);
or U141 (N_141,In_1134,In_235);
xor U142 (N_142,In_1358,In_1700);
and U143 (N_143,In_865,In_1379);
nor U144 (N_144,In_1257,In_914);
and U145 (N_145,In_1107,In_1056);
or U146 (N_146,In_317,In_309);
and U147 (N_147,In_401,In_697);
and U148 (N_148,In_1016,In_100);
and U149 (N_149,In_633,In_1138);
and U150 (N_150,In_1439,In_1917);
and U151 (N_151,In_1127,In_1302);
or U152 (N_152,In_1147,In_1370);
and U153 (N_153,In_1214,In_1374);
xnor U154 (N_154,In_302,In_463);
nand U155 (N_155,In_1810,In_951);
nand U156 (N_156,In_944,In_1024);
and U157 (N_157,In_101,In_330);
nor U158 (N_158,In_193,In_521);
xor U159 (N_159,In_563,In_30);
nand U160 (N_160,In_1567,In_1536);
nand U161 (N_161,In_1052,In_1491);
xnor U162 (N_162,In_1509,In_1198);
nand U163 (N_163,In_1125,In_773);
xor U164 (N_164,In_1566,In_1221);
nor U165 (N_165,In_824,In_1351);
xor U166 (N_166,In_594,In_1992);
nor U167 (N_167,In_715,In_776);
or U168 (N_168,In_1971,In_875);
or U169 (N_169,In_1708,In_743);
nor U170 (N_170,In_972,In_1534);
or U171 (N_171,In_1692,In_812);
xnor U172 (N_172,In_1684,In_995);
and U173 (N_173,In_1565,In_9);
and U174 (N_174,In_724,In_1817);
xnor U175 (N_175,In_754,In_1913);
nand U176 (N_176,In_1606,In_1400);
nor U177 (N_177,In_800,In_959);
xnor U178 (N_178,In_1256,In_1990);
and U179 (N_179,In_723,In_88);
or U180 (N_180,In_305,In_1396);
and U181 (N_181,In_1892,In_440);
and U182 (N_182,In_1930,In_1441);
xnor U183 (N_183,In_1101,In_1083);
nor U184 (N_184,In_902,In_1978);
nor U185 (N_185,In_1502,In_350);
xnor U186 (N_186,In_424,In_885);
xnor U187 (N_187,In_792,In_864);
nor U188 (N_188,In_640,In_1939);
xor U189 (N_189,In_1630,In_169);
or U190 (N_190,In_841,In_1665);
or U191 (N_191,In_1312,In_706);
and U192 (N_192,In_1182,In_1364);
or U193 (N_193,In_1757,In_1246);
xnor U194 (N_194,In_1924,In_712);
or U195 (N_195,In_652,In_1552);
and U196 (N_196,In_1017,In_231);
nand U197 (N_197,In_1158,In_1888);
nor U198 (N_198,In_1993,In_1513);
or U199 (N_199,In_246,In_1850);
xor U200 (N_200,In_1047,In_43);
nor U201 (N_201,In_491,In_1640);
or U202 (N_202,In_442,In_436);
xnor U203 (N_203,In_1874,In_541);
nor U204 (N_204,In_1478,In_308);
and U205 (N_205,In_1135,In_946);
nand U206 (N_206,In_85,In_747);
or U207 (N_207,In_1883,In_1995);
or U208 (N_208,In_202,In_549);
or U209 (N_209,In_150,In_799);
nor U210 (N_210,In_273,In_10);
xnor U211 (N_211,In_1964,In_1558);
nor U212 (N_212,In_64,In_1404);
and U213 (N_213,In_778,In_255);
nand U214 (N_214,In_1716,In_1959);
xnor U215 (N_215,In_685,In_227);
and U216 (N_216,In_785,In_1271);
or U217 (N_217,In_347,In_1972);
or U218 (N_218,In_166,In_274);
and U219 (N_219,In_365,In_1553);
nand U220 (N_220,In_1336,In_1376);
xnor U221 (N_221,In_1864,In_20);
nand U222 (N_222,In_46,In_782);
or U223 (N_223,In_887,In_1207);
or U224 (N_224,In_37,In_410);
nor U225 (N_225,In_70,In_1848);
or U226 (N_226,In_1087,In_810);
or U227 (N_227,In_757,In_1782);
and U228 (N_228,In_1638,In_1564);
and U229 (N_229,In_1189,In_62);
xor U230 (N_230,In_1977,In_1932);
and U231 (N_231,In_1822,In_733);
or U232 (N_232,In_825,In_716);
nand U233 (N_233,In_206,In_1201);
xor U234 (N_234,In_1745,In_1480);
nand U235 (N_235,In_203,In_1410);
nor U236 (N_236,In_379,In_1806);
and U237 (N_237,In_300,In_543);
nor U238 (N_238,In_1239,In_265);
xnor U239 (N_239,In_691,In_795);
and U240 (N_240,In_1460,In_1865);
nor U241 (N_241,In_1798,In_1761);
and U242 (N_242,In_862,In_1279);
nor U243 (N_243,In_1783,In_1092);
nor U244 (N_244,In_1003,In_1412);
nor U245 (N_245,In_1472,In_1753);
xnor U246 (N_246,In_1751,In_1582);
nand U247 (N_247,In_1734,In_1928);
and U248 (N_248,In_1973,In_1738);
or U249 (N_249,In_953,In_1590);
or U250 (N_250,In_831,In_1356);
and U251 (N_251,In_1834,In_1766);
nor U252 (N_252,In_994,In_16);
and U253 (N_253,In_403,In_1710);
nor U254 (N_254,In_1855,In_1646);
nor U255 (N_255,In_781,In_1961);
and U256 (N_256,In_1197,In_1369);
xor U257 (N_257,In_266,In_730);
nand U258 (N_258,In_1916,In_963);
nor U259 (N_259,In_901,In_1584);
nor U260 (N_260,In_806,In_31);
or U261 (N_261,In_532,In_574);
and U262 (N_262,In_667,In_870);
or U263 (N_263,In_1512,In_1330);
and U264 (N_264,In_1267,In_278);
nor U265 (N_265,In_1905,In_448);
nand U266 (N_266,In_394,In_13);
or U267 (N_267,In_1704,In_1516);
or U268 (N_268,In_1471,In_1657);
nand U269 (N_269,In_1556,In_515);
nand U270 (N_270,In_506,In_343);
nand U271 (N_271,In_1880,In_1998);
nand U272 (N_272,In_1694,In_1611);
xnor U273 (N_273,In_1175,In_1307);
or U274 (N_274,In_1316,In_1332);
xnor U275 (N_275,In_1896,In_973);
nand U276 (N_276,In_961,In_236);
nor U277 (N_277,In_1272,In_414);
xor U278 (N_278,In_608,In_112);
and U279 (N_279,In_1762,In_1212);
xor U280 (N_280,In_1130,In_669);
nand U281 (N_281,In_1679,In_505);
nor U282 (N_282,In_774,In_1457);
or U283 (N_283,In_1299,In_1579);
and U284 (N_284,In_1820,In_61);
and U285 (N_285,In_923,In_107);
xor U286 (N_286,In_839,In_614);
and U287 (N_287,In_1845,In_1402);
or U288 (N_288,In_1161,In_607);
nand U289 (N_289,In_1688,In_876);
and U290 (N_290,In_1222,In_1597);
xor U291 (N_291,In_1194,In_1927);
xor U292 (N_292,In_270,In_497);
or U293 (N_293,In_513,In_1284);
nor U294 (N_294,In_1444,In_163);
and U295 (N_295,In_299,In_307);
nand U296 (N_296,In_1349,In_1686);
and U297 (N_297,In_935,In_1075);
nor U298 (N_298,In_1142,In_547);
xor U299 (N_299,In_1970,In_1520);
nand U300 (N_300,In_1721,In_420);
nand U301 (N_301,In_670,In_892);
or U302 (N_302,In_1873,In_1608);
xnor U303 (N_303,In_867,In_1859);
or U304 (N_304,In_1758,In_63);
nand U305 (N_305,In_1372,In_1904);
or U306 (N_306,In_272,In_157);
nor U307 (N_307,In_51,In_284);
nand U308 (N_308,In_113,In_1421);
or U309 (N_309,In_82,In_1278);
and U310 (N_310,In_528,In_609);
and U311 (N_311,In_671,In_151);
or U312 (N_312,In_1533,In_1238);
and U313 (N_313,In_285,In_861);
nor U314 (N_314,In_344,In_1088);
nor U315 (N_315,In_445,In_630);
or U316 (N_316,In_53,In_753);
xnor U317 (N_317,In_1581,In_1141);
or U318 (N_318,In_750,In_282);
xor U319 (N_319,In_675,In_144);
nor U320 (N_320,In_1096,In_1754);
or U321 (N_321,In_1368,In_807);
or U322 (N_322,In_1521,In_1414);
xnor U323 (N_323,In_73,In_531);
nor U324 (N_324,In_1765,In_1609);
nand U325 (N_325,In_1732,In_650);
or U326 (N_326,In_1922,In_805);
and U327 (N_327,In_295,In_1759);
nand U328 (N_328,In_539,In_1151);
nor U329 (N_329,In_341,In_1792);
or U330 (N_330,In_749,In_1954);
and U331 (N_331,In_955,In_949);
or U332 (N_332,In_334,In_60);
xnor U333 (N_333,In_1018,In_472);
xor U334 (N_334,In_1086,In_1388);
and U335 (N_335,In_1706,In_184);
nor U336 (N_336,In_120,In_1663);
or U337 (N_337,In_1829,In_1601);
nor U338 (N_338,In_544,In_1363);
nand U339 (N_339,In_311,In_1795);
or U340 (N_340,In_851,In_1729);
nand U341 (N_341,In_1339,In_1997);
xnor U342 (N_342,In_576,In_1854);
and U343 (N_343,In_352,In_687);
nor U344 (N_344,In_1132,In_899);
nor U345 (N_345,In_558,In_1539);
xnor U346 (N_346,In_1907,In_920);
and U347 (N_347,In_1031,In_1220);
nor U348 (N_348,In_551,In_1683);
nand U349 (N_349,In_87,In_1867);
nand U350 (N_350,In_1498,In_358);
nand U351 (N_351,In_1697,In_1001);
xor U352 (N_352,In_599,In_755);
or U353 (N_353,In_1436,In_889);
nand U354 (N_354,In_1228,In_72);
nand U355 (N_355,In_1994,In_522);
nor U356 (N_356,In_1607,In_1171);
or U357 (N_357,In_674,In_1140);
or U358 (N_358,In_592,In_952);
nand U359 (N_359,In_1411,In_931);
xnor U360 (N_360,In_446,In_699);
nor U361 (N_361,In_1375,In_245);
xor U362 (N_362,In_187,In_1519);
or U363 (N_363,In_1023,In_1285);
and U364 (N_364,In_182,In_1595);
xnor U365 (N_365,In_385,In_1106);
and U366 (N_366,In_499,In_1730);
nand U367 (N_367,In_1204,In_911);
xnor U368 (N_368,In_1658,In_535);
nand U369 (N_369,In_140,In_1676);
nand U370 (N_370,In_1099,In_840);
and U371 (N_371,In_1026,In_1020);
nor U372 (N_372,In_229,In_976);
or U373 (N_373,In_84,In_617);
nor U374 (N_374,In_79,In_27);
and U375 (N_375,In_226,In_925);
nor U376 (N_376,In_254,In_433);
or U377 (N_377,In_573,In_1976);
or U378 (N_378,In_537,In_1965);
or U379 (N_379,In_353,In_1244);
nor U380 (N_380,In_924,In_791);
or U381 (N_381,In_984,In_622);
nor U382 (N_382,In_1853,In_1011);
nor U383 (N_383,In_1046,In_748);
nand U384 (N_384,In_779,In_593);
xnor U385 (N_385,In_216,In_483);
nand U386 (N_386,In_438,In_486);
or U387 (N_387,In_1517,In_1529);
nor U388 (N_388,In_1165,In_1470);
xnor U389 (N_389,In_982,In_1723);
or U390 (N_390,In_1982,In_1860);
and U391 (N_391,In_826,In_1505);
xor U392 (N_392,In_183,In_577);
or U393 (N_393,In_816,In_1852);
or U394 (N_394,In_1184,In_915);
xor U395 (N_395,In_1423,In_507);
and U396 (N_396,In_1722,In_249);
or U397 (N_397,In_1461,In_377);
and U398 (N_398,In_1213,In_1602);
and U399 (N_399,In_588,In_196);
nand U400 (N_400,In_1469,In_837);
nor U401 (N_401,In_1826,In_1474);
nand U402 (N_402,In_252,In_415);
nor U403 (N_403,In_1545,In_222);
nand U404 (N_404,In_1719,In_956);
and U405 (N_405,In_703,In_1172);
xor U406 (N_406,In_1345,In_803);
xnor U407 (N_407,In_1588,In_1709);
xnor U408 (N_408,In_1068,In_766);
or U409 (N_409,In_704,In_798);
or U410 (N_410,In_843,In_1170);
or U411 (N_411,In_1079,In_854);
xnor U412 (N_412,In_1095,In_1191);
xor U413 (N_413,In_1029,In_941);
nand U414 (N_414,In_134,In_751);
nor U415 (N_415,In_681,In_314);
xor U416 (N_416,In_303,In_555);
xnor U417 (N_417,In_1043,In_315);
or U418 (N_418,In_584,In_1360);
and U419 (N_419,In_1381,In_1527);
nor U420 (N_420,In_1615,In_595);
and U421 (N_421,In_1416,In_1986);
and U422 (N_422,In_1265,In_34);
or U423 (N_423,In_185,In_1217);
xor U424 (N_424,In_1196,In_1442);
and U425 (N_425,In_1583,In_1780);
and U426 (N_426,In_1202,In_1877);
xor U427 (N_427,In_628,In_680);
nand U428 (N_428,In_734,In_1731);
nor U429 (N_429,In_65,In_370);
nor U430 (N_430,In_1809,In_852);
and U431 (N_431,In_672,In_1484);
nor U432 (N_432,In_1561,In_280);
xor U433 (N_433,In_1743,In_210);
nor U434 (N_434,In_1053,In_668);
or U435 (N_435,In_550,In_204);
nor U436 (N_436,In_676,In_1249);
xnor U437 (N_437,In_1210,In_1240);
xor U438 (N_438,In_1531,In_1090);
xor U439 (N_439,In_408,In_732);
nor U440 (N_440,In_989,In_1572);
xnor U441 (N_441,In_1702,In_626);
xor U442 (N_442,In_906,In_649);
nand U443 (N_443,In_1462,In_937);
or U444 (N_444,In_772,In_2);
and U445 (N_445,In_742,In_1070);
xnor U446 (N_446,In_39,In_1174);
and U447 (N_447,In_1577,In_664);
nand U448 (N_448,In_1286,In_639);
xor U449 (N_449,In_1091,In_690);
nor U450 (N_450,In_1645,In_139);
nand U451 (N_451,In_700,In_225);
nor U452 (N_452,In_1144,In_375);
or U453 (N_453,In_606,In_1183);
xor U454 (N_454,In_1633,In_289);
or U455 (N_455,In_1799,In_1979);
nor U456 (N_456,In_26,In_1574);
nand U457 (N_457,In_488,In_1812);
xor U458 (N_458,In_1185,In_1503);
or U459 (N_459,In_897,In_1985);
or U460 (N_460,In_128,In_36);
and U461 (N_461,In_679,In_1061);
and U462 (N_462,In_1340,In_570);
xnor U463 (N_463,In_1488,In_692);
xor U464 (N_464,In_1825,In_1551);
nor U465 (N_465,In_376,In_1387);
nand U466 (N_466,In_1308,In_1073);
or U467 (N_467,In_1452,In_1084);
and U468 (N_468,In_1464,In_1785);
and U469 (N_469,In_287,In_1724);
xnor U470 (N_470,In_1789,In_1310);
nand U471 (N_471,In_355,In_817);
nand U472 (N_472,In_1055,In_1705);
and U473 (N_473,In_1557,In_98);
and U474 (N_474,In_1080,In_1294);
nor U475 (N_475,In_660,In_1319);
xnor U476 (N_476,In_809,In_999);
and U477 (N_477,In_580,In_1245);
and U478 (N_478,In_1739,In_1912);
and U479 (N_479,In_371,In_1477);
xor U480 (N_480,In_611,In_947);
xnor U481 (N_481,In_1415,In_1868);
nand U482 (N_482,In_1968,In_165);
nand U483 (N_483,In_1578,In_1508);
xnor U484 (N_484,In_1050,In_1129);
and U485 (N_485,In_1664,In_1241);
or U486 (N_486,In_1875,In_1377);
or U487 (N_487,In_1224,In_1323);
and U488 (N_488,In_819,In_1670);
nand U489 (N_489,In_554,In_1453);
nor U490 (N_490,In_658,In_1274);
or U491 (N_491,In_1116,In_845);
and U492 (N_492,In_1966,In_1494);
nand U493 (N_493,In_888,In_1941);
nand U494 (N_494,In_1996,In_1625);
nor U495 (N_495,In_545,In_28);
nand U496 (N_496,In_1764,In_168);
xnor U497 (N_497,In_1815,In_1098);
xnor U498 (N_498,In_223,In_1248);
and U499 (N_499,In_1025,In_869);
nor U500 (N_500,In_1305,In_397);
nor U501 (N_501,In_866,In_253);
and U502 (N_502,In_1348,In_279);
nand U503 (N_503,In_1908,In_883);
xnor U504 (N_504,In_321,In_1938);
xnor U505 (N_505,In_244,In_138);
nand U506 (N_506,In_1082,In_1235);
xnor U507 (N_507,In_719,In_564);
or U508 (N_508,In_237,In_207);
nand U509 (N_509,In_1433,In_416);
and U510 (N_510,In_1015,In_1057);
nor U511 (N_511,In_164,In_1479);
and U512 (N_512,In_133,In_985);
and U513 (N_513,In_1290,In_233);
and U514 (N_514,In_15,In_927);
and U515 (N_515,In_1655,In_1380);
xnor U516 (N_516,In_8,In_452);
nand U517 (N_517,In_735,In_306);
or U518 (N_518,In_979,In_934);
and U519 (N_519,In_908,In_143);
or U520 (N_520,In_533,In_1767);
nand U521 (N_521,In_1591,In_1619);
nand U522 (N_522,In_293,In_1504);
xor U523 (N_523,In_616,In_821);
nor U524 (N_524,In_1422,In_1247);
xor U525 (N_525,In_103,In_1604);
nand U526 (N_526,In_858,In_158);
nand U527 (N_527,In_991,In_455);
and U528 (N_528,In_895,In_678);
or U529 (N_529,In_411,In_604);
nor U530 (N_530,In_276,In_154);
or U531 (N_531,In_1639,In_468);
and U532 (N_532,In_1392,In_1218);
or U533 (N_533,In_1642,In_1813);
nand U534 (N_534,In_1447,In_1603);
and U535 (N_535,In_1044,In_450);
nor U536 (N_536,In_964,In_56);
or U537 (N_537,In_938,In_1324);
or U538 (N_538,In_40,In_1231);
xnor U539 (N_539,In_171,In_406);
nand U540 (N_540,In_419,In_970);
or U541 (N_541,In_860,In_1303);
xor U542 (N_542,In_382,In_797);
or U543 (N_543,In_1776,In_578);
and U544 (N_544,In_1311,In_1251);
nand U545 (N_545,In_1293,In_465);
and U546 (N_546,In_631,In_1805);
nand U547 (N_547,In_1987,In_1651);
xor U548 (N_548,In_197,In_1839);
nand U549 (N_549,In_1955,In_68);
and U550 (N_550,In_1081,In_1242);
nand U551 (N_551,In_590,In_907);
xor U552 (N_552,In_1981,In_257);
nand U553 (N_553,In_627,In_1975);
xnor U554 (N_554,In_1746,In_1592);
xor U555 (N_555,In_1983,In_1252);
and U556 (N_556,In_1699,In_1656);
nor U557 (N_557,In_1653,In_1921);
xor U558 (N_558,In_1910,In_1629);
nor U559 (N_559,In_1033,In_33);
nor U560 (N_560,In_707,In_1876);
nor U561 (N_561,In_836,In_597);
nand U562 (N_562,In_1787,In_291);
or U563 (N_563,In_1838,In_966);
nand U564 (N_564,In_1117,In_1771);
or U565 (N_565,In_1902,In_1355);
or U566 (N_566,In_1773,In_527);
xnor U567 (N_567,In_504,In_346);
and U568 (N_568,In_213,In_1282);
nor U569 (N_569,In_432,In_1136);
and U570 (N_570,In_12,In_705);
nor U571 (N_571,In_1689,In_517);
and U572 (N_572,In_1895,In_155);
or U573 (N_573,In_1,In_844);
and U574 (N_574,In_1300,In_1858);
or U575 (N_575,In_214,In_218);
xnor U576 (N_576,In_500,In_1550);
and U577 (N_577,In_161,In_48);
and U578 (N_578,In_600,In_624);
and U579 (N_579,In_96,In_1911);
nand U580 (N_580,In_1901,In_1587);
and U581 (N_581,In_808,In_116);
nand U582 (N_582,In_1403,In_975);
and U583 (N_583,In_1225,In_153);
nand U584 (N_584,In_1538,In_1847);
and U585 (N_585,In_1643,In_651);
and U586 (N_586,In_7,In_1008);
and U587 (N_587,In_613,In_893);
and U588 (N_588,In_1641,In_1331);
nor U589 (N_589,In_1109,In_1923);
xor U590 (N_590,In_180,In_1100);
nand U591 (N_591,In_1897,In_457);
xnor U592 (N_592,In_1291,In_1179);
xnor U593 (N_593,In_263,In_359);
nand U594 (N_594,In_471,In_362);
and U595 (N_595,In_1094,In_1391);
or U596 (N_596,In_1371,In_695);
xor U597 (N_597,In_1701,In_489);
nand U598 (N_598,In_756,In_1361);
and U599 (N_599,In_1672,In_737);
nor U600 (N_600,In_1832,In_814);
xor U601 (N_601,In_718,In_215);
and U602 (N_602,In_1931,In_992);
nor U603 (N_603,In_1680,In_1071);
or U604 (N_604,In_378,In_760);
or U605 (N_605,In_114,In_247);
or U606 (N_606,In_417,In_1543);
nor U607 (N_607,In_603,In_1675);
xor U608 (N_608,In_1429,In_1489);
nor U609 (N_609,In_1862,In_632);
nand U610 (N_610,In_1264,In_746);
nor U611 (N_611,In_1703,In_1012);
nand U612 (N_612,In_1542,In_859);
and U613 (N_613,In_297,In_1846);
xnor U614 (N_614,In_364,In_383);
and U615 (N_615,In_89,In_148);
nand U616 (N_616,In_1164,In_412);
nor U617 (N_617,In_954,In_1674);
nor U618 (N_618,In_762,In_1818);
and U619 (N_619,In_978,In_423);
nor U620 (N_620,In_1943,In_1203);
and U621 (N_621,In_903,In_159);
and U622 (N_622,In_968,In_456);
xnor U623 (N_623,In_1540,In_898);
nor U624 (N_624,In_1952,In_610);
and U625 (N_625,In_645,In_1162);
nor U626 (N_626,In_950,In_1051);
nor U627 (N_627,In_1511,In_682);
or U628 (N_628,In_269,In_1333);
nand U629 (N_629,In_525,In_502);
and U630 (N_630,In_1951,In_1920);
nor U631 (N_631,In_1678,In_683);
nor U632 (N_632,In_913,In_115);
or U633 (N_633,In_476,In_572);
nor U634 (N_634,In_922,In_1443);
or U635 (N_635,In_1960,In_1097);
nor U636 (N_636,In_1654,In_1263);
or U637 (N_637,In_1695,In_42);
nand U638 (N_638,In_1337,In_1485);
xnor U639 (N_639,In_1777,In_1315);
nand U640 (N_640,In_50,In_1696);
xor U641 (N_641,In_1475,In_1693);
nor U642 (N_642,In_793,In_1435);
or U643 (N_643,In_477,In_1153);
or U644 (N_644,In_1576,In_661);
nor U645 (N_645,In_636,In_71);
or U646 (N_646,In_846,In_66);
and U647 (N_647,In_86,In_1934);
nor U648 (N_648,In_1596,In_1173);
and U649 (N_649,In_351,In_1811);
nand U650 (N_650,In_1317,In_981);
or U651 (N_651,In_264,In_5);
nand U652 (N_652,In_1069,In_396);
nor U653 (N_653,In_1523,In_234);
and U654 (N_654,In_360,In_863);
and U655 (N_655,In_243,In_1048);
nor U656 (N_656,In_1473,In_1497);
xnor U657 (N_657,In_444,In_936);
nor U658 (N_658,In_1373,In_820);
nor U659 (N_659,In_1510,In_1559);
xnor U660 (N_660,In_1181,In_21);
nand U661 (N_661,In_1028,In_721);
or U662 (N_662,In_1903,In_1808);
or U663 (N_663,In_1295,In_1156);
or U664 (N_664,In_1385,In_1649);
or U665 (N_665,In_538,In_794);
nor U666 (N_666,In_1169,In_1104);
and U667 (N_667,In_1631,In_1463);
or U668 (N_668,In_1119,In_1886);
nor U669 (N_669,In_1660,In_1287);
nor U670 (N_670,In_648,In_1707);
xor U671 (N_671,In_1717,In_162);
or U672 (N_672,In_1570,In_248);
or U673 (N_673,In_546,In_1796);
or U674 (N_674,In_635,In_891);
and U675 (N_675,In_856,In_1483);
and U676 (N_676,In_1108,In_195);
nand U677 (N_677,In_172,In_374);
and U678 (N_678,In_1237,In_105);
nor U679 (N_679,In_1085,In_557);
nand U680 (N_680,In_1541,In_1999);
nor U681 (N_681,In_1668,In_1049);
or U682 (N_682,In_1725,In_316);
xnor U683 (N_683,In_1065,In_1727);
and U684 (N_684,In_1467,In_1857);
nand U685 (N_685,In_1329,In_523);
nand U686 (N_686,In_815,In_1763);
nor U687 (N_687,In_1569,In_69);
nor U688 (N_688,In_582,In_129);
nor U689 (N_689,In_1045,In_1713);
or U690 (N_690,In_59,In_1112);
or U691 (N_691,In_1227,In_1563);
xor U692 (N_692,In_929,In_1748);
xnor U693 (N_693,In_1180,In_559);
or U694 (N_694,In_1522,In_1314);
xor U695 (N_695,In_1113,In_240);
xnor U696 (N_696,In_1382,In_621);
xor U697 (N_697,In_1788,In_702);
nand U698 (N_698,In_409,In_1004);
and U699 (N_699,In_1942,In_1365);
and U700 (N_700,In_759,In_1159);
nand U701 (N_701,In_1790,In_761);
and U702 (N_702,In_1801,In_1163);
or U703 (N_703,In_1940,In_1131);
and U704 (N_704,In_1882,In_1493);
or U705 (N_705,In_95,In_980);
nor U706 (N_706,In_1666,In_147);
nand U707 (N_707,In_1525,In_1009);
and U708 (N_708,In_479,In_1233);
and U709 (N_709,In_833,In_224);
or U710 (N_710,In_524,In_460);
and U711 (N_711,In_335,In_1843);
nand U712 (N_712,In_1465,In_77);
xnor U713 (N_713,In_131,In_1344);
or U714 (N_714,In_777,In_829);
nor U715 (N_715,In_369,In_744);
xnor U716 (N_716,In_847,In_1114);
xnor U717 (N_717,In_250,In_32);
nor U718 (N_718,In_470,In_404);
or U719 (N_719,In_850,In_1791);
xor U720 (N_720,In_318,In_1118);
nand U721 (N_721,In_583,In_1667);
and U722 (N_722,In_1544,In_286);
nor U723 (N_723,In_1918,In_117);
or U724 (N_724,In_536,In_124);
nor U725 (N_725,In_996,In_1733);
nand U726 (N_726,In_18,In_1623);
nand U727 (N_727,In_1814,In_1537);
nand U728 (N_728,In_1755,In_1750);
nor U729 (N_729,In_896,In_451);
xnor U730 (N_730,In_1851,In_349);
or U731 (N_731,In_880,In_426);
and U732 (N_732,In_1885,In_1121);
and U733 (N_733,In_830,In_877);
or U734 (N_734,In_1555,In_258);
xor U735 (N_735,In_585,In_890);
nand U736 (N_736,In_725,In_492);
or U737 (N_737,In_834,In_1634);
xnor U738 (N_738,In_1390,In_1919);
nor U739 (N_739,In_835,In_1105);
nor U740 (N_740,In_109,In_173);
or U741 (N_741,In_1176,In_189);
and U742 (N_742,In_1661,In_1599);
nor U743 (N_743,In_1756,In_780);
nor U744 (N_744,In_1455,In_83);
and U745 (N_745,In_312,In_209);
or U746 (N_746,In_1154,In_1448);
and U747 (N_747,In_1648,In_437);
nand U748 (N_748,In_1833,In_1438);
or U749 (N_749,In_398,In_1636);
and U750 (N_750,In_827,In_998);
nor U751 (N_751,In_413,In_122);
and U752 (N_752,In_1626,In_1937);
xor U753 (N_753,In_495,In_983);
or U754 (N_754,In_1562,In_1898);
or U755 (N_755,In_17,In_602);
and U756 (N_756,In_1318,In_262);
xor U757 (N_757,In_127,In_405);
xor U758 (N_758,In_722,In_764);
xnor U759 (N_759,In_986,In_1844);
nor U760 (N_760,In_568,In_1167);
and U761 (N_761,In_790,In_1866);
xor U762 (N_762,In_1157,In_1989);
nor U763 (N_763,In_1712,In_219);
nand U764 (N_764,In_962,In_1650);
nor U765 (N_765,In_102,In_1205);
nand U766 (N_766,In_1378,In_283);
nand U767 (N_767,In_1137,In_177);
nand U768 (N_768,In_1744,In_259);
and U769 (N_769,In_1021,In_106);
xor U770 (N_770,In_1747,In_729);
or U771 (N_771,In_221,In_587);
and U772 (N_772,In_119,In_228);
xor U773 (N_773,In_1769,In_342);
or U774 (N_774,In_1816,In_1321);
or U775 (N_775,In_1884,In_945);
nor U776 (N_776,In_238,In_188);
nor U777 (N_777,In_801,In_842);
nand U778 (N_778,In_1362,In_388);
nand U779 (N_779,In_1518,In_261);
and U780 (N_780,In_1027,In_511);
nand U781 (N_781,In_868,In_1594);
xnor U782 (N_782,In_530,In_361);
nand U783 (N_783,In_693,In_711);
or U784 (N_784,In_393,In_1036);
and U785 (N_785,In_1102,In_80);
and U786 (N_786,In_1681,In_1288);
and U787 (N_787,In_1507,In_1620);
nand U788 (N_788,In_271,In_881);
xor U789 (N_789,In_694,In_714);
nand U790 (N_790,In_1326,In_1232);
or U791 (N_791,In_717,In_1334);
nor U792 (N_792,In_428,In_1010);
nand U793 (N_793,In_1685,In_918);
xor U794 (N_794,In_1617,In_615);
xnor U795 (N_795,In_1698,In_175);
or U796 (N_796,In_1495,In_1405);
nor U797 (N_797,In_1346,In_141);
and U798 (N_798,In_418,In_381);
nor U799 (N_799,In_1573,In_1468);
or U800 (N_800,In_137,In_191);
or U801 (N_801,In_1831,In_23);
or U802 (N_802,In_1948,In_1740);
or U803 (N_803,In_855,In_217);
xor U804 (N_804,In_1589,In_736);
nor U805 (N_805,In_1089,In_230);
xor U806 (N_806,In_1002,In_1889);
and U807 (N_807,In_104,In_1007);
xor U808 (N_808,In_1714,In_320);
xnor U809 (N_809,In_1819,In_1500);
nor U810 (N_810,In_1741,In_178);
and U811 (N_811,In_752,In_1936);
and U812 (N_812,In_1243,In_387);
xor U813 (N_813,In_490,In_1394);
nand U814 (N_814,In_569,In_1530);
nand U815 (N_815,In_629,In_1450);
xnor U816 (N_816,In_878,In_1887);
nor U817 (N_817,In_1258,In_389);
nor U818 (N_818,In_435,In_1445);
or U819 (N_819,In_1427,In_1253);
xnor U820 (N_820,In_1419,In_698);
nand U821 (N_821,In_526,In_93);
or U822 (N_822,In_823,In_1434);
and U823 (N_823,In_1881,In_395);
and U824 (N_824,In_1837,In_392);
nand U825 (N_825,In_482,In_1869);
nand U826 (N_826,In_1216,In_1546);
nand U827 (N_827,In_1298,In_462);
xnor U828 (N_828,In_1490,In_313);
nor U829 (N_829,In_654,In_1019);
or U830 (N_830,In_909,In_294);
and U831 (N_831,In_1208,In_1528);
and U832 (N_832,In_713,In_1496);
nand U833 (N_833,In_220,In_327);
nor U834 (N_834,In_1146,In_1752);
nor U835 (N_835,In_1255,In_1988);
and U836 (N_836,In_739,In_1915);
and U837 (N_837,In_290,In_260);
nand U838 (N_838,In_571,In_575);
nand U839 (N_839,In_1652,In_1320);
and U840 (N_840,In_534,In_1187);
xnor U841 (N_841,In_990,In_1199);
nor U842 (N_842,In_181,In_461);
nor U843 (N_843,In_81,In_666);
or U844 (N_844,In_123,In_1353);
nand U845 (N_845,In_386,In_696);
and U846 (N_846,In_402,In_1532);
or U847 (N_847,In_194,In_1067);
nand U848 (N_848,In_145,In_333);
or U849 (N_849,In_52,In_1804);
xnor U850 (N_850,In_466,In_328);
and U851 (N_851,In_501,In_1549);
and U852 (N_852,In_356,In_1190);
and U853 (N_853,In_656,In_905);
nor U854 (N_854,In_1408,In_338);
nand U855 (N_855,In_1343,In_372);
and U856 (N_856,In_1515,In_0);
nand U857 (N_857,In_848,In_677);
xor U858 (N_858,In_553,In_566);
and U859 (N_859,In_1234,In_1359);
nor U860 (N_860,In_1428,In_1659);
nand U861 (N_861,In_1409,In_1836);
or U862 (N_862,In_1350,In_1425);
nand U863 (N_863,In_1935,In_1778);
nor U864 (N_864,In_118,In_1166);
or U865 (N_865,In_449,In_1206);
nor U866 (N_866,In_1143,In_601);
xor U867 (N_867,In_977,In_1289);
xor U868 (N_868,In_663,In_589);
and U869 (N_869,In_348,In_478);
xor U870 (N_870,In_1383,In_662);
xor U871 (N_871,In_1451,In_464);
nor U872 (N_872,In_625,In_19);
or U873 (N_873,In_1925,In_1150);
xor U874 (N_874,In_1041,In_1835);
xor U875 (N_875,In_726,In_1335);
or U876 (N_876,In_1426,In_1177);
nor U877 (N_877,In_1437,In_1548);
nand U878 (N_878,In_146,In_1226);
nor U879 (N_879,In_132,In_1624);
or U880 (N_880,In_1580,In_1062);
nor U881 (N_881,In_1040,In_174);
and U882 (N_882,In_25,In_268);
nor U883 (N_883,In_1458,In_1186);
and U884 (N_884,In_857,In_1793);
nor U885 (N_885,In_1749,In_1030);
nor U886 (N_886,In_458,In_1535);
xor U887 (N_887,In_1644,In_1283);
or U888 (N_888,In_390,In_1760);
nand U889 (N_889,In_367,In_556);
nor U890 (N_890,In_1063,In_769);
nor U891 (N_891,In_494,In_1120);
nand U892 (N_892,In_1946,In_520);
xor U893 (N_893,In_443,In_1292);
nor U894 (N_894,In_212,In_1673);
nand U895 (N_895,In_1524,In_201);
nand U896 (N_896,In_942,In_1014);
nor U897 (N_897,In_634,In_58);
nor U898 (N_898,In_655,In_399);
xnor U899 (N_899,In_993,In_41);
xnor U900 (N_900,In_431,In_1613);
xnor U901 (N_901,In_1691,In_1342);
nand U902 (N_902,In_267,In_510);
nand U903 (N_903,In_1476,In_943);
nand U904 (N_904,In_516,In_1802);
nor U905 (N_905,In_612,In_688);
or U906 (N_906,In_1635,In_1393);
or U907 (N_907,In_1807,In_1870);
nor U908 (N_908,In_1726,In_1259);
or U909 (N_909,In_1456,In_1418);
and U910 (N_910,In_1297,In_384);
nor U911 (N_911,In_1616,In_135);
xor U912 (N_912,In_813,In_1840);
and U913 (N_913,In_1406,In_1499);
nand U914 (N_914,In_514,In_1022);
or U915 (N_915,In_828,In_474);
nand U916 (N_916,In_1671,In_838);
or U917 (N_917,In_1275,In_770);
and U918 (N_918,In_1306,In_1037);
and U919 (N_919,In_1236,In_1407);
nand U920 (N_920,In_22,In_1327);
nand U921 (N_921,In_1209,In_804);
nor U922 (N_922,In_673,In_1800);
nor U923 (N_923,In_1149,In_643);
nor U924 (N_924,In_1894,In_1779);
and U925 (N_925,In_917,In_1268);
and U926 (N_926,In_4,In_1454);
nor U927 (N_927,In_49,In_1647);
nand U928 (N_928,In_560,In_933);
or U929 (N_929,In_1775,In_1856);
and U930 (N_930,In_659,In_1863);
and U931 (N_931,In_1841,In_727);
or U932 (N_932,In_391,In_509);
or U933 (N_933,In_1958,In_484);
or U934 (N_934,In_620,In_1389);
nand U935 (N_935,In_336,In_644);
nand U936 (N_936,In_1139,In_1560);
and U937 (N_937,In_292,In_1013);
or U938 (N_938,In_872,In_298);
nand U939 (N_939,In_156,In_200);
or U940 (N_940,In_789,In_684);
nand U941 (N_941,In_1039,In_1148);
and U942 (N_942,In_366,In_928);
nor U943 (N_943,In_775,In_1547);
or U944 (N_944,In_1962,In_641);
and U945 (N_945,In_1466,In_1093);
xor U946 (N_946,In_605,In_480);
or U947 (N_947,In_447,In_686);
or U948 (N_948,In_745,In_459);
and U949 (N_949,In_125,In_332);
or U950 (N_950,In_811,In_1849);
and U951 (N_951,In_498,In_1276);
nand U952 (N_952,In_967,In_1963);
nand U953 (N_953,In_1230,In_400);
xor U954 (N_954,In_211,In_618);
xor U955 (N_955,In_1397,In_441);
nor U956 (N_956,In_930,In_916);
nor U957 (N_957,In_422,In_368);
xor U958 (N_958,In_24,In_579);
nor U959 (N_959,In_1612,In_1842);
or U960 (N_960,In_323,In_1060);
nand U961 (N_961,In_1824,In_1035);
and U962 (N_962,In_454,In_822);
or U963 (N_963,In_1301,In_882);
nand U964 (N_964,In_1266,In_912);
and U965 (N_965,In_784,In_1413);
nand U966 (N_966,In_1774,In_1632);
nor U967 (N_967,In_1687,In_1155);
nor U968 (N_968,In_304,In_251);
or U969 (N_969,In_765,In_873);
and U970 (N_970,In_242,In_1280);
nand U971 (N_971,In_1341,In_1618);
xor U972 (N_972,In_241,In_1006);
and U973 (N_973,In_540,In_1950);
and U974 (N_974,In_939,In_1728);
xor U975 (N_975,In_1281,In_894);
nand U976 (N_976,In_1059,In_874);
nand U977 (N_977,In_1501,In_1947);
nand U978 (N_978,In_586,In_728);
nand U979 (N_979,In_179,In_1398);
nor U980 (N_980,In_14,In_1446);
and U981 (N_981,In_55,In_818);
and U982 (N_982,In_1900,In_1506);
xor U983 (N_983,In_919,In_638);
or U984 (N_984,In_1034,In_731);
or U985 (N_985,In_1828,In_709);
xor U986 (N_986,In_310,In_900);
nand U987 (N_987,In_940,In_1269);
nor U988 (N_988,In_75,In_529);
or U989 (N_989,In_512,In_6);
or U990 (N_990,In_1586,In_1417);
nor U991 (N_991,In_1610,In_1956);
xnor U992 (N_992,In_47,In_1200);
xor U993 (N_993,In_1354,In_879);
nand U994 (N_994,In_1211,In_1737);
and U995 (N_995,In_1929,In_44);
and U996 (N_996,In_190,In_1133);
and U997 (N_997,In_1042,In_561);
nor U998 (N_998,In_1058,In_1637);
nor U999 (N_999,In_35,In_1893);
and U1000 (N_1000,N_198,N_514);
or U1001 (N_1001,N_875,N_94);
and U1002 (N_1002,N_114,N_453);
xnor U1003 (N_1003,N_745,N_278);
nand U1004 (N_1004,N_771,N_392);
and U1005 (N_1005,N_192,N_911);
xnor U1006 (N_1006,N_426,N_787);
nor U1007 (N_1007,N_471,N_482);
xnor U1008 (N_1008,N_21,N_661);
nor U1009 (N_1009,N_690,N_165);
nor U1010 (N_1010,N_579,N_190);
or U1011 (N_1011,N_971,N_552);
and U1012 (N_1012,N_731,N_646);
or U1013 (N_1013,N_536,N_334);
or U1014 (N_1014,N_166,N_587);
xor U1015 (N_1015,N_513,N_721);
or U1016 (N_1016,N_119,N_649);
nor U1017 (N_1017,N_885,N_125);
and U1018 (N_1018,N_358,N_491);
or U1019 (N_1019,N_857,N_889);
nor U1020 (N_1020,N_707,N_765);
xnor U1021 (N_1021,N_312,N_995);
nand U1022 (N_1022,N_264,N_769);
or U1023 (N_1023,N_757,N_935);
nand U1024 (N_1024,N_624,N_922);
or U1025 (N_1025,N_508,N_997);
nor U1026 (N_1026,N_152,N_148);
or U1027 (N_1027,N_977,N_778);
or U1028 (N_1028,N_147,N_728);
xor U1029 (N_1029,N_770,N_446);
xnor U1030 (N_1030,N_395,N_283);
nand U1031 (N_1031,N_443,N_989);
nor U1032 (N_1032,N_247,N_293);
and U1033 (N_1033,N_355,N_274);
xnor U1034 (N_1034,N_241,N_343);
or U1035 (N_1035,N_478,N_159);
or U1036 (N_1036,N_724,N_651);
xor U1037 (N_1037,N_946,N_973);
and U1038 (N_1038,N_258,N_527);
nor U1039 (N_1039,N_52,N_703);
and U1040 (N_1040,N_434,N_479);
xor U1041 (N_1041,N_883,N_128);
nand U1042 (N_1042,N_506,N_149);
nor U1043 (N_1043,N_562,N_43);
or U1044 (N_1044,N_77,N_755);
xnor U1045 (N_1045,N_687,N_341);
or U1046 (N_1046,N_79,N_408);
and U1047 (N_1047,N_447,N_678);
xor U1048 (N_1048,N_591,N_254);
or U1049 (N_1049,N_75,N_457);
and U1050 (N_1050,N_277,N_713);
xor U1051 (N_1051,N_608,N_390);
xnor U1052 (N_1052,N_620,N_310);
or U1053 (N_1053,N_958,N_715);
nand U1054 (N_1054,N_982,N_1);
xnor U1055 (N_1055,N_581,N_841);
nand U1056 (N_1056,N_679,N_511);
and U1057 (N_1057,N_378,N_336);
nor U1058 (N_1058,N_969,N_618);
xnor U1059 (N_1059,N_73,N_898);
xnor U1060 (N_1060,N_311,N_349);
and U1061 (N_1061,N_696,N_637);
nor U1062 (N_1062,N_409,N_531);
or U1063 (N_1063,N_486,N_196);
nor U1064 (N_1064,N_689,N_641);
or U1065 (N_1065,N_464,N_570);
nand U1066 (N_1066,N_782,N_229);
or U1067 (N_1067,N_932,N_677);
nand U1068 (N_1068,N_671,N_961);
nor U1069 (N_1069,N_580,N_490);
and U1070 (N_1070,N_811,N_203);
and U1071 (N_1071,N_298,N_427);
xnor U1072 (N_1072,N_297,N_156);
nor U1073 (N_1073,N_122,N_786);
or U1074 (N_1074,N_146,N_880);
nand U1075 (N_1075,N_112,N_217);
and U1076 (N_1076,N_548,N_628);
nor U1077 (N_1077,N_215,N_741);
or U1078 (N_1078,N_947,N_442);
and U1079 (N_1079,N_107,N_137);
or U1080 (N_1080,N_444,N_80);
nand U1081 (N_1081,N_567,N_10);
and U1082 (N_1082,N_424,N_8);
and U1083 (N_1083,N_586,N_981);
or U1084 (N_1084,N_597,N_924);
nand U1085 (N_1085,N_960,N_894);
nand U1086 (N_1086,N_403,N_759);
or U1087 (N_1087,N_899,N_55);
xnor U1088 (N_1088,N_244,N_131);
nand U1089 (N_1089,N_228,N_539);
and U1090 (N_1090,N_81,N_465);
and U1091 (N_1091,N_942,N_940);
and U1092 (N_1092,N_939,N_36);
xnor U1093 (N_1093,N_472,N_74);
or U1094 (N_1094,N_111,N_124);
nor U1095 (N_1095,N_136,N_705);
nor U1096 (N_1096,N_344,N_384);
and U1097 (N_1097,N_139,N_154);
nor U1098 (N_1098,N_595,N_550);
xnor U1099 (N_1099,N_379,N_884);
nand U1100 (N_1100,N_207,N_510);
nand U1101 (N_1101,N_991,N_351);
xor U1102 (N_1102,N_406,N_420);
xor U1103 (N_1103,N_907,N_616);
and U1104 (N_1104,N_369,N_199);
and U1105 (N_1105,N_126,N_176);
xor U1106 (N_1106,N_342,N_585);
nor U1107 (N_1107,N_463,N_633);
nand U1108 (N_1108,N_200,N_415);
nor U1109 (N_1109,N_321,N_142);
xor U1110 (N_1110,N_615,N_121);
xnor U1111 (N_1111,N_610,N_487);
and U1112 (N_1112,N_520,N_996);
and U1113 (N_1113,N_90,N_402);
and U1114 (N_1114,N_167,N_993);
or U1115 (N_1115,N_812,N_727);
or U1116 (N_1116,N_57,N_507);
nand U1117 (N_1117,N_662,N_239);
and U1118 (N_1118,N_557,N_632);
or U1119 (N_1119,N_177,N_326);
nand U1120 (N_1120,N_938,N_454);
xor U1121 (N_1121,N_668,N_599);
nand U1122 (N_1122,N_819,N_927);
xor U1123 (N_1123,N_323,N_452);
or U1124 (N_1124,N_364,N_459);
or U1125 (N_1125,N_584,N_158);
or U1126 (N_1126,N_855,N_639);
nand U1127 (N_1127,N_861,N_19);
or U1128 (N_1128,N_40,N_596);
nand U1129 (N_1129,N_157,N_746);
or U1130 (N_1130,N_951,N_505);
xor U1131 (N_1131,N_860,N_84);
nor U1132 (N_1132,N_308,N_399);
and U1133 (N_1133,N_280,N_685);
or U1134 (N_1134,N_161,N_774);
nor U1135 (N_1135,N_743,N_181);
and U1136 (N_1136,N_231,N_856);
and U1137 (N_1137,N_734,N_357);
nand U1138 (N_1138,N_46,N_617);
nor U1139 (N_1139,N_120,N_163);
nand U1140 (N_1140,N_523,N_791);
nand U1141 (N_1141,N_793,N_162);
or U1142 (N_1142,N_0,N_448);
nor U1143 (N_1143,N_692,N_260);
nor U1144 (N_1144,N_495,N_317);
and U1145 (N_1145,N_914,N_598);
nor U1146 (N_1146,N_423,N_389);
nand U1147 (N_1147,N_847,N_698);
nand U1148 (N_1148,N_288,N_96);
nand U1149 (N_1149,N_381,N_56);
nor U1150 (N_1150,N_890,N_422);
or U1151 (N_1151,N_645,N_895);
nand U1152 (N_1152,N_467,N_886);
and U1153 (N_1153,N_612,N_909);
xnor U1154 (N_1154,N_71,N_603);
xnor U1155 (N_1155,N_469,N_930);
and U1156 (N_1156,N_761,N_391);
xnor U1157 (N_1157,N_450,N_413);
or U1158 (N_1158,N_42,N_974);
xnor U1159 (N_1159,N_566,N_695);
nand U1160 (N_1160,N_493,N_220);
or U1161 (N_1161,N_376,N_301);
and U1162 (N_1162,N_213,N_431);
nand U1163 (N_1163,N_943,N_556);
xnor U1164 (N_1164,N_150,N_929);
xnor U1165 (N_1165,N_65,N_955);
or U1166 (N_1166,N_540,N_754);
xor U1167 (N_1167,N_904,N_848);
or U1168 (N_1168,N_265,N_809);
nor U1169 (N_1169,N_22,N_606);
xor U1170 (N_1170,N_717,N_370);
and U1171 (N_1171,N_232,N_750);
and U1172 (N_1172,N_625,N_913);
or U1173 (N_1173,N_551,N_103);
nand U1174 (N_1174,N_691,N_99);
nor U1175 (N_1175,N_656,N_998);
xnor U1176 (N_1176,N_307,N_908);
or U1177 (N_1177,N_416,N_327);
xor U1178 (N_1178,N_316,N_115);
nor U1179 (N_1179,N_795,N_218);
or U1180 (N_1180,N_693,N_180);
or U1181 (N_1181,N_186,N_708);
nand U1182 (N_1182,N_638,N_840);
xnor U1183 (N_1183,N_257,N_63);
or U1184 (N_1184,N_172,N_964);
and U1185 (N_1185,N_132,N_843);
nand U1186 (N_1186,N_936,N_484);
and U1187 (N_1187,N_365,N_817);
nand U1188 (N_1188,N_674,N_322);
or U1189 (N_1189,N_397,N_398);
and U1190 (N_1190,N_534,N_498);
and U1191 (N_1191,N_50,N_533);
and U1192 (N_1192,N_794,N_91);
nor U1193 (N_1193,N_779,N_345);
nand U1194 (N_1194,N_752,N_474);
nor U1195 (N_1195,N_572,N_171);
or U1196 (N_1196,N_286,N_78);
or U1197 (N_1197,N_396,N_489);
nand U1198 (N_1198,N_235,N_460);
and U1199 (N_1199,N_151,N_699);
nand U1200 (N_1200,N_204,N_517);
or U1201 (N_1201,N_711,N_667);
xor U1202 (N_1202,N_101,N_823);
xnor U1203 (N_1203,N_243,N_836);
nor U1204 (N_1204,N_944,N_375);
nor U1205 (N_1205,N_3,N_990);
and U1206 (N_1206,N_648,N_335);
and U1207 (N_1207,N_437,N_829);
and U1208 (N_1208,N_828,N_411);
or U1209 (N_1209,N_141,N_547);
nor U1210 (N_1210,N_97,N_653);
xnor U1211 (N_1211,N_810,N_503);
nor U1212 (N_1212,N_887,N_155);
or U1213 (N_1213,N_593,N_354);
nand U1214 (N_1214,N_796,N_783);
or U1215 (N_1215,N_153,N_558);
or U1216 (N_1216,N_4,N_762);
or U1217 (N_1217,N_109,N_480);
xor U1218 (N_1218,N_643,N_33);
xor U1219 (N_1219,N_462,N_330);
nand U1220 (N_1220,N_234,N_306);
nor U1221 (N_1221,N_549,N_401);
and U1222 (N_1222,N_455,N_35);
or U1223 (N_1223,N_532,N_135);
nand U1224 (N_1224,N_882,N_704);
or U1225 (N_1225,N_921,N_193);
xor U1226 (N_1226,N_528,N_304);
or U1227 (N_1227,N_920,N_838);
and U1228 (N_1228,N_631,N_582);
or U1229 (N_1229,N_85,N_225);
xnor U1230 (N_1230,N_105,N_282);
or U1231 (N_1231,N_377,N_979);
or U1232 (N_1232,N_339,N_303);
and U1233 (N_1233,N_952,N_576);
or U1234 (N_1234,N_594,N_877);
nand U1235 (N_1235,N_729,N_833);
nand U1236 (N_1236,N_451,N_976);
xor U1237 (N_1237,N_32,N_133);
nor U1238 (N_1238,N_26,N_834);
nor U1239 (N_1239,N_499,N_227);
xor U1240 (N_1240,N_792,N_205);
nand U1241 (N_1241,N_476,N_751);
nand U1242 (N_1242,N_660,N_160);
nand U1243 (N_1243,N_799,N_360);
or U1244 (N_1244,N_92,N_440);
nand U1245 (N_1245,N_170,N_98);
or U1246 (N_1246,N_9,N_983);
and U1247 (N_1247,N_429,N_726);
nand U1248 (N_1248,N_688,N_577);
xnor U1249 (N_1249,N_915,N_337);
xor U1250 (N_1250,N_530,N_30);
nand U1251 (N_1251,N_305,N_901);
nor U1252 (N_1252,N_134,N_54);
and U1253 (N_1253,N_820,N_24);
nor U1254 (N_1254,N_972,N_916);
nor U1255 (N_1255,N_742,N_845);
nor U1256 (N_1256,N_607,N_421);
and U1257 (N_1257,N_12,N_201);
and U1258 (N_1258,N_965,N_826);
nand U1259 (N_1259,N_801,N_574);
and U1260 (N_1260,N_87,N_553);
xor U1261 (N_1261,N_872,N_363);
and U1262 (N_1262,N_108,N_412);
xor U1263 (N_1263,N_832,N_18);
xor U1264 (N_1264,N_373,N_256);
xor U1265 (N_1265,N_937,N_435);
nand U1266 (N_1266,N_623,N_439);
or U1267 (N_1267,N_502,N_723);
nand U1268 (N_1268,N_953,N_980);
xnor U1269 (N_1269,N_143,N_208);
nand U1270 (N_1270,N_737,N_481);
nand U1271 (N_1271,N_571,N_544);
nand U1272 (N_1272,N_388,N_758);
nand U1273 (N_1273,N_252,N_332);
or U1274 (N_1274,N_892,N_814);
and U1275 (N_1275,N_117,N_34);
and U1276 (N_1276,N_621,N_684);
nor U1277 (N_1277,N_28,N_417);
and U1278 (N_1278,N_554,N_372);
or U1279 (N_1279,N_945,N_869);
xnor U1280 (N_1280,N_784,N_39);
or U1281 (N_1281,N_211,N_605);
or U1282 (N_1282,N_863,N_565);
xnor U1283 (N_1283,N_483,N_338);
nand U1284 (N_1284,N_449,N_138);
and U1285 (N_1285,N_988,N_957);
nor U1286 (N_1286,N_197,N_106);
xor U1287 (N_1287,N_477,N_261);
nor U1288 (N_1288,N_492,N_44);
nor U1289 (N_1289,N_642,N_233);
or U1290 (N_1290,N_910,N_816);
or U1291 (N_1291,N_60,N_858);
nand U1292 (N_1292,N_179,N_735);
and U1293 (N_1293,N_622,N_800);
nor U1294 (N_1294,N_184,N_352);
xnor U1295 (N_1295,N_174,N_785);
and U1296 (N_1296,N_905,N_670);
and U1297 (N_1297,N_51,N_775);
xnor U1298 (N_1298,N_798,N_468);
xor U1299 (N_1299,N_564,N_130);
or U1300 (N_1300,N_314,N_64);
nor U1301 (N_1301,N_985,N_777);
nand U1302 (N_1302,N_366,N_309);
xor U1303 (N_1303,N_246,N_226);
nor U1304 (N_1304,N_903,N_780);
or U1305 (N_1305,N_830,N_318);
nand U1306 (N_1306,N_747,N_221);
nor U1307 (N_1307,N_831,N_986);
or U1308 (N_1308,N_665,N_569);
or U1309 (N_1309,N_730,N_815);
and U1310 (N_1310,N_521,N_331);
nand U1311 (N_1311,N_488,N_340);
xnor U1312 (N_1312,N_613,N_419);
or U1313 (N_1313,N_725,N_145);
xnor U1314 (N_1314,N_404,N_509);
nor U1315 (N_1315,N_950,N_763);
or U1316 (N_1316,N_249,N_191);
nor U1317 (N_1317,N_206,N_425);
nand U1318 (N_1318,N_825,N_850);
nor U1319 (N_1319,N_876,N_718);
xnor U1320 (N_1320,N_635,N_299);
or U1321 (N_1321,N_776,N_268);
xor U1322 (N_1322,N_676,N_854);
nor U1323 (N_1323,N_900,N_13);
and U1324 (N_1324,N_432,N_31);
xor U1325 (N_1325,N_879,N_797);
nand U1326 (N_1326,N_292,N_53);
xnor U1327 (N_1327,N_393,N_978);
and U1328 (N_1328,N_948,N_118);
nand U1329 (N_1329,N_526,N_933);
or U1330 (N_1330,N_712,N_822);
nand U1331 (N_1331,N_14,N_560);
and U1332 (N_1332,N_716,N_680);
xnor U1333 (N_1333,N_546,N_970);
and U1334 (N_1334,N_251,N_466);
nand U1335 (N_1335,N_319,N_963);
and U1336 (N_1336,N_385,N_592);
xor U1337 (N_1337,N_663,N_931);
nor U1338 (N_1338,N_275,N_273);
and U1339 (N_1339,N_89,N_7);
nand U1340 (N_1340,N_458,N_756);
and U1341 (N_1341,N_753,N_368);
nor U1342 (N_1342,N_992,N_868);
nand U1343 (N_1343,N_238,N_290);
and U1344 (N_1344,N_512,N_324);
xor U1345 (N_1345,N_348,N_543);
nand U1346 (N_1346,N_764,N_700);
xor U1347 (N_1347,N_430,N_906);
nor U1348 (N_1348,N_714,N_110);
xor U1349 (N_1349,N_654,N_789);
xnor U1350 (N_1350,N_966,N_561);
xor U1351 (N_1351,N_896,N_169);
xor U1352 (N_1352,N_237,N_709);
and U1353 (N_1353,N_697,N_760);
and U1354 (N_1354,N_144,N_949);
and U1355 (N_1355,N_767,N_296);
nor U1356 (N_1356,N_294,N_445);
nor U1357 (N_1357,N_563,N_600);
or U1358 (N_1358,N_140,N_362);
nand U1359 (N_1359,N_62,N_583);
xnor U1360 (N_1360,N_804,N_897);
nor U1361 (N_1361,N_164,N_5);
xnor U1362 (N_1362,N_320,N_891);
nor U1363 (N_1363,N_76,N_371);
nand U1364 (N_1364,N_281,N_744);
xor U1365 (N_1365,N_655,N_524);
xnor U1366 (N_1366,N_58,N_329);
or U1367 (N_1367,N_23,N_436);
xor U1368 (N_1368,N_954,N_934);
xor U1369 (N_1369,N_248,N_518);
and U1370 (N_1370,N_888,N_456);
nor U1371 (N_1371,N_129,N_739);
or U1372 (N_1372,N_15,N_195);
nand U1373 (N_1373,N_941,N_788);
nor U1374 (N_1374,N_808,N_470);
xnor U1375 (N_1375,N_473,N_367);
nor U1376 (N_1376,N_236,N_485);
nand U1377 (N_1377,N_844,N_640);
nor U1378 (N_1378,N_6,N_300);
and U1379 (N_1379,N_578,N_383);
or U1380 (N_1380,N_346,N_70);
nand U1381 (N_1381,N_59,N_504);
or U1382 (N_1382,N_515,N_636);
nor U1383 (N_1383,N_188,N_289);
and U1384 (N_1384,N_912,N_644);
xnor U1385 (N_1385,N_394,N_223);
xor U1386 (N_1386,N_67,N_871);
and U1387 (N_1387,N_266,N_202);
xor U1388 (N_1388,N_555,N_183);
or U1389 (N_1389,N_573,N_538);
nand U1390 (N_1390,N_189,N_500);
nand U1391 (N_1391,N_347,N_842);
nor U1392 (N_1392,N_720,N_999);
and U1393 (N_1393,N_272,N_328);
nor U1394 (N_1394,N_82,N_602);
and U1395 (N_1395,N_864,N_240);
nor U1396 (N_1396,N_497,N_611);
or U1397 (N_1397,N_433,N_102);
nor U1398 (N_1398,N_182,N_187);
xor U1399 (N_1399,N_925,N_919);
nor U1400 (N_1400,N_589,N_849);
or U1401 (N_1401,N_20,N_772);
nor U1402 (N_1402,N_738,N_496);
and U1403 (N_1403,N_859,N_669);
or U1404 (N_1404,N_287,N_262);
nor U1405 (N_1405,N_873,N_893);
or U1406 (N_1406,N_994,N_219);
or U1407 (N_1407,N_410,N_284);
xnor U1408 (N_1408,N_866,N_673);
or U1409 (N_1409,N_270,N_253);
and U1410 (N_1410,N_870,N_61);
or U1411 (N_1411,N_69,N_86);
nand U1412 (N_1412,N_387,N_874);
xor U1413 (N_1413,N_100,N_359);
or U1414 (N_1414,N_382,N_194);
nand U1415 (N_1415,N_768,N_17);
or U1416 (N_1416,N_749,N_630);
xnor U1417 (N_1417,N_271,N_400);
nor U1418 (N_1418,N_353,N_962);
and U1419 (N_1419,N_923,N_719);
nand U1420 (N_1420,N_88,N_881);
nor U1421 (N_1421,N_604,N_535);
nor U1422 (N_1422,N_173,N_45);
nor U1423 (N_1423,N_926,N_918);
xnor U1424 (N_1424,N_230,N_113);
or U1425 (N_1425,N_380,N_350);
or U1426 (N_1426,N_806,N_259);
nand U1427 (N_1427,N_537,N_790);
xnor U1428 (N_1428,N_250,N_66);
and U1429 (N_1429,N_706,N_659);
or U1430 (N_1430,N_210,N_650);
and U1431 (N_1431,N_839,N_501);
xnor U1432 (N_1432,N_116,N_601);
nor U1433 (N_1433,N_276,N_852);
xnor U1434 (N_1434,N_519,N_575);
nand U1435 (N_1435,N_862,N_878);
nand U1436 (N_1436,N_686,N_522);
nand U1437 (N_1437,N_732,N_682);
xor U1438 (N_1438,N_2,N_475);
xor U1439 (N_1439,N_414,N_529);
nand U1440 (N_1440,N_123,N_701);
and U1441 (N_1441,N_104,N_984);
nor U1442 (N_1442,N_694,N_867);
or U1443 (N_1443,N_333,N_629);
nor U1444 (N_1444,N_302,N_652);
nand U1445 (N_1445,N_16,N_541);
and U1446 (N_1446,N_48,N_559);
xnor U1447 (N_1447,N_619,N_975);
nand U1448 (N_1448,N_956,N_657);
nor U1449 (N_1449,N_245,N_545);
xor U1450 (N_1450,N_733,N_588);
nand U1451 (N_1451,N_664,N_647);
nand U1452 (N_1452,N_313,N_865);
and U1453 (N_1453,N_29,N_178);
or U1454 (N_1454,N_710,N_813);
or U1455 (N_1455,N_25,N_407);
xnor U1456 (N_1456,N_47,N_827);
or U1457 (N_1457,N_285,N_295);
and U1458 (N_1458,N_279,N_95);
nor U1459 (N_1459,N_291,N_525);
nand U1460 (N_1460,N_837,N_807);
nor U1461 (N_1461,N_766,N_516);
nand U1462 (N_1462,N_242,N_568);
and U1463 (N_1463,N_818,N_93);
nor U1464 (N_1464,N_267,N_803);
and U1465 (N_1465,N_418,N_781);
and U1466 (N_1466,N_185,N_11);
and U1467 (N_1467,N_325,N_967);
nor U1468 (N_1468,N_805,N_672);
xor U1469 (N_1469,N_851,N_374);
nand U1470 (N_1470,N_683,N_494);
and U1471 (N_1471,N_209,N_386);
nand U1472 (N_1472,N_255,N_987);
xnor U1473 (N_1473,N_461,N_917);
nand U1474 (N_1474,N_175,N_216);
and U1475 (N_1475,N_835,N_315);
or U1476 (N_1476,N_405,N_38);
and U1477 (N_1477,N_853,N_72);
nand U1478 (N_1478,N_675,N_748);
and U1479 (N_1479,N_658,N_37);
or U1480 (N_1480,N_928,N_168);
nand U1481 (N_1481,N_361,N_356);
nor U1482 (N_1482,N_773,N_740);
nor U1483 (N_1483,N_736,N_821);
xnor U1484 (N_1484,N_959,N_634);
nand U1485 (N_1485,N_27,N_127);
xor U1486 (N_1486,N_83,N_41);
xnor U1487 (N_1487,N_681,N_68);
and U1488 (N_1488,N_428,N_438);
xnor U1489 (N_1489,N_441,N_590);
xnor U1490 (N_1490,N_666,N_846);
nand U1491 (N_1491,N_224,N_626);
nor U1492 (N_1492,N_269,N_614);
nor U1493 (N_1493,N_609,N_542);
or U1494 (N_1494,N_702,N_627);
xor U1495 (N_1495,N_222,N_802);
xor U1496 (N_1496,N_263,N_968);
xor U1497 (N_1497,N_49,N_902);
nand U1498 (N_1498,N_824,N_722);
or U1499 (N_1499,N_212,N_214);
or U1500 (N_1500,N_304,N_563);
nor U1501 (N_1501,N_307,N_60);
nand U1502 (N_1502,N_606,N_519);
or U1503 (N_1503,N_173,N_416);
or U1504 (N_1504,N_225,N_669);
and U1505 (N_1505,N_993,N_245);
nand U1506 (N_1506,N_566,N_692);
and U1507 (N_1507,N_129,N_313);
xor U1508 (N_1508,N_328,N_781);
xnor U1509 (N_1509,N_809,N_948);
and U1510 (N_1510,N_801,N_571);
xnor U1511 (N_1511,N_740,N_651);
and U1512 (N_1512,N_488,N_552);
nand U1513 (N_1513,N_902,N_225);
nand U1514 (N_1514,N_809,N_678);
nor U1515 (N_1515,N_40,N_397);
nor U1516 (N_1516,N_353,N_415);
nor U1517 (N_1517,N_188,N_366);
or U1518 (N_1518,N_331,N_180);
nand U1519 (N_1519,N_854,N_640);
or U1520 (N_1520,N_74,N_813);
nand U1521 (N_1521,N_453,N_626);
and U1522 (N_1522,N_337,N_29);
xor U1523 (N_1523,N_873,N_423);
or U1524 (N_1524,N_659,N_373);
nand U1525 (N_1525,N_795,N_394);
nor U1526 (N_1526,N_223,N_902);
xor U1527 (N_1527,N_273,N_206);
xnor U1528 (N_1528,N_670,N_260);
nor U1529 (N_1529,N_349,N_744);
and U1530 (N_1530,N_805,N_614);
or U1531 (N_1531,N_432,N_847);
nor U1532 (N_1532,N_117,N_670);
xor U1533 (N_1533,N_797,N_211);
and U1534 (N_1534,N_842,N_185);
and U1535 (N_1535,N_678,N_880);
and U1536 (N_1536,N_594,N_802);
xnor U1537 (N_1537,N_227,N_267);
nor U1538 (N_1538,N_132,N_441);
or U1539 (N_1539,N_909,N_239);
xor U1540 (N_1540,N_749,N_1);
nor U1541 (N_1541,N_751,N_671);
or U1542 (N_1542,N_8,N_124);
nand U1543 (N_1543,N_954,N_601);
xor U1544 (N_1544,N_921,N_285);
nor U1545 (N_1545,N_650,N_892);
xor U1546 (N_1546,N_952,N_126);
nor U1547 (N_1547,N_519,N_677);
nand U1548 (N_1548,N_316,N_646);
and U1549 (N_1549,N_859,N_751);
nor U1550 (N_1550,N_543,N_689);
and U1551 (N_1551,N_810,N_51);
nor U1552 (N_1552,N_684,N_659);
nand U1553 (N_1553,N_577,N_24);
nand U1554 (N_1554,N_933,N_468);
nor U1555 (N_1555,N_705,N_132);
and U1556 (N_1556,N_117,N_323);
nand U1557 (N_1557,N_32,N_574);
xor U1558 (N_1558,N_905,N_910);
nor U1559 (N_1559,N_274,N_263);
xor U1560 (N_1560,N_311,N_741);
or U1561 (N_1561,N_164,N_832);
or U1562 (N_1562,N_24,N_739);
nand U1563 (N_1563,N_971,N_696);
xor U1564 (N_1564,N_960,N_225);
or U1565 (N_1565,N_537,N_931);
and U1566 (N_1566,N_88,N_925);
nand U1567 (N_1567,N_915,N_289);
nand U1568 (N_1568,N_978,N_766);
xnor U1569 (N_1569,N_148,N_648);
or U1570 (N_1570,N_489,N_334);
xnor U1571 (N_1571,N_186,N_227);
xnor U1572 (N_1572,N_629,N_464);
xnor U1573 (N_1573,N_720,N_135);
xor U1574 (N_1574,N_149,N_101);
and U1575 (N_1575,N_26,N_949);
nor U1576 (N_1576,N_671,N_828);
xnor U1577 (N_1577,N_637,N_127);
and U1578 (N_1578,N_646,N_130);
or U1579 (N_1579,N_499,N_550);
xnor U1580 (N_1580,N_179,N_214);
xor U1581 (N_1581,N_12,N_765);
or U1582 (N_1582,N_314,N_121);
and U1583 (N_1583,N_672,N_191);
and U1584 (N_1584,N_547,N_629);
or U1585 (N_1585,N_344,N_398);
or U1586 (N_1586,N_676,N_104);
xor U1587 (N_1587,N_588,N_756);
or U1588 (N_1588,N_715,N_780);
xor U1589 (N_1589,N_603,N_266);
and U1590 (N_1590,N_725,N_759);
and U1591 (N_1591,N_817,N_497);
xor U1592 (N_1592,N_325,N_289);
or U1593 (N_1593,N_443,N_877);
and U1594 (N_1594,N_30,N_365);
or U1595 (N_1595,N_882,N_393);
and U1596 (N_1596,N_21,N_655);
or U1597 (N_1597,N_625,N_449);
nand U1598 (N_1598,N_404,N_278);
xor U1599 (N_1599,N_613,N_281);
nor U1600 (N_1600,N_372,N_336);
xnor U1601 (N_1601,N_175,N_387);
xor U1602 (N_1602,N_614,N_134);
or U1603 (N_1603,N_497,N_228);
and U1604 (N_1604,N_312,N_943);
nand U1605 (N_1605,N_554,N_841);
nor U1606 (N_1606,N_455,N_662);
or U1607 (N_1607,N_211,N_546);
nor U1608 (N_1608,N_638,N_817);
and U1609 (N_1609,N_487,N_995);
or U1610 (N_1610,N_194,N_996);
or U1611 (N_1611,N_647,N_522);
nand U1612 (N_1612,N_193,N_526);
and U1613 (N_1613,N_477,N_843);
and U1614 (N_1614,N_141,N_520);
or U1615 (N_1615,N_109,N_714);
nor U1616 (N_1616,N_815,N_676);
xnor U1617 (N_1617,N_300,N_345);
xor U1618 (N_1618,N_65,N_109);
nor U1619 (N_1619,N_84,N_82);
and U1620 (N_1620,N_876,N_86);
nor U1621 (N_1621,N_667,N_565);
nor U1622 (N_1622,N_193,N_501);
nand U1623 (N_1623,N_77,N_917);
xnor U1624 (N_1624,N_741,N_184);
nor U1625 (N_1625,N_255,N_213);
xor U1626 (N_1626,N_837,N_657);
nor U1627 (N_1627,N_928,N_16);
and U1628 (N_1628,N_168,N_96);
xor U1629 (N_1629,N_328,N_803);
nand U1630 (N_1630,N_612,N_614);
or U1631 (N_1631,N_828,N_770);
nand U1632 (N_1632,N_772,N_736);
xor U1633 (N_1633,N_464,N_893);
xor U1634 (N_1634,N_72,N_419);
nand U1635 (N_1635,N_17,N_763);
or U1636 (N_1636,N_667,N_70);
and U1637 (N_1637,N_833,N_936);
or U1638 (N_1638,N_176,N_632);
nor U1639 (N_1639,N_249,N_454);
xnor U1640 (N_1640,N_285,N_179);
and U1641 (N_1641,N_738,N_541);
nor U1642 (N_1642,N_994,N_845);
nand U1643 (N_1643,N_18,N_47);
nor U1644 (N_1644,N_129,N_536);
and U1645 (N_1645,N_83,N_334);
nor U1646 (N_1646,N_887,N_800);
nor U1647 (N_1647,N_480,N_551);
nand U1648 (N_1648,N_957,N_92);
xnor U1649 (N_1649,N_635,N_813);
or U1650 (N_1650,N_582,N_276);
xnor U1651 (N_1651,N_18,N_890);
xnor U1652 (N_1652,N_633,N_367);
or U1653 (N_1653,N_854,N_155);
nand U1654 (N_1654,N_575,N_6);
or U1655 (N_1655,N_472,N_48);
and U1656 (N_1656,N_0,N_339);
nand U1657 (N_1657,N_951,N_133);
nor U1658 (N_1658,N_233,N_850);
or U1659 (N_1659,N_778,N_891);
and U1660 (N_1660,N_184,N_621);
xor U1661 (N_1661,N_139,N_685);
and U1662 (N_1662,N_919,N_670);
or U1663 (N_1663,N_239,N_514);
xnor U1664 (N_1664,N_808,N_872);
nor U1665 (N_1665,N_924,N_968);
xnor U1666 (N_1666,N_303,N_672);
and U1667 (N_1667,N_999,N_951);
nor U1668 (N_1668,N_368,N_73);
xnor U1669 (N_1669,N_626,N_481);
nand U1670 (N_1670,N_398,N_626);
or U1671 (N_1671,N_189,N_71);
or U1672 (N_1672,N_137,N_40);
or U1673 (N_1673,N_48,N_655);
nor U1674 (N_1674,N_127,N_743);
and U1675 (N_1675,N_180,N_569);
and U1676 (N_1676,N_375,N_140);
nand U1677 (N_1677,N_563,N_32);
nor U1678 (N_1678,N_338,N_484);
or U1679 (N_1679,N_140,N_128);
and U1680 (N_1680,N_670,N_525);
nand U1681 (N_1681,N_631,N_942);
xnor U1682 (N_1682,N_287,N_627);
nor U1683 (N_1683,N_358,N_762);
xor U1684 (N_1684,N_132,N_975);
nand U1685 (N_1685,N_738,N_359);
nand U1686 (N_1686,N_884,N_517);
nor U1687 (N_1687,N_29,N_368);
or U1688 (N_1688,N_422,N_138);
and U1689 (N_1689,N_145,N_277);
xnor U1690 (N_1690,N_916,N_50);
nor U1691 (N_1691,N_941,N_170);
nand U1692 (N_1692,N_866,N_0);
nor U1693 (N_1693,N_964,N_813);
xnor U1694 (N_1694,N_532,N_580);
nor U1695 (N_1695,N_697,N_474);
nand U1696 (N_1696,N_67,N_986);
and U1697 (N_1697,N_596,N_322);
or U1698 (N_1698,N_733,N_494);
or U1699 (N_1699,N_158,N_247);
xnor U1700 (N_1700,N_435,N_15);
or U1701 (N_1701,N_698,N_619);
or U1702 (N_1702,N_242,N_396);
nor U1703 (N_1703,N_137,N_305);
nand U1704 (N_1704,N_448,N_929);
nand U1705 (N_1705,N_862,N_144);
nand U1706 (N_1706,N_6,N_611);
and U1707 (N_1707,N_609,N_865);
or U1708 (N_1708,N_25,N_970);
or U1709 (N_1709,N_646,N_886);
and U1710 (N_1710,N_359,N_736);
and U1711 (N_1711,N_317,N_47);
xnor U1712 (N_1712,N_378,N_172);
or U1713 (N_1713,N_52,N_485);
xnor U1714 (N_1714,N_892,N_224);
nand U1715 (N_1715,N_38,N_302);
nor U1716 (N_1716,N_26,N_682);
nor U1717 (N_1717,N_203,N_532);
nand U1718 (N_1718,N_413,N_995);
xor U1719 (N_1719,N_282,N_50);
nor U1720 (N_1720,N_31,N_146);
or U1721 (N_1721,N_937,N_29);
and U1722 (N_1722,N_22,N_492);
or U1723 (N_1723,N_73,N_136);
nand U1724 (N_1724,N_533,N_15);
xnor U1725 (N_1725,N_496,N_511);
or U1726 (N_1726,N_23,N_997);
xnor U1727 (N_1727,N_682,N_133);
xor U1728 (N_1728,N_95,N_904);
or U1729 (N_1729,N_730,N_44);
or U1730 (N_1730,N_568,N_107);
nor U1731 (N_1731,N_684,N_498);
and U1732 (N_1732,N_582,N_59);
and U1733 (N_1733,N_478,N_391);
nand U1734 (N_1734,N_721,N_546);
nor U1735 (N_1735,N_741,N_940);
nor U1736 (N_1736,N_395,N_574);
nor U1737 (N_1737,N_650,N_700);
and U1738 (N_1738,N_771,N_549);
nor U1739 (N_1739,N_875,N_366);
xor U1740 (N_1740,N_273,N_229);
or U1741 (N_1741,N_821,N_894);
xnor U1742 (N_1742,N_369,N_342);
xnor U1743 (N_1743,N_98,N_115);
xnor U1744 (N_1744,N_857,N_276);
nand U1745 (N_1745,N_207,N_313);
xor U1746 (N_1746,N_809,N_534);
or U1747 (N_1747,N_466,N_738);
and U1748 (N_1748,N_138,N_181);
nor U1749 (N_1749,N_984,N_882);
nor U1750 (N_1750,N_506,N_765);
and U1751 (N_1751,N_834,N_297);
nand U1752 (N_1752,N_357,N_801);
nor U1753 (N_1753,N_497,N_74);
and U1754 (N_1754,N_503,N_366);
nand U1755 (N_1755,N_189,N_422);
xnor U1756 (N_1756,N_117,N_493);
xnor U1757 (N_1757,N_223,N_909);
nand U1758 (N_1758,N_346,N_432);
nor U1759 (N_1759,N_872,N_396);
or U1760 (N_1760,N_923,N_393);
or U1761 (N_1761,N_905,N_440);
nand U1762 (N_1762,N_665,N_515);
or U1763 (N_1763,N_213,N_849);
nand U1764 (N_1764,N_220,N_277);
or U1765 (N_1765,N_840,N_702);
or U1766 (N_1766,N_570,N_763);
and U1767 (N_1767,N_978,N_982);
nand U1768 (N_1768,N_489,N_868);
nand U1769 (N_1769,N_95,N_27);
nor U1770 (N_1770,N_231,N_632);
xor U1771 (N_1771,N_22,N_329);
nand U1772 (N_1772,N_820,N_884);
nor U1773 (N_1773,N_127,N_662);
or U1774 (N_1774,N_862,N_783);
or U1775 (N_1775,N_501,N_322);
and U1776 (N_1776,N_700,N_279);
xnor U1777 (N_1777,N_250,N_260);
nand U1778 (N_1778,N_719,N_167);
nor U1779 (N_1779,N_902,N_756);
xor U1780 (N_1780,N_750,N_682);
xor U1781 (N_1781,N_366,N_101);
or U1782 (N_1782,N_732,N_194);
nor U1783 (N_1783,N_928,N_188);
nand U1784 (N_1784,N_885,N_900);
nor U1785 (N_1785,N_914,N_320);
or U1786 (N_1786,N_671,N_680);
and U1787 (N_1787,N_995,N_196);
xor U1788 (N_1788,N_510,N_842);
or U1789 (N_1789,N_19,N_338);
xnor U1790 (N_1790,N_416,N_538);
nand U1791 (N_1791,N_273,N_739);
and U1792 (N_1792,N_807,N_148);
nor U1793 (N_1793,N_17,N_443);
xor U1794 (N_1794,N_355,N_582);
and U1795 (N_1795,N_80,N_520);
or U1796 (N_1796,N_212,N_284);
nor U1797 (N_1797,N_459,N_224);
and U1798 (N_1798,N_493,N_726);
or U1799 (N_1799,N_595,N_686);
and U1800 (N_1800,N_322,N_960);
xnor U1801 (N_1801,N_8,N_519);
nor U1802 (N_1802,N_420,N_72);
nor U1803 (N_1803,N_326,N_372);
and U1804 (N_1804,N_405,N_80);
xnor U1805 (N_1805,N_694,N_611);
and U1806 (N_1806,N_965,N_434);
or U1807 (N_1807,N_267,N_680);
xor U1808 (N_1808,N_175,N_483);
or U1809 (N_1809,N_810,N_266);
or U1810 (N_1810,N_24,N_804);
and U1811 (N_1811,N_539,N_431);
nor U1812 (N_1812,N_912,N_973);
and U1813 (N_1813,N_115,N_409);
nor U1814 (N_1814,N_296,N_399);
xor U1815 (N_1815,N_701,N_632);
nand U1816 (N_1816,N_753,N_670);
nand U1817 (N_1817,N_810,N_838);
nand U1818 (N_1818,N_409,N_429);
nand U1819 (N_1819,N_103,N_844);
xor U1820 (N_1820,N_739,N_73);
nor U1821 (N_1821,N_715,N_711);
xor U1822 (N_1822,N_518,N_594);
nor U1823 (N_1823,N_390,N_521);
nand U1824 (N_1824,N_949,N_356);
and U1825 (N_1825,N_671,N_316);
or U1826 (N_1826,N_127,N_709);
nand U1827 (N_1827,N_291,N_321);
or U1828 (N_1828,N_344,N_276);
nor U1829 (N_1829,N_739,N_523);
and U1830 (N_1830,N_209,N_499);
nand U1831 (N_1831,N_643,N_613);
xnor U1832 (N_1832,N_361,N_126);
and U1833 (N_1833,N_688,N_190);
nand U1834 (N_1834,N_403,N_653);
nand U1835 (N_1835,N_936,N_314);
nor U1836 (N_1836,N_648,N_577);
or U1837 (N_1837,N_217,N_224);
or U1838 (N_1838,N_319,N_622);
xnor U1839 (N_1839,N_449,N_626);
xnor U1840 (N_1840,N_672,N_603);
or U1841 (N_1841,N_893,N_144);
nor U1842 (N_1842,N_608,N_67);
nor U1843 (N_1843,N_641,N_358);
nand U1844 (N_1844,N_218,N_627);
and U1845 (N_1845,N_627,N_459);
nand U1846 (N_1846,N_486,N_801);
or U1847 (N_1847,N_307,N_489);
nand U1848 (N_1848,N_227,N_604);
nor U1849 (N_1849,N_43,N_105);
xnor U1850 (N_1850,N_587,N_832);
nand U1851 (N_1851,N_970,N_824);
xnor U1852 (N_1852,N_556,N_226);
nand U1853 (N_1853,N_580,N_275);
xnor U1854 (N_1854,N_491,N_479);
and U1855 (N_1855,N_393,N_591);
nor U1856 (N_1856,N_838,N_890);
xnor U1857 (N_1857,N_64,N_407);
nor U1858 (N_1858,N_3,N_434);
or U1859 (N_1859,N_115,N_469);
xnor U1860 (N_1860,N_960,N_684);
nand U1861 (N_1861,N_215,N_595);
nor U1862 (N_1862,N_296,N_978);
nand U1863 (N_1863,N_275,N_372);
nand U1864 (N_1864,N_42,N_225);
nor U1865 (N_1865,N_691,N_839);
or U1866 (N_1866,N_310,N_171);
or U1867 (N_1867,N_687,N_973);
or U1868 (N_1868,N_272,N_188);
nor U1869 (N_1869,N_234,N_355);
nand U1870 (N_1870,N_953,N_918);
xor U1871 (N_1871,N_337,N_505);
and U1872 (N_1872,N_512,N_377);
nor U1873 (N_1873,N_29,N_378);
or U1874 (N_1874,N_586,N_265);
xor U1875 (N_1875,N_48,N_477);
nor U1876 (N_1876,N_985,N_231);
and U1877 (N_1877,N_388,N_832);
and U1878 (N_1878,N_512,N_31);
and U1879 (N_1879,N_527,N_927);
or U1880 (N_1880,N_732,N_613);
nor U1881 (N_1881,N_208,N_367);
nor U1882 (N_1882,N_858,N_987);
or U1883 (N_1883,N_436,N_209);
nor U1884 (N_1884,N_166,N_198);
and U1885 (N_1885,N_917,N_436);
xnor U1886 (N_1886,N_948,N_22);
and U1887 (N_1887,N_20,N_667);
xor U1888 (N_1888,N_809,N_766);
xor U1889 (N_1889,N_981,N_767);
xor U1890 (N_1890,N_504,N_774);
nor U1891 (N_1891,N_755,N_947);
nor U1892 (N_1892,N_44,N_472);
nor U1893 (N_1893,N_937,N_738);
xnor U1894 (N_1894,N_90,N_543);
and U1895 (N_1895,N_710,N_369);
nor U1896 (N_1896,N_780,N_585);
or U1897 (N_1897,N_96,N_799);
nor U1898 (N_1898,N_878,N_463);
and U1899 (N_1899,N_923,N_189);
xor U1900 (N_1900,N_124,N_11);
or U1901 (N_1901,N_75,N_490);
or U1902 (N_1902,N_66,N_280);
xor U1903 (N_1903,N_952,N_76);
nor U1904 (N_1904,N_70,N_799);
or U1905 (N_1905,N_428,N_898);
xnor U1906 (N_1906,N_568,N_753);
nand U1907 (N_1907,N_299,N_998);
nor U1908 (N_1908,N_493,N_675);
or U1909 (N_1909,N_480,N_176);
or U1910 (N_1910,N_55,N_445);
and U1911 (N_1911,N_814,N_117);
and U1912 (N_1912,N_444,N_98);
or U1913 (N_1913,N_522,N_153);
nand U1914 (N_1914,N_308,N_515);
nor U1915 (N_1915,N_932,N_946);
and U1916 (N_1916,N_402,N_604);
and U1917 (N_1917,N_934,N_290);
nor U1918 (N_1918,N_248,N_768);
and U1919 (N_1919,N_746,N_224);
xnor U1920 (N_1920,N_452,N_442);
or U1921 (N_1921,N_296,N_571);
nor U1922 (N_1922,N_692,N_972);
nand U1923 (N_1923,N_662,N_839);
or U1924 (N_1924,N_822,N_995);
nor U1925 (N_1925,N_855,N_340);
or U1926 (N_1926,N_837,N_912);
or U1927 (N_1927,N_465,N_688);
or U1928 (N_1928,N_792,N_106);
or U1929 (N_1929,N_835,N_679);
nor U1930 (N_1930,N_648,N_44);
and U1931 (N_1931,N_428,N_88);
nor U1932 (N_1932,N_291,N_280);
nand U1933 (N_1933,N_937,N_502);
nand U1934 (N_1934,N_198,N_644);
or U1935 (N_1935,N_743,N_985);
and U1936 (N_1936,N_218,N_874);
and U1937 (N_1937,N_39,N_734);
or U1938 (N_1938,N_447,N_957);
nand U1939 (N_1939,N_326,N_812);
and U1940 (N_1940,N_624,N_557);
nor U1941 (N_1941,N_247,N_665);
xnor U1942 (N_1942,N_883,N_433);
xnor U1943 (N_1943,N_27,N_501);
and U1944 (N_1944,N_428,N_320);
or U1945 (N_1945,N_781,N_436);
and U1946 (N_1946,N_726,N_403);
or U1947 (N_1947,N_50,N_624);
nand U1948 (N_1948,N_402,N_605);
or U1949 (N_1949,N_510,N_87);
nor U1950 (N_1950,N_287,N_219);
xnor U1951 (N_1951,N_645,N_730);
nand U1952 (N_1952,N_848,N_825);
nor U1953 (N_1953,N_338,N_124);
nor U1954 (N_1954,N_256,N_317);
xor U1955 (N_1955,N_482,N_478);
nand U1956 (N_1956,N_362,N_898);
or U1957 (N_1957,N_260,N_785);
xnor U1958 (N_1958,N_326,N_520);
xnor U1959 (N_1959,N_10,N_232);
or U1960 (N_1960,N_685,N_174);
or U1961 (N_1961,N_259,N_366);
nand U1962 (N_1962,N_150,N_370);
nor U1963 (N_1963,N_905,N_60);
nand U1964 (N_1964,N_73,N_290);
or U1965 (N_1965,N_782,N_402);
xnor U1966 (N_1966,N_426,N_467);
nand U1967 (N_1967,N_935,N_672);
xor U1968 (N_1968,N_125,N_192);
nor U1969 (N_1969,N_86,N_345);
nand U1970 (N_1970,N_383,N_321);
nand U1971 (N_1971,N_80,N_582);
or U1972 (N_1972,N_666,N_479);
and U1973 (N_1973,N_962,N_160);
and U1974 (N_1974,N_932,N_423);
and U1975 (N_1975,N_471,N_638);
xnor U1976 (N_1976,N_775,N_465);
and U1977 (N_1977,N_705,N_232);
xnor U1978 (N_1978,N_62,N_991);
or U1979 (N_1979,N_186,N_213);
nor U1980 (N_1980,N_736,N_897);
xnor U1981 (N_1981,N_918,N_965);
xor U1982 (N_1982,N_593,N_275);
xor U1983 (N_1983,N_399,N_866);
nand U1984 (N_1984,N_54,N_779);
or U1985 (N_1985,N_111,N_427);
or U1986 (N_1986,N_843,N_333);
nand U1987 (N_1987,N_133,N_651);
nand U1988 (N_1988,N_961,N_807);
and U1989 (N_1989,N_146,N_282);
xor U1990 (N_1990,N_617,N_873);
nor U1991 (N_1991,N_139,N_521);
and U1992 (N_1992,N_472,N_828);
and U1993 (N_1993,N_63,N_268);
or U1994 (N_1994,N_279,N_907);
or U1995 (N_1995,N_308,N_306);
nor U1996 (N_1996,N_446,N_942);
xor U1997 (N_1997,N_322,N_731);
nand U1998 (N_1998,N_311,N_246);
nand U1999 (N_1999,N_189,N_610);
and U2000 (N_2000,N_1202,N_1739);
and U2001 (N_2001,N_1995,N_1776);
nand U2002 (N_2002,N_1966,N_1632);
and U2003 (N_2003,N_1023,N_1317);
and U2004 (N_2004,N_1914,N_1200);
and U2005 (N_2005,N_1439,N_1127);
nor U2006 (N_2006,N_1700,N_1828);
or U2007 (N_2007,N_1203,N_1495);
nand U2008 (N_2008,N_1989,N_1781);
nand U2009 (N_2009,N_1770,N_1189);
or U2010 (N_2010,N_1680,N_1937);
and U2011 (N_2011,N_1179,N_1606);
nor U2012 (N_2012,N_1983,N_1492);
nor U2013 (N_2013,N_1283,N_1244);
and U2014 (N_2014,N_1086,N_1126);
nor U2015 (N_2015,N_1480,N_1798);
xnor U2016 (N_2016,N_1663,N_1526);
nand U2017 (N_2017,N_1140,N_1326);
or U2018 (N_2018,N_1251,N_1953);
or U2019 (N_2019,N_1155,N_1794);
nor U2020 (N_2020,N_1684,N_1404);
and U2021 (N_2021,N_1812,N_1925);
or U2022 (N_2022,N_1911,N_1508);
or U2023 (N_2023,N_1182,N_1012);
xnor U2024 (N_2024,N_1305,N_1751);
nor U2025 (N_2025,N_1912,N_1071);
nor U2026 (N_2026,N_1947,N_1855);
and U2027 (N_2027,N_1981,N_1138);
xor U2028 (N_2028,N_1550,N_1698);
and U2029 (N_2029,N_1859,N_1790);
or U2030 (N_2030,N_1627,N_1758);
or U2031 (N_2031,N_1481,N_1585);
nand U2032 (N_2032,N_1486,N_1544);
xor U2033 (N_2033,N_1059,N_1458);
and U2034 (N_2034,N_1690,N_1729);
nand U2035 (N_2035,N_1494,N_1287);
xor U2036 (N_2036,N_1027,N_1873);
xor U2037 (N_2037,N_1341,N_1659);
or U2038 (N_2038,N_1493,N_1269);
nand U2039 (N_2039,N_1637,N_1805);
or U2040 (N_2040,N_1516,N_1788);
nor U2041 (N_2041,N_1377,N_1471);
nor U2042 (N_2042,N_1276,N_1513);
nor U2043 (N_2043,N_1025,N_1594);
or U2044 (N_2044,N_1675,N_1514);
xor U2045 (N_2045,N_1384,N_1730);
nand U2046 (N_2046,N_1157,N_1304);
nor U2047 (N_2047,N_1357,N_1642);
xnor U2048 (N_2048,N_1685,N_1498);
or U2049 (N_2049,N_1964,N_1372);
xnor U2050 (N_2050,N_1766,N_1451);
nand U2051 (N_2051,N_1863,N_1803);
xnor U2052 (N_2052,N_1406,N_1078);
xnor U2053 (N_2053,N_1978,N_1804);
nand U2054 (N_2054,N_1329,N_1191);
nor U2055 (N_2055,N_1418,N_1407);
nand U2056 (N_2056,N_1125,N_1009);
and U2057 (N_2057,N_1643,N_1576);
nor U2058 (N_2058,N_1166,N_1993);
xor U2059 (N_2059,N_1586,N_1614);
nor U2060 (N_2060,N_1882,N_1255);
xor U2061 (N_2061,N_1783,N_1742);
nor U2062 (N_2062,N_1216,N_1561);
nand U2063 (N_2063,N_1485,N_1262);
nor U2064 (N_2064,N_1535,N_1950);
nand U2065 (N_2065,N_1152,N_1218);
nor U2066 (N_2066,N_1633,N_1780);
nand U2067 (N_2067,N_1691,N_1162);
nor U2068 (N_2068,N_1253,N_1075);
nand U2069 (N_2069,N_1462,N_1967);
xnor U2070 (N_2070,N_1099,N_1907);
xnor U2071 (N_2071,N_1196,N_1610);
and U2072 (N_2072,N_1673,N_1667);
nand U2073 (N_2073,N_1006,N_1677);
nor U2074 (N_2074,N_1440,N_1817);
nor U2075 (N_2075,N_1625,N_1823);
or U2076 (N_2076,N_1844,N_1135);
or U2077 (N_2077,N_1419,N_1399);
nor U2078 (N_2078,N_1756,N_1646);
xnor U2079 (N_2079,N_1603,N_1593);
nor U2080 (N_2080,N_1024,N_1866);
nor U2081 (N_2081,N_1497,N_1917);
and U2082 (N_2082,N_1104,N_1233);
and U2083 (N_2083,N_1749,N_1062);
nand U2084 (N_2084,N_1592,N_1300);
nor U2085 (N_2085,N_1861,N_1611);
and U2086 (N_2086,N_1306,N_1320);
nor U2087 (N_2087,N_1987,N_1521);
and U2088 (N_2088,N_1323,N_1076);
or U2089 (N_2089,N_1132,N_1052);
xor U2090 (N_2090,N_1327,N_1468);
and U2091 (N_2091,N_1734,N_1797);
or U2092 (N_2092,N_1792,N_1778);
and U2093 (N_2093,N_1807,N_1137);
nand U2094 (N_2094,N_1892,N_1999);
and U2095 (N_2095,N_1414,N_1428);
xnor U2096 (N_2096,N_1392,N_1924);
or U2097 (N_2097,N_1904,N_1957);
and U2098 (N_2098,N_1029,N_1156);
or U2099 (N_2099,N_1442,N_1353);
and U2100 (N_2100,N_1768,N_1648);
and U2101 (N_2101,N_1187,N_1765);
nor U2102 (N_2102,N_1026,N_1204);
nor U2103 (N_2103,N_1374,N_1644);
xnor U2104 (N_2104,N_1965,N_1281);
xor U2105 (N_2105,N_1296,N_1650);
and U2106 (N_2106,N_1932,N_1895);
or U2107 (N_2107,N_1032,N_1990);
and U2108 (N_2108,N_1148,N_1877);
and U2109 (N_2109,N_1149,N_1120);
xnor U2110 (N_2110,N_1901,N_1411);
nor U2111 (N_2111,N_1186,N_1049);
xnor U2112 (N_2112,N_1194,N_1446);
nor U2113 (N_2113,N_1097,N_1040);
xnor U2114 (N_2114,N_1867,N_1813);
xor U2115 (N_2115,N_1985,N_1755);
and U2116 (N_2116,N_1143,N_1369);
xor U2117 (N_2117,N_1332,N_1333);
or U2118 (N_2118,N_1284,N_1915);
nand U2119 (N_2119,N_1034,N_1266);
xnor U2120 (N_2120,N_1010,N_1299);
nor U2121 (N_2121,N_1031,N_1821);
nand U2122 (N_2122,N_1172,N_1436);
nand U2123 (N_2123,N_1786,N_1397);
or U2124 (N_2124,N_1998,N_1686);
and U2125 (N_2125,N_1709,N_1146);
xor U2126 (N_2126,N_1130,N_1519);
nand U2127 (N_2127,N_1112,N_1587);
and U2128 (N_2128,N_1349,N_1619);
xnor U2129 (N_2129,N_1242,N_1295);
and U2130 (N_2130,N_1081,N_1158);
and U2131 (N_2131,N_1342,N_1389);
and U2132 (N_2132,N_1772,N_1575);
nand U2133 (N_2133,N_1115,N_1209);
xnor U2134 (N_2134,N_1843,N_1634);
xor U2135 (N_2135,N_1558,N_1356);
or U2136 (N_2136,N_1976,N_1618);
nor U2137 (N_2137,N_1640,N_1687);
nor U2138 (N_2138,N_1628,N_1896);
nor U2139 (N_2139,N_1929,N_1580);
or U2140 (N_2140,N_1973,N_1566);
nand U2141 (N_2141,N_1702,N_1394);
nor U2142 (N_2142,N_1703,N_1744);
xnor U2143 (N_2143,N_1609,N_1482);
nor U2144 (N_2144,N_1565,N_1583);
xor U2145 (N_2145,N_1588,N_1693);
and U2146 (N_2146,N_1910,N_1825);
xor U2147 (N_2147,N_1762,N_1641);
xor U2148 (N_2148,N_1154,N_1551);
xor U2149 (N_2149,N_1639,N_1651);
and U2150 (N_2150,N_1815,N_1229);
nor U2151 (N_2151,N_1236,N_1211);
nand U2152 (N_2152,N_1946,N_1017);
nand U2153 (N_2153,N_1883,N_1291);
nand U2154 (N_2154,N_1933,N_1653);
or U2155 (N_2155,N_1941,N_1980);
nor U2156 (N_2156,N_1908,N_1810);
and U2157 (N_2157,N_1952,N_1072);
nor U2158 (N_2158,N_1534,N_1227);
or U2159 (N_2159,N_1197,N_1920);
nand U2160 (N_2160,N_1692,N_1832);
or U2161 (N_2161,N_1316,N_1248);
and U2162 (N_2162,N_1100,N_1145);
nand U2163 (N_2163,N_1708,N_1909);
and U2164 (N_2164,N_1022,N_1752);
and U2165 (N_2165,N_1678,N_1977);
and U2166 (N_2166,N_1577,N_1930);
nand U2167 (N_2167,N_1718,N_1199);
xor U2168 (N_2168,N_1288,N_1180);
nor U2169 (N_2169,N_1707,N_1490);
or U2170 (N_2170,N_1533,N_1169);
or U2171 (N_2171,N_1556,N_1874);
nor U2172 (N_2172,N_1122,N_1626);
or U2173 (N_2173,N_1705,N_1385);
nor U2174 (N_2174,N_1721,N_1339);
nand U2175 (N_2175,N_1310,N_1465);
nand U2176 (N_2176,N_1164,N_1613);
nor U2177 (N_2177,N_1808,N_1740);
and U2178 (N_2178,N_1717,N_1694);
nor U2179 (N_2179,N_1363,N_1738);
or U2180 (N_2180,N_1129,N_1567);
nor U2181 (N_2181,N_1880,N_1923);
and U2182 (N_2182,N_1105,N_1171);
or U2183 (N_2183,N_1258,N_1000);
or U2184 (N_2184,N_1728,N_1053);
xor U2185 (N_2185,N_1117,N_1926);
xnor U2186 (N_2186,N_1102,N_1715);
nor U2187 (N_2187,N_1390,N_1144);
nand U2188 (N_2188,N_1972,N_1777);
xor U2189 (N_2189,N_1150,N_1015);
xor U2190 (N_2190,N_1789,N_1979);
xor U2191 (N_2191,N_1520,N_1417);
nor U2192 (N_2192,N_1210,N_1589);
and U2193 (N_2193,N_1224,N_1898);
nand U2194 (N_2194,N_1019,N_1857);
and U2195 (N_2195,N_1506,N_1991);
and U2196 (N_2196,N_1886,N_1225);
xnor U2197 (N_2197,N_1077,N_1970);
xnor U2198 (N_2198,N_1563,N_1185);
and U2199 (N_2199,N_1597,N_1038);
or U2200 (N_2200,N_1699,N_1340);
nor U2201 (N_2201,N_1381,N_1934);
nand U2202 (N_2202,N_1870,N_1540);
or U2203 (N_2203,N_1106,N_1652);
and U2204 (N_2204,N_1261,N_1278);
or U2205 (N_2205,N_1927,N_1095);
and U2206 (N_2206,N_1775,N_1615);
nand U2207 (N_2207,N_1885,N_1665);
and U2208 (N_2208,N_1443,N_1359);
nand U2209 (N_2209,N_1101,N_1219);
nor U2210 (N_2210,N_1975,N_1552);
nand U2211 (N_2211,N_1878,N_1959);
and U2212 (N_2212,N_1386,N_1163);
nand U2213 (N_2213,N_1664,N_1512);
or U2214 (N_2214,N_1726,N_1467);
or U2215 (N_2215,N_1065,N_1669);
nand U2216 (N_2216,N_1461,N_1475);
and U2217 (N_2217,N_1711,N_1568);
or U2218 (N_2218,N_1846,N_1408);
or U2219 (N_2219,N_1319,N_1396);
nand U2220 (N_2220,N_1884,N_1887);
xnor U2221 (N_2221,N_1335,N_1502);
or U2222 (N_2222,N_1548,N_1916);
nand U2223 (N_2223,N_1159,N_1437);
or U2224 (N_2224,N_1827,N_1949);
xnor U2225 (N_2225,N_1388,N_1134);
nand U2226 (N_2226,N_1982,N_1324);
nand U2227 (N_2227,N_1487,N_1352);
and U2228 (N_2228,N_1367,N_1271);
nor U2229 (N_2229,N_1448,N_1259);
xnor U2230 (N_2230,N_1434,N_1221);
and U2231 (N_2231,N_1806,N_1572);
xor U2232 (N_2232,N_1286,N_1802);
nor U2233 (N_2233,N_1042,N_1060);
and U2234 (N_2234,N_1464,N_1936);
or U2235 (N_2235,N_1033,N_1379);
or U2236 (N_2236,N_1782,N_1181);
nand U2237 (N_2237,N_1541,N_1057);
and U2238 (N_2238,N_1315,N_1167);
nor U2239 (N_2239,N_1091,N_1234);
and U2240 (N_2240,N_1328,N_1165);
nand U2241 (N_2241,N_1141,N_1849);
or U2242 (N_2242,N_1838,N_1647);
or U2243 (N_2243,N_1064,N_1241);
nand U2244 (N_2244,N_1007,N_1674);
nand U2245 (N_2245,N_1013,N_1268);
nand U2246 (N_2246,N_1226,N_1252);
and U2247 (N_2247,N_1562,N_1198);
xor U2248 (N_2248,N_1212,N_1139);
and U2249 (N_2249,N_1491,N_1472);
or U2250 (N_2250,N_1265,N_1507);
xor U2251 (N_2251,N_1913,N_1517);
nor U2252 (N_2252,N_1837,N_1061);
xor U2253 (N_2253,N_1668,N_1899);
or U2254 (N_2254,N_1881,N_1463);
xor U2255 (N_2255,N_1872,N_1041);
nand U2256 (N_2256,N_1303,N_1621);
and U2257 (N_2257,N_1871,N_1438);
or U2258 (N_2258,N_1530,N_1596);
and U2259 (N_2259,N_1293,N_1488);
nor U2260 (N_2260,N_1956,N_1791);
or U2261 (N_2261,N_1160,N_1661);
nor U2262 (N_2262,N_1347,N_1719);
nor U2263 (N_2263,N_1282,N_1174);
and U2264 (N_2264,N_1409,N_1249);
nand U2265 (N_2265,N_1853,N_1918);
or U2266 (N_2266,N_1107,N_1215);
or U2267 (N_2267,N_1955,N_1662);
or U2268 (N_2268,N_1733,N_1831);
nor U2269 (N_2269,N_1176,N_1503);
xnor U2270 (N_2270,N_1168,N_1570);
or U2271 (N_2271,N_1745,N_1222);
or U2272 (N_2272,N_1787,N_1205);
and U2273 (N_2273,N_1795,N_1084);
or U2274 (N_2274,N_1444,N_1054);
nor U2275 (N_2275,N_1591,N_1852);
and U2276 (N_2276,N_1557,N_1869);
xnor U2277 (N_2277,N_1931,N_1764);
and U2278 (N_2278,N_1048,N_1943);
xnor U2279 (N_2279,N_1193,N_1454);
or U2280 (N_2280,N_1645,N_1090);
nor U2281 (N_2281,N_1584,N_1903);
nand U2282 (N_2282,N_1096,N_1935);
nor U2283 (N_2283,N_1243,N_1254);
nor U2284 (N_2284,N_1312,N_1759);
nor U2285 (N_2285,N_1047,N_1539);
or U2286 (N_2286,N_1500,N_1043);
or U2287 (N_2287,N_1582,N_1522);
or U2288 (N_2288,N_1382,N_1456);
and U2289 (N_2289,N_1416,N_1706);
nand U2290 (N_2290,N_1429,N_1747);
or U2291 (N_2291,N_1771,N_1875);
xor U2292 (N_2292,N_1401,N_1037);
or U2293 (N_2293,N_1161,N_1368);
or U2294 (N_2294,N_1239,N_1942);
nand U2295 (N_2295,N_1525,N_1400);
or U2296 (N_2296,N_1532,N_1051);
or U2297 (N_2297,N_1969,N_1876);
nand U2298 (N_2298,N_1536,N_1919);
or U2299 (N_2299,N_1631,N_1004);
nor U2300 (N_2300,N_1608,N_1297);
and U2301 (N_2301,N_1748,N_1554);
nand U2302 (N_2302,N_1195,N_1238);
and U2303 (N_2303,N_1842,N_1681);
nand U2304 (N_2304,N_1961,N_1449);
or U2305 (N_2305,N_1649,N_1689);
or U2306 (N_2306,N_1088,N_1799);
nand U2307 (N_2307,N_1063,N_1206);
xor U2308 (N_2308,N_1214,N_1131);
or U2309 (N_2309,N_1067,N_1109);
nand U2310 (N_2310,N_1779,N_1085);
or U2311 (N_2311,N_1294,N_1201);
nand U2312 (N_2312,N_1922,N_1793);
or U2313 (N_2313,N_1850,N_1499);
nor U2314 (N_2314,N_1579,N_1424);
and U2315 (N_2315,N_1289,N_1420);
nor U2316 (N_2316,N_1422,N_1476);
nand U2317 (N_2317,N_1002,N_1590);
xor U2318 (N_2318,N_1360,N_1055);
and U2319 (N_2319,N_1014,N_1380);
nand U2320 (N_2320,N_1290,N_1250);
nor U2321 (N_2321,N_1346,N_1058);
or U2322 (N_2322,N_1992,N_1403);
nand U2323 (N_2323,N_1720,N_1736);
nand U2324 (N_2324,N_1302,N_1398);
nand U2325 (N_2325,N_1345,N_1840);
or U2326 (N_2326,N_1655,N_1110);
or U2327 (N_2327,N_1361,N_1070);
xor U2328 (N_2328,N_1971,N_1116);
and U2329 (N_2329,N_1636,N_1879);
or U2330 (N_2330,N_1528,N_1858);
xnor U2331 (N_2331,N_1121,N_1724);
and U2332 (N_2332,N_1814,N_1905);
xor U2333 (N_2333,N_1028,N_1103);
or U2334 (N_2334,N_1108,N_1089);
nand U2335 (N_2335,N_1050,N_1604);
nor U2336 (N_2336,N_1030,N_1545);
and U2337 (N_2337,N_1093,N_1553);
nor U2338 (N_2338,N_1413,N_1713);
nand U2339 (N_2339,N_1834,N_1489);
and U2340 (N_2340,N_1314,N_1841);
nor U2341 (N_2341,N_1569,N_1046);
and U2342 (N_2342,N_1509,N_1761);
xnor U2343 (N_2343,N_1263,N_1391);
nor U2344 (N_2344,N_1954,N_1722);
or U2345 (N_2345,N_1123,N_1426);
nand U2346 (N_2346,N_1602,N_1275);
or U2347 (N_2347,N_1183,N_1737);
nand U2348 (N_2348,N_1524,N_1811);
xnor U2349 (N_2349,N_1240,N_1018);
or U2350 (N_2350,N_1743,N_1723);
nor U2351 (N_2351,N_1547,N_1245);
or U2352 (N_2352,N_1231,N_1003);
nor U2353 (N_2353,N_1331,N_1405);
nand U2354 (N_2354,N_1616,N_1839);
or U2355 (N_2355,N_1321,N_1682);
nor U2356 (N_2356,N_1410,N_1546);
xnor U2357 (N_2357,N_1732,N_1036);
xnor U2358 (N_2358,N_1620,N_1450);
nor U2359 (N_2359,N_1531,N_1460);
nand U2360 (N_2360,N_1940,N_1994);
or U2361 (N_2361,N_1432,N_1988);
nand U2362 (N_2362,N_1835,N_1082);
or U2363 (N_2363,N_1868,N_1505);
or U2364 (N_2364,N_1270,N_1119);
or U2365 (N_2365,N_1617,N_1826);
nor U2366 (N_2366,N_1845,N_1383);
nor U2367 (N_2367,N_1336,N_1478);
or U2368 (N_2368,N_1773,N_1153);
or U2369 (N_2369,N_1020,N_1453);
nand U2370 (N_2370,N_1555,N_1571);
xor U2371 (N_2371,N_1848,N_1601);
and U2372 (N_2372,N_1725,N_1769);
xor U2373 (N_2373,N_1371,N_1069);
or U2374 (N_2374,N_1011,N_1754);
nor U2375 (N_2375,N_1595,N_1142);
or U2376 (N_2376,N_1986,N_1862);
and U2377 (N_2377,N_1433,N_1133);
nand U2378 (N_2378,N_1607,N_1308);
nor U2379 (N_2379,N_1656,N_1113);
or U2380 (N_2380,N_1688,N_1948);
or U2381 (N_2381,N_1044,N_1958);
and U2382 (N_2382,N_1274,N_1763);
nand U2383 (N_2383,N_1466,N_1860);
nor U2384 (N_2384,N_1441,N_1318);
nor U2385 (N_2385,N_1136,N_1474);
nand U2386 (N_2386,N_1889,N_1629);
nor U2387 (N_2387,N_1056,N_1151);
or U2388 (N_2388,N_1549,N_1175);
and U2389 (N_2389,N_1395,N_1247);
or U2390 (N_2390,N_1622,N_1573);
nand U2391 (N_2391,N_1753,N_1897);
nor U2392 (N_2392,N_1430,N_1537);
nor U2393 (N_2393,N_1350,N_1750);
nand U2394 (N_2394,N_1996,N_1035);
nor U2395 (N_2395,N_1272,N_1114);
xnor U2396 (N_2396,N_1727,N_1230);
or U2397 (N_2397,N_1279,N_1496);
xnor U2398 (N_2398,N_1358,N_1008);
nand U2399 (N_2399,N_1654,N_1818);
nand U2400 (N_2400,N_1459,N_1301);
and U2401 (N_2401,N_1260,N_1370);
xor U2402 (N_2402,N_1173,N_1757);
xnor U2403 (N_2403,N_1307,N_1188);
nand U2404 (N_2404,N_1455,N_1731);
nand U2405 (N_2405,N_1170,N_1423);
nand U2406 (N_2406,N_1376,N_1425);
nor U2407 (N_2407,N_1962,N_1984);
nor U2408 (N_2408,N_1974,N_1068);
nand U2409 (N_2409,N_1285,N_1894);
nor U2410 (N_2410,N_1313,N_1623);
or U2411 (N_2411,N_1264,N_1111);
nor U2412 (N_2412,N_1311,N_1638);
and U2413 (N_2413,N_1348,N_1473);
or U2414 (N_2414,N_1147,N_1208);
or U2415 (N_2415,N_1670,N_1207);
nor U2416 (N_2416,N_1256,N_1900);
nor U2417 (N_2417,N_1518,N_1073);
nor U2418 (N_2418,N_1944,N_1469);
nand U2419 (N_2419,N_1847,N_1819);
nor U2420 (N_2420,N_1362,N_1504);
xor U2421 (N_2421,N_1128,N_1666);
and U2422 (N_2422,N_1774,N_1343);
or U2423 (N_2423,N_1511,N_1671);
or U2424 (N_2424,N_1672,N_1581);
xor U2425 (N_2425,N_1267,N_1351);
and U2426 (N_2426,N_1337,N_1564);
and U2427 (N_2427,N_1767,N_1997);
nor U2428 (N_2428,N_1016,N_1893);
xor U2429 (N_2429,N_1373,N_1741);
or U2430 (N_2430,N_1630,N_1083);
or U2431 (N_2431,N_1710,N_1366);
and U2432 (N_2432,N_1298,N_1080);
and U2433 (N_2433,N_1612,N_1246);
nor U2434 (N_2434,N_1829,N_1697);
nor U2435 (N_2435,N_1412,N_1824);
nor U2436 (N_2436,N_1683,N_1542);
or U2437 (N_2437,N_1421,N_1960);
nor U2438 (N_2438,N_1074,N_1851);
and U2439 (N_2439,N_1830,N_1220);
or U2440 (N_2440,N_1746,N_1635);
nand U2441 (N_2441,N_1510,N_1235);
or U2442 (N_2442,N_1325,N_1696);
or U2443 (N_2443,N_1445,N_1477);
nor U2444 (N_2444,N_1714,N_1001);
nor U2445 (N_2445,N_1599,N_1079);
nor U2446 (N_2446,N_1538,N_1322);
and U2447 (N_2447,N_1796,N_1387);
xor U2448 (N_2448,N_1515,N_1330);
or U2449 (N_2449,N_1816,N_1760);
and U2450 (N_2450,N_1177,N_1273);
nor U2451 (N_2451,N_1005,N_1701);
or U2452 (N_2452,N_1415,N_1213);
xor U2453 (N_2453,N_1543,N_1364);
nor U2454 (N_2454,N_1921,N_1560);
nand U2455 (N_2455,N_1968,N_1232);
nand U2456 (N_2456,N_1679,N_1178);
xnor U2457 (N_2457,N_1484,N_1735);
and U2458 (N_2458,N_1906,N_1605);
xnor U2459 (N_2459,N_1292,N_1431);
nand U2460 (N_2460,N_1427,N_1470);
xnor U2461 (N_2461,N_1021,N_1864);
nand U2462 (N_2462,N_1452,N_1228);
and U2463 (N_2463,N_1658,N_1865);
xor U2464 (N_2464,N_1820,N_1624);
or U2465 (N_2465,N_1704,N_1822);
and U2466 (N_2466,N_1523,N_1712);
nor U2467 (N_2467,N_1217,N_1716);
and U2468 (N_2468,N_1280,N_1365);
xnor U2469 (N_2469,N_1598,N_1574);
and U2470 (N_2470,N_1257,N_1277);
nor U2471 (N_2471,N_1695,N_1527);
nor U2472 (N_2472,N_1784,N_1833);
and U2473 (N_2473,N_1939,N_1928);
xnor U2474 (N_2474,N_1902,N_1501);
nor U2475 (N_2475,N_1338,N_1891);
and U2476 (N_2476,N_1856,N_1354);
and U2477 (N_2477,N_1529,N_1355);
and U2478 (N_2478,N_1092,N_1963);
nor U2479 (N_2479,N_1836,N_1190);
nor U2480 (N_2480,N_1660,N_1801);
nand U2481 (N_2481,N_1066,N_1483);
xor U2482 (N_2482,N_1098,N_1559);
or U2483 (N_2483,N_1809,N_1785);
xnor U2484 (N_2484,N_1334,N_1854);
nor U2485 (N_2485,N_1039,N_1435);
or U2486 (N_2486,N_1951,N_1888);
nand U2487 (N_2487,N_1890,N_1309);
nor U2488 (N_2488,N_1578,N_1237);
xor U2489 (N_2489,N_1378,N_1938);
xnor U2490 (N_2490,N_1447,N_1375);
or U2491 (N_2491,N_1118,N_1676);
xor U2492 (N_2492,N_1457,N_1600);
xor U2493 (N_2493,N_1124,N_1945);
nor U2494 (N_2494,N_1657,N_1479);
nor U2495 (N_2495,N_1393,N_1344);
nand U2496 (N_2496,N_1223,N_1184);
xnor U2497 (N_2497,N_1402,N_1192);
nand U2498 (N_2498,N_1087,N_1094);
and U2499 (N_2499,N_1045,N_1800);
nand U2500 (N_2500,N_1003,N_1059);
and U2501 (N_2501,N_1352,N_1296);
xnor U2502 (N_2502,N_1035,N_1907);
nor U2503 (N_2503,N_1501,N_1598);
or U2504 (N_2504,N_1597,N_1604);
xor U2505 (N_2505,N_1771,N_1717);
or U2506 (N_2506,N_1120,N_1903);
and U2507 (N_2507,N_1741,N_1525);
and U2508 (N_2508,N_1984,N_1934);
xnor U2509 (N_2509,N_1304,N_1364);
nor U2510 (N_2510,N_1595,N_1206);
and U2511 (N_2511,N_1428,N_1765);
nor U2512 (N_2512,N_1204,N_1887);
or U2513 (N_2513,N_1548,N_1033);
and U2514 (N_2514,N_1288,N_1306);
xnor U2515 (N_2515,N_1419,N_1855);
or U2516 (N_2516,N_1670,N_1764);
nor U2517 (N_2517,N_1500,N_1818);
nor U2518 (N_2518,N_1297,N_1894);
and U2519 (N_2519,N_1470,N_1938);
or U2520 (N_2520,N_1018,N_1248);
or U2521 (N_2521,N_1956,N_1001);
or U2522 (N_2522,N_1846,N_1935);
and U2523 (N_2523,N_1744,N_1005);
or U2524 (N_2524,N_1548,N_1268);
and U2525 (N_2525,N_1976,N_1400);
or U2526 (N_2526,N_1164,N_1239);
and U2527 (N_2527,N_1566,N_1933);
xor U2528 (N_2528,N_1740,N_1637);
or U2529 (N_2529,N_1243,N_1492);
nand U2530 (N_2530,N_1561,N_1300);
and U2531 (N_2531,N_1493,N_1743);
nor U2532 (N_2532,N_1674,N_1491);
nand U2533 (N_2533,N_1040,N_1536);
nor U2534 (N_2534,N_1921,N_1384);
nor U2535 (N_2535,N_1422,N_1361);
nand U2536 (N_2536,N_1714,N_1212);
and U2537 (N_2537,N_1512,N_1106);
nand U2538 (N_2538,N_1163,N_1243);
xnor U2539 (N_2539,N_1241,N_1352);
nor U2540 (N_2540,N_1626,N_1875);
nand U2541 (N_2541,N_1153,N_1548);
xor U2542 (N_2542,N_1318,N_1491);
nor U2543 (N_2543,N_1979,N_1049);
or U2544 (N_2544,N_1655,N_1963);
nor U2545 (N_2545,N_1941,N_1435);
nor U2546 (N_2546,N_1235,N_1023);
xnor U2547 (N_2547,N_1840,N_1616);
nand U2548 (N_2548,N_1263,N_1865);
nand U2549 (N_2549,N_1396,N_1562);
nor U2550 (N_2550,N_1777,N_1673);
nand U2551 (N_2551,N_1994,N_1508);
nand U2552 (N_2552,N_1235,N_1232);
and U2553 (N_2553,N_1748,N_1822);
xor U2554 (N_2554,N_1127,N_1586);
nor U2555 (N_2555,N_1372,N_1475);
or U2556 (N_2556,N_1319,N_1142);
nand U2557 (N_2557,N_1295,N_1096);
nor U2558 (N_2558,N_1906,N_1473);
nand U2559 (N_2559,N_1980,N_1309);
or U2560 (N_2560,N_1188,N_1636);
nand U2561 (N_2561,N_1953,N_1724);
or U2562 (N_2562,N_1428,N_1028);
nand U2563 (N_2563,N_1508,N_1081);
nor U2564 (N_2564,N_1974,N_1118);
xor U2565 (N_2565,N_1779,N_1569);
and U2566 (N_2566,N_1865,N_1214);
nor U2567 (N_2567,N_1823,N_1238);
nand U2568 (N_2568,N_1846,N_1003);
and U2569 (N_2569,N_1937,N_1138);
nor U2570 (N_2570,N_1146,N_1406);
nand U2571 (N_2571,N_1795,N_1378);
or U2572 (N_2572,N_1714,N_1783);
and U2573 (N_2573,N_1355,N_1445);
and U2574 (N_2574,N_1907,N_1040);
or U2575 (N_2575,N_1070,N_1057);
and U2576 (N_2576,N_1706,N_1684);
xor U2577 (N_2577,N_1631,N_1121);
or U2578 (N_2578,N_1219,N_1706);
and U2579 (N_2579,N_1542,N_1032);
or U2580 (N_2580,N_1111,N_1529);
nor U2581 (N_2581,N_1247,N_1255);
xor U2582 (N_2582,N_1096,N_1560);
nand U2583 (N_2583,N_1013,N_1442);
nand U2584 (N_2584,N_1805,N_1793);
or U2585 (N_2585,N_1719,N_1597);
xor U2586 (N_2586,N_1728,N_1689);
or U2587 (N_2587,N_1857,N_1004);
or U2588 (N_2588,N_1288,N_1538);
nand U2589 (N_2589,N_1929,N_1176);
or U2590 (N_2590,N_1016,N_1845);
or U2591 (N_2591,N_1201,N_1267);
xnor U2592 (N_2592,N_1256,N_1184);
nand U2593 (N_2593,N_1030,N_1167);
nor U2594 (N_2594,N_1576,N_1899);
nand U2595 (N_2595,N_1763,N_1541);
and U2596 (N_2596,N_1266,N_1298);
or U2597 (N_2597,N_1653,N_1018);
nand U2598 (N_2598,N_1776,N_1366);
nor U2599 (N_2599,N_1772,N_1682);
or U2600 (N_2600,N_1139,N_1420);
xnor U2601 (N_2601,N_1844,N_1870);
nor U2602 (N_2602,N_1172,N_1922);
or U2603 (N_2603,N_1340,N_1827);
nand U2604 (N_2604,N_1611,N_1185);
and U2605 (N_2605,N_1176,N_1810);
or U2606 (N_2606,N_1755,N_1092);
nor U2607 (N_2607,N_1287,N_1222);
nand U2608 (N_2608,N_1672,N_1660);
or U2609 (N_2609,N_1682,N_1976);
or U2610 (N_2610,N_1545,N_1579);
nor U2611 (N_2611,N_1476,N_1298);
or U2612 (N_2612,N_1021,N_1840);
nor U2613 (N_2613,N_1029,N_1282);
nor U2614 (N_2614,N_1786,N_1623);
xor U2615 (N_2615,N_1729,N_1486);
nor U2616 (N_2616,N_1880,N_1577);
nor U2617 (N_2617,N_1742,N_1921);
nor U2618 (N_2618,N_1223,N_1857);
xnor U2619 (N_2619,N_1081,N_1406);
nand U2620 (N_2620,N_1509,N_1973);
nor U2621 (N_2621,N_1609,N_1649);
nand U2622 (N_2622,N_1323,N_1600);
nor U2623 (N_2623,N_1970,N_1870);
or U2624 (N_2624,N_1779,N_1831);
and U2625 (N_2625,N_1844,N_1204);
xor U2626 (N_2626,N_1519,N_1536);
xor U2627 (N_2627,N_1298,N_1064);
nor U2628 (N_2628,N_1679,N_1740);
nand U2629 (N_2629,N_1131,N_1951);
or U2630 (N_2630,N_1546,N_1720);
or U2631 (N_2631,N_1744,N_1082);
nor U2632 (N_2632,N_1453,N_1873);
and U2633 (N_2633,N_1969,N_1643);
and U2634 (N_2634,N_1560,N_1088);
nand U2635 (N_2635,N_1849,N_1298);
xor U2636 (N_2636,N_1670,N_1129);
and U2637 (N_2637,N_1337,N_1880);
xnor U2638 (N_2638,N_1282,N_1871);
nor U2639 (N_2639,N_1345,N_1852);
and U2640 (N_2640,N_1291,N_1661);
nor U2641 (N_2641,N_1943,N_1150);
nand U2642 (N_2642,N_1898,N_1105);
xnor U2643 (N_2643,N_1107,N_1922);
and U2644 (N_2644,N_1444,N_1767);
or U2645 (N_2645,N_1775,N_1950);
nor U2646 (N_2646,N_1241,N_1790);
and U2647 (N_2647,N_1447,N_1439);
xnor U2648 (N_2648,N_1479,N_1410);
nand U2649 (N_2649,N_1988,N_1486);
or U2650 (N_2650,N_1366,N_1902);
nand U2651 (N_2651,N_1689,N_1145);
nand U2652 (N_2652,N_1761,N_1558);
or U2653 (N_2653,N_1479,N_1769);
or U2654 (N_2654,N_1498,N_1129);
and U2655 (N_2655,N_1050,N_1802);
and U2656 (N_2656,N_1263,N_1196);
nor U2657 (N_2657,N_1034,N_1810);
or U2658 (N_2658,N_1308,N_1284);
nor U2659 (N_2659,N_1580,N_1709);
and U2660 (N_2660,N_1838,N_1047);
xnor U2661 (N_2661,N_1048,N_1042);
or U2662 (N_2662,N_1462,N_1914);
or U2663 (N_2663,N_1507,N_1168);
or U2664 (N_2664,N_1643,N_1649);
nor U2665 (N_2665,N_1329,N_1994);
or U2666 (N_2666,N_1552,N_1619);
or U2667 (N_2667,N_1140,N_1872);
and U2668 (N_2668,N_1530,N_1234);
xor U2669 (N_2669,N_1368,N_1402);
nand U2670 (N_2670,N_1551,N_1038);
nor U2671 (N_2671,N_1437,N_1158);
nor U2672 (N_2672,N_1760,N_1891);
nand U2673 (N_2673,N_1293,N_1322);
xnor U2674 (N_2674,N_1142,N_1588);
xnor U2675 (N_2675,N_1259,N_1904);
or U2676 (N_2676,N_1239,N_1555);
or U2677 (N_2677,N_1746,N_1222);
nand U2678 (N_2678,N_1210,N_1133);
xor U2679 (N_2679,N_1101,N_1001);
and U2680 (N_2680,N_1138,N_1870);
or U2681 (N_2681,N_1964,N_1485);
or U2682 (N_2682,N_1223,N_1409);
and U2683 (N_2683,N_1891,N_1227);
and U2684 (N_2684,N_1922,N_1516);
nor U2685 (N_2685,N_1500,N_1332);
or U2686 (N_2686,N_1759,N_1995);
or U2687 (N_2687,N_1335,N_1402);
or U2688 (N_2688,N_1754,N_1972);
nand U2689 (N_2689,N_1979,N_1368);
or U2690 (N_2690,N_1493,N_1366);
xor U2691 (N_2691,N_1546,N_1800);
or U2692 (N_2692,N_1912,N_1476);
nor U2693 (N_2693,N_1377,N_1038);
xnor U2694 (N_2694,N_1074,N_1056);
xor U2695 (N_2695,N_1531,N_1038);
or U2696 (N_2696,N_1906,N_1637);
nand U2697 (N_2697,N_1461,N_1764);
nand U2698 (N_2698,N_1350,N_1369);
nand U2699 (N_2699,N_1550,N_1567);
nand U2700 (N_2700,N_1079,N_1521);
or U2701 (N_2701,N_1015,N_1393);
and U2702 (N_2702,N_1704,N_1234);
nor U2703 (N_2703,N_1792,N_1994);
xnor U2704 (N_2704,N_1451,N_1264);
nor U2705 (N_2705,N_1006,N_1441);
nor U2706 (N_2706,N_1957,N_1821);
or U2707 (N_2707,N_1282,N_1122);
xor U2708 (N_2708,N_1930,N_1230);
nand U2709 (N_2709,N_1337,N_1356);
nor U2710 (N_2710,N_1473,N_1314);
xor U2711 (N_2711,N_1680,N_1333);
and U2712 (N_2712,N_1034,N_1444);
xnor U2713 (N_2713,N_1602,N_1953);
nand U2714 (N_2714,N_1531,N_1380);
nor U2715 (N_2715,N_1381,N_1929);
xnor U2716 (N_2716,N_1119,N_1100);
or U2717 (N_2717,N_1023,N_1804);
or U2718 (N_2718,N_1409,N_1778);
xnor U2719 (N_2719,N_1945,N_1307);
and U2720 (N_2720,N_1598,N_1119);
nor U2721 (N_2721,N_1583,N_1032);
and U2722 (N_2722,N_1644,N_1654);
nand U2723 (N_2723,N_1310,N_1831);
nand U2724 (N_2724,N_1443,N_1114);
and U2725 (N_2725,N_1834,N_1977);
nor U2726 (N_2726,N_1915,N_1875);
or U2727 (N_2727,N_1239,N_1207);
nand U2728 (N_2728,N_1622,N_1194);
nand U2729 (N_2729,N_1807,N_1558);
or U2730 (N_2730,N_1141,N_1957);
nor U2731 (N_2731,N_1532,N_1805);
xor U2732 (N_2732,N_1639,N_1190);
or U2733 (N_2733,N_1842,N_1926);
nand U2734 (N_2734,N_1784,N_1685);
nor U2735 (N_2735,N_1424,N_1800);
nand U2736 (N_2736,N_1126,N_1908);
nor U2737 (N_2737,N_1659,N_1391);
xnor U2738 (N_2738,N_1228,N_1914);
and U2739 (N_2739,N_1337,N_1037);
nor U2740 (N_2740,N_1505,N_1439);
and U2741 (N_2741,N_1000,N_1661);
and U2742 (N_2742,N_1740,N_1642);
or U2743 (N_2743,N_1707,N_1742);
and U2744 (N_2744,N_1325,N_1213);
nand U2745 (N_2745,N_1595,N_1984);
and U2746 (N_2746,N_1125,N_1611);
or U2747 (N_2747,N_1221,N_1165);
or U2748 (N_2748,N_1786,N_1193);
and U2749 (N_2749,N_1141,N_1362);
nor U2750 (N_2750,N_1763,N_1748);
xnor U2751 (N_2751,N_1880,N_1401);
and U2752 (N_2752,N_1278,N_1409);
and U2753 (N_2753,N_1871,N_1589);
or U2754 (N_2754,N_1309,N_1275);
xnor U2755 (N_2755,N_1669,N_1748);
or U2756 (N_2756,N_1070,N_1076);
or U2757 (N_2757,N_1258,N_1237);
or U2758 (N_2758,N_1205,N_1530);
nand U2759 (N_2759,N_1840,N_1516);
and U2760 (N_2760,N_1125,N_1059);
and U2761 (N_2761,N_1444,N_1754);
nor U2762 (N_2762,N_1864,N_1503);
or U2763 (N_2763,N_1806,N_1917);
or U2764 (N_2764,N_1848,N_1751);
nand U2765 (N_2765,N_1612,N_1398);
xnor U2766 (N_2766,N_1884,N_1520);
nand U2767 (N_2767,N_1370,N_1409);
nor U2768 (N_2768,N_1705,N_1927);
nand U2769 (N_2769,N_1522,N_1920);
nand U2770 (N_2770,N_1714,N_1389);
xnor U2771 (N_2771,N_1683,N_1952);
nand U2772 (N_2772,N_1133,N_1733);
xnor U2773 (N_2773,N_1801,N_1590);
xnor U2774 (N_2774,N_1734,N_1431);
nand U2775 (N_2775,N_1732,N_1359);
or U2776 (N_2776,N_1655,N_1354);
and U2777 (N_2777,N_1607,N_1547);
or U2778 (N_2778,N_1233,N_1467);
or U2779 (N_2779,N_1175,N_1883);
nor U2780 (N_2780,N_1820,N_1164);
xor U2781 (N_2781,N_1093,N_1904);
nand U2782 (N_2782,N_1606,N_1950);
and U2783 (N_2783,N_1422,N_1095);
nor U2784 (N_2784,N_1119,N_1787);
nand U2785 (N_2785,N_1394,N_1039);
xor U2786 (N_2786,N_1422,N_1972);
or U2787 (N_2787,N_1534,N_1654);
nor U2788 (N_2788,N_1070,N_1981);
and U2789 (N_2789,N_1489,N_1875);
xnor U2790 (N_2790,N_1079,N_1090);
and U2791 (N_2791,N_1361,N_1223);
nand U2792 (N_2792,N_1135,N_1940);
or U2793 (N_2793,N_1766,N_1636);
nand U2794 (N_2794,N_1888,N_1878);
xor U2795 (N_2795,N_1708,N_1684);
nor U2796 (N_2796,N_1456,N_1393);
and U2797 (N_2797,N_1010,N_1538);
and U2798 (N_2798,N_1044,N_1330);
nor U2799 (N_2799,N_1290,N_1821);
nand U2800 (N_2800,N_1395,N_1015);
nor U2801 (N_2801,N_1736,N_1978);
and U2802 (N_2802,N_1316,N_1198);
nor U2803 (N_2803,N_1726,N_1821);
nor U2804 (N_2804,N_1557,N_1289);
xor U2805 (N_2805,N_1765,N_1053);
xor U2806 (N_2806,N_1863,N_1241);
and U2807 (N_2807,N_1111,N_1184);
and U2808 (N_2808,N_1464,N_1435);
and U2809 (N_2809,N_1171,N_1304);
nand U2810 (N_2810,N_1409,N_1651);
or U2811 (N_2811,N_1331,N_1794);
nor U2812 (N_2812,N_1582,N_1128);
xor U2813 (N_2813,N_1266,N_1364);
nor U2814 (N_2814,N_1342,N_1028);
and U2815 (N_2815,N_1512,N_1451);
xor U2816 (N_2816,N_1990,N_1639);
and U2817 (N_2817,N_1839,N_1605);
nand U2818 (N_2818,N_1712,N_1144);
or U2819 (N_2819,N_1594,N_1962);
nand U2820 (N_2820,N_1093,N_1928);
and U2821 (N_2821,N_1088,N_1862);
xnor U2822 (N_2822,N_1867,N_1368);
nand U2823 (N_2823,N_1103,N_1451);
or U2824 (N_2824,N_1554,N_1302);
xnor U2825 (N_2825,N_1401,N_1855);
xor U2826 (N_2826,N_1565,N_1523);
nor U2827 (N_2827,N_1934,N_1655);
and U2828 (N_2828,N_1256,N_1629);
nor U2829 (N_2829,N_1957,N_1968);
or U2830 (N_2830,N_1649,N_1984);
nor U2831 (N_2831,N_1853,N_1155);
and U2832 (N_2832,N_1499,N_1177);
and U2833 (N_2833,N_1974,N_1871);
xor U2834 (N_2834,N_1322,N_1511);
and U2835 (N_2835,N_1760,N_1459);
or U2836 (N_2836,N_1706,N_1526);
and U2837 (N_2837,N_1182,N_1306);
and U2838 (N_2838,N_1098,N_1872);
or U2839 (N_2839,N_1163,N_1676);
and U2840 (N_2840,N_1910,N_1661);
and U2841 (N_2841,N_1914,N_1491);
nor U2842 (N_2842,N_1834,N_1684);
nor U2843 (N_2843,N_1432,N_1914);
nand U2844 (N_2844,N_1968,N_1358);
nand U2845 (N_2845,N_1671,N_1664);
nand U2846 (N_2846,N_1528,N_1636);
and U2847 (N_2847,N_1162,N_1258);
xor U2848 (N_2848,N_1498,N_1290);
and U2849 (N_2849,N_1049,N_1790);
and U2850 (N_2850,N_1457,N_1385);
and U2851 (N_2851,N_1117,N_1931);
nor U2852 (N_2852,N_1470,N_1576);
or U2853 (N_2853,N_1685,N_1451);
xor U2854 (N_2854,N_1884,N_1080);
xnor U2855 (N_2855,N_1240,N_1641);
xor U2856 (N_2856,N_1508,N_1525);
and U2857 (N_2857,N_1319,N_1489);
nor U2858 (N_2858,N_1215,N_1230);
nor U2859 (N_2859,N_1506,N_1894);
xor U2860 (N_2860,N_1754,N_1085);
and U2861 (N_2861,N_1077,N_1152);
nand U2862 (N_2862,N_1612,N_1147);
nand U2863 (N_2863,N_1134,N_1839);
or U2864 (N_2864,N_1896,N_1129);
nand U2865 (N_2865,N_1665,N_1084);
xor U2866 (N_2866,N_1114,N_1337);
xor U2867 (N_2867,N_1056,N_1439);
nand U2868 (N_2868,N_1293,N_1552);
or U2869 (N_2869,N_1715,N_1529);
nand U2870 (N_2870,N_1801,N_1667);
nor U2871 (N_2871,N_1971,N_1914);
nand U2872 (N_2872,N_1662,N_1102);
or U2873 (N_2873,N_1190,N_1172);
and U2874 (N_2874,N_1413,N_1266);
nor U2875 (N_2875,N_1074,N_1184);
nor U2876 (N_2876,N_1653,N_1931);
and U2877 (N_2877,N_1862,N_1315);
xnor U2878 (N_2878,N_1222,N_1062);
nand U2879 (N_2879,N_1465,N_1563);
and U2880 (N_2880,N_1225,N_1794);
and U2881 (N_2881,N_1194,N_1574);
and U2882 (N_2882,N_1387,N_1986);
nor U2883 (N_2883,N_1468,N_1329);
xor U2884 (N_2884,N_1895,N_1466);
nand U2885 (N_2885,N_1377,N_1046);
and U2886 (N_2886,N_1233,N_1002);
or U2887 (N_2887,N_1867,N_1937);
and U2888 (N_2888,N_1771,N_1822);
or U2889 (N_2889,N_1051,N_1899);
and U2890 (N_2890,N_1936,N_1034);
xnor U2891 (N_2891,N_1693,N_1093);
nand U2892 (N_2892,N_1315,N_1116);
or U2893 (N_2893,N_1811,N_1172);
xor U2894 (N_2894,N_1444,N_1518);
or U2895 (N_2895,N_1168,N_1370);
nor U2896 (N_2896,N_1897,N_1725);
xnor U2897 (N_2897,N_1039,N_1156);
xor U2898 (N_2898,N_1079,N_1833);
and U2899 (N_2899,N_1117,N_1205);
nand U2900 (N_2900,N_1532,N_1867);
nand U2901 (N_2901,N_1715,N_1580);
xor U2902 (N_2902,N_1948,N_1924);
and U2903 (N_2903,N_1557,N_1504);
or U2904 (N_2904,N_1717,N_1020);
nor U2905 (N_2905,N_1003,N_1700);
nand U2906 (N_2906,N_1899,N_1445);
or U2907 (N_2907,N_1876,N_1170);
xor U2908 (N_2908,N_1663,N_1670);
xor U2909 (N_2909,N_1575,N_1439);
xnor U2910 (N_2910,N_1881,N_1467);
xor U2911 (N_2911,N_1653,N_1989);
or U2912 (N_2912,N_1263,N_1287);
and U2913 (N_2913,N_1548,N_1177);
nand U2914 (N_2914,N_1036,N_1305);
nor U2915 (N_2915,N_1684,N_1723);
or U2916 (N_2916,N_1211,N_1826);
and U2917 (N_2917,N_1360,N_1615);
or U2918 (N_2918,N_1317,N_1640);
nand U2919 (N_2919,N_1563,N_1236);
nor U2920 (N_2920,N_1729,N_1501);
and U2921 (N_2921,N_1582,N_1146);
and U2922 (N_2922,N_1086,N_1232);
nor U2923 (N_2923,N_1839,N_1881);
and U2924 (N_2924,N_1355,N_1211);
nand U2925 (N_2925,N_1889,N_1300);
or U2926 (N_2926,N_1428,N_1720);
nor U2927 (N_2927,N_1847,N_1280);
xor U2928 (N_2928,N_1060,N_1788);
xor U2929 (N_2929,N_1277,N_1325);
or U2930 (N_2930,N_1255,N_1089);
or U2931 (N_2931,N_1379,N_1160);
and U2932 (N_2932,N_1904,N_1263);
nand U2933 (N_2933,N_1403,N_1061);
and U2934 (N_2934,N_1639,N_1629);
xor U2935 (N_2935,N_1463,N_1803);
nand U2936 (N_2936,N_1158,N_1974);
nor U2937 (N_2937,N_1856,N_1919);
and U2938 (N_2938,N_1839,N_1630);
nand U2939 (N_2939,N_1824,N_1708);
xnor U2940 (N_2940,N_1363,N_1173);
xor U2941 (N_2941,N_1735,N_1573);
or U2942 (N_2942,N_1143,N_1911);
and U2943 (N_2943,N_1274,N_1645);
nand U2944 (N_2944,N_1849,N_1898);
nor U2945 (N_2945,N_1028,N_1369);
nand U2946 (N_2946,N_1351,N_1848);
and U2947 (N_2947,N_1231,N_1831);
nor U2948 (N_2948,N_1645,N_1335);
nor U2949 (N_2949,N_1622,N_1830);
and U2950 (N_2950,N_1885,N_1601);
xor U2951 (N_2951,N_1348,N_1490);
or U2952 (N_2952,N_1451,N_1106);
nand U2953 (N_2953,N_1824,N_1538);
or U2954 (N_2954,N_1575,N_1520);
and U2955 (N_2955,N_1426,N_1859);
xnor U2956 (N_2956,N_1460,N_1946);
nor U2957 (N_2957,N_1641,N_1323);
and U2958 (N_2958,N_1897,N_1517);
and U2959 (N_2959,N_1627,N_1897);
and U2960 (N_2960,N_1585,N_1393);
and U2961 (N_2961,N_1870,N_1600);
or U2962 (N_2962,N_1515,N_1990);
and U2963 (N_2963,N_1090,N_1657);
xor U2964 (N_2964,N_1497,N_1710);
or U2965 (N_2965,N_1056,N_1260);
xnor U2966 (N_2966,N_1661,N_1964);
xor U2967 (N_2967,N_1506,N_1791);
nor U2968 (N_2968,N_1718,N_1160);
and U2969 (N_2969,N_1342,N_1684);
xor U2970 (N_2970,N_1480,N_1978);
or U2971 (N_2971,N_1729,N_1388);
nand U2972 (N_2972,N_1062,N_1150);
nand U2973 (N_2973,N_1977,N_1536);
xor U2974 (N_2974,N_1616,N_1157);
nand U2975 (N_2975,N_1133,N_1816);
and U2976 (N_2976,N_1480,N_1187);
xor U2977 (N_2977,N_1342,N_1871);
nor U2978 (N_2978,N_1535,N_1781);
or U2979 (N_2979,N_1121,N_1059);
and U2980 (N_2980,N_1269,N_1641);
and U2981 (N_2981,N_1829,N_1239);
or U2982 (N_2982,N_1527,N_1178);
and U2983 (N_2983,N_1758,N_1077);
nor U2984 (N_2984,N_1522,N_1118);
nand U2985 (N_2985,N_1108,N_1903);
xnor U2986 (N_2986,N_1960,N_1766);
and U2987 (N_2987,N_1024,N_1847);
and U2988 (N_2988,N_1546,N_1730);
or U2989 (N_2989,N_1728,N_1439);
nor U2990 (N_2990,N_1558,N_1720);
or U2991 (N_2991,N_1706,N_1465);
or U2992 (N_2992,N_1226,N_1820);
or U2993 (N_2993,N_1480,N_1203);
and U2994 (N_2994,N_1578,N_1364);
xnor U2995 (N_2995,N_1822,N_1245);
nand U2996 (N_2996,N_1277,N_1047);
or U2997 (N_2997,N_1699,N_1175);
or U2998 (N_2998,N_1408,N_1856);
xnor U2999 (N_2999,N_1701,N_1898);
xnor U3000 (N_3000,N_2487,N_2965);
nand U3001 (N_3001,N_2462,N_2898);
and U3002 (N_3002,N_2019,N_2452);
and U3003 (N_3003,N_2698,N_2821);
nor U3004 (N_3004,N_2252,N_2928);
nand U3005 (N_3005,N_2245,N_2447);
xnor U3006 (N_3006,N_2064,N_2617);
nor U3007 (N_3007,N_2827,N_2998);
xnor U3008 (N_3008,N_2396,N_2646);
nor U3009 (N_3009,N_2306,N_2107);
or U3010 (N_3010,N_2254,N_2630);
xor U3011 (N_3011,N_2048,N_2959);
and U3012 (N_3012,N_2446,N_2061);
and U3013 (N_3013,N_2903,N_2268);
nand U3014 (N_3014,N_2927,N_2093);
nor U3015 (N_3015,N_2278,N_2382);
nand U3016 (N_3016,N_2942,N_2349);
nor U3017 (N_3017,N_2970,N_2614);
nand U3018 (N_3018,N_2392,N_2830);
or U3019 (N_3019,N_2526,N_2621);
nand U3020 (N_3020,N_2146,N_2096);
and U3021 (N_3021,N_2424,N_2340);
nor U3022 (N_3022,N_2595,N_2983);
or U3023 (N_3023,N_2894,N_2869);
xnor U3024 (N_3024,N_2173,N_2732);
or U3025 (N_3025,N_2347,N_2601);
xor U3026 (N_3026,N_2355,N_2774);
nand U3027 (N_3027,N_2914,N_2425);
xnor U3028 (N_3028,N_2228,N_2012);
nor U3029 (N_3029,N_2844,N_2443);
nand U3030 (N_3030,N_2422,N_2657);
nand U3031 (N_3031,N_2257,N_2559);
or U3032 (N_3032,N_2592,N_2563);
nor U3033 (N_3033,N_2302,N_2641);
and U3034 (N_3034,N_2517,N_2231);
nand U3035 (N_3035,N_2969,N_2880);
nor U3036 (N_3036,N_2263,N_2238);
xor U3037 (N_3037,N_2185,N_2739);
nand U3038 (N_3038,N_2217,N_2095);
and U3039 (N_3039,N_2461,N_2674);
nor U3040 (N_3040,N_2301,N_2471);
nor U3041 (N_3041,N_2673,N_2459);
nor U3042 (N_3042,N_2489,N_2594);
nand U3043 (N_3043,N_2444,N_2530);
or U3044 (N_3044,N_2862,N_2362);
nor U3045 (N_3045,N_2016,N_2442);
nand U3046 (N_3046,N_2693,N_2399);
nor U3047 (N_3047,N_2464,N_2256);
nand U3048 (N_3048,N_2220,N_2551);
or U3049 (N_3049,N_2529,N_2935);
or U3050 (N_3050,N_2280,N_2125);
and U3051 (N_3051,N_2651,N_2549);
or U3052 (N_3052,N_2977,N_2162);
xnor U3053 (N_3053,N_2250,N_2802);
xnor U3054 (N_3054,N_2097,N_2138);
nand U3055 (N_3055,N_2864,N_2719);
nor U3056 (N_3056,N_2578,N_2961);
or U3057 (N_3057,N_2397,N_2099);
or U3058 (N_3058,N_2648,N_2121);
and U3059 (N_3059,N_2438,N_2090);
and U3060 (N_3060,N_2724,N_2418);
nand U3061 (N_3061,N_2351,N_2044);
nand U3062 (N_3062,N_2571,N_2834);
nand U3063 (N_3063,N_2117,N_2502);
or U3064 (N_3064,N_2825,N_2335);
nor U3065 (N_3065,N_2457,N_2807);
nor U3066 (N_3066,N_2264,N_2475);
nand U3067 (N_3067,N_2429,N_2276);
xnor U3068 (N_3068,N_2144,N_2359);
nor U3069 (N_3069,N_2607,N_2040);
xnor U3070 (N_3070,N_2790,N_2971);
nor U3071 (N_3071,N_2770,N_2671);
xnor U3072 (N_3072,N_2714,N_2199);
xor U3073 (N_3073,N_2750,N_2449);
xnor U3074 (N_3074,N_2161,N_2658);
nor U3075 (N_3075,N_2356,N_2796);
nor U3076 (N_3076,N_2391,N_2158);
nor U3077 (N_3077,N_2386,N_2157);
nand U3078 (N_3078,N_2988,N_2182);
nor U3079 (N_3079,N_2792,N_2833);
nor U3080 (N_3080,N_2331,N_2100);
and U3081 (N_3081,N_2017,N_2111);
nor U3082 (N_3082,N_2288,N_2177);
and U3083 (N_3083,N_2987,N_2664);
xor U3084 (N_3084,N_2877,N_2950);
xnor U3085 (N_3085,N_2700,N_2136);
nand U3086 (N_3086,N_2723,N_2067);
xor U3087 (N_3087,N_2179,N_2769);
nand U3088 (N_3088,N_2932,N_2900);
nand U3089 (N_3089,N_2532,N_2326);
nand U3090 (N_3090,N_2685,N_2148);
and U3091 (N_3091,N_2180,N_2902);
xnor U3092 (N_3092,N_2477,N_2929);
nand U3093 (N_3093,N_2063,N_2883);
nand U3094 (N_3094,N_2272,N_2696);
nor U3095 (N_3095,N_2773,N_2011);
and U3096 (N_3096,N_2856,N_2266);
or U3097 (N_3097,N_2817,N_2695);
nand U3098 (N_3098,N_2938,N_2101);
or U3099 (N_3099,N_2577,N_2677);
nor U3100 (N_3100,N_2564,N_2828);
and U3101 (N_3101,N_2163,N_2992);
and U3102 (N_3102,N_2388,N_2749);
or U3103 (N_3103,N_2921,N_2203);
nand U3104 (N_3104,N_2520,N_2643);
and U3105 (N_3105,N_2247,N_2077);
nor U3106 (N_3106,N_2324,N_2704);
or U3107 (N_3107,N_2416,N_2383);
nor U3108 (N_3108,N_2450,N_2645);
and U3109 (N_3109,N_2210,N_2219);
xor U3110 (N_3110,N_2133,N_2752);
xnor U3111 (N_3111,N_2015,N_2200);
and U3112 (N_3112,N_2634,N_2178);
xor U3113 (N_3113,N_2958,N_2370);
nor U3114 (N_3114,N_2801,N_2406);
and U3115 (N_3115,N_2761,N_2066);
or U3116 (N_3116,N_2859,N_2400);
xor U3117 (N_3117,N_2493,N_2947);
nand U3118 (N_3118,N_2610,N_2080);
or U3119 (N_3119,N_2389,N_2135);
xnor U3120 (N_3120,N_2013,N_2069);
xor U3121 (N_3121,N_2627,N_2169);
or U3122 (N_3122,N_2765,N_2020);
or U3123 (N_3123,N_2312,N_2613);
xnor U3124 (N_3124,N_2296,N_2835);
or U3125 (N_3125,N_2249,N_2281);
nand U3126 (N_3126,N_2141,N_2183);
xor U3127 (N_3127,N_2165,N_2378);
xor U3128 (N_3128,N_2027,N_2137);
nand U3129 (N_3129,N_2419,N_2838);
and U3130 (N_3130,N_2103,N_2758);
and U3131 (N_3131,N_2891,N_2271);
nand U3132 (N_3132,N_2995,N_2994);
or U3133 (N_3133,N_2244,N_2084);
or U3134 (N_3134,N_2376,N_2516);
nand U3135 (N_3135,N_2236,N_2171);
and U3136 (N_3136,N_2031,N_2556);
nor U3137 (N_3137,N_2939,N_2046);
and U3138 (N_3138,N_2497,N_2919);
xnor U3139 (N_3139,N_2408,N_2650);
and U3140 (N_3140,N_2336,N_2628);
xnor U3141 (N_3141,N_2709,N_2604);
nand U3142 (N_3142,N_2726,N_2809);
nand U3143 (N_3143,N_2925,N_2846);
and U3144 (N_3144,N_2706,N_2277);
nand U3145 (N_3145,N_2991,N_2813);
nand U3146 (N_3146,N_2678,N_2832);
nand U3147 (N_3147,N_2579,N_2500);
and U3148 (N_3148,N_2889,N_2829);
xor U3149 (N_3149,N_2690,N_2780);
nand U3150 (N_3150,N_2956,N_2218);
nor U3151 (N_3151,N_2523,N_2365);
or U3152 (N_3152,N_2711,N_2273);
nor U3153 (N_3153,N_2666,N_2297);
xnor U3154 (N_3154,N_2837,N_2025);
nand U3155 (N_3155,N_2779,N_2703);
nand U3156 (N_3156,N_2812,N_2744);
nor U3157 (N_3157,N_2030,N_2075);
xor U3158 (N_3158,N_2062,N_2002);
or U3159 (N_3159,N_2304,N_2985);
xnor U3160 (N_3160,N_2901,N_2831);
or U3161 (N_3161,N_2207,N_2633);
nor U3162 (N_3162,N_2583,N_2699);
nand U3163 (N_3163,N_2608,N_2049);
nand U3164 (N_3164,N_2167,N_2401);
or U3165 (N_3165,N_2842,N_2728);
nand U3166 (N_3166,N_2174,N_2753);
xor U3167 (N_3167,N_2113,N_2495);
or U3168 (N_3168,N_2688,N_2420);
nand U3169 (N_3169,N_2404,N_2629);
or U3170 (N_3170,N_2552,N_2763);
nand U3171 (N_3171,N_2885,N_2211);
nand U3172 (N_3172,N_2963,N_2521);
nand U3173 (N_3173,N_2308,N_2073);
nor U3174 (N_3174,N_2996,N_2631);
xnor U3175 (N_3175,N_2968,N_2981);
or U3176 (N_3176,N_2887,N_2267);
or U3177 (N_3177,N_2525,N_2072);
or U3178 (N_3178,N_2313,N_2081);
nand U3179 (N_3179,N_2599,N_2348);
nor U3180 (N_3180,N_2531,N_2733);
or U3181 (N_3181,N_2213,N_2960);
nand U3182 (N_3182,N_2691,N_2702);
nor U3183 (N_3183,N_2060,N_2852);
or U3184 (N_3184,N_2976,N_2307);
nand U3185 (N_3185,N_2474,N_2716);
and U3186 (N_3186,N_2858,N_2059);
xor U3187 (N_3187,N_2541,N_2374);
nand U3188 (N_3188,N_2022,N_2708);
nor U3189 (N_3189,N_2056,N_2786);
or U3190 (N_3190,N_2237,N_2897);
and U3191 (N_3191,N_2955,N_2147);
xnor U3192 (N_3192,N_2032,N_2488);
and U3193 (N_3193,N_2352,N_2116);
nand U3194 (N_3194,N_2941,N_2934);
xnor U3195 (N_3195,N_2819,N_2198);
or U3196 (N_3196,N_2204,N_2377);
and U3197 (N_3197,N_2553,N_2655);
or U3198 (N_3198,N_2870,N_2888);
nor U3199 (N_3199,N_2661,N_2142);
xnor U3200 (N_3200,N_2893,N_2395);
and U3201 (N_3201,N_2468,N_2155);
nor U3202 (N_3202,N_2094,N_2262);
nor U3203 (N_3203,N_2944,N_2620);
nor U3204 (N_3204,N_2980,N_2482);
or U3205 (N_3205,N_2293,N_2381);
or U3206 (N_3206,N_2164,N_2041);
nand U3207 (N_3207,N_2029,N_2582);
and U3208 (N_3208,N_2943,N_2734);
nand U3209 (N_3209,N_2189,N_2122);
xor U3210 (N_3210,N_2130,N_2717);
or U3211 (N_3211,N_2289,N_2490);
xor U3212 (N_3212,N_2637,N_2496);
or U3213 (N_3213,N_2258,N_2239);
or U3214 (N_3214,N_2149,N_2907);
or U3215 (N_3215,N_2322,N_2320);
nand U3216 (N_3216,N_2172,N_2848);
nor U3217 (N_3217,N_2342,N_2546);
or U3218 (N_3218,N_2283,N_2920);
xor U3219 (N_3219,N_2713,N_2675);
or U3220 (N_3220,N_2115,N_2091);
nor U3221 (N_3221,N_2587,N_2682);
nand U3222 (N_3222,N_2550,N_2315);
xnor U3223 (N_3223,N_2491,N_2818);
xor U3224 (N_3224,N_2334,N_2636);
nor U3225 (N_3225,N_2930,N_2451);
or U3226 (N_3226,N_2318,N_2330);
or U3227 (N_3227,N_2760,N_2465);
xor U3228 (N_3228,N_2603,N_2727);
and U3229 (N_3229,N_2363,N_2777);
and U3230 (N_3230,N_2413,N_2260);
nand U3231 (N_3231,N_2248,N_2951);
nor U3232 (N_3232,N_2403,N_2052);
nand U3233 (N_3233,N_2311,N_2622);
nand U3234 (N_3234,N_2722,N_2479);
nor U3235 (N_3235,N_2701,N_2865);
nor U3236 (N_3236,N_2205,N_2104);
and U3237 (N_3237,N_2566,N_2145);
nand U3238 (N_3238,N_2667,N_2843);
xnor U3239 (N_3239,N_2319,N_2784);
nor U3240 (N_3240,N_2088,N_2439);
xor U3241 (N_3241,N_2229,N_2473);
nor U3242 (N_3242,N_2906,N_2624);
nor U3243 (N_3243,N_2740,N_2937);
nand U3244 (N_3244,N_2776,N_2087);
or U3245 (N_3245,N_2954,N_2948);
xnor U3246 (N_3246,N_2193,N_2332);
and U3247 (N_3247,N_2861,N_2092);
xnor U3248 (N_3248,N_2979,N_2875);
or U3249 (N_3249,N_2772,N_2949);
and U3250 (N_3250,N_2082,N_2261);
nor U3251 (N_3251,N_2153,N_2242);
or U3252 (N_3252,N_2741,N_2508);
xor U3253 (N_3253,N_2507,N_2751);
xnor U3254 (N_3254,N_2569,N_2151);
nor U3255 (N_3255,N_2840,N_2933);
xnor U3256 (N_3256,N_2476,N_2923);
and U3257 (N_3257,N_2639,N_2454);
xnor U3258 (N_3258,N_2323,N_2366);
nand U3259 (N_3259,N_2557,N_2611);
and U3260 (N_3260,N_2787,N_2814);
nor U3261 (N_3261,N_2554,N_2710);
xor U3262 (N_3262,N_2572,N_2884);
or U3263 (N_3263,N_2874,N_2816);
nand U3264 (N_3264,N_2808,N_2547);
and U3265 (N_3265,N_2574,N_2748);
or U3266 (N_3266,N_2453,N_2668);
and U3267 (N_3267,N_2918,N_2102);
or U3268 (N_3268,N_2371,N_2086);
and U3269 (N_3269,N_2768,N_2385);
nor U3270 (N_3270,N_2882,N_2119);
or U3271 (N_3271,N_2509,N_2154);
xor U3272 (N_3272,N_2168,N_2513);
nand U3273 (N_3273,N_2600,N_2209);
and U3274 (N_3274,N_2738,N_2568);
xor U3275 (N_3275,N_2851,N_2054);
nor U3276 (N_3276,N_2384,N_2434);
nand U3277 (N_3277,N_2070,N_2916);
nand U3278 (N_3278,N_2803,N_2999);
nand U3279 (N_3279,N_2871,N_2501);
xor U3280 (N_3280,N_2591,N_2841);
or U3281 (N_3281,N_2896,N_2008);
or U3282 (N_3282,N_2310,N_2417);
nor U3283 (N_3283,N_2437,N_2612);
and U3284 (N_3284,N_2783,N_2043);
and U3285 (N_3285,N_2192,N_2292);
and U3286 (N_3286,N_2705,N_2047);
xor U3287 (N_3287,N_2576,N_2618);
or U3288 (N_3288,N_2033,N_2373);
xor U3289 (N_3289,N_2057,N_2390);
and U3290 (N_3290,N_2079,N_2867);
or U3291 (N_3291,N_2876,N_2873);
nor U3292 (N_3292,N_2333,N_2616);
and U3293 (N_3293,N_2632,N_2051);
nor U3294 (N_3294,N_2317,N_2227);
and U3295 (N_3295,N_2215,N_2364);
or U3296 (N_3296,N_2681,N_2234);
nand U3297 (N_3297,N_2156,N_2793);
and U3298 (N_3298,N_2899,N_2683);
or U3299 (N_3299,N_2360,N_2190);
nor U3300 (N_3300,N_2160,N_2527);
or U3301 (N_3301,N_2644,N_2432);
and U3302 (N_3302,N_2367,N_2623);
nand U3303 (N_3303,N_2849,N_2514);
and U3304 (N_3304,N_2068,N_2638);
nand U3305 (N_3305,N_2275,N_2625);
and U3306 (N_3306,N_2868,N_2026);
nor U3307 (N_3307,N_2565,N_2201);
or U3308 (N_3308,N_2372,N_2253);
or U3309 (N_3309,N_2109,N_2820);
nand U3310 (N_3310,N_2021,N_2036);
nand U3311 (N_3311,N_2660,N_2469);
and U3312 (N_3312,N_2926,N_2427);
xnor U3313 (N_3313,N_2872,N_2143);
xor U3314 (N_3314,N_2309,N_2795);
nor U3315 (N_3315,N_2619,N_2435);
nor U3316 (N_3316,N_2375,N_2120);
and U3317 (N_3317,N_2615,N_2050);
nand U3318 (N_3318,N_2196,N_2756);
xor U3319 (N_3319,N_2353,N_2184);
or U3320 (N_3320,N_2410,N_2522);
nor U3321 (N_3321,N_2314,N_2393);
or U3322 (N_3322,N_2775,N_2078);
nand U3323 (N_3323,N_2720,N_2878);
or U3324 (N_3324,N_2892,N_2537);
nand U3325 (N_3325,N_2361,N_2484);
and U3326 (N_3326,N_2506,N_2098);
and U3327 (N_3327,N_2555,N_2847);
nor U3328 (N_3328,N_2656,N_2166);
or U3329 (N_3329,N_2762,N_2483);
or U3330 (N_3330,N_2575,N_2039);
and U3331 (N_3331,N_2782,N_2560);
nand U3332 (N_3332,N_2584,N_2186);
and U3333 (N_3333,N_2232,N_2216);
nand U3334 (N_3334,N_2561,N_2511);
nand U3335 (N_3335,N_2692,N_2823);
and U3336 (N_3336,N_2542,N_2910);
or U3337 (N_3337,N_2518,N_2684);
nor U3338 (N_3338,N_2222,N_2535);
or U3339 (N_3339,N_2754,N_2853);
or U3340 (N_3340,N_2368,N_2387);
or U3341 (N_3341,N_2291,N_2037);
xnor U3342 (N_3342,N_2570,N_2197);
and U3343 (N_3343,N_2966,N_2676);
nor U3344 (N_3344,N_2824,N_2414);
and U3345 (N_3345,N_2225,N_2339);
nor U3346 (N_3346,N_2472,N_2598);
and U3347 (N_3347,N_2771,N_2904);
nand U3348 (N_3348,N_2735,N_2799);
xor U3349 (N_3349,N_2815,N_2499);
nand U3350 (N_3350,N_2839,N_2195);
nand U3351 (N_3351,N_2441,N_2863);
nor U3352 (N_3352,N_2781,N_2159);
and U3353 (N_3353,N_2321,N_2759);
or U3354 (N_3354,N_2010,N_2652);
or U3355 (N_3355,N_2132,N_2058);
nand U3356 (N_3356,N_2004,N_2085);
nor U3357 (N_3357,N_2456,N_2394);
or U3358 (N_3358,N_2640,N_2035);
or U3359 (N_3359,N_2328,N_2785);
or U3360 (N_3360,N_2743,N_2076);
or U3361 (N_3361,N_2845,N_2797);
and U3362 (N_3362,N_2074,N_2953);
nor U3363 (N_3363,N_2492,N_2533);
nand U3364 (N_3364,N_2654,N_2409);
xnor U3365 (N_3365,N_2718,N_2007);
or U3366 (N_3366,N_2562,N_2590);
nand U3367 (N_3367,N_2505,N_2028);
and U3368 (N_3368,N_2265,N_2504);
xnor U3369 (N_3369,N_2285,N_2984);
nor U3370 (N_3370,N_2665,N_2972);
xor U3371 (N_3371,N_2905,N_2712);
and U3372 (N_3372,N_2379,N_2338);
nand U3373 (N_3373,N_2226,N_2246);
xor U3374 (N_3374,N_2567,N_2746);
nand U3375 (N_3375,N_2548,N_2014);
or U3376 (N_3376,N_2045,N_2663);
xnor U3377 (N_3377,N_2042,N_2512);
nand U3378 (N_3378,N_2118,N_2881);
nor U3379 (N_3379,N_2912,N_2680);
nand U3380 (N_3380,N_2642,N_2936);
nor U3381 (N_3381,N_2486,N_2662);
or U3382 (N_3382,N_2240,N_2343);
and U3383 (N_3383,N_2745,N_2053);
nand U3384 (N_3384,N_2689,N_2672);
nor U3385 (N_3385,N_2973,N_2911);
and U3386 (N_3386,N_2747,N_2931);
or U3387 (N_3387,N_2398,N_2152);
nand U3388 (N_3388,N_2202,N_2055);
nand U3389 (N_3389,N_2433,N_2445);
nand U3390 (N_3390,N_2649,N_2114);
or U3391 (N_3391,N_2485,N_2975);
nor U3392 (N_3392,N_2860,N_2494);
nor U3393 (N_3393,N_2299,N_2669);
nand U3394 (N_3394,N_2997,N_2290);
and U3395 (N_3395,N_2009,N_2071);
or U3396 (N_3396,N_2804,N_2778);
or U3397 (N_3397,N_2105,N_2791);
and U3398 (N_3398,N_2503,N_2806);
nand U3399 (N_3399,N_2725,N_2127);
or U3400 (N_3400,N_2659,N_2805);
or U3401 (N_3401,N_2543,N_2380);
and U3402 (N_3402,N_2593,N_2284);
and U3403 (N_3403,N_2034,N_2194);
nor U3404 (N_3404,N_2811,N_2766);
nor U3405 (N_3405,N_2697,N_2346);
xor U3406 (N_3406,N_2337,N_2524);
xor U3407 (N_3407,N_2989,N_2005);
xnor U3408 (N_3408,N_2810,N_2269);
nand U3409 (N_3409,N_2890,N_2915);
or U3410 (N_3410,N_2407,N_2440);
nand U3411 (N_3411,N_2128,N_2606);
or U3412 (N_3412,N_2428,N_2255);
or U3413 (N_3413,N_2964,N_2126);
or U3414 (N_3414,N_2478,N_2235);
nor U3415 (N_3415,N_2913,N_2498);
or U3416 (N_3416,N_2350,N_2946);
or U3417 (N_3417,N_2251,N_2731);
xor U3418 (N_3418,N_2515,N_2139);
nor U3419 (N_3419,N_2836,N_2679);
or U3420 (N_3420,N_2986,N_2962);
nand U3421 (N_3421,N_2279,N_2586);
and U3422 (N_3422,N_2917,N_2305);
nand U3423 (N_3423,N_2895,N_2123);
xnor U3424 (N_3424,N_2589,N_2794);
nor U3425 (N_3425,N_2857,N_2581);
and U3426 (N_3426,N_2083,N_2585);
or U3427 (N_3427,N_2952,N_2241);
nor U3428 (N_3428,N_2140,N_2191);
and U3429 (N_3429,N_2850,N_2647);
and U3430 (N_3430,N_2089,N_2412);
or U3431 (N_3431,N_2957,N_2580);
xor U3432 (N_3432,N_2737,N_2736);
nor U3433 (N_3433,N_2539,N_2065);
xnor U3434 (N_3434,N_2221,N_2327);
xnor U3435 (N_3435,N_2430,N_2423);
nor U3436 (N_3436,N_2609,N_2908);
nor U3437 (N_3437,N_2448,N_2481);
or U3438 (N_3438,N_2480,N_2329);
nand U3439 (N_3439,N_2879,N_2798);
nand U3440 (N_3440,N_2206,N_2295);
nor U3441 (N_3441,N_2274,N_2181);
and U3442 (N_3442,N_2993,N_2715);
nand U3443 (N_3443,N_2538,N_2558);
and U3444 (N_3444,N_2764,N_2303);
nor U3445 (N_3445,N_2001,N_2259);
and U3446 (N_3446,N_2131,N_2730);
or U3447 (N_3447,N_2024,N_2967);
xor U3448 (N_3448,N_2826,N_2940);
nor U3449 (N_3449,N_2038,N_2978);
nand U3450 (N_3450,N_2855,N_2170);
nor U3451 (N_3451,N_2415,N_2573);
nor U3452 (N_3452,N_2341,N_2411);
or U3453 (N_3453,N_2458,N_2605);
nor U3454 (N_3454,N_2286,N_2534);
nand U3455 (N_3455,N_2544,N_2421);
nand U3456 (N_3456,N_2528,N_2540);
nor U3457 (N_3457,N_2018,N_2006);
nand U3458 (N_3458,N_2208,N_2886);
nor U3459 (N_3459,N_2510,N_2223);
nand U3460 (N_3460,N_2922,N_2129);
and U3461 (N_3461,N_2023,N_2990);
nand U3462 (N_3462,N_2402,N_2405);
or U3463 (N_3463,N_2270,N_2982);
xnor U3464 (N_3464,N_2767,N_2742);
or U3465 (N_3465,N_2316,N_2467);
nor U3466 (N_3466,N_2626,N_2150);
nand U3467 (N_3467,N_2670,N_2003);
and U3468 (N_3468,N_2354,N_2188);
nor U3469 (N_3469,N_2909,N_2325);
and U3470 (N_3470,N_2463,N_2588);
nand U3471 (N_3471,N_2460,N_2597);
and U3472 (N_3472,N_2545,N_2431);
and U3473 (N_3473,N_2187,N_2224);
nand U3474 (N_3474,N_2000,N_2854);
nor U3475 (N_3475,N_2687,N_2602);
nor U3476 (N_3476,N_2466,N_2243);
and U3477 (N_3477,N_2344,N_2233);
or U3478 (N_3478,N_2369,N_2470);
nor U3479 (N_3479,N_2124,N_2357);
or U3480 (N_3480,N_2686,N_2214);
or U3481 (N_3481,N_2924,N_2108);
and U3482 (N_3482,N_2282,N_2974);
nand U3483 (N_3483,N_2212,N_2294);
nor U3484 (N_3484,N_2707,N_2945);
nor U3485 (N_3485,N_2436,N_2300);
and U3486 (N_3486,N_2298,N_2287);
nor U3487 (N_3487,N_2800,N_2345);
xnor U3488 (N_3488,N_2757,N_2176);
or U3489 (N_3489,N_2721,N_2175);
or U3490 (N_3490,N_2426,N_2755);
and U3491 (N_3491,N_2596,N_2358);
nor U3492 (N_3492,N_2822,N_2519);
or U3493 (N_3493,N_2866,N_2106);
and U3494 (N_3494,N_2455,N_2110);
nand U3495 (N_3495,N_2230,N_2536);
nor U3496 (N_3496,N_2729,N_2694);
xor U3497 (N_3497,N_2134,N_2788);
xor U3498 (N_3498,N_2635,N_2653);
xor U3499 (N_3499,N_2789,N_2112);
xor U3500 (N_3500,N_2435,N_2054);
xor U3501 (N_3501,N_2494,N_2283);
and U3502 (N_3502,N_2831,N_2292);
and U3503 (N_3503,N_2811,N_2218);
nand U3504 (N_3504,N_2498,N_2920);
nand U3505 (N_3505,N_2911,N_2439);
or U3506 (N_3506,N_2663,N_2310);
xnor U3507 (N_3507,N_2333,N_2859);
and U3508 (N_3508,N_2523,N_2736);
and U3509 (N_3509,N_2373,N_2035);
and U3510 (N_3510,N_2698,N_2680);
nand U3511 (N_3511,N_2491,N_2852);
or U3512 (N_3512,N_2257,N_2408);
nor U3513 (N_3513,N_2914,N_2399);
or U3514 (N_3514,N_2527,N_2045);
nor U3515 (N_3515,N_2878,N_2806);
nand U3516 (N_3516,N_2440,N_2877);
xor U3517 (N_3517,N_2780,N_2160);
nor U3518 (N_3518,N_2054,N_2522);
and U3519 (N_3519,N_2641,N_2831);
and U3520 (N_3520,N_2648,N_2169);
or U3521 (N_3521,N_2942,N_2935);
nand U3522 (N_3522,N_2240,N_2994);
nor U3523 (N_3523,N_2377,N_2371);
or U3524 (N_3524,N_2043,N_2309);
or U3525 (N_3525,N_2258,N_2796);
nand U3526 (N_3526,N_2808,N_2334);
or U3527 (N_3527,N_2583,N_2069);
or U3528 (N_3528,N_2978,N_2925);
nand U3529 (N_3529,N_2825,N_2584);
or U3530 (N_3530,N_2059,N_2545);
xnor U3531 (N_3531,N_2994,N_2226);
and U3532 (N_3532,N_2009,N_2214);
nand U3533 (N_3533,N_2652,N_2977);
xnor U3534 (N_3534,N_2201,N_2032);
or U3535 (N_3535,N_2055,N_2699);
or U3536 (N_3536,N_2584,N_2291);
and U3537 (N_3537,N_2351,N_2497);
nand U3538 (N_3538,N_2568,N_2601);
and U3539 (N_3539,N_2382,N_2378);
and U3540 (N_3540,N_2727,N_2645);
xnor U3541 (N_3541,N_2684,N_2321);
xor U3542 (N_3542,N_2655,N_2283);
nor U3543 (N_3543,N_2578,N_2248);
xnor U3544 (N_3544,N_2955,N_2159);
and U3545 (N_3545,N_2637,N_2822);
xor U3546 (N_3546,N_2584,N_2219);
nor U3547 (N_3547,N_2658,N_2546);
and U3548 (N_3548,N_2696,N_2752);
nor U3549 (N_3549,N_2370,N_2598);
or U3550 (N_3550,N_2839,N_2772);
xor U3551 (N_3551,N_2244,N_2208);
or U3552 (N_3552,N_2166,N_2140);
or U3553 (N_3553,N_2066,N_2558);
and U3554 (N_3554,N_2132,N_2888);
xnor U3555 (N_3555,N_2228,N_2523);
nor U3556 (N_3556,N_2935,N_2908);
and U3557 (N_3557,N_2234,N_2701);
and U3558 (N_3558,N_2998,N_2727);
xnor U3559 (N_3559,N_2409,N_2296);
and U3560 (N_3560,N_2847,N_2984);
nand U3561 (N_3561,N_2263,N_2339);
xnor U3562 (N_3562,N_2444,N_2004);
nor U3563 (N_3563,N_2362,N_2682);
nand U3564 (N_3564,N_2847,N_2435);
or U3565 (N_3565,N_2522,N_2655);
and U3566 (N_3566,N_2633,N_2116);
and U3567 (N_3567,N_2133,N_2868);
or U3568 (N_3568,N_2632,N_2970);
nor U3569 (N_3569,N_2867,N_2735);
nand U3570 (N_3570,N_2225,N_2826);
nor U3571 (N_3571,N_2523,N_2522);
or U3572 (N_3572,N_2659,N_2347);
nor U3573 (N_3573,N_2753,N_2199);
nand U3574 (N_3574,N_2111,N_2900);
xnor U3575 (N_3575,N_2785,N_2511);
nor U3576 (N_3576,N_2612,N_2002);
and U3577 (N_3577,N_2228,N_2213);
and U3578 (N_3578,N_2719,N_2927);
xor U3579 (N_3579,N_2187,N_2839);
and U3580 (N_3580,N_2883,N_2317);
xnor U3581 (N_3581,N_2625,N_2410);
xor U3582 (N_3582,N_2250,N_2912);
xor U3583 (N_3583,N_2613,N_2690);
and U3584 (N_3584,N_2819,N_2140);
or U3585 (N_3585,N_2820,N_2498);
nand U3586 (N_3586,N_2233,N_2200);
nand U3587 (N_3587,N_2960,N_2482);
nor U3588 (N_3588,N_2285,N_2140);
xor U3589 (N_3589,N_2304,N_2252);
and U3590 (N_3590,N_2807,N_2531);
nor U3591 (N_3591,N_2583,N_2657);
xnor U3592 (N_3592,N_2479,N_2468);
or U3593 (N_3593,N_2151,N_2865);
nor U3594 (N_3594,N_2551,N_2341);
nor U3595 (N_3595,N_2089,N_2846);
xnor U3596 (N_3596,N_2297,N_2745);
nand U3597 (N_3597,N_2257,N_2060);
xor U3598 (N_3598,N_2610,N_2484);
and U3599 (N_3599,N_2819,N_2264);
xnor U3600 (N_3600,N_2781,N_2851);
nor U3601 (N_3601,N_2281,N_2770);
xnor U3602 (N_3602,N_2741,N_2607);
nor U3603 (N_3603,N_2210,N_2619);
nand U3604 (N_3604,N_2632,N_2713);
or U3605 (N_3605,N_2208,N_2564);
and U3606 (N_3606,N_2489,N_2988);
or U3607 (N_3607,N_2710,N_2967);
or U3608 (N_3608,N_2723,N_2121);
xnor U3609 (N_3609,N_2662,N_2982);
and U3610 (N_3610,N_2304,N_2697);
or U3611 (N_3611,N_2000,N_2085);
xnor U3612 (N_3612,N_2315,N_2841);
and U3613 (N_3613,N_2875,N_2232);
or U3614 (N_3614,N_2318,N_2296);
xnor U3615 (N_3615,N_2515,N_2300);
and U3616 (N_3616,N_2988,N_2491);
xor U3617 (N_3617,N_2008,N_2330);
and U3618 (N_3618,N_2739,N_2689);
nor U3619 (N_3619,N_2079,N_2683);
and U3620 (N_3620,N_2040,N_2856);
or U3621 (N_3621,N_2840,N_2144);
and U3622 (N_3622,N_2252,N_2048);
xor U3623 (N_3623,N_2249,N_2547);
nor U3624 (N_3624,N_2607,N_2363);
and U3625 (N_3625,N_2705,N_2839);
or U3626 (N_3626,N_2571,N_2177);
nand U3627 (N_3627,N_2764,N_2827);
or U3628 (N_3628,N_2943,N_2030);
or U3629 (N_3629,N_2644,N_2359);
nor U3630 (N_3630,N_2280,N_2138);
xor U3631 (N_3631,N_2567,N_2356);
xor U3632 (N_3632,N_2090,N_2121);
xnor U3633 (N_3633,N_2465,N_2559);
xor U3634 (N_3634,N_2729,N_2833);
or U3635 (N_3635,N_2573,N_2919);
xnor U3636 (N_3636,N_2518,N_2280);
xnor U3637 (N_3637,N_2477,N_2664);
nor U3638 (N_3638,N_2291,N_2466);
or U3639 (N_3639,N_2377,N_2537);
and U3640 (N_3640,N_2155,N_2713);
and U3641 (N_3641,N_2936,N_2201);
and U3642 (N_3642,N_2975,N_2946);
nor U3643 (N_3643,N_2619,N_2516);
nand U3644 (N_3644,N_2334,N_2399);
or U3645 (N_3645,N_2271,N_2538);
and U3646 (N_3646,N_2932,N_2690);
nor U3647 (N_3647,N_2946,N_2887);
and U3648 (N_3648,N_2330,N_2776);
nor U3649 (N_3649,N_2125,N_2131);
nand U3650 (N_3650,N_2551,N_2681);
xnor U3651 (N_3651,N_2128,N_2704);
xor U3652 (N_3652,N_2008,N_2309);
xor U3653 (N_3653,N_2671,N_2819);
nor U3654 (N_3654,N_2530,N_2416);
and U3655 (N_3655,N_2886,N_2688);
xor U3656 (N_3656,N_2918,N_2161);
nor U3657 (N_3657,N_2225,N_2972);
and U3658 (N_3658,N_2177,N_2703);
or U3659 (N_3659,N_2922,N_2716);
nor U3660 (N_3660,N_2933,N_2771);
and U3661 (N_3661,N_2779,N_2731);
or U3662 (N_3662,N_2702,N_2430);
xnor U3663 (N_3663,N_2808,N_2253);
xnor U3664 (N_3664,N_2531,N_2553);
or U3665 (N_3665,N_2054,N_2389);
xor U3666 (N_3666,N_2433,N_2281);
nand U3667 (N_3667,N_2523,N_2548);
xor U3668 (N_3668,N_2574,N_2290);
or U3669 (N_3669,N_2965,N_2892);
nor U3670 (N_3670,N_2510,N_2069);
nand U3671 (N_3671,N_2540,N_2713);
or U3672 (N_3672,N_2539,N_2087);
nor U3673 (N_3673,N_2551,N_2644);
nand U3674 (N_3674,N_2000,N_2579);
or U3675 (N_3675,N_2723,N_2117);
nand U3676 (N_3676,N_2795,N_2064);
and U3677 (N_3677,N_2084,N_2999);
nor U3678 (N_3678,N_2921,N_2244);
xor U3679 (N_3679,N_2489,N_2131);
and U3680 (N_3680,N_2688,N_2868);
nand U3681 (N_3681,N_2391,N_2005);
and U3682 (N_3682,N_2948,N_2791);
and U3683 (N_3683,N_2136,N_2805);
or U3684 (N_3684,N_2088,N_2736);
or U3685 (N_3685,N_2152,N_2035);
nand U3686 (N_3686,N_2868,N_2792);
or U3687 (N_3687,N_2937,N_2840);
nor U3688 (N_3688,N_2752,N_2801);
and U3689 (N_3689,N_2252,N_2984);
and U3690 (N_3690,N_2430,N_2931);
nor U3691 (N_3691,N_2659,N_2729);
or U3692 (N_3692,N_2950,N_2659);
or U3693 (N_3693,N_2005,N_2067);
xnor U3694 (N_3694,N_2086,N_2611);
xor U3695 (N_3695,N_2958,N_2909);
xnor U3696 (N_3696,N_2823,N_2427);
or U3697 (N_3697,N_2861,N_2789);
and U3698 (N_3698,N_2214,N_2365);
nand U3699 (N_3699,N_2749,N_2635);
xor U3700 (N_3700,N_2754,N_2504);
nor U3701 (N_3701,N_2745,N_2460);
and U3702 (N_3702,N_2002,N_2362);
nand U3703 (N_3703,N_2199,N_2376);
xnor U3704 (N_3704,N_2630,N_2677);
nor U3705 (N_3705,N_2182,N_2799);
or U3706 (N_3706,N_2537,N_2686);
nor U3707 (N_3707,N_2259,N_2448);
or U3708 (N_3708,N_2999,N_2165);
nor U3709 (N_3709,N_2696,N_2948);
and U3710 (N_3710,N_2303,N_2105);
nand U3711 (N_3711,N_2966,N_2352);
and U3712 (N_3712,N_2324,N_2950);
and U3713 (N_3713,N_2621,N_2173);
or U3714 (N_3714,N_2174,N_2958);
nand U3715 (N_3715,N_2665,N_2108);
xor U3716 (N_3716,N_2822,N_2708);
nand U3717 (N_3717,N_2738,N_2849);
nand U3718 (N_3718,N_2506,N_2973);
nand U3719 (N_3719,N_2515,N_2319);
xnor U3720 (N_3720,N_2095,N_2657);
nand U3721 (N_3721,N_2866,N_2388);
and U3722 (N_3722,N_2779,N_2267);
xnor U3723 (N_3723,N_2535,N_2542);
xnor U3724 (N_3724,N_2368,N_2577);
and U3725 (N_3725,N_2250,N_2885);
or U3726 (N_3726,N_2628,N_2118);
nor U3727 (N_3727,N_2892,N_2010);
nand U3728 (N_3728,N_2425,N_2094);
nor U3729 (N_3729,N_2555,N_2805);
nand U3730 (N_3730,N_2961,N_2003);
or U3731 (N_3731,N_2291,N_2976);
nand U3732 (N_3732,N_2777,N_2201);
or U3733 (N_3733,N_2847,N_2866);
or U3734 (N_3734,N_2588,N_2145);
nand U3735 (N_3735,N_2992,N_2052);
nand U3736 (N_3736,N_2025,N_2581);
nand U3737 (N_3737,N_2295,N_2765);
and U3738 (N_3738,N_2803,N_2308);
and U3739 (N_3739,N_2589,N_2208);
xnor U3740 (N_3740,N_2715,N_2603);
nor U3741 (N_3741,N_2601,N_2308);
nand U3742 (N_3742,N_2209,N_2386);
nand U3743 (N_3743,N_2018,N_2180);
nand U3744 (N_3744,N_2051,N_2272);
nand U3745 (N_3745,N_2666,N_2300);
nand U3746 (N_3746,N_2654,N_2799);
and U3747 (N_3747,N_2125,N_2168);
or U3748 (N_3748,N_2809,N_2377);
xor U3749 (N_3749,N_2086,N_2214);
nand U3750 (N_3750,N_2849,N_2432);
nor U3751 (N_3751,N_2582,N_2976);
nor U3752 (N_3752,N_2735,N_2433);
nor U3753 (N_3753,N_2985,N_2747);
and U3754 (N_3754,N_2263,N_2362);
xor U3755 (N_3755,N_2498,N_2081);
xnor U3756 (N_3756,N_2890,N_2865);
or U3757 (N_3757,N_2961,N_2329);
xnor U3758 (N_3758,N_2806,N_2203);
nor U3759 (N_3759,N_2403,N_2570);
nand U3760 (N_3760,N_2451,N_2682);
nor U3761 (N_3761,N_2156,N_2766);
nor U3762 (N_3762,N_2373,N_2426);
xor U3763 (N_3763,N_2496,N_2386);
xnor U3764 (N_3764,N_2970,N_2862);
nor U3765 (N_3765,N_2880,N_2420);
nand U3766 (N_3766,N_2749,N_2931);
or U3767 (N_3767,N_2057,N_2293);
nand U3768 (N_3768,N_2413,N_2088);
or U3769 (N_3769,N_2857,N_2816);
nor U3770 (N_3770,N_2274,N_2382);
xnor U3771 (N_3771,N_2988,N_2860);
nor U3772 (N_3772,N_2978,N_2882);
and U3773 (N_3773,N_2165,N_2911);
or U3774 (N_3774,N_2399,N_2448);
or U3775 (N_3775,N_2984,N_2996);
nand U3776 (N_3776,N_2495,N_2323);
xnor U3777 (N_3777,N_2695,N_2784);
nand U3778 (N_3778,N_2911,N_2192);
xnor U3779 (N_3779,N_2468,N_2621);
or U3780 (N_3780,N_2712,N_2818);
and U3781 (N_3781,N_2411,N_2612);
nand U3782 (N_3782,N_2065,N_2106);
nor U3783 (N_3783,N_2543,N_2234);
or U3784 (N_3784,N_2468,N_2832);
or U3785 (N_3785,N_2154,N_2313);
xor U3786 (N_3786,N_2088,N_2597);
xor U3787 (N_3787,N_2911,N_2907);
nand U3788 (N_3788,N_2175,N_2642);
xor U3789 (N_3789,N_2502,N_2213);
nand U3790 (N_3790,N_2859,N_2040);
nand U3791 (N_3791,N_2150,N_2476);
or U3792 (N_3792,N_2983,N_2711);
nand U3793 (N_3793,N_2186,N_2538);
nor U3794 (N_3794,N_2612,N_2599);
nor U3795 (N_3795,N_2391,N_2275);
and U3796 (N_3796,N_2224,N_2733);
and U3797 (N_3797,N_2102,N_2529);
xnor U3798 (N_3798,N_2900,N_2236);
and U3799 (N_3799,N_2492,N_2785);
nor U3800 (N_3800,N_2606,N_2689);
nand U3801 (N_3801,N_2481,N_2716);
and U3802 (N_3802,N_2008,N_2144);
nor U3803 (N_3803,N_2698,N_2732);
or U3804 (N_3804,N_2410,N_2352);
or U3805 (N_3805,N_2041,N_2104);
nor U3806 (N_3806,N_2718,N_2732);
and U3807 (N_3807,N_2948,N_2237);
nor U3808 (N_3808,N_2682,N_2591);
or U3809 (N_3809,N_2283,N_2056);
nand U3810 (N_3810,N_2751,N_2245);
xor U3811 (N_3811,N_2719,N_2189);
and U3812 (N_3812,N_2940,N_2763);
nand U3813 (N_3813,N_2939,N_2943);
xor U3814 (N_3814,N_2275,N_2806);
xor U3815 (N_3815,N_2026,N_2172);
or U3816 (N_3816,N_2602,N_2648);
nor U3817 (N_3817,N_2620,N_2348);
or U3818 (N_3818,N_2774,N_2533);
nor U3819 (N_3819,N_2838,N_2881);
nor U3820 (N_3820,N_2510,N_2632);
or U3821 (N_3821,N_2260,N_2530);
nor U3822 (N_3822,N_2337,N_2527);
nor U3823 (N_3823,N_2507,N_2649);
or U3824 (N_3824,N_2022,N_2178);
xor U3825 (N_3825,N_2436,N_2786);
or U3826 (N_3826,N_2840,N_2783);
or U3827 (N_3827,N_2768,N_2693);
or U3828 (N_3828,N_2682,N_2293);
and U3829 (N_3829,N_2151,N_2470);
nand U3830 (N_3830,N_2952,N_2494);
xor U3831 (N_3831,N_2958,N_2100);
nand U3832 (N_3832,N_2174,N_2013);
nor U3833 (N_3833,N_2886,N_2188);
or U3834 (N_3834,N_2909,N_2123);
nand U3835 (N_3835,N_2828,N_2265);
nor U3836 (N_3836,N_2838,N_2114);
nor U3837 (N_3837,N_2486,N_2860);
and U3838 (N_3838,N_2948,N_2962);
or U3839 (N_3839,N_2412,N_2970);
nand U3840 (N_3840,N_2757,N_2977);
or U3841 (N_3841,N_2195,N_2407);
or U3842 (N_3842,N_2457,N_2407);
or U3843 (N_3843,N_2154,N_2990);
or U3844 (N_3844,N_2597,N_2520);
xor U3845 (N_3845,N_2410,N_2172);
xnor U3846 (N_3846,N_2589,N_2213);
and U3847 (N_3847,N_2658,N_2487);
or U3848 (N_3848,N_2561,N_2276);
nor U3849 (N_3849,N_2101,N_2171);
nor U3850 (N_3850,N_2085,N_2150);
and U3851 (N_3851,N_2959,N_2513);
nand U3852 (N_3852,N_2587,N_2261);
nand U3853 (N_3853,N_2197,N_2910);
or U3854 (N_3854,N_2899,N_2890);
and U3855 (N_3855,N_2245,N_2272);
xor U3856 (N_3856,N_2037,N_2242);
or U3857 (N_3857,N_2435,N_2423);
nor U3858 (N_3858,N_2430,N_2216);
and U3859 (N_3859,N_2222,N_2219);
and U3860 (N_3860,N_2705,N_2372);
nor U3861 (N_3861,N_2872,N_2479);
xnor U3862 (N_3862,N_2318,N_2212);
xor U3863 (N_3863,N_2433,N_2285);
nand U3864 (N_3864,N_2130,N_2289);
and U3865 (N_3865,N_2827,N_2396);
and U3866 (N_3866,N_2616,N_2708);
nor U3867 (N_3867,N_2378,N_2725);
and U3868 (N_3868,N_2979,N_2528);
nor U3869 (N_3869,N_2672,N_2452);
and U3870 (N_3870,N_2907,N_2112);
nor U3871 (N_3871,N_2793,N_2401);
and U3872 (N_3872,N_2466,N_2323);
xor U3873 (N_3873,N_2654,N_2226);
xnor U3874 (N_3874,N_2830,N_2619);
or U3875 (N_3875,N_2807,N_2857);
or U3876 (N_3876,N_2702,N_2719);
nor U3877 (N_3877,N_2054,N_2877);
xnor U3878 (N_3878,N_2085,N_2619);
nor U3879 (N_3879,N_2411,N_2298);
nor U3880 (N_3880,N_2354,N_2599);
or U3881 (N_3881,N_2816,N_2548);
nand U3882 (N_3882,N_2113,N_2594);
or U3883 (N_3883,N_2330,N_2549);
nor U3884 (N_3884,N_2194,N_2790);
xnor U3885 (N_3885,N_2734,N_2691);
nor U3886 (N_3886,N_2844,N_2220);
and U3887 (N_3887,N_2745,N_2476);
nor U3888 (N_3888,N_2730,N_2355);
nor U3889 (N_3889,N_2203,N_2780);
nor U3890 (N_3890,N_2177,N_2163);
or U3891 (N_3891,N_2632,N_2161);
or U3892 (N_3892,N_2182,N_2484);
and U3893 (N_3893,N_2606,N_2637);
nor U3894 (N_3894,N_2549,N_2544);
xor U3895 (N_3895,N_2326,N_2792);
and U3896 (N_3896,N_2506,N_2461);
and U3897 (N_3897,N_2201,N_2477);
nand U3898 (N_3898,N_2621,N_2559);
nor U3899 (N_3899,N_2482,N_2657);
or U3900 (N_3900,N_2716,N_2315);
or U3901 (N_3901,N_2026,N_2682);
and U3902 (N_3902,N_2929,N_2412);
nand U3903 (N_3903,N_2512,N_2579);
xnor U3904 (N_3904,N_2152,N_2198);
or U3905 (N_3905,N_2069,N_2245);
and U3906 (N_3906,N_2499,N_2424);
and U3907 (N_3907,N_2160,N_2815);
and U3908 (N_3908,N_2853,N_2147);
or U3909 (N_3909,N_2246,N_2739);
nand U3910 (N_3910,N_2467,N_2571);
nand U3911 (N_3911,N_2587,N_2558);
xnor U3912 (N_3912,N_2914,N_2876);
and U3913 (N_3913,N_2607,N_2605);
nor U3914 (N_3914,N_2113,N_2886);
nor U3915 (N_3915,N_2722,N_2407);
nor U3916 (N_3916,N_2003,N_2784);
nor U3917 (N_3917,N_2228,N_2667);
or U3918 (N_3918,N_2930,N_2519);
and U3919 (N_3919,N_2255,N_2228);
or U3920 (N_3920,N_2436,N_2753);
or U3921 (N_3921,N_2331,N_2134);
nand U3922 (N_3922,N_2830,N_2482);
nand U3923 (N_3923,N_2088,N_2404);
and U3924 (N_3924,N_2021,N_2524);
nor U3925 (N_3925,N_2314,N_2536);
xnor U3926 (N_3926,N_2463,N_2277);
or U3927 (N_3927,N_2399,N_2115);
xor U3928 (N_3928,N_2818,N_2009);
nand U3929 (N_3929,N_2613,N_2820);
xnor U3930 (N_3930,N_2317,N_2429);
nor U3931 (N_3931,N_2975,N_2338);
or U3932 (N_3932,N_2870,N_2124);
nand U3933 (N_3933,N_2189,N_2726);
nand U3934 (N_3934,N_2606,N_2767);
nand U3935 (N_3935,N_2037,N_2074);
xnor U3936 (N_3936,N_2413,N_2343);
and U3937 (N_3937,N_2194,N_2427);
nand U3938 (N_3938,N_2453,N_2141);
or U3939 (N_3939,N_2951,N_2191);
nor U3940 (N_3940,N_2840,N_2317);
or U3941 (N_3941,N_2919,N_2302);
nor U3942 (N_3942,N_2855,N_2779);
xor U3943 (N_3943,N_2953,N_2586);
nand U3944 (N_3944,N_2762,N_2747);
and U3945 (N_3945,N_2630,N_2685);
nand U3946 (N_3946,N_2824,N_2172);
and U3947 (N_3947,N_2141,N_2390);
or U3948 (N_3948,N_2681,N_2626);
xor U3949 (N_3949,N_2197,N_2686);
nand U3950 (N_3950,N_2304,N_2040);
nor U3951 (N_3951,N_2160,N_2272);
or U3952 (N_3952,N_2664,N_2117);
and U3953 (N_3953,N_2420,N_2496);
and U3954 (N_3954,N_2165,N_2624);
and U3955 (N_3955,N_2074,N_2446);
and U3956 (N_3956,N_2622,N_2660);
or U3957 (N_3957,N_2190,N_2200);
nand U3958 (N_3958,N_2196,N_2881);
xor U3959 (N_3959,N_2912,N_2810);
and U3960 (N_3960,N_2514,N_2727);
xor U3961 (N_3961,N_2559,N_2053);
and U3962 (N_3962,N_2588,N_2009);
or U3963 (N_3963,N_2040,N_2943);
nand U3964 (N_3964,N_2804,N_2405);
nor U3965 (N_3965,N_2497,N_2661);
or U3966 (N_3966,N_2836,N_2391);
and U3967 (N_3967,N_2155,N_2824);
nor U3968 (N_3968,N_2133,N_2044);
and U3969 (N_3969,N_2467,N_2596);
xor U3970 (N_3970,N_2586,N_2043);
xnor U3971 (N_3971,N_2672,N_2723);
nor U3972 (N_3972,N_2857,N_2693);
or U3973 (N_3973,N_2742,N_2263);
and U3974 (N_3974,N_2743,N_2206);
nor U3975 (N_3975,N_2475,N_2584);
nand U3976 (N_3976,N_2395,N_2596);
and U3977 (N_3977,N_2717,N_2362);
or U3978 (N_3978,N_2228,N_2295);
or U3979 (N_3979,N_2030,N_2764);
or U3980 (N_3980,N_2060,N_2020);
nor U3981 (N_3981,N_2181,N_2537);
xor U3982 (N_3982,N_2652,N_2578);
or U3983 (N_3983,N_2450,N_2489);
nand U3984 (N_3984,N_2805,N_2688);
nor U3985 (N_3985,N_2447,N_2395);
and U3986 (N_3986,N_2482,N_2524);
or U3987 (N_3987,N_2141,N_2667);
or U3988 (N_3988,N_2814,N_2746);
nand U3989 (N_3989,N_2478,N_2656);
or U3990 (N_3990,N_2434,N_2550);
xnor U3991 (N_3991,N_2641,N_2709);
and U3992 (N_3992,N_2548,N_2335);
xor U3993 (N_3993,N_2440,N_2821);
nand U3994 (N_3994,N_2581,N_2348);
nand U3995 (N_3995,N_2869,N_2992);
xor U3996 (N_3996,N_2113,N_2628);
xnor U3997 (N_3997,N_2749,N_2443);
nand U3998 (N_3998,N_2150,N_2321);
xor U3999 (N_3999,N_2770,N_2767);
or U4000 (N_4000,N_3621,N_3061);
xor U4001 (N_4001,N_3678,N_3471);
nor U4002 (N_4002,N_3766,N_3472);
xnor U4003 (N_4003,N_3223,N_3431);
nand U4004 (N_4004,N_3566,N_3434);
nor U4005 (N_4005,N_3830,N_3167);
xor U4006 (N_4006,N_3054,N_3803);
nor U4007 (N_4007,N_3522,N_3119);
nor U4008 (N_4008,N_3609,N_3599);
nor U4009 (N_4009,N_3221,N_3245);
nor U4010 (N_4010,N_3401,N_3352);
nor U4011 (N_4011,N_3982,N_3478);
xnor U4012 (N_4012,N_3856,N_3600);
and U4013 (N_4013,N_3244,N_3706);
xnor U4014 (N_4014,N_3376,N_3709);
xor U4015 (N_4015,N_3584,N_3332);
xnor U4016 (N_4016,N_3820,N_3722);
nor U4017 (N_4017,N_3065,N_3737);
nand U4018 (N_4018,N_3092,N_3105);
nand U4019 (N_4019,N_3439,N_3504);
and U4020 (N_4020,N_3035,N_3901);
xnor U4021 (N_4021,N_3057,N_3157);
or U4022 (N_4022,N_3151,N_3549);
and U4023 (N_4023,N_3028,N_3844);
and U4024 (N_4024,N_3289,N_3932);
or U4025 (N_4025,N_3337,N_3104);
and U4026 (N_4026,N_3215,N_3581);
or U4027 (N_4027,N_3835,N_3476);
or U4028 (N_4028,N_3624,N_3146);
nand U4029 (N_4029,N_3630,N_3275);
nor U4030 (N_4030,N_3214,N_3338);
nand U4031 (N_4031,N_3196,N_3456);
nand U4032 (N_4032,N_3865,N_3144);
or U4033 (N_4033,N_3169,N_3891);
nor U4034 (N_4034,N_3907,N_3642);
nor U4035 (N_4035,N_3479,N_3674);
xor U4036 (N_4036,N_3102,N_3178);
xor U4037 (N_4037,N_3062,N_3985);
nor U4038 (N_4038,N_3586,N_3738);
or U4039 (N_4039,N_3287,N_3646);
xor U4040 (N_4040,N_3895,N_3975);
nand U4041 (N_4041,N_3809,N_3233);
and U4042 (N_4042,N_3792,N_3121);
or U4043 (N_4043,N_3790,N_3445);
nand U4044 (N_4044,N_3539,N_3681);
nand U4045 (N_4045,N_3515,N_3429);
nor U4046 (N_4046,N_3415,N_3644);
and U4047 (N_4047,N_3817,N_3661);
or U4048 (N_4048,N_3075,N_3977);
xor U4049 (N_4049,N_3654,N_3371);
nand U4050 (N_4050,N_3968,N_3322);
xor U4051 (N_4051,N_3921,N_3508);
or U4052 (N_4052,N_3085,N_3055);
and U4053 (N_4053,N_3155,N_3514);
xnor U4054 (N_4054,N_3935,N_3220);
or U4055 (N_4055,N_3548,N_3318);
xnor U4056 (N_4056,N_3730,N_3695);
nand U4057 (N_4057,N_3484,N_3947);
and U4058 (N_4058,N_3779,N_3771);
or U4059 (N_4059,N_3818,N_3927);
xnor U4060 (N_4060,N_3353,N_3098);
and U4061 (N_4061,N_3474,N_3745);
and U4062 (N_4062,N_3978,N_3083);
xnor U4063 (N_4063,N_3093,N_3103);
or U4064 (N_4064,N_3385,N_3117);
or U4065 (N_4065,N_3726,N_3411);
nor U4066 (N_4066,N_3534,N_3242);
or U4067 (N_4067,N_3191,N_3870);
nor U4068 (N_4068,N_3410,N_3911);
nand U4069 (N_4069,N_3791,N_3127);
nor U4070 (N_4070,N_3979,N_3395);
nand U4071 (N_4071,N_3457,N_3109);
nand U4072 (N_4072,N_3056,N_3896);
nor U4073 (N_4073,N_3235,N_3816);
xor U4074 (N_4074,N_3645,N_3773);
xor U4075 (N_4075,N_3269,N_3443);
nor U4076 (N_4076,N_3620,N_3733);
nor U4077 (N_4077,N_3114,N_3304);
nor U4078 (N_4078,N_3789,N_3370);
nor U4079 (N_4079,N_3194,N_3461);
nor U4080 (N_4080,N_3604,N_3232);
nor U4081 (N_4081,N_3836,N_3675);
or U4082 (N_4082,N_3752,N_3428);
xnor U4083 (N_4083,N_3123,N_3750);
nor U4084 (N_4084,N_3349,N_3996);
or U4085 (N_4085,N_3305,N_3038);
nor U4086 (N_4086,N_3740,N_3128);
and U4087 (N_4087,N_3024,N_3329);
and U4088 (N_4088,N_3036,N_3639);
xor U4089 (N_4089,N_3552,N_3217);
or U4090 (N_4090,N_3433,N_3778);
nand U4091 (N_4091,N_3048,N_3701);
and U4092 (N_4092,N_3611,N_3783);
nor U4093 (N_4093,N_3717,N_3568);
xor U4094 (N_4094,N_3131,N_3142);
and U4095 (N_4095,N_3209,N_3689);
nand U4096 (N_4096,N_3130,N_3081);
and U4097 (N_4097,N_3828,N_3161);
xor U4098 (N_4098,N_3775,N_3523);
nor U4099 (N_4099,N_3893,N_3561);
xnor U4100 (N_4100,N_3704,N_3004);
xnor U4101 (N_4101,N_3833,N_3078);
nor U4102 (N_4102,N_3690,N_3501);
and U4103 (N_4103,N_3255,N_3852);
xnor U4104 (N_4104,N_3317,N_3197);
or U4105 (N_4105,N_3653,N_3832);
or U4106 (N_4106,N_3917,N_3139);
xnor U4107 (N_4107,N_3859,N_3010);
nor U4108 (N_4108,N_3551,N_3897);
nand U4109 (N_4109,N_3276,N_3188);
and U4110 (N_4110,N_3596,N_3403);
or U4111 (N_4111,N_3281,N_3475);
xnor U4112 (N_4112,N_3133,N_3166);
nor U4113 (N_4113,N_3040,N_3570);
or U4114 (N_4114,N_3351,N_3077);
xnor U4115 (N_4115,N_3041,N_3498);
nor U4116 (N_4116,N_3718,N_3741);
nor U4117 (N_4117,N_3212,N_3321);
xnor U4118 (N_4118,N_3615,N_3894);
or U4119 (N_4119,N_3601,N_3686);
nand U4120 (N_4120,N_3455,N_3361);
nor U4121 (N_4121,N_3770,N_3003);
xor U4122 (N_4122,N_3398,N_3268);
nand U4123 (N_4123,N_3988,N_3186);
or U4124 (N_4124,N_3889,N_3112);
xor U4125 (N_4125,N_3294,N_3619);
nor U4126 (N_4126,N_3559,N_3251);
or U4127 (N_4127,N_3617,N_3406);
or U4128 (N_4128,N_3152,N_3288);
nand U4129 (N_4129,N_3387,N_3449);
nor U4130 (N_4130,N_3134,N_3802);
nand U4131 (N_4131,N_3195,N_3684);
and U4132 (N_4132,N_3184,N_3796);
or U4133 (N_4133,N_3824,N_3165);
and U4134 (N_4134,N_3204,N_3373);
nor U4135 (N_4135,N_3107,N_3864);
or U4136 (N_4136,N_3125,N_3224);
or U4137 (N_4137,N_3392,N_3122);
xor U4138 (N_4138,N_3341,N_3282);
nor U4139 (N_4139,N_3538,N_3058);
nand U4140 (N_4140,N_3017,N_3583);
and U4141 (N_4141,N_3307,N_3231);
nand U4142 (N_4142,N_3437,N_3211);
nand U4143 (N_4143,N_3354,N_3997);
nor U4144 (N_4144,N_3399,N_3090);
nor U4145 (N_4145,N_3571,N_3120);
nand U4146 (N_4146,N_3272,N_3805);
xor U4147 (N_4147,N_3867,N_3569);
xor U4148 (N_4148,N_3416,N_3939);
or U4149 (N_4149,N_3525,N_3074);
or U4150 (N_4150,N_3958,N_3441);
or U4151 (N_4151,N_3814,N_3080);
xnor U4152 (N_4152,N_3933,N_3995);
xnor U4153 (N_4153,N_3340,N_3810);
nand U4154 (N_4154,N_3168,N_3452);
xnor U4155 (N_4155,N_3595,N_3407);
xnor U4156 (N_4156,N_3736,N_3855);
xnor U4157 (N_4157,N_3612,N_3831);
nand U4158 (N_4158,N_3762,N_3145);
and U4159 (N_4159,N_3348,N_3453);
xor U4160 (N_4160,N_3396,N_3821);
and U4161 (N_4161,N_3222,N_3488);
and U4162 (N_4162,N_3256,N_3328);
and U4163 (N_4163,N_3842,N_3823);
nand U4164 (N_4164,N_3034,N_3293);
nand U4165 (N_4165,N_3544,N_3362);
nor U4166 (N_4166,N_3862,N_3438);
nor U4167 (N_4167,N_3379,N_3528);
and U4168 (N_4168,N_3138,N_3286);
nor U4169 (N_4169,N_3170,N_3252);
or U4170 (N_4170,N_3193,N_3800);
nor U4171 (N_4171,N_3336,N_3537);
and U4172 (N_4172,N_3380,N_3598);
nor U4173 (N_4173,N_3798,N_3365);
or U4174 (N_4174,N_3384,N_3388);
and U4175 (N_4175,N_3160,N_3647);
xnor U4176 (N_4176,N_3719,N_3776);
and U4177 (N_4177,N_3210,N_3412);
xnor U4178 (N_4178,N_3531,N_3141);
and U4179 (N_4179,N_3749,N_3974);
nand U4180 (N_4180,N_3826,N_3914);
and U4181 (N_4181,N_3938,N_3989);
and U4182 (N_4182,N_3545,N_3807);
xnor U4183 (N_4183,N_3044,N_3285);
and U4184 (N_4184,N_3099,N_3442);
nand U4185 (N_4185,N_3963,N_3780);
xnor U4186 (N_4186,N_3393,N_3676);
xor U4187 (N_4187,N_3973,N_3339);
xor U4188 (N_4188,N_3192,N_3883);
or U4189 (N_4189,N_3553,N_3547);
nand U4190 (N_4190,N_3853,N_3582);
nand U4191 (N_4191,N_3513,N_3758);
or U4192 (N_4192,N_3179,N_3477);
or U4193 (N_4193,N_3705,N_3091);
nand U4194 (N_4194,N_3660,N_3019);
and U4195 (N_4195,N_3636,N_3880);
xor U4196 (N_4196,N_3970,N_3208);
nor U4197 (N_4197,N_3001,N_3687);
nand U4198 (N_4198,N_3665,N_3887);
or U4199 (N_4199,N_3769,N_3633);
nor U4200 (N_4200,N_3971,N_3774);
nand U4201 (N_4201,N_3804,N_3734);
and U4202 (N_4202,N_3651,N_3126);
nand U4203 (N_4203,N_3277,N_3900);
nand U4204 (N_4204,N_3436,N_3366);
or U4205 (N_4205,N_3858,N_3143);
nor U4206 (N_4206,N_3587,N_3378);
or U4207 (N_4207,N_3009,N_3301);
or U4208 (N_4208,N_3696,N_3190);
xnor U4209 (N_4209,N_3014,N_3068);
xnor U4210 (N_4210,N_3786,N_3180);
xor U4211 (N_4211,N_3657,N_3246);
xor U4212 (N_4212,N_3987,N_3567);
and U4213 (N_4213,N_3664,N_3331);
nand U4214 (N_4214,N_3735,N_3115);
xnor U4215 (N_4215,N_3391,N_3829);
xor U4216 (N_4216,N_3497,N_3714);
nand U4217 (N_4217,N_3618,N_3767);
nand U4218 (N_4218,N_3519,N_3656);
nor U4219 (N_4219,N_3259,N_3448);
or U4220 (N_4220,N_3808,N_3037);
and U4221 (N_4221,N_3755,N_3154);
nand U4222 (N_4222,N_3492,N_3863);
or U4223 (N_4223,N_3725,N_3482);
and U4224 (N_4224,N_3228,N_3173);
nand U4225 (N_4225,N_3147,N_3782);
and U4226 (N_4226,N_3822,N_3230);
and U4227 (N_4227,N_3781,N_3554);
and U4228 (N_4228,N_3266,N_3417);
xor U4229 (N_4229,N_3851,N_3811);
and U4230 (N_4230,N_3878,N_3008);
and U4231 (N_4231,N_3565,N_3588);
xor U4232 (N_4232,N_3465,N_3797);
nor U4233 (N_4233,N_3931,N_3011);
or U4234 (N_4234,N_3327,N_3953);
or U4235 (N_4235,N_3032,N_3861);
nor U4236 (N_4236,N_3291,N_3536);
nand U4237 (N_4237,N_3637,N_3788);
nand U4238 (N_4238,N_3206,N_3924);
and U4239 (N_4239,N_3335,N_3960);
or U4240 (N_4240,N_3980,N_3616);
or U4241 (N_4241,N_3319,N_3234);
xor U4242 (N_4242,N_3400,N_3659);
and U4243 (N_4243,N_3998,N_3350);
nand U4244 (N_4244,N_3849,N_3025);
or U4245 (N_4245,N_3007,N_3652);
and U4246 (N_4246,N_3892,N_3467);
xnor U4247 (N_4247,N_3540,N_3713);
nor U4248 (N_4248,N_3535,N_3423);
xor U4249 (N_4249,N_3840,N_3969);
nand U4250 (N_4250,N_3592,N_3261);
xnor U4251 (N_4251,N_3984,N_3238);
nand U4252 (N_4252,N_3216,N_3372);
and U4253 (N_4253,N_3941,N_3715);
or U4254 (N_4254,N_3493,N_3623);
nor U4255 (N_4255,N_3876,N_3203);
nor U4256 (N_4256,N_3723,N_3326);
and U4257 (N_4257,N_3521,N_3520);
xor U4258 (N_4258,N_3576,N_3382);
nand U4259 (N_4259,N_3063,N_3702);
nor U4260 (N_4260,N_3967,N_3156);
or U4261 (N_4261,N_3283,N_3346);
and U4262 (N_4262,N_3881,N_3879);
nand U4263 (N_4263,N_3280,N_3655);
and U4264 (N_4264,N_3869,N_3064);
xnor U4265 (N_4265,N_3033,N_3240);
nand U4266 (N_4266,N_3846,N_3672);
and U4267 (N_4267,N_3250,N_3763);
or U4268 (N_4268,N_3993,N_3700);
or U4269 (N_4269,N_3356,N_3377);
nand U4270 (N_4270,N_3183,N_3972);
or U4271 (N_4271,N_3005,N_3043);
or U4272 (N_4272,N_3765,N_3627);
nor U4273 (N_4273,N_3920,N_3854);
nor U4274 (N_4274,N_3267,N_3042);
or U4275 (N_4275,N_3450,N_3751);
nor U4276 (N_4276,N_3720,N_3868);
and U4277 (N_4277,N_3402,N_3589);
nor U4278 (N_4278,N_3698,N_3466);
xnor U4279 (N_4279,N_3628,N_3030);
nand U4280 (N_4280,N_3950,N_3047);
nor U4281 (N_4281,N_3296,N_3721);
and U4282 (N_4282,N_3097,N_3909);
xnor U4283 (N_4283,N_3526,N_3018);
xor U4284 (N_4284,N_3158,N_3490);
or U4285 (N_4285,N_3239,N_3507);
nand U4286 (N_4286,N_3787,N_3885);
nand U4287 (N_4287,N_3679,N_3111);
or U4288 (N_4288,N_3961,N_3839);
and U4289 (N_4289,N_3499,N_3952);
and U4290 (N_4290,N_3866,N_3594);
nor U4291 (N_4291,N_3946,N_3991);
xor U4292 (N_4292,N_3084,N_3913);
and U4293 (N_4293,N_3237,N_3243);
nand U4294 (N_4294,N_3638,N_3819);
or U4295 (N_4295,N_3279,N_3563);
nand U4296 (N_4296,N_3925,N_3505);
or U4297 (N_4297,N_3915,N_3494);
or U4298 (N_4298,N_3648,N_3013);
or U4299 (N_4299,N_3051,N_3650);
nand U4300 (N_4300,N_3470,N_3607);
nor U4301 (N_4301,N_3857,N_3330);
xnor U4302 (N_4302,N_3527,N_3390);
xor U4303 (N_4303,N_3405,N_3045);
nor U4304 (N_4304,N_3744,N_3027);
and U4305 (N_4305,N_3579,N_3124);
or U4306 (N_4306,N_3543,N_3550);
and U4307 (N_4307,N_3067,N_3573);
xor U4308 (N_4308,N_3945,N_3295);
and U4309 (N_4309,N_3608,N_3825);
nand U4310 (N_4310,N_3585,N_3072);
nand U4311 (N_4311,N_3426,N_3748);
or U4312 (N_4312,N_3070,N_3087);
and U4313 (N_4313,N_3605,N_3355);
nor U4314 (N_4314,N_3236,N_3937);
nor U4315 (N_4315,N_3556,N_3631);
nor U4316 (N_4316,N_3606,N_3760);
nand U4317 (N_4317,N_3089,N_3023);
nor U4318 (N_4318,N_3954,N_3205);
or U4319 (N_4319,N_3512,N_3136);
nor U4320 (N_4320,N_3575,N_3172);
or U4321 (N_4321,N_3884,N_3533);
nand U4322 (N_4322,N_3118,N_3308);
or U4323 (N_4323,N_3424,N_3936);
xnor U4324 (N_4324,N_3772,N_3274);
or U4325 (N_4325,N_3956,N_3200);
and U4326 (N_4326,N_3517,N_3872);
and U4327 (N_4327,N_3850,N_3218);
and U4328 (N_4328,N_3066,N_3847);
nand U4329 (N_4329,N_3688,N_3316);
or U4330 (N_4330,N_3060,N_3964);
nand U4331 (N_4331,N_3306,N_3368);
nand U4332 (N_4332,N_3207,N_3910);
and U4333 (N_4333,N_3082,N_3187);
and U4334 (N_4334,N_3496,N_3626);
and U4335 (N_4335,N_3100,N_3747);
nor U4336 (N_4336,N_3313,N_3990);
or U4337 (N_4337,N_3342,N_3464);
xnor U4338 (N_4338,N_3182,N_3634);
xor U4339 (N_4339,N_3271,N_3153);
nand U4340 (N_4340,N_3440,N_3603);
nor U4341 (N_4341,N_3577,N_3860);
and U4342 (N_4342,N_3164,N_3069);
or U4343 (N_4343,N_3462,N_3530);
nor U4344 (N_4344,N_3420,N_3999);
nand U4345 (N_4345,N_3265,N_3315);
and U4346 (N_4346,N_3247,N_3632);
nand U4347 (N_4347,N_3181,N_3677);
and U4348 (N_4348,N_3692,N_3270);
and U4349 (N_4349,N_3459,N_3957);
xnor U4350 (N_4350,N_3903,N_3454);
xor U4351 (N_4351,N_3290,N_3263);
and U4352 (N_4352,N_3435,N_3981);
nand U4353 (N_4353,N_3059,N_3140);
nand U4354 (N_4354,N_3959,N_3662);
nor U4355 (N_4355,N_3794,N_3345);
xnor U4356 (N_4356,N_3314,N_3591);
and U4357 (N_4357,N_3303,N_3712);
nand U4358 (N_4358,N_3463,N_3397);
xnor U4359 (N_4359,N_3815,N_3258);
xor U4360 (N_4360,N_3580,N_3095);
nor U4361 (N_4361,N_3015,N_3487);
nand U4362 (N_4362,N_3088,N_3837);
and U4363 (N_4363,N_3716,N_3310);
or U4364 (N_4364,N_3602,N_3202);
or U4365 (N_4365,N_3753,N_3162);
nor U4366 (N_4366,N_3694,N_3106);
nor U4367 (N_4367,N_3699,N_3229);
xor U4368 (N_4368,N_3572,N_3198);
or U4369 (N_4369,N_3046,N_3943);
or U4370 (N_4370,N_3666,N_3469);
and U4371 (N_4371,N_3050,N_3759);
and U4372 (N_4372,N_3079,N_3425);
xor U4373 (N_4373,N_3367,N_3020);
or U4374 (N_4374,N_3213,N_3300);
nand U4375 (N_4375,N_3890,N_3670);
and U4376 (N_4376,N_3076,N_3177);
and U4377 (N_4377,N_3578,N_3323);
and U4378 (N_4378,N_3249,N_3827);
or U4379 (N_4379,N_3635,N_3710);
xor U4380 (N_4380,N_3557,N_3026);
or U4381 (N_4381,N_3756,N_3312);
nand U4382 (N_4382,N_3375,N_3574);
or U4383 (N_4383,N_3622,N_3728);
or U4384 (N_4384,N_3148,N_3260);
or U4385 (N_4385,N_3625,N_3486);
nand U4386 (N_4386,N_3685,N_3359);
or U4387 (N_4387,N_3511,N_3297);
xor U4388 (N_4388,N_3386,N_3481);
nor U4389 (N_4389,N_3383,N_3813);
and U4390 (N_4390,N_3613,N_3944);
xnor U4391 (N_4391,N_3691,N_3006);
or U4392 (N_4392,N_3189,N_3875);
nand U4393 (N_4393,N_3558,N_3916);
and U4394 (N_4394,N_3962,N_3176);
nor U4395 (N_4395,N_3643,N_3649);
nand U4396 (N_4396,N_3668,N_3473);
or U4397 (N_4397,N_3500,N_3273);
and U4398 (N_4398,N_3149,N_3966);
xnor U4399 (N_4399,N_3309,N_3381);
xor U4400 (N_4400,N_3029,N_3711);
nor U4401 (N_4401,N_3754,N_3524);
xor U4402 (N_4402,N_3427,N_3793);
or U4403 (N_4403,N_3052,N_3311);
or U4404 (N_4404,N_3302,N_3784);
and U4405 (N_4405,N_3022,N_3801);
xnor U4406 (N_4406,N_3480,N_3697);
and U4407 (N_4407,N_3873,N_3510);
nor U4408 (N_4408,N_3983,N_3739);
nand U4409 (N_4409,N_3926,N_3389);
xor U4410 (N_4410,N_3732,N_3882);
nand U4411 (N_4411,N_3347,N_3845);
and U4412 (N_4412,N_3795,N_3363);
nand U4413 (N_4413,N_3923,N_3529);
and U4414 (N_4414,N_3799,N_3422);
nor U4415 (N_4415,N_3432,N_3680);
nand U4416 (N_4416,N_3053,N_3135);
nand U4417 (N_4417,N_3163,N_3000);
and U4418 (N_4418,N_3727,N_3408);
and U4419 (N_4419,N_3421,N_3409);
or U4420 (N_4420,N_3502,N_3226);
nor U4421 (N_4421,N_3564,N_3489);
nand U4422 (N_4422,N_3506,N_3159);
nor U4423 (N_4423,N_3743,N_3324);
or U4424 (N_4424,N_3418,N_3491);
xnor U4425 (N_4425,N_3468,N_3364);
nor U4426 (N_4426,N_3934,N_3344);
and U4427 (N_4427,N_3299,N_3451);
xor U4428 (N_4428,N_3369,N_3284);
or U4429 (N_4429,N_3278,N_3994);
and U4430 (N_4430,N_3404,N_3746);
nor U4431 (N_4431,N_3071,N_3012);
and U4432 (N_4432,N_3888,N_3485);
xor U4433 (N_4433,N_3460,N_3049);
nand U4434 (N_4434,N_3812,N_3227);
nand U4435 (N_4435,N_3641,N_3495);
nand U4436 (N_4436,N_3199,N_3593);
nor U4437 (N_4437,N_3039,N_3742);
xor U4438 (N_4438,N_3785,N_3683);
or U4439 (N_4439,N_3253,N_3663);
nor U4440 (N_4440,N_3262,N_3912);
nor U4441 (N_4441,N_3930,N_3562);
and U4442 (N_4442,N_3298,N_3871);
and U4443 (N_4443,N_3546,N_3016);
and U4444 (N_4444,N_3886,N_3116);
xor U4445 (N_4445,N_3841,N_3874);
xnor U4446 (N_4446,N_3357,N_3414);
or U4447 (N_4447,N_3419,N_3629);
and U4448 (N_4448,N_3877,N_3682);
nand U4449 (N_4449,N_3673,N_3949);
or U4450 (N_4450,N_3761,N_3174);
and U4451 (N_4451,N_3908,N_3031);
nor U4452 (N_4452,N_3986,N_3137);
or U4453 (N_4453,N_3708,N_3757);
and U4454 (N_4454,N_3768,N_3693);
nand U4455 (N_4455,N_3703,N_3320);
xor U4456 (N_4456,N_3430,N_3241);
nor U4457 (N_4457,N_3902,N_3671);
nand U4458 (N_4458,N_3248,N_3334);
and U4459 (N_4459,N_3110,N_3899);
nand U4460 (N_4460,N_3929,N_3948);
nand U4461 (N_4461,N_3976,N_3838);
nor U4462 (N_4462,N_3965,N_3132);
nand U4463 (N_4463,N_3094,N_3942);
xnor U4464 (N_4464,N_3992,N_3483);
and U4465 (N_4465,N_3928,N_3669);
xnor U4466 (N_4466,N_3590,N_3898);
nand U4467 (N_4467,N_3171,N_3843);
xnor U4468 (N_4468,N_3360,N_3560);
xor U4469 (N_4469,N_3518,N_3101);
nand U4470 (N_4470,N_3597,N_3904);
or U4471 (N_4471,N_3458,N_3185);
nor U4472 (N_4472,N_3922,N_3254);
nor U4473 (N_4473,N_3509,N_3096);
or U4474 (N_4474,N_3021,N_3150);
xor U4475 (N_4475,N_3358,N_3667);
and U4476 (N_4476,N_3731,N_3764);
and U4477 (N_4477,N_3175,N_3905);
nor U4478 (N_4478,N_3264,N_3325);
xnor U4479 (N_4479,N_3086,N_3918);
or U4480 (N_4480,N_3257,N_3541);
and U4481 (N_4481,N_3532,N_3446);
xor U4482 (N_4482,N_3940,N_3555);
nand U4483 (N_4483,N_3333,N_3729);
nand U4484 (N_4484,N_3129,N_3444);
and U4485 (N_4485,N_3503,N_3073);
nor U4486 (N_4486,N_3394,N_3919);
xnor U4487 (N_4487,N_3955,N_3834);
nor U4488 (N_4488,N_3951,N_3640);
xor U4489 (N_4489,N_3374,N_3658);
xor U4490 (N_4490,N_3542,N_3777);
or U4491 (N_4491,N_3002,N_3906);
and U4492 (N_4492,N_3113,N_3724);
nand U4493 (N_4493,N_3343,N_3516);
nand U4494 (N_4494,N_3806,N_3707);
or U4495 (N_4495,N_3848,N_3292);
xnor U4496 (N_4496,N_3201,N_3219);
nor U4497 (N_4497,N_3610,N_3108);
nand U4498 (N_4498,N_3225,N_3447);
nor U4499 (N_4499,N_3413,N_3614);
nor U4500 (N_4500,N_3402,N_3342);
or U4501 (N_4501,N_3733,N_3559);
nand U4502 (N_4502,N_3022,N_3562);
or U4503 (N_4503,N_3872,N_3185);
nor U4504 (N_4504,N_3072,N_3861);
nand U4505 (N_4505,N_3747,N_3316);
nor U4506 (N_4506,N_3579,N_3002);
or U4507 (N_4507,N_3558,N_3122);
nor U4508 (N_4508,N_3481,N_3652);
nand U4509 (N_4509,N_3441,N_3885);
and U4510 (N_4510,N_3000,N_3050);
nor U4511 (N_4511,N_3419,N_3692);
nand U4512 (N_4512,N_3857,N_3703);
xor U4513 (N_4513,N_3929,N_3895);
nor U4514 (N_4514,N_3520,N_3788);
xor U4515 (N_4515,N_3178,N_3903);
nand U4516 (N_4516,N_3293,N_3800);
nor U4517 (N_4517,N_3685,N_3658);
xnor U4518 (N_4518,N_3454,N_3132);
or U4519 (N_4519,N_3552,N_3560);
or U4520 (N_4520,N_3990,N_3987);
nand U4521 (N_4521,N_3816,N_3920);
or U4522 (N_4522,N_3931,N_3808);
xor U4523 (N_4523,N_3662,N_3696);
xor U4524 (N_4524,N_3803,N_3851);
nor U4525 (N_4525,N_3352,N_3533);
nand U4526 (N_4526,N_3659,N_3889);
and U4527 (N_4527,N_3353,N_3230);
and U4528 (N_4528,N_3684,N_3107);
nand U4529 (N_4529,N_3634,N_3206);
nor U4530 (N_4530,N_3887,N_3000);
nand U4531 (N_4531,N_3186,N_3420);
and U4532 (N_4532,N_3088,N_3907);
or U4533 (N_4533,N_3438,N_3085);
or U4534 (N_4534,N_3238,N_3792);
nor U4535 (N_4535,N_3375,N_3484);
nor U4536 (N_4536,N_3929,N_3610);
nand U4537 (N_4537,N_3700,N_3635);
nor U4538 (N_4538,N_3108,N_3998);
nand U4539 (N_4539,N_3488,N_3677);
or U4540 (N_4540,N_3949,N_3179);
nor U4541 (N_4541,N_3567,N_3859);
nor U4542 (N_4542,N_3265,N_3126);
xnor U4543 (N_4543,N_3800,N_3861);
xnor U4544 (N_4544,N_3595,N_3164);
and U4545 (N_4545,N_3750,N_3451);
nand U4546 (N_4546,N_3492,N_3596);
and U4547 (N_4547,N_3367,N_3350);
or U4548 (N_4548,N_3921,N_3997);
nor U4549 (N_4549,N_3886,N_3897);
and U4550 (N_4550,N_3854,N_3626);
or U4551 (N_4551,N_3793,N_3885);
nor U4552 (N_4552,N_3966,N_3672);
or U4553 (N_4553,N_3964,N_3755);
nand U4554 (N_4554,N_3136,N_3435);
xor U4555 (N_4555,N_3254,N_3965);
xnor U4556 (N_4556,N_3360,N_3673);
nor U4557 (N_4557,N_3293,N_3305);
nor U4558 (N_4558,N_3122,N_3195);
or U4559 (N_4559,N_3803,N_3536);
nor U4560 (N_4560,N_3451,N_3821);
nand U4561 (N_4561,N_3218,N_3723);
nand U4562 (N_4562,N_3308,N_3718);
or U4563 (N_4563,N_3825,N_3175);
nand U4564 (N_4564,N_3451,N_3418);
and U4565 (N_4565,N_3234,N_3165);
nand U4566 (N_4566,N_3444,N_3581);
or U4567 (N_4567,N_3544,N_3013);
xor U4568 (N_4568,N_3952,N_3676);
or U4569 (N_4569,N_3793,N_3705);
xor U4570 (N_4570,N_3723,N_3890);
xnor U4571 (N_4571,N_3297,N_3641);
nor U4572 (N_4572,N_3862,N_3470);
nand U4573 (N_4573,N_3942,N_3694);
nand U4574 (N_4574,N_3250,N_3805);
nand U4575 (N_4575,N_3386,N_3422);
nand U4576 (N_4576,N_3392,N_3226);
and U4577 (N_4577,N_3061,N_3579);
or U4578 (N_4578,N_3591,N_3013);
nand U4579 (N_4579,N_3486,N_3161);
or U4580 (N_4580,N_3134,N_3044);
nor U4581 (N_4581,N_3556,N_3261);
xor U4582 (N_4582,N_3341,N_3819);
or U4583 (N_4583,N_3605,N_3377);
nor U4584 (N_4584,N_3989,N_3863);
or U4585 (N_4585,N_3408,N_3774);
and U4586 (N_4586,N_3613,N_3209);
xor U4587 (N_4587,N_3381,N_3825);
or U4588 (N_4588,N_3688,N_3590);
xnor U4589 (N_4589,N_3275,N_3299);
nand U4590 (N_4590,N_3190,N_3987);
xnor U4591 (N_4591,N_3735,N_3753);
nand U4592 (N_4592,N_3421,N_3284);
nand U4593 (N_4593,N_3615,N_3318);
nor U4594 (N_4594,N_3980,N_3776);
and U4595 (N_4595,N_3293,N_3585);
and U4596 (N_4596,N_3188,N_3389);
and U4597 (N_4597,N_3792,N_3132);
or U4598 (N_4598,N_3267,N_3552);
and U4599 (N_4599,N_3398,N_3219);
and U4600 (N_4600,N_3474,N_3040);
xor U4601 (N_4601,N_3334,N_3546);
nand U4602 (N_4602,N_3673,N_3645);
nand U4603 (N_4603,N_3151,N_3413);
nor U4604 (N_4604,N_3533,N_3902);
nor U4605 (N_4605,N_3401,N_3218);
and U4606 (N_4606,N_3664,N_3830);
nand U4607 (N_4607,N_3742,N_3275);
and U4608 (N_4608,N_3029,N_3203);
xor U4609 (N_4609,N_3525,N_3581);
nor U4610 (N_4610,N_3673,N_3038);
nor U4611 (N_4611,N_3241,N_3912);
and U4612 (N_4612,N_3294,N_3618);
xor U4613 (N_4613,N_3709,N_3247);
and U4614 (N_4614,N_3076,N_3009);
nand U4615 (N_4615,N_3292,N_3463);
nand U4616 (N_4616,N_3545,N_3038);
or U4617 (N_4617,N_3078,N_3746);
nand U4618 (N_4618,N_3638,N_3439);
nand U4619 (N_4619,N_3059,N_3519);
xor U4620 (N_4620,N_3609,N_3185);
nand U4621 (N_4621,N_3313,N_3655);
nor U4622 (N_4622,N_3040,N_3008);
nor U4623 (N_4623,N_3783,N_3498);
or U4624 (N_4624,N_3831,N_3217);
nor U4625 (N_4625,N_3557,N_3340);
xor U4626 (N_4626,N_3278,N_3870);
nand U4627 (N_4627,N_3620,N_3827);
or U4628 (N_4628,N_3047,N_3728);
nand U4629 (N_4629,N_3558,N_3205);
or U4630 (N_4630,N_3020,N_3863);
xnor U4631 (N_4631,N_3891,N_3503);
nand U4632 (N_4632,N_3500,N_3289);
nand U4633 (N_4633,N_3622,N_3243);
xor U4634 (N_4634,N_3868,N_3555);
and U4635 (N_4635,N_3734,N_3662);
xnor U4636 (N_4636,N_3354,N_3512);
and U4637 (N_4637,N_3344,N_3227);
nand U4638 (N_4638,N_3364,N_3056);
and U4639 (N_4639,N_3686,N_3703);
xnor U4640 (N_4640,N_3048,N_3053);
and U4641 (N_4641,N_3932,N_3122);
and U4642 (N_4642,N_3290,N_3102);
nor U4643 (N_4643,N_3680,N_3585);
nor U4644 (N_4644,N_3418,N_3940);
nand U4645 (N_4645,N_3387,N_3819);
nor U4646 (N_4646,N_3388,N_3833);
nand U4647 (N_4647,N_3874,N_3628);
and U4648 (N_4648,N_3035,N_3308);
xor U4649 (N_4649,N_3931,N_3580);
or U4650 (N_4650,N_3634,N_3468);
nor U4651 (N_4651,N_3275,N_3185);
or U4652 (N_4652,N_3375,N_3120);
and U4653 (N_4653,N_3413,N_3385);
nor U4654 (N_4654,N_3132,N_3353);
xor U4655 (N_4655,N_3788,N_3638);
nor U4656 (N_4656,N_3761,N_3255);
nor U4657 (N_4657,N_3100,N_3689);
nor U4658 (N_4658,N_3882,N_3183);
and U4659 (N_4659,N_3225,N_3998);
and U4660 (N_4660,N_3074,N_3655);
and U4661 (N_4661,N_3569,N_3922);
nand U4662 (N_4662,N_3672,N_3274);
and U4663 (N_4663,N_3239,N_3488);
nand U4664 (N_4664,N_3493,N_3873);
nor U4665 (N_4665,N_3530,N_3005);
and U4666 (N_4666,N_3021,N_3419);
or U4667 (N_4667,N_3780,N_3602);
nand U4668 (N_4668,N_3572,N_3382);
xnor U4669 (N_4669,N_3495,N_3365);
and U4670 (N_4670,N_3321,N_3627);
xnor U4671 (N_4671,N_3017,N_3902);
xor U4672 (N_4672,N_3516,N_3980);
or U4673 (N_4673,N_3560,N_3257);
or U4674 (N_4674,N_3515,N_3093);
xnor U4675 (N_4675,N_3661,N_3885);
nor U4676 (N_4676,N_3892,N_3748);
nand U4677 (N_4677,N_3855,N_3349);
and U4678 (N_4678,N_3154,N_3370);
and U4679 (N_4679,N_3874,N_3402);
or U4680 (N_4680,N_3123,N_3292);
xor U4681 (N_4681,N_3588,N_3359);
and U4682 (N_4682,N_3214,N_3456);
nand U4683 (N_4683,N_3095,N_3783);
or U4684 (N_4684,N_3862,N_3783);
or U4685 (N_4685,N_3781,N_3030);
or U4686 (N_4686,N_3060,N_3349);
xor U4687 (N_4687,N_3808,N_3153);
and U4688 (N_4688,N_3401,N_3577);
and U4689 (N_4689,N_3359,N_3159);
nand U4690 (N_4690,N_3794,N_3109);
xnor U4691 (N_4691,N_3101,N_3745);
nand U4692 (N_4692,N_3006,N_3202);
and U4693 (N_4693,N_3705,N_3305);
nand U4694 (N_4694,N_3306,N_3936);
xnor U4695 (N_4695,N_3202,N_3846);
nand U4696 (N_4696,N_3709,N_3627);
xnor U4697 (N_4697,N_3618,N_3408);
and U4698 (N_4698,N_3164,N_3756);
or U4699 (N_4699,N_3982,N_3174);
nand U4700 (N_4700,N_3341,N_3782);
xnor U4701 (N_4701,N_3759,N_3636);
and U4702 (N_4702,N_3809,N_3616);
xor U4703 (N_4703,N_3392,N_3611);
or U4704 (N_4704,N_3226,N_3775);
nand U4705 (N_4705,N_3573,N_3887);
nand U4706 (N_4706,N_3265,N_3783);
or U4707 (N_4707,N_3528,N_3164);
or U4708 (N_4708,N_3507,N_3260);
or U4709 (N_4709,N_3343,N_3660);
and U4710 (N_4710,N_3697,N_3232);
nand U4711 (N_4711,N_3979,N_3750);
nand U4712 (N_4712,N_3579,N_3762);
and U4713 (N_4713,N_3614,N_3990);
nor U4714 (N_4714,N_3680,N_3019);
and U4715 (N_4715,N_3513,N_3304);
nor U4716 (N_4716,N_3954,N_3877);
nor U4717 (N_4717,N_3244,N_3981);
xor U4718 (N_4718,N_3292,N_3183);
and U4719 (N_4719,N_3507,N_3179);
nand U4720 (N_4720,N_3260,N_3937);
and U4721 (N_4721,N_3998,N_3901);
and U4722 (N_4722,N_3110,N_3936);
or U4723 (N_4723,N_3729,N_3209);
nor U4724 (N_4724,N_3515,N_3131);
nand U4725 (N_4725,N_3357,N_3313);
and U4726 (N_4726,N_3507,N_3232);
nor U4727 (N_4727,N_3272,N_3861);
or U4728 (N_4728,N_3754,N_3703);
and U4729 (N_4729,N_3889,N_3002);
and U4730 (N_4730,N_3306,N_3891);
xnor U4731 (N_4731,N_3134,N_3942);
nor U4732 (N_4732,N_3014,N_3995);
xor U4733 (N_4733,N_3792,N_3874);
nor U4734 (N_4734,N_3674,N_3401);
nor U4735 (N_4735,N_3222,N_3441);
nor U4736 (N_4736,N_3738,N_3184);
or U4737 (N_4737,N_3021,N_3998);
and U4738 (N_4738,N_3349,N_3319);
nor U4739 (N_4739,N_3878,N_3762);
xnor U4740 (N_4740,N_3064,N_3893);
nor U4741 (N_4741,N_3125,N_3884);
xnor U4742 (N_4742,N_3891,N_3579);
and U4743 (N_4743,N_3178,N_3675);
nand U4744 (N_4744,N_3758,N_3337);
nor U4745 (N_4745,N_3899,N_3483);
xor U4746 (N_4746,N_3309,N_3154);
nand U4747 (N_4747,N_3879,N_3595);
nor U4748 (N_4748,N_3957,N_3555);
or U4749 (N_4749,N_3270,N_3646);
or U4750 (N_4750,N_3490,N_3655);
or U4751 (N_4751,N_3251,N_3341);
nor U4752 (N_4752,N_3261,N_3120);
nand U4753 (N_4753,N_3819,N_3002);
nor U4754 (N_4754,N_3140,N_3362);
nand U4755 (N_4755,N_3240,N_3142);
nor U4756 (N_4756,N_3275,N_3658);
nand U4757 (N_4757,N_3481,N_3522);
nand U4758 (N_4758,N_3196,N_3014);
and U4759 (N_4759,N_3857,N_3092);
nor U4760 (N_4760,N_3226,N_3901);
nor U4761 (N_4761,N_3667,N_3155);
and U4762 (N_4762,N_3958,N_3654);
or U4763 (N_4763,N_3772,N_3601);
nand U4764 (N_4764,N_3212,N_3391);
xnor U4765 (N_4765,N_3544,N_3454);
nand U4766 (N_4766,N_3522,N_3900);
nand U4767 (N_4767,N_3152,N_3835);
xnor U4768 (N_4768,N_3879,N_3863);
nor U4769 (N_4769,N_3388,N_3004);
xor U4770 (N_4770,N_3864,N_3318);
xor U4771 (N_4771,N_3771,N_3984);
and U4772 (N_4772,N_3530,N_3145);
nor U4773 (N_4773,N_3900,N_3406);
or U4774 (N_4774,N_3587,N_3960);
nor U4775 (N_4775,N_3583,N_3169);
nor U4776 (N_4776,N_3255,N_3529);
and U4777 (N_4777,N_3226,N_3168);
nor U4778 (N_4778,N_3457,N_3104);
and U4779 (N_4779,N_3160,N_3862);
nand U4780 (N_4780,N_3946,N_3339);
xnor U4781 (N_4781,N_3216,N_3718);
nand U4782 (N_4782,N_3321,N_3426);
nand U4783 (N_4783,N_3770,N_3448);
nor U4784 (N_4784,N_3668,N_3020);
and U4785 (N_4785,N_3995,N_3065);
xor U4786 (N_4786,N_3467,N_3861);
and U4787 (N_4787,N_3630,N_3357);
or U4788 (N_4788,N_3779,N_3609);
or U4789 (N_4789,N_3564,N_3348);
nand U4790 (N_4790,N_3657,N_3121);
nand U4791 (N_4791,N_3692,N_3326);
or U4792 (N_4792,N_3172,N_3881);
and U4793 (N_4793,N_3696,N_3576);
or U4794 (N_4794,N_3278,N_3630);
or U4795 (N_4795,N_3411,N_3037);
or U4796 (N_4796,N_3414,N_3691);
and U4797 (N_4797,N_3722,N_3501);
xor U4798 (N_4798,N_3531,N_3881);
or U4799 (N_4799,N_3462,N_3715);
nor U4800 (N_4800,N_3017,N_3252);
xnor U4801 (N_4801,N_3541,N_3235);
xor U4802 (N_4802,N_3474,N_3556);
nor U4803 (N_4803,N_3831,N_3868);
xor U4804 (N_4804,N_3896,N_3458);
nor U4805 (N_4805,N_3355,N_3912);
nor U4806 (N_4806,N_3639,N_3616);
and U4807 (N_4807,N_3899,N_3902);
xnor U4808 (N_4808,N_3164,N_3072);
and U4809 (N_4809,N_3257,N_3150);
nor U4810 (N_4810,N_3336,N_3255);
nor U4811 (N_4811,N_3427,N_3645);
nor U4812 (N_4812,N_3621,N_3995);
xor U4813 (N_4813,N_3492,N_3514);
xor U4814 (N_4814,N_3339,N_3830);
nor U4815 (N_4815,N_3613,N_3471);
xnor U4816 (N_4816,N_3914,N_3699);
nand U4817 (N_4817,N_3246,N_3096);
nand U4818 (N_4818,N_3100,N_3995);
and U4819 (N_4819,N_3195,N_3307);
nor U4820 (N_4820,N_3095,N_3921);
xor U4821 (N_4821,N_3125,N_3999);
nand U4822 (N_4822,N_3029,N_3177);
nor U4823 (N_4823,N_3829,N_3725);
xor U4824 (N_4824,N_3764,N_3889);
xnor U4825 (N_4825,N_3886,N_3492);
nand U4826 (N_4826,N_3624,N_3026);
and U4827 (N_4827,N_3349,N_3372);
or U4828 (N_4828,N_3474,N_3828);
and U4829 (N_4829,N_3462,N_3714);
xor U4830 (N_4830,N_3346,N_3144);
or U4831 (N_4831,N_3755,N_3553);
or U4832 (N_4832,N_3698,N_3981);
and U4833 (N_4833,N_3535,N_3367);
and U4834 (N_4834,N_3970,N_3665);
or U4835 (N_4835,N_3304,N_3321);
nor U4836 (N_4836,N_3132,N_3488);
or U4837 (N_4837,N_3429,N_3836);
nor U4838 (N_4838,N_3908,N_3729);
nor U4839 (N_4839,N_3938,N_3347);
nand U4840 (N_4840,N_3341,N_3887);
or U4841 (N_4841,N_3090,N_3001);
and U4842 (N_4842,N_3418,N_3317);
nor U4843 (N_4843,N_3650,N_3958);
nor U4844 (N_4844,N_3926,N_3316);
xor U4845 (N_4845,N_3852,N_3922);
nor U4846 (N_4846,N_3680,N_3102);
nand U4847 (N_4847,N_3476,N_3348);
and U4848 (N_4848,N_3851,N_3116);
nor U4849 (N_4849,N_3659,N_3777);
nor U4850 (N_4850,N_3110,N_3237);
nand U4851 (N_4851,N_3650,N_3901);
xor U4852 (N_4852,N_3870,N_3190);
and U4853 (N_4853,N_3295,N_3100);
nand U4854 (N_4854,N_3708,N_3495);
nand U4855 (N_4855,N_3035,N_3565);
xnor U4856 (N_4856,N_3352,N_3136);
nand U4857 (N_4857,N_3509,N_3319);
xnor U4858 (N_4858,N_3807,N_3216);
xor U4859 (N_4859,N_3492,N_3079);
nor U4860 (N_4860,N_3560,N_3060);
nor U4861 (N_4861,N_3522,N_3953);
xor U4862 (N_4862,N_3560,N_3182);
nor U4863 (N_4863,N_3588,N_3461);
and U4864 (N_4864,N_3631,N_3468);
xor U4865 (N_4865,N_3283,N_3997);
nand U4866 (N_4866,N_3515,N_3996);
xnor U4867 (N_4867,N_3041,N_3241);
xnor U4868 (N_4868,N_3889,N_3629);
and U4869 (N_4869,N_3856,N_3480);
and U4870 (N_4870,N_3794,N_3863);
nand U4871 (N_4871,N_3913,N_3027);
or U4872 (N_4872,N_3730,N_3655);
nand U4873 (N_4873,N_3486,N_3110);
or U4874 (N_4874,N_3585,N_3825);
and U4875 (N_4875,N_3334,N_3407);
nor U4876 (N_4876,N_3426,N_3799);
or U4877 (N_4877,N_3004,N_3961);
and U4878 (N_4878,N_3297,N_3670);
and U4879 (N_4879,N_3857,N_3631);
nor U4880 (N_4880,N_3806,N_3402);
or U4881 (N_4881,N_3491,N_3420);
and U4882 (N_4882,N_3193,N_3958);
xor U4883 (N_4883,N_3761,N_3418);
and U4884 (N_4884,N_3217,N_3878);
or U4885 (N_4885,N_3395,N_3313);
xnor U4886 (N_4886,N_3086,N_3148);
xnor U4887 (N_4887,N_3748,N_3225);
and U4888 (N_4888,N_3588,N_3042);
or U4889 (N_4889,N_3123,N_3487);
nor U4890 (N_4890,N_3005,N_3993);
or U4891 (N_4891,N_3147,N_3508);
nand U4892 (N_4892,N_3491,N_3615);
or U4893 (N_4893,N_3685,N_3553);
nand U4894 (N_4894,N_3750,N_3367);
nand U4895 (N_4895,N_3916,N_3123);
xnor U4896 (N_4896,N_3813,N_3232);
xnor U4897 (N_4897,N_3261,N_3527);
and U4898 (N_4898,N_3730,N_3684);
xnor U4899 (N_4899,N_3002,N_3411);
and U4900 (N_4900,N_3776,N_3771);
xnor U4901 (N_4901,N_3666,N_3163);
nand U4902 (N_4902,N_3516,N_3878);
nand U4903 (N_4903,N_3084,N_3931);
and U4904 (N_4904,N_3464,N_3116);
nor U4905 (N_4905,N_3421,N_3066);
or U4906 (N_4906,N_3577,N_3774);
nand U4907 (N_4907,N_3320,N_3051);
xor U4908 (N_4908,N_3994,N_3908);
and U4909 (N_4909,N_3708,N_3037);
xnor U4910 (N_4910,N_3088,N_3612);
xnor U4911 (N_4911,N_3459,N_3904);
and U4912 (N_4912,N_3185,N_3364);
xnor U4913 (N_4913,N_3898,N_3970);
nand U4914 (N_4914,N_3166,N_3282);
or U4915 (N_4915,N_3882,N_3743);
and U4916 (N_4916,N_3671,N_3456);
and U4917 (N_4917,N_3311,N_3062);
and U4918 (N_4918,N_3033,N_3628);
xor U4919 (N_4919,N_3711,N_3555);
xnor U4920 (N_4920,N_3039,N_3130);
and U4921 (N_4921,N_3781,N_3525);
xor U4922 (N_4922,N_3660,N_3209);
xnor U4923 (N_4923,N_3376,N_3247);
or U4924 (N_4924,N_3066,N_3566);
nor U4925 (N_4925,N_3328,N_3978);
or U4926 (N_4926,N_3545,N_3662);
or U4927 (N_4927,N_3295,N_3988);
nor U4928 (N_4928,N_3464,N_3432);
nor U4929 (N_4929,N_3725,N_3234);
nor U4930 (N_4930,N_3427,N_3058);
and U4931 (N_4931,N_3249,N_3578);
or U4932 (N_4932,N_3783,N_3232);
or U4933 (N_4933,N_3204,N_3134);
and U4934 (N_4934,N_3979,N_3325);
nand U4935 (N_4935,N_3307,N_3610);
or U4936 (N_4936,N_3502,N_3629);
xnor U4937 (N_4937,N_3684,N_3716);
xor U4938 (N_4938,N_3209,N_3226);
and U4939 (N_4939,N_3741,N_3610);
and U4940 (N_4940,N_3236,N_3520);
xnor U4941 (N_4941,N_3264,N_3814);
or U4942 (N_4942,N_3334,N_3622);
nor U4943 (N_4943,N_3019,N_3323);
nor U4944 (N_4944,N_3346,N_3366);
and U4945 (N_4945,N_3809,N_3647);
nand U4946 (N_4946,N_3084,N_3832);
and U4947 (N_4947,N_3888,N_3296);
or U4948 (N_4948,N_3749,N_3366);
xor U4949 (N_4949,N_3271,N_3047);
nand U4950 (N_4950,N_3079,N_3212);
xnor U4951 (N_4951,N_3836,N_3814);
nor U4952 (N_4952,N_3732,N_3008);
and U4953 (N_4953,N_3229,N_3611);
nor U4954 (N_4954,N_3735,N_3913);
or U4955 (N_4955,N_3751,N_3935);
or U4956 (N_4956,N_3033,N_3737);
or U4957 (N_4957,N_3093,N_3461);
xor U4958 (N_4958,N_3221,N_3087);
and U4959 (N_4959,N_3163,N_3126);
nor U4960 (N_4960,N_3104,N_3734);
and U4961 (N_4961,N_3810,N_3931);
xnor U4962 (N_4962,N_3839,N_3723);
xor U4963 (N_4963,N_3493,N_3398);
nor U4964 (N_4964,N_3514,N_3322);
or U4965 (N_4965,N_3892,N_3220);
nand U4966 (N_4966,N_3301,N_3234);
nor U4967 (N_4967,N_3429,N_3350);
xor U4968 (N_4968,N_3306,N_3457);
and U4969 (N_4969,N_3259,N_3619);
or U4970 (N_4970,N_3736,N_3983);
and U4971 (N_4971,N_3182,N_3781);
nor U4972 (N_4972,N_3642,N_3334);
nand U4973 (N_4973,N_3478,N_3727);
xnor U4974 (N_4974,N_3105,N_3144);
and U4975 (N_4975,N_3457,N_3801);
or U4976 (N_4976,N_3265,N_3782);
and U4977 (N_4977,N_3732,N_3055);
nor U4978 (N_4978,N_3469,N_3981);
and U4979 (N_4979,N_3480,N_3661);
nor U4980 (N_4980,N_3073,N_3207);
nor U4981 (N_4981,N_3153,N_3617);
or U4982 (N_4982,N_3826,N_3313);
nand U4983 (N_4983,N_3719,N_3342);
nor U4984 (N_4984,N_3413,N_3880);
nor U4985 (N_4985,N_3476,N_3496);
nand U4986 (N_4986,N_3007,N_3399);
xor U4987 (N_4987,N_3046,N_3242);
nor U4988 (N_4988,N_3664,N_3418);
or U4989 (N_4989,N_3883,N_3661);
xnor U4990 (N_4990,N_3184,N_3467);
and U4991 (N_4991,N_3541,N_3272);
and U4992 (N_4992,N_3357,N_3574);
and U4993 (N_4993,N_3135,N_3503);
nand U4994 (N_4994,N_3442,N_3918);
nand U4995 (N_4995,N_3355,N_3059);
nand U4996 (N_4996,N_3554,N_3650);
nand U4997 (N_4997,N_3857,N_3117);
and U4998 (N_4998,N_3993,N_3417);
nor U4999 (N_4999,N_3314,N_3876);
xor U5000 (N_5000,N_4889,N_4663);
nand U5001 (N_5001,N_4035,N_4400);
nor U5002 (N_5002,N_4947,N_4188);
xnor U5003 (N_5003,N_4315,N_4955);
nor U5004 (N_5004,N_4182,N_4245);
or U5005 (N_5005,N_4166,N_4980);
xor U5006 (N_5006,N_4375,N_4202);
or U5007 (N_5007,N_4384,N_4687);
nand U5008 (N_5008,N_4366,N_4819);
nand U5009 (N_5009,N_4354,N_4149);
and U5010 (N_5010,N_4544,N_4521);
or U5011 (N_5011,N_4279,N_4068);
nand U5012 (N_5012,N_4714,N_4923);
xor U5013 (N_5013,N_4434,N_4455);
xor U5014 (N_5014,N_4535,N_4514);
nor U5015 (N_5015,N_4566,N_4957);
nor U5016 (N_5016,N_4837,N_4284);
and U5017 (N_5017,N_4854,N_4715);
or U5018 (N_5018,N_4700,N_4849);
nor U5019 (N_5019,N_4757,N_4492);
xnor U5020 (N_5020,N_4822,N_4355);
nand U5021 (N_5021,N_4960,N_4285);
or U5022 (N_5022,N_4786,N_4417);
xnor U5023 (N_5023,N_4193,N_4563);
nand U5024 (N_5024,N_4716,N_4790);
xnor U5025 (N_5025,N_4495,N_4728);
and U5026 (N_5026,N_4327,N_4292);
nor U5027 (N_5027,N_4989,N_4684);
or U5028 (N_5028,N_4802,N_4922);
or U5029 (N_5029,N_4621,N_4964);
or U5030 (N_5030,N_4228,N_4640);
and U5031 (N_5031,N_4737,N_4456);
xnor U5032 (N_5032,N_4598,N_4224);
and U5033 (N_5033,N_4209,N_4704);
or U5034 (N_5034,N_4868,N_4530);
and U5035 (N_5035,N_4606,N_4734);
xnor U5036 (N_5036,N_4860,N_4576);
nor U5037 (N_5037,N_4558,N_4498);
xor U5038 (N_5038,N_4537,N_4690);
and U5039 (N_5039,N_4471,N_4447);
nand U5040 (N_5040,N_4472,N_4045);
xor U5041 (N_5041,N_4438,N_4759);
nor U5042 (N_5042,N_4599,N_4641);
or U5043 (N_5043,N_4446,N_4985);
nor U5044 (N_5044,N_4042,N_4454);
or U5045 (N_5045,N_4164,N_4928);
xor U5046 (N_5046,N_4775,N_4741);
nand U5047 (N_5047,N_4114,N_4143);
nand U5048 (N_5048,N_4970,N_4835);
and U5049 (N_5049,N_4177,N_4738);
nor U5050 (N_5050,N_4256,N_4672);
xor U5051 (N_5051,N_4811,N_4482);
and U5052 (N_5052,N_4917,N_4317);
nor U5053 (N_5053,N_4264,N_4605);
xor U5054 (N_5054,N_4887,N_4688);
or U5055 (N_5055,N_4910,N_4953);
xor U5056 (N_5056,N_4705,N_4581);
and U5057 (N_5057,N_4654,N_4797);
or U5058 (N_5058,N_4394,N_4773);
or U5059 (N_5059,N_4286,N_4020);
xnor U5060 (N_5060,N_4069,N_4719);
and U5061 (N_5061,N_4280,N_4548);
nor U5062 (N_5062,N_4866,N_4150);
nand U5063 (N_5063,N_4679,N_4274);
or U5064 (N_5064,N_4230,N_4508);
xor U5065 (N_5065,N_4639,N_4263);
nand U5066 (N_5066,N_4401,N_4404);
or U5067 (N_5067,N_4695,N_4983);
nor U5068 (N_5068,N_4670,N_4380);
and U5069 (N_5069,N_4839,N_4706);
nand U5070 (N_5070,N_4457,N_4419);
or U5071 (N_5071,N_4927,N_4736);
xor U5072 (N_5072,N_4485,N_4374);
or U5073 (N_5073,N_4332,N_4435);
nand U5074 (N_5074,N_4626,N_4818);
nor U5075 (N_5075,N_4016,N_4179);
or U5076 (N_5076,N_4678,N_4160);
xnor U5077 (N_5077,N_4119,N_4258);
or U5078 (N_5078,N_4403,N_4727);
or U5079 (N_5079,N_4386,N_4013);
and U5080 (N_5080,N_4395,N_4021);
nor U5081 (N_5081,N_4081,N_4667);
or U5082 (N_5082,N_4210,N_4600);
or U5083 (N_5083,N_4616,N_4359);
nand U5084 (N_5084,N_4565,N_4223);
xor U5085 (N_5085,N_4681,N_4270);
or U5086 (N_5086,N_4437,N_4466);
and U5087 (N_5087,N_4049,N_4615);
and U5088 (N_5088,N_4992,N_4052);
xnor U5089 (N_5089,N_4310,N_4560);
or U5090 (N_5090,N_4618,N_4763);
nand U5091 (N_5091,N_4542,N_4623);
xor U5092 (N_5092,N_4901,N_4844);
xnor U5093 (N_5093,N_4717,N_4314);
nor U5094 (N_5094,N_4668,N_4662);
nand U5095 (N_5095,N_4468,N_4268);
and U5096 (N_5096,N_4415,N_4793);
nor U5097 (N_5097,N_4489,N_4774);
and U5098 (N_5098,N_4307,N_4720);
xnor U5099 (N_5099,N_4702,N_4554);
nor U5100 (N_5100,N_4283,N_4557);
nor U5101 (N_5101,N_4147,N_4628);
nand U5102 (N_5102,N_4078,N_4969);
xnor U5103 (N_5103,N_4102,N_4750);
and U5104 (N_5104,N_4301,N_4219);
xor U5105 (N_5105,N_4298,N_4841);
or U5106 (N_5106,N_4816,N_4065);
nor U5107 (N_5107,N_4007,N_4490);
xnor U5108 (N_5108,N_4347,N_4361);
xor U5109 (N_5109,N_4154,N_4429);
xor U5110 (N_5110,N_4194,N_4171);
and U5111 (N_5111,N_4729,N_4241);
and U5112 (N_5112,N_4026,N_4523);
nor U5113 (N_5113,N_4879,N_4617);
or U5114 (N_5114,N_4784,N_4755);
nor U5115 (N_5115,N_4915,N_4853);
xor U5116 (N_5116,N_4445,N_4813);
nor U5117 (N_5117,N_4838,N_4464);
and U5118 (N_5118,N_4778,N_4877);
or U5119 (N_5119,N_4261,N_4764);
or U5120 (N_5120,N_4961,N_4918);
or U5121 (N_5121,N_4041,N_4897);
and U5122 (N_5122,N_4036,N_4357);
nand U5123 (N_5123,N_4269,N_4063);
or U5124 (N_5124,N_4372,N_4249);
xnor U5125 (N_5125,N_4772,N_4232);
nor U5126 (N_5126,N_4422,N_4547);
nand U5127 (N_5127,N_4836,N_4847);
nand U5128 (N_5128,N_4136,N_4226);
nor U5129 (N_5129,N_4010,N_4963);
nor U5130 (N_5130,N_4597,N_4892);
nand U5131 (N_5131,N_4899,N_4411);
and U5132 (N_5132,N_4723,N_4760);
nand U5133 (N_5133,N_4048,N_4396);
and U5134 (N_5134,N_4885,N_4005);
nor U5135 (N_5135,N_4766,N_4101);
nor U5136 (N_5136,N_4197,N_4423);
nand U5137 (N_5137,N_4333,N_4941);
or U5138 (N_5138,N_4478,N_4135);
and U5139 (N_5139,N_4770,N_4612);
xnor U5140 (N_5140,N_4912,N_4730);
xor U5141 (N_5141,N_4832,N_4904);
xnor U5142 (N_5142,N_4526,N_4011);
xnor U5143 (N_5143,N_4096,N_4677);
and U5144 (N_5144,N_4481,N_4296);
nand U5145 (N_5145,N_4319,N_4754);
nand U5146 (N_5146,N_4273,N_4751);
or U5147 (N_5147,N_4064,N_4082);
nor U5148 (N_5148,N_4338,N_4093);
nor U5149 (N_5149,N_4682,N_4003);
xor U5150 (N_5150,N_4475,N_4743);
nor U5151 (N_5151,N_4528,N_4044);
nand U5152 (N_5152,N_4831,N_4659);
and U5153 (N_5153,N_4848,N_4609);
nor U5154 (N_5154,N_4158,N_4480);
and U5155 (N_5155,N_4692,N_4780);
nor U5156 (N_5156,N_4825,N_4178);
xor U5157 (N_5157,N_4204,N_4024);
or U5158 (N_5158,N_4184,N_4876);
and U5159 (N_5159,N_4630,N_4324);
nor U5160 (N_5160,N_4342,N_4595);
nand U5161 (N_5161,N_4788,N_4805);
or U5162 (N_5162,N_4246,N_4894);
or U5163 (N_5163,N_4488,N_4130);
xor U5164 (N_5164,N_4546,N_4686);
and U5165 (N_5165,N_4893,N_4017);
nand U5166 (N_5166,N_4919,N_4954);
nand U5167 (N_5167,N_4425,N_4066);
or U5168 (N_5168,N_4936,N_4591);
nor U5169 (N_5169,N_4553,N_4823);
nand U5170 (N_5170,N_4951,N_4603);
nand U5171 (N_5171,N_4602,N_4556);
nand U5172 (N_5172,N_4931,N_4175);
nand U5173 (N_5173,N_4995,N_4207);
nor U5174 (N_5174,N_4588,N_4449);
nand U5175 (N_5175,N_4161,N_4453);
or U5176 (N_5176,N_4721,N_4900);
xnor U5177 (N_5177,N_4646,N_4532);
nor U5178 (N_5178,N_4765,N_4229);
nor U5179 (N_5179,N_4829,N_4085);
nand U5180 (N_5180,N_4213,N_4845);
or U5181 (N_5181,N_4781,N_4196);
or U5182 (N_5182,N_4504,N_4255);
or U5183 (N_5183,N_4474,N_4914);
or U5184 (N_5184,N_4262,N_4337);
xnor U5185 (N_5185,N_4070,N_4982);
or U5186 (N_5186,N_4758,N_4260);
nor U5187 (N_5187,N_4058,N_4994);
nand U5188 (N_5188,N_4015,N_4125);
nand U5189 (N_5189,N_4392,N_4067);
xor U5190 (N_5190,N_4511,N_4810);
nor U5191 (N_5191,N_4611,N_4402);
nor U5192 (N_5192,N_4830,N_4133);
nand U5193 (N_5193,N_4451,N_4227);
and U5194 (N_5194,N_4809,N_4545);
or U5195 (N_5195,N_4469,N_4625);
or U5196 (N_5196,N_4022,N_4250);
and U5197 (N_5197,N_4276,N_4124);
or U5198 (N_5198,N_4363,N_4567);
or U5199 (N_5199,N_4183,N_4608);
nor U5200 (N_5200,N_4054,N_4079);
nor U5201 (N_5201,N_4432,N_4903);
nand U5202 (N_5202,N_4346,N_4747);
nor U5203 (N_5203,N_4950,N_4944);
and U5204 (N_5204,N_4517,N_4939);
nand U5205 (N_5205,N_4574,N_4962);
nand U5206 (N_5206,N_4115,N_4585);
and U5207 (N_5207,N_4691,N_4515);
or U5208 (N_5208,N_4379,N_4840);
nand U5209 (N_5209,N_4390,N_4050);
nor U5210 (N_5210,N_4051,N_4420);
xnor U5211 (N_5211,N_4607,N_4956);
nor U5212 (N_5212,N_4025,N_4381);
and U5213 (N_5213,N_4142,N_4155);
or U5214 (N_5214,N_4398,N_4745);
xor U5215 (N_5215,N_4586,N_4973);
nor U5216 (N_5216,N_4002,N_4855);
xnor U5217 (N_5217,N_4113,N_4393);
xor U5218 (N_5218,N_4859,N_4593);
xor U5219 (N_5219,N_4858,N_4494);
or U5220 (N_5220,N_4653,N_4683);
xnor U5221 (N_5221,N_4414,N_4685);
nor U5222 (N_5222,N_4167,N_4305);
or U5223 (N_5223,N_4126,N_4159);
nand U5224 (N_5224,N_4047,N_4933);
nand U5225 (N_5225,N_4857,N_4929);
and U5226 (N_5226,N_4867,N_4938);
xor U5227 (N_5227,N_4075,N_4222);
and U5228 (N_5228,N_4046,N_4708);
or U5229 (N_5229,N_4525,N_4215);
nor U5230 (N_5230,N_4031,N_4092);
and U5231 (N_5231,N_4666,N_4012);
nand U5232 (N_5232,N_4698,N_4644);
or U5233 (N_5233,N_4531,N_4176);
or U5234 (N_5234,N_4740,N_4507);
or U5235 (N_5235,N_4986,N_4582);
and U5236 (N_5236,N_4975,N_4820);
xnor U5237 (N_5237,N_4689,N_4742);
nand U5238 (N_5238,N_4669,N_4295);
or U5239 (N_5239,N_4629,N_4584);
xnor U5240 (N_5240,N_4105,N_4088);
nor U5241 (N_5241,N_4496,N_4930);
nor U5242 (N_5242,N_4339,N_4601);
xnor U5243 (N_5243,N_4146,N_4416);
nor U5244 (N_5244,N_4103,N_4779);
and U5245 (N_5245,N_4712,N_4871);
nand U5246 (N_5246,N_4440,N_4173);
nor U5247 (N_5247,N_4972,N_4293);
nand U5248 (N_5248,N_4552,N_4157);
or U5249 (N_5249,N_4756,N_4127);
xor U5250 (N_5250,N_4856,N_4925);
or U5251 (N_5251,N_4680,N_4039);
and U5252 (N_5252,N_4412,N_4299);
or U5253 (N_5253,N_4144,N_4106);
xnor U5254 (N_5254,N_4658,N_4713);
xnor U5255 (N_5255,N_4886,N_4100);
and U5256 (N_5256,N_4038,N_4789);
nand U5257 (N_5257,N_4536,N_4703);
nand U5258 (N_5258,N_4664,N_4863);
and U5259 (N_5259,N_4564,N_4834);
and U5260 (N_5260,N_4128,N_4699);
and U5261 (N_5261,N_4444,N_4405);
nor U5262 (N_5262,N_4345,N_4470);
nor U5263 (N_5263,N_4649,N_4524);
xnor U5264 (N_5264,N_4978,N_4367);
and U5265 (N_5265,N_4350,N_4921);
nor U5266 (N_5266,N_4138,N_4519);
xnor U5267 (N_5267,N_4502,N_4221);
nand U5268 (N_5268,N_4244,N_4259);
nor U5269 (N_5269,N_4053,N_4240);
and U5270 (N_5270,N_4580,N_4200);
nand U5271 (N_5271,N_4477,N_4181);
nand U5272 (N_5272,N_4225,N_4675);
nand U5273 (N_5273,N_4217,N_4997);
nand U5274 (N_5274,N_4371,N_4083);
or U5275 (N_5275,N_4726,N_4798);
or U5276 (N_5276,N_4418,N_4578);
and U5277 (N_5277,N_4272,N_4330);
or U5278 (N_5278,N_4739,N_4843);
or U5279 (N_5279,N_4817,N_4001);
or U5280 (N_5280,N_4231,N_4169);
nand U5281 (N_5281,N_4325,N_4235);
nor U5282 (N_5282,N_4627,N_4851);
nor U5283 (N_5283,N_4833,N_4503);
xor U5284 (N_5284,N_4694,N_4028);
or U5285 (N_5285,N_4761,N_4660);
xnor U5286 (N_5286,N_4097,N_4527);
xnor U5287 (N_5287,N_4624,N_4465);
nor U5288 (N_5288,N_4724,N_4619);
or U5289 (N_5289,N_4121,N_4657);
nor U5290 (N_5290,N_4874,N_4343);
nand U5291 (N_5291,N_4369,N_4673);
nand U5292 (N_5292,N_4777,N_4186);
and U5293 (N_5293,N_4577,N_4302);
and U5294 (N_5294,N_4785,N_4771);
or U5295 (N_5295,N_4300,N_4134);
and U5296 (N_5296,N_4201,N_4674);
or U5297 (N_5297,N_4562,N_4852);
or U5298 (N_5298,N_4387,N_4008);
or U5299 (N_5299,N_4275,N_4632);
xnor U5300 (N_5300,N_4029,N_4436);
nor U5301 (N_5301,N_4192,N_4095);
or U5302 (N_5302,N_4073,N_4696);
xnor U5303 (N_5303,N_4501,N_4665);
or U5304 (N_5304,N_4570,N_4631);
and U5305 (N_5305,N_4034,N_4212);
or U5306 (N_5306,N_4410,N_4098);
nand U5307 (N_5307,N_4145,N_4568);
or U5308 (N_5308,N_4592,N_4397);
and U5309 (N_5309,N_4266,N_4247);
and U5310 (N_5310,N_4483,N_4122);
and U5311 (N_5311,N_4792,N_4306);
and U5312 (N_5312,N_4216,N_4676);
and U5313 (N_5313,N_4991,N_4541);
xor U5314 (N_5314,N_4004,N_4864);
and U5315 (N_5315,N_4278,N_4123);
or U5316 (N_5316,N_4373,N_4170);
nor U5317 (N_5317,N_4977,N_4006);
nor U5318 (N_5318,N_4151,N_4311);
xor U5319 (N_5319,N_4055,N_4808);
or U5320 (N_5320,N_4252,N_4370);
xor U5321 (N_5321,N_4180,N_4647);
nor U5322 (N_5322,N_4710,N_4378);
and U5323 (N_5323,N_4165,N_4239);
nand U5324 (N_5324,N_4473,N_4642);
xnor U5325 (N_5325,N_4439,N_4875);
and U5326 (N_5326,N_4237,N_4460);
and U5327 (N_5327,N_4814,N_4981);
nand U5328 (N_5328,N_4932,N_4783);
nor U5329 (N_5329,N_4934,N_4984);
nor U5330 (N_5330,N_4952,N_4303);
nor U5331 (N_5331,N_4862,N_4433);
or U5332 (N_5332,N_4336,N_4799);
xor U5333 (N_5333,N_4313,N_4104);
nor U5334 (N_5334,N_4023,N_4806);
nand U5335 (N_5335,N_4516,N_4059);
nor U5336 (N_5336,N_4803,N_4604);
or U5337 (N_5337,N_4804,N_4056);
nor U5338 (N_5338,N_4368,N_4152);
or U5339 (N_5339,N_4948,N_4538);
nand U5340 (N_5340,N_4711,N_4132);
and U5341 (N_5341,N_4413,N_4060);
nor U5342 (N_5342,N_4966,N_4842);
xnor U5343 (N_5343,N_4030,N_4238);
nand U5344 (N_5344,N_4137,N_4828);
nor U5345 (N_5345,N_4195,N_4522);
nand U5346 (N_5346,N_4162,N_4131);
and U5347 (N_5347,N_4282,N_4328);
nand U5348 (N_5348,N_4360,N_4596);
xor U5349 (N_5349,N_4076,N_4140);
and U5350 (N_5350,N_4652,N_4141);
nor U5351 (N_5351,N_4731,N_4815);
nand U5352 (N_5352,N_4935,N_4637);
and U5353 (N_5353,N_4094,N_4009);
or U5354 (N_5354,N_4945,N_4826);
or U5355 (N_5355,N_4409,N_4873);
nand U5356 (N_5356,N_4476,N_4579);
or U5357 (N_5357,N_4529,N_4884);
or U5358 (N_5358,N_4421,N_4072);
nor U5359 (N_5359,N_4571,N_4746);
and U5360 (N_5360,N_4462,N_4205);
or U5361 (N_5361,N_4513,N_4163);
nand U5362 (N_5362,N_4878,N_4895);
nor U5363 (N_5363,N_4812,N_4865);
and U5364 (N_5364,N_4351,N_4987);
xnor U5365 (N_5365,N_4572,N_4540);
and U5366 (N_5366,N_4356,N_4909);
nor U5367 (N_5367,N_4043,N_4443);
xor U5368 (N_5368,N_4318,N_4074);
nand U5369 (N_5369,N_4880,N_4883);
and U5370 (N_5370,N_4718,N_4385);
and U5371 (N_5371,N_4748,N_4458);
and U5372 (N_5372,N_4116,N_4294);
and U5373 (N_5373,N_4291,N_4911);
or U5374 (N_5374,N_4290,N_4265);
nand U5375 (N_5375,N_4861,N_4650);
or U5376 (N_5376,N_4622,N_4377);
and U5377 (N_5377,N_4084,N_4320);
or U5378 (N_5378,N_4118,N_4019);
and U5379 (N_5379,N_4499,N_4924);
or U5380 (N_5380,N_4220,N_4424);
nor U5381 (N_5381,N_4243,N_4080);
xor U5382 (N_5382,N_4129,N_4725);
nor U5383 (N_5383,N_4329,N_4287);
nand U5384 (N_5384,N_4099,N_4189);
xnor U5385 (N_5385,N_4309,N_4208);
nand U5386 (N_5386,N_4655,N_4500);
or U5387 (N_5387,N_4087,N_4316);
or U5388 (N_5388,N_4614,N_4236);
or U5389 (N_5389,N_4732,N_4958);
nor U5390 (N_5390,N_4156,N_4108);
nor U5391 (N_5391,N_4391,N_4061);
xnor U5392 (N_5392,N_4583,N_4497);
xnor U5393 (N_5393,N_4733,N_4827);
and U5394 (N_5394,N_4388,N_4993);
or U5395 (N_5395,N_4461,N_4248);
and U5396 (N_5396,N_4251,N_4040);
nand U5397 (N_5397,N_4362,N_4331);
and U5398 (N_5398,N_4898,N_4768);
and U5399 (N_5399,N_4551,N_4946);
and U5400 (N_5400,N_4870,N_4408);
and U5401 (N_5401,N_4965,N_4920);
nor U5402 (N_5402,N_4942,N_4634);
xor U5403 (N_5403,N_4086,N_4032);
nor U5404 (N_5404,N_4253,N_4559);
xor U5405 (N_5405,N_4512,N_4364);
or U5406 (N_5406,N_4510,N_4800);
nor U5407 (N_5407,N_4467,N_4312);
nor U5408 (N_5408,N_4636,N_4139);
nand U5409 (N_5409,N_4594,N_4902);
xor U5410 (N_5410,N_4613,N_4575);
or U5411 (N_5411,N_4555,N_4491);
or U5412 (N_5412,N_4693,N_4821);
xnor U5413 (N_5413,N_4426,N_4089);
nor U5414 (N_5414,N_4120,N_4796);
and U5415 (N_5415,N_4620,N_4976);
nor U5416 (N_5416,N_4762,N_4257);
xor U5417 (N_5417,N_4633,N_4281);
xor U5418 (N_5418,N_4543,N_4486);
and U5419 (N_5419,N_4441,N_4233);
xor U5420 (N_5420,N_4153,N_4908);
xnor U5421 (N_5421,N_4335,N_4890);
xnor U5422 (N_5422,N_4709,N_4431);
nand U5423 (N_5423,N_4561,N_4168);
or U5424 (N_5424,N_4077,N_4974);
or U5425 (N_5425,N_4707,N_4109);
nand U5426 (N_5426,N_4214,N_4999);
or U5427 (N_5427,N_4971,N_4891);
nand U5428 (N_5428,N_4321,N_4277);
xnor U5429 (N_5429,N_4807,N_4430);
or U5430 (N_5430,N_4289,N_4869);
and U5431 (N_5431,N_4479,N_4062);
nor U5432 (N_5432,N_4907,N_4509);
xor U5433 (N_5433,N_4506,N_4267);
xnor U5434 (N_5434,N_4033,N_4881);
and U5435 (N_5435,N_4749,N_4071);
xnor U5436 (N_5436,N_4365,N_4988);
nor U5437 (N_5437,N_4520,N_4211);
nand U5438 (N_5438,N_4722,N_4518);
xor U5439 (N_5439,N_4701,N_4744);
nand U5440 (N_5440,N_4174,N_4487);
xnor U5441 (N_5441,N_4000,N_4308);
nand U5442 (N_5442,N_4353,N_4791);
or U5443 (N_5443,N_4589,N_4376);
nor U5444 (N_5444,N_4697,N_4590);
nand U5445 (N_5445,N_4428,N_4172);
or U5446 (N_5446,N_4767,N_4322);
or U5447 (N_5447,N_4288,N_4199);
or U5448 (N_5448,N_4505,N_4407);
or U5449 (N_5449,N_4916,N_4794);
nor U5450 (N_5450,N_4795,N_4406);
nor U5451 (N_5451,N_4091,N_4661);
nor U5452 (N_5452,N_4906,N_4656);
or U5453 (N_5453,N_4297,N_4979);
xnor U5454 (N_5454,N_4484,N_4967);
xnor U5455 (N_5455,N_4242,N_4389);
nand U5456 (N_5456,N_4112,N_4573);
xnor U5457 (N_5457,N_4752,N_4671);
nand U5458 (N_5458,N_4254,N_4610);
and U5459 (N_5459,N_4648,N_4198);
and U5460 (N_5460,N_4782,N_4190);
nand U5461 (N_5461,N_4905,N_4651);
and U5462 (N_5462,N_4018,N_4352);
xor U5463 (N_5463,N_4940,N_4888);
or U5464 (N_5464,N_4107,N_4533);
and U5465 (N_5465,N_4090,N_4539);
nor U5466 (N_5466,N_4635,N_4117);
and U5467 (N_5467,N_4493,N_4846);
or U5468 (N_5468,N_4037,N_4206);
and U5469 (N_5469,N_4304,N_4027);
xnor U5470 (N_5470,N_4014,N_4996);
nor U5471 (N_5471,N_4937,N_4358);
xor U5472 (N_5472,N_4110,N_4452);
or U5473 (N_5473,N_4735,N_4459);
xnor U5474 (N_5474,N_4382,N_4753);
or U5475 (N_5475,N_4187,N_4057);
nand U5476 (N_5476,N_4949,N_4638);
xnor U5477 (N_5477,N_4534,N_4399);
and U5478 (N_5478,N_4148,N_4998);
nand U5479 (N_5479,N_4218,N_4801);
or U5480 (N_5480,N_4442,N_4550);
nand U5481 (N_5481,N_4882,N_4569);
xor U5482 (N_5482,N_4340,N_4943);
nand U5483 (N_5483,N_4587,N_4348);
or U5484 (N_5484,N_4349,N_4341);
nor U5485 (N_5485,N_4463,N_4111);
xor U5486 (N_5486,N_4896,N_4850);
and U5487 (N_5487,N_4643,N_4334);
nand U5488 (N_5488,N_4448,N_4450);
and U5489 (N_5489,N_4383,N_4427);
xnor U5490 (N_5490,N_4990,N_4959);
xor U5491 (N_5491,N_4913,N_4645);
nor U5492 (N_5492,N_4203,N_4824);
xnor U5493 (N_5493,N_4549,N_4344);
or U5494 (N_5494,N_4326,N_4234);
xnor U5495 (N_5495,N_4769,N_4323);
and U5496 (N_5496,N_4968,N_4872);
or U5497 (N_5497,N_4776,N_4926);
xnor U5498 (N_5498,N_4271,N_4185);
xor U5499 (N_5499,N_4191,N_4787);
and U5500 (N_5500,N_4047,N_4953);
nand U5501 (N_5501,N_4885,N_4006);
nand U5502 (N_5502,N_4570,N_4618);
and U5503 (N_5503,N_4709,N_4395);
nand U5504 (N_5504,N_4196,N_4788);
nor U5505 (N_5505,N_4863,N_4994);
nor U5506 (N_5506,N_4343,N_4499);
xnor U5507 (N_5507,N_4574,N_4156);
nand U5508 (N_5508,N_4724,N_4078);
nand U5509 (N_5509,N_4702,N_4482);
xnor U5510 (N_5510,N_4798,N_4267);
nor U5511 (N_5511,N_4732,N_4011);
nor U5512 (N_5512,N_4450,N_4561);
nor U5513 (N_5513,N_4427,N_4944);
and U5514 (N_5514,N_4326,N_4619);
and U5515 (N_5515,N_4928,N_4945);
nor U5516 (N_5516,N_4676,N_4816);
nand U5517 (N_5517,N_4194,N_4147);
nor U5518 (N_5518,N_4115,N_4217);
and U5519 (N_5519,N_4193,N_4269);
and U5520 (N_5520,N_4161,N_4368);
xnor U5521 (N_5521,N_4508,N_4782);
xor U5522 (N_5522,N_4676,N_4368);
and U5523 (N_5523,N_4271,N_4234);
or U5524 (N_5524,N_4141,N_4519);
xnor U5525 (N_5525,N_4040,N_4408);
and U5526 (N_5526,N_4482,N_4822);
and U5527 (N_5527,N_4312,N_4377);
xnor U5528 (N_5528,N_4760,N_4188);
or U5529 (N_5529,N_4009,N_4179);
or U5530 (N_5530,N_4167,N_4691);
nand U5531 (N_5531,N_4592,N_4434);
nand U5532 (N_5532,N_4491,N_4189);
xnor U5533 (N_5533,N_4547,N_4697);
xor U5534 (N_5534,N_4673,N_4852);
xnor U5535 (N_5535,N_4853,N_4268);
nand U5536 (N_5536,N_4917,N_4875);
nand U5537 (N_5537,N_4351,N_4431);
xor U5538 (N_5538,N_4099,N_4386);
nor U5539 (N_5539,N_4822,N_4929);
and U5540 (N_5540,N_4061,N_4938);
nor U5541 (N_5541,N_4827,N_4413);
xnor U5542 (N_5542,N_4649,N_4503);
nor U5543 (N_5543,N_4702,N_4520);
nor U5544 (N_5544,N_4258,N_4664);
nor U5545 (N_5545,N_4585,N_4086);
or U5546 (N_5546,N_4522,N_4482);
nand U5547 (N_5547,N_4741,N_4585);
and U5548 (N_5548,N_4975,N_4705);
and U5549 (N_5549,N_4062,N_4680);
and U5550 (N_5550,N_4767,N_4908);
xnor U5551 (N_5551,N_4169,N_4506);
or U5552 (N_5552,N_4593,N_4773);
xor U5553 (N_5553,N_4513,N_4784);
and U5554 (N_5554,N_4078,N_4128);
or U5555 (N_5555,N_4677,N_4152);
and U5556 (N_5556,N_4049,N_4296);
or U5557 (N_5557,N_4820,N_4180);
nor U5558 (N_5558,N_4699,N_4484);
and U5559 (N_5559,N_4413,N_4233);
xnor U5560 (N_5560,N_4334,N_4853);
xor U5561 (N_5561,N_4154,N_4927);
nand U5562 (N_5562,N_4203,N_4672);
or U5563 (N_5563,N_4867,N_4889);
xor U5564 (N_5564,N_4706,N_4272);
nor U5565 (N_5565,N_4786,N_4005);
xor U5566 (N_5566,N_4386,N_4598);
nand U5567 (N_5567,N_4464,N_4611);
and U5568 (N_5568,N_4219,N_4908);
or U5569 (N_5569,N_4792,N_4990);
and U5570 (N_5570,N_4382,N_4087);
xor U5571 (N_5571,N_4442,N_4759);
nor U5572 (N_5572,N_4850,N_4948);
and U5573 (N_5573,N_4099,N_4098);
nor U5574 (N_5574,N_4985,N_4670);
nand U5575 (N_5575,N_4784,N_4071);
nor U5576 (N_5576,N_4414,N_4935);
and U5577 (N_5577,N_4544,N_4228);
and U5578 (N_5578,N_4116,N_4796);
nand U5579 (N_5579,N_4938,N_4041);
xnor U5580 (N_5580,N_4115,N_4312);
nor U5581 (N_5581,N_4715,N_4052);
and U5582 (N_5582,N_4767,N_4696);
or U5583 (N_5583,N_4623,N_4675);
and U5584 (N_5584,N_4235,N_4575);
nor U5585 (N_5585,N_4104,N_4663);
and U5586 (N_5586,N_4313,N_4422);
or U5587 (N_5587,N_4840,N_4489);
nor U5588 (N_5588,N_4099,N_4371);
nand U5589 (N_5589,N_4165,N_4454);
nand U5590 (N_5590,N_4398,N_4090);
nand U5591 (N_5591,N_4834,N_4989);
nor U5592 (N_5592,N_4742,N_4290);
nor U5593 (N_5593,N_4460,N_4034);
nor U5594 (N_5594,N_4305,N_4209);
or U5595 (N_5595,N_4924,N_4349);
and U5596 (N_5596,N_4897,N_4277);
xor U5597 (N_5597,N_4620,N_4349);
nor U5598 (N_5598,N_4114,N_4085);
or U5599 (N_5599,N_4708,N_4143);
nand U5600 (N_5600,N_4686,N_4259);
xnor U5601 (N_5601,N_4699,N_4379);
and U5602 (N_5602,N_4303,N_4585);
nand U5603 (N_5603,N_4370,N_4580);
nor U5604 (N_5604,N_4428,N_4967);
xor U5605 (N_5605,N_4000,N_4081);
nor U5606 (N_5606,N_4154,N_4626);
or U5607 (N_5607,N_4065,N_4196);
nand U5608 (N_5608,N_4694,N_4434);
nand U5609 (N_5609,N_4820,N_4863);
and U5610 (N_5610,N_4420,N_4247);
xor U5611 (N_5611,N_4452,N_4265);
nand U5612 (N_5612,N_4289,N_4770);
and U5613 (N_5613,N_4325,N_4987);
nand U5614 (N_5614,N_4948,N_4692);
nor U5615 (N_5615,N_4115,N_4055);
nand U5616 (N_5616,N_4162,N_4126);
nand U5617 (N_5617,N_4574,N_4421);
nor U5618 (N_5618,N_4223,N_4333);
or U5619 (N_5619,N_4617,N_4888);
and U5620 (N_5620,N_4935,N_4631);
and U5621 (N_5621,N_4008,N_4949);
xnor U5622 (N_5622,N_4192,N_4069);
nand U5623 (N_5623,N_4722,N_4571);
nor U5624 (N_5624,N_4935,N_4733);
nand U5625 (N_5625,N_4415,N_4815);
and U5626 (N_5626,N_4022,N_4564);
or U5627 (N_5627,N_4165,N_4829);
nand U5628 (N_5628,N_4053,N_4500);
xnor U5629 (N_5629,N_4272,N_4413);
and U5630 (N_5630,N_4431,N_4133);
xnor U5631 (N_5631,N_4582,N_4987);
nand U5632 (N_5632,N_4549,N_4188);
xor U5633 (N_5633,N_4844,N_4750);
nand U5634 (N_5634,N_4722,N_4888);
xor U5635 (N_5635,N_4911,N_4695);
nand U5636 (N_5636,N_4724,N_4035);
or U5637 (N_5637,N_4460,N_4028);
or U5638 (N_5638,N_4332,N_4838);
nor U5639 (N_5639,N_4968,N_4306);
xnor U5640 (N_5640,N_4917,N_4688);
nor U5641 (N_5641,N_4036,N_4923);
or U5642 (N_5642,N_4217,N_4370);
nand U5643 (N_5643,N_4120,N_4813);
nor U5644 (N_5644,N_4376,N_4485);
xnor U5645 (N_5645,N_4836,N_4468);
and U5646 (N_5646,N_4343,N_4816);
xnor U5647 (N_5647,N_4485,N_4850);
nand U5648 (N_5648,N_4673,N_4051);
nor U5649 (N_5649,N_4954,N_4785);
nand U5650 (N_5650,N_4915,N_4799);
nor U5651 (N_5651,N_4412,N_4392);
xor U5652 (N_5652,N_4441,N_4654);
nand U5653 (N_5653,N_4041,N_4676);
and U5654 (N_5654,N_4356,N_4987);
or U5655 (N_5655,N_4770,N_4673);
and U5656 (N_5656,N_4320,N_4770);
nor U5657 (N_5657,N_4741,N_4405);
xnor U5658 (N_5658,N_4330,N_4607);
nand U5659 (N_5659,N_4367,N_4550);
xnor U5660 (N_5660,N_4138,N_4832);
xor U5661 (N_5661,N_4541,N_4004);
nor U5662 (N_5662,N_4947,N_4557);
nand U5663 (N_5663,N_4055,N_4908);
or U5664 (N_5664,N_4056,N_4608);
xnor U5665 (N_5665,N_4102,N_4696);
nand U5666 (N_5666,N_4895,N_4320);
and U5667 (N_5667,N_4089,N_4236);
xnor U5668 (N_5668,N_4159,N_4052);
xnor U5669 (N_5669,N_4552,N_4207);
or U5670 (N_5670,N_4931,N_4988);
nor U5671 (N_5671,N_4421,N_4954);
nor U5672 (N_5672,N_4085,N_4191);
nand U5673 (N_5673,N_4365,N_4863);
and U5674 (N_5674,N_4679,N_4292);
nor U5675 (N_5675,N_4007,N_4650);
and U5676 (N_5676,N_4772,N_4713);
or U5677 (N_5677,N_4536,N_4446);
xnor U5678 (N_5678,N_4070,N_4728);
nand U5679 (N_5679,N_4201,N_4490);
and U5680 (N_5680,N_4510,N_4977);
and U5681 (N_5681,N_4523,N_4090);
nor U5682 (N_5682,N_4492,N_4354);
nand U5683 (N_5683,N_4078,N_4248);
nand U5684 (N_5684,N_4107,N_4302);
nand U5685 (N_5685,N_4802,N_4594);
and U5686 (N_5686,N_4118,N_4660);
and U5687 (N_5687,N_4332,N_4951);
xnor U5688 (N_5688,N_4384,N_4167);
or U5689 (N_5689,N_4149,N_4546);
nand U5690 (N_5690,N_4113,N_4037);
nor U5691 (N_5691,N_4734,N_4039);
nor U5692 (N_5692,N_4291,N_4948);
nand U5693 (N_5693,N_4978,N_4753);
nand U5694 (N_5694,N_4213,N_4630);
xnor U5695 (N_5695,N_4299,N_4449);
nor U5696 (N_5696,N_4105,N_4389);
and U5697 (N_5697,N_4810,N_4858);
and U5698 (N_5698,N_4622,N_4944);
nand U5699 (N_5699,N_4420,N_4153);
xnor U5700 (N_5700,N_4587,N_4527);
xnor U5701 (N_5701,N_4293,N_4335);
or U5702 (N_5702,N_4943,N_4142);
nor U5703 (N_5703,N_4494,N_4384);
or U5704 (N_5704,N_4515,N_4912);
or U5705 (N_5705,N_4377,N_4883);
xor U5706 (N_5706,N_4418,N_4514);
xor U5707 (N_5707,N_4505,N_4706);
or U5708 (N_5708,N_4546,N_4380);
and U5709 (N_5709,N_4761,N_4428);
nand U5710 (N_5710,N_4063,N_4109);
or U5711 (N_5711,N_4166,N_4286);
xor U5712 (N_5712,N_4899,N_4554);
and U5713 (N_5713,N_4549,N_4021);
nand U5714 (N_5714,N_4764,N_4613);
and U5715 (N_5715,N_4936,N_4610);
nand U5716 (N_5716,N_4077,N_4096);
or U5717 (N_5717,N_4894,N_4663);
nor U5718 (N_5718,N_4544,N_4908);
or U5719 (N_5719,N_4462,N_4143);
nor U5720 (N_5720,N_4332,N_4912);
or U5721 (N_5721,N_4589,N_4494);
or U5722 (N_5722,N_4779,N_4405);
and U5723 (N_5723,N_4095,N_4986);
nand U5724 (N_5724,N_4828,N_4151);
nor U5725 (N_5725,N_4136,N_4034);
and U5726 (N_5726,N_4216,N_4733);
nand U5727 (N_5727,N_4562,N_4120);
or U5728 (N_5728,N_4252,N_4055);
and U5729 (N_5729,N_4646,N_4196);
nor U5730 (N_5730,N_4908,N_4793);
and U5731 (N_5731,N_4736,N_4227);
or U5732 (N_5732,N_4371,N_4273);
xor U5733 (N_5733,N_4517,N_4720);
xnor U5734 (N_5734,N_4458,N_4871);
or U5735 (N_5735,N_4903,N_4975);
nor U5736 (N_5736,N_4358,N_4091);
nor U5737 (N_5737,N_4858,N_4531);
xnor U5738 (N_5738,N_4797,N_4097);
or U5739 (N_5739,N_4621,N_4207);
nand U5740 (N_5740,N_4832,N_4906);
or U5741 (N_5741,N_4882,N_4186);
nor U5742 (N_5742,N_4513,N_4579);
and U5743 (N_5743,N_4563,N_4657);
xor U5744 (N_5744,N_4602,N_4125);
nor U5745 (N_5745,N_4154,N_4096);
xnor U5746 (N_5746,N_4327,N_4367);
and U5747 (N_5747,N_4546,N_4347);
nor U5748 (N_5748,N_4818,N_4594);
nand U5749 (N_5749,N_4986,N_4985);
xor U5750 (N_5750,N_4623,N_4726);
nand U5751 (N_5751,N_4519,N_4008);
nor U5752 (N_5752,N_4845,N_4913);
nor U5753 (N_5753,N_4185,N_4539);
or U5754 (N_5754,N_4029,N_4704);
and U5755 (N_5755,N_4440,N_4560);
and U5756 (N_5756,N_4415,N_4723);
nand U5757 (N_5757,N_4296,N_4963);
xor U5758 (N_5758,N_4815,N_4173);
or U5759 (N_5759,N_4243,N_4612);
xnor U5760 (N_5760,N_4824,N_4382);
nor U5761 (N_5761,N_4487,N_4480);
or U5762 (N_5762,N_4422,N_4128);
xnor U5763 (N_5763,N_4440,N_4494);
and U5764 (N_5764,N_4209,N_4275);
or U5765 (N_5765,N_4471,N_4015);
nand U5766 (N_5766,N_4845,N_4899);
nand U5767 (N_5767,N_4277,N_4259);
xnor U5768 (N_5768,N_4971,N_4774);
nor U5769 (N_5769,N_4550,N_4130);
xnor U5770 (N_5770,N_4678,N_4382);
and U5771 (N_5771,N_4228,N_4410);
nor U5772 (N_5772,N_4291,N_4549);
nor U5773 (N_5773,N_4233,N_4731);
xor U5774 (N_5774,N_4174,N_4447);
nand U5775 (N_5775,N_4326,N_4717);
nor U5776 (N_5776,N_4438,N_4566);
nand U5777 (N_5777,N_4831,N_4218);
nand U5778 (N_5778,N_4260,N_4929);
and U5779 (N_5779,N_4880,N_4189);
and U5780 (N_5780,N_4477,N_4888);
nand U5781 (N_5781,N_4328,N_4692);
and U5782 (N_5782,N_4153,N_4890);
and U5783 (N_5783,N_4752,N_4350);
or U5784 (N_5784,N_4384,N_4844);
nor U5785 (N_5785,N_4344,N_4407);
or U5786 (N_5786,N_4537,N_4704);
or U5787 (N_5787,N_4213,N_4664);
or U5788 (N_5788,N_4277,N_4769);
nand U5789 (N_5789,N_4892,N_4420);
nand U5790 (N_5790,N_4387,N_4541);
or U5791 (N_5791,N_4733,N_4649);
nor U5792 (N_5792,N_4650,N_4137);
and U5793 (N_5793,N_4024,N_4397);
nor U5794 (N_5794,N_4179,N_4883);
nor U5795 (N_5795,N_4597,N_4249);
nor U5796 (N_5796,N_4963,N_4086);
and U5797 (N_5797,N_4952,N_4880);
or U5798 (N_5798,N_4907,N_4609);
and U5799 (N_5799,N_4263,N_4760);
nor U5800 (N_5800,N_4751,N_4888);
xor U5801 (N_5801,N_4749,N_4295);
xor U5802 (N_5802,N_4006,N_4546);
xnor U5803 (N_5803,N_4691,N_4198);
or U5804 (N_5804,N_4646,N_4459);
and U5805 (N_5805,N_4553,N_4234);
nor U5806 (N_5806,N_4043,N_4882);
nor U5807 (N_5807,N_4596,N_4641);
nor U5808 (N_5808,N_4576,N_4662);
and U5809 (N_5809,N_4651,N_4902);
nand U5810 (N_5810,N_4375,N_4115);
or U5811 (N_5811,N_4668,N_4883);
xor U5812 (N_5812,N_4631,N_4844);
xnor U5813 (N_5813,N_4711,N_4779);
nor U5814 (N_5814,N_4228,N_4620);
nor U5815 (N_5815,N_4061,N_4335);
nand U5816 (N_5816,N_4682,N_4480);
nor U5817 (N_5817,N_4539,N_4380);
nand U5818 (N_5818,N_4701,N_4976);
and U5819 (N_5819,N_4147,N_4626);
nor U5820 (N_5820,N_4875,N_4894);
xnor U5821 (N_5821,N_4499,N_4494);
and U5822 (N_5822,N_4499,N_4443);
nor U5823 (N_5823,N_4873,N_4157);
or U5824 (N_5824,N_4104,N_4815);
nand U5825 (N_5825,N_4508,N_4017);
xor U5826 (N_5826,N_4985,N_4621);
and U5827 (N_5827,N_4036,N_4762);
nor U5828 (N_5828,N_4890,N_4964);
and U5829 (N_5829,N_4541,N_4975);
xor U5830 (N_5830,N_4642,N_4827);
and U5831 (N_5831,N_4584,N_4437);
nor U5832 (N_5832,N_4001,N_4458);
nand U5833 (N_5833,N_4030,N_4425);
nand U5834 (N_5834,N_4854,N_4383);
xnor U5835 (N_5835,N_4763,N_4640);
and U5836 (N_5836,N_4960,N_4145);
nand U5837 (N_5837,N_4659,N_4081);
nor U5838 (N_5838,N_4234,N_4661);
nand U5839 (N_5839,N_4532,N_4347);
nor U5840 (N_5840,N_4691,N_4665);
and U5841 (N_5841,N_4717,N_4125);
nor U5842 (N_5842,N_4855,N_4638);
nand U5843 (N_5843,N_4846,N_4740);
nor U5844 (N_5844,N_4722,N_4982);
nor U5845 (N_5845,N_4939,N_4512);
xor U5846 (N_5846,N_4377,N_4485);
or U5847 (N_5847,N_4601,N_4243);
xor U5848 (N_5848,N_4611,N_4552);
nand U5849 (N_5849,N_4591,N_4573);
nor U5850 (N_5850,N_4525,N_4557);
nor U5851 (N_5851,N_4390,N_4107);
and U5852 (N_5852,N_4270,N_4743);
nand U5853 (N_5853,N_4371,N_4653);
nor U5854 (N_5854,N_4727,N_4492);
xnor U5855 (N_5855,N_4988,N_4839);
nor U5856 (N_5856,N_4122,N_4061);
nor U5857 (N_5857,N_4115,N_4006);
xnor U5858 (N_5858,N_4065,N_4026);
xor U5859 (N_5859,N_4872,N_4415);
nor U5860 (N_5860,N_4340,N_4409);
and U5861 (N_5861,N_4749,N_4292);
and U5862 (N_5862,N_4093,N_4218);
nor U5863 (N_5863,N_4816,N_4230);
or U5864 (N_5864,N_4147,N_4076);
xnor U5865 (N_5865,N_4614,N_4339);
nor U5866 (N_5866,N_4559,N_4891);
xor U5867 (N_5867,N_4473,N_4856);
nand U5868 (N_5868,N_4351,N_4622);
and U5869 (N_5869,N_4490,N_4523);
nor U5870 (N_5870,N_4671,N_4600);
nand U5871 (N_5871,N_4766,N_4262);
nor U5872 (N_5872,N_4539,N_4089);
or U5873 (N_5873,N_4165,N_4727);
or U5874 (N_5874,N_4166,N_4855);
nand U5875 (N_5875,N_4905,N_4165);
or U5876 (N_5876,N_4395,N_4205);
and U5877 (N_5877,N_4359,N_4611);
nand U5878 (N_5878,N_4518,N_4840);
and U5879 (N_5879,N_4562,N_4367);
nor U5880 (N_5880,N_4867,N_4770);
nor U5881 (N_5881,N_4995,N_4933);
and U5882 (N_5882,N_4734,N_4475);
nand U5883 (N_5883,N_4758,N_4125);
nor U5884 (N_5884,N_4724,N_4089);
nand U5885 (N_5885,N_4939,N_4306);
xor U5886 (N_5886,N_4567,N_4082);
nand U5887 (N_5887,N_4948,N_4392);
or U5888 (N_5888,N_4102,N_4336);
nor U5889 (N_5889,N_4486,N_4421);
or U5890 (N_5890,N_4994,N_4383);
or U5891 (N_5891,N_4385,N_4503);
or U5892 (N_5892,N_4561,N_4597);
nand U5893 (N_5893,N_4801,N_4136);
xor U5894 (N_5894,N_4039,N_4024);
nor U5895 (N_5895,N_4908,N_4620);
or U5896 (N_5896,N_4997,N_4135);
nor U5897 (N_5897,N_4835,N_4621);
xnor U5898 (N_5898,N_4327,N_4108);
and U5899 (N_5899,N_4456,N_4242);
or U5900 (N_5900,N_4769,N_4692);
nand U5901 (N_5901,N_4238,N_4770);
and U5902 (N_5902,N_4941,N_4887);
nor U5903 (N_5903,N_4328,N_4494);
xnor U5904 (N_5904,N_4484,N_4286);
or U5905 (N_5905,N_4950,N_4141);
nand U5906 (N_5906,N_4384,N_4309);
xnor U5907 (N_5907,N_4746,N_4036);
and U5908 (N_5908,N_4224,N_4553);
and U5909 (N_5909,N_4812,N_4154);
xnor U5910 (N_5910,N_4752,N_4457);
and U5911 (N_5911,N_4647,N_4760);
or U5912 (N_5912,N_4104,N_4150);
nor U5913 (N_5913,N_4818,N_4550);
and U5914 (N_5914,N_4740,N_4742);
or U5915 (N_5915,N_4445,N_4002);
nand U5916 (N_5916,N_4324,N_4135);
xor U5917 (N_5917,N_4813,N_4442);
nand U5918 (N_5918,N_4167,N_4427);
or U5919 (N_5919,N_4001,N_4480);
xor U5920 (N_5920,N_4340,N_4129);
or U5921 (N_5921,N_4567,N_4176);
nand U5922 (N_5922,N_4643,N_4326);
xor U5923 (N_5923,N_4299,N_4174);
nor U5924 (N_5924,N_4552,N_4687);
or U5925 (N_5925,N_4376,N_4037);
nand U5926 (N_5926,N_4948,N_4085);
nor U5927 (N_5927,N_4260,N_4809);
or U5928 (N_5928,N_4812,N_4226);
nor U5929 (N_5929,N_4017,N_4600);
nor U5930 (N_5930,N_4400,N_4235);
or U5931 (N_5931,N_4472,N_4672);
xor U5932 (N_5932,N_4917,N_4366);
nor U5933 (N_5933,N_4130,N_4128);
and U5934 (N_5934,N_4876,N_4421);
xnor U5935 (N_5935,N_4212,N_4353);
and U5936 (N_5936,N_4059,N_4729);
nand U5937 (N_5937,N_4913,N_4640);
or U5938 (N_5938,N_4153,N_4672);
or U5939 (N_5939,N_4988,N_4965);
nand U5940 (N_5940,N_4535,N_4367);
or U5941 (N_5941,N_4051,N_4906);
and U5942 (N_5942,N_4914,N_4964);
nand U5943 (N_5943,N_4281,N_4885);
nor U5944 (N_5944,N_4067,N_4810);
nor U5945 (N_5945,N_4276,N_4446);
nand U5946 (N_5946,N_4970,N_4056);
and U5947 (N_5947,N_4889,N_4792);
xnor U5948 (N_5948,N_4399,N_4544);
nor U5949 (N_5949,N_4487,N_4974);
xor U5950 (N_5950,N_4295,N_4386);
nand U5951 (N_5951,N_4179,N_4594);
nand U5952 (N_5952,N_4910,N_4208);
nor U5953 (N_5953,N_4992,N_4897);
xnor U5954 (N_5954,N_4404,N_4370);
nor U5955 (N_5955,N_4334,N_4503);
nor U5956 (N_5956,N_4128,N_4302);
nor U5957 (N_5957,N_4207,N_4042);
and U5958 (N_5958,N_4759,N_4183);
nor U5959 (N_5959,N_4442,N_4499);
xor U5960 (N_5960,N_4939,N_4363);
xnor U5961 (N_5961,N_4000,N_4680);
or U5962 (N_5962,N_4797,N_4045);
xor U5963 (N_5963,N_4789,N_4798);
nand U5964 (N_5964,N_4755,N_4990);
xnor U5965 (N_5965,N_4835,N_4209);
nor U5966 (N_5966,N_4607,N_4766);
or U5967 (N_5967,N_4868,N_4614);
or U5968 (N_5968,N_4011,N_4090);
or U5969 (N_5969,N_4644,N_4940);
xnor U5970 (N_5970,N_4197,N_4652);
or U5971 (N_5971,N_4651,N_4176);
or U5972 (N_5972,N_4656,N_4987);
nand U5973 (N_5973,N_4820,N_4378);
xor U5974 (N_5974,N_4173,N_4057);
or U5975 (N_5975,N_4262,N_4653);
xor U5976 (N_5976,N_4234,N_4290);
nor U5977 (N_5977,N_4875,N_4701);
xnor U5978 (N_5978,N_4031,N_4094);
nand U5979 (N_5979,N_4343,N_4222);
nand U5980 (N_5980,N_4212,N_4735);
nand U5981 (N_5981,N_4669,N_4348);
or U5982 (N_5982,N_4370,N_4559);
nand U5983 (N_5983,N_4306,N_4232);
or U5984 (N_5984,N_4697,N_4078);
nor U5985 (N_5985,N_4974,N_4236);
or U5986 (N_5986,N_4470,N_4471);
nor U5987 (N_5987,N_4189,N_4396);
or U5988 (N_5988,N_4721,N_4564);
and U5989 (N_5989,N_4309,N_4847);
and U5990 (N_5990,N_4194,N_4842);
xnor U5991 (N_5991,N_4256,N_4253);
nand U5992 (N_5992,N_4698,N_4078);
nand U5993 (N_5993,N_4859,N_4990);
or U5994 (N_5994,N_4228,N_4682);
or U5995 (N_5995,N_4591,N_4169);
xnor U5996 (N_5996,N_4744,N_4649);
and U5997 (N_5997,N_4396,N_4242);
or U5998 (N_5998,N_4164,N_4222);
or U5999 (N_5999,N_4614,N_4523);
nor U6000 (N_6000,N_5801,N_5598);
nor U6001 (N_6001,N_5919,N_5485);
xnor U6002 (N_6002,N_5241,N_5912);
nor U6003 (N_6003,N_5905,N_5233);
and U6004 (N_6004,N_5833,N_5131);
nor U6005 (N_6005,N_5248,N_5047);
nand U6006 (N_6006,N_5627,N_5298);
nand U6007 (N_6007,N_5489,N_5743);
nand U6008 (N_6008,N_5755,N_5917);
or U6009 (N_6009,N_5266,N_5630);
or U6010 (N_6010,N_5192,N_5349);
nor U6011 (N_6011,N_5484,N_5009);
nor U6012 (N_6012,N_5375,N_5786);
xor U6013 (N_6013,N_5441,N_5898);
xor U6014 (N_6014,N_5623,N_5978);
and U6015 (N_6015,N_5715,N_5215);
xnor U6016 (N_6016,N_5619,N_5190);
xor U6017 (N_6017,N_5799,N_5189);
and U6018 (N_6018,N_5566,N_5274);
xor U6019 (N_6019,N_5038,N_5726);
or U6020 (N_6020,N_5197,N_5153);
xnor U6021 (N_6021,N_5582,N_5121);
and U6022 (N_6022,N_5350,N_5065);
nand U6023 (N_6023,N_5272,N_5909);
nor U6024 (N_6024,N_5175,N_5240);
nand U6025 (N_6025,N_5820,N_5367);
or U6026 (N_6026,N_5525,N_5452);
and U6027 (N_6027,N_5933,N_5147);
nand U6028 (N_6028,N_5053,N_5980);
nand U6029 (N_6029,N_5827,N_5171);
and U6030 (N_6030,N_5507,N_5208);
or U6031 (N_6031,N_5366,N_5376);
or U6032 (N_6032,N_5615,N_5050);
nor U6033 (N_6033,N_5934,N_5889);
xnor U6034 (N_6034,N_5915,N_5168);
or U6035 (N_6035,N_5590,N_5094);
nor U6036 (N_6036,N_5652,N_5579);
or U6037 (N_6037,N_5079,N_5541);
nor U6038 (N_6038,N_5389,N_5112);
or U6039 (N_6039,N_5993,N_5339);
xor U6040 (N_6040,N_5870,N_5026);
nand U6041 (N_6041,N_5460,N_5132);
xnor U6042 (N_6042,N_5767,N_5692);
xor U6043 (N_6043,N_5676,N_5849);
and U6044 (N_6044,N_5105,N_5231);
nand U6045 (N_6045,N_5989,N_5365);
and U6046 (N_6046,N_5016,N_5639);
and U6047 (N_6047,N_5247,N_5137);
xor U6048 (N_6048,N_5729,N_5650);
or U6049 (N_6049,N_5311,N_5420);
nand U6050 (N_6050,N_5698,N_5635);
or U6051 (N_6051,N_5254,N_5696);
or U6052 (N_6052,N_5569,N_5480);
nand U6053 (N_6053,N_5000,N_5516);
nor U6054 (N_6054,N_5161,N_5323);
xnor U6055 (N_6055,N_5888,N_5526);
xnor U6056 (N_6056,N_5229,N_5900);
or U6057 (N_6057,N_5005,N_5822);
nor U6058 (N_6058,N_5290,N_5007);
and U6059 (N_6059,N_5914,N_5275);
or U6060 (N_6060,N_5391,N_5720);
and U6061 (N_6061,N_5707,N_5501);
nor U6062 (N_6062,N_5351,N_5456);
or U6063 (N_6063,N_5417,N_5641);
nor U6064 (N_6064,N_5775,N_5879);
xor U6065 (N_6065,N_5219,N_5087);
xor U6066 (N_6066,N_5562,N_5405);
nand U6067 (N_6067,N_5477,N_5803);
nor U6068 (N_6068,N_5437,N_5776);
or U6069 (N_6069,N_5515,N_5436);
nand U6070 (N_6070,N_5884,N_5172);
and U6071 (N_6071,N_5249,N_5622);
nor U6072 (N_6072,N_5142,N_5856);
and U6073 (N_6073,N_5487,N_5727);
xor U6074 (N_6074,N_5874,N_5394);
nor U6075 (N_6075,N_5300,N_5403);
and U6076 (N_6076,N_5586,N_5740);
and U6077 (N_6077,N_5925,N_5072);
or U6078 (N_6078,N_5910,N_5442);
and U6079 (N_6079,N_5447,N_5647);
nor U6080 (N_6080,N_5689,N_5908);
xor U6081 (N_6081,N_5844,N_5415);
xnor U6082 (N_6082,N_5816,N_5322);
xnor U6083 (N_6083,N_5002,N_5400);
xor U6084 (N_6084,N_5426,N_5140);
xnor U6085 (N_6085,N_5631,N_5629);
nand U6086 (N_6086,N_5202,N_5327);
and U6087 (N_6087,N_5319,N_5469);
nor U6088 (N_6088,N_5330,N_5279);
xor U6089 (N_6089,N_5329,N_5228);
and U6090 (N_6090,N_5694,N_5760);
xor U6091 (N_6091,N_5014,N_5714);
or U6092 (N_6092,N_5939,N_5281);
nand U6093 (N_6093,N_5494,N_5320);
and U6094 (N_6094,N_5089,N_5158);
nor U6095 (N_6095,N_5560,N_5283);
nand U6096 (N_6096,N_5781,N_5035);
nor U6097 (N_6097,N_5991,N_5658);
or U6098 (N_6098,N_5739,N_5163);
or U6099 (N_6099,N_5663,N_5178);
nor U6100 (N_6100,N_5445,N_5444);
or U6101 (N_6101,N_5704,N_5924);
xor U6102 (N_6102,N_5069,N_5620);
or U6103 (N_6103,N_5837,N_5962);
xnor U6104 (N_6104,N_5056,N_5601);
and U6105 (N_6105,N_5062,N_5798);
nor U6106 (N_6106,N_5738,N_5113);
xnor U6107 (N_6107,N_5921,N_5397);
nor U6108 (N_6108,N_5768,N_5093);
xor U6109 (N_6109,N_5258,N_5474);
or U6110 (N_6110,N_5999,N_5855);
or U6111 (N_6111,N_5270,N_5173);
or U6112 (N_6112,N_5644,N_5773);
nor U6113 (N_6113,N_5162,N_5481);
or U6114 (N_6114,N_5237,N_5745);
nor U6115 (N_6115,N_5116,N_5675);
xnor U6116 (N_6116,N_5091,N_5335);
nor U6117 (N_6117,N_5911,N_5842);
xor U6118 (N_6118,N_5957,N_5027);
and U6119 (N_6119,N_5883,N_5595);
nand U6120 (N_6120,N_5122,N_5559);
xor U6121 (N_6121,N_5699,N_5554);
xnor U6122 (N_6122,N_5592,N_5572);
and U6123 (N_6123,N_5220,N_5536);
xnor U6124 (N_6124,N_5829,N_5066);
or U6125 (N_6125,N_5728,N_5363);
xor U6126 (N_6126,N_5078,N_5287);
nor U6127 (N_6127,N_5128,N_5204);
nand U6128 (N_6128,N_5134,N_5511);
nand U6129 (N_6129,N_5333,N_5661);
nand U6130 (N_6130,N_5857,N_5733);
xor U6131 (N_6131,N_5555,N_5503);
nand U6132 (N_6132,N_5968,N_5302);
nor U6133 (N_6133,N_5778,N_5257);
or U6134 (N_6134,N_5668,N_5373);
xnor U6135 (N_6135,N_5763,N_5731);
and U6136 (N_6136,N_5199,N_5434);
xnor U6137 (N_6137,N_5086,N_5826);
nor U6138 (N_6138,N_5787,N_5549);
and U6139 (N_6139,N_5930,N_5467);
or U6140 (N_6140,N_5383,N_5607);
nand U6141 (N_6141,N_5783,N_5265);
nor U6142 (N_6142,N_5682,N_5677);
nand U6143 (N_6143,N_5651,N_5625);
nand U6144 (N_6144,N_5095,N_5824);
xor U6145 (N_6145,N_5479,N_5929);
nand U6146 (N_6146,N_5044,N_5749);
or U6147 (N_6147,N_5736,N_5368);
nand U6148 (N_6148,N_5036,N_5893);
xor U6149 (N_6149,N_5211,N_5491);
nand U6150 (N_6150,N_5193,N_5818);
or U6151 (N_6151,N_5815,N_5359);
nor U6152 (N_6152,N_5847,N_5422);
and U6153 (N_6153,N_5107,N_5340);
or U6154 (N_6154,N_5186,N_5049);
and U6155 (N_6155,N_5100,N_5697);
nor U6156 (N_6156,N_5156,N_5573);
xor U6157 (N_6157,N_5166,N_5780);
nor U6158 (N_6158,N_5315,N_5975);
or U6159 (N_6159,N_5372,N_5721);
or U6160 (N_6160,N_5440,N_5344);
or U6161 (N_6161,N_5965,N_5077);
and U6162 (N_6162,N_5753,N_5180);
or U6163 (N_6163,N_5756,N_5409);
xnor U6164 (N_6164,N_5244,N_5752);
xnor U6165 (N_6165,N_5075,N_5135);
and U6166 (N_6166,N_5332,N_5458);
or U6167 (N_6167,N_5061,N_5292);
and U6168 (N_6168,N_5927,N_5291);
and U6169 (N_6169,N_5343,N_5098);
xor U6170 (N_6170,N_5746,N_5609);
nand U6171 (N_6171,N_5854,N_5765);
nand U6172 (N_6172,N_5695,N_5613);
nor U6173 (N_6173,N_5490,N_5297);
or U6174 (N_6174,N_5782,N_5424);
xor U6175 (N_6175,N_5722,N_5981);
nor U6176 (N_6176,N_5769,N_5051);
or U6177 (N_6177,N_5341,N_5115);
and U6178 (N_6178,N_5621,N_5596);
xor U6179 (N_6179,N_5942,N_5608);
nor U6180 (N_6180,N_5127,N_5179);
xor U6181 (N_6181,N_5779,N_5788);
or U6182 (N_6182,N_5187,N_5809);
xor U6183 (N_6183,N_5513,N_5169);
nor U6184 (N_6184,N_5662,N_5529);
nand U6185 (N_6185,N_5149,N_5982);
nand U6186 (N_6186,N_5561,N_5239);
or U6187 (N_6187,N_5468,N_5386);
nor U6188 (N_6188,N_5324,N_5589);
and U6189 (N_6189,N_5741,N_5170);
and U6190 (N_6190,N_5730,N_5548);
nor U6191 (N_6191,N_5144,N_5402);
or U6192 (N_6192,N_5584,N_5364);
nand U6193 (N_6193,N_5509,N_5508);
xor U6194 (N_6194,N_5438,N_5146);
nor U6195 (N_6195,N_5500,N_5719);
nand U6196 (N_6196,N_5977,N_5793);
xnor U6197 (N_6197,N_5421,N_5308);
nor U6198 (N_6198,N_5578,N_5869);
xor U6199 (N_6199,N_5159,N_5316);
nand U6200 (N_6200,N_5843,N_5284);
or U6201 (N_6201,N_5744,N_5819);
or U6202 (N_6202,N_5232,N_5309);
xor U6203 (N_6203,N_5686,N_5011);
xor U6204 (N_6204,N_5129,N_5935);
xor U6205 (N_6205,N_5439,N_5519);
or U6206 (N_6206,N_5304,N_5797);
and U6207 (N_6207,N_5902,N_5737);
nand U6208 (N_6208,N_5659,N_5286);
xor U6209 (N_6209,N_5952,N_5611);
nor U6210 (N_6210,N_5633,N_5416);
or U6211 (N_6211,N_5814,N_5425);
nor U6212 (N_6212,N_5392,N_5583);
or U6213 (N_6213,N_5209,N_5587);
nor U6214 (N_6214,N_5985,N_5546);
nand U6215 (N_6215,N_5638,N_5015);
nor U6216 (N_6216,N_5345,N_5045);
nand U6217 (N_6217,N_5461,N_5064);
xor U6218 (N_6218,N_5030,N_5138);
nor U6219 (N_6219,N_5412,N_5514);
or U6220 (N_6220,N_5222,N_5070);
or U6221 (N_6221,N_5916,N_5101);
and U6222 (N_6222,N_5922,N_5471);
nand U6223 (N_6223,N_5387,N_5691);
nand U6224 (N_6224,N_5221,N_5382);
xnor U6225 (N_6225,N_5565,N_5654);
or U6226 (N_6226,N_5716,N_5591);
nor U6227 (N_6227,N_5881,N_5873);
and U6228 (N_6228,N_5557,N_5314);
nor U6229 (N_6229,N_5260,N_5664);
nand U6230 (N_6230,N_5154,N_5111);
and U6231 (N_6231,N_5360,N_5834);
or U6232 (N_6232,N_5032,N_5648);
nand U6233 (N_6233,N_5785,N_5758);
xor U6234 (N_6234,N_5057,N_5810);
nor U6235 (N_6235,N_5994,N_5451);
nand U6236 (N_6236,N_5423,N_5362);
xnor U6237 (N_6237,N_5058,N_5210);
nand U6238 (N_6238,N_5090,N_5564);
or U6239 (N_6239,N_5357,N_5846);
and U6240 (N_6240,N_5031,N_5454);
and U6241 (N_6241,N_5264,N_5742);
and U6242 (N_6242,N_5504,N_5606);
or U6243 (N_6243,N_5577,N_5242);
nor U6244 (N_6244,N_5342,N_5540);
and U6245 (N_6245,N_5380,N_5983);
nand U6246 (N_6246,N_5996,N_5570);
xor U6247 (N_6247,N_5836,N_5688);
and U6248 (N_6248,N_5667,N_5023);
or U6249 (N_6249,N_5282,N_5462);
nor U6250 (N_6250,N_5823,N_5196);
and U6251 (N_6251,N_5871,N_5407);
nor U6252 (N_6252,N_5643,N_5995);
or U6253 (N_6253,N_5499,N_5528);
nor U6254 (N_6254,N_5096,N_5390);
nand U6255 (N_6255,N_5640,N_5896);
and U6256 (N_6256,N_5931,N_5547);
and U6257 (N_6257,N_5612,N_5894);
and U6258 (N_6258,N_5301,N_5936);
and U6259 (N_6259,N_5892,N_5711);
or U6260 (N_6260,N_5259,N_5317);
nor U6261 (N_6261,N_5618,N_5724);
nor U6262 (N_6262,N_5414,N_5396);
or U6263 (N_6263,N_5273,N_5478);
nor U6264 (N_6264,N_5940,N_5551);
nand U6265 (N_6265,N_5533,N_5568);
xor U6266 (N_6266,N_5886,N_5959);
nand U6267 (N_6267,N_5832,N_5255);
nor U6268 (N_6268,N_5218,N_5603);
nor U6269 (N_6269,N_5791,N_5294);
xor U6270 (N_6270,N_5806,N_5794);
nor U6271 (N_6271,N_5450,N_5945);
and U6272 (N_6272,N_5401,N_5191);
nor U6273 (N_6273,N_5073,N_5076);
nand U6274 (N_6274,N_5493,N_5251);
and U6275 (N_6275,N_5971,N_5545);
nand U6276 (N_6276,N_5862,N_5998);
nor U6277 (N_6277,N_5148,N_5899);
and U6278 (N_6278,N_5880,N_5448);
or U6279 (N_6279,N_5762,N_5097);
xor U6280 (N_6280,N_5817,N_5961);
and U6281 (N_6281,N_5708,N_5923);
and U6282 (N_6282,N_5628,N_5106);
nor U6283 (N_6283,N_5712,N_5216);
xnor U6284 (N_6284,N_5904,N_5067);
xor U6285 (N_6285,N_5130,N_5379);
nand U6286 (N_6286,N_5771,N_5475);
nand U6287 (N_6287,N_5404,N_5831);
and U6288 (N_6288,N_5864,N_5679);
xnor U6289 (N_6289,N_5054,N_5060);
nor U6290 (N_6290,N_5271,N_5670);
and U6291 (N_6291,N_5920,N_5710);
or U6292 (N_6292,N_5807,N_5845);
nor U6293 (N_6293,N_5512,N_5534);
nand U6294 (N_6294,N_5331,N_5151);
or U6295 (N_6295,N_5988,N_5687);
xor U6296 (N_6296,N_5152,N_5653);
or U6297 (N_6297,N_5885,N_5976);
nor U6298 (N_6298,N_5074,N_5759);
nor U6299 (N_6299,N_5206,N_5969);
or U6300 (N_6300,N_5732,N_5784);
xnor U6301 (N_6301,N_5010,N_5878);
xor U6302 (N_6302,N_5001,N_5223);
and U6303 (N_6303,N_5347,N_5388);
xnor U6304 (N_6304,N_5684,N_5796);
nand U6305 (N_6305,N_5019,N_5928);
or U6306 (N_6306,N_5234,N_5553);
and U6307 (N_6307,N_5944,N_5427);
or U6308 (N_6308,N_5226,N_5895);
or U6309 (N_6309,N_5435,N_5262);
and U6310 (N_6310,N_5860,N_5167);
and U6311 (N_6311,N_5446,N_5757);
or U6312 (N_6312,N_5616,N_5039);
nor U6313 (N_6313,N_5043,N_5483);
nand U6314 (N_6314,N_5808,N_5970);
nor U6315 (N_6315,N_5012,N_5120);
xnor U6316 (N_6316,N_5486,N_5839);
nand U6317 (N_6317,N_5141,N_5046);
and U6318 (N_6318,N_5498,N_5430);
xnor U6319 (N_6319,N_5354,N_5906);
nor U6320 (N_6320,N_5681,N_5747);
nor U6321 (N_6321,N_5033,N_5393);
nor U6322 (N_6322,N_5600,N_5418);
and U6323 (N_6323,N_5201,N_5979);
and U6324 (N_6324,N_5353,N_5212);
nand U6325 (N_6325,N_5177,N_5602);
nand U6326 (N_6326,N_5092,N_5718);
nand U6327 (N_6327,N_5558,N_5157);
and U6328 (N_6328,N_5109,N_5850);
nand U6329 (N_6329,N_5104,N_5766);
nor U6330 (N_6330,N_5048,N_5571);
or U6331 (N_6331,N_5133,N_5725);
nor U6332 (N_6332,N_5838,N_5610);
nand U6333 (N_6333,N_5813,N_5358);
nand U6334 (N_6334,N_5812,N_5029);
nor U6335 (N_6335,N_5110,N_5642);
xnor U6336 (N_6336,N_5953,N_5574);
nand U6337 (N_6337,N_5346,N_5901);
nand U6338 (N_6338,N_5443,N_5693);
or U6339 (N_6339,N_5059,N_5851);
and U6340 (N_6340,N_5750,N_5160);
and U6341 (N_6341,N_5374,N_5950);
and U6342 (N_6342,N_5713,N_5099);
and U6343 (N_6343,N_5195,N_5102);
or U6344 (N_6344,N_5108,N_5626);
or U6345 (N_6345,N_5371,N_5470);
xor U6346 (N_6346,N_5080,N_5868);
nor U6347 (N_6347,N_5634,N_5188);
xnor U6348 (N_6348,N_5419,N_5800);
or U6349 (N_6349,N_5941,N_5355);
xnor U6350 (N_6350,N_5224,N_5947);
xnor U6351 (N_6351,N_5071,N_5268);
xor U6352 (N_6352,N_5466,N_5293);
nand U6353 (N_6353,N_5325,N_5482);
nand U6354 (N_6354,N_5198,N_5966);
xnor U6355 (N_6355,N_5025,N_5041);
nand U6356 (N_6356,N_5225,N_5084);
and U6357 (N_6357,N_5537,N_5337);
xor U6358 (N_6358,N_5535,N_5789);
or U6359 (N_6359,N_5476,N_5948);
and U6360 (N_6360,N_5717,N_5361);
and U6361 (N_6361,N_5336,N_5990);
nand U6362 (N_6362,N_5182,N_5835);
and U6363 (N_6363,N_5926,N_5656);
nor U6364 (N_6364,N_5024,N_5987);
xnor U6365 (N_6365,N_5770,N_5865);
and U6366 (N_6366,N_5636,N_5280);
nand U6367 (N_6367,N_5655,N_5665);
xnor U6368 (N_6368,N_5124,N_5986);
nor U6369 (N_6369,N_5520,N_5413);
or U6370 (N_6370,N_5021,N_5811);
xnor U6371 (N_6371,N_5126,N_5754);
xor U6372 (N_6372,N_5938,N_5666);
nor U6373 (N_6373,N_5683,N_5243);
or U6374 (N_6374,N_5804,N_5575);
or U6375 (N_6375,N_5082,N_5709);
or U6376 (N_6376,N_5118,N_5453);
or U6377 (N_6377,N_5949,N_5830);
xnor U6378 (N_6378,N_5701,N_5624);
nand U6379 (N_6379,N_5312,N_5411);
nor U6380 (N_6380,N_5326,N_5518);
nand U6381 (N_6381,N_5457,N_5594);
or U6382 (N_6382,N_5020,N_5278);
xnor U6383 (N_6383,N_5524,N_5303);
nand U6384 (N_6384,N_5081,N_5703);
xnor U6385 (N_6385,N_5828,N_5492);
nor U6386 (N_6386,N_5805,N_5205);
and U6387 (N_6387,N_5334,N_5772);
and U6388 (N_6388,N_5013,N_5338);
nor U6389 (N_6389,N_5370,N_5907);
and U6390 (N_6390,N_5495,N_5245);
or U6391 (N_6391,N_5532,N_5252);
xor U6392 (N_6392,N_5552,N_5381);
nor U6393 (N_6393,N_5256,N_5685);
and U6394 (N_6394,N_5867,N_5841);
or U6395 (N_6395,N_5992,N_5285);
xnor U6396 (N_6396,N_5406,N_5429);
nor U6397 (N_6397,N_5165,N_5877);
xnor U6398 (N_6398,N_5531,N_5250);
xnor U6399 (N_6399,N_5673,N_5734);
xor U6400 (N_6400,N_5802,N_5550);
and U6401 (N_6401,N_5184,N_5008);
nand U6402 (N_6402,N_5085,N_5542);
and U6403 (N_6403,N_5496,N_5506);
and U6404 (N_6404,N_5660,N_5706);
nor U6405 (N_6405,N_5876,N_5003);
xnor U6406 (N_6406,N_5777,N_5764);
or U6407 (N_6407,N_5428,N_5034);
nand U6408 (N_6408,N_5897,N_5863);
nor U6409 (N_6409,N_5891,N_5185);
or U6410 (N_6410,N_5678,N_5181);
nor U6411 (N_6411,N_5748,N_5527);
nand U6412 (N_6412,N_5974,N_5645);
or U6413 (N_6413,N_5866,N_5859);
and U6414 (N_6414,N_5544,N_5472);
nor U6415 (N_6415,N_5117,N_5702);
nor U6416 (N_6416,N_5269,N_5580);
and U6417 (N_6417,N_5700,N_5114);
nand U6418 (N_6418,N_5964,N_5581);
or U6419 (N_6419,N_5517,N_5313);
nand U6420 (N_6420,N_5649,N_5530);
xor U6421 (N_6421,N_5261,N_5539);
and U6422 (N_6422,N_5617,N_5604);
and U6423 (N_6423,N_5143,N_5236);
nor U6424 (N_6424,N_5194,N_5006);
nor U6425 (N_6425,N_5088,N_5022);
or U6426 (N_6426,N_5852,N_5318);
nor U6427 (N_6427,N_5473,N_5328);
and U6428 (N_6428,N_5882,N_5465);
and U6429 (N_6429,N_5488,N_5671);
xor U6430 (N_6430,N_5213,N_5253);
nand U6431 (N_6431,N_5352,N_5395);
nand U6432 (N_6432,N_5004,N_5605);
and U6433 (N_6433,N_5585,N_5183);
nand U6434 (N_6434,N_5235,N_5593);
and U6435 (N_6435,N_5522,N_5464);
nor U6436 (N_6436,N_5378,N_5433);
nand U6437 (N_6437,N_5954,N_5176);
and U6438 (N_6438,N_5848,N_5875);
and U6439 (N_6439,N_5267,N_5960);
and U6440 (N_6440,N_5853,N_5538);
and U6441 (N_6441,N_5657,N_5646);
nor U6442 (N_6442,N_5040,N_5028);
xnor U6443 (N_6443,N_5761,N_5125);
nand U6444 (N_6444,N_5083,N_5321);
nand U6445 (N_6445,N_5399,N_5356);
nand U6446 (N_6446,N_5913,N_5563);
nor U6447 (N_6447,N_5972,N_5967);
or U6448 (N_6448,N_5018,N_5795);
nand U6449 (N_6449,N_5890,N_5432);
or U6450 (N_6450,N_5672,N_5576);
and U6451 (N_6451,N_5690,N_5230);
nor U6452 (N_6452,N_5774,N_5103);
xnor U6453 (N_6453,N_5246,N_5145);
and U6454 (N_6454,N_5455,N_5307);
and U6455 (N_6455,N_5825,N_5932);
xor U6456 (N_6456,N_5119,N_5597);
nand U6457 (N_6457,N_5288,N_5567);
nor U6458 (N_6458,N_5956,N_5042);
xor U6459 (N_6459,N_5521,N_5973);
nor U6460 (N_6460,N_5858,N_5276);
and U6461 (N_6461,N_5459,N_5463);
or U6462 (N_6462,N_5958,N_5903);
xor U6463 (N_6463,N_5277,N_5946);
or U6464 (N_6464,N_5037,N_5385);
and U6465 (N_6465,N_5306,N_5497);
nor U6466 (N_6466,N_5068,N_5289);
nand U6467 (N_6467,N_5735,N_5510);
or U6468 (N_6468,N_5155,N_5150);
nor U6469 (N_6469,N_5310,N_5431);
xnor U6470 (N_6470,N_5556,N_5203);
or U6471 (N_6471,N_5887,N_5123);
and U6472 (N_6472,N_5055,N_5227);
xor U6473 (N_6473,N_5410,N_5017);
nand U6474 (N_6474,N_5543,N_5792);
or U6475 (N_6475,N_5296,N_5937);
nand U6476 (N_6476,N_5052,N_5214);
xnor U6477 (N_6477,N_5614,N_5790);
or U6478 (N_6478,N_5872,N_5502);
nor U6479 (N_6479,N_5139,N_5369);
or U6480 (N_6480,N_5305,N_5723);
and U6481 (N_6481,N_5200,N_5751);
xor U6482 (N_6482,N_5705,N_5377);
nor U6483 (N_6483,N_5299,N_5637);
xor U6484 (N_6484,N_5955,N_5669);
xor U6485 (N_6485,N_5963,N_5063);
xnor U6486 (N_6486,N_5384,N_5238);
nand U6487 (N_6487,N_5295,N_5348);
or U6488 (N_6488,N_5398,N_5680);
nor U6489 (N_6489,N_5632,N_5821);
and U6490 (N_6490,N_5207,N_5588);
or U6491 (N_6491,N_5918,N_5217);
nor U6492 (N_6492,N_5861,N_5984);
and U6493 (N_6493,N_5505,N_5523);
nand U6494 (N_6494,N_5599,N_5174);
nand U6495 (N_6495,N_5263,N_5951);
or U6496 (N_6496,N_5943,N_5674);
nand U6497 (N_6497,N_5449,N_5408);
nand U6498 (N_6498,N_5136,N_5164);
nand U6499 (N_6499,N_5997,N_5840);
or U6500 (N_6500,N_5385,N_5594);
nand U6501 (N_6501,N_5072,N_5223);
nand U6502 (N_6502,N_5883,N_5076);
or U6503 (N_6503,N_5498,N_5936);
nand U6504 (N_6504,N_5358,N_5209);
nand U6505 (N_6505,N_5315,N_5852);
nor U6506 (N_6506,N_5352,N_5599);
or U6507 (N_6507,N_5222,N_5104);
xnor U6508 (N_6508,N_5009,N_5084);
xnor U6509 (N_6509,N_5410,N_5890);
nand U6510 (N_6510,N_5644,N_5647);
xor U6511 (N_6511,N_5018,N_5719);
and U6512 (N_6512,N_5738,N_5529);
xor U6513 (N_6513,N_5826,N_5430);
and U6514 (N_6514,N_5657,N_5980);
or U6515 (N_6515,N_5199,N_5995);
and U6516 (N_6516,N_5742,N_5692);
nand U6517 (N_6517,N_5543,N_5168);
xnor U6518 (N_6518,N_5120,N_5053);
or U6519 (N_6519,N_5375,N_5021);
nor U6520 (N_6520,N_5733,N_5752);
nand U6521 (N_6521,N_5644,N_5837);
nand U6522 (N_6522,N_5354,N_5628);
nor U6523 (N_6523,N_5159,N_5092);
xor U6524 (N_6524,N_5941,N_5589);
and U6525 (N_6525,N_5386,N_5185);
xnor U6526 (N_6526,N_5965,N_5034);
and U6527 (N_6527,N_5910,N_5526);
xnor U6528 (N_6528,N_5150,N_5730);
and U6529 (N_6529,N_5830,N_5282);
and U6530 (N_6530,N_5527,N_5719);
nor U6531 (N_6531,N_5386,N_5237);
or U6532 (N_6532,N_5447,N_5905);
or U6533 (N_6533,N_5262,N_5107);
and U6534 (N_6534,N_5365,N_5664);
or U6535 (N_6535,N_5984,N_5279);
xnor U6536 (N_6536,N_5584,N_5051);
and U6537 (N_6537,N_5080,N_5006);
xor U6538 (N_6538,N_5050,N_5321);
nand U6539 (N_6539,N_5761,N_5129);
nor U6540 (N_6540,N_5740,N_5455);
nor U6541 (N_6541,N_5879,N_5893);
nor U6542 (N_6542,N_5492,N_5959);
or U6543 (N_6543,N_5520,N_5574);
xor U6544 (N_6544,N_5504,N_5888);
xor U6545 (N_6545,N_5764,N_5197);
or U6546 (N_6546,N_5510,N_5084);
nor U6547 (N_6547,N_5722,N_5325);
nand U6548 (N_6548,N_5049,N_5328);
or U6549 (N_6549,N_5581,N_5518);
xor U6550 (N_6550,N_5516,N_5715);
and U6551 (N_6551,N_5934,N_5960);
or U6552 (N_6552,N_5287,N_5092);
and U6553 (N_6553,N_5677,N_5789);
or U6554 (N_6554,N_5504,N_5524);
nand U6555 (N_6555,N_5358,N_5384);
or U6556 (N_6556,N_5115,N_5011);
nor U6557 (N_6557,N_5813,N_5462);
nand U6558 (N_6558,N_5421,N_5037);
and U6559 (N_6559,N_5499,N_5663);
xnor U6560 (N_6560,N_5078,N_5055);
and U6561 (N_6561,N_5467,N_5596);
or U6562 (N_6562,N_5297,N_5312);
xor U6563 (N_6563,N_5307,N_5196);
xor U6564 (N_6564,N_5914,N_5520);
nor U6565 (N_6565,N_5679,N_5232);
nand U6566 (N_6566,N_5059,N_5550);
xor U6567 (N_6567,N_5020,N_5701);
nand U6568 (N_6568,N_5774,N_5802);
xor U6569 (N_6569,N_5179,N_5051);
nand U6570 (N_6570,N_5072,N_5121);
or U6571 (N_6571,N_5127,N_5526);
nor U6572 (N_6572,N_5052,N_5999);
nand U6573 (N_6573,N_5813,N_5341);
nand U6574 (N_6574,N_5726,N_5453);
and U6575 (N_6575,N_5562,N_5242);
xnor U6576 (N_6576,N_5212,N_5871);
or U6577 (N_6577,N_5303,N_5733);
nand U6578 (N_6578,N_5813,N_5756);
xor U6579 (N_6579,N_5796,N_5219);
xnor U6580 (N_6580,N_5206,N_5144);
and U6581 (N_6581,N_5680,N_5068);
and U6582 (N_6582,N_5944,N_5398);
nor U6583 (N_6583,N_5237,N_5096);
nor U6584 (N_6584,N_5993,N_5479);
or U6585 (N_6585,N_5043,N_5883);
nand U6586 (N_6586,N_5427,N_5683);
xnor U6587 (N_6587,N_5995,N_5933);
xor U6588 (N_6588,N_5880,N_5153);
and U6589 (N_6589,N_5696,N_5881);
and U6590 (N_6590,N_5857,N_5310);
nor U6591 (N_6591,N_5408,N_5349);
xor U6592 (N_6592,N_5730,N_5780);
nand U6593 (N_6593,N_5875,N_5902);
or U6594 (N_6594,N_5676,N_5835);
nand U6595 (N_6595,N_5773,N_5137);
or U6596 (N_6596,N_5532,N_5727);
nor U6597 (N_6597,N_5076,N_5934);
nand U6598 (N_6598,N_5151,N_5399);
nand U6599 (N_6599,N_5166,N_5617);
and U6600 (N_6600,N_5537,N_5843);
and U6601 (N_6601,N_5067,N_5546);
and U6602 (N_6602,N_5211,N_5532);
nor U6603 (N_6603,N_5083,N_5757);
nand U6604 (N_6604,N_5154,N_5770);
and U6605 (N_6605,N_5664,N_5318);
and U6606 (N_6606,N_5181,N_5251);
xnor U6607 (N_6607,N_5874,N_5964);
nor U6608 (N_6608,N_5242,N_5943);
and U6609 (N_6609,N_5532,N_5908);
nor U6610 (N_6610,N_5248,N_5453);
and U6611 (N_6611,N_5816,N_5514);
and U6612 (N_6612,N_5070,N_5627);
and U6613 (N_6613,N_5621,N_5912);
and U6614 (N_6614,N_5405,N_5549);
or U6615 (N_6615,N_5932,N_5826);
or U6616 (N_6616,N_5008,N_5049);
nor U6617 (N_6617,N_5062,N_5324);
nand U6618 (N_6618,N_5496,N_5932);
or U6619 (N_6619,N_5073,N_5910);
or U6620 (N_6620,N_5689,N_5286);
nand U6621 (N_6621,N_5846,N_5380);
and U6622 (N_6622,N_5496,N_5007);
and U6623 (N_6623,N_5143,N_5272);
nor U6624 (N_6624,N_5287,N_5966);
or U6625 (N_6625,N_5820,N_5658);
xnor U6626 (N_6626,N_5235,N_5976);
nand U6627 (N_6627,N_5985,N_5876);
nor U6628 (N_6628,N_5946,N_5742);
nor U6629 (N_6629,N_5610,N_5972);
nor U6630 (N_6630,N_5284,N_5659);
and U6631 (N_6631,N_5612,N_5564);
or U6632 (N_6632,N_5242,N_5254);
nand U6633 (N_6633,N_5453,N_5688);
and U6634 (N_6634,N_5468,N_5560);
xor U6635 (N_6635,N_5197,N_5128);
or U6636 (N_6636,N_5115,N_5420);
and U6637 (N_6637,N_5685,N_5468);
nor U6638 (N_6638,N_5302,N_5520);
and U6639 (N_6639,N_5147,N_5270);
or U6640 (N_6640,N_5916,N_5052);
xnor U6641 (N_6641,N_5729,N_5593);
or U6642 (N_6642,N_5678,N_5061);
nand U6643 (N_6643,N_5619,N_5489);
nand U6644 (N_6644,N_5234,N_5984);
or U6645 (N_6645,N_5964,N_5296);
and U6646 (N_6646,N_5510,N_5680);
xnor U6647 (N_6647,N_5471,N_5667);
nor U6648 (N_6648,N_5588,N_5442);
nand U6649 (N_6649,N_5600,N_5288);
or U6650 (N_6650,N_5297,N_5232);
nor U6651 (N_6651,N_5659,N_5141);
and U6652 (N_6652,N_5251,N_5692);
and U6653 (N_6653,N_5612,N_5887);
nand U6654 (N_6654,N_5482,N_5690);
and U6655 (N_6655,N_5102,N_5072);
nand U6656 (N_6656,N_5766,N_5038);
nor U6657 (N_6657,N_5738,N_5315);
nor U6658 (N_6658,N_5573,N_5496);
or U6659 (N_6659,N_5226,N_5097);
and U6660 (N_6660,N_5608,N_5105);
or U6661 (N_6661,N_5240,N_5885);
xor U6662 (N_6662,N_5591,N_5101);
or U6663 (N_6663,N_5467,N_5599);
and U6664 (N_6664,N_5502,N_5547);
nor U6665 (N_6665,N_5635,N_5445);
or U6666 (N_6666,N_5882,N_5632);
nand U6667 (N_6667,N_5066,N_5902);
nand U6668 (N_6668,N_5169,N_5956);
and U6669 (N_6669,N_5868,N_5182);
and U6670 (N_6670,N_5419,N_5370);
and U6671 (N_6671,N_5276,N_5767);
xor U6672 (N_6672,N_5505,N_5922);
and U6673 (N_6673,N_5247,N_5376);
nor U6674 (N_6674,N_5876,N_5634);
and U6675 (N_6675,N_5839,N_5429);
or U6676 (N_6676,N_5884,N_5314);
and U6677 (N_6677,N_5912,N_5355);
xnor U6678 (N_6678,N_5210,N_5012);
and U6679 (N_6679,N_5172,N_5164);
nand U6680 (N_6680,N_5530,N_5923);
nand U6681 (N_6681,N_5575,N_5326);
or U6682 (N_6682,N_5414,N_5332);
or U6683 (N_6683,N_5091,N_5723);
xor U6684 (N_6684,N_5114,N_5135);
or U6685 (N_6685,N_5826,N_5222);
nand U6686 (N_6686,N_5863,N_5939);
xnor U6687 (N_6687,N_5783,N_5073);
nor U6688 (N_6688,N_5883,N_5127);
nor U6689 (N_6689,N_5677,N_5982);
and U6690 (N_6690,N_5401,N_5651);
or U6691 (N_6691,N_5787,N_5258);
nor U6692 (N_6692,N_5648,N_5763);
nand U6693 (N_6693,N_5064,N_5660);
nor U6694 (N_6694,N_5577,N_5200);
and U6695 (N_6695,N_5811,N_5817);
nand U6696 (N_6696,N_5859,N_5156);
xor U6697 (N_6697,N_5666,N_5863);
nand U6698 (N_6698,N_5729,N_5841);
or U6699 (N_6699,N_5637,N_5314);
nor U6700 (N_6700,N_5900,N_5756);
and U6701 (N_6701,N_5892,N_5425);
nor U6702 (N_6702,N_5506,N_5821);
and U6703 (N_6703,N_5225,N_5625);
nand U6704 (N_6704,N_5469,N_5597);
nor U6705 (N_6705,N_5733,N_5539);
and U6706 (N_6706,N_5737,N_5371);
nor U6707 (N_6707,N_5987,N_5564);
nor U6708 (N_6708,N_5874,N_5568);
xnor U6709 (N_6709,N_5689,N_5679);
nand U6710 (N_6710,N_5370,N_5834);
nor U6711 (N_6711,N_5248,N_5865);
xor U6712 (N_6712,N_5595,N_5532);
or U6713 (N_6713,N_5834,N_5979);
nor U6714 (N_6714,N_5695,N_5657);
and U6715 (N_6715,N_5873,N_5443);
xor U6716 (N_6716,N_5496,N_5636);
and U6717 (N_6717,N_5186,N_5047);
or U6718 (N_6718,N_5023,N_5235);
nor U6719 (N_6719,N_5027,N_5570);
or U6720 (N_6720,N_5083,N_5705);
and U6721 (N_6721,N_5180,N_5784);
nand U6722 (N_6722,N_5545,N_5523);
xnor U6723 (N_6723,N_5550,N_5245);
or U6724 (N_6724,N_5960,N_5823);
nor U6725 (N_6725,N_5336,N_5903);
xnor U6726 (N_6726,N_5163,N_5904);
xor U6727 (N_6727,N_5140,N_5191);
nand U6728 (N_6728,N_5823,N_5400);
and U6729 (N_6729,N_5558,N_5465);
nor U6730 (N_6730,N_5377,N_5711);
and U6731 (N_6731,N_5111,N_5547);
or U6732 (N_6732,N_5901,N_5413);
nand U6733 (N_6733,N_5270,N_5409);
nand U6734 (N_6734,N_5014,N_5924);
nand U6735 (N_6735,N_5324,N_5765);
or U6736 (N_6736,N_5973,N_5853);
nor U6737 (N_6737,N_5098,N_5164);
xnor U6738 (N_6738,N_5249,N_5654);
xor U6739 (N_6739,N_5393,N_5791);
xnor U6740 (N_6740,N_5723,N_5238);
xor U6741 (N_6741,N_5280,N_5966);
and U6742 (N_6742,N_5249,N_5594);
nand U6743 (N_6743,N_5687,N_5005);
xnor U6744 (N_6744,N_5025,N_5722);
nand U6745 (N_6745,N_5678,N_5039);
or U6746 (N_6746,N_5202,N_5402);
and U6747 (N_6747,N_5032,N_5624);
nand U6748 (N_6748,N_5110,N_5175);
xnor U6749 (N_6749,N_5866,N_5377);
nor U6750 (N_6750,N_5011,N_5969);
or U6751 (N_6751,N_5642,N_5104);
and U6752 (N_6752,N_5812,N_5042);
nand U6753 (N_6753,N_5361,N_5686);
nor U6754 (N_6754,N_5432,N_5776);
nand U6755 (N_6755,N_5768,N_5877);
nor U6756 (N_6756,N_5905,N_5907);
nor U6757 (N_6757,N_5692,N_5794);
and U6758 (N_6758,N_5134,N_5096);
and U6759 (N_6759,N_5741,N_5768);
nor U6760 (N_6760,N_5916,N_5463);
or U6761 (N_6761,N_5958,N_5990);
and U6762 (N_6762,N_5491,N_5362);
nor U6763 (N_6763,N_5473,N_5181);
and U6764 (N_6764,N_5081,N_5814);
nor U6765 (N_6765,N_5392,N_5389);
nand U6766 (N_6766,N_5194,N_5054);
or U6767 (N_6767,N_5056,N_5503);
or U6768 (N_6768,N_5547,N_5489);
and U6769 (N_6769,N_5647,N_5387);
nor U6770 (N_6770,N_5874,N_5841);
nand U6771 (N_6771,N_5726,N_5718);
xnor U6772 (N_6772,N_5182,N_5620);
nand U6773 (N_6773,N_5460,N_5640);
nand U6774 (N_6774,N_5008,N_5718);
or U6775 (N_6775,N_5628,N_5525);
nand U6776 (N_6776,N_5793,N_5011);
nand U6777 (N_6777,N_5601,N_5668);
xor U6778 (N_6778,N_5403,N_5107);
or U6779 (N_6779,N_5613,N_5832);
xor U6780 (N_6780,N_5292,N_5013);
and U6781 (N_6781,N_5482,N_5036);
or U6782 (N_6782,N_5743,N_5415);
nor U6783 (N_6783,N_5508,N_5684);
xor U6784 (N_6784,N_5821,N_5415);
nor U6785 (N_6785,N_5016,N_5184);
nand U6786 (N_6786,N_5921,N_5889);
nand U6787 (N_6787,N_5935,N_5671);
nand U6788 (N_6788,N_5461,N_5373);
and U6789 (N_6789,N_5360,N_5196);
nand U6790 (N_6790,N_5678,N_5109);
nor U6791 (N_6791,N_5457,N_5890);
xor U6792 (N_6792,N_5031,N_5709);
nand U6793 (N_6793,N_5196,N_5901);
nor U6794 (N_6794,N_5529,N_5217);
and U6795 (N_6795,N_5117,N_5108);
and U6796 (N_6796,N_5485,N_5019);
or U6797 (N_6797,N_5525,N_5483);
xor U6798 (N_6798,N_5646,N_5954);
xor U6799 (N_6799,N_5225,N_5855);
nand U6800 (N_6800,N_5979,N_5764);
or U6801 (N_6801,N_5217,N_5880);
xor U6802 (N_6802,N_5320,N_5850);
nor U6803 (N_6803,N_5195,N_5520);
nor U6804 (N_6804,N_5653,N_5585);
nand U6805 (N_6805,N_5376,N_5673);
xor U6806 (N_6806,N_5486,N_5378);
or U6807 (N_6807,N_5421,N_5720);
and U6808 (N_6808,N_5517,N_5209);
nand U6809 (N_6809,N_5383,N_5910);
xnor U6810 (N_6810,N_5023,N_5476);
or U6811 (N_6811,N_5855,N_5748);
and U6812 (N_6812,N_5558,N_5111);
nand U6813 (N_6813,N_5976,N_5710);
nor U6814 (N_6814,N_5249,N_5003);
nor U6815 (N_6815,N_5797,N_5315);
xor U6816 (N_6816,N_5211,N_5179);
xnor U6817 (N_6817,N_5116,N_5744);
nand U6818 (N_6818,N_5719,N_5910);
and U6819 (N_6819,N_5851,N_5265);
nor U6820 (N_6820,N_5530,N_5116);
and U6821 (N_6821,N_5342,N_5450);
xor U6822 (N_6822,N_5532,N_5875);
xor U6823 (N_6823,N_5487,N_5443);
or U6824 (N_6824,N_5358,N_5677);
xor U6825 (N_6825,N_5148,N_5222);
or U6826 (N_6826,N_5996,N_5766);
nand U6827 (N_6827,N_5513,N_5610);
and U6828 (N_6828,N_5230,N_5176);
nor U6829 (N_6829,N_5377,N_5687);
xnor U6830 (N_6830,N_5321,N_5745);
or U6831 (N_6831,N_5128,N_5744);
nand U6832 (N_6832,N_5118,N_5876);
nor U6833 (N_6833,N_5989,N_5070);
nand U6834 (N_6834,N_5582,N_5717);
xnor U6835 (N_6835,N_5972,N_5306);
and U6836 (N_6836,N_5801,N_5016);
and U6837 (N_6837,N_5257,N_5834);
or U6838 (N_6838,N_5635,N_5542);
nor U6839 (N_6839,N_5586,N_5574);
nand U6840 (N_6840,N_5668,N_5357);
nand U6841 (N_6841,N_5570,N_5660);
xnor U6842 (N_6842,N_5034,N_5174);
and U6843 (N_6843,N_5284,N_5468);
xnor U6844 (N_6844,N_5679,N_5885);
xnor U6845 (N_6845,N_5340,N_5460);
xor U6846 (N_6846,N_5407,N_5501);
nor U6847 (N_6847,N_5250,N_5545);
or U6848 (N_6848,N_5383,N_5975);
nor U6849 (N_6849,N_5377,N_5978);
xnor U6850 (N_6850,N_5990,N_5459);
or U6851 (N_6851,N_5798,N_5357);
or U6852 (N_6852,N_5139,N_5904);
nand U6853 (N_6853,N_5999,N_5628);
and U6854 (N_6854,N_5682,N_5580);
or U6855 (N_6855,N_5628,N_5865);
and U6856 (N_6856,N_5800,N_5054);
nand U6857 (N_6857,N_5084,N_5325);
or U6858 (N_6858,N_5350,N_5997);
and U6859 (N_6859,N_5191,N_5848);
xnor U6860 (N_6860,N_5387,N_5456);
nor U6861 (N_6861,N_5720,N_5521);
nand U6862 (N_6862,N_5370,N_5623);
and U6863 (N_6863,N_5780,N_5078);
or U6864 (N_6864,N_5156,N_5368);
xor U6865 (N_6865,N_5395,N_5899);
or U6866 (N_6866,N_5791,N_5079);
or U6867 (N_6867,N_5881,N_5009);
nand U6868 (N_6868,N_5669,N_5985);
and U6869 (N_6869,N_5234,N_5730);
or U6870 (N_6870,N_5269,N_5569);
nor U6871 (N_6871,N_5331,N_5391);
nor U6872 (N_6872,N_5701,N_5145);
xnor U6873 (N_6873,N_5575,N_5826);
and U6874 (N_6874,N_5342,N_5333);
and U6875 (N_6875,N_5201,N_5806);
xor U6876 (N_6876,N_5517,N_5766);
nor U6877 (N_6877,N_5809,N_5986);
or U6878 (N_6878,N_5349,N_5596);
or U6879 (N_6879,N_5454,N_5447);
nand U6880 (N_6880,N_5728,N_5309);
nand U6881 (N_6881,N_5999,N_5104);
xnor U6882 (N_6882,N_5609,N_5820);
nor U6883 (N_6883,N_5868,N_5383);
or U6884 (N_6884,N_5134,N_5989);
xor U6885 (N_6885,N_5917,N_5419);
xnor U6886 (N_6886,N_5534,N_5429);
nor U6887 (N_6887,N_5635,N_5549);
nor U6888 (N_6888,N_5868,N_5796);
nor U6889 (N_6889,N_5850,N_5709);
and U6890 (N_6890,N_5767,N_5566);
nor U6891 (N_6891,N_5486,N_5748);
xnor U6892 (N_6892,N_5246,N_5778);
and U6893 (N_6893,N_5408,N_5068);
and U6894 (N_6894,N_5325,N_5362);
and U6895 (N_6895,N_5064,N_5155);
or U6896 (N_6896,N_5840,N_5687);
and U6897 (N_6897,N_5811,N_5207);
or U6898 (N_6898,N_5613,N_5017);
or U6899 (N_6899,N_5447,N_5903);
or U6900 (N_6900,N_5400,N_5972);
nand U6901 (N_6901,N_5739,N_5563);
nor U6902 (N_6902,N_5459,N_5918);
and U6903 (N_6903,N_5336,N_5454);
xnor U6904 (N_6904,N_5995,N_5304);
nand U6905 (N_6905,N_5751,N_5371);
nand U6906 (N_6906,N_5000,N_5821);
nor U6907 (N_6907,N_5249,N_5117);
xnor U6908 (N_6908,N_5691,N_5165);
nor U6909 (N_6909,N_5626,N_5482);
xor U6910 (N_6910,N_5803,N_5124);
or U6911 (N_6911,N_5928,N_5673);
or U6912 (N_6912,N_5983,N_5500);
or U6913 (N_6913,N_5221,N_5188);
xor U6914 (N_6914,N_5214,N_5138);
nand U6915 (N_6915,N_5026,N_5926);
xnor U6916 (N_6916,N_5962,N_5450);
nand U6917 (N_6917,N_5607,N_5274);
or U6918 (N_6918,N_5876,N_5776);
xor U6919 (N_6919,N_5150,N_5453);
and U6920 (N_6920,N_5880,N_5384);
xor U6921 (N_6921,N_5657,N_5384);
nor U6922 (N_6922,N_5848,N_5699);
and U6923 (N_6923,N_5794,N_5637);
xnor U6924 (N_6924,N_5257,N_5959);
xor U6925 (N_6925,N_5068,N_5719);
and U6926 (N_6926,N_5503,N_5435);
and U6927 (N_6927,N_5779,N_5532);
nor U6928 (N_6928,N_5752,N_5143);
xnor U6929 (N_6929,N_5098,N_5011);
xnor U6930 (N_6930,N_5119,N_5430);
xor U6931 (N_6931,N_5955,N_5484);
nor U6932 (N_6932,N_5808,N_5726);
nor U6933 (N_6933,N_5507,N_5398);
or U6934 (N_6934,N_5227,N_5002);
nor U6935 (N_6935,N_5256,N_5692);
nand U6936 (N_6936,N_5888,N_5847);
and U6937 (N_6937,N_5555,N_5591);
or U6938 (N_6938,N_5959,N_5486);
xor U6939 (N_6939,N_5834,N_5107);
or U6940 (N_6940,N_5512,N_5424);
nand U6941 (N_6941,N_5573,N_5741);
and U6942 (N_6942,N_5549,N_5158);
xor U6943 (N_6943,N_5345,N_5009);
xnor U6944 (N_6944,N_5248,N_5694);
nor U6945 (N_6945,N_5340,N_5055);
or U6946 (N_6946,N_5580,N_5083);
nand U6947 (N_6947,N_5741,N_5540);
and U6948 (N_6948,N_5233,N_5502);
or U6949 (N_6949,N_5644,N_5662);
and U6950 (N_6950,N_5192,N_5705);
nand U6951 (N_6951,N_5445,N_5779);
xnor U6952 (N_6952,N_5256,N_5445);
and U6953 (N_6953,N_5587,N_5348);
nor U6954 (N_6954,N_5588,N_5834);
nor U6955 (N_6955,N_5125,N_5481);
and U6956 (N_6956,N_5807,N_5830);
or U6957 (N_6957,N_5125,N_5573);
nand U6958 (N_6958,N_5751,N_5416);
or U6959 (N_6959,N_5209,N_5839);
or U6960 (N_6960,N_5060,N_5962);
and U6961 (N_6961,N_5845,N_5070);
and U6962 (N_6962,N_5061,N_5029);
and U6963 (N_6963,N_5248,N_5377);
nor U6964 (N_6964,N_5893,N_5183);
nor U6965 (N_6965,N_5712,N_5373);
nand U6966 (N_6966,N_5617,N_5388);
nand U6967 (N_6967,N_5076,N_5766);
xnor U6968 (N_6968,N_5691,N_5931);
nand U6969 (N_6969,N_5931,N_5483);
nor U6970 (N_6970,N_5835,N_5144);
nor U6971 (N_6971,N_5447,N_5397);
or U6972 (N_6972,N_5308,N_5162);
xnor U6973 (N_6973,N_5368,N_5331);
nand U6974 (N_6974,N_5179,N_5160);
nor U6975 (N_6975,N_5232,N_5311);
xnor U6976 (N_6976,N_5272,N_5954);
or U6977 (N_6977,N_5525,N_5588);
and U6978 (N_6978,N_5149,N_5261);
or U6979 (N_6979,N_5126,N_5704);
xnor U6980 (N_6980,N_5272,N_5058);
and U6981 (N_6981,N_5006,N_5011);
nand U6982 (N_6982,N_5695,N_5245);
nand U6983 (N_6983,N_5113,N_5569);
nand U6984 (N_6984,N_5759,N_5928);
or U6985 (N_6985,N_5667,N_5147);
and U6986 (N_6986,N_5025,N_5823);
xor U6987 (N_6987,N_5878,N_5514);
nand U6988 (N_6988,N_5027,N_5857);
nor U6989 (N_6989,N_5701,N_5933);
or U6990 (N_6990,N_5434,N_5304);
nor U6991 (N_6991,N_5018,N_5625);
and U6992 (N_6992,N_5576,N_5285);
and U6993 (N_6993,N_5758,N_5988);
and U6994 (N_6994,N_5208,N_5949);
and U6995 (N_6995,N_5542,N_5717);
or U6996 (N_6996,N_5592,N_5629);
nand U6997 (N_6997,N_5094,N_5166);
nor U6998 (N_6998,N_5911,N_5823);
and U6999 (N_6999,N_5222,N_5675);
or U7000 (N_7000,N_6625,N_6524);
or U7001 (N_7001,N_6035,N_6835);
nand U7002 (N_7002,N_6620,N_6659);
nand U7003 (N_7003,N_6675,N_6962);
or U7004 (N_7004,N_6742,N_6305);
or U7005 (N_7005,N_6853,N_6705);
nand U7006 (N_7006,N_6817,N_6345);
xor U7007 (N_7007,N_6757,N_6665);
nand U7008 (N_7008,N_6952,N_6315);
nor U7009 (N_7009,N_6358,N_6143);
xnor U7010 (N_7010,N_6619,N_6974);
or U7011 (N_7011,N_6445,N_6095);
xnor U7012 (N_7012,N_6046,N_6566);
nand U7013 (N_7013,N_6339,N_6890);
xor U7014 (N_7014,N_6282,N_6258);
xnor U7015 (N_7015,N_6654,N_6780);
and U7016 (N_7016,N_6068,N_6500);
xor U7017 (N_7017,N_6804,N_6114);
or U7018 (N_7018,N_6873,N_6082);
xnor U7019 (N_7019,N_6111,N_6145);
nand U7020 (N_7020,N_6755,N_6929);
nand U7021 (N_7021,N_6493,N_6264);
xor U7022 (N_7022,N_6970,N_6115);
xnor U7023 (N_7023,N_6181,N_6255);
or U7024 (N_7024,N_6470,N_6295);
or U7025 (N_7025,N_6256,N_6939);
and U7026 (N_7026,N_6628,N_6006);
and U7027 (N_7027,N_6541,N_6584);
nor U7028 (N_7028,N_6877,N_6026);
nor U7029 (N_7029,N_6013,N_6866);
nor U7030 (N_7030,N_6951,N_6465);
or U7031 (N_7031,N_6056,N_6100);
or U7032 (N_7032,N_6471,N_6474);
xnor U7033 (N_7033,N_6395,N_6996);
and U7034 (N_7034,N_6191,N_6435);
and U7035 (N_7035,N_6613,N_6271);
nand U7036 (N_7036,N_6463,N_6079);
xnor U7037 (N_7037,N_6257,N_6049);
and U7038 (N_7038,N_6723,N_6727);
xor U7039 (N_7039,N_6652,N_6765);
xnor U7040 (N_7040,N_6534,N_6883);
nor U7041 (N_7041,N_6270,N_6022);
xor U7042 (N_7042,N_6975,N_6531);
or U7043 (N_7043,N_6569,N_6643);
or U7044 (N_7044,N_6856,N_6074);
and U7045 (N_7045,N_6381,N_6807);
nand U7046 (N_7046,N_6629,N_6878);
xnor U7047 (N_7047,N_6405,N_6144);
xor U7048 (N_7048,N_6547,N_6546);
nand U7049 (N_7049,N_6741,N_6525);
nor U7050 (N_7050,N_6801,N_6104);
nor U7051 (N_7051,N_6651,N_6172);
and U7052 (N_7052,N_6568,N_6812);
or U7053 (N_7053,N_6598,N_6323);
nand U7054 (N_7054,N_6484,N_6863);
and U7055 (N_7055,N_6333,N_6288);
nand U7056 (N_7056,N_6960,N_6580);
xnor U7057 (N_7057,N_6707,N_6177);
and U7058 (N_7058,N_6131,N_6389);
nor U7059 (N_7059,N_6262,N_6815);
and U7060 (N_7060,N_6066,N_6123);
nand U7061 (N_7061,N_6422,N_6153);
and U7062 (N_7062,N_6609,N_6868);
xnor U7063 (N_7063,N_6062,N_6110);
nor U7064 (N_7064,N_6876,N_6036);
nor U7065 (N_7065,N_6229,N_6505);
xor U7066 (N_7066,N_6045,N_6926);
xor U7067 (N_7067,N_6591,N_6605);
or U7068 (N_7068,N_6922,N_6942);
and U7069 (N_7069,N_6735,N_6363);
nand U7070 (N_7070,N_6535,N_6284);
and U7071 (N_7071,N_6135,N_6134);
or U7072 (N_7072,N_6925,N_6479);
and U7073 (N_7073,N_6320,N_6290);
xor U7074 (N_7074,N_6176,N_6206);
nor U7075 (N_7075,N_6697,N_6461);
and U7076 (N_7076,N_6239,N_6915);
or U7077 (N_7077,N_6109,N_6771);
or U7078 (N_7078,N_6203,N_6120);
and U7079 (N_7079,N_6881,N_6453);
nor U7080 (N_7080,N_6517,N_6141);
nand U7081 (N_7081,N_6025,N_6767);
or U7082 (N_7082,N_6084,N_6164);
and U7083 (N_7083,N_6442,N_6934);
nand U7084 (N_7084,N_6720,N_6956);
and U7085 (N_7085,N_6979,N_6486);
or U7086 (N_7086,N_6336,N_6946);
or U7087 (N_7087,N_6857,N_6269);
nand U7088 (N_7088,N_6273,N_6051);
or U7089 (N_7089,N_6630,N_6984);
nor U7090 (N_7090,N_6018,N_6579);
or U7091 (N_7091,N_6912,N_6214);
nand U7092 (N_7092,N_6673,N_6538);
nand U7093 (N_7093,N_6379,N_6512);
nor U7094 (N_7094,N_6828,N_6642);
or U7095 (N_7095,N_6370,N_6210);
and U7096 (N_7096,N_6749,N_6808);
xnor U7097 (N_7097,N_6454,N_6017);
nor U7098 (N_7098,N_6884,N_6986);
or U7099 (N_7099,N_6513,N_6039);
and U7100 (N_7100,N_6748,N_6738);
nor U7101 (N_7101,N_6124,N_6614);
nand U7102 (N_7102,N_6932,N_6947);
nand U7103 (N_7103,N_6796,N_6390);
or U7104 (N_7104,N_6433,N_6162);
nand U7105 (N_7105,N_6964,N_6662);
xor U7106 (N_7106,N_6632,N_6849);
nor U7107 (N_7107,N_6001,N_6692);
nand U7108 (N_7108,N_6684,N_6216);
nand U7109 (N_7109,N_6014,N_6289);
and U7110 (N_7110,N_6187,N_6814);
nor U7111 (N_7111,N_6699,N_6155);
or U7112 (N_7112,N_6447,N_6657);
and U7113 (N_7113,N_6940,N_6369);
and U7114 (N_7114,N_6587,N_6848);
nand U7115 (N_7115,N_6448,N_6365);
nand U7116 (N_7116,N_6417,N_6610);
nor U7117 (N_7117,N_6054,N_6337);
xnor U7118 (N_7118,N_6838,N_6421);
xor U7119 (N_7119,N_6910,N_6069);
nor U7120 (N_7120,N_6174,N_6927);
xnor U7121 (N_7121,N_6166,N_6373);
and U7122 (N_7122,N_6411,N_6261);
or U7123 (N_7123,N_6416,N_6887);
and U7124 (N_7124,N_6567,N_6382);
xor U7125 (N_7125,N_6576,N_6016);
nand U7126 (N_7126,N_6059,N_6129);
or U7127 (N_7127,N_6754,N_6093);
nand U7128 (N_7128,N_6081,N_6639);
or U7129 (N_7129,N_6434,N_6317);
nand U7130 (N_7130,N_6800,N_6357);
nand U7131 (N_7131,N_6444,N_6329);
xor U7132 (N_7132,N_6297,N_6739);
xnor U7133 (N_7133,N_6980,N_6840);
or U7134 (N_7134,N_6543,N_6763);
nand U7135 (N_7135,N_6518,N_6238);
nor U7136 (N_7136,N_6497,N_6773);
xor U7137 (N_7137,N_6151,N_6918);
xor U7138 (N_7138,N_6420,N_6943);
nor U7139 (N_7139,N_6539,N_6170);
and U7140 (N_7140,N_6564,N_6717);
xnor U7141 (N_7141,N_6799,N_6752);
and U7142 (N_7142,N_6080,N_6136);
and U7143 (N_7143,N_6944,N_6190);
or U7144 (N_7144,N_6585,N_6087);
or U7145 (N_7145,N_6060,N_6899);
nand U7146 (N_7146,N_6184,N_6839);
xor U7147 (N_7147,N_6169,N_6274);
or U7148 (N_7148,N_6552,N_6489);
nor U7149 (N_7149,N_6803,N_6075);
xor U7150 (N_7150,N_6595,N_6307);
nor U7151 (N_7151,N_6981,N_6052);
xnor U7152 (N_7152,N_6142,N_6237);
nor U7153 (N_7153,N_6427,N_6233);
and U7154 (N_7154,N_6885,N_6851);
and U7155 (N_7155,N_6232,N_6355);
nand U7156 (N_7156,N_6199,N_6354);
nor U7157 (N_7157,N_6293,N_6419);
nor U7158 (N_7158,N_6235,N_6396);
xor U7159 (N_7159,N_6350,N_6408);
and U7160 (N_7160,N_6965,N_6321);
nor U7161 (N_7161,N_6043,N_6053);
nor U7162 (N_7162,N_6725,N_6924);
xnor U7163 (N_7163,N_6356,N_6055);
xnor U7164 (N_7164,N_6963,N_6935);
nand U7165 (N_7165,N_6615,N_6196);
or U7166 (N_7166,N_6776,N_6178);
xnor U7167 (N_7167,N_6253,N_6572);
xnor U7168 (N_7168,N_6532,N_6030);
and U7169 (N_7169,N_6248,N_6275);
and U7170 (N_7170,N_6607,N_6446);
nand U7171 (N_7171,N_6303,N_6718);
nor U7172 (N_7172,N_6548,N_6971);
nand U7173 (N_7173,N_6976,N_6666);
nor U7174 (N_7174,N_6360,N_6917);
xnor U7175 (N_7175,N_6452,N_6252);
or U7176 (N_7176,N_6677,N_6770);
and U7177 (N_7177,N_6823,N_6793);
nor U7178 (N_7178,N_6914,N_6653);
and U7179 (N_7179,N_6475,N_6913);
nor U7180 (N_7180,N_6700,N_6246);
or U7181 (N_7181,N_6186,N_6743);
nor U7182 (N_7182,N_6509,N_6714);
and U7183 (N_7183,N_6327,N_6234);
and U7184 (N_7184,N_6772,N_6762);
nand U7185 (N_7185,N_6343,N_6788);
nor U7186 (N_7186,N_6734,N_6460);
nand U7187 (N_7187,N_6729,N_6462);
nor U7188 (N_7188,N_6318,N_6496);
xnor U7189 (N_7189,N_6312,N_6311);
xnor U7190 (N_7190,N_6894,N_6280);
and U7191 (N_7191,N_6820,N_6761);
nand U7192 (N_7192,N_6845,N_6331);
xnor U7193 (N_7193,N_6418,N_6528);
nand U7194 (N_7194,N_6310,N_6693);
and U7195 (N_7195,N_6414,N_6031);
nor U7196 (N_7196,N_6994,N_6871);
xnor U7197 (N_7197,N_6067,N_6027);
and U7198 (N_7198,N_6266,N_6362);
xor U7199 (N_7199,N_6634,N_6933);
nand U7200 (N_7200,N_6160,N_6314);
and U7201 (N_7201,N_6867,N_6818);
nor U7202 (N_7202,N_6483,N_6608);
nand U7203 (N_7203,N_6244,N_6973);
nor U7204 (N_7204,N_6374,N_6415);
and U7205 (N_7205,N_6854,N_6148);
nor U7206 (N_7206,N_6254,N_6167);
and U7207 (N_7207,N_6106,N_6565);
xnor U7208 (N_7208,N_6626,N_6602);
nand U7209 (N_7209,N_6477,N_6459);
and U7210 (N_7210,N_6431,N_6575);
xor U7211 (N_7211,N_6002,N_6751);
nand U7212 (N_7212,N_6152,N_6750);
nor U7213 (N_7213,N_6805,N_6536);
and U7214 (N_7214,N_6102,N_6746);
and U7215 (N_7215,N_6968,N_6126);
or U7216 (N_7216,N_6703,N_6071);
nor U7217 (N_7217,N_6737,N_6954);
and U7218 (N_7218,N_6989,N_6473);
or U7219 (N_7219,N_6590,N_6300);
or U7220 (N_7220,N_6826,N_6798);
xnor U7221 (N_7221,N_6432,N_6861);
and U7222 (N_7222,N_6923,N_6830);
xnor U7223 (N_7223,N_6180,N_6384);
xnor U7224 (N_7224,N_6810,N_6819);
or U7225 (N_7225,N_6132,N_6545);
xor U7226 (N_7226,N_6637,N_6335);
or U7227 (N_7227,N_6011,N_6292);
nand U7228 (N_7228,N_6032,N_6636);
or U7229 (N_7229,N_6685,N_6201);
nor U7230 (N_7230,N_6574,N_6519);
nand U7231 (N_7231,N_6426,N_6501);
and U7232 (N_7232,N_6249,N_6641);
or U7233 (N_7233,N_6193,N_6090);
or U7234 (N_7234,N_6958,N_6859);
and U7235 (N_7235,N_6691,N_6516);
nand U7236 (N_7236,N_6900,N_6862);
nand U7237 (N_7237,N_6351,N_6676);
nor U7238 (N_7238,N_6514,N_6251);
or U7239 (N_7239,N_6400,N_6596);
or U7240 (N_7240,N_6661,N_6385);
xnor U7241 (N_7241,N_6230,N_6078);
or U7242 (N_7242,N_6044,N_6306);
and U7243 (N_7243,N_6101,N_6359);
nor U7244 (N_7244,N_6842,N_6557);
xor U7245 (N_7245,N_6756,N_6977);
nor U7246 (N_7246,N_6852,N_6347);
and U7247 (N_7247,N_6554,N_6860);
nor U7248 (N_7248,N_6711,N_6037);
or U7249 (N_7249,N_6481,N_6349);
or U7250 (N_7250,N_6399,N_6119);
nand U7251 (N_7251,N_6740,N_6386);
xnor U7252 (N_7252,N_6578,N_6904);
xnor U7253 (N_7253,N_6834,N_6809);
and U7254 (N_7254,N_6726,N_6897);
and U7255 (N_7255,N_6905,N_6077);
and U7256 (N_7256,N_6133,N_6466);
nand U7257 (N_7257,N_6209,N_6222);
nor U7258 (N_7258,N_6589,N_6437);
nand U7259 (N_7259,N_6594,N_6383);
xor U7260 (N_7260,N_6212,N_6482);
nor U7261 (N_7261,N_6103,N_6844);
or U7262 (N_7262,N_6781,N_6736);
and U7263 (N_7263,N_6361,N_6831);
nor U7264 (N_7264,N_6806,N_6301);
xor U7265 (N_7265,N_6858,N_6791);
nand U7266 (N_7266,N_6438,N_6122);
nand U7267 (N_7267,N_6945,N_6789);
or U7268 (N_7268,N_6019,N_6021);
nor U7269 (N_7269,N_6091,N_6458);
nand U7270 (N_7270,N_6635,N_6154);
or U7271 (N_7271,N_6616,N_6268);
or U7272 (N_7272,N_6003,N_6058);
nor U7273 (N_7273,N_6029,N_6367);
xnor U7274 (N_7274,N_6753,N_6227);
and U7275 (N_7275,N_6494,N_6825);
nor U7276 (N_7276,N_6072,N_6423);
xor U7277 (N_7277,N_6701,N_6577);
xor U7278 (N_7278,N_6468,N_6498);
nor U7279 (N_7279,N_6766,N_6888);
and U7280 (N_7280,N_6436,N_6183);
and U7281 (N_7281,N_6224,N_6338);
or U7282 (N_7282,N_6603,N_6950);
and U7283 (N_7283,N_6380,N_6560);
nand U7284 (N_7284,N_6715,N_6724);
xnor U7285 (N_7285,N_6679,N_6957);
or U7286 (N_7286,N_6217,N_6606);
nor U7287 (N_7287,N_6961,N_6646);
or U7288 (N_7288,N_6198,N_6621);
xor U7289 (N_7289,N_6397,N_6540);
and U7290 (N_7290,N_6682,N_6503);
and U7291 (N_7291,N_6938,N_6833);
or U7292 (N_7292,N_6687,N_6330);
and U7293 (N_7293,N_6065,N_6245);
xor U7294 (N_7294,N_6695,N_6604);
nor U7295 (N_7295,N_6112,N_6732);
xor U7296 (N_7296,N_6401,N_6664);
xnor U7297 (N_7297,N_6864,N_6992);
and U7298 (N_7298,N_6378,N_6782);
or U7299 (N_7299,N_6777,N_6197);
xnor U7300 (N_7300,N_6722,N_6207);
nor U7301 (N_7301,N_6012,N_6640);
nand U7302 (N_7302,N_6972,N_6127);
or U7303 (N_7303,N_6645,N_6393);
and U7304 (N_7304,N_6869,N_6319);
or U7305 (N_7305,N_6507,N_6571);
xor U7306 (N_7306,N_6403,N_6404);
nand U7307 (N_7307,N_6702,N_6332);
nand U7308 (N_7308,N_6520,N_6712);
nor U7309 (N_7309,N_6556,N_6076);
and U7310 (N_7310,N_6672,N_6392);
or U7311 (N_7311,N_6202,N_6523);
nor U7312 (N_7312,N_6694,N_6121);
nor U7313 (N_7313,N_6582,N_6930);
xnor U7314 (N_7314,N_6138,N_6147);
nor U7315 (N_7315,N_6424,N_6953);
nand U7316 (N_7316,N_6730,N_6240);
xor U7317 (N_7317,N_6982,N_6627);
or U7318 (N_7318,N_6009,N_6158);
nor U7319 (N_7319,N_6710,N_6522);
nand U7320 (N_7320,N_6430,N_6099);
xnor U7321 (N_7321,N_6061,N_6034);
or U7322 (N_7322,N_6267,N_6488);
nand U7323 (N_7323,N_6792,N_6125);
nor U7324 (N_7324,N_6822,N_6936);
and U7325 (N_7325,N_6218,N_6324);
nor U7326 (N_7326,N_6683,N_6787);
xor U7327 (N_7327,N_6891,N_6991);
xnor U7328 (N_7328,N_6504,N_6117);
xnor U7329 (N_7329,N_6279,N_6412);
nand U7330 (N_7330,N_6921,N_6200);
xnor U7331 (N_7331,N_6993,N_6092);
or U7332 (N_7332,N_6213,N_6220);
or U7333 (N_7333,N_6149,N_6583);
nand U7334 (N_7334,N_6816,N_6308);
and U7335 (N_7335,N_6686,N_6478);
and U7336 (N_7336,N_6708,N_6449);
nor U7337 (N_7337,N_6189,N_6005);
and U7338 (N_7338,N_6719,N_6173);
and U7339 (N_7339,N_6491,N_6850);
nor U7340 (N_7340,N_6259,N_6786);
nand U7341 (N_7341,N_6283,N_6802);
nor U7342 (N_7342,N_6004,N_6247);
nand U7343 (N_7343,N_6794,N_6228);
and U7344 (N_7344,N_6502,N_6836);
nand U7345 (N_7345,N_6492,N_6024);
or U7346 (N_7346,N_6413,N_6304);
nor U7347 (N_7347,N_6456,N_6529);
or U7348 (N_7348,N_6085,N_6108);
nor U7349 (N_7349,N_6678,N_6185);
xor U7350 (N_7350,N_6428,N_6041);
nand U7351 (N_7351,N_6882,N_6558);
xnor U7352 (N_7352,N_6829,N_6778);
and U7353 (N_7353,N_6033,N_6241);
and U7354 (N_7354,N_6759,N_6376);
and U7355 (N_7355,N_6113,N_6118);
nand U7356 (N_7356,N_6624,N_6916);
nand U7357 (N_7357,N_6020,N_6731);
nand U7358 (N_7358,N_6325,N_6690);
nor U7359 (N_7359,N_6983,N_6713);
and U7360 (N_7360,N_6163,N_6451);
xor U7361 (N_7361,N_6000,N_6334);
or U7362 (N_7362,N_6941,N_6889);
and U7363 (N_7363,N_6784,N_6480);
or U7364 (N_7364,N_6611,N_6893);
and U7365 (N_7365,N_6843,N_6250);
or U7366 (N_7366,N_6219,N_6073);
xnor U7367 (N_7367,N_6455,N_6137);
nand U7368 (N_7368,N_6597,N_6188);
or U7369 (N_7369,N_6783,N_6865);
xor U7370 (N_7370,N_6660,N_6495);
or U7371 (N_7371,N_6667,N_6116);
xnor U7372 (N_7372,N_6105,N_6588);
nor U7373 (N_7373,N_6140,N_6168);
nor U7374 (N_7374,N_6511,N_6995);
and U7375 (N_7375,N_6847,N_6559);
or U7376 (N_7376,N_6561,N_6903);
and U7377 (N_7377,N_6902,N_6182);
or U7378 (N_7378,N_6985,N_6716);
nand U7379 (N_7379,N_6394,N_6837);
xor U7380 (N_7380,N_6161,N_6895);
nand U7381 (N_7381,N_6827,N_6909);
or U7382 (N_7382,N_6341,N_6128);
nor U7383 (N_7383,N_6409,N_6706);
and U7384 (N_7384,N_6194,N_6928);
and U7385 (N_7385,N_6506,N_6875);
and U7386 (N_7386,N_6439,N_6328);
nand U7387 (N_7387,N_6959,N_6457);
xor U7388 (N_7388,N_6824,N_6008);
or U7389 (N_7389,N_6467,N_6352);
or U7390 (N_7390,N_6955,N_6709);
nand U7391 (N_7391,N_6375,N_6515);
nand U7392 (N_7392,N_6286,N_6299);
and U7393 (N_7393,N_6083,N_6047);
and U7394 (N_7394,N_6285,N_6195);
nand U7395 (N_7395,N_6015,N_6728);
nor U7396 (N_7396,N_6570,N_6669);
and U7397 (N_7397,N_6366,N_6906);
or U7398 (N_7398,N_6464,N_6485);
nor U7399 (N_7399,N_6919,N_6745);
nand U7400 (N_7400,N_6038,N_6130);
nand U7401 (N_7401,N_6171,N_6521);
nor U7402 (N_7402,N_6175,N_6760);
or U7403 (N_7403,N_6931,N_6680);
xor U7404 (N_7404,N_6967,N_6050);
and U7405 (N_7405,N_6581,N_6322);
nand U7406 (N_7406,N_6348,N_6880);
or U7407 (N_7407,N_6042,N_6872);
or U7408 (N_7408,N_6907,N_6098);
or U7409 (N_7409,N_6159,N_6948);
xor U7410 (N_7410,N_6698,N_6832);
or U7411 (N_7411,N_6088,N_6165);
or U7412 (N_7412,N_6920,N_6593);
nor U7413 (N_7413,N_6443,N_6276);
or U7414 (N_7414,N_6785,N_6874);
or U7415 (N_7415,N_6998,N_6377);
xnor U7416 (N_7416,N_6987,N_6551);
or U7417 (N_7417,N_6287,N_6094);
and U7418 (N_7418,N_6744,N_6544);
nand U7419 (N_7419,N_6663,N_6097);
and U7420 (N_7420,N_6302,N_6990);
nor U7421 (N_7421,N_6215,N_6550);
nand U7422 (N_7422,N_6096,N_6908);
nor U7423 (N_7423,N_6139,N_6542);
nor U7424 (N_7424,N_6674,N_6221);
xor U7425 (N_7425,N_6064,N_6313);
xor U7426 (N_7426,N_6562,N_6797);
nor U7427 (N_7427,N_6278,N_6549);
nor U7428 (N_7428,N_6721,N_6107);
xnor U7429 (N_7429,N_6696,N_6655);
nand U7430 (N_7430,N_6368,N_6656);
or U7431 (N_7431,N_6670,N_6425);
and U7432 (N_7432,N_6225,N_6911);
nor U7433 (N_7433,N_6537,N_6398);
nand U7434 (N_7434,N_6638,N_6242);
nand U7435 (N_7435,N_6841,N_6526);
nor U7436 (N_7436,N_6999,N_6353);
or U7437 (N_7437,N_6855,N_6949);
or U7438 (N_7438,N_6371,N_6402);
nor U7439 (N_7439,N_6648,N_6344);
nor U7440 (N_7440,N_6407,N_6192);
xnor U7441 (N_7441,N_6530,N_6688);
and U7442 (N_7442,N_6758,N_6294);
nand U7443 (N_7443,N_6527,N_6440);
or U7444 (N_7444,N_6966,N_6689);
or U7445 (N_7445,N_6291,N_6450);
nand U7446 (N_7446,N_6764,N_6790);
or U7447 (N_7447,N_6372,N_6775);
nand U7448 (N_7448,N_6063,N_6340);
xnor U7449 (N_7449,N_6007,N_6671);
nor U7450 (N_7450,N_6410,N_6316);
nor U7451 (N_7451,N_6179,N_6487);
and U7452 (N_7452,N_6057,N_6040);
nand U7453 (N_7453,N_6901,N_6892);
xnor U7454 (N_7454,N_6988,N_6631);
nor U7455 (N_7455,N_6846,N_6272);
xor U7456 (N_7456,N_6644,N_6070);
xnor U7457 (N_7457,N_6555,N_6429);
xor U7458 (N_7458,N_6342,N_6647);
or U7459 (N_7459,N_6622,N_6668);
nor U7460 (N_7460,N_6811,N_6813);
or U7461 (N_7461,N_6086,N_6795);
nand U7462 (N_7462,N_6612,N_6769);
nor U7463 (N_7463,N_6150,N_6969);
xnor U7464 (N_7464,N_6633,N_6553);
xnor U7465 (N_7465,N_6649,N_6472);
nor U7466 (N_7466,N_6260,N_6243);
and U7467 (N_7467,N_6231,N_6978);
and U7468 (N_7468,N_6733,N_6156);
or U7469 (N_7469,N_6208,N_6157);
or U7470 (N_7470,N_6028,N_6508);
nand U7471 (N_7471,N_6277,N_6623);
or U7472 (N_7472,N_6469,N_6618);
nor U7473 (N_7473,N_6586,N_6896);
xnor U7474 (N_7474,N_6886,N_6265);
xnor U7475 (N_7475,N_6747,N_6779);
and U7476 (N_7476,N_6010,N_6499);
nor U7477 (N_7477,N_6600,N_6821);
and U7478 (N_7478,N_6599,N_6298);
or U7479 (N_7479,N_6309,N_6211);
xnor U7480 (N_7480,N_6387,N_6898);
and U7481 (N_7481,N_6205,N_6681);
and U7482 (N_7482,N_6997,N_6204);
nor U7483 (N_7483,N_6510,N_6768);
and U7484 (N_7484,N_6563,N_6870);
nor U7485 (N_7485,N_6223,N_6226);
nor U7486 (N_7486,N_6774,N_6592);
nor U7487 (N_7487,N_6490,N_6658);
and U7488 (N_7488,N_6089,N_6406);
nor U7489 (N_7489,N_6573,N_6263);
or U7490 (N_7490,N_6346,N_6146);
or U7491 (N_7491,N_6879,N_6441);
xnor U7492 (N_7492,N_6023,N_6281);
nor U7493 (N_7493,N_6704,N_6048);
and U7494 (N_7494,N_6326,N_6236);
and U7495 (N_7495,N_6601,N_6533);
and U7496 (N_7496,N_6391,N_6476);
nand U7497 (N_7497,N_6388,N_6650);
nor U7498 (N_7498,N_6617,N_6296);
nor U7499 (N_7499,N_6364,N_6937);
nand U7500 (N_7500,N_6153,N_6497);
and U7501 (N_7501,N_6706,N_6107);
or U7502 (N_7502,N_6612,N_6005);
nand U7503 (N_7503,N_6064,N_6082);
xnor U7504 (N_7504,N_6816,N_6386);
or U7505 (N_7505,N_6300,N_6545);
xnor U7506 (N_7506,N_6142,N_6015);
and U7507 (N_7507,N_6440,N_6293);
nand U7508 (N_7508,N_6643,N_6046);
or U7509 (N_7509,N_6835,N_6060);
and U7510 (N_7510,N_6576,N_6875);
xor U7511 (N_7511,N_6254,N_6507);
and U7512 (N_7512,N_6289,N_6898);
and U7513 (N_7513,N_6936,N_6103);
or U7514 (N_7514,N_6385,N_6605);
and U7515 (N_7515,N_6349,N_6637);
and U7516 (N_7516,N_6300,N_6481);
and U7517 (N_7517,N_6341,N_6718);
xnor U7518 (N_7518,N_6655,N_6725);
and U7519 (N_7519,N_6943,N_6509);
nor U7520 (N_7520,N_6269,N_6852);
and U7521 (N_7521,N_6994,N_6082);
xnor U7522 (N_7522,N_6133,N_6938);
nor U7523 (N_7523,N_6695,N_6981);
nand U7524 (N_7524,N_6154,N_6145);
and U7525 (N_7525,N_6900,N_6391);
xnor U7526 (N_7526,N_6484,N_6489);
nand U7527 (N_7527,N_6213,N_6310);
nand U7528 (N_7528,N_6911,N_6564);
or U7529 (N_7529,N_6271,N_6052);
or U7530 (N_7530,N_6643,N_6368);
nand U7531 (N_7531,N_6567,N_6262);
nor U7532 (N_7532,N_6122,N_6784);
and U7533 (N_7533,N_6225,N_6781);
or U7534 (N_7534,N_6553,N_6724);
and U7535 (N_7535,N_6462,N_6469);
or U7536 (N_7536,N_6321,N_6796);
or U7537 (N_7537,N_6610,N_6794);
xor U7538 (N_7538,N_6263,N_6253);
and U7539 (N_7539,N_6107,N_6693);
and U7540 (N_7540,N_6381,N_6986);
nand U7541 (N_7541,N_6206,N_6366);
nor U7542 (N_7542,N_6328,N_6694);
or U7543 (N_7543,N_6338,N_6986);
nor U7544 (N_7544,N_6204,N_6830);
nand U7545 (N_7545,N_6940,N_6988);
nand U7546 (N_7546,N_6156,N_6794);
or U7547 (N_7547,N_6743,N_6823);
nand U7548 (N_7548,N_6974,N_6024);
or U7549 (N_7549,N_6865,N_6819);
nor U7550 (N_7550,N_6619,N_6489);
and U7551 (N_7551,N_6296,N_6960);
nand U7552 (N_7552,N_6085,N_6632);
xor U7553 (N_7553,N_6667,N_6573);
nor U7554 (N_7554,N_6594,N_6084);
nor U7555 (N_7555,N_6436,N_6338);
nand U7556 (N_7556,N_6135,N_6410);
nor U7557 (N_7557,N_6632,N_6998);
nor U7558 (N_7558,N_6323,N_6534);
nor U7559 (N_7559,N_6913,N_6999);
nor U7560 (N_7560,N_6203,N_6887);
nand U7561 (N_7561,N_6194,N_6434);
nand U7562 (N_7562,N_6432,N_6021);
and U7563 (N_7563,N_6324,N_6812);
or U7564 (N_7564,N_6421,N_6207);
nor U7565 (N_7565,N_6787,N_6514);
nand U7566 (N_7566,N_6157,N_6724);
nand U7567 (N_7567,N_6223,N_6867);
xor U7568 (N_7568,N_6971,N_6643);
xor U7569 (N_7569,N_6572,N_6359);
nor U7570 (N_7570,N_6461,N_6531);
or U7571 (N_7571,N_6050,N_6697);
or U7572 (N_7572,N_6210,N_6102);
or U7573 (N_7573,N_6399,N_6029);
or U7574 (N_7574,N_6904,N_6941);
and U7575 (N_7575,N_6189,N_6986);
and U7576 (N_7576,N_6123,N_6801);
or U7577 (N_7577,N_6667,N_6953);
nor U7578 (N_7578,N_6020,N_6062);
nand U7579 (N_7579,N_6137,N_6402);
nand U7580 (N_7580,N_6420,N_6210);
nand U7581 (N_7581,N_6209,N_6165);
nand U7582 (N_7582,N_6449,N_6548);
and U7583 (N_7583,N_6900,N_6880);
and U7584 (N_7584,N_6101,N_6659);
and U7585 (N_7585,N_6650,N_6599);
and U7586 (N_7586,N_6283,N_6813);
xnor U7587 (N_7587,N_6539,N_6615);
xor U7588 (N_7588,N_6157,N_6005);
or U7589 (N_7589,N_6347,N_6376);
and U7590 (N_7590,N_6219,N_6258);
xor U7591 (N_7591,N_6263,N_6984);
and U7592 (N_7592,N_6737,N_6869);
and U7593 (N_7593,N_6151,N_6114);
or U7594 (N_7594,N_6175,N_6484);
xnor U7595 (N_7595,N_6320,N_6298);
nor U7596 (N_7596,N_6639,N_6133);
nor U7597 (N_7597,N_6731,N_6039);
nand U7598 (N_7598,N_6921,N_6013);
nand U7599 (N_7599,N_6500,N_6072);
nand U7600 (N_7600,N_6282,N_6578);
nor U7601 (N_7601,N_6230,N_6139);
and U7602 (N_7602,N_6125,N_6086);
nor U7603 (N_7603,N_6145,N_6810);
xor U7604 (N_7604,N_6785,N_6727);
xor U7605 (N_7605,N_6864,N_6695);
nor U7606 (N_7606,N_6000,N_6714);
nor U7607 (N_7607,N_6580,N_6230);
nand U7608 (N_7608,N_6982,N_6086);
xor U7609 (N_7609,N_6757,N_6192);
nand U7610 (N_7610,N_6957,N_6777);
nand U7611 (N_7611,N_6579,N_6319);
xnor U7612 (N_7612,N_6205,N_6136);
xnor U7613 (N_7613,N_6478,N_6687);
nand U7614 (N_7614,N_6589,N_6766);
and U7615 (N_7615,N_6228,N_6098);
xnor U7616 (N_7616,N_6916,N_6351);
or U7617 (N_7617,N_6421,N_6291);
nand U7618 (N_7618,N_6161,N_6823);
or U7619 (N_7619,N_6934,N_6350);
xnor U7620 (N_7620,N_6575,N_6372);
nor U7621 (N_7621,N_6789,N_6577);
and U7622 (N_7622,N_6671,N_6010);
or U7623 (N_7623,N_6930,N_6274);
and U7624 (N_7624,N_6420,N_6290);
nand U7625 (N_7625,N_6232,N_6018);
and U7626 (N_7626,N_6624,N_6128);
xnor U7627 (N_7627,N_6994,N_6124);
xor U7628 (N_7628,N_6791,N_6933);
nor U7629 (N_7629,N_6999,N_6323);
and U7630 (N_7630,N_6059,N_6120);
xnor U7631 (N_7631,N_6853,N_6330);
or U7632 (N_7632,N_6591,N_6733);
xnor U7633 (N_7633,N_6915,N_6575);
nor U7634 (N_7634,N_6961,N_6901);
or U7635 (N_7635,N_6599,N_6505);
or U7636 (N_7636,N_6108,N_6933);
nor U7637 (N_7637,N_6843,N_6278);
xnor U7638 (N_7638,N_6027,N_6776);
xnor U7639 (N_7639,N_6757,N_6203);
nor U7640 (N_7640,N_6075,N_6066);
nor U7641 (N_7641,N_6415,N_6070);
nor U7642 (N_7642,N_6694,N_6717);
nand U7643 (N_7643,N_6929,N_6253);
nor U7644 (N_7644,N_6539,N_6215);
nand U7645 (N_7645,N_6773,N_6096);
or U7646 (N_7646,N_6940,N_6944);
or U7647 (N_7647,N_6265,N_6101);
and U7648 (N_7648,N_6358,N_6191);
or U7649 (N_7649,N_6380,N_6931);
or U7650 (N_7650,N_6877,N_6630);
nand U7651 (N_7651,N_6920,N_6894);
nand U7652 (N_7652,N_6032,N_6570);
xnor U7653 (N_7653,N_6038,N_6804);
or U7654 (N_7654,N_6180,N_6804);
xor U7655 (N_7655,N_6480,N_6036);
nand U7656 (N_7656,N_6016,N_6126);
and U7657 (N_7657,N_6744,N_6022);
or U7658 (N_7658,N_6742,N_6476);
and U7659 (N_7659,N_6798,N_6869);
or U7660 (N_7660,N_6638,N_6212);
nor U7661 (N_7661,N_6464,N_6647);
xnor U7662 (N_7662,N_6679,N_6572);
and U7663 (N_7663,N_6264,N_6354);
or U7664 (N_7664,N_6748,N_6374);
or U7665 (N_7665,N_6284,N_6634);
nor U7666 (N_7666,N_6795,N_6028);
nand U7667 (N_7667,N_6357,N_6339);
nor U7668 (N_7668,N_6961,N_6482);
nand U7669 (N_7669,N_6835,N_6919);
nor U7670 (N_7670,N_6163,N_6524);
and U7671 (N_7671,N_6930,N_6999);
nand U7672 (N_7672,N_6134,N_6754);
or U7673 (N_7673,N_6043,N_6566);
and U7674 (N_7674,N_6992,N_6340);
and U7675 (N_7675,N_6776,N_6741);
or U7676 (N_7676,N_6363,N_6189);
nand U7677 (N_7677,N_6862,N_6521);
nor U7678 (N_7678,N_6841,N_6756);
nor U7679 (N_7679,N_6499,N_6290);
and U7680 (N_7680,N_6250,N_6904);
nand U7681 (N_7681,N_6638,N_6769);
nor U7682 (N_7682,N_6061,N_6314);
nand U7683 (N_7683,N_6392,N_6629);
or U7684 (N_7684,N_6603,N_6666);
nor U7685 (N_7685,N_6372,N_6121);
and U7686 (N_7686,N_6786,N_6468);
and U7687 (N_7687,N_6217,N_6968);
or U7688 (N_7688,N_6147,N_6861);
and U7689 (N_7689,N_6335,N_6470);
or U7690 (N_7690,N_6519,N_6424);
and U7691 (N_7691,N_6747,N_6729);
and U7692 (N_7692,N_6234,N_6712);
and U7693 (N_7693,N_6397,N_6630);
and U7694 (N_7694,N_6296,N_6429);
nor U7695 (N_7695,N_6295,N_6993);
and U7696 (N_7696,N_6544,N_6384);
or U7697 (N_7697,N_6210,N_6374);
nand U7698 (N_7698,N_6984,N_6051);
or U7699 (N_7699,N_6229,N_6414);
nand U7700 (N_7700,N_6445,N_6400);
and U7701 (N_7701,N_6010,N_6066);
xor U7702 (N_7702,N_6556,N_6725);
and U7703 (N_7703,N_6308,N_6482);
and U7704 (N_7704,N_6936,N_6421);
xor U7705 (N_7705,N_6364,N_6404);
nor U7706 (N_7706,N_6345,N_6472);
xnor U7707 (N_7707,N_6881,N_6634);
xor U7708 (N_7708,N_6514,N_6134);
xnor U7709 (N_7709,N_6441,N_6657);
xor U7710 (N_7710,N_6308,N_6999);
and U7711 (N_7711,N_6182,N_6352);
and U7712 (N_7712,N_6087,N_6565);
nand U7713 (N_7713,N_6980,N_6930);
nor U7714 (N_7714,N_6495,N_6173);
or U7715 (N_7715,N_6968,N_6111);
nor U7716 (N_7716,N_6879,N_6351);
nand U7717 (N_7717,N_6873,N_6876);
and U7718 (N_7718,N_6859,N_6339);
and U7719 (N_7719,N_6966,N_6465);
xor U7720 (N_7720,N_6118,N_6461);
nor U7721 (N_7721,N_6319,N_6671);
nand U7722 (N_7722,N_6181,N_6410);
and U7723 (N_7723,N_6212,N_6437);
and U7724 (N_7724,N_6995,N_6994);
or U7725 (N_7725,N_6314,N_6319);
xor U7726 (N_7726,N_6295,N_6972);
and U7727 (N_7727,N_6133,N_6559);
nor U7728 (N_7728,N_6049,N_6006);
and U7729 (N_7729,N_6524,N_6271);
nor U7730 (N_7730,N_6036,N_6559);
and U7731 (N_7731,N_6156,N_6267);
or U7732 (N_7732,N_6196,N_6176);
xnor U7733 (N_7733,N_6293,N_6627);
xor U7734 (N_7734,N_6273,N_6964);
nor U7735 (N_7735,N_6450,N_6434);
xnor U7736 (N_7736,N_6452,N_6767);
and U7737 (N_7737,N_6126,N_6319);
nand U7738 (N_7738,N_6110,N_6647);
nor U7739 (N_7739,N_6440,N_6836);
xor U7740 (N_7740,N_6580,N_6220);
or U7741 (N_7741,N_6710,N_6345);
nand U7742 (N_7742,N_6571,N_6691);
or U7743 (N_7743,N_6125,N_6666);
and U7744 (N_7744,N_6352,N_6258);
nand U7745 (N_7745,N_6106,N_6060);
xnor U7746 (N_7746,N_6935,N_6186);
and U7747 (N_7747,N_6326,N_6105);
and U7748 (N_7748,N_6940,N_6344);
and U7749 (N_7749,N_6361,N_6658);
nor U7750 (N_7750,N_6743,N_6436);
nor U7751 (N_7751,N_6105,N_6202);
nand U7752 (N_7752,N_6418,N_6604);
and U7753 (N_7753,N_6949,N_6026);
nor U7754 (N_7754,N_6404,N_6323);
xnor U7755 (N_7755,N_6503,N_6987);
or U7756 (N_7756,N_6763,N_6116);
or U7757 (N_7757,N_6590,N_6351);
and U7758 (N_7758,N_6598,N_6666);
and U7759 (N_7759,N_6932,N_6210);
nor U7760 (N_7760,N_6906,N_6516);
and U7761 (N_7761,N_6464,N_6065);
or U7762 (N_7762,N_6914,N_6860);
nor U7763 (N_7763,N_6080,N_6526);
and U7764 (N_7764,N_6516,N_6324);
nor U7765 (N_7765,N_6969,N_6073);
and U7766 (N_7766,N_6391,N_6012);
and U7767 (N_7767,N_6127,N_6306);
xnor U7768 (N_7768,N_6400,N_6204);
xnor U7769 (N_7769,N_6113,N_6184);
or U7770 (N_7770,N_6607,N_6424);
xnor U7771 (N_7771,N_6058,N_6228);
nand U7772 (N_7772,N_6021,N_6453);
nand U7773 (N_7773,N_6886,N_6302);
xnor U7774 (N_7774,N_6885,N_6419);
or U7775 (N_7775,N_6812,N_6625);
xnor U7776 (N_7776,N_6016,N_6307);
and U7777 (N_7777,N_6519,N_6196);
xnor U7778 (N_7778,N_6224,N_6435);
and U7779 (N_7779,N_6691,N_6290);
xnor U7780 (N_7780,N_6645,N_6896);
xor U7781 (N_7781,N_6031,N_6586);
nor U7782 (N_7782,N_6942,N_6027);
xnor U7783 (N_7783,N_6837,N_6228);
nor U7784 (N_7784,N_6384,N_6949);
and U7785 (N_7785,N_6298,N_6110);
nor U7786 (N_7786,N_6560,N_6809);
or U7787 (N_7787,N_6052,N_6756);
and U7788 (N_7788,N_6926,N_6180);
or U7789 (N_7789,N_6948,N_6727);
nor U7790 (N_7790,N_6311,N_6287);
or U7791 (N_7791,N_6582,N_6783);
or U7792 (N_7792,N_6819,N_6708);
xor U7793 (N_7793,N_6047,N_6812);
nand U7794 (N_7794,N_6153,N_6165);
or U7795 (N_7795,N_6547,N_6494);
nor U7796 (N_7796,N_6495,N_6234);
and U7797 (N_7797,N_6793,N_6618);
and U7798 (N_7798,N_6255,N_6842);
xnor U7799 (N_7799,N_6161,N_6805);
nand U7800 (N_7800,N_6950,N_6639);
and U7801 (N_7801,N_6357,N_6108);
nor U7802 (N_7802,N_6230,N_6000);
xnor U7803 (N_7803,N_6465,N_6942);
and U7804 (N_7804,N_6821,N_6921);
nor U7805 (N_7805,N_6915,N_6552);
nand U7806 (N_7806,N_6825,N_6103);
xnor U7807 (N_7807,N_6998,N_6651);
or U7808 (N_7808,N_6894,N_6530);
and U7809 (N_7809,N_6855,N_6934);
nor U7810 (N_7810,N_6668,N_6481);
and U7811 (N_7811,N_6142,N_6865);
and U7812 (N_7812,N_6861,N_6741);
and U7813 (N_7813,N_6889,N_6579);
nor U7814 (N_7814,N_6687,N_6683);
nor U7815 (N_7815,N_6278,N_6934);
nor U7816 (N_7816,N_6684,N_6470);
xor U7817 (N_7817,N_6429,N_6888);
nand U7818 (N_7818,N_6743,N_6054);
and U7819 (N_7819,N_6919,N_6894);
nand U7820 (N_7820,N_6358,N_6008);
xor U7821 (N_7821,N_6270,N_6405);
or U7822 (N_7822,N_6824,N_6815);
or U7823 (N_7823,N_6383,N_6664);
or U7824 (N_7824,N_6629,N_6100);
and U7825 (N_7825,N_6934,N_6660);
or U7826 (N_7826,N_6785,N_6293);
xor U7827 (N_7827,N_6234,N_6461);
and U7828 (N_7828,N_6704,N_6163);
nand U7829 (N_7829,N_6440,N_6475);
or U7830 (N_7830,N_6185,N_6086);
xor U7831 (N_7831,N_6938,N_6309);
nand U7832 (N_7832,N_6808,N_6512);
nand U7833 (N_7833,N_6890,N_6949);
xnor U7834 (N_7834,N_6954,N_6970);
xnor U7835 (N_7835,N_6479,N_6202);
and U7836 (N_7836,N_6199,N_6691);
nand U7837 (N_7837,N_6959,N_6706);
nand U7838 (N_7838,N_6933,N_6635);
nor U7839 (N_7839,N_6947,N_6216);
nor U7840 (N_7840,N_6691,N_6353);
or U7841 (N_7841,N_6513,N_6238);
or U7842 (N_7842,N_6073,N_6268);
or U7843 (N_7843,N_6519,N_6404);
or U7844 (N_7844,N_6817,N_6872);
nand U7845 (N_7845,N_6201,N_6611);
xnor U7846 (N_7846,N_6512,N_6316);
or U7847 (N_7847,N_6141,N_6346);
and U7848 (N_7848,N_6856,N_6100);
or U7849 (N_7849,N_6867,N_6660);
nand U7850 (N_7850,N_6544,N_6976);
nor U7851 (N_7851,N_6823,N_6951);
nor U7852 (N_7852,N_6110,N_6843);
and U7853 (N_7853,N_6564,N_6363);
or U7854 (N_7854,N_6047,N_6001);
nand U7855 (N_7855,N_6218,N_6556);
or U7856 (N_7856,N_6185,N_6776);
xnor U7857 (N_7857,N_6091,N_6119);
and U7858 (N_7858,N_6111,N_6300);
xnor U7859 (N_7859,N_6973,N_6022);
nor U7860 (N_7860,N_6891,N_6003);
and U7861 (N_7861,N_6085,N_6983);
xnor U7862 (N_7862,N_6285,N_6010);
nand U7863 (N_7863,N_6928,N_6491);
nor U7864 (N_7864,N_6097,N_6530);
and U7865 (N_7865,N_6663,N_6382);
xor U7866 (N_7866,N_6443,N_6486);
xnor U7867 (N_7867,N_6532,N_6314);
xor U7868 (N_7868,N_6263,N_6601);
nor U7869 (N_7869,N_6938,N_6670);
nand U7870 (N_7870,N_6733,N_6165);
nor U7871 (N_7871,N_6331,N_6346);
nor U7872 (N_7872,N_6729,N_6439);
or U7873 (N_7873,N_6046,N_6013);
and U7874 (N_7874,N_6417,N_6568);
nand U7875 (N_7875,N_6961,N_6797);
and U7876 (N_7876,N_6524,N_6195);
or U7877 (N_7877,N_6037,N_6548);
xnor U7878 (N_7878,N_6754,N_6119);
nand U7879 (N_7879,N_6960,N_6246);
xor U7880 (N_7880,N_6476,N_6556);
xnor U7881 (N_7881,N_6318,N_6144);
nand U7882 (N_7882,N_6245,N_6881);
nand U7883 (N_7883,N_6982,N_6152);
nand U7884 (N_7884,N_6311,N_6132);
and U7885 (N_7885,N_6224,N_6174);
nor U7886 (N_7886,N_6004,N_6940);
and U7887 (N_7887,N_6078,N_6192);
xor U7888 (N_7888,N_6983,N_6990);
nand U7889 (N_7889,N_6626,N_6489);
and U7890 (N_7890,N_6098,N_6785);
nor U7891 (N_7891,N_6504,N_6892);
or U7892 (N_7892,N_6141,N_6324);
nand U7893 (N_7893,N_6382,N_6211);
nor U7894 (N_7894,N_6038,N_6711);
and U7895 (N_7895,N_6263,N_6153);
or U7896 (N_7896,N_6830,N_6596);
and U7897 (N_7897,N_6887,N_6561);
and U7898 (N_7898,N_6960,N_6890);
nor U7899 (N_7899,N_6984,N_6810);
xnor U7900 (N_7900,N_6578,N_6750);
nand U7901 (N_7901,N_6450,N_6078);
xnor U7902 (N_7902,N_6515,N_6038);
xor U7903 (N_7903,N_6058,N_6386);
nor U7904 (N_7904,N_6147,N_6387);
nand U7905 (N_7905,N_6717,N_6527);
xor U7906 (N_7906,N_6206,N_6791);
nand U7907 (N_7907,N_6061,N_6694);
or U7908 (N_7908,N_6454,N_6263);
nor U7909 (N_7909,N_6719,N_6836);
nand U7910 (N_7910,N_6323,N_6240);
nand U7911 (N_7911,N_6560,N_6889);
nor U7912 (N_7912,N_6042,N_6575);
nor U7913 (N_7913,N_6610,N_6854);
or U7914 (N_7914,N_6198,N_6451);
nor U7915 (N_7915,N_6974,N_6177);
nand U7916 (N_7916,N_6042,N_6780);
nor U7917 (N_7917,N_6026,N_6744);
or U7918 (N_7918,N_6421,N_6458);
or U7919 (N_7919,N_6238,N_6123);
or U7920 (N_7920,N_6544,N_6359);
or U7921 (N_7921,N_6008,N_6577);
xnor U7922 (N_7922,N_6737,N_6939);
nand U7923 (N_7923,N_6584,N_6399);
xnor U7924 (N_7924,N_6372,N_6381);
nand U7925 (N_7925,N_6519,N_6205);
nand U7926 (N_7926,N_6557,N_6315);
nor U7927 (N_7927,N_6591,N_6584);
nor U7928 (N_7928,N_6867,N_6126);
nor U7929 (N_7929,N_6571,N_6287);
and U7930 (N_7930,N_6192,N_6194);
nand U7931 (N_7931,N_6828,N_6912);
or U7932 (N_7932,N_6094,N_6837);
and U7933 (N_7933,N_6825,N_6321);
nand U7934 (N_7934,N_6040,N_6790);
and U7935 (N_7935,N_6584,N_6819);
nand U7936 (N_7936,N_6106,N_6945);
xnor U7937 (N_7937,N_6661,N_6122);
or U7938 (N_7938,N_6796,N_6605);
nand U7939 (N_7939,N_6424,N_6473);
xnor U7940 (N_7940,N_6727,N_6605);
nand U7941 (N_7941,N_6457,N_6044);
nand U7942 (N_7942,N_6371,N_6734);
and U7943 (N_7943,N_6733,N_6258);
nand U7944 (N_7944,N_6628,N_6844);
or U7945 (N_7945,N_6861,N_6929);
and U7946 (N_7946,N_6017,N_6315);
xor U7947 (N_7947,N_6397,N_6857);
nor U7948 (N_7948,N_6075,N_6961);
xnor U7949 (N_7949,N_6538,N_6515);
or U7950 (N_7950,N_6648,N_6958);
and U7951 (N_7951,N_6394,N_6477);
nand U7952 (N_7952,N_6835,N_6049);
or U7953 (N_7953,N_6457,N_6718);
and U7954 (N_7954,N_6568,N_6788);
and U7955 (N_7955,N_6073,N_6353);
xor U7956 (N_7956,N_6036,N_6308);
or U7957 (N_7957,N_6186,N_6700);
nand U7958 (N_7958,N_6238,N_6033);
nand U7959 (N_7959,N_6927,N_6662);
nand U7960 (N_7960,N_6506,N_6774);
or U7961 (N_7961,N_6853,N_6990);
nand U7962 (N_7962,N_6693,N_6977);
and U7963 (N_7963,N_6524,N_6540);
xor U7964 (N_7964,N_6678,N_6124);
xnor U7965 (N_7965,N_6641,N_6282);
nor U7966 (N_7966,N_6427,N_6123);
nand U7967 (N_7967,N_6155,N_6832);
and U7968 (N_7968,N_6892,N_6215);
xnor U7969 (N_7969,N_6071,N_6662);
and U7970 (N_7970,N_6876,N_6085);
nor U7971 (N_7971,N_6905,N_6786);
nor U7972 (N_7972,N_6250,N_6254);
nand U7973 (N_7973,N_6282,N_6463);
nor U7974 (N_7974,N_6788,N_6602);
xnor U7975 (N_7975,N_6098,N_6218);
nor U7976 (N_7976,N_6843,N_6849);
and U7977 (N_7977,N_6842,N_6601);
or U7978 (N_7978,N_6887,N_6734);
nor U7979 (N_7979,N_6111,N_6997);
and U7980 (N_7980,N_6208,N_6050);
and U7981 (N_7981,N_6884,N_6367);
nor U7982 (N_7982,N_6739,N_6981);
xnor U7983 (N_7983,N_6236,N_6224);
nand U7984 (N_7984,N_6125,N_6733);
or U7985 (N_7985,N_6025,N_6947);
nor U7986 (N_7986,N_6359,N_6942);
or U7987 (N_7987,N_6235,N_6513);
and U7988 (N_7988,N_6996,N_6807);
nand U7989 (N_7989,N_6357,N_6744);
and U7990 (N_7990,N_6367,N_6187);
nand U7991 (N_7991,N_6009,N_6146);
nand U7992 (N_7992,N_6401,N_6253);
nor U7993 (N_7993,N_6770,N_6349);
and U7994 (N_7994,N_6566,N_6522);
nor U7995 (N_7995,N_6421,N_6367);
nand U7996 (N_7996,N_6821,N_6533);
or U7997 (N_7997,N_6953,N_6442);
xnor U7998 (N_7998,N_6685,N_6592);
and U7999 (N_7999,N_6827,N_6694);
or U8000 (N_8000,N_7131,N_7296);
xnor U8001 (N_8001,N_7850,N_7054);
xor U8002 (N_8002,N_7437,N_7786);
nor U8003 (N_8003,N_7022,N_7723);
and U8004 (N_8004,N_7954,N_7771);
nor U8005 (N_8005,N_7543,N_7338);
and U8006 (N_8006,N_7980,N_7959);
or U8007 (N_8007,N_7649,N_7453);
nor U8008 (N_8008,N_7204,N_7128);
and U8009 (N_8009,N_7216,N_7645);
and U8010 (N_8010,N_7059,N_7000);
xor U8011 (N_8011,N_7307,N_7776);
xor U8012 (N_8012,N_7225,N_7475);
nand U8013 (N_8013,N_7541,N_7501);
xor U8014 (N_8014,N_7751,N_7125);
and U8015 (N_8015,N_7246,N_7197);
nor U8016 (N_8016,N_7862,N_7934);
xnor U8017 (N_8017,N_7393,N_7871);
and U8018 (N_8018,N_7895,N_7271);
xnor U8019 (N_8019,N_7029,N_7426);
nor U8020 (N_8020,N_7117,N_7242);
and U8021 (N_8021,N_7889,N_7123);
nand U8022 (N_8022,N_7268,N_7989);
or U8023 (N_8023,N_7406,N_7354);
nand U8024 (N_8024,N_7876,N_7181);
xor U8025 (N_8025,N_7510,N_7162);
or U8026 (N_8026,N_7542,N_7223);
nor U8027 (N_8027,N_7262,N_7208);
or U8028 (N_8028,N_7695,N_7798);
xnor U8029 (N_8029,N_7352,N_7928);
nor U8030 (N_8030,N_7791,N_7859);
nor U8031 (N_8031,N_7881,N_7624);
xor U8032 (N_8032,N_7807,N_7300);
and U8033 (N_8033,N_7089,N_7970);
or U8034 (N_8034,N_7962,N_7425);
nand U8035 (N_8035,N_7444,N_7714);
xnor U8036 (N_8036,N_7210,N_7343);
xnor U8037 (N_8037,N_7294,N_7825);
and U8038 (N_8038,N_7056,N_7500);
or U8039 (N_8039,N_7953,N_7068);
and U8040 (N_8040,N_7212,N_7449);
nand U8041 (N_8041,N_7183,N_7906);
nand U8042 (N_8042,N_7536,N_7037);
and U8043 (N_8043,N_7978,N_7486);
xnor U8044 (N_8044,N_7764,N_7076);
nand U8045 (N_8045,N_7824,N_7707);
xor U8046 (N_8046,N_7885,N_7992);
nor U8047 (N_8047,N_7255,N_7991);
and U8048 (N_8048,N_7739,N_7321);
nand U8049 (N_8049,N_7839,N_7579);
xnor U8050 (N_8050,N_7247,N_7091);
xnor U8051 (N_8051,N_7062,N_7166);
xor U8052 (N_8052,N_7506,N_7362);
nand U8053 (N_8053,N_7176,N_7511);
nand U8054 (N_8054,N_7842,N_7150);
nor U8055 (N_8055,N_7921,N_7400);
nor U8056 (N_8056,N_7974,N_7904);
or U8057 (N_8057,N_7168,N_7256);
or U8058 (N_8058,N_7941,N_7588);
nor U8059 (N_8059,N_7907,N_7872);
xnor U8060 (N_8060,N_7985,N_7388);
and U8061 (N_8061,N_7323,N_7113);
or U8062 (N_8062,N_7621,N_7823);
and U8063 (N_8063,N_7404,N_7005);
nor U8064 (N_8064,N_7502,N_7121);
nor U8065 (N_8065,N_7287,N_7283);
nor U8066 (N_8066,N_7900,N_7844);
and U8067 (N_8067,N_7046,N_7464);
or U8068 (N_8068,N_7526,N_7996);
or U8069 (N_8069,N_7401,N_7447);
xor U8070 (N_8070,N_7908,N_7341);
or U8071 (N_8071,N_7164,N_7157);
and U8072 (N_8072,N_7568,N_7703);
nor U8073 (N_8073,N_7747,N_7259);
nand U8074 (N_8074,N_7892,N_7186);
and U8075 (N_8075,N_7680,N_7976);
or U8076 (N_8076,N_7184,N_7828);
nand U8077 (N_8077,N_7705,N_7538);
nor U8078 (N_8078,N_7377,N_7968);
xor U8079 (N_8079,N_7518,N_7810);
nor U8080 (N_8080,N_7522,N_7493);
nand U8081 (N_8081,N_7656,N_7965);
nand U8082 (N_8082,N_7671,N_7334);
xor U8083 (N_8083,N_7863,N_7491);
xor U8084 (N_8084,N_7883,N_7407);
and U8085 (N_8085,N_7455,N_7398);
nand U8086 (N_8086,N_7483,N_7295);
nor U8087 (N_8087,N_7207,N_7653);
nor U8088 (N_8088,N_7039,N_7547);
and U8089 (N_8089,N_7152,N_7815);
xnor U8090 (N_8090,N_7631,N_7231);
or U8091 (N_8091,N_7233,N_7086);
nor U8092 (N_8092,N_7413,N_7610);
nand U8093 (N_8093,N_7877,N_7441);
nand U8094 (N_8094,N_7726,N_7608);
xnor U8095 (N_8095,N_7744,N_7688);
xor U8096 (N_8096,N_7137,N_7912);
and U8097 (N_8097,N_7894,N_7622);
xnor U8098 (N_8098,N_7279,N_7067);
nand U8099 (N_8099,N_7971,N_7618);
xor U8100 (N_8100,N_7571,N_7517);
or U8101 (N_8101,N_7848,N_7161);
xor U8102 (N_8102,N_7053,N_7069);
or U8103 (N_8103,N_7209,N_7276);
and U8104 (N_8104,N_7265,N_7213);
nor U8105 (N_8105,N_7781,N_7837);
nor U8106 (N_8106,N_7675,N_7008);
xor U8107 (N_8107,N_7336,N_7898);
and U8108 (N_8108,N_7301,N_7014);
xnor U8109 (N_8109,N_7679,N_7901);
nor U8110 (N_8110,N_7326,N_7512);
nand U8111 (N_8111,N_7686,N_7106);
xnor U8112 (N_8112,N_7796,N_7221);
xor U8113 (N_8113,N_7473,N_7016);
and U8114 (N_8114,N_7869,N_7293);
nor U8115 (N_8115,N_7580,N_7327);
or U8116 (N_8116,N_7690,N_7964);
and U8117 (N_8117,N_7487,N_7760);
and U8118 (N_8118,N_7499,N_7017);
nor U8119 (N_8119,N_7820,N_7100);
nor U8120 (N_8120,N_7396,N_7290);
or U8121 (N_8121,N_7075,N_7155);
nand U8122 (N_8122,N_7597,N_7103);
xor U8123 (N_8123,N_7361,N_7915);
nand U8124 (N_8124,N_7419,N_7598);
and U8125 (N_8125,N_7972,N_7110);
nor U8126 (N_8126,N_7582,N_7732);
or U8127 (N_8127,N_7034,N_7277);
xnor U8128 (N_8128,N_7789,N_7566);
and U8129 (N_8129,N_7381,N_7083);
nor U8130 (N_8130,N_7725,N_7812);
and U8131 (N_8131,N_7599,N_7006);
nand U8132 (N_8132,N_7389,N_7572);
nor U8133 (N_8133,N_7120,N_7535);
xnor U8134 (N_8134,N_7662,N_7809);
xnor U8135 (N_8135,N_7460,N_7569);
nor U8136 (N_8136,N_7590,N_7643);
or U8137 (N_8137,N_7663,N_7811);
or U8138 (N_8138,N_7281,N_7678);
and U8139 (N_8139,N_7145,N_7981);
or U8140 (N_8140,N_7498,N_7350);
xor U8141 (N_8141,N_7768,N_7891);
or U8142 (N_8142,N_7485,N_7430);
xor U8143 (N_8143,N_7717,N_7418);
or U8144 (N_8144,N_7021,N_7530);
nand U8145 (N_8145,N_7840,N_7387);
and U8146 (N_8146,N_7759,N_7031);
xor U8147 (N_8147,N_7278,N_7190);
or U8148 (N_8148,N_7490,N_7911);
nor U8149 (N_8149,N_7559,N_7966);
and U8150 (N_8150,N_7456,N_7836);
nor U8151 (N_8151,N_7045,N_7557);
xnor U8152 (N_8152,N_7886,N_7697);
or U8153 (N_8153,N_7097,N_7357);
xnor U8154 (N_8154,N_7689,N_7058);
nand U8155 (N_8155,N_7537,N_7470);
and U8156 (N_8156,N_7332,N_7769);
and U8157 (N_8157,N_7269,N_7292);
or U8158 (N_8158,N_7636,N_7369);
and U8159 (N_8159,N_7451,N_7267);
xor U8160 (N_8160,N_7040,N_7665);
and U8161 (N_8161,N_7193,N_7392);
nand U8162 (N_8162,N_7520,N_7140);
nor U8163 (N_8163,N_7821,N_7731);
or U8164 (N_8164,N_7803,N_7750);
or U8165 (N_8165,N_7880,N_7394);
and U8166 (N_8166,N_7578,N_7122);
xnor U8167 (N_8167,N_7669,N_7195);
or U8168 (N_8168,N_7468,N_7047);
or U8169 (N_8169,N_7755,N_7084);
nor U8170 (N_8170,N_7007,N_7232);
and U8171 (N_8171,N_7317,N_7135);
and U8172 (N_8172,N_7777,N_7462);
or U8173 (N_8173,N_7275,N_7693);
or U8174 (N_8174,N_7129,N_7217);
nand U8175 (N_8175,N_7312,N_7030);
nand U8176 (N_8176,N_7314,N_7860);
xnor U8177 (N_8177,N_7364,N_7534);
xor U8178 (N_8178,N_7710,N_7998);
nor U8179 (N_8179,N_7923,N_7814);
and U8180 (N_8180,N_7325,N_7527);
xor U8181 (N_8181,N_7476,N_7395);
and U8182 (N_8182,N_7228,N_7523);
or U8183 (N_8183,N_7153,N_7435);
and U8184 (N_8184,N_7728,N_7893);
nor U8185 (N_8185,N_7639,N_7514);
xor U8186 (N_8186,N_7788,N_7593);
xnor U8187 (N_8187,N_7932,N_7497);
xnor U8188 (N_8188,N_7422,N_7933);
and U8189 (N_8189,N_7920,N_7177);
or U8190 (N_8190,N_7730,N_7549);
xor U8191 (N_8191,N_7298,N_7148);
or U8192 (N_8192,N_7185,N_7757);
and U8193 (N_8193,N_7105,N_7215);
and U8194 (N_8194,N_7107,N_7875);
and U8195 (N_8195,N_7489,N_7592);
and U8196 (N_8196,N_7994,N_7507);
and U8197 (N_8197,N_7924,N_7719);
and U8198 (N_8198,N_7940,N_7019);
and U8199 (N_8199,N_7074,N_7218);
xnor U8200 (N_8200,N_7052,N_7041);
and U8201 (N_8201,N_7613,N_7482);
nor U8202 (N_8202,N_7124,N_7554);
xnor U8203 (N_8203,N_7315,N_7160);
and U8204 (N_8204,N_7254,N_7480);
nand U8205 (N_8205,N_7372,N_7651);
or U8206 (N_8206,N_7712,N_7002);
nand U8207 (N_8207,N_7085,N_7257);
nor U8208 (N_8208,N_7127,N_7439);
nor U8209 (N_8209,N_7635,N_7577);
nand U8210 (N_8210,N_7311,N_7556);
and U8211 (N_8211,N_7594,N_7260);
xnor U8212 (N_8212,N_7250,N_7179);
or U8213 (N_8213,N_7513,N_7503);
xor U8214 (N_8214,N_7531,N_7383);
nor U8215 (N_8215,N_7385,N_7943);
nand U8216 (N_8216,N_7775,N_7787);
and U8217 (N_8217,N_7214,N_7095);
and U8218 (N_8218,N_7676,N_7716);
nand U8219 (N_8219,N_7013,N_7371);
or U8220 (N_8220,N_7375,N_7586);
and U8221 (N_8221,N_7248,N_7852);
or U8222 (N_8222,N_7263,N_7887);
xnor U8223 (N_8223,N_7222,N_7648);
or U8224 (N_8224,N_7691,N_7038);
nand U8225 (N_8225,N_7333,N_7025);
nor U8226 (N_8226,N_7525,N_7958);
or U8227 (N_8227,N_7251,N_7012);
or U8228 (N_8228,N_7191,N_7303);
nand U8229 (N_8229,N_7754,N_7144);
nor U8230 (N_8230,N_7339,N_7802);
and U8231 (N_8231,N_7200,N_7328);
xnor U8232 (N_8232,N_7685,N_7558);
and U8233 (N_8233,N_7093,N_7082);
nor U8234 (N_8234,N_7956,N_7727);
nand U8235 (N_8235,N_7938,N_7515);
nor U8236 (N_8236,N_7443,N_7795);
nand U8237 (N_8237,N_7196,N_7602);
nand U8238 (N_8238,N_7858,N_7785);
or U8239 (N_8239,N_7702,N_7826);
nand U8240 (N_8240,N_7829,N_7118);
and U8241 (N_8241,N_7611,N_7841);
and U8242 (N_8242,N_7681,N_7199);
nor U8243 (N_8243,N_7734,N_7565);
nor U8244 (N_8244,N_7987,N_7851);
xor U8245 (N_8245,N_7182,N_7316);
xor U8246 (N_8246,N_7092,N_7450);
nor U8247 (N_8247,N_7818,N_7947);
or U8248 (N_8248,N_7386,N_7674);
xor U8249 (N_8249,N_7553,N_7477);
nor U8250 (N_8250,N_7461,N_7696);
nand U8251 (N_8251,N_7718,N_7666);
or U8252 (N_8252,N_7655,N_7711);
or U8253 (N_8253,N_7607,N_7736);
or U8254 (N_8254,N_7353,N_7471);
nor U8255 (N_8255,N_7431,N_7806);
nor U8256 (N_8256,N_7741,N_7945);
or U8257 (N_8257,N_7359,N_7104);
and U8258 (N_8258,N_7416,N_7027);
and U8259 (N_8259,N_7993,N_7935);
and U8260 (N_8260,N_7562,N_7567);
nor U8261 (N_8261,N_7835,N_7308);
or U8262 (N_8262,N_7746,N_7799);
or U8263 (N_8263,N_7999,N_7832);
xnor U8264 (N_8264,N_7733,N_7884);
or U8265 (N_8265,N_7819,N_7412);
or U8266 (N_8266,N_7600,N_7310);
and U8267 (N_8267,N_7245,N_7949);
and U8268 (N_8268,N_7201,N_7478);
nor U8269 (N_8269,N_7304,N_7952);
nand U8270 (N_8270,N_7855,N_7094);
nor U8271 (N_8271,N_7220,N_7903);
nor U8272 (N_8272,N_7004,N_7454);
xor U8273 (N_8273,N_7149,N_7939);
nand U8274 (N_8274,N_7459,N_7202);
xnor U8275 (N_8275,N_7780,N_7172);
nor U8276 (N_8276,N_7291,N_7864);
nand U8277 (N_8277,N_7043,N_7738);
nor U8278 (N_8278,N_7763,N_7615);
xor U8279 (N_8279,N_7355,N_7857);
xnor U8280 (N_8280,N_7948,N_7324);
xor U8281 (N_8281,N_7380,N_7146);
nor U8282 (N_8282,N_7946,N_7023);
nor U8283 (N_8283,N_7772,N_7761);
nand U8284 (N_8284,N_7440,N_7575);
xnor U8285 (N_8285,N_7720,N_7982);
xor U8286 (N_8286,N_7365,N_7488);
xor U8287 (N_8287,N_7770,N_7061);
nor U8288 (N_8288,N_7042,N_7423);
and U8289 (N_8289,N_7944,N_7274);
nor U8290 (N_8290,N_7629,N_7758);
and U8291 (N_8291,N_7874,N_7415);
nand U8292 (N_8292,N_7630,N_7158);
and U8293 (N_8293,N_7505,N_7638);
and U8294 (N_8294,N_7099,N_7853);
xor U8295 (N_8295,N_7227,N_7329);
nor U8296 (N_8296,N_7018,N_7767);
nand U8297 (N_8297,N_7986,N_7130);
xor U8298 (N_8298,N_7918,N_7701);
nor U8299 (N_8299,N_7692,N_7282);
xnor U8300 (N_8300,N_7410,N_7253);
nor U8301 (N_8301,N_7936,N_7897);
or U8302 (N_8302,N_7673,N_7438);
or U8303 (N_8303,N_7408,N_7109);
xor U8304 (N_8304,N_7838,N_7240);
nor U8305 (N_8305,N_7374,N_7126);
nor U8306 (N_8306,N_7044,N_7114);
and U8307 (N_8307,N_7188,N_7899);
and U8308 (N_8308,N_7942,N_7830);
nand U8309 (N_8309,N_7721,N_7171);
and U8310 (N_8310,N_7226,N_7286);
nor U8311 (N_8311,N_7805,N_7737);
nand U8312 (N_8312,N_7102,N_7509);
nor U8313 (N_8313,N_7816,N_7573);
xor U8314 (N_8314,N_7141,N_7927);
and U8315 (N_8315,N_7762,N_7951);
nor U8316 (N_8316,N_7448,N_7132);
and U8317 (N_8317,N_7793,N_7545);
xnor U8318 (N_8318,N_7847,N_7187);
and U8319 (N_8319,N_7910,N_7672);
nand U8320 (N_8320,N_7765,N_7194);
xor U8321 (N_8321,N_7108,N_7048);
or U8322 (N_8322,N_7896,N_7390);
xor U8323 (N_8323,N_7417,N_7403);
or U8324 (N_8324,N_7516,N_7722);
nor U8325 (N_8325,N_7589,N_7474);
and U8326 (N_8326,N_7591,N_7784);
nor U8327 (N_8327,N_7873,N_7612);
nand U8328 (N_8328,N_7698,N_7159);
or U8329 (N_8329,N_7112,N_7211);
or U8330 (N_8330,N_7133,N_7345);
xnor U8331 (N_8331,N_7077,N_7646);
and U8332 (N_8332,N_7072,N_7684);
and U8333 (N_8333,N_7467,N_7309);
xor U8334 (N_8334,N_7609,N_7879);
nor U8335 (N_8335,N_7682,N_7306);
nor U8336 (N_8336,N_7272,N_7521);
and U8337 (N_8337,N_7337,N_7929);
nor U8338 (N_8338,N_7561,N_7640);
or U8339 (N_8339,N_7654,N_7800);
nor U8340 (N_8340,N_7090,N_7601);
nand U8341 (N_8341,N_7484,N_7289);
or U8342 (N_8342,N_7313,N_7614);
xnor U8343 (N_8343,N_7078,N_7351);
or U8344 (N_8344,N_7529,N_7111);
and U8345 (N_8345,N_7551,N_7165);
nand U8346 (N_8346,N_7546,N_7748);
nor U8347 (N_8347,N_7683,N_7931);
nand U8348 (N_8348,N_7713,N_7657);
nor U8349 (N_8349,N_7280,N_7011);
nor U8350 (N_8350,N_7913,N_7424);
nor U8351 (N_8351,N_7540,N_7555);
or U8352 (N_8352,N_7234,N_7865);
and U8353 (N_8353,N_7180,N_7930);
nand U8354 (N_8354,N_7270,N_7032);
or U8355 (N_8355,N_7596,N_7797);
nand U8356 (N_8356,N_7584,N_7349);
nor U8357 (N_8357,N_7409,N_7977);
nand U8358 (N_8358,N_7028,N_7519);
nand U8359 (N_8359,N_7560,N_7318);
nor U8360 (N_8360,N_7634,N_7302);
xor U8361 (N_8361,N_7378,N_7147);
nor U8362 (N_8362,N_7495,N_7020);
xor U8363 (N_8363,N_7975,N_7660);
nand U8364 (N_8364,N_7340,N_7376);
xor U8365 (N_8365,N_7436,N_7687);
nand U8366 (N_8366,N_7652,N_7670);
xor U8367 (N_8367,N_7319,N_7466);
nor U8368 (N_8368,N_7442,N_7729);
or U8369 (N_8369,N_7492,N_7967);
nand U8370 (N_8370,N_7742,N_7632);
and U8371 (N_8371,N_7065,N_7370);
nor U8372 (N_8372,N_7330,N_7647);
nand U8373 (N_8373,N_7134,N_7363);
nor U8374 (N_8374,N_7890,N_7576);
and U8375 (N_8375,N_7241,N_7969);
and U8376 (N_8376,N_7914,N_7642);
or U8377 (N_8377,N_7446,N_7868);
nor U8378 (N_8378,N_7595,N_7659);
xor U8379 (N_8379,N_7382,N_7445);
nor U8380 (N_8380,N_7817,N_7342);
xnor U8381 (N_8381,N_7834,N_7055);
and U8382 (N_8382,N_7205,N_7979);
or U8383 (N_8383,N_7533,N_7249);
nand U8384 (N_8384,N_7548,N_7585);
nand U8385 (N_8385,N_7922,N_7237);
nand U8386 (N_8386,N_7532,N_7175);
xnor U8387 (N_8387,N_7285,N_7570);
xor U8388 (N_8388,N_7650,N_7743);
xnor U8389 (N_8389,N_7957,N_7917);
nand U8390 (N_8390,N_7997,N_7051);
nand U8391 (N_8391,N_7229,N_7539);
nor U8392 (N_8392,N_7366,N_7288);
nor U8393 (N_8393,N_7098,N_7358);
and U8394 (N_8394,N_7955,N_7322);
nor U8395 (N_8395,N_7888,N_7224);
and U8396 (N_8396,N_7273,N_7628);
nor U8397 (N_8397,N_7411,N_7709);
and U8398 (N_8398,N_7715,N_7902);
nand U8399 (N_8399,N_7178,N_7472);
nand U8400 (N_8400,N_7668,N_7866);
and U8401 (N_8401,N_7049,N_7804);
and U8402 (N_8402,N_7988,N_7552);
or U8403 (N_8403,N_7479,N_7015);
nor U8404 (N_8404,N_7606,N_7481);
xor U8405 (N_8405,N_7783,N_7524);
xnor U8406 (N_8406,N_7603,N_7916);
xnor U8407 (N_8407,N_7457,N_7399);
and U8408 (N_8408,N_7173,N_7036);
or U8409 (N_8409,N_7667,N_7658);
and U8410 (N_8410,N_7604,N_7119);
nand U8411 (N_8411,N_7633,N_7427);
xor U8412 (N_8412,N_7238,N_7574);
xnor U8413 (N_8413,N_7235,N_7854);
and U8414 (N_8414,N_7347,N_7790);
or U8415 (N_8415,N_7139,N_7833);
or U8416 (N_8416,N_7845,N_7073);
xor U8417 (N_8417,N_7623,N_7071);
and U8418 (N_8418,N_7026,N_7626);
or U8419 (N_8419,N_7230,N_7661);
nor U8420 (N_8420,N_7849,N_7878);
nor U8421 (N_8421,N_7244,N_7414);
xor U8422 (N_8422,N_7432,N_7961);
xnor U8423 (N_8423,N_7239,N_7391);
or U8424 (N_8424,N_7050,N_7033);
nor U8425 (N_8425,N_7344,N_7143);
and U8426 (N_8426,N_7081,N_7984);
and U8427 (N_8427,N_7779,N_7297);
or U8428 (N_8428,N_7960,N_7236);
and U8429 (N_8429,N_7360,N_7079);
and U8430 (N_8430,N_7792,N_7116);
xor U8431 (N_8431,N_7174,N_7243);
or U8432 (N_8432,N_7627,N_7001);
xnor U8433 (N_8433,N_7060,N_7937);
xor U8434 (N_8434,N_7420,N_7368);
nand U8435 (N_8435,N_7831,N_7331);
and U8436 (N_8436,N_7990,N_7066);
or U8437 (N_8437,N_7167,N_7384);
xnor U8438 (N_8438,N_7995,N_7528);
xnor U8439 (N_8439,N_7808,N_7198);
and U8440 (N_8440,N_7169,N_7973);
xor U8441 (N_8441,N_7861,N_7694);
nor U8442 (N_8442,N_7756,N_7773);
nor U8443 (N_8443,N_7919,N_7465);
nor U8444 (N_8444,N_7284,N_7494);
or U8445 (N_8445,N_7402,N_7469);
or U8446 (N_8446,N_7320,N_7782);
or U8447 (N_8447,N_7496,N_7905);
and U8448 (N_8448,N_7142,N_7843);
nor U8449 (N_8449,N_7348,N_7813);
nor U8450 (N_8450,N_7063,N_7356);
and U8451 (N_8451,N_7266,N_7827);
and U8452 (N_8452,N_7421,N_7963);
nand U8453 (N_8453,N_7637,N_7138);
nand U8454 (N_8454,N_7677,N_7070);
nand U8455 (N_8455,N_7508,N_7189);
nand U8456 (N_8456,N_7644,N_7064);
or U8457 (N_8457,N_7305,N_7700);
nand U8458 (N_8458,N_7463,N_7379);
and U8459 (N_8459,N_7080,N_7088);
nor U8460 (N_8460,N_7620,N_7335);
nand U8461 (N_8461,N_7010,N_7587);
nand U8462 (N_8462,N_7009,N_7616);
xor U8463 (N_8463,N_7544,N_7154);
or U8464 (N_8464,N_7428,N_7170);
xor U8465 (N_8465,N_7774,N_7219);
nor U8466 (N_8466,N_7724,N_7504);
and U8467 (N_8467,N_7101,N_7035);
and U8468 (N_8468,N_7822,N_7429);
or U8469 (N_8469,N_7664,N_7752);
and U8470 (N_8470,N_7264,N_7151);
nor U8471 (N_8471,N_7926,N_7096);
and U8472 (N_8472,N_7983,N_7882);
and U8473 (N_8473,N_7346,N_7405);
xnor U8474 (N_8474,N_7909,N_7057);
nor U8475 (N_8475,N_7706,N_7625);
xnor U8476 (N_8476,N_7699,N_7745);
or U8477 (N_8477,N_7550,N_7753);
nor U8478 (N_8478,N_7749,N_7452);
nor U8479 (N_8479,N_7641,N_7708);
nor U8480 (N_8480,N_7870,N_7203);
or U8481 (N_8481,N_7024,N_7740);
xor U8482 (N_8482,N_7704,N_7581);
and U8483 (N_8483,N_7867,N_7617);
nor U8484 (N_8484,N_7563,N_7299);
nor U8485 (N_8485,N_7766,N_7605);
nand U8486 (N_8486,N_7735,N_7846);
or U8487 (N_8487,N_7087,N_7258);
xor U8488 (N_8488,N_7564,N_7252);
and U8489 (N_8489,N_7192,N_7950);
and U8490 (N_8490,N_7156,N_7373);
nor U8491 (N_8491,N_7003,N_7619);
xor U8492 (N_8492,N_7115,N_7136);
nand U8493 (N_8493,N_7261,N_7433);
and U8494 (N_8494,N_7397,N_7458);
nand U8495 (N_8495,N_7778,N_7583);
nand U8496 (N_8496,N_7794,N_7163);
xnor U8497 (N_8497,N_7801,N_7206);
and U8498 (N_8498,N_7434,N_7367);
and U8499 (N_8499,N_7856,N_7925);
xor U8500 (N_8500,N_7112,N_7117);
and U8501 (N_8501,N_7954,N_7783);
or U8502 (N_8502,N_7321,N_7531);
nor U8503 (N_8503,N_7510,N_7937);
nor U8504 (N_8504,N_7701,N_7743);
nor U8505 (N_8505,N_7776,N_7240);
and U8506 (N_8506,N_7357,N_7192);
nand U8507 (N_8507,N_7513,N_7574);
and U8508 (N_8508,N_7719,N_7016);
nand U8509 (N_8509,N_7588,N_7388);
xor U8510 (N_8510,N_7274,N_7965);
xor U8511 (N_8511,N_7860,N_7353);
or U8512 (N_8512,N_7306,N_7378);
nand U8513 (N_8513,N_7240,N_7183);
nor U8514 (N_8514,N_7848,N_7988);
nand U8515 (N_8515,N_7510,N_7547);
and U8516 (N_8516,N_7591,N_7831);
or U8517 (N_8517,N_7186,N_7215);
xnor U8518 (N_8518,N_7644,N_7459);
and U8519 (N_8519,N_7070,N_7337);
or U8520 (N_8520,N_7714,N_7947);
nor U8521 (N_8521,N_7931,N_7620);
nand U8522 (N_8522,N_7340,N_7741);
nor U8523 (N_8523,N_7203,N_7070);
nand U8524 (N_8524,N_7584,N_7936);
nor U8525 (N_8525,N_7333,N_7091);
xor U8526 (N_8526,N_7988,N_7745);
or U8527 (N_8527,N_7676,N_7599);
or U8528 (N_8528,N_7307,N_7702);
nand U8529 (N_8529,N_7769,N_7854);
or U8530 (N_8530,N_7409,N_7925);
or U8531 (N_8531,N_7220,N_7063);
nor U8532 (N_8532,N_7151,N_7964);
nand U8533 (N_8533,N_7957,N_7720);
or U8534 (N_8534,N_7727,N_7673);
nor U8535 (N_8535,N_7814,N_7514);
and U8536 (N_8536,N_7831,N_7380);
xor U8537 (N_8537,N_7805,N_7101);
nor U8538 (N_8538,N_7005,N_7816);
xor U8539 (N_8539,N_7481,N_7117);
nand U8540 (N_8540,N_7693,N_7670);
xor U8541 (N_8541,N_7388,N_7542);
and U8542 (N_8542,N_7435,N_7189);
and U8543 (N_8543,N_7691,N_7377);
and U8544 (N_8544,N_7762,N_7022);
nand U8545 (N_8545,N_7761,N_7109);
and U8546 (N_8546,N_7446,N_7544);
nand U8547 (N_8547,N_7300,N_7956);
nor U8548 (N_8548,N_7241,N_7903);
and U8549 (N_8549,N_7069,N_7398);
nor U8550 (N_8550,N_7647,N_7838);
or U8551 (N_8551,N_7161,N_7890);
and U8552 (N_8552,N_7108,N_7683);
nand U8553 (N_8553,N_7653,N_7178);
nand U8554 (N_8554,N_7342,N_7602);
xor U8555 (N_8555,N_7945,N_7477);
and U8556 (N_8556,N_7761,N_7660);
xor U8557 (N_8557,N_7772,N_7214);
and U8558 (N_8558,N_7554,N_7081);
and U8559 (N_8559,N_7237,N_7766);
nor U8560 (N_8560,N_7008,N_7232);
nor U8561 (N_8561,N_7167,N_7529);
and U8562 (N_8562,N_7274,N_7679);
nand U8563 (N_8563,N_7098,N_7736);
nand U8564 (N_8564,N_7560,N_7559);
nor U8565 (N_8565,N_7684,N_7948);
xnor U8566 (N_8566,N_7539,N_7380);
and U8567 (N_8567,N_7124,N_7959);
nor U8568 (N_8568,N_7676,N_7210);
nor U8569 (N_8569,N_7003,N_7115);
xnor U8570 (N_8570,N_7531,N_7091);
nand U8571 (N_8571,N_7158,N_7604);
or U8572 (N_8572,N_7809,N_7484);
nor U8573 (N_8573,N_7272,N_7434);
or U8574 (N_8574,N_7555,N_7889);
nor U8575 (N_8575,N_7756,N_7671);
or U8576 (N_8576,N_7128,N_7979);
and U8577 (N_8577,N_7778,N_7454);
nand U8578 (N_8578,N_7455,N_7559);
xor U8579 (N_8579,N_7046,N_7422);
nor U8580 (N_8580,N_7078,N_7856);
and U8581 (N_8581,N_7313,N_7649);
xor U8582 (N_8582,N_7953,N_7134);
or U8583 (N_8583,N_7652,N_7281);
and U8584 (N_8584,N_7701,N_7417);
nand U8585 (N_8585,N_7444,N_7170);
nor U8586 (N_8586,N_7168,N_7244);
or U8587 (N_8587,N_7670,N_7444);
xor U8588 (N_8588,N_7137,N_7697);
or U8589 (N_8589,N_7485,N_7665);
nand U8590 (N_8590,N_7951,N_7687);
nand U8591 (N_8591,N_7235,N_7955);
xnor U8592 (N_8592,N_7045,N_7856);
nor U8593 (N_8593,N_7697,N_7332);
and U8594 (N_8594,N_7053,N_7961);
nand U8595 (N_8595,N_7653,N_7020);
xnor U8596 (N_8596,N_7071,N_7636);
nor U8597 (N_8597,N_7545,N_7252);
or U8598 (N_8598,N_7820,N_7111);
nor U8599 (N_8599,N_7798,N_7379);
or U8600 (N_8600,N_7599,N_7093);
and U8601 (N_8601,N_7251,N_7476);
or U8602 (N_8602,N_7283,N_7093);
nor U8603 (N_8603,N_7550,N_7922);
xnor U8604 (N_8604,N_7038,N_7569);
or U8605 (N_8605,N_7603,N_7033);
nor U8606 (N_8606,N_7101,N_7511);
or U8607 (N_8607,N_7163,N_7276);
nor U8608 (N_8608,N_7950,N_7187);
or U8609 (N_8609,N_7161,N_7533);
nor U8610 (N_8610,N_7901,N_7297);
or U8611 (N_8611,N_7821,N_7878);
nand U8612 (N_8612,N_7178,N_7081);
xor U8613 (N_8613,N_7961,N_7298);
xor U8614 (N_8614,N_7808,N_7648);
nor U8615 (N_8615,N_7132,N_7838);
xor U8616 (N_8616,N_7539,N_7098);
nand U8617 (N_8617,N_7561,N_7426);
and U8618 (N_8618,N_7254,N_7119);
nand U8619 (N_8619,N_7812,N_7310);
xor U8620 (N_8620,N_7245,N_7416);
xnor U8621 (N_8621,N_7202,N_7927);
and U8622 (N_8622,N_7485,N_7164);
or U8623 (N_8623,N_7005,N_7317);
nor U8624 (N_8624,N_7114,N_7817);
or U8625 (N_8625,N_7104,N_7989);
and U8626 (N_8626,N_7533,N_7350);
nor U8627 (N_8627,N_7942,N_7131);
nand U8628 (N_8628,N_7608,N_7839);
nand U8629 (N_8629,N_7627,N_7459);
xor U8630 (N_8630,N_7133,N_7948);
and U8631 (N_8631,N_7633,N_7942);
xor U8632 (N_8632,N_7741,N_7067);
xor U8633 (N_8633,N_7335,N_7592);
nor U8634 (N_8634,N_7075,N_7862);
nand U8635 (N_8635,N_7776,N_7115);
or U8636 (N_8636,N_7812,N_7869);
nand U8637 (N_8637,N_7394,N_7875);
xnor U8638 (N_8638,N_7044,N_7231);
and U8639 (N_8639,N_7526,N_7168);
xor U8640 (N_8640,N_7954,N_7503);
xnor U8641 (N_8641,N_7901,N_7692);
and U8642 (N_8642,N_7599,N_7987);
xnor U8643 (N_8643,N_7963,N_7779);
nand U8644 (N_8644,N_7600,N_7274);
xor U8645 (N_8645,N_7044,N_7597);
xnor U8646 (N_8646,N_7449,N_7247);
and U8647 (N_8647,N_7733,N_7020);
and U8648 (N_8648,N_7574,N_7611);
nor U8649 (N_8649,N_7609,N_7633);
xnor U8650 (N_8650,N_7867,N_7263);
nand U8651 (N_8651,N_7558,N_7159);
or U8652 (N_8652,N_7522,N_7559);
xor U8653 (N_8653,N_7894,N_7799);
or U8654 (N_8654,N_7742,N_7066);
xor U8655 (N_8655,N_7210,N_7943);
or U8656 (N_8656,N_7268,N_7029);
xor U8657 (N_8657,N_7718,N_7753);
or U8658 (N_8658,N_7397,N_7412);
and U8659 (N_8659,N_7201,N_7122);
and U8660 (N_8660,N_7719,N_7029);
and U8661 (N_8661,N_7211,N_7137);
or U8662 (N_8662,N_7754,N_7058);
xor U8663 (N_8663,N_7180,N_7145);
xnor U8664 (N_8664,N_7775,N_7864);
nor U8665 (N_8665,N_7450,N_7857);
or U8666 (N_8666,N_7301,N_7001);
and U8667 (N_8667,N_7068,N_7272);
and U8668 (N_8668,N_7498,N_7298);
nand U8669 (N_8669,N_7628,N_7119);
xor U8670 (N_8670,N_7510,N_7914);
xnor U8671 (N_8671,N_7440,N_7626);
and U8672 (N_8672,N_7860,N_7808);
nor U8673 (N_8673,N_7055,N_7954);
xor U8674 (N_8674,N_7509,N_7201);
nor U8675 (N_8675,N_7514,N_7541);
nor U8676 (N_8676,N_7605,N_7830);
nor U8677 (N_8677,N_7162,N_7647);
and U8678 (N_8678,N_7245,N_7095);
nand U8679 (N_8679,N_7836,N_7179);
or U8680 (N_8680,N_7536,N_7720);
or U8681 (N_8681,N_7857,N_7056);
and U8682 (N_8682,N_7777,N_7910);
or U8683 (N_8683,N_7232,N_7670);
nor U8684 (N_8684,N_7630,N_7426);
and U8685 (N_8685,N_7227,N_7391);
nor U8686 (N_8686,N_7679,N_7310);
nor U8687 (N_8687,N_7120,N_7650);
and U8688 (N_8688,N_7008,N_7491);
nor U8689 (N_8689,N_7225,N_7884);
nand U8690 (N_8690,N_7861,N_7568);
and U8691 (N_8691,N_7508,N_7672);
xnor U8692 (N_8692,N_7471,N_7062);
nand U8693 (N_8693,N_7836,N_7821);
xnor U8694 (N_8694,N_7617,N_7530);
nand U8695 (N_8695,N_7526,N_7158);
xnor U8696 (N_8696,N_7431,N_7239);
xor U8697 (N_8697,N_7270,N_7568);
nand U8698 (N_8698,N_7011,N_7458);
xnor U8699 (N_8699,N_7417,N_7580);
and U8700 (N_8700,N_7155,N_7236);
and U8701 (N_8701,N_7723,N_7809);
xnor U8702 (N_8702,N_7812,N_7791);
nand U8703 (N_8703,N_7366,N_7189);
nor U8704 (N_8704,N_7432,N_7044);
xor U8705 (N_8705,N_7609,N_7230);
or U8706 (N_8706,N_7310,N_7691);
nor U8707 (N_8707,N_7185,N_7007);
nor U8708 (N_8708,N_7434,N_7092);
nor U8709 (N_8709,N_7352,N_7334);
xnor U8710 (N_8710,N_7386,N_7587);
or U8711 (N_8711,N_7276,N_7215);
xor U8712 (N_8712,N_7351,N_7859);
xor U8713 (N_8713,N_7264,N_7727);
and U8714 (N_8714,N_7808,N_7304);
xor U8715 (N_8715,N_7027,N_7495);
and U8716 (N_8716,N_7151,N_7971);
and U8717 (N_8717,N_7107,N_7334);
xor U8718 (N_8718,N_7399,N_7354);
xor U8719 (N_8719,N_7058,N_7248);
xnor U8720 (N_8720,N_7758,N_7991);
nand U8721 (N_8721,N_7993,N_7215);
and U8722 (N_8722,N_7843,N_7436);
nand U8723 (N_8723,N_7841,N_7714);
and U8724 (N_8724,N_7282,N_7680);
xor U8725 (N_8725,N_7259,N_7198);
nand U8726 (N_8726,N_7085,N_7130);
or U8727 (N_8727,N_7586,N_7252);
nor U8728 (N_8728,N_7253,N_7165);
or U8729 (N_8729,N_7157,N_7249);
nor U8730 (N_8730,N_7756,N_7472);
or U8731 (N_8731,N_7815,N_7817);
nand U8732 (N_8732,N_7508,N_7154);
nor U8733 (N_8733,N_7539,N_7264);
nand U8734 (N_8734,N_7138,N_7928);
nor U8735 (N_8735,N_7650,N_7609);
xnor U8736 (N_8736,N_7665,N_7249);
nor U8737 (N_8737,N_7823,N_7273);
nor U8738 (N_8738,N_7286,N_7178);
nor U8739 (N_8739,N_7348,N_7590);
or U8740 (N_8740,N_7892,N_7381);
and U8741 (N_8741,N_7410,N_7905);
xor U8742 (N_8742,N_7767,N_7927);
nor U8743 (N_8743,N_7273,N_7332);
or U8744 (N_8744,N_7755,N_7650);
or U8745 (N_8745,N_7757,N_7740);
xor U8746 (N_8746,N_7143,N_7463);
or U8747 (N_8747,N_7177,N_7418);
and U8748 (N_8748,N_7064,N_7258);
nand U8749 (N_8749,N_7103,N_7257);
or U8750 (N_8750,N_7525,N_7255);
and U8751 (N_8751,N_7352,N_7660);
nor U8752 (N_8752,N_7289,N_7114);
xnor U8753 (N_8753,N_7507,N_7230);
xnor U8754 (N_8754,N_7953,N_7204);
nor U8755 (N_8755,N_7460,N_7048);
nor U8756 (N_8756,N_7489,N_7776);
xor U8757 (N_8757,N_7480,N_7293);
nand U8758 (N_8758,N_7976,N_7186);
nand U8759 (N_8759,N_7503,N_7679);
or U8760 (N_8760,N_7848,N_7826);
xnor U8761 (N_8761,N_7780,N_7997);
nand U8762 (N_8762,N_7676,N_7190);
nand U8763 (N_8763,N_7158,N_7571);
nand U8764 (N_8764,N_7906,N_7591);
and U8765 (N_8765,N_7876,N_7228);
nor U8766 (N_8766,N_7180,N_7419);
and U8767 (N_8767,N_7490,N_7960);
and U8768 (N_8768,N_7078,N_7210);
or U8769 (N_8769,N_7060,N_7211);
nand U8770 (N_8770,N_7447,N_7525);
xor U8771 (N_8771,N_7228,N_7299);
nand U8772 (N_8772,N_7004,N_7077);
or U8773 (N_8773,N_7493,N_7255);
nand U8774 (N_8774,N_7310,N_7996);
nor U8775 (N_8775,N_7003,N_7620);
and U8776 (N_8776,N_7324,N_7373);
or U8777 (N_8777,N_7447,N_7611);
xor U8778 (N_8778,N_7729,N_7362);
or U8779 (N_8779,N_7810,N_7949);
nand U8780 (N_8780,N_7963,N_7805);
nor U8781 (N_8781,N_7897,N_7611);
xor U8782 (N_8782,N_7264,N_7290);
xnor U8783 (N_8783,N_7615,N_7415);
xor U8784 (N_8784,N_7170,N_7997);
and U8785 (N_8785,N_7469,N_7178);
xnor U8786 (N_8786,N_7372,N_7676);
nor U8787 (N_8787,N_7457,N_7924);
and U8788 (N_8788,N_7851,N_7874);
nor U8789 (N_8789,N_7899,N_7598);
nor U8790 (N_8790,N_7242,N_7055);
nor U8791 (N_8791,N_7531,N_7755);
nor U8792 (N_8792,N_7531,N_7633);
xnor U8793 (N_8793,N_7242,N_7241);
or U8794 (N_8794,N_7402,N_7959);
and U8795 (N_8795,N_7508,N_7214);
xor U8796 (N_8796,N_7982,N_7232);
nand U8797 (N_8797,N_7305,N_7189);
and U8798 (N_8798,N_7911,N_7936);
xor U8799 (N_8799,N_7335,N_7031);
nand U8800 (N_8800,N_7772,N_7328);
nor U8801 (N_8801,N_7534,N_7745);
and U8802 (N_8802,N_7963,N_7812);
xnor U8803 (N_8803,N_7124,N_7964);
xor U8804 (N_8804,N_7376,N_7200);
and U8805 (N_8805,N_7559,N_7037);
nor U8806 (N_8806,N_7042,N_7704);
nor U8807 (N_8807,N_7763,N_7307);
xnor U8808 (N_8808,N_7900,N_7339);
nand U8809 (N_8809,N_7964,N_7160);
nor U8810 (N_8810,N_7183,N_7662);
and U8811 (N_8811,N_7262,N_7935);
nand U8812 (N_8812,N_7454,N_7047);
nand U8813 (N_8813,N_7866,N_7917);
xnor U8814 (N_8814,N_7051,N_7819);
or U8815 (N_8815,N_7517,N_7498);
or U8816 (N_8816,N_7470,N_7607);
xor U8817 (N_8817,N_7523,N_7011);
and U8818 (N_8818,N_7782,N_7993);
or U8819 (N_8819,N_7418,N_7818);
xnor U8820 (N_8820,N_7749,N_7715);
nor U8821 (N_8821,N_7194,N_7519);
xor U8822 (N_8822,N_7128,N_7378);
nor U8823 (N_8823,N_7434,N_7063);
nand U8824 (N_8824,N_7700,N_7470);
or U8825 (N_8825,N_7385,N_7143);
nor U8826 (N_8826,N_7452,N_7557);
nand U8827 (N_8827,N_7427,N_7503);
xor U8828 (N_8828,N_7663,N_7944);
nor U8829 (N_8829,N_7708,N_7378);
xnor U8830 (N_8830,N_7830,N_7173);
or U8831 (N_8831,N_7488,N_7974);
and U8832 (N_8832,N_7971,N_7865);
nor U8833 (N_8833,N_7128,N_7066);
and U8834 (N_8834,N_7872,N_7725);
nor U8835 (N_8835,N_7360,N_7403);
nor U8836 (N_8836,N_7519,N_7442);
nand U8837 (N_8837,N_7286,N_7869);
nand U8838 (N_8838,N_7115,N_7210);
nand U8839 (N_8839,N_7331,N_7555);
or U8840 (N_8840,N_7990,N_7524);
xnor U8841 (N_8841,N_7046,N_7845);
nor U8842 (N_8842,N_7432,N_7943);
nor U8843 (N_8843,N_7942,N_7880);
nor U8844 (N_8844,N_7534,N_7149);
or U8845 (N_8845,N_7336,N_7433);
nor U8846 (N_8846,N_7331,N_7683);
or U8847 (N_8847,N_7435,N_7976);
or U8848 (N_8848,N_7626,N_7727);
and U8849 (N_8849,N_7332,N_7922);
nand U8850 (N_8850,N_7908,N_7529);
and U8851 (N_8851,N_7674,N_7219);
nand U8852 (N_8852,N_7900,N_7413);
nor U8853 (N_8853,N_7535,N_7949);
xor U8854 (N_8854,N_7348,N_7860);
and U8855 (N_8855,N_7470,N_7270);
nor U8856 (N_8856,N_7720,N_7442);
or U8857 (N_8857,N_7592,N_7537);
nor U8858 (N_8858,N_7539,N_7638);
nor U8859 (N_8859,N_7701,N_7080);
and U8860 (N_8860,N_7230,N_7361);
xor U8861 (N_8861,N_7590,N_7298);
or U8862 (N_8862,N_7868,N_7357);
nor U8863 (N_8863,N_7235,N_7146);
and U8864 (N_8864,N_7114,N_7116);
nor U8865 (N_8865,N_7321,N_7029);
and U8866 (N_8866,N_7389,N_7024);
nand U8867 (N_8867,N_7307,N_7149);
and U8868 (N_8868,N_7709,N_7028);
or U8869 (N_8869,N_7655,N_7289);
xnor U8870 (N_8870,N_7146,N_7803);
nor U8871 (N_8871,N_7443,N_7551);
or U8872 (N_8872,N_7619,N_7651);
and U8873 (N_8873,N_7010,N_7217);
and U8874 (N_8874,N_7561,N_7063);
xnor U8875 (N_8875,N_7556,N_7636);
nor U8876 (N_8876,N_7392,N_7989);
and U8877 (N_8877,N_7301,N_7666);
or U8878 (N_8878,N_7185,N_7455);
nor U8879 (N_8879,N_7852,N_7597);
nor U8880 (N_8880,N_7752,N_7411);
nand U8881 (N_8881,N_7003,N_7002);
and U8882 (N_8882,N_7093,N_7680);
and U8883 (N_8883,N_7242,N_7854);
nor U8884 (N_8884,N_7919,N_7443);
xor U8885 (N_8885,N_7279,N_7852);
or U8886 (N_8886,N_7259,N_7342);
and U8887 (N_8887,N_7085,N_7455);
nor U8888 (N_8888,N_7217,N_7588);
and U8889 (N_8889,N_7058,N_7656);
nor U8890 (N_8890,N_7454,N_7415);
and U8891 (N_8891,N_7127,N_7179);
and U8892 (N_8892,N_7835,N_7067);
nor U8893 (N_8893,N_7569,N_7133);
nor U8894 (N_8894,N_7987,N_7016);
and U8895 (N_8895,N_7690,N_7992);
or U8896 (N_8896,N_7212,N_7383);
and U8897 (N_8897,N_7558,N_7041);
nor U8898 (N_8898,N_7069,N_7027);
xnor U8899 (N_8899,N_7997,N_7668);
nand U8900 (N_8900,N_7400,N_7824);
xnor U8901 (N_8901,N_7932,N_7107);
and U8902 (N_8902,N_7855,N_7742);
nor U8903 (N_8903,N_7110,N_7869);
nand U8904 (N_8904,N_7691,N_7374);
xnor U8905 (N_8905,N_7045,N_7596);
and U8906 (N_8906,N_7109,N_7123);
nor U8907 (N_8907,N_7832,N_7764);
xor U8908 (N_8908,N_7346,N_7920);
and U8909 (N_8909,N_7488,N_7076);
xnor U8910 (N_8910,N_7431,N_7467);
or U8911 (N_8911,N_7183,N_7164);
nor U8912 (N_8912,N_7416,N_7070);
or U8913 (N_8913,N_7474,N_7206);
nand U8914 (N_8914,N_7845,N_7265);
xnor U8915 (N_8915,N_7748,N_7447);
or U8916 (N_8916,N_7075,N_7257);
and U8917 (N_8917,N_7988,N_7627);
xor U8918 (N_8918,N_7622,N_7947);
nor U8919 (N_8919,N_7864,N_7209);
and U8920 (N_8920,N_7864,N_7549);
and U8921 (N_8921,N_7327,N_7510);
or U8922 (N_8922,N_7264,N_7511);
nor U8923 (N_8923,N_7934,N_7483);
nand U8924 (N_8924,N_7538,N_7316);
and U8925 (N_8925,N_7610,N_7090);
nand U8926 (N_8926,N_7687,N_7203);
and U8927 (N_8927,N_7794,N_7773);
xnor U8928 (N_8928,N_7429,N_7253);
xor U8929 (N_8929,N_7778,N_7888);
nand U8930 (N_8930,N_7550,N_7652);
nor U8931 (N_8931,N_7376,N_7281);
and U8932 (N_8932,N_7204,N_7820);
and U8933 (N_8933,N_7051,N_7410);
xor U8934 (N_8934,N_7847,N_7593);
or U8935 (N_8935,N_7283,N_7167);
nand U8936 (N_8936,N_7413,N_7021);
nand U8937 (N_8937,N_7167,N_7931);
xnor U8938 (N_8938,N_7535,N_7471);
nand U8939 (N_8939,N_7991,N_7152);
xor U8940 (N_8940,N_7296,N_7390);
or U8941 (N_8941,N_7279,N_7316);
nand U8942 (N_8942,N_7200,N_7382);
xnor U8943 (N_8943,N_7910,N_7143);
nor U8944 (N_8944,N_7289,N_7680);
nand U8945 (N_8945,N_7197,N_7845);
or U8946 (N_8946,N_7885,N_7089);
xor U8947 (N_8947,N_7258,N_7629);
or U8948 (N_8948,N_7696,N_7264);
xnor U8949 (N_8949,N_7567,N_7492);
nor U8950 (N_8950,N_7906,N_7847);
and U8951 (N_8951,N_7479,N_7901);
nor U8952 (N_8952,N_7362,N_7265);
xnor U8953 (N_8953,N_7069,N_7461);
nor U8954 (N_8954,N_7846,N_7513);
nor U8955 (N_8955,N_7815,N_7823);
or U8956 (N_8956,N_7599,N_7625);
xor U8957 (N_8957,N_7173,N_7041);
nand U8958 (N_8958,N_7487,N_7847);
and U8959 (N_8959,N_7065,N_7829);
nor U8960 (N_8960,N_7010,N_7331);
or U8961 (N_8961,N_7496,N_7061);
nand U8962 (N_8962,N_7914,N_7901);
nand U8963 (N_8963,N_7506,N_7088);
or U8964 (N_8964,N_7553,N_7351);
or U8965 (N_8965,N_7984,N_7071);
nor U8966 (N_8966,N_7871,N_7623);
or U8967 (N_8967,N_7799,N_7253);
and U8968 (N_8968,N_7119,N_7891);
xor U8969 (N_8969,N_7661,N_7457);
or U8970 (N_8970,N_7832,N_7218);
or U8971 (N_8971,N_7613,N_7793);
or U8972 (N_8972,N_7143,N_7477);
nand U8973 (N_8973,N_7456,N_7304);
xor U8974 (N_8974,N_7775,N_7220);
nand U8975 (N_8975,N_7615,N_7806);
nor U8976 (N_8976,N_7037,N_7915);
and U8977 (N_8977,N_7255,N_7477);
and U8978 (N_8978,N_7256,N_7631);
xor U8979 (N_8979,N_7787,N_7765);
nand U8980 (N_8980,N_7339,N_7154);
xor U8981 (N_8981,N_7901,N_7489);
and U8982 (N_8982,N_7958,N_7021);
and U8983 (N_8983,N_7081,N_7473);
xor U8984 (N_8984,N_7584,N_7590);
or U8985 (N_8985,N_7784,N_7794);
or U8986 (N_8986,N_7599,N_7910);
or U8987 (N_8987,N_7271,N_7728);
and U8988 (N_8988,N_7551,N_7630);
nor U8989 (N_8989,N_7540,N_7326);
nand U8990 (N_8990,N_7880,N_7269);
or U8991 (N_8991,N_7287,N_7929);
xnor U8992 (N_8992,N_7407,N_7968);
nand U8993 (N_8993,N_7238,N_7035);
xnor U8994 (N_8994,N_7200,N_7456);
and U8995 (N_8995,N_7707,N_7188);
nor U8996 (N_8996,N_7148,N_7088);
or U8997 (N_8997,N_7388,N_7477);
xor U8998 (N_8998,N_7858,N_7035);
nand U8999 (N_8999,N_7231,N_7999);
or U9000 (N_9000,N_8937,N_8474);
xor U9001 (N_9001,N_8734,N_8404);
and U9002 (N_9002,N_8019,N_8493);
or U9003 (N_9003,N_8290,N_8747);
xnor U9004 (N_9004,N_8247,N_8731);
xor U9005 (N_9005,N_8720,N_8228);
xor U9006 (N_9006,N_8346,N_8817);
nand U9007 (N_9007,N_8125,N_8451);
xor U9008 (N_9008,N_8210,N_8438);
nor U9009 (N_9009,N_8171,N_8163);
or U9010 (N_9010,N_8291,N_8337);
and U9011 (N_9011,N_8356,N_8636);
and U9012 (N_9012,N_8002,N_8830);
and U9013 (N_9013,N_8053,N_8484);
nor U9014 (N_9014,N_8508,N_8314);
nand U9015 (N_9015,N_8049,N_8539);
or U9016 (N_9016,N_8591,N_8323);
and U9017 (N_9017,N_8032,N_8600);
or U9018 (N_9018,N_8961,N_8098);
nor U9019 (N_9019,N_8864,N_8602);
and U9020 (N_9020,N_8753,N_8453);
nand U9021 (N_9021,N_8728,N_8795);
or U9022 (N_9022,N_8472,N_8899);
or U9023 (N_9023,N_8353,N_8202);
or U9024 (N_9024,N_8796,N_8820);
nor U9025 (N_9025,N_8026,N_8266);
or U9026 (N_9026,N_8471,N_8548);
or U9027 (N_9027,N_8354,N_8216);
and U9028 (N_9028,N_8188,N_8248);
or U9029 (N_9029,N_8803,N_8643);
and U9030 (N_9030,N_8827,N_8856);
nand U9031 (N_9031,N_8117,N_8645);
xnor U9032 (N_9032,N_8811,N_8981);
nor U9033 (N_9033,N_8782,N_8449);
nor U9034 (N_9034,N_8520,N_8271);
or U9035 (N_9035,N_8191,N_8751);
and U9036 (N_9036,N_8040,N_8273);
and U9037 (N_9037,N_8554,N_8615);
or U9038 (N_9038,N_8324,N_8081);
nand U9039 (N_9039,N_8298,N_8208);
xor U9040 (N_9040,N_8141,N_8544);
or U9041 (N_9041,N_8686,N_8009);
xnor U9042 (N_9042,N_8612,N_8244);
and U9043 (N_9043,N_8936,N_8810);
nand U9044 (N_9044,N_8999,N_8183);
xnor U9045 (N_9045,N_8109,N_8322);
and U9046 (N_9046,N_8545,N_8625);
nor U9047 (N_9047,N_8560,N_8572);
nand U9048 (N_9048,N_8714,N_8024);
or U9049 (N_9049,N_8088,N_8789);
and U9050 (N_9050,N_8411,N_8058);
or U9051 (N_9051,N_8589,N_8694);
nor U9052 (N_9052,N_8931,N_8083);
xor U9053 (N_9053,N_8950,N_8985);
nor U9054 (N_9054,N_8061,N_8529);
and U9055 (N_9055,N_8689,N_8569);
xnor U9056 (N_9056,N_8491,N_8166);
xor U9057 (N_9057,N_8003,N_8349);
nor U9058 (N_9058,N_8730,N_8701);
nor U9059 (N_9059,N_8086,N_8194);
and U9060 (N_9060,N_8719,N_8587);
xor U9061 (N_9061,N_8388,N_8558);
nor U9062 (N_9062,N_8433,N_8499);
xnor U9063 (N_9063,N_8492,N_8175);
nor U9064 (N_9064,N_8684,N_8860);
xnor U9065 (N_9065,N_8055,N_8070);
and U9066 (N_9066,N_8829,N_8465);
xor U9067 (N_9067,N_8181,N_8609);
or U9068 (N_9068,N_8561,N_8954);
or U9069 (N_9069,N_8408,N_8564);
nand U9070 (N_9070,N_8599,N_8173);
and U9071 (N_9071,N_8229,N_8749);
nand U9072 (N_9072,N_8987,N_8306);
nor U9073 (N_9073,N_8787,N_8267);
nor U9074 (N_9074,N_8580,N_8697);
nor U9075 (N_9075,N_8104,N_8670);
and U9076 (N_9076,N_8613,N_8847);
and U9077 (N_9077,N_8761,N_8674);
and U9078 (N_9078,N_8716,N_8718);
xor U9079 (N_9079,N_8967,N_8436);
or U9080 (N_9080,N_8938,N_8839);
nand U9081 (N_9081,N_8851,N_8164);
or U9082 (N_9082,N_8087,N_8984);
or U9083 (N_9083,N_8254,N_8755);
and U9084 (N_9084,N_8380,N_8628);
or U9085 (N_9085,N_8340,N_8970);
nor U9086 (N_9086,N_8343,N_8373);
or U9087 (N_9087,N_8547,N_8555);
xnor U9088 (N_9088,N_8148,N_8011);
nand U9089 (N_9089,N_8956,N_8902);
nor U9090 (N_9090,N_8543,N_8176);
xnor U9091 (N_9091,N_8489,N_8246);
nand U9092 (N_9092,N_8533,N_8683);
nand U9093 (N_9093,N_8137,N_8754);
or U9094 (N_9094,N_8966,N_8690);
xnor U9095 (N_9095,N_8868,N_8307);
nor U9096 (N_9096,N_8804,N_8170);
and U9097 (N_9097,N_8387,N_8506);
and U9098 (N_9098,N_8159,N_8382);
nor U9099 (N_9099,N_8583,N_8317);
nor U9100 (N_9100,N_8918,N_8235);
or U9101 (N_9101,N_8769,N_8809);
and U9102 (N_9102,N_8496,N_8319);
or U9103 (N_9103,N_8883,N_8671);
nand U9104 (N_9104,N_8524,N_8022);
or U9105 (N_9105,N_8712,N_8010);
and U9106 (N_9106,N_8124,N_8487);
xor U9107 (N_9107,N_8197,N_8696);
nor U9108 (N_9108,N_8930,N_8515);
xor U9109 (N_9109,N_8080,N_8189);
xor U9110 (N_9110,N_8205,N_8993);
nand U9111 (N_9111,N_8468,N_8403);
and U9112 (N_9112,N_8252,N_8845);
or U9113 (N_9113,N_8917,N_8893);
nor U9114 (N_9114,N_8897,N_8604);
nand U9115 (N_9115,N_8452,N_8635);
nor U9116 (N_9116,N_8103,N_8046);
xor U9117 (N_9117,N_8112,N_8910);
and U9118 (N_9118,N_8834,N_8018);
xnor U9119 (N_9119,N_8959,N_8974);
nand U9120 (N_9120,N_8495,N_8552);
nor U9121 (N_9121,N_8106,N_8100);
nand U9122 (N_9122,N_8700,N_8763);
xor U9123 (N_9123,N_8315,N_8919);
nand U9124 (N_9124,N_8486,N_8299);
nor U9125 (N_9125,N_8001,N_8313);
nand U9126 (N_9126,N_8145,N_8309);
and U9127 (N_9127,N_8578,N_8488);
nor U9128 (N_9128,N_8691,N_8818);
or U9129 (N_9129,N_8146,N_8178);
xnor U9130 (N_9130,N_8446,N_8607);
nand U9131 (N_9131,N_8000,N_8998);
nor U9132 (N_9132,N_8633,N_8051);
or U9133 (N_9133,N_8951,N_8126);
or U9134 (N_9134,N_8370,N_8581);
xor U9135 (N_9135,N_8321,N_8814);
and U9136 (N_9136,N_8614,N_8756);
nor U9137 (N_9137,N_8375,N_8287);
nor U9138 (N_9138,N_8085,N_8479);
xnor U9139 (N_9139,N_8733,N_8577);
nand U9140 (N_9140,N_8417,N_8477);
or U9141 (N_9141,N_8646,N_8182);
xnor U9142 (N_9142,N_8652,N_8147);
or U9143 (N_9143,N_8603,N_8360);
nor U9144 (N_9144,N_8835,N_8185);
or U9145 (N_9145,N_8757,N_8187);
or U9146 (N_9146,N_8736,N_8741);
or U9147 (N_9147,N_8036,N_8160);
or U9148 (N_9148,N_8485,N_8406);
and U9149 (N_9149,N_8157,N_8294);
nand U9150 (N_9150,N_8074,N_8791);
and U9151 (N_9151,N_8685,N_8447);
xnor U9152 (N_9152,N_8828,N_8792);
and U9153 (N_9153,N_8677,N_8429);
and U9154 (N_9154,N_8859,N_8768);
xnor U9155 (N_9155,N_8457,N_8698);
nor U9156 (N_9156,N_8812,N_8132);
or U9157 (N_9157,N_8213,N_8348);
and U9158 (N_9158,N_8089,N_8470);
nor U9159 (N_9159,N_8710,N_8220);
and U9160 (N_9160,N_8546,N_8441);
nor U9161 (N_9161,N_8758,N_8881);
xor U9162 (N_9162,N_8608,N_8898);
or U9163 (N_9163,N_8932,N_8318);
and U9164 (N_9164,N_8156,N_8034);
or U9165 (N_9165,N_8443,N_8084);
and U9166 (N_9166,N_8655,N_8415);
nand U9167 (N_9167,N_8878,N_8177);
nor U9168 (N_9168,N_8855,N_8514);
nor U9169 (N_9169,N_8102,N_8507);
and U9170 (N_9170,N_8704,N_8234);
xnor U9171 (N_9171,N_8301,N_8707);
nand U9172 (N_9172,N_8639,N_8190);
xor U9173 (N_9173,N_8432,N_8651);
or U9174 (N_9174,N_8043,N_8798);
xor U9175 (N_9175,N_8550,N_8774);
xnor U9176 (N_9176,N_8045,N_8342);
and U9177 (N_9177,N_8647,N_8218);
or U9178 (N_9178,N_8350,N_8393);
or U9179 (N_9179,N_8588,N_8551);
xnor U9180 (N_9180,N_8584,N_8838);
nand U9181 (N_9181,N_8631,N_8161);
xor U9182 (N_9182,N_8502,N_8371);
xnor U9183 (N_9183,N_8624,N_8662);
or U9184 (N_9184,N_8421,N_8642);
nor U9185 (N_9185,N_8900,N_8179);
or U9186 (N_9186,N_8279,N_8044);
and U9187 (N_9187,N_8896,N_8894);
nand U9188 (N_9188,N_8225,N_8122);
xor U9189 (N_9189,N_8933,N_8861);
nor U9190 (N_9190,N_8922,N_8399);
and U9191 (N_9191,N_8195,N_8152);
nand U9192 (N_9192,N_8420,N_8935);
or U9193 (N_9193,N_8873,N_8767);
nor U9194 (N_9194,N_8735,N_8724);
nor U9195 (N_9195,N_8014,N_8131);
or U9196 (N_9196,N_8882,N_8217);
and U9197 (N_9197,N_8243,N_8473);
nor U9198 (N_9198,N_8801,N_8364);
nand U9199 (N_9199,N_8312,N_8067);
xor U9200 (N_9200,N_8511,N_8017);
nor U9201 (N_9201,N_8331,N_8211);
or U9202 (N_9202,N_8027,N_8732);
xor U9203 (N_9203,N_8250,N_8605);
or U9204 (N_9204,N_8108,N_8887);
nand U9205 (N_9205,N_8326,N_8585);
or U9206 (N_9206,N_8392,N_8991);
nand U9207 (N_9207,N_8850,N_8711);
or U9208 (N_9208,N_8316,N_8778);
nor U9209 (N_9209,N_8852,N_8562);
and U9210 (N_9210,N_8806,N_8596);
or U9211 (N_9211,N_8021,N_8105);
nor U9212 (N_9212,N_8142,N_8862);
nor U9213 (N_9213,N_8286,N_8007);
nand U9214 (N_9214,N_8214,N_8542);
nor U9215 (N_9215,N_8407,N_8903);
xor U9216 (N_9216,N_8586,N_8526);
xor U9217 (N_9217,N_8110,N_8888);
xnor U9218 (N_9218,N_8119,N_8345);
xnor U9219 (N_9219,N_8831,N_8260);
xor U9220 (N_9220,N_8426,N_8750);
nand U9221 (N_9221,N_8460,N_8962);
nor U9222 (N_9222,N_8875,N_8475);
or U9223 (N_9223,N_8944,N_8076);
and U9224 (N_9224,N_8934,N_8781);
xor U9225 (N_9225,N_8527,N_8239);
or U9226 (N_9226,N_8050,N_8952);
nand U9227 (N_9227,N_8872,N_8198);
nor U9228 (N_9228,N_8302,N_8169);
xor U9229 (N_9229,N_8971,N_8006);
xnor U9230 (N_9230,N_8069,N_8759);
nor U9231 (N_9231,N_8630,N_8275);
and U9232 (N_9232,N_8965,N_8154);
and U9233 (N_9233,N_8231,N_8238);
or U9234 (N_9234,N_8269,N_8245);
or U9235 (N_9235,N_8430,N_8400);
xor U9236 (N_9236,N_8155,N_8620);
and U9237 (N_9237,N_8192,N_8553);
xor U9238 (N_9238,N_8826,N_8448);
nand U9239 (N_9239,N_8120,N_8300);
nand U9240 (N_9240,N_8595,N_8390);
and U9241 (N_9241,N_8992,N_8740);
or U9242 (N_9242,N_8540,N_8770);
and U9243 (N_9243,N_8994,N_8303);
and U9244 (N_9244,N_8840,N_8090);
nor U9245 (N_9245,N_8619,N_8819);
xor U9246 (N_9246,N_8258,N_8361);
nor U9247 (N_9247,N_8101,N_8920);
xnor U9248 (N_9248,N_8706,N_8115);
nand U9249 (N_9249,N_8895,N_8632);
xor U9250 (N_9250,N_8232,N_8909);
nand U9251 (N_9251,N_8212,N_8982);
or U9252 (N_9252,N_8901,N_8359);
nand U9253 (N_9253,N_8012,N_8270);
nor U9254 (N_9254,N_8648,N_8140);
nor U9255 (N_9255,N_8825,N_8413);
nor U9256 (N_9256,N_8530,N_8478);
and U9257 (N_9257,N_8111,N_8093);
nand U9258 (N_9258,N_8841,N_8094);
nand U9259 (N_9259,N_8374,N_8737);
xnor U9260 (N_9260,N_8594,N_8510);
or U9261 (N_9261,N_8644,N_8573);
xor U9262 (N_9262,N_8422,N_8699);
or U9263 (N_9263,N_8016,N_8005);
xor U9264 (N_9264,N_8242,N_8945);
and U9265 (N_9265,N_8365,N_8305);
or U9266 (N_9266,N_8256,N_8459);
and U9267 (N_9267,N_8531,N_8114);
nor U9268 (N_9268,N_8601,N_8066);
nand U9269 (N_9269,N_8654,N_8536);
or U9270 (N_9270,N_8611,N_8667);
nor U9271 (N_9271,N_8023,N_8249);
and U9272 (N_9272,N_8263,N_8219);
and U9273 (N_9273,N_8889,N_8236);
and U9274 (N_9274,N_8742,N_8802);
nand U9275 (N_9275,N_8230,N_8186);
nand U9276 (N_9276,N_8516,N_8138);
or U9277 (N_9277,N_8963,N_8566);
nor U9278 (N_9278,N_8385,N_8772);
nand U9279 (N_9279,N_8541,N_8418);
xor U9280 (N_9280,N_8693,N_8377);
or U9281 (N_9281,N_8462,N_8505);
xor U9282 (N_9282,N_8983,N_8790);
and U9283 (N_9283,N_8854,N_8281);
nand U9284 (N_9284,N_8869,N_8015);
xor U9285 (N_9285,N_8977,N_8501);
xor U9286 (N_9286,N_8203,N_8261);
nor U9287 (N_9287,N_8622,N_8297);
or U9288 (N_9288,N_8989,N_8092);
nand U9289 (N_9289,N_8968,N_8362);
or U9290 (N_9290,N_8091,N_8412);
nor U9291 (N_9291,N_8037,N_8455);
nor U9292 (N_9292,N_8064,N_8174);
or U9293 (N_9293,N_8785,N_8773);
nand U9294 (N_9294,N_8033,N_8383);
and U9295 (N_9295,N_8638,N_8660);
nand U9296 (N_9296,N_8549,N_8409);
and U9297 (N_9297,N_8884,N_8357);
nand U9298 (N_9298,N_8890,N_8870);
nand U9299 (N_9299,N_8130,N_8942);
nor U9300 (N_9300,N_8634,N_8571);
and U9301 (N_9301,N_8597,N_8042);
nand U9302 (N_9302,N_8363,N_8347);
or U9303 (N_9303,N_8669,N_8771);
or U9304 (N_9304,N_8445,N_8762);
and U9305 (N_9305,N_8863,N_8574);
xor U9306 (N_9306,N_8657,N_8973);
or U9307 (N_9307,N_8004,N_8209);
nor U9308 (N_9308,N_8240,N_8456);
or U9309 (N_9309,N_8886,N_8498);
and U9310 (N_9310,N_8518,N_8367);
and U9311 (N_9311,N_8410,N_8915);
and U9312 (N_9312,N_8149,N_8593);
or U9313 (N_9313,N_8416,N_8262);
or U9314 (N_9314,N_8206,N_8077);
xor U9315 (N_9315,N_8955,N_8320);
nand U9316 (N_9316,N_8439,N_8059);
or U9317 (N_9317,N_8695,N_8062);
nand U9318 (N_9318,N_8675,N_8682);
or U9319 (N_9319,N_8525,N_8912);
and U9320 (N_9320,N_8681,N_8640);
nor U9321 (N_9321,N_8853,N_8723);
nor U9322 (N_9322,N_8797,N_8929);
nand U9323 (N_9323,N_8904,N_8168);
nand U9324 (N_9324,N_8738,N_8143);
or U9325 (N_9325,N_8776,N_8123);
or U9326 (N_9326,N_8128,N_8162);
nor U9327 (N_9327,N_8133,N_8204);
and U9328 (N_9328,N_8095,N_8423);
xnor U9329 (N_9329,N_8729,N_8995);
or U9330 (N_9330,N_8394,N_8874);
and U9331 (N_9331,N_8858,N_8978);
xor U9332 (N_9332,N_8031,N_8121);
xor U9333 (N_9333,N_8268,N_8029);
nor U9334 (N_9334,N_8490,N_8226);
nor U9335 (N_9335,N_8025,N_8512);
xor U9336 (N_9336,N_8284,N_8866);
nor U9337 (N_9337,N_8038,N_8867);
xor U9338 (N_9338,N_8107,N_8964);
nand U9339 (N_9339,N_8435,N_8567);
and U9340 (N_9340,N_8292,N_8172);
nor U9341 (N_9341,N_8405,N_8833);
nor U9342 (N_9342,N_8442,N_8521);
nor U9343 (N_9343,N_8805,N_8799);
and U9344 (N_9344,N_8215,N_8150);
xnor U9345 (N_9345,N_8463,N_8030);
nand U9346 (N_9346,N_8783,N_8891);
or U9347 (N_9347,N_8779,N_8708);
or U9348 (N_9348,N_8253,N_8280);
nor U9349 (N_9349,N_8293,N_8715);
and U9350 (N_9350,N_8672,N_8200);
xor U9351 (N_9351,N_8800,N_8816);
nand U9352 (N_9352,N_8264,N_8467);
nor U9353 (N_9353,N_8713,N_8285);
nor U9354 (N_9354,N_8621,N_8310);
xnor U9355 (N_9355,N_8913,N_8338);
xor U9356 (N_9356,N_8047,N_8461);
or U9357 (N_9357,N_8135,N_8822);
xnor U9358 (N_9358,N_8905,N_8788);
nor U9359 (N_9359,N_8389,N_8165);
nor U9360 (N_9360,N_8519,N_8656);
and U9361 (N_9361,N_8241,N_8274);
and U9362 (N_9362,N_8289,N_8760);
xor U9363 (N_9363,N_8946,N_8748);
nand U9364 (N_9364,N_8118,N_8641);
and U9365 (N_9365,N_8048,N_8391);
nand U9366 (N_9366,N_8237,N_8916);
nand U9367 (N_9367,N_8673,N_8764);
nand U9368 (N_9368,N_8368,N_8666);
nand U9369 (N_9369,N_8440,N_8617);
nand U9370 (N_9370,N_8606,N_8134);
nand U9371 (N_9371,N_8687,N_8509);
nand U9372 (N_9372,N_8196,N_8227);
or U9373 (N_9373,N_8907,N_8953);
or U9374 (N_9374,N_8351,N_8568);
nor U9375 (N_9375,N_8923,N_8610);
or U9376 (N_9376,N_8892,N_8464);
nand U9377 (N_9377,N_8914,N_8688);
nand U9378 (N_9378,N_8592,N_8582);
xnor U9379 (N_9379,N_8482,N_8557);
nor U9380 (N_9380,N_8824,N_8793);
and U9381 (N_9381,N_8665,N_8381);
nand U9382 (N_9382,N_8949,N_8637);
nand U9383 (N_9383,N_8846,N_8207);
nand U9384 (N_9384,N_8650,N_8065);
nor U9385 (N_9385,N_8096,N_8997);
and U9386 (N_9386,N_8054,N_8837);
xor U9387 (N_9387,N_8726,N_8288);
or U9388 (N_9388,N_8616,N_8328);
nand U9389 (N_9389,N_8127,N_8481);
nand U9390 (N_9390,N_8376,N_8575);
or U9391 (N_9391,N_8522,N_8099);
and U9392 (N_9392,N_8259,N_8958);
xnor U9393 (N_9393,N_8379,N_8927);
and U9394 (N_9394,N_8336,N_8908);
or U9395 (N_9395,N_8703,N_8702);
and U9396 (N_9396,N_8466,N_8794);
or U9397 (N_9397,N_8335,N_8559);
or U9398 (N_9398,N_8765,N_8570);
nor U9399 (N_9399,N_8957,N_8784);
nand U9400 (N_9400,N_8330,N_8948);
nand U9401 (N_9401,N_8590,N_8849);
or U9402 (N_9402,N_8283,N_8813);
nor U9403 (N_9403,N_8073,N_8661);
nand U9404 (N_9404,N_8960,N_8517);
and U9405 (N_9405,N_8692,N_8871);
and U9406 (N_9406,N_8668,N_8535);
or U9407 (N_9407,N_8251,N_8402);
and U9408 (N_9408,N_8663,N_8969);
or U9409 (N_9409,N_8911,N_8068);
nor U9410 (N_9410,N_8311,N_8151);
nand U9411 (N_9411,N_8180,N_8020);
nor U9412 (N_9412,N_8184,N_8678);
nand U9413 (N_9413,N_8523,N_8906);
xor U9414 (N_9414,N_8339,N_8384);
xor U9415 (N_9415,N_8325,N_8943);
nor U9416 (N_9416,N_8424,N_8780);
and U9417 (N_9417,N_8265,N_8534);
and U9418 (N_9418,N_8352,N_8082);
and U9419 (N_9419,N_8947,N_8513);
or U9420 (N_9420,N_8623,N_8885);
xnor U9421 (N_9421,N_8832,N_8556);
nand U9422 (N_9422,N_8329,N_8928);
nand U9423 (N_9423,N_8295,N_8414);
or U9424 (N_9424,N_8679,N_8139);
or U9425 (N_9425,N_8334,N_8664);
or U9426 (N_9426,N_8745,N_8308);
xnor U9427 (N_9427,N_8113,N_8427);
nand U9428 (N_9428,N_8836,N_8848);
or U9429 (N_9429,N_8497,N_8476);
xor U9430 (N_9430,N_8052,N_8876);
nor U9431 (N_9431,N_8976,N_8941);
nor U9432 (N_9432,N_8158,N_8167);
nor U9433 (N_9433,N_8815,N_8437);
nor U9434 (N_9434,N_8395,N_8786);
nand U9435 (N_9435,N_8344,N_8727);
or U9436 (N_9436,N_8221,N_8940);
and U9437 (N_9437,N_8709,N_8972);
xor U9438 (N_9438,N_8717,N_8705);
nand U9439 (N_9439,N_8565,N_8277);
or U9440 (N_9440,N_8013,N_8450);
nor U9441 (N_9441,N_8939,N_8746);
and U9442 (N_9442,N_8223,N_8454);
xnor U9443 (N_9443,N_8041,N_8458);
xor U9444 (N_9444,N_8056,N_8035);
or U9445 (N_9445,N_8743,N_8807);
xor U9446 (N_9446,N_8378,N_8879);
nor U9447 (N_9447,N_8332,N_8257);
and U9448 (N_9448,N_8877,N_8008);
xnor U9449 (N_9449,N_8079,N_8649);
nor U9450 (N_9450,N_8372,N_8304);
or U9451 (N_9451,N_8658,N_8428);
nor U9452 (N_9452,N_8333,N_8282);
nor U9453 (N_9453,N_8193,N_8136);
or U9454 (N_9454,N_8469,N_8341);
or U9455 (N_9455,N_8752,N_8725);
nand U9456 (N_9456,N_8224,N_8659);
xor U9457 (N_9457,N_8296,N_8653);
nor U9458 (N_9458,N_8996,N_8823);
or U9459 (N_9459,N_8057,N_8028);
nand U9460 (N_9460,N_8366,N_8480);
nor U9461 (N_9461,N_8201,N_8865);
xnor U9462 (N_9462,N_8097,N_8975);
nor U9463 (N_9463,N_8627,N_8071);
and U9464 (N_9464,N_8039,N_8739);
or U9465 (N_9465,N_8494,N_8144);
or U9466 (N_9466,N_8926,N_8434);
xnor U9467 (N_9467,N_8222,N_8386);
nand U9468 (N_9468,N_8598,N_8925);
and U9469 (N_9469,N_8444,N_8880);
and U9470 (N_9470,N_8327,N_8680);
nor U9471 (N_9471,N_8777,N_8821);
nand U9472 (N_9472,N_8921,N_8116);
and U9473 (N_9473,N_8538,N_8990);
nor U9474 (N_9474,N_8844,N_8072);
xnor U9475 (N_9475,N_8808,N_8060);
and U9476 (N_9476,N_8857,N_8629);
and U9477 (N_9477,N_8078,N_8766);
xor U9478 (N_9478,N_8278,N_8626);
nand U9479 (N_9479,N_8483,N_8355);
and U9480 (N_9480,N_8419,N_8924);
nand U9481 (N_9481,N_8576,N_8425);
xnor U9482 (N_9482,N_8276,N_8986);
xnor U9483 (N_9483,N_8843,N_8722);
nor U9484 (N_9484,N_8579,N_8398);
or U9485 (N_9485,N_8721,N_8075);
or U9486 (N_9486,N_8153,N_8988);
or U9487 (N_9487,N_8528,N_8532);
nand U9488 (N_9488,N_8063,N_8676);
xnor U9489 (N_9489,N_8431,N_8358);
xnor U9490 (N_9490,N_8980,N_8369);
nor U9491 (N_9491,N_8842,N_8618);
or U9492 (N_9492,N_8744,N_8979);
and U9493 (N_9493,N_8775,N_8397);
nor U9494 (N_9494,N_8504,N_8503);
nor U9495 (N_9495,N_8233,N_8255);
xor U9496 (N_9496,N_8537,N_8272);
xnor U9497 (N_9497,N_8500,N_8129);
nand U9498 (N_9498,N_8199,N_8396);
nor U9499 (N_9499,N_8401,N_8563);
xor U9500 (N_9500,N_8730,N_8739);
nor U9501 (N_9501,N_8402,N_8236);
nand U9502 (N_9502,N_8535,N_8063);
nand U9503 (N_9503,N_8855,N_8371);
or U9504 (N_9504,N_8138,N_8189);
xor U9505 (N_9505,N_8434,N_8270);
and U9506 (N_9506,N_8077,N_8154);
nor U9507 (N_9507,N_8040,N_8943);
or U9508 (N_9508,N_8636,N_8531);
xor U9509 (N_9509,N_8244,N_8214);
or U9510 (N_9510,N_8734,N_8785);
and U9511 (N_9511,N_8889,N_8379);
or U9512 (N_9512,N_8982,N_8996);
nor U9513 (N_9513,N_8970,N_8067);
xnor U9514 (N_9514,N_8931,N_8994);
xnor U9515 (N_9515,N_8115,N_8217);
and U9516 (N_9516,N_8625,N_8876);
nand U9517 (N_9517,N_8324,N_8452);
nand U9518 (N_9518,N_8402,N_8943);
nor U9519 (N_9519,N_8581,N_8620);
or U9520 (N_9520,N_8039,N_8311);
nand U9521 (N_9521,N_8211,N_8439);
nand U9522 (N_9522,N_8000,N_8829);
and U9523 (N_9523,N_8601,N_8184);
or U9524 (N_9524,N_8378,N_8040);
nor U9525 (N_9525,N_8319,N_8842);
or U9526 (N_9526,N_8289,N_8978);
xnor U9527 (N_9527,N_8575,N_8638);
xnor U9528 (N_9528,N_8685,N_8702);
nand U9529 (N_9529,N_8642,N_8710);
nor U9530 (N_9530,N_8716,N_8261);
xnor U9531 (N_9531,N_8156,N_8663);
or U9532 (N_9532,N_8586,N_8116);
and U9533 (N_9533,N_8373,N_8565);
nand U9534 (N_9534,N_8218,N_8682);
and U9535 (N_9535,N_8940,N_8043);
and U9536 (N_9536,N_8715,N_8093);
and U9537 (N_9537,N_8607,N_8214);
and U9538 (N_9538,N_8519,N_8551);
and U9539 (N_9539,N_8642,N_8817);
and U9540 (N_9540,N_8102,N_8696);
xnor U9541 (N_9541,N_8786,N_8011);
nor U9542 (N_9542,N_8045,N_8626);
xor U9543 (N_9543,N_8402,N_8573);
and U9544 (N_9544,N_8813,N_8095);
or U9545 (N_9545,N_8430,N_8625);
and U9546 (N_9546,N_8840,N_8595);
nand U9547 (N_9547,N_8984,N_8077);
or U9548 (N_9548,N_8292,N_8897);
or U9549 (N_9549,N_8536,N_8052);
nor U9550 (N_9550,N_8228,N_8327);
nor U9551 (N_9551,N_8240,N_8463);
nor U9552 (N_9552,N_8502,N_8600);
and U9553 (N_9553,N_8401,N_8606);
or U9554 (N_9554,N_8947,N_8666);
nand U9555 (N_9555,N_8321,N_8008);
and U9556 (N_9556,N_8531,N_8051);
xnor U9557 (N_9557,N_8683,N_8667);
nor U9558 (N_9558,N_8452,N_8602);
nand U9559 (N_9559,N_8104,N_8056);
xor U9560 (N_9560,N_8463,N_8714);
nand U9561 (N_9561,N_8628,N_8007);
nor U9562 (N_9562,N_8152,N_8659);
xnor U9563 (N_9563,N_8310,N_8164);
and U9564 (N_9564,N_8504,N_8023);
xnor U9565 (N_9565,N_8308,N_8675);
nand U9566 (N_9566,N_8978,N_8035);
and U9567 (N_9567,N_8593,N_8444);
nand U9568 (N_9568,N_8639,N_8312);
nor U9569 (N_9569,N_8612,N_8414);
or U9570 (N_9570,N_8543,N_8105);
or U9571 (N_9571,N_8378,N_8589);
nor U9572 (N_9572,N_8541,N_8618);
nand U9573 (N_9573,N_8894,N_8046);
or U9574 (N_9574,N_8326,N_8361);
or U9575 (N_9575,N_8600,N_8559);
xnor U9576 (N_9576,N_8248,N_8166);
xor U9577 (N_9577,N_8029,N_8924);
nor U9578 (N_9578,N_8568,N_8453);
xnor U9579 (N_9579,N_8096,N_8279);
xnor U9580 (N_9580,N_8260,N_8453);
or U9581 (N_9581,N_8952,N_8052);
xnor U9582 (N_9582,N_8870,N_8456);
and U9583 (N_9583,N_8342,N_8512);
nor U9584 (N_9584,N_8485,N_8276);
and U9585 (N_9585,N_8930,N_8270);
nand U9586 (N_9586,N_8077,N_8771);
and U9587 (N_9587,N_8027,N_8423);
and U9588 (N_9588,N_8141,N_8571);
xor U9589 (N_9589,N_8980,N_8057);
and U9590 (N_9590,N_8815,N_8424);
nand U9591 (N_9591,N_8865,N_8204);
or U9592 (N_9592,N_8016,N_8135);
nor U9593 (N_9593,N_8735,N_8625);
or U9594 (N_9594,N_8620,N_8762);
nand U9595 (N_9595,N_8456,N_8598);
and U9596 (N_9596,N_8463,N_8877);
xnor U9597 (N_9597,N_8206,N_8739);
nor U9598 (N_9598,N_8671,N_8815);
xor U9599 (N_9599,N_8233,N_8891);
or U9600 (N_9600,N_8614,N_8383);
or U9601 (N_9601,N_8152,N_8365);
and U9602 (N_9602,N_8231,N_8082);
and U9603 (N_9603,N_8808,N_8884);
nand U9604 (N_9604,N_8854,N_8948);
xnor U9605 (N_9605,N_8371,N_8737);
xor U9606 (N_9606,N_8383,N_8821);
nand U9607 (N_9607,N_8666,N_8239);
and U9608 (N_9608,N_8332,N_8680);
nor U9609 (N_9609,N_8370,N_8165);
nand U9610 (N_9610,N_8624,N_8687);
nand U9611 (N_9611,N_8927,N_8213);
or U9612 (N_9612,N_8647,N_8968);
xnor U9613 (N_9613,N_8566,N_8452);
nand U9614 (N_9614,N_8739,N_8554);
and U9615 (N_9615,N_8851,N_8236);
xnor U9616 (N_9616,N_8054,N_8739);
nand U9617 (N_9617,N_8950,N_8514);
nor U9618 (N_9618,N_8620,N_8307);
nand U9619 (N_9619,N_8542,N_8660);
and U9620 (N_9620,N_8691,N_8528);
nand U9621 (N_9621,N_8797,N_8216);
and U9622 (N_9622,N_8371,N_8382);
xnor U9623 (N_9623,N_8241,N_8531);
xor U9624 (N_9624,N_8561,N_8620);
nor U9625 (N_9625,N_8931,N_8187);
or U9626 (N_9626,N_8390,N_8984);
and U9627 (N_9627,N_8000,N_8542);
nand U9628 (N_9628,N_8899,N_8867);
nor U9629 (N_9629,N_8995,N_8461);
or U9630 (N_9630,N_8801,N_8498);
and U9631 (N_9631,N_8644,N_8560);
xor U9632 (N_9632,N_8256,N_8194);
nand U9633 (N_9633,N_8891,N_8672);
nor U9634 (N_9634,N_8613,N_8536);
nand U9635 (N_9635,N_8635,N_8351);
or U9636 (N_9636,N_8885,N_8382);
nand U9637 (N_9637,N_8755,N_8408);
and U9638 (N_9638,N_8290,N_8730);
nand U9639 (N_9639,N_8264,N_8561);
nor U9640 (N_9640,N_8212,N_8791);
xor U9641 (N_9641,N_8857,N_8611);
xnor U9642 (N_9642,N_8526,N_8205);
and U9643 (N_9643,N_8911,N_8767);
nor U9644 (N_9644,N_8013,N_8351);
or U9645 (N_9645,N_8405,N_8547);
xnor U9646 (N_9646,N_8902,N_8390);
and U9647 (N_9647,N_8219,N_8268);
and U9648 (N_9648,N_8017,N_8719);
xor U9649 (N_9649,N_8782,N_8221);
or U9650 (N_9650,N_8101,N_8159);
nand U9651 (N_9651,N_8780,N_8975);
nor U9652 (N_9652,N_8010,N_8367);
nand U9653 (N_9653,N_8241,N_8277);
nor U9654 (N_9654,N_8112,N_8517);
or U9655 (N_9655,N_8458,N_8459);
or U9656 (N_9656,N_8246,N_8757);
and U9657 (N_9657,N_8855,N_8584);
nor U9658 (N_9658,N_8885,N_8440);
nor U9659 (N_9659,N_8070,N_8325);
nor U9660 (N_9660,N_8515,N_8093);
nand U9661 (N_9661,N_8634,N_8896);
nand U9662 (N_9662,N_8975,N_8739);
or U9663 (N_9663,N_8148,N_8178);
nor U9664 (N_9664,N_8077,N_8280);
and U9665 (N_9665,N_8922,N_8698);
nand U9666 (N_9666,N_8416,N_8312);
or U9667 (N_9667,N_8305,N_8860);
and U9668 (N_9668,N_8413,N_8086);
and U9669 (N_9669,N_8324,N_8849);
xnor U9670 (N_9670,N_8592,N_8167);
xnor U9671 (N_9671,N_8737,N_8498);
or U9672 (N_9672,N_8960,N_8135);
nor U9673 (N_9673,N_8179,N_8831);
xnor U9674 (N_9674,N_8900,N_8951);
nand U9675 (N_9675,N_8886,N_8188);
nor U9676 (N_9676,N_8582,N_8066);
xor U9677 (N_9677,N_8067,N_8394);
and U9678 (N_9678,N_8136,N_8312);
nor U9679 (N_9679,N_8938,N_8735);
or U9680 (N_9680,N_8080,N_8375);
xor U9681 (N_9681,N_8094,N_8173);
and U9682 (N_9682,N_8397,N_8760);
or U9683 (N_9683,N_8940,N_8215);
xor U9684 (N_9684,N_8864,N_8873);
nor U9685 (N_9685,N_8958,N_8427);
xnor U9686 (N_9686,N_8952,N_8817);
xor U9687 (N_9687,N_8838,N_8278);
nand U9688 (N_9688,N_8879,N_8913);
and U9689 (N_9689,N_8873,N_8081);
nor U9690 (N_9690,N_8031,N_8531);
xnor U9691 (N_9691,N_8568,N_8363);
nand U9692 (N_9692,N_8303,N_8402);
nor U9693 (N_9693,N_8083,N_8900);
nor U9694 (N_9694,N_8835,N_8664);
or U9695 (N_9695,N_8774,N_8860);
nand U9696 (N_9696,N_8953,N_8355);
or U9697 (N_9697,N_8198,N_8705);
or U9698 (N_9698,N_8264,N_8564);
nand U9699 (N_9699,N_8219,N_8790);
nor U9700 (N_9700,N_8974,N_8329);
nor U9701 (N_9701,N_8405,N_8366);
xor U9702 (N_9702,N_8330,N_8235);
or U9703 (N_9703,N_8178,N_8593);
nand U9704 (N_9704,N_8496,N_8279);
xor U9705 (N_9705,N_8007,N_8443);
xnor U9706 (N_9706,N_8462,N_8739);
nand U9707 (N_9707,N_8333,N_8677);
and U9708 (N_9708,N_8763,N_8548);
nor U9709 (N_9709,N_8915,N_8805);
and U9710 (N_9710,N_8739,N_8231);
or U9711 (N_9711,N_8013,N_8426);
or U9712 (N_9712,N_8678,N_8160);
nand U9713 (N_9713,N_8675,N_8595);
or U9714 (N_9714,N_8802,N_8383);
nor U9715 (N_9715,N_8611,N_8803);
xor U9716 (N_9716,N_8690,N_8926);
or U9717 (N_9717,N_8804,N_8428);
or U9718 (N_9718,N_8387,N_8605);
xor U9719 (N_9719,N_8964,N_8132);
and U9720 (N_9720,N_8452,N_8165);
nand U9721 (N_9721,N_8620,N_8074);
xnor U9722 (N_9722,N_8323,N_8732);
nor U9723 (N_9723,N_8942,N_8931);
and U9724 (N_9724,N_8162,N_8571);
xor U9725 (N_9725,N_8836,N_8475);
nor U9726 (N_9726,N_8689,N_8505);
nor U9727 (N_9727,N_8400,N_8946);
nand U9728 (N_9728,N_8632,N_8511);
nand U9729 (N_9729,N_8767,N_8309);
nor U9730 (N_9730,N_8369,N_8715);
nand U9731 (N_9731,N_8985,N_8091);
and U9732 (N_9732,N_8275,N_8160);
nor U9733 (N_9733,N_8991,N_8934);
and U9734 (N_9734,N_8735,N_8910);
nor U9735 (N_9735,N_8429,N_8840);
nor U9736 (N_9736,N_8135,N_8346);
nor U9737 (N_9737,N_8110,N_8714);
or U9738 (N_9738,N_8387,N_8691);
nand U9739 (N_9739,N_8160,N_8007);
xor U9740 (N_9740,N_8512,N_8142);
nor U9741 (N_9741,N_8287,N_8810);
nor U9742 (N_9742,N_8087,N_8361);
nand U9743 (N_9743,N_8474,N_8123);
and U9744 (N_9744,N_8834,N_8811);
xor U9745 (N_9745,N_8488,N_8684);
nor U9746 (N_9746,N_8044,N_8382);
nand U9747 (N_9747,N_8763,N_8556);
xor U9748 (N_9748,N_8281,N_8591);
nor U9749 (N_9749,N_8565,N_8834);
and U9750 (N_9750,N_8503,N_8299);
xnor U9751 (N_9751,N_8035,N_8481);
nor U9752 (N_9752,N_8928,N_8663);
xnor U9753 (N_9753,N_8017,N_8902);
nor U9754 (N_9754,N_8159,N_8140);
nand U9755 (N_9755,N_8088,N_8587);
xnor U9756 (N_9756,N_8358,N_8702);
nand U9757 (N_9757,N_8824,N_8840);
or U9758 (N_9758,N_8627,N_8901);
nor U9759 (N_9759,N_8955,N_8951);
or U9760 (N_9760,N_8692,N_8445);
nand U9761 (N_9761,N_8860,N_8322);
nand U9762 (N_9762,N_8063,N_8304);
nor U9763 (N_9763,N_8726,N_8927);
nor U9764 (N_9764,N_8409,N_8189);
nand U9765 (N_9765,N_8138,N_8077);
or U9766 (N_9766,N_8073,N_8452);
or U9767 (N_9767,N_8023,N_8372);
xor U9768 (N_9768,N_8784,N_8998);
xor U9769 (N_9769,N_8081,N_8555);
xnor U9770 (N_9770,N_8819,N_8988);
nor U9771 (N_9771,N_8051,N_8589);
nor U9772 (N_9772,N_8629,N_8980);
or U9773 (N_9773,N_8862,N_8787);
or U9774 (N_9774,N_8855,N_8341);
xnor U9775 (N_9775,N_8565,N_8142);
nand U9776 (N_9776,N_8120,N_8233);
xor U9777 (N_9777,N_8640,N_8331);
xor U9778 (N_9778,N_8778,N_8710);
nand U9779 (N_9779,N_8064,N_8577);
nand U9780 (N_9780,N_8299,N_8252);
and U9781 (N_9781,N_8073,N_8685);
nand U9782 (N_9782,N_8519,N_8671);
or U9783 (N_9783,N_8024,N_8833);
or U9784 (N_9784,N_8154,N_8899);
nor U9785 (N_9785,N_8645,N_8241);
and U9786 (N_9786,N_8065,N_8731);
and U9787 (N_9787,N_8430,N_8207);
and U9788 (N_9788,N_8270,N_8235);
xor U9789 (N_9789,N_8483,N_8414);
or U9790 (N_9790,N_8657,N_8471);
nand U9791 (N_9791,N_8115,N_8789);
or U9792 (N_9792,N_8731,N_8666);
nand U9793 (N_9793,N_8230,N_8039);
nor U9794 (N_9794,N_8412,N_8288);
xor U9795 (N_9795,N_8645,N_8695);
nor U9796 (N_9796,N_8444,N_8260);
or U9797 (N_9797,N_8512,N_8046);
or U9798 (N_9798,N_8378,N_8047);
nand U9799 (N_9799,N_8587,N_8465);
xor U9800 (N_9800,N_8413,N_8991);
or U9801 (N_9801,N_8049,N_8800);
nor U9802 (N_9802,N_8241,N_8619);
nand U9803 (N_9803,N_8303,N_8543);
or U9804 (N_9804,N_8474,N_8101);
xor U9805 (N_9805,N_8289,N_8627);
and U9806 (N_9806,N_8161,N_8839);
and U9807 (N_9807,N_8061,N_8301);
nand U9808 (N_9808,N_8646,N_8131);
and U9809 (N_9809,N_8243,N_8089);
or U9810 (N_9810,N_8887,N_8619);
and U9811 (N_9811,N_8588,N_8638);
or U9812 (N_9812,N_8117,N_8005);
nand U9813 (N_9813,N_8915,N_8765);
nor U9814 (N_9814,N_8542,N_8752);
nor U9815 (N_9815,N_8196,N_8977);
nor U9816 (N_9816,N_8582,N_8188);
nand U9817 (N_9817,N_8726,N_8819);
or U9818 (N_9818,N_8661,N_8746);
xor U9819 (N_9819,N_8806,N_8587);
and U9820 (N_9820,N_8674,N_8529);
and U9821 (N_9821,N_8567,N_8189);
xor U9822 (N_9822,N_8733,N_8904);
and U9823 (N_9823,N_8236,N_8928);
and U9824 (N_9824,N_8457,N_8658);
and U9825 (N_9825,N_8230,N_8300);
xor U9826 (N_9826,N_8848,N_8660);
or U9827 (N_9827,N_8017,N_8881);
or U9828 (N_9828,N_8733,N_8421);
nor U9829 (N_9829,N_8601,N_8672);
and U9830 (N_9830,N_8638,N_8719);
nand U9831 (N_9831,N_8981,N_8607);
xnor U9832 (N_9832,N_8927,N_8285);
xnor U9833 (N_9833,N_8610,N_8235);
and U9834 (N_9834,N_8417,N_8682);
nor U9835 (N_9835,N_8316,N_8300);
or U9836 (N_9836,N_8795,N_8171);
and U9837 (N_9837,N_8109,N_8098);
nor U9838 (N_9838,N_8867,N_8904);
or U9839 (N_9839,N_8127,N_8868);
nor U9840 (N_9840,N_8354,N_8684);
nor U9841 (N_9841,N_8499,N_8266);
nor U9842 (N_9842,N_8456,N_8597);
nand U9843 (N_9843,N_8385,N_8397);
or U9844 (N_9844,N_8515,N_8688);
nor U9845 (N_9845,N_8924,N_8552);
xnor U9846 (N_9846,N_8466,N_8490);
nor U9847 (N_9847,N_8656,N_8453);
or U9848 (N_9848,N_8707,N_8845);
xnor U9849 (N_9849,N_8871,N_8353);
and U9850 (N_9850,N_8517,N_8524);
nand U9851 (N_9851,N_8445,N_8768);
xor U9852 (N_9852,N_8265,N_8852);
nand U9853 (N_9853,N_8588,N_8440);
and U9854 (N_9854,N_8983,N_8760);
and U9855 (N_9855,N_8014,N_8230);
or U9856 (N_9856,N_8208,N_8673);
and U9857 (N_9857,N_8798,N_8370);
and U9858 (N_9858,N_8171,N_8576);
xnor U9859 (N_9859,N_8628,N_8451);
nor U9860 (N_9860,N_8031,N_8700);
xnor U9861 (N_9861,N_8347,N_8659);
nand U9862 (N_9862,N_8584,N_8316);
xor U9863 (N_9863,N_8368,N_8023);
or U9864 (N_9864,N_8719,N_8281);
xnor U9865 (N_9865,N_8309,N_8409);
and U9866 (N_9866,N_8233,N_8276);
and U9867 (N_9867,N_8944,N_8666);
xnor U9868 (N_9868,N_8406,N_8673);
or U9869 (N_9869,N_8198,N_8636);
nand U9870 (N_9870,N_8282,N_8763);
and U9871 (N_9871,N_8077,N_8639);
or U9872 (N_9872,N_8776,N_8656);
xnor U9873 (N_9873,N_8021,N_8295);
or U9874 (N_9874,N_8980,N_8858);
nand U9875 (N_9875,N_8103,N_8309);
nor U9876 (N_9876,N_8114,N_8789);
and U9877 (N_9877,N_8448,N_8677);
nand U9878 (N_9878,N_8096,N_8966);
or U9879 (N_9879,N_8631,N_8405);
xor U9880 (N_9880,N_8363,N_8295);
or U9881 (N_9881,N_8066,N_8239);
and U9882 (N_9882,N_8924,N_8320);
nand U9883 (N_9883,N_8682,N_8325);
nand U9884 (N_9884,N_8787,N_8784);
nand U9885 (N_9885,N_8141,N_8240);
nand U9886 (N_9886,N_8893,N_8273);
or U9887 (N_9887,N_8693,N_8280);
xnor U9888 (N_9888,N_8882,N_8168);
nand U9889 (N_9889,N_8481,N_8662);
xor U9890 (N_9890,N_8434,N_8166);
or U9891 (N_9891,N_8185,N_8098);
nand U9892 (N_9892,N_8228,N_8628);
nor U9893 (N_9893,N_8004,N_8428);
and U9894 (N_9894,N_8426,N_8268);
nor U9895 (N_9895,N_8846,N_8049);
and U9896 (N_9896,N_8490,N_8508);
or U9897 (N_9897,N_8037,N_8224);
nand U9898 (N_9898,N_8656,N_8150);
or U9899 (N_9899,N_8677,N_8325);
nor U9900 (N_9900,N_8547,N_8958);
nand U9901 (N_9901,N_8540,N_8565);
xor U9902 (N_9902,N_8214,N_8703);
or U9903 (N_9903,N_8668,N_8152);
and U9904 (N_9904,N_8057,N_8216);
or U9905 (N_9905,N_8652,N_8442);
nand U9906 (N_9906,N_8214,N_8291);
or U9907 (N_9907,N_8977,N_8048);
nor U9908 (N_9908,N_8985,N_8203);
nor U9909 (N_9909,N_8236,N_8502);
or U9910 (N_9910,N_8867,N_8535);
nand U9911 (N_9911,N_8794,N_8259);
nand U9912 (N_9912,N_8663,N_8145);
nand U9913 (N_9913,N_8142,N_8838);
nand U9914 (N_9914,N_8883,N_8090);
nor U9915 (N_9915,N_8257,N_8053);
xor U9916 (N_9916,N_8218,N_8014);
and U9917 (N_9917,N_8326,N_8145);
xnor U9918 (N_9918,N_8721,N_8470);
or U9919 (N_9919,N_8659,N_8898);
and U9920 (N_9920,N_8105,N_8425);
nor U9921 (N_9921,N_8901,N_8485);
or U9922 (N_9922,N_8568,N_8848);
or U9923 (N_9923,N_8722,N_8314);
xnor U9924 (N_9924,N_8288,N_8833);
nand U9925 (N_9925,N_8253,N_8439);
xnor U9926 (N_9926,N_8023,N_8743);
or U9927 (N_9927,N_8764,N_8147);
or U9928 (N_9928,N_8444,N_8899);
nor U9929 (N_9929,N_8805,N_8020);
or U9930 (N_9930,N_8148,N_8786);
or U9931 (N_9931,N_8077,N_8863);
or U9932 (N_9932,N_8230,N_8785);
nand U9933 (N_9933,N_8983,N_8063);
xnor U9934 (N_9934,N_8804,N_8321);
or U9935 (N_9935,N_8915,N_8668);
and U9936 (N_9936,N_8619,N_8048);
xnor U9937 (N_9937,N_8555,N_8878);
or U9938 (N_9938,N_8623,N_8110);
or U9939 (N_9939,N_8633,N_8553);
nor U9940 (N_9940,N_8771,N_8686);
nor U9941 (N_9941,N_8150,N_8903);
xor U9942 (N_9942,N_8720,N_8041);
or U9943 (N_9943,N_8554,N_8682);
xnor U9944 (N_9944,N_8978,N_8965);
or U9945 (N_9945,N_8989,N_8403);
or U9946 (N_9946,N_8930,N_8938);
nor U9947 (N_9947,N_8421,N_8590);
and U9948 (N_9948,N_8988,N_8117);
nor U9949 (N_9949,N_8871,N_8751);
nor U9950 (N_9950,N_8638,N_8668);
xor U9951 (N_9951,N_8794,N_8617);
and U9952 (N_9952,N_8675,N_8282);
or U9953 (N_9953,N_8252,N_8539);
or U9954 (N_9954,N_8709,N_8301);
xnor U9955 (N_9955,N_8919,N_8554);
nor U9956 (N_9956,N_8035,N_8927);
xnor U9957 (N_9957,N_8522,N_8813);
and U9958 (N_9958,N_8584,N_8252);
nor U9959 (N_9959,N_8735,N_8817);
and U9960 (N_9960,N_8264,N_8146);
nor U9961 (N_9961,N_8425,N_8511);
nand U9962 (N_9962,N_8737,N_8160);
nand U9963 (N_9963,N_8705,N_8310);
nand U9964 (N_9964,N_8658,N_8901);
nor U9965 (N_9965,N_8731,N_8018);
nand U9966 (N_9966,N_8136,N_8331);
nor U9967 (N_9967,N_8967,N_8722);
and U9968 (N_9968,N_8473,N_8301);
nor U9969 (N_9969,N_8817,N_8621);
nor U9970 (N_9970,N_8923,N_8392);
xnor U9971 (N_9971,N_8284,N_8766);
nand U9972 (N_9972,N_8408,N_8667);
nor U9973 (N_9973,N_8759,N_8077);
nor U9974 (N_9974,N_8518,N_8901);
xnor U9975 (N_9975,N_8534,N_8984);
nand U9976 (N_9976,N_8742,N_8271);
xnor U9977 (N_9977,N_8479,N_8232);
or U9978 (N_9978,N_8853,N_8400);
nand U9979 (N_9979,N_8671,N_8086);
nor U9980 (N_9980,N_8637,N_8056);
nor U9981 (N_9981,N_8573,N_8872);
and U9982 (N_9982,N_8102,N_8748);
and U9983 (N_9983,N_8435,N_8767);
and U9984 (N_9984,N_8139,N_8706);
xnor U9985 (N_9985,N_8361,N_8320);
and U9986 (N_9986,N_8969,N_8556);
nand U9987 (N_9987,N_8870,N_8485);
or U9988 (N_9988,N_8224,N_8541);
xnor U9989 (N_9989,N_8120,N_8847);
and U9990 (N_9990,N_8836,N_8782);
nand U9991 (N_9991,N_8030,N_8520);
nor U9992 (N_9992,N_8155,N_8214);
nand U9993 (N_9993,N_8462,N_8114);
xor U9994 (N_9994,N_8330,N_8165);
nand U9995 (N_9995,N_8739,N_8595);
nor U9996 (N_9996,N_8230,N_8475);
nand U9997 (N_9997,N_8900,N_8018);
nor U9998 (N_9998,N_8367,N_8385);
xor U9999 (N_9999,N_8190,N_8999);
nor U10000 (N_10000,N_9771,N_9468);
xor U10001 (N_10001,N_9688,N_9635);
xor U10002 (N_10002,N_9415,N_9428);
nand U10003 (N_10003,N_9593,N_9937);
nand U10004 (N_10004,N_9904,N_9375);
and U10005 (N_10005,N_9551,N_9436);
and U10006 (N_10006,N_9684,N_9470);
xor U10007 (N_10007,N_9558,N_9977);
xor U10008 (N_10008,N_9751,N_9836);
nand U10009 (N_10009,N_9474,N_9589);
nand U10010 (N_10010,N_9034,N_9199);
or U10011 (N_10011,N_9946,N_9228);
nand U10012 (N_10012,N_9685,N_9732);
and U10013 (N_10013,N_9661,N_9260);
xnor U10014 (N_10014,N_9716,N_9959);
xnor U10015 (N_10015,N_9484,N_9234);
or U10016 (N_10016,N_9888,N_9837);
xor U10017 (N_10017,N_9682,N_9278);
nor U10018 (N_10018,N_9312,N_9958);
nand U10019 (N_10019,N_9962,N_9868);
nand U10020 (N_10020,N_9820,N_9177);
nor U10021 (N_10021,N_9392,N_9862);
and U10022 (N_10022,N_9048,N_9898);
or U10023 (N_10023,N_9262,N_9750);
and U10024 (N_10024,N_9204,N_9102);
or U10025 (N_10025,N_9662,N_9604);
nand U10026 (N_10026,N_9487,N_9001);
or U10027 (N_10027,N_9063,N_9207);
nand U10028 (N_10028,N_9779,N_9710);
xor U10029 (N_10029,N_9988,N_9208);
or U10030 (N_10030,N_9914,N_9894);
and U10031 (N_10031,N_9726,N_9320);
and U10032 (N_10032,N_9215,N_9179);
xnor U10033 (N_10033,N_9957,N_9284);
and U10034 (N_10034,N_9654,N_9292);
nor U10035 (N_10035,N_9683,N_9706);
xor U10036 (N_10036,N_9818,N_9606);
and U10037 (N_10037,N_9964,N_9287);
or U10038 (N_10038,N_9446,N_9056);
xor U10039 (N_10039,N_9037,N_9809);
nor U10040 (N_10040,N_9273,N_9697);
nand U10041 (N_10041,N_9121,N_9972);
xnor U10042 (N_10042,N_9305,N_9354);
and U10043 (N_10043,N_9867,N_9229);
nor U10044 (N_10044,N_9376,N_9736);
nand U10045 (N_10045,N_9197,N_9326);
or U10046 (N_10046,N_9586,N_9950);
nand U10047 (N_10047,N_9335,N_9250);
nor U10048 (N_10048,N_9703,N_9276);
nand U10049 (N_10049,N_9955,N_9473);
nor U10050 (N_10050,N_9355,N_9641);
nor U10051 (N_10051,N_9587,N_9910);
or U10052 (N_10052,N_9164,N_9310);
xor U10053 (N_10053,N_9852,N_9406);
xnor U10054 (N_10054,N_9351,N_9761);
nor U10055 (N_10055,N_9297,N_9347);
nand U10056 (N_10056,N_9731,N_9833);
and U10057 (N_10057,N_9525,N_9924);
nor U10058 (N_10058,N_9848,N_9511);
xnor U10059 (N_10059,N_9502,N_9985);
xor U10060 (N_10060,N_9785,N_9159);
xnor U10061 (N_10061,N_9166,N_9669);
and U10062 (N_10062,N_9879,N_9546);
xor U10063 (N_10063,N_9110,N_9188);
nand U10064 (N_10064,N_9876,N_9532);
nor U10065 (N_10065,N_9040,N_9900);
nor U10066 (N_10066,N_9651,N_9658);
nand U10067 (N_10067,N_9482,N_9097);
nor U10068 (N_10068,N_9638,N_9120);
nand U10069 (N_10069,N_9352,N_9481);
or U10070 (N_10070,N_9861,N_9570);
and U10071 (N_10071,N_9004,N_9382);
nand U10072 (N_10072,N_9644,N_9308);
and U10073 (N_10073,N_9098,N_9686);
and U10074 (N_10074,N_9711,N_9655);
nand U10075 (N_10075,N_9007,N_9117);
xor U10076 (N_10076,N_9242,N_9559);
nor U10077 (N_10077,N_9438,N_9887);
or U10078 (N_10078,N_9170,N_9776);
nor U10079 (N_10079,N_9115,N_9877);
nor U10080 (N_10080,N_9562,N_9423);
or U10081 (N_10081,N_9829,N_9368);
and U10082 (N_10082,N_9344,N_9766);
or U10083 (N_10083,N_9530,N_9025);
nand U10084 (N_10084,N_9053,N_9636);
or U10085 (N_10085,N_9783,N_9496);
or U10086 (N_10086,N_9555,N_9134);
nand U10087 (N_10087,N_9968,N_9533);
or U10088 (N_10088,N_9652,N_9595);
nand U10089 (N_10089,N_9236,N_9384);
and U10090 (N_10090,N_9031,N_9218);
or U10091 (N_10091,N_9069,N_9360);
and U10092 (N_10092,N_9495,N_9026);
xnor U10093 (N_10093,N_9377,N_9926);
or U10094 (N_10094,N_9065,N_9183);
and U10095 (N_10095,N_9461,N_9526);
and U10096 (N_10096,N_9426,N_9801);
nor U10097 (N_10097,N_9138,N_9032);
nor U10098 (N_10098,N_9216,N_9005);
nor U10099 (N_10099,N_9890,N_9393);
xor U10100 (N_10100,N_9489,N_9047);
nand U10101 (N_10101,N_9286,N_9568);
nand U10102 (N_10102,N_9573,N_9788);
xnor U10103 (N_10103,N_9497,N_9980);
nand U10104 (N_10104,N_9918,N_9067);
or U10105 (N_10105,N_9011,N_9509);
and U10106 (N_10106,N_9319,N_9510);
or U10107 (N_10107,N_9214,N_9906);
nand U10108 (N_10108,N_9127,N_9572);
and U10109 (N_10109,N_9927,N_9182);
and U10110 (N_10110,N_9947,N_9363);
nor U10111 (N_10111,N_9830,N_9431);
nor U10112 (N_10112,N_9288,N_9013);
nor U10113 (N_10113,N_9095,N_9444);
xnor U10114 (N_10114,N_9755,N_9154);
xnor U10115 (N_10115,N_9791,N_9739);
nor U10116 (N_10116,N_9306,N_9519);
and U10117 (N_10117,N_9539,N_9342);
or U10118 (N_10118,N_9404,N_9463);
and U10119 (N_10119,N_9349,N_9488);
xnor U10120 (N_10120,N_9581,N_9498);
nand U10121 (N_10121,N_9969,N_9590);
or U10122 (N_10122,N_9709,N_9677);
xnor U10123 (N_10123,N_9209,N_9321);
and U10124 (N_10124,N_9564,N_9049);
nor U10125 (N_10125,N_9241,N_9608);
or U10126 (N_10126,N_9781,N_9029);
or U10127 (N_10127,N_9387,N_9883);
nand U10128 (N_10128,N_9398,N_9812);
nor U10129 (N_10129,N_9113,N_9458);
xnor U10130 (N_10130,N_9621,N_9014);
or U10131 (N_10131,N_9986,N_9615);
xor U10132 (N_10132,N_9094,N_9884);
xnor U10133 (N_10133,N_9309,N_9079);
and U10134 (N_10134,N_9612,N_9540);
and U10135 (N_10135,N_9239,N_9361);
nor U10136 (N_10136,N_9637,N_9022);
xnor U10137 (N_10137,N_9885,N_9493);
xnor U10138 (N_10138,N_9993,N_9777);
xor U10139 (N_10139,N_9831,N_9858);
nand U10140 (N_10140,N_9994,N_9729);
nand U10141 (N_10141,N_9003,N_9583);
nor U10142 (N_10142,N_9220,N_9018);
xnor U10143 (N_10143,N_9191,N_9718);
xor U10144 (N_10144,N_9720,N_9506);
and U10145 (N_10145,N_9388,N_9650);
nor U10146 (N_10146,N_9698,N_9329);
nor U10147 (N_10147,N_9042,N_9293);
nand U10148 (N_10148,N_9936,N_9033);
and U10149 (N_10149,N_9841,N_9690);
and U10150 (N_10150,N_9941,N_9563);
and U10151 (N_10151,N_9476,N_9456);
and U10152 (N_10152,N_9804,N_9060);
nor U10153 (N_10153,N_9092,N_9405);
nand U10154 (N_10154,N_9261,N_9624);
nor U10155 (N_10155,N_9920,N_9106);
nor U10156 (N_10156,N_9847,N_9002);
or U10157 (N_10157,N_9210,N_9998);
or U10158 (N_10158,N_9246,N_9571);
and U10159 (N_10159,N_9547,N_9141);
and U10160 (N_10160,N_9737,N_9850);
xnor U10161 (N_10161,N_9317,N_9853);
nor U10162 (N_10162,N_9648,N_9917);
nand U10163 (N_10163,N_9350,N_9940);
xor U10164 (N_10164,N_9325,N_9348);
and U10165 (N_10165,N_9765,N_9882);
xnor U10166 (N_10166,N_9613,N_9130);
xnor U10167 (N_10167,N_9915,N_9815);
nand U10168 (N_10168,N_9125,N_9870);
xor U10169 (N_10169,N_9365,N_9548);
or U10170 (N_10170,N_9758,N_9992);
nand U10171 (N_10171,N_9921,N_9948);
or U10172 (N_10172,N_9327,N_9507);
nor U10173 (N_10173,N_9514,N_9660);
and U10174 (N_10174,N_9235,N_9000);
nand U10175 (N_10175,N_9640,N_9932);
nor U10176 (N_10176,N_9741,N_9006);
nand U10177 (N_10177,N_9696,N_9826);
nor U10178 (N_10178,N_9078,N_9735);
nand U10179 (N_10179,N_9421,N_9175);
nand U10180 (N_10180,N_9895,N_9753);
or U10181 (N_10181,N_9050,N_9453);
xor U10182 (N_10182,N_9338,N_9978);
xnor U10183 (N_10183,N_9919,N_9222);
nand U10184 (N_10184,N_9395,N_9550);
xor U10185 (N_10185,N_9083,N_9171);
xor U10186 (N_10186,N_9096,N_9332);
nand U10187 (N_10187,N_9517,N_9605);
xnor U10188 (N_10188,N_9925,N_9633);
nor U10189 (N_10189,N_9093,N_9074);
or U10190 (N_10190,N_9903,N_9762);
or U10191 (N_10191,N_9422,N_9574);
xor U10192 (N_10192,N_9524,N_9201);
nor U10193 (N_10193,N_9816,N_9668);
nor U10194 (N_10194,N_9128,N_9723);
or U10195 (N_10195,N_9435,N_9109);
nand U10196 (N_10196,N_9975,N_9080);
or U10197 (N_10197,N_9410,N_9963);
xnor U10198 (N_10198,N_9237,N_9800);
and U10199 (N_10199,N_9880,N_9614);
xor U10200 (N_10200,N_9872,N_9869);
nand U10201 (N_10201,N_9359,N_9675);
nand U10202 (N_10202,N_9591,N_9749);
nor U10203 (N_10203,N_9203,N_9967);
nand U10204 (N_10204,N_9643,N_9299);
xnor U10205 (N_10205,N_9202,N_9694);
and U10206 (N_10206,N_9036,N_9270);
or U10207 (N_10207,N_9930,N_9784);
nand U10208 (N_10208,N_9943,N_9667);
and U10209 (N_10209,N_9631,N_9206);
nand U10210 (N_10210,N_9137,N_9369);
xor U10211 (N_10211,N_9730,N_9534);
or U10212 (N_10212,N_9748,N_9970);
nor U10213 (N_10213,N_9854,N_9584);
nor U10214 (N_10214,N_9195,N_9399);
nand U10215 (N_10215,N_9371,N_9200);
and U10216 (N_10216,N_9440,N_9027);
nand U10217 (N_10217,N_9066,N_9795);
or U10218 (N_10218,N_9126,N_9073);
and U10219 (N_10219,N_9501,N_9623);
or U10220 (N_10220,N_9044,N_9782);
nand U10221 (N_10221,N_9923,N_9545);
nor U10222 (N_10222,N_9577,N_9827);
xor U10223 (N_10223,N_9905,N_9775);
nand U10224 (N_10224,N_9646,N_9708);
nor U10225 (N_10225,N_9588,N_9521);
nand U10226 (N_10226,N_9580,N_9717);
nand U10227 (N_10227,N_9185,N_9911);
xnor U10228 (N_10228,N_9275,N_9017);
nor U10229 (N_10229,N_9151,N_9433);
xnor U10230 (N_10230,N_9780,N_9045);
nor U10231 (N_10231,N_9023,N_9855);
nor U10232 (N_10232,N_9322,N_9454);
nand U10233 (N_10233,N_9089,N_9626);
xor U10234 (N_10234,N_9238,N_9483);
and U10235 (N_10235,N_9806,N_9609);
xor U10236 (N_10236,N_9617,N_9944);
nor U10237 (N_10237,N_9192,N_9908);
nand U10238 (N_10238,N_9180,N_9010);
and U10239 (N_10239,N_9754,N_9328);
xor U10240 (N_10240,N_9418,N_9679);
nand U10241 (N_10241,N_9653,N_9929);
and U10242 (N_10242,N_9362,N_9490);
xor U10243 (N_10243,N_9528,N_9657);
and U10244 (N_10244,N_9071,N_9249);
xnor U10245 (N_10245,N_9851,N_9860);
nor U10246 (N_10246,N_9835,N_9727);
and U10247 (N_10247,N_9448,N_9971);
xor U10248 (N_10248,N_9162,N_9107);
xnor U10249 (N_10249,N_9274,N_9099);
nor U10250 (N_10250,N_9401,N_9465);
and U10251 (N_10251,N_9757,N_9557);
nor U10252 (N_10252,N_9380,N_9337);
nand U10253 (N_10253,N_9466,N_9692);
nand U10254 (N_10254,N_9952,N_9233);
and U10255 (N_10255,N_9687,N_9263);
nand U10256 (N_10256,N_9085,N_9913);
and U10257 (N_10257,N_9336,N_9316);
nand U10258 (N_10258,N_9021,N_9302);
or U10259 (N_10259,N_9663,N_9184);
and U10260 (N_10260,N_9909,N_9928);
xor U10261 (N_10261,N_9700,N_9279);
nand U10262 (N_10262,N_9907,N_9062);
nand U10263 (N_10263,N_9015,N_9665);
or U10264 (N_10264,N_9719,N_9020);
xor U10265 (N_10265,N_9585,N_9370);
and U10266 (N_10266,N_9445,N_9224);
and U10267 (N_10267,N_9459,N_9298);
nand U10268 (N_10268,N_9267,N_9429);
nor U10269 (N_10269,N_9172,N_9659);
xor U10270 (N_10270,N_9627,N_9983);
nor U10271 (N_10271,N_9645,N_9118);
nor U10272 (N_10272,N_9596,N_9979);
nor U10273 (N_10273,N_9756,N_9542);
and U10274 (N_10274,N_9272,N_9999);
xor U10275 (N_10275,N_9255,N_9133);
or U10276 (N_10276,N_9916,N_9119);
nor U10277 (N_10277,N_9701,N_9714);
xnor U10278 (N_10278,N_9632,N_9642);
or U10279 (N_10279,N_9902,N_9949);
and U10280 (N_10280,N_9283,N_9226);
nor U10281 (N_10281,N_9285,N_9464);
nor U10282 (N_10282,N_9715,N_9733);
and U10283 (N_10283,N_9523,N_9467);
and U10284 (N_10284,N_9770,N_9565);
nand U10285 (N_10285,N_9313,N_9265);
nor U10286 (N_10286,N_9213,N_9124);
or U10287 (N_10287,N_9190,N_9300);
and U10288 (N_10288,N_9742,N_9939);
and U10289 (N_10289,N_9394,N_9691);
xnor U10290 (N_10290,N_9019,N_9449);
or U10291 (N_10291,N_9039,N_9560);
and U10292 (N_10292,N_9374,N_9075);
or U10293 (N_10293,N_9081,N_9807);
and U10294 (N_10294,N_9747,N_9146);
or U10295 (N_10295,N_9030,N_9024);
and U10296 (N_10296,N_9432,N_9251);
nor U10297 (N_10297,N_9630,N_9656);
and U10298 (N_10298,N_9439,N_9379);
nand U10299 (N_10299,N_9383,N_9984);
and U10300 (N_10300,N_9499,N_9543);
nand U10301 (N_10301,N_9174,N_9427);
or U10302 (N_10302,N_9520,N_9148);
and U10303 (N_10303,N_9114,N_9341);
xnor U10304 (N_10304,N_9028,N_9061);
and U10305 (N_10305,N_9161,N_9554);
nand U10306 (N_10306,N_9789,N_9689);
xor U10307 (N_10307,N_9649,N_9212);
xor U10308 (N_10308,N_9430,N_9043);
and U10309 (N_10309,N_9610,N_9152);
nor U10310 (N_10310,N_9976,N_9728);
nand U10311 (N_10311,N_9378,N_9457);
xor U10312 (N_10312,N_9960,N_9803);
xor U10313 (N_10313,N_9280,N_9712);
or U10314 (N_10314,N_9996,N_9536);
nor U10315 (N_10315,N_9527,N_9419);
or U10316 (N_10316,N_9258,N_9620);
or U10317 (N_10317,N_9230,N_9254);
and U10318 (N_10318,N_9893,N_9296);
xnor U10319 (N_10319,N_9752,N_9538);
nor U10320 (N_10320,N_9938,N_9289);
xnor U10321 (N_10321,N_9139,N_9147);
or U10322 (N_10322,N_9515,N_9556);
or U10323 (N_10323,N_9386,N_9391);
xnor U10324 (N_10324,N_9157,N_9385);
xnor U10325 (N_10325,N_9790,N_9169);
nor U10326 (N_10326,N_9366,N_9345);
nor U10327 (N_10327,N_9541,N_9492);
nand U10328 (N_10328,N_9009,N_9318);
or U10329 (N_10329,N_9769,N_9232);
xor U10330 (N_10330,N_9598,N_9512);
and U10331 (N_10331,N_9480,N_9567);
nor U10332 (N_10332,N_9264,N_9412);
xnor U10333 (N_10333,N_9603,N_9140);
xor U10334 (N_10334,N_9695,N_9135);
nand U10335 (N_10335,N_9674,N_9934);
xor U10336 (N_10336,N_9403,N_9734);
nor U10337 (N_10337,N_9068,N_9805);
nor U10338 (N_10338,N_9167,N_9504);
and U10339 (N_10339,N_9822,N_9054);
and U10340 (N_10340,N_9997,N_9186);
xnor U10341 (N_10341,N_9123,N_9301);
nand U10342 (N_10342,N_9721,N_9076);
nand U10343 (N_10343,N_9221,N_9447);
and U10344 (N_10344,N_9163,N_9874);
or U10345 (N_10345,N_9173,N_9295);
or U10346 (N_10346,N_9500,N_9840);
nor U10347 (N_10347,N_9477,N_9865);
or U10348 (N_10348,N_9103,N_9266);
or U10349 (N_10349,N_9244,N_9535);
or U10350 (N_10350,N_9472,N_9856);
xor U10351 (N_10351,N_9602,N_9839);
xor U10352 (N_10352,N_9973,N_9823);
and U10353 (N_10353,N_9672,N_9304);
and U10354 (N_10354,N_9743,N_9843);
or U10355 (N_10355,N_9475,N_9100);
and U10356 (N_10356,N_9012,N_9390);
and U10357 (N_10357,N_9844,N_9082);
nand U10358 (N_10358,N_9131,N_9248);
xor U10359 (N_10359,N_9271,N_9931);
and U10360 (N_10360,N_9413,N_9252);
xnor U10361 (N_10361,N_9494,N_9101);
nor U10362 (N_10362,N_9838,N_9607);
or U10363 (N_10363,N_9340,N_9866);
xnor U10364 (N_10364,N_9323,N_9176);
and U10365 (N_10365,N_9425,N_9767);
nor U10366 (N_10366,N_9051,N_9486);
nor U10367 (N_10367,N_9673,N_9343);
nor U10368 (N_10368,N_9995,N_9257);
and U10369 (N_10369,N_9451,N_9824);
nor U10370 (N_10370,N_9090,N_9745);
or U10371 (N_10371,N_9738,N_9629);
xor U10372 (N_10372,N_9108,N_9143);
nand U10373 (N_10373,N_9664,N_9281);
xnor U10374 (N_10374,N_9294,N_9205);
or U10375 (N_10375,N_9849,N_9578);
or U10376 (N_10376,N_9953,N_9112);
or U10377 (N_10377,N_9819,N_9569);
and U10378 (N_10378,N_9954,N_9277);
xnor U10379 (N_10379,N_9896,N_9981);
nor U10380 (N_10380,N_9334,N_9680);
and U10381 (N_10381,N_9508,N_9240);
or U10382 (N_10382,N_9307,N_9544);
nor U10383 (N_10383,N_9989,N_9786);
or U10384 (N_10384,N_9724,N_9740);
nand U10385 (N_10385,N_9942,N_9291);
xnor U10386 (N_10386,N_9424,N_9619);
xor U10387 (N_10387,N_9084,N_9821);
nor U10388 (N_10388,N_9671,N_9798);
nand U10389 (N_10389,N_9759,N_9808);
or U10390 (N_10390,N_9441,N_9611);
xor U10391 (N_10391,N_9773,N_9945);
nor U10392 (N_10392,N_9817,N_9647);
and U10393 (N_10393,N_9705,N_9764);
and U10394 (N_10394,N_9871,N_9016);
xor U10395 (N_10395,N_9485,N_9358);
xnor U10396 (N_10396,N_9503,N_9217);
nand U10397 (N_10397,N_9537,N_9058);
or U10398 (N_10398,N_9522,N_9707);
xnor U10399 (N_10399,N_9966,N_9746);
xor U10400 (N_10400,N_9402,N_9518);
nand U10401 (N_10401,N_9892,N_9303);
xor U10402 (N_10402,N_9846,N_9878);
nand U10403 (N_10403,N_9597,N_9478);
xor U10404 (N_10404,N_9064,N_9414);
nand U10405 (N_10405,N_9057,N_9132);
and U10406 (N_10406,N_9797,N_9987);
nor U10407 (N_10407,N_9832,N_9153);
and U10408 (N_10408,N_9396,N_9437);
xor U10409 (N_10409,N_9149,N_9859);
and U10410 (N_10410,N_9666,N_9549);
xnor U10411 (N_10411,N_9223,N_9256);
and U10412 (N_10412,N_9253,N_9160);
xnor U10413 (N_10413,N_9863,N_9702);
and U10414 (N_10414,N_9196,N_9901);
or U10415 (N_10415,N_9634,N_9330);
and U10416 (N_10416,N_9982,N_9794);
or U10417 (N_10417,N_9531,N_9052);
and U10418 (N_10418,N_9247,N_9193);
nor U10419 (N_10419,N_9834,N_9129);
nand U10420 (N_10420,N_9802,N_9144);
xor U10421 (N_10421,N_9625,N_9787);
and U10422 (N_10422,N_9181,N_9864);
nor U10423 (N_10423,N_9462,N_9156);
nand U10424 (N_10424,N_9411,N_9744);
xor U10425 (N_10425,N_9842,N_9678);
and U10426 (N_10426,N_9077,N_9813);
nand U10427 (N_10427,N_9793,N_9145);
nand U10428 (N_10428,N_9091,N_9409);
nand U10429 (N_10429,N_9814,N_9713);
or U10430 (N_10430,N_9951,N_9346);
xnor U10431 (N_10431,N_9245,N_9087);
and U10432 (N_10432,N_9616,N_9990);
nand U10433 (N_10433,N_9356,N_9269);
and U10434 (N_10434,N_9136,N_9035);
nand U10435 (N_10435,N_9873,N_9227);
xnor U10436 (N_10436,N_9104,N_9886);
and U10437 (N_10437,N_9857,N_9072);
nor U10438 (N_10438,N_9553,N_9367);
nor U10439 (N_10439,N_9243,N_9935);
nor U10440 (N_10440,N_9059,N_9116);
nand U10441 (N_10441,N_9845,N_9529);
and U10442 (N_10442,N_9704,N_9225);
and U10443 (N_10443,N_9774,N_9443);
or U10444 (N_10444,N_9991,N_9324);
nand U10445 (N_10445,N_9142,N_9282);
nor U10446 (N_10446,N_9956,N_9416);
nand U10447 (N_10447,N_9639,N_9922);
xnor U10448 (N_10448,N_9592,N_9357);
and U10449 (N_10449,N_9420,N_9155);
and U10450 (N_10450,N_9974,N_9491);
nand U10451 (N_10451,N_9471,N_9772);
or U10452 (N_10452,N_9768,N_9189);
or U10453 (N_10453,N_9055,N_9889);
xor U10454 (N_10454,N_9372,N_9618);
or U10455 (N_10455,N_9046,N_9796);
or U10456 (N_10456,N_9373,N_9198);
nand U10457 (N_10457,N_9314,N_9600);
nor U10458 (N_10458,N_9601,N_9778);
xnor U10459 (N_10459,N_9070,N_9582);
xor U10460 (N_10460,N_9259,N_9961);
and U10461 (N_10461,N_9579,N_9008);
xor U10462 (N_10462,N_9168,N_9455);
and U10463 (N_10463,N_9933,N_9041);
or U10464 (N_10464,N_9158,N_9799);
or U10465 (N_10465,N_9333,N_9194);
and U10466 (N_10466,N_9760,N_9460);
and U10467 (N_10467,N_9912,N_9311);
nor U10468 (N_10468,N_9407,N_9965);
and U10469 (N_10469,N_9792,N_9479);
nor U10470 (N_10470,N_9725,N_9561);
and U10471 (N_10471,N_9400,N_9122);
nor U10472 (N_10472,N_9450,N_9881);
nor U10473 (N_10473,N_9628,N_9088);
xnor U10474 (N_10474,N_9331,N_9187);
or U10475 (N_10475,N_9875,N_9576);
and U10476 (N_10476,N_9676,N_9290);
and U10477 (N_10477,N_9594,N_9353);
and U10478 (N_10478,N_9452,N_9505);
or U10479 (N_10479,N_9165,N_9825);
xor U10480 (N_10480,N_9811,N_9566);
or U10481 (N_10481,N_9899,N_9086);
or U10482 (N_10482,N_9513,N_9891);
xor U10483 (N_10483,N_9417,N_9810);
nor U10484 (N_10484,N_9516,N_9693);
and U10485 (N_10485,N_9178,N_9268);
or U10486 (N_10486,N_9231,N_9389);
nand U10487 (N_10487,N_9599,N_9681);
nor U10488 (N_10488,N_9670,N_9828);
nor U10489 (N_10489,N_9897,N_9397);
or U10490 (N_10490,N_9763,N_9364);
nor U10491 (N_10491,N_9211,N_9105);
xor U10492 (N_10492,N_9552,N_9219);
nand U10493 (N_10493,N_9150,N_9111);
xor U10494 (N_10494,N_9315,N_9722);
and U10495 (N_10495,N_9381,N_9469);
xor U10496 (N_10496,N_9408,N_9038);
nand U10497 (N_10497,N_9442,N_9575);
and U10498 (N_10498,N_9434,N_9339);
nor U10499 (N_10499,N_9622,N_9699);
nand U10500 (N_10500,N_9828,N_9620);
nand U10501 (N_10501,N_9123,N_9080);
xnor U10502 (N_10502,N_9782,N_9646);
and U10503 (N_10503,N_9684,N_9258);
and U10504 (N_10504,N_9331,N_9929);
nor U10505 (N_10505,N_9392,N_9082);
nor U10506 (N_10506,N_9400,N_9376);
or U10507 (N_10507,N_9253,N_9868);
nand U10508 (N_10508,N_9714,N_9824);
nor U10509 (N_10509,N_9142,N_9457);
xnor U10510 (N_10510,N_9516,N_9387);
xor U10511 (N_10511,N_9153,N_9909);
nand U10512 (N_10512,N_9206,N_9637);
or U10513 (N_10513,N_9939,N_9032);
or U10514 (N_10514,N_9482,N_9750);
nand U10515 (N_10515,N_9578,N_9865);
and U10516 (N_10516,N_9748,N_9062);
or U10517 (N_10517,N_9488,N_9163);
nand U10518 (N_10518,N_9304,N_9039);
or U10519 (N_10519,N_9092,N_9530);
and U10520 (N_10520,N_9011,N_9165);
xnor U10521 (N_10521,N_9967,N_9692);
and U10522 (N_10522,N_9397,N_9768);
xnor U10523 (N_10523,N_9255,N_9413);
xor U10524 (N_10524,N_9400,N_9430);
or U10525 (N_10525,N_9307,N_9572);
xnor U10526 (N_10526,N_9457,N_9323);
or U10527 (N_10527,N_9215,N_9305);
nor U10528 (N_10528,N_9999,N_9238);
nor U10529 (N_10529,N_9590,N_9055);
nor U10530 (N_10530,N_9240,N_9995);
or U10531 (N_10531,N_9450,N_9135);
xnor U10532 (N_10532,N_9418,N_9609);
or U10533 (N_10533,N_9428,N_9404);
nor U10534 (N_10534,N_9913,N_9719);
nor U10535 (N_10535,N_9512,N_9750);
and U10536 (N_10536,N_9662,N_9590);
xor U10537 (N_10537,N_9750,N_9552);
nand U10538 (N_10538,N_9343,N_9410);
nand U10539 (N_10539,N_9261,N_9063);
xor U10540 (N_10540,N_9760,N_9932);
and U10541 (N_10541,N_9369,N_9269);
and U10542 (N_10542,N_9934,N_9636);
nand U10543 (N_10543,N_9273,N_9275);
and U10544 (N_10544,N_9596,N_9861);
nor U10545 (N_10545,N_9396,N_9525);
or U10546 (N_10546,N_9634,N_9389);
nand U10547 (N_10547,N_9424,N_9975);
nor U10548 (N_10548,N_9084,N_9962);
nand U10549 (N_10549,N_9528,N_9610);
and U10550 (N_10550,N_9346,N_9669);
or U10551 (N_10551,N_9555,N_9028);
and U10552 (N_10552,N_9374,N_9237);
nand U10553 (N_10553,N_9105,N_9528);
xor U10554 (N_10554,N_9424,N_9066);
and U10555 (N_10555,N_9022,N_9557);
xor U10556 (N_10556,N_9327,N_9841);
xor U10557 (N_10557,N_9011,N_9500);
nand U10558 (N_10558,N_9052,N_9165);
xor U10559 (N_10559,N_9785,N_9801);
nand U10560 (N_10560,N_9539,N_9493);
or U10561 (N_10561,N_9606,N_9577);
or U10562 (N_10562,N_9762,N_9788);
and U10563 (N_10563,N_9865,N_9112);
nor U10564 (N_10564,N_9941,N_9666);
nor U10565 (N_10565,N_9226,N_9322);
xnor U10566 (N_10566,N_9797,N_9320);
or U10567 (N_10567,N_9490,N_9599);
xor U10568 (N_10568,N_9549,N_9915);
and U10569 (N_10569,N_9908,N_9088);
nand U10570 (N_10570,N_9282,N_9268);
nand U10571 (N_10571,N_9159,N_9216);
xnor U10572 (N_10572,N_9161,N_9331);
xnor U10573 (N_10573,N_9928,N_9224);
and U10574 (N_10574,N_9719,N_9124);
and U10575 (N_10575,N_9244,N_9731);
or U10576 (N_10576,N_9394,N_9695);
xnor U10577 (N_10577,N_9871,N_9664);
xnor U10578 (N_10578,N_9496,N_9736);
xor U10579 (N_10579,N_9824,N_9616);
and U10580 (N_10580,N_9296,N_9725);
nor U10581 (N_10581,N_9798,N_9329);
and U10582 (N_10582,N_9801,N_9664);
or U10583 (N_10583,N_9266,N_9496);
nor U10584 (N_10584,N_9380,N_9017);
and U10585 (N_10585,N_9139,N_9562);
nor U10586 (N_10586,N_9884,N_9095);
nor U10587 (N_10587,N_9370,N_9787);
nand U10588 (N_10588,N_9974,N_9261);
xor U10589 (N_10589,N_9822,N_9853);
or U10590 (N_10590,N_9989,N_9534);
nand U10591 (N_10591,N_9158,N_9914);
or U10592 (N_10592,N_9025,N_9885);
or U10593 (N_10593,N_9787,N_9096);
and U10594 (N_10594,N_9894,N_9000);
nor U10595 (N_10595,N_9742,N_9795);
nor U10596 (N_10596,N_9257,N_9395);
xnor U10597 (N_10597,N_9809,N_9803);
and U10598 (N_10598,N_9004,N_9707);
and U10599 (N_10599,N_9005,N_9489);
nand U10600 (N_10600,N_9755,N_9396);
nand U10601 (N_10601,N_9497,N_9496);
nor U10602 (N_10602,N_9709,N_9894);
and U10603 (N_10603,N_9114,N_9454);
and U10604 (N_10604,N_9422,N_9712);
xor U10605 (N_10605,N_9515,N_9557);
or U10606 (N_10606,N_9198,N_9524);
xor U10607 (N_10607,N_9422,N_9276);
or U10608 (N_10608,N_9468,N_9583);
nand U10609 (N_10609,N_9076,N_9288);
xor U10610 (N_10610,N_9009,N_9350);
nand U10611 (N_10611,N_9256,N_9333);
xnor U10612 (N_10612,N_9405,N_9381);
nand U10613 (N_10613,N_9634,N_9540);
xor U10614 (N_10614,N_9843,N_9858);
nor U10615 (N_10615,N_9629,N_9632);
and U10616 (N_10616,N_9737,N_9300);
nor U10617 (N_10617,N_9451,N_9650);
xnor U10618 (N_10618,N_9458,N_9626);
or U10619 (N_10619,N_9301,N_9270);
nor U10620 (N_10620,N_9901,N_9940);
nand U10621 (N_10621,N_9072,N_9964);
xor U10622 (N_10622,N_9779,N_9926);
xor U10623 (N_10623,N_9605,N_9315);
nand U10624 (N_10624,N_9352,N_9615);
xor U10625 (N_10625,N_9856,N_9065);
and U10626 (N_10626,N_9775,N_9572);
xnor U10627 (N_10627,N_9003,N_9223);
nor U10628 (N_10628,N_9929,N_9369);
nor U10629 (N_10629,N_9448,N_9240);
xnor U10630 (N_10630,N_9935,N_9902);
and U10631 (N_10631,N_9661,N_9206);
xnor U10632 (N_10632,N_9165,N_9307);
nor U10633 (N_10633,N_9529,N_9829);
and U10634 (N_10634,N_9079,N_9857);
xnor U10635 (N_10635,N_9657,N_9390);
nor U10636 (N_10636,N_9330,N_9671);
nor U10637 (N_10637,N_9574,N_9286);
nand U10638 (N_10638,N_9120,N_9394);
nor U10639 (N_10639,N_9077,N_9508);
or U10640 (N_10640,N_9449,N_9260);
or U10641 (N_10641,N_9323,N_9377);
xor U10642 (N_10642,N_9346,N_9439);
and U10643 (N_10643,N_9995,N_9455);
nand U10644 (N_10644,N_9269,N_9532);
and U10645 (N_10645,N_9644,N_9869);
nand U10646 (N_10646,N_9920,N_9313);
or U10647 (N_10647,N_9337,N_9238);
and U10648 (N_10648,N_9300,N_9802);
and U10649 (N_10649,N_9119,N_9395);
and U10650 (N_10650,N_9817,N_9041);
or U10651 (N_10651,N_9248,N_9466);
nor U10652 (N_10652,N_9274,N_9813);
and U10653 (N_10653,N_9392,N_9419);
and U10654 (N_10654,N_9397,N_9882);
nor U10655 (N_10655,N_9962,N_9250);
xor U10656 (N_10656,N_9629,N_9854);
nor U10657 (N_10657,N_9059,N_9970);
and U10658 (N_10658,N_9984,N_9244);
xnor U10659 (N_10659,N_9181,N_9894);
xor U10660 (N_10660,N_9099,N_9182);
nand U10661 (N_10661,N_9022,N_9754);
nor U10662 (N_10662,N_9240,N_9237);
nor U10663 (N_10663,N_9841,N_9823);
nand U10664 (N_10664,N_9953,N_9586);
and U10665 (N_10665,N_9893,N_9676);
nand U10666 (N_10666,N_9199,N_9985);
or U10667 (N_10667,N_9364,N_9347);
nor U10668 (N_10668,N_9019,N_9536);
nand U10669 (N_10669,N_9782,N_9418);
nor U10670 (N_10670,N_9124,N_9649);
nor U10671 (N_10671,N_9517,N_9726);
or U10672 (N_10672,N_9278,N_9895);
xor U10673 (N_10673,N_9289,N_9103);
nand U10674 (N_10674,N_9615,N_9029);
nor U10675 (N_10675,N_9403,N_9301);
nor U10676 (N_10676,N_9851,N_9388);
nand U10677 (N_10677,N_9387,N_9223);
and U10678 (N_10678,N_9521,N_9256);
nand U10679 (N_10679,N_9311,N_9341);
and U10680 (N_10680,N_9592,N_9582);
nor U10681 (N_10681,N_9463,N_9015);
nor U10682 (N_10682,N_9149,N_9915);
xnor U10683 (N_10683,N_9256,N_9230);
nor U10684 (N_10684,N_9001,N_9884);
nand U10685 (N_10685,N_9568,N_9980);
and U10686 (N_10686,N_9078,N_9229);
and U10687 (N_10687,N_9096,N_9870);
nand U10688 (N_10688,N_9774,N_9580);
and U10689 (N_10689,N_9621,N_9866);
nor U10690 (N_10690,N_9482,N_9099);
nor U10691 (N_10691,N_9673,N_9517);
nor U10692 (N_10692,N_9413,N_9908);
or U10693 (N_10693,N_9757,N_9896);
xnor U10694 (N_10694,N_9187,N_9994);
nor U10695 (N_10695,N_9033,N_9285);
nor U10696 (N_10696,N_9010,N_9737);
nor U10697 (N_10697,N_9780,N_9474);
nor U10698 (N_10698,N_9366,N_9807);
nand U10699 (N_10699,N_9328,N_9024);
nor U10700 (N_10700,N_9775,N_9314);
or U10701 (N_10701,N_9945,N_9389);
or U10702 (N_10702,N_9127,N_9370);
nor U10703 (N_10703,N_9407,N_9563);
and U10704 (N_10704,N_9469,N_9730);
or U10705 (N_10705,N_9341,N_9006);
and U10706 (N_10706,N_9195,N_9529);
or U10707 (N_10707,N_9052,N_9897);
nor U10708 (N_10708,N_9650,N_9630);
or U10709 (N_10709,N_9455,N_9447);
nor U10710 (N_10710,N_9852,N_9280);
nor U10711 (N_10711,N_9866,N_9733);
nand U10712 (N_10712,N_9442,N_9457);
nor U10713 (N_10713,N_9682,N_9275);
and U10714 (N_10714,N_9882,N_9304);
nor U10715 (N_10715,N_9364,N_9781);
nor U10716 (N_10716,N_9069,N_9479);
nor U10717 (N_10717,N_9910,N_9353);
nor U10718 (N_10718,N_9618,N_9308);
nand U10719 (N_10719,N_9203,N_9417);
nand U10720 (N_10720,N_9601,N_9551);
xor U10721 (N_10721,N_9241,N_9342);
and U10722 (N_10722,N_9227,N_9349);
and U10723 (N_10723,N_9212,N_9485);
or U10724 (N_10724,N_9303,N_9451);
and U10725 (N_10725,N_9124,N_9358);
nor U10726 (N_10726,N_9215,N_9258);
nor U10727 (N_10727,N_9203,N_9950);
or U10728 (N_10728,N_9876,N_9133);
or U10729 (N_10729,N_9883,N_9832);
or U10730 (N_10730,N_9481,N_9091);
or U10731 (N_10731,N_9291,N_9259);
xor U10732 (N_10732,N_9372,N_9759);
or U10733 (N_10733,N_9999,N_9091);
xnor U10734 (N_10734,N_9136,N_9585);
and U10735 (N_10735,N_9131,N_9890);
or U10736 (N_10736,N_9463,N_9246);
nor U10737 (N_10737,N_9919,N_9193);
xnor U10738 (N_10738,N_9329,N_9321);
or U10739 (N_10739,N_9724,N_9109);
and U10740 (N_10740,N_9308,N_9245);
nor U10741 (N_10741,N_9164,N_9884);
nor U10742 (N_10742,N_9517,N_9520);
or U10743 (N_10743,N_9298,N_9301);
or U10744 (N_10744,N_9120,N_9448);
and U10745 (N_10745,N_9579,N_9375);
nand U10746 (N_10746,N_9622,N_9452);
nand U10747 (N_10747,N_9548,N_9020);
nor U10748 (N_10748,N_9939,N_9407);
and U10749 (N_10749,N_9639,N_9551);
xnor U10750 (N_10750,N_9168,N_9339);
xor U10751 (N_10751,N_9417,N_9303);
xor U10752 (N_10752,N_9177,N_9973);
and U10753 (N_10753,N_9780,N_9772);
nor U10754 (N_10754,N_9221,N_9784);
nor U10755 (N_10755,N_9629,N_9759);
nand U10756 (N_10756,N_9565,N_9260);
or U10757 (N_10757,N_9953,N_9703);
or U10758 (N_10758,N_9328,N_9305);
and U10759 (N_10759,N_9657,N_9663);
or U10760 (N_10760,N_9615,N_9654);
nor U10761 (N_10761,N_9629,N_9760);
nor U10762 (N_10762,N_9110,N_9598);
or U10763 (N_10763,N_9228,N_9775);
or U10764 (N_10764,N_9881,N_9393);
and U10765 (N_10765,N_9514,N_9231);
and U10766 (N_10766,N_9400,N_9782);
nand U10767 (N_10767,N_9985,N_9729);
nor U10768 (N_10768,N_9994,N_9349);
nand U10769 (N_10769,N_9391,N_9370);
and U10770 (N_10770,N_9339,N_9609);
or U10771 (N_10771,N_9921,N_9870);
nand U10772 (N_10772,N_9410,N_9385);
or U10773 (N_10773,N_9125,N_9749);
nor U10774 (N_10774,N_9394,N_9959);
nand U10775 (N_10775,N_9355,N_9282);
or U10776 (N_10776,N_9566,N_9830);
nor U10777 (N_10777,N_9684,N_9183);
nand U10778 (N_10778,N_9744,N_9537);
xor U10779 (N_10779,N_9966,N_9082);
nand U10780 (N_10780,N_9042,N_9858);
xor U10781 (N_10781,N_9767,N_9995);
and U10782 (N_10782,N_9905,N_9850);
nor U10783 (N_10783,N_9387,N_9272);
and U10784 (N_10784,N_9060,N_9563);
nor U10785 (N_10785,N_9879,N_9923);
and U10786 (N_10786,N_9921,N_9997);
nand U10787 (N_10787,N_9386,N_9653);
nand U10788 (N_10788,N_9276,N_9000);
nand U10789 (N_10789,N_9030,N_9438);
and U10790 (N_10790,N_9057,N_9318);
and U10791 (N_10791,N_9156,N_9065);
nor U10792 (N_10792,N_9358,N_9457);
xor U10793 (N_10793,N_9673,N_9912);
xnor U10794 (N_10794,N_9472,N_9637);
xor U10795 (N_10795,N_9682,N_9087);
or U10796 (N_10796,N_9418,N_9167);
nand U10797 (N_10797,N_9020,N_9094);
or U10798 (N_10798,N_9609,N_9075);
and U10799 (N_10799,N_9047,N_9334);
or U10800 (N_10800,N_9624,N_9802);
xor U10801 (N_10801,N_9287,N_9799);
nor U10802 (N_10802,N_9763,N_9670);
or U10803 (N_10803,N_9639,N_9605);
or U10804 (N_10804,N_9128,N_9087);
xnor U10805 (N_10805,N_9191,N_9523);
and U10806 (N_10806,N_9258,N_9519);
or U10807 (N_10807,N_9348,N_9262);
nand U10808 (N_10808,N_9202,N_9168);
nand U10809 (N_10809,N_9132,N_9429);
and U10810 (N_10810,N_9242,N_9537);
nand U10811 (N_10811,N_9076,N_9010);
xnor U10812 (N_10812,N_9611,N_9775);
and U10813 (N_10813,N_9074,N_9801);
xor U10814 (N_10814,N_9367,N_9655);
or U10815 (N_10815,N_9421,N_9075);
nand U10816 (N_10816,N_9289,N_9726);
nor U10817 (N_10817,N_9122,N_9137);
nand U10818 (N_10818,N_9603,N_9618);
and U10819 (N_10819,N_9963,N_9264);
nand U10820 (N_10820,N_9683,N_9075);
nand U10821 (N_10821,N_9721,N_9221);
xor U10822 (N_10822,N_9853,N_9344);
and U10823 (N_10823,N_9217,N_9226);
nand U10824 (N_10824,N_9659,N_9208);
xor U10825 (N_10825,N_9074,N_9827);
nand U10826 (N_10826,N_9439,N_9367);
nand U10827 (N_10827,N_9040,N_9660);
nand U10828 (N_10828,N_9616,N_9482);
nor U10829 (N_10829,N_9637,N_9014);
nor U10830 (N_10830,N_9761,N_9524);
and U10831 (N_10831,N_9093,N_9108);
nand U10832 (N_10832,N_9505,N_9126);
or U10833 (N_10833,N_9752,N_9101);
or U10834 (N_10834,N_9956,N_9409);
xnor U10835 (N_10835,N_9941,N_9539);
nor U10836 (N_10836,N_9033,N_9901);
nand U10837 (N_10837,N_9609,N_9151);
xor U10838 (N_10838,N_9668,N_9813);
nand U10839 (N_10839,N_9133,N_9968);
nor U10840 (N_10840,N_9724,N_9837);
or U10841 (N_10841,N_9517,N_9337);
xor U10842 (N_10842,N_9407,N_9924);
or U10843 (N_10843,N_9395,N_9824);
nand U10844 (N_10844,N_9447,N_9011);
xnor U10845 (N_10845,N_9330,N_9086);
and U10846 (N_10846,N_9495,N_9505);
and U10847 (N_10847,N_9974,N_9900);
or U10848 (N_10848,N_9418,N_9727);
or U10849 (N_10849,N_9336,N_9026);
nor U10850 (N_10850,N_9269,N_9135);
nor U10851 (N_10851,N_9908,N_9223);
nor U10852 (N_10852,N_9782,N_9394);
xor U10853 (N_10853,N_9041,N_9245);
xor U10854 (N_10854,N_9973,N_9682);
or U10855 (N_10855,N_9163,N_9954);
or U10856 (N_10856,N_9598,N_9859);
and U10857 (N_10857,N_9586,N_9604);
and U10858 (N_10858,N_9118,N_9741);
and U10859 (N_10859,N_9947,N_9876);
and U10860 (N_10860,N_9228,N_9672);
nor U10861 (N_10861,N_9868,N_9165);
nor U10862 (N_10862,N_9614,N_9998);
and U10863 (N_10863,N_9015,N_9010);
and U10864 (N_10864,N_9240,N_9189);
and U10865 (N_10865,N_9304,N_9517);
and U10866 (N_10866,N_9952,N_9064);
nor U10867 (N_10867,N_9058,N_9782);
nor U10868 (N_10868,N_9570,N_9744);
nand U10869 (N_10869,N_9509,N_9706);
nor U10870 (N_10870,N_9074,N_9154);
nor U10871 (N_10871,N_9050,N_9585);
nor U10872 (N_10872,N_9628,N_9851);
or U10873 (N_10873,N_9199,N_9459);
or U10874 (N_10874,N_9137,N_9731);
or U10875 (N_10875,N_9544,N_9616);
nor U10876 (N_10876,N_9857,N_9171);
nand U10877 (N_10877,N_9967,N_9750);
nand U10878 (N_10878,N_9672,N_9026);
or U10879 (N_10879,N_9792,N_9047);
or U10880 (N_10880,N_9546,N_9176);
or U10881 (N_10881,N_9821,N_9312);
and U10882 (N_10882,N_9573,N_9347);
nor U10883 (N_10883,N_9439,N_9324);
nor U10884 (N_10884,N_9643,N_9837);
nand U10885 (N_10885,N_9732,N_9854);
nand U10886 (N_10886,N_9394,N_9009);
xnor U10887 (N_10887,N_9365,N_9895);
and U10888 (N_10888,N_9780,N_9267);
and U10889 (N_10889,N_9587,N_9162);
nand U10890 (N_10890,N_9379,N_9020);
and U10891 (N_10891,N_9514,N_9995);
xor U10892 (N_10892,N_9886,N_9435);
and U10893 (N_10893,N_9321,N_9796);
and U10894 (N_10894,N_9898,N_9396);
or U10895 (N_10895,N_9922,N_9705);
xnor U10896 (N_10896,N_9602,N_9109);
or U10897 (N_10897,N_9206,N_9652);
xor U10898 (N_10898,N_9229,N_9580);
xor U10899 (N_10899,N_9555,N_9144);
xnor U10900 (N_10900,N_9582,N_9727);
xor U10901 (N_10901,N_9176,N_9263);
or U10902 (N_10902,N_9564,N_9728);
or U10903 (N_10903,N_9680,N_9142);
xnor U10904 (N_10904,N_9306,N_9666);
nor U10905 (N_10905,N_9481,N_9742);
nor U10906 (N_10906,N_9722,N_9319);
nand U10907 (N_10907,N_9742,N_9565);
xnor U10908 (N_10908,N_9593,N_9922);
and U10909 (N_10909,N_9000,N_9876);
or U10910 (N_10910,N_9760,N_9350);
xor U10911 (N_10911,N_9513,N_9093);
nand U10912 (N_10912,N_9942,N_9357);
xnor U10913 (N_10913,N_9007,N_9941);
nand U10914 (N_10914,N_9495,N_9247);
nand U10915 (N_10915,N_9493,N_9720);
or U10916 (N_10916,N_9601,N_9666);
or U10917 (N_10917,N_9723,N_9135);
nand U10918 (N_10918,N_9846,N_9868);
nand U10919 (N_10919,N_9544,N_9277);
nor U10920 (N_10920,N_9673,N_9216);
and U10921 (N_10921,N_9070,N_9466);
xnor U10922 (N_10922,N_9435,N_9444);
nand U10923 (N_10923,N_9907,N_9414);
nand U10924 (N_10924,N_9646,N_9963);
nor U10925 (N_10925,N_9730,N_9657);
nor U10926 (N_10926,N_9352,N_9146);
xnor U10927 (N_10927,N_9573,N_9607);
and U10928 (N_10928,N_9635,N_9199);
nor U10929 (N_10929,N_9116,N_9055);
and U10930 (N_10930,N_9970,N_9026);
nand U10931 (N_10931,N_9051,N_9291);
and U10932 (N_10932,N_9804,N_9328);
nand U10933 (N_10933,N_9750,N_9703);
and U10934 (N_10934,N_9053,N_9500);
nand U10935 (N_10935,N_9317,N_9293);
nor U10936 (N_10936,N_9644,N_9251);
or U10937 (N_10937,N_9016,N_9017);
or U10938 (N_10938,N_9854,N_9845);
xor U10939 (N_10939,N_9203,N_9954);
xor U10940 (N_10940,N_9519,N_9130);
xnor U10941 (N_10941,N_9747,N_9103);
xnor U10942 (N_10942,N_9280,N_9845);
or U10943 (N_10943,N_9952,N_9970);
and U10944 (N_10944,N_9621,N_9020);
nand U10945 (N_10945,N_9044,N_9445);
or U10946 (N_10946,N_9210,N_9905);
nor U10947 (N_10947,N_9661,N_9346);
or U10948 (N_10948,N_9586,N_9596);
nand U10949 (N_10949,N_9791,N_9400);
nor U10950 (N_10950,N_9522,N_9861);
xor U10951 (N_10951,N_9095,N_9789);
and U10952 (N_10952,N_9614,N_9565);
nor U10953 (N_10953,N_9289,N_9535);
xnor U10954 (N_10954,N_9899,N_9574);
nor U10955 (N_10955,N_9306,N_9532);
nand U10956 (N_10956,N_9511,N_9275);
nand U10957 (N_10957,N_9980,N_9080);
nand U10958 (N_10958,N_9984,N_9428);
nand U10959 (N_10959,N_9398,N_9907);
or U10960 (N_10960,N_9431,N_9104);
nand U10961 (N_10961,N_9702,N_9950);
and U10962 (N_10962,N_9861,N_9929);
and U10963 (N_10963,N_9433,N_9874);
and U10964 (N_10964,N_9819,N_9632);
nand U10965 (N_10965,N_9260,N_9819);
and U10966 (N_10966,N_9636,N_9169);
nor U10967 (N_10967,N_9678,N_9139);
or U10968 (N_10968,N_9827,N_9413);
and U10969 (N_10969,N_9851,N_9397);
or U10970 (N_10970,N_9994,N_9031);
nand U10971 (N_10971,N_9838,N_9457);
and U10972 (N_10972,N_9755,N_9776);
nand U10973 (N_10973,N_9649,N_9276);
nor U10974 (N_10974,N_9279,N_9192);
xor U10975 (N_10975,N_9466,N_9262);
xnor U10976 (N_10976,N_9293,N_9915);
nand U10977 (N_10977,N_9458,N_9608);
or U10978 (N_10978,N_9701,N_9983);
xnor U10979 (N_10979,N_9757,N_9852);
nor U10980 (N_10980,N_9650,N_9224);
xnor U10981 (N_10981,N_9122,N_9101);
and U10982 (N_10982,N_9446,N_9974);
nand U10983 (N_10983,N_9512,N_9520);
and U10984 (N_10984,N_9140,N_9393);
and U10985 (N_10985,N_9347,N_9060);
xor U10986 (N_10986,N_9574,N_9219);
or U10987 (N_10987,N_9547,N_9942);
and U10988 (N_10988,N_9340,N_9115);
xnor U10989 (N_10989,N_9381,N_9171);
nand U10990 (N_10990,N_9702,N_9221);
or U10991 (N_10991,N_9437,N_9123);
nor U10992 (N_10992,N_9086,N_9249);
nor U10993 (N_10993,N_9801,N_9778);
nand U10994 (N_10994,N_9583,N_9991);
or U10995 (N_10995,N_9632,N_9805);
nand U10996 (N_10996,N_9290,N_9079);
nand U10997 (N_10997,N_9383,N_9053);
xnor U10998 (N_10998,N_9575,N_9036);
and U10999 (N_10999,N_9121,N_9932);
and U11000 (N_11000,N_10826,N_10943);
xor U11001 (N_11001,N_10131,N_10992);
or U11002 (N_11002,N_10337,N_10734);
nor U11003 (N_11003,N_10580,N_10909);
nor U11004 (N_11004,N_10209,N_10723);
nand U11005 (N_11005,N_10850,N_10170);
and U11006 (N_11006,N_10299,N_10304);
xnor U11007 (N_11007,N_10585,N_10387);
nand U11008 (N_11008,N_10285,N_10417);
nand U11009 (N_11009,N_10410,N_10265);
or U11010 (N_11010,N_10748,N_10957);
xor U11011 (N_11011,N_10628,N_10513);
nor U11012 (N_11012,N_10276,N_10956);
and U11013 (N_11013,N_10418,N_10253);
or U11014 (N_11014,N_10964,N_10538);
xor U11015 (N_11015,N_10504,N_10042);
nand U11016 (N_11016,N_10548,N_10078);
nor U11017 (N_11017,N_10446,N_10901);
xor U11018 (N_11018,N_10604,N_10981);
and U11019 (N_11019,N_10185,N_10004);
or U11020 (N_11020,N_10737,N_10799);
nand U11021 (N_11021,N_10949,N_10771);
nor U11022 (N_11022,N_10411,N_10512);
nor U11023 (N_11023,N_10983,N_10684);
nor U11024 (N_11024,N_10573,N_10184);
nor U11025 (N_11025,N_10447,N_10026);
nand U11026 (N_11026,N_10007,N_10867);
and U11027 (N_11027,N_10180,N_10136);
nor U11028 (N_11028,N_10827,N_10062);
nand U11029 (N_11029,N_10646,N_10414);
xor U11030 (N_11030,N_10287,N_10741);
nand U11031 (N_11031,N_10950,N_10670);
or U11032 (N_11032,N_10899,N_10219);
or U11033 (N_11033,N_10444,N_10743);
nor U11034 (N_11034,N_10961,N_10437);
xor U11035 (N_11035,N_10478,N_10526);
nor U11036 (N_11036,N_10313,N_10627);
nor U11037 (N_11037,N_10134,N_10652);
nor U11038 (N_11038,N_10671,N_10699);
nand U11039 (N_11039,N_10858,N_10532);
or U11040 (N_11040,N_10255,N_10631);
and U11041 (N_11041,N_10552,N_10896);
or U11042 (N_11042,N_10404,N_10861);
and U11043 (N_11043,N_10075,N_10354);
xnor U11044 (N_11044,N_10519,N_10084);
and U11045 (N_11045,N_10231,N_10856);
xor U11046 (N_11046,N_10929,N_10874);
nand U11047 (N_11047,N_10505,N_10844);
xor U11048 (N_11048,N_10939,N_10716);
nand U11049 (N_11049,N_10173,N_10675);
nor U11050 (N_11050,N_10308,N_10088);
xor U11051 (N_11051,N_10830,N_10800);
nor U11052 (N_11052,N_10987,N_10686);
and U11053 (N_11053,N_10730,N_10360);
nand U11054 (N_11054,N_10434,N_10306);
and U11055 (N_11055,N_10566,N_10539);
and U11056 (N_11056,N_10297,N_10208);
or U11057 (N_11057,N_10782,N_10727);
nand U11058 (N_11058,N_10973,N_10791);
nand U11059 (N_11059,N_10935,N_10216);
and U11060 (N_11060,N_10873,N_10608);
and U11061 (N_11061,N_10009,N_10419);
nor U11062 (N_11062,N_10919,N_10128);
or U11063 (N_11063,N_10379,N_10839);
or U11064 (N_11064,N_10768,N_10402);
or U11065 (N_11065,N_10393,N_10481);
or U11066 (N_11066,N_10385,N_10784);
xnor U11067 (N_11067,N_10897,N_10930);
xnor U11068 (N_11068,N_10609,N_10192);
nand U11069 (N_11069,N_10661,N_10408);
nor U11070 (N_11070,N_10559,N_10579);
nand U11071 (N_11071,N_10963,N_10266);
nand U11072 (N_11072,N_10605,N_10491);
nand U11073 (N_11073,N_10178,N_10698);
nand U11074 (N_11074,N_10564,N_10642);
or U11075 (N_11075,N_10857,N_10917);
and U11076 (N_11076,N_10483,N_10130);
nor U11077 (N_11077,N_10141,N_10568);
or U11078 (N_11078,N_10112,N_10468);
and U11079 (N_11079,N_10195,N_10588);
xnor U11080 (N_11080,N_10091,N_10116);
nor U11081 (N_11081,N_10341,N_10429);
xnor U11082 (N_11082,N_10061,N_10168);
or U11083 (N_11083,N_10347,N_10140);
nand U11084 (N_11084,N_10601,N_10327);
and U11085 (N_11085,N_10912,N_10904);
nor U11086 (N_11086,N_10531,N_10701);
or U11087 (N_11087,N_10704,N_10119);
or U11088 (N_11088,N_10056,N_10537);
xnor U11089 (N_11089,N_10754,N_10355);
and U11090 (N_11090,N_10106,N_10103);
or U11091 (N_11091,N_10044,N_10794);
nor U11092 (N_11092,N_10320,N_10878);
or U11093 (N_11093,N_10480,N_10043);
nand U11094 (N_11094,N_10953,N_10148);
nand U11095 (N_11095,N_10045,N_10174);
nand U11096 (N_11096,N_10616,N_10895);
nor U11097 (N_11097,N_10490,N_10375);
or U11098 (N_11098,N_10825,N_10651);
nand U11099 (N_11099,N_10779,N_10450);
nand U11100 (N_11100,N_10115,N_10703);
nor U11101 (N_11101,N_10251,N_10037);
xor U11102 (N_11102,N_10584,N_10028);
and U11103 (N_11103,N_10016,N_10254);
nand U11104 (N_11104,N_10332,N_10127);
nor U11105 (N_11105,N_10546,N_10525);
nand U11106 (N_11106,N_10558,N_10259);
nand U11107 (N_11107,N_10169,N_10882);
nor U11108 (N_11108,N_10193,N_10911);
and U11109 (N_11109,N_10612,N_10098);
nor U11110 (N_11110,N_10465,N_10994);
or U11111 (N_11111,N_10625,N_10866);
or U11112 (N_11112,N_10053,N_10638);
and U11113 (N_11113,N_10773,N_10440);
or U11114 (N_11114,N_10654,N_10680);
nor U11115 (N_11115,N_10070,N_10795);
nor U11116 (N_11116,N_10475,N_10836);
or U11117 (N_11117,N_10808,N_10221);
and U11118 (N_11118,N_10906,N_10439);
nor U11119 (N_11119,N_10790,N_10988);
and U11120 (N_11120,N_10035,N_10213);
nand U11121 (N_11121,N_10373,N_10067);
nand U11122 (N_11122,N_10821,N_10818);
and U11123 (N_11123,N_10555,N_10143);
or U11124 (N_11124,N_10835,N_10346);
nor U11125 (N_11125,N_10606,N_10298);
or U11126 (N_11126,N_10740,N_10416);
xnor U11127 (N_11127,N_10838,N_10382);
xor U11128 (N_11128,N_10508,N_10712);
or U11129 (N_11129,N_10139,N_10977);
and U11130 (N_11130,N_10217,N_10095);
nor U11131 (N_11131,N_10931,N_10292);
nor U11132 (N_11132,N_10990,N_10649);
xnor U11133 (N_11133,N_10235,N_10146);
xnor U11134 (N_11134,N_10218,N_10717);
xnor U11135 (N_11135,N_10695,N_10284);
nand U11136 (N_11136,N_10430,N_10557);
xor U11137 (N_11137,N_10370,N_10516);
and U11138 (N_11138,N_10186,N_10828);
xnor U11139 (N_11139,N_10226,N_10592);
or U11140 (N_11140,N_10694,N_10772);
or U11141 (N_11141,N_10003,N_10029);
nor U11142 (N_11142,N_10805,N_10980);
nand U11143 (N_11143,N_10995,N_10693);
or U11144 (N_11144,N_10275,N_10248);
xor U11145 (N_11145,N_10300,N_10732);
nor U11146 (N_11146,N_10747,N_10665);
nor U11147 (N_11147,N_10421,N_10842);
or U11148 (N_11148,N_10560,N_10542);
nand U11149 (N_11149,N_10764,N_10073);
xnor U11150 (N_11150,N_10510,N_10877);
nand U11151 (N_11151,N_10780,N_10362);
nor U11152 (N_11152,N_10735,N_10643);
and U11153 (N_11153,N_10966,N_10984);
xor U11154 (N_11154,N_10600,N_10775);
xor U11155 (N_11155,N_10426,N_10239);
nor U11156 (N_11156,N_10569,N_10249);
and U11157 (N_11157,N_10309,N_10707);
and U11158 (N_11158,N_10294,N_10114);
or U11159 (N_11159,N_10025,N_10286);
xnor U11160 (N_11160,N_10348,N_10484);
nor U11161 (N_11161,N_10677,N_10145);
nor U11162 (N_11162,N_10664,N_10894);
nand U11163 (N_11163,N_10345,N_10824);
nor U11164 (N_11164,N_10224,N_10590);
and U11165 (N_11165,N_10296,N_10445);
xor U11166 (N_11166,N_10455,N_10024);
nor U11167 (N_11167,N_10496,N_10083);
xor U11168 (N_11168,N_10229,N_10926);
or U11169 (N_11169,N_10371,N_10859);
nand U11170 (N_11170,N_10036,N_10910);
nor U11171 (N_11171,N_10972,N_10692);
or U11172 (N_11172,N_10968,N_10122);
and U11173 (N_11173,N_10562,N_10241);
xor U11174 (N_11174,N_10970,N_10498);
xnor U11175 (N_11175,N_10602,N_10637);
nor U11176 (N_11176,N_10100,N_10689);
or U11177 (N_11177,N_10936,N_10524);
and U11178 (N_11178,N_10204,N_10428);
xor U11179 (N_11179,N_10520,N_10399);
or U11180 (N_11180,N_10001,N_10094);
nor U11181 (N_11181,N_10817,N_10583);
and U11182 (N_11182,N_10365,N_10745);
nor U11183 (N_11183,N_10515,N_10788);
and U11184 (N_11184,N_10215,N_10565);
nor U11185 (N_11185,N_10381,N_10395);
xnor U11186 (N_11186,N_10948,N_10924);
nand U11187 (N_11187,N_10998,N_10305);
nor U11188 (N_11188,N_10974,N_10205);
xor U11189 (N_11189,N_10540,N_10242);
nand U11190 (N_11190,N_10080,N_10914);
nand U11191 (N_11191,N_10787,N_10182);
or U11192 (N_11192,N_10349,N_10572);
and U11193 (N_11193,N_10645,N_10617);
nand U11194 (N_11194,N_10576,N_10700);
nor U11195 (N_11195,N_10211,N_10751);
xnor U11196 (N_11196,N_10847,N_10040);
nor U11197 (N_11197,N_10815,N_10641);
nand U11198 (N_11198,N_10702,N_10422);
and U11199 (N_11199,N_10372,N_10786);
nand U11200 (N_11200,N_10006,N_10511);
nor U11201 (N_11201,N_10487,N_10685);
or U11202 (N_11202,N_10636,N_10884);
nor U11203 (N_11203,N_10340,N_10622);
or U11204 (N_11204,N_10763,N_10769);
xor U11205 (N_11205,N_10027,N_10172);
nand U11206 (N_11206,N_10030,N_10472);
xor U11207 (N_11207,N_10368,N_10944);
nand U11208 (N_11208,N_10879,N_10262);
and U11209 (N_11209,N_10753,N_10158);
nor U11210 (N_11210,N_10367,N_10869);
xnor U11211 (N_11211,N_10117,N_10733);
xor U11212 (N_11212,N_10766,N_10054);
xnor U11213 (N_11213,N_10055,N_10196);
xor U11214 (N_11214,N_10156,N_10999);
nor U11215 (N_11215,N_10234,N_10626);
nor U11216 (N_11216,N_10384,N_10840);
xor U11217 (N_11217,N_10683,N_10060);
nand U11218 (N_11218,N_10871,N_10603);
or U11219 (N_11219,N_10497,N_10749);
nor U11220 (N_11220,N_10263,N_10005);
and U11221 (N_11221,N_10507,N_10150);
xor U11222 (N_11222,N_10473,N_10377);
xnor U11223 (N_11223,N_10587,N_10048);
xor U11224 (N_11224,N_10339,N_10523);
nor U11225 (N_11225,N_10288,N_10389);
or U11226 (N_11226,N_10104,N_10407);
xor U11227 (N_11227,N_10233,N_10462);
and U11228 (N_11228,N_10778,N_10971);
or U11229 (N_11229,N_10765,N_10880);
and U11230 (N_11230,N_10783,N_10570);
nor U11231 (N_11231,N_10102,N_10726);
xnor U11232 (N_11232,N_10635,N_10925);
and U11233 (N_11233,N_10049,N_10915);
nor U11234 (N_11234,N_10967,N_10489);
or U11235 (N_11235,N_10464,N_10181);
nor U11236 (N_11236,N_10798,N_10191);
nand U11237 (N_11237,N_10085,N_10619);
nand U11238 (N_11238,N_10829,N_10744);
xnor U11239 (N_11239,N_10503,N_10492);
xor U11240 (N_11240,N_10868,N_10722);
and U11241 (N_11241,N_10357,N_10133);
and U11242 (N_11242,N_10438,N_10920);
nor U11243 (N_11243,N_10678,N_10290);
nor U11244 (N_11244,N_10656,N_10281);
and U11245 (N_11245,N_10162,N_10068);
or U11246 (N_11246,N_10841,N_10057);
nor U11247 (N_11247,N_10323,N_10586);
or U11248 (N_11248,N_10846,N_10237);
nor U11249 (N_11249,N_10853,N_10900);
and U11250 (N_11250,N_10796,N_10789);
and U11251 (N_11251,N_10982,N_10463);
nor U11252 (N_11252,N_10289,N_10738);
xnor U11253 (N_11253,N_10750,N_10940);
or U11254 (N_11254,N_10731,N_10223);
and U11255 (N_11255,N_10330,N_10965);
xnor U11256 (N_11256,N_10301,N_10849);
xnor U11257 (N_11257,N_10653,N_10500);
nand U11258 (N_11258,N_10630,N_10436);
or U11259 (N_11259,N_10351,N_10757);
and U11260 (N_11260,N_10659,N_10321);
xnor U11261 (N_11261,N_10124,N_10812);
nor U11262 (N_11262,N_10166,N_10177);
or U11263 (N_11263,N_10724,N_10081);
or U11264 (N_11264,N_10008,N_10629);
nor U11265 (N_11265,N_10050,N_10711);
xor U11266 (N_11266,N_10872,N_10891);
nor U11267 (N_11267,N_10898,N_10495);
and U11268 (N_11268,N_10942,N_10014);
xor U11269 (N_11269,N_10441,N_10502);
or U11270 (N_11270,N_10640,N_10390);
nor U11271 (N_11271,N_10614,N_10041);
or U11272 (N_11272,N_10230,N_10012);
nand U11273 (N_11273,N_10530,N_10454);
or U11274 (N_11274,N_10848,N_10681);
nand U11275 (N_11275,N_10203,N_10739);
and U11276 (N_11276,N_10047,N_10257);
and U11277 (N_11277,N_10620,N_10535);
xnor U11278 (N_11278,N_10383,N_10427);
nand U11279 (N_11279,N_10220,N_10243);
nand U11280 (N_11280,N_10250,N_10096);
or U11281 (N_11281,N_10344,N_10819);
or U11282 (N_11282,N_10244,N_10621);
xor U11283 (N_11283,N_10425,N_10352);
nor U11284 (N_11284,N_10975,N_10493);
nand U11285 (N_11285,N_10946,N_10907);
nor U11286 (N_11286,N_10563,N_10415);
and U11287 (N_11287,N_10167,N_10721);
and U11288 (N_11288,N_10142,N_10655);
nor U11289 (N_11289,N_10138,N_10593);
nor U11290 (N_11290,N_10669,N_10863);
or U11291 (N_11291,N_10792,N_10713);
nand U11292 (N_11292,N_10623,N_10589);
or U11293 (N_11293,N_10715,N_10212);
and U11294 (N_11294,N_10129,N_10277);
nor U11295 (N_11295,N_10577,N_10801);
nor U11296 (N_11296,N_10160,N_10811);
nor U11297 (N_11297,N_10802,N_10804);
or U11298 (N_11298,N_10273,N_10561);
or U11299 (N_11299,N_10860,N_10916);
or U11300 (N_11300,N_10256,N_10082);
xnor U11301 (N_11301,N_10820,N_10864);
xor U11302 (N_11302,N_10756,N_10709);
xnor U11303 (N_11303,N_10110,N_10401);
nor U11304 (N_11304,N_10315,N_10391);
and U11305 (N_11305,N_10065,N_10159);
or U11306 (N_11306,N_10807,N_10350);
or U11307 (N_11307,N_10227,N_10282);
nand U11308 (N_11308,N_10663,N_10163);
nand U11309 (N_11309,N_10574,N_10528);
nand U11310 (N_11310,N_10550,N_10118);
or U11311 (N_11311,N_10696,N_10245);
xor U11312 (N_11312,N_10232,N_10071);
nand U11313 (N_11313,N_10010,N_10658);
nor U11314 (N_11314,N_10509,N_10597);
xnor U11315 (N_11315,N_10400,N_10571);
nand U11316 (N_11316,N_10615,N_10985);
or U11317 (N_11317,N_10499,N_10039);
nor U11318 (N_11318,N_10596,N_10072);
nor U11319 (N_11319,N_10816,N_10144);
or U11320 (N_11320,N_10189,N_10923);
nand U11321 (N_11321,N_10137,N_10889);
nand U11322 (N_11322,N_10222,N_10545);
nand U11323 (N_11323,N_10761,N_10632);
xnor U11324 (N_11324,N_10161,N_10945);
and U11325 (N_11325,N_10890,N_10918);
nand U11326 (N_11326,N_10870,N_10153);
or U11327 (N_11327,N_10011,N_10022);
and U11328 (N_11328,N_10435,N_10312);
nor U11329 (N_11329,N_10618,N_10363);
and U11330 (N_11330,N_10554,N_10742);
xnor U11331 (N_11331,N_10886,N_10902);
nor U11332 (N_11332,N_10852,N_10020);
nand U11333 (N_11333,N_10679,N_10536);
nand U11334 (N_11334,N_10947,N_10470);
and U11335 (N_11335,N_10278,N_10113);
nor U11336 (N_11336,N_10392,N_10591);
nor U11337 (N_11337,N_10398,N_10431);
xor U11338 (N_11338,N_10674,N_10486);
or U11339 (N_11339,N_10171,N_10449);
nor U11340 (N_11340,N_10806,N_10522);
nor U11341 (N_11341,N_10461,N_10595);
nor U11342 (N_11342,N_10017,N_10214);
nor U11343 (N_11343,N_10729,N_10302);
nor U11344 (N_11344,N_10506,N_10667);
and U11345 (N_11345,N_10720,N_10610);
and U11346 (N_11346,N_10776,N_10228);
and U11347 (N_11347,N_10324,N_10932);
nand U11348 (N_11348,N_10823,N_10314);
nand U11349 (N_11349,N_10079,N_10076);
xnor U11350 (N_11350,N_10543,N_10388);
xnor U11351 (N_11351,N_10814,N_10272);
or U11352 (N_11352,N_10018,N_10225);
xnor U11353 (N_11353,N_10032,N_10969);
and U11354 (N_11354,N_10803,N_10760);
and U11355 (N_11355,N_10708,N_10316);
nand U11356 (N_11356,N_10238,N_10594);
nand U11357 (N_11357,N_10941,N_10951);
nor U11358 (N_11358,N_10993,N_10329);
nand U11359 (N_11359,N_10295,N_10291);
nand U11360 (N_11360,N_10364,N_10485);
or U11361 (N_11361,N_10903,N_10333);
or U11362 (N_11362,N_10705,N_10855);
nand U11363 (N_11363,N_10267,N_10002);
nand U11364 (N_11364,N_10752,N_10567);
or U11365 (N_11365,N_10876,N_10187);
or U11366 (N_11366,N_10905,N_10200);
nand U11367 (N_11367,N_10443,N_10885);
and U11368 (N_11368,N_10660,N_10319);
xor U11369 (N_11369,N_10527,N_10843);
nor U11370 (N_11370,N_10466,N_10013);
and U11371 (N_11371,N_10544,N_10063);
nand U11372 (N_11372,N_10714,N_10471);
or U11373 (N_11373,N_10353,N_10413);
nand U11374 (N_11374,N_10922,N_10101);
or U11375 (N_11375,N_10240,N_10976);
and U11376 (N_11376,N_10000,N_10270);
nor U11377 (N_11377,N_10832,N_10328);
and U11378 (N_11378,N_10342,N_10376);
xnor U11379 (N_11379,N_10386,N_10672);
and U11380 (N_11380,N_10962,N_10958);
nor U11381 (N_11381,N_10599,N_10706);
xor U11382 (N_11382,N_10448,N_10725);
nand U11383 (N_11383,N_10074,N_10986);
or U11384 (N_11384,N_10322,N_10433);
xor U11385 (N_11385,N_10154,N_10152);
and U11386 (N_11386,N_10837,N_10865);
and U11387 (N_11387,N_10318,N_10822);
and U11388 (N_11388,N_10774,N_10378);
nor U11389 (N_11389,N_10303,N_10335);
xor U11390 (N_11390,N_10126,N_10607);
nor U11391 (N_11391,N_10657,N_10058);
nand U11392 (N_11392,N_10533,N_10111);
nor U11393 (N_11393,N_10691,N_10165);
nor U11394 (N_11394,N_10147,N_10633);
and U11395 (N_11395,N_10650,N_10469);
or U11396 (N_11396,N_10467,N_10666);
nor U11397 (N_11397,N_10356,N_10274);
nor U11398 (N_11398,N_10097,N_10477);
nor U11399 (N_11399,N_10934,N_10207);
and U11400 (N_11400,N_10718,N_10412);
xnor U11401 (N_11401,N_10258,N_10598);
nand U11402 (N_11402,N_10668,N_10135);
and U11403 (N_11403,N_10210,N_10662);
nand U11404 (N_11404,N_10206,N_10246);
xnor U11405 (N_11405,N_10514,N_10394);
or U11406 (N_11406,N_10123,N_10893);
or U11407 (N_11407,N_10978,N_10359);
nor U11408 (N_11408,N_10758,N_10268);
nor U11409 (N_11409,N_10746,N_10881);
nand U11410 (N_11410,N_10613,N_10781);
nor U11411 (N_11411,N_10959,N_10052);
nand U11412 (N_11412,N_10845,N_10770);
or U11413 (N_11413,N_10336,N_10397);
or U11414 (N_11414,N_10201,N_10093);
nor U11415 (N_11415,N_10575,N_10374);
nand U11416 (N_11416,N_10019,N_10451);
xnor U11417 (N_11417,N_10883,N_10927);
or U11418 (N_11418,N_10199,N_10938);
or U11419 (N_11419,N_10979,N_10611);
xor U11420 (N_11420,N_10908,N_10405);
and U11421 (N_11421,N_10190,N_10236);
nand U11422 (N_11422,N_10547,N_10033);
xnor U11423 (N_11423,N_10458,N_10380);
and U11424 (N_11424,N_10120,N_10090);
or U11425 (N_11425,N_10283,N_10494);
and U11426 (N_11426,N_10697,N_10247);
or U11427 (N_11427,N_10317,N_10517);
and U11428 (N_11428,N_10719,N_10409);
nor U11429 (N_11429,N_10797,N_10423);
and U11430 (N_11430,N_10762,N_10155);
xor U11431 (N_11431,N_10534,N_10997);
or U11432 (N_11432,N_10457,N_10887);
or U11433 (N_11433,N_10260,N_10459);
nor U11434 (N_11434,N_10366,N_10077);
and U11435 (N_11435,N_10064,N_10179);
and U11436 (N_11436,N_10676,N_10086);
and U11437 (N_11437,N_10673,N_10046);
or U11438 (N_11438,N_10755,N_10479);
or U11439 (N_11439,N_10269,N_10125);
and U11440 (N_11440,N_10687,N_10518);
or U11441 (N_11441,N_10087,N_10183);
xor U11442 (N_11442,N_10913,N_10813);
and U11443 (N_11443,N_10474,N_10157);
or U11444 (N_11444,N_10488,N_10928);
and U11445 (N_11445,N_10059,N_10264);
or U11446 (N_11446,N_10175,N_10460);
nand U11447 (N_11447,N_10151,N_10293);
or U11448 (N_11448,N_10767,N_10176);
or U11449 (N_11449,N_10015,N_10326);
nor U11450 (N_11450,N_10482,N_10875);
and U11451 (N_11451,N_10279,N_10785);
nor U11452 (N_11452,N_10777,N_10476);
or U11453 (N_11453,N_10862,N_10952);
or U11454 (N_11454,N_10442,N_10271);
and U11455 (N_11455,N_10107,N_10325);
nor U11456 (N_11456,N_10810,N_10023);
and U11457 (N_11457,N_10149,N_10452);
nand U11458 (N_11458,N_10338,N_10954);
nand U11459 (N_11459,N_10736,N_10644);
nor U11460 (N_11460,N_10038,N_10834);
nor U11461 (N_11461,N_10202,N_10021);
xor U11462 (N_11462,N_10682,N_10089);
or U11463 (N_11463,N_10501,N_10541);
or U11464 (N_11464,N_10759,N_10034);
nor U11465 (N_11465,N_10937,N_10578);
or U11466 (N_11466,N_10261,N_10582);
or U11467 (N_11467,N_10099,N_10809);
or U11468 (N_11468,N_10647,N_10996);
xor U11469 (N_11469,N_10358,N_10854);
nand U11470 (N_11470,N_10132,N_10311);
nor U11471 (N_11471,N_10690,N_10793);
and U11472 (N_11472,N_10551,N_10553);
xor U11473 (N_11473,N_10432,N_10105);
nand U11474 (N_11474,N_10066,N_10403);
nor U11475 (N_11475,N_10710,N_10989);
nand U11476 (N_11476,N_10197,N_10307);
nor U11477 (N_11477,N_10092,N_10648);
xor U11478 (N_11478,N_10198,N_10639);
or U11479 (N_11479,N_10406,N_10833);
and U11480 (N_11480,N_10343,N_10556);
and U11481 (N_11481,N_10194,N_10334);
or U11482 (N_11482,N_10188,N_10121);
or U11483 (N_11483,N_10361,N_10831);
or U11484 (N_11484,N_10109,N_10420);
nand U11485 (N_11485,N_10521,N_10252);
nor U11486 (N_11486,N_10634,N_10921);
xor U11487 (N_11487,N_10955,N_10456);
xor U11488 (N_11488,N_10331,N_10892);
and U11489 (N_11489,N_10728,N_10164);
or U11490 (N_11490,N_10529,N_10688);
nor U11491 (N_11491,N_10624,N_10108);
xnor U11492 (N_11492,N_10310,N_10888);
xnor U11493 (N_11493,N_10396,N_10453);
or U11494 (N_11494,N_10424,N_10991);
xor U11495 (N_11495,N_10933,N_10280);
and U11496 (N_11496,N_10851,N_10069);
or U11497 (N_11497,N_10051,N_10549);
and U11498 (N_11498,N_10369,N_10581);
nand U11499 (N_11499,N_10960,N_10031);
or U11500 (N_11500,N_10107,N_10441);
xor U11501 (N_11501,N_10986,N_10377);
xor U11502 (N_11502,N_10713,N_10377);
and U11503 (N_11503,N_10261,N_10186);
and U11504 (N_11504,N_10451,N_10875);
nand U11505 (N_11505,N_10454,N_10607);
nor U11506 (N_11506,N_10178,N_10021);
or U11507 (N_11507,N_10651,N_10119);
nand U11508 (N_11508,N_10587,N_10701);
nor U11509 (N_11509,N_10089,N_10185);
nand U11510 (N_11510,N_10110,N_10511);
nor U11511 (N_11511,N_10521,N_10606);
or U11512 (N_11512,N_10932,N_10668);
or U11513 (N_11513,N_10263,N_10814);
nand U11514 (N_11514,N_10593,N_10754);
nand U11515 (N_11515,N_10346,N_10554);
xnor U11516 (N_11516,N_10643,N_10219);
xor U11517 (N_11517,N_10789,N_10774);
or U11518 (N_11518,N_10870,N_10439);
xor U11519 (N_11519,N_10326,N_10116);
and U11520 (N_11520,N_10551,N_10795);
and U11521 (N_11521,N_10678,N_10861);
xor U11522 (N_11522,N_10112,N_10244);
nand U11523 (N_11523,N_10874,N_10188);
nand U11524 (N_11524,N_10132,N_10978);
nand U11525 (N_11525,N_10740,N_10493);
nand U11526 (N_11526,N_10234,N_10479);
or U11527 (N_11527,N_10588,N_10657);
or U11528 (N_11528,N_10205,N_10694);
nand U11529 (N_11529,N_10856,N_10620);
xnor U11530 (N_11530,N_10640,N_10909);
nor U11531 (N_11531,N_10855,N_10160);
xnor U11532 (N_11532,N_10310,N_10520);
and U11533 (N_11533,N_10016,N_10998);
and U11534 (N_11534,N_10091,N_10819);
nand U11535 (N_11535,N_10084,N_10766);
or U11536 (N_11536,N_10707,N_10749);
xor U11537 (N_11537,N_10359,N_10314);
xnor U11538 (N_11538,N_10707,N_10759);
and U11539 (N_11539,N_10846,N_10946);
xnor U11540 (N_11540,N_10648,N_10205);
nor U11541 (N_11541,N_10363,N_10447);
nor U11542 (N_11542,N_10913,N_10194);
nor U11543 (N_11543,N_10044,N_10184);
nand U11544 (N_11544,N_10366,N_10432);
nand U11545 (N_11545,N_10972,N_10015);
nor U11546 (N_11546,N_10343,N_10188);
nand U11547 (N_11547,N_10310,N_10457);
and U11548 (N_11548,N_10494,N_10127);
nor U11549 (N_11549,N_10180,N_10934);
nor U11550 (N_11550,N_10648,N_10118);
xnor U11551 (N_11551,N_10779,N_10550);
nor U11552 (N_11552,N_10737,N_10111);
nand U11553 (N_11553,N_10862,N_10961);
or U11554 (N_11554,N_10218,N_10800);
nor U11555 (N_11555,N_10400,N_10157);
nand U11556 (N_11556,N_10502,N_10075);
or U11557 (N_11557,N_10273,N_10150);
and U11558 (N_11558,N_10005,N_10872);
xor U11559 (N_11559,N_10575,N_10748);
nand U11560 (N_11560,N_10508,N_10565);
and U11561 (N_11561,N_10251,N_10970);
xnor U11562 (N_11562,N_10526,N_10032);
nor U11563 (N_11563,N_10435,N_10674);
or U11564 (N_11564,N_10153,N_10260);
nor U11565 (N_11565,N_10259,N_10625);
or U11566 (N_11566,N_10754,N_10606);
xnor U11567 (N_11567,N_10066,N_10994);
xor U11568 (N_11568,N_10662,N_10990);
nor U11569 (N_11569,N_10129,N_10992);
or U11570 (N_11570,N_10339,N_10234);
nand U11571 (N_11571,N_10699,N_10141);
or U11572 (N_11572,N_10584,N_10394);
xnor U11573 (N_11573,N_10819,N_10037);
nor U11574 (N_11574,N_10874,N_10526);
and U11575 (N_11575,N_10913,N_10999);
nand U11576 (N_11576,N_10876,N_10605);
xnor U11577 (N_11577,N_10409,N_10991);
xnor U11578 (N_11578,N_10191,N_10613);
or U11579 (N_11579,N_10976,N_10282);
nor U11580 (N_11580,N_10306,N_10325);
nor U11581 (N_11581,N_10824,N_10417);
nand U11582 (N_11582,N_10894,N_10817);
nand U11583 (N_11583,N_10891,N_10869);
or U11584 (N_11584,N_10482,N_10232);
nand U11585 (N_11585,N_10102,N_10793);
and U11586 (N_11586,N_10007,N_10653);
nand U11587 (N_11587,N_10096,N_10187);
or U11588 (N_11588,N_10790,N_10673);
nand U11589 (N_11589,N_10536,N_10293);
xor U11590 (N_11590,N_10072,N_10444);
nand U11591 (N_11591,N_10290,N_10885);
or U11592 (N_11592,N_10745,N_10309);
and U11593 (N_11593,N_10919,N_10289);
xor U11594 (N_11594,N_10409,N_10277);
xnor U11595 (N_11595,N_10959,N_10593);
xor U11596 (N_11596,N_10098,N_10686);
nand U11597 (N_11597,N_10854,N_10256);
xor U11598 (N_11598,N_10567,N_10612);
or U11599 (N_11599,N_10188,N_10756);
nor U11600 (N_11600,N_10796,N_10079);
xnor U11601 (N_11601,N_10043,N_10798);
nand U11602 (N_11602,N_10844,N_10653);
xnor U11603 (N_11603,N_10416,N_10863);
nor U11604 (N_11604,N_10116,N_10042);
nor U11605 (N_11605,N_10273,N_10501);
and U11606 (N_11606,N_10760,N_10857);
xnor U11607 (N_11607,N_10434,N_10524);
and U11608 (N_11608,N_10026,N_10210);
nor U11609 (N_11609,N_10842,N_10534);
nand U11610 (N_11610,N_10387,N_10431);
xor U11611 (N_11611,N_10158,N_10066);
nand U11612 (N_11612,N_10702,N_10563);
xor U11613 (N_11613,N_10001,N_10713);
nor U11614 (N_11614,N_10518,N_10045);
or U11615 (N_11615,N_10245,N_10388);
xnor U11616 (N_11616,N_10316,N_10423);
nor U11617 (N_11617,N_10464,N_10706);
xor U11618 (N_11618,N_10460,N_10392);
or U11619 (N_11619,N_10934,N_10223);
xnor U11620 (N_11620,N_10583,N_10596);
or U11621 (N_11621,N_10666,N_10672);
nand U11622 (N_11622,N_10766,N_10541);
xnor U11623 (N_11623,N_10784,N_10064);
nand U11624 (N_11624,N_10168,N_10893);
or U11625 (N_11625,N_10706,N_10517);
and U11626 (N_11626,N_10728,N_10989);
nand U11627 (N_11627,N_10251,N_10573);
nand U11628 (N_11628,N_10136,N_10893);
and U11629 (N_11629,N_10086,N_10404);
and U11630 (N_11630,N_10328,N_10194);
xnor U11631 (N_11631,N_10686,N_10339);
nor U11632 (N_11632,N_10689,N_10524);
xor U11633 (N_11633,N_10943,N_10279);
nand U11634 (N_11634,N_10470,N_10116);
xnor U11635 (N_11635,N_10006,N_10409);
or U11636 (N_11636,N_10943,N_10730);
or U11637 (N_11637,N_10649,N_10316);
nand U11638 (N_11638,N_10433,N_10809);
xnor U11639 (N_11639,N_10232,N_10444);
nand U11640 (N_11640,N_10597,N_10469);
nand U11641 (N_11641,N_10587,N_10851);
xor U11642 (N_11642,N_10916,N_10263);
or U11643 (N_11643,N_10504,N_10701);
or U11644 (N_11644,N_10803,N_10211);
xnor U11645 (N_11645,N_10946,N_10532);
nand U11646 (N_11646,N_10096,N_10138);
or U11647 (N_11647,N_10701,N_10942);
nor U11648 (N_11648,N_10240,N_10790);
xor U11649 (N_11649,N_10111,N_10984);
nand U11650 (N_11650,N_10096,N_10453);
or U11651 (N_11651,N_10240,N_10261);
nand U11652 (N_11652,N_10367,N_10313);
nand U11653 (N_11653,N_10192,N_10104);
or U11654 (N_11654,N_10481,N_10734);
or U11655 (N_11655,N_10448,N_10729);
xor U11656 (N_11656,N_10072,N_10797);
nand U11657 (N_11657,N_10194,N_10873);
nand U11658 (N_11658,N_10093,N_10237);
and U11659 (N_11659,N_10332,N_10248);
xnor U11660 (N_11660,N_10168,N_10221);
nand U11661 (N_11661,N_10308,N_10856);
and U11662 (N_11662,N_10751,N_10266);
and U11663 (N_11663,N_10449,N_10288);
and U11664 (N_11664,N_10926,N_10075);
or U11665 (N_11665,N_10713,N_10890);
nand U11666 (N_11666,N_10643,N_10733);
and U11667 (N_11667,N_10809,N_10326);
nand U11668 (N_11668,N_10200,N_10892);
or U11669 (N_11669,N_10584,N_10421);
xnor U11670 (N_11670,N_10502,N_10276);
xor U11671 (N_11671,N_10665,N_10293);
and U11672 (N_11672,N_10553,N_10396);
and U11673 (N_11673,N_10722,N_10715);
nand U11674 (N_11674,N_10441,N_10718);
nand U11675 (N_11675,N_10171,N_10835);
nor U11676 (N_11676,N_10962,N_10287);
xor U11677 (N_11677,N_10386,N_10437);
or U11678 (N_11678,N_10286,N_10023);
and U11679 (N_11679,N_10779,N_10545);
xor U11680 (N_11680,N_10287,N_10793);
and U11681 (N_11681,N_10213,N_10986);
xor U11682 (N_11682,N_10613,N_10599);
nor U11683 (N_11683,N_10454,N_10884);
xnor U11684 (N_11684,N_10971,N_10590);
nor U11685 (N_11685,N_10947,N_10621);
nor U11686 (N_11686,N_10235,N_10504);
and U11687 (N_11687,N_10672,N_10653);
nor U11688 (N_11688,N_10008,N_10045);
nand U11689 (N_11689,N_10083,N_10673);
nor U11690 (N_11690,N_10057,N_10898);
nor U11691 (N_11691,N_10162,N_10537);
xnor U11692 (N_11692,N_10222,N_10383);
or U11693 (N_11693,N_10366,N_10920);
or U11694 (N_11694,N_10634,N_10660);
nor U11695 (N_11695,N_10227,N_10754);
xor U11696 (N_11696,N_10941,N_10025);
xnor U11697 (N_11697,N_10015,N_10897);
nor U11698 (N_11698,N_10119,N_10250);
and U11699 (N_11699,N_10602,N_10431);
and U11700 (N_11700,N_10478,N_10439);
xor U11701 (N_11701,N_10545,N_10930);
or U11702 (N_11702,N_10107,N_10609);
nand U11703 (N_11703,N_10874,N_10529);
nand U11704 (N_11704,N_10009,N_10608);
xor U11705 (N_11705,N_10245,N_10047);
xnor U11706 (N_11706,N_10257,N_10540);
xor U11707 (N_11707,N_10533,N_10701);
nor U11708 (N_11708,N_10073,N_10779);
and U11709 (N_11709,N_10368,N_10355);
or U11710 (N_11710,N_10763,N_10053);
or U11711 (N_11711,N_10156,N_10482);
xor U11712 (N_11712,N_10247,N_10569);
or U11713 (N_11713,N_10986,N_10710);
and U11714 (N_11714,N_10861,N_10478);
and U11715 (N_11715,N_10412,N_10706);
nand U11716 (N_11716,N_10666,N_10920);
or U11717 (N_11717,N_10004,N_10802);
nand U11718 (N_11718,N_10783,N_10896);
xor U11719 (N_11719,N_10726,N_10817);
nor U11720 (N_11720,N_10759,N_10309);
and U11721 (N_11721,N_10663,N_10418);
or U11722 (N_11722,N_10910,N_10136);
xnor U11723 (N_11723,N_10017,N_10071);
nor U11724 (N_11724,N_10641,N_10229);
nand U11725 (N_11725,N_10650,N_10414);
xor U11726 (N_11726,N_10147,N_10163);
xor U11727 (N_11727,N_10990,N_10701);
or U11728 (N_11728,N_10591,N_10340);
or U11729 (N_11729,N_10715,N_10942);
and U11730 (N_11730,N_10823,N_10926);
nand U11731 (N_11731,N_10544,N_10552);
and U11732 (N_11732,N_10838,N_10585);
and U11733 (N_11733,N_10581,N_10413);
and U11734 (N_11734,N_10580,N_10945);
nand U11735 (N_11735,N_10190,N_10958);
or U11736 (N_11736,N_10840,N_10827);
or U11737 (N_11737,N_10795,N_10760);
nand U11738 (N_11738,N_10499,N_10395);
or U11739 (N_11739,N_10190,N_10805);
xor U11740 (N_11740,N_10568,N_10979);
nor U11741 (N_11741,N_10379,N_10362);
nor U11742 (N_11742,N_10749,N_10615);
xnor U11743 (N_11743,N_10126,N_10756);
and U11744 (N_11744,N_10189,N_10913);
or U11745 (N_11745,N_10595,N_10736);
nand U11746 (N_11746,N_10196,N_10077);
nor U11747 (N_11747,N_10690,N_10988);
nand U11748 (N_11748,N_10282,N_10831);
nor U11749 (N_11749,N_10991,N_10681);
or U11750 (N_11750,N_10898,N_10713);
nor U11751 (N_11751,N_10948,N_10159);
or U11752 (N_11752,N_10167,N_10967);
nand U11753 (N_11753,N_10040,N_10932);
nand U11754 (N_11754,N_10195,N_10087);
or U11755 (N_11755,N_10174,N_10755);
nor U11756 (N_11756,N_10519,N_10109);
and U11757 (N_11757,N_10963,N_10102);
xnor U11758 (N_11758,N_10700,N_10923);
and U11759 (N_11759,N_10782,N_10443);
nand U11760 (N_11760,N_10643,N_10065);
xor U11761 (N_11761,N_10593,N_10319);
or U11762 (N_11762,N_10559,N_10729);
nor U11763 (N_11763,N_10954,N_10242);
nand U11764 (N_11764,N_10783,N_10687);
nand U11765 (N_11765,N_10785,N_10164);
or U11766 (N_11766,N_10702,N_10588);
or U11767 (N_11767,N_10126,N_10114);
or U11768 (N_11768,N_10056,N_10020);
xnor U11769 (N_11769,N_10370,N_10878);
or U11770 (N_11770,N_10662,N_10062);
or U11771 (N_11771,N_10309,N_10689);
or U11772 (N_11772,N_10109,N_10360);
or U11773 (N_11773,N_10671,N_10189);
or U11774 (N_11774,N_10366,N_10963);
nand U11775 (N_11775,N_10387,N_10056);
nor U11776 (N_11776,N_10526,N_10522);
nor U11777 (N_11777,N_10501,N_10174);
or U11778 (N_11778,N_10771,N_10090);
and U11779 (N_11779,N_10884,N_10970);
nor U11780 (N_11780,N_10781,N_10407);
nor U11781 (N_11781,N_10926,N_10657);
and U11782 (N_11782,N_10191,N_10080);
and U11783 (N_11783,N_10468,N_10961);
nand U11784 (N_11784,N_10522,N_10464);
nand U11785 (N_11785,N_10024,N_10866);
or U11786 (N_11786,N_10238,N_10127);
nor U11787 (N_11787,N_10177,N_10531);
or U11788 (N_11788,N_10318,N_10722);
and U11789 (N_11789,N_10235,N_10917);
or U11790 (N_11790,N_10176,N_10413);
and U11791 (N_11791,N_10883,N_10107);
nor U11792 (N_11792,N_10464,N_10973);
and U11793 (N_11793,N_10490,N_10099);
nand U11794 (N_11794,N_10520,N_10358);
nand U11795 (N_11795,N_10288,N_10930);
nand U11796 (N_11796,N_10913,N_10616);
and U11797 (N_11797,N_10211,N_10554);
nand U11798 (N_11798,N_10227,N_10318);
and U11799 (N_11799,N_10465,N_10154);
nor U11800 (N_11800,N_10874,N_10890);
and U11801 (N_11801,N_10789,N_10752);
xor U11802 (N_11802,N_10133,N_10293);
xor U11803 (N_11803,N_10816,N_10449);
nand U11804 (N_11804,N_10452,N_10087);
or U11805 (N_11805,N_10385,N_10566);
xnor U11806 (N_11806,N_10592,N_10696);
or U11807 (N_11807,N_10388,N_10686);
nor U11808 (N_11808,N_10040,N_10944);
and U11809 (N_11809,N_10802,N_10438);
or U11810 (N_11810,N_10295,N_10450);
nand U11811 (N_11811,N_10942,N_10659);
nand U11812 (N_11812,N_10049,N_10256);
nand U11813 (N_11813,N_10568,N_10212);
or U11814 (N_11814,N_10410,N_10178);
nand U11815 (N_11815,N_10104,N_10708);
nor U11816 (N_11816,N_10388,N_10437);
or U11817 (N_11817,N_10232,N_10723);
and U11818 (N_11818,N_10114,N_10488);
nor U11819 (N_11819,N_10507,N_10679);
or U11820 (N_11820,N_10929,N_10274);
and U11821 (N_11821,N_10345,N_10788);
nand U11822 (N_11822,N_10742,N_10345);
xor U11823 (N_11823,N_10424,N_10768);
or U11824 (N_11824,N_10646,N_10561);
nor U11825 (N_11825,N_10024,N_10009);
and U11826 (N_11826,N_10897,N_10097);
or U11827 (N_11827,N_10895,N_10730);
nor U11828 (N_11828,N_10050,N_10403);
or U11829 (N_11829,N_10649,N_10874);
nor U11830 (N_11830,N_10163,N_10213);
and U11831 (N_11831,N_10674,N_10868);
nand U11832 (N_11832,N_10155,N_10514);
and U11833 (N_11833,N_10040,N_10693);
nand U11834 (N_11834,N_10303,N_10884);
xnor U11835 (N_11835,N_10345,N_10063);
or U11836 (N_11836,N_10511,N_10406);
or U11837 (N_11837,N_10348,N_10894);
nand U11838 (N_11838,N_10878,N_10188);
or U11839 (N_11839,N_10952,N_10355);
and U11840 (N_11840,N_10424,N_10001);
nand U11841 (N_11841,N_10231,N_10708);
nor U11842 (N_11842,N_10696,N_10573);
nand U11843 (N_11843,N_10814,N_10027);
nor U11844 (N_11844,N_10786,N_10888);
or U11845 (N_11845,N_10031,N_10016);
nand U11846 (N_11846,N_10235,N_10609);
xor U11847 (N_11847,N_10885,N_10489);
or U11848 (N_11848,N_10891,N_10487);
nor U11849 (N_11849,N_10652,N_10256);
xor U11850 (N_11850,N_10974,N_10654);
xnor U11851 (N_11851,N_10032,N_10530);
nor U11852 (N_11852,N_10071,N_10895);
and U11853 (N_11853,N_10683,N_10998);
nand U11854 (N_11854,N_10494,N_10181);
and U11855 (N_11855,N_10312,N_10358);
or U11856 (N_11856,N_10248,N_10777);
or U11857 (N_11857,N_10197,N_10814);
nor U11858 (N_11858,N_10283,N_10153);
xor U11859 (N_11859,N_10133,N_10234);
nand U11860 (N_11860,N_10272,N_10030);
xnor U11861 (N_11861,N_10847,N_10417);
xor U11862 (N_11862,N_10274,N_10575);
and U11863 (N_11863,N_10569,N_10428);
or U11864 (N_11864,N_10283,N_10750);
xnor U11865 (N_11865,N_10190,N_10434);
or U11866 (N_11866,N_10907,N_10123);
nor U11867 (N_11867,N_10515,N_10901);
or U11868 (N_11868,N_10595,N_10168);
xor U11869 (N_11869,N_10898,N_10186);
or U11870 (N_11870,N_10312,N_10723);
and U11871 (N_11871,N_10289,N_10151);
nand U11872 (N_11872,N_10870,N_10967);
nand U11873 (N_11873,N_10442,N_10860);
nor U11874 (N_11874,N_10431,N_10391);
or U11875 (N_11875,N_10745,N_10542);
or U11876 (N_11876,N_10961,N_10956);
or U11877 (N_11877,N_10808,N_10790);
or U11878 (N_11878,N_10069,N_10232);
or U11879 (N_11879,N_10473,N_10481);
and U11880 (N_11880,N_10270,N_10674);
and U11881 (N_11881,N_10971,N_10095);
nand U11882 (N_11882,N_10270,N_10029);
and U11883 (N_11883,N_10775,N_10708);
and U11884 (N_11884,N_10315,N_10072);
nand U11885 (N_11885,N_10307,N_10709);
or U11886 (N_11886,N_10310,N_10935);
or U11887 (N_11887,N_10150,N_10317);
xnor U11888 (N_11888,N_10513,N_10460);
nand U11889 (N_11889,N_10678,N_10770);
and U11890 (N_11890,N_10780,N_10640);
nand U11891 (N_11891,N_10449,N_10700);
nand U11892 (N_11892,N_10359,N_10368);
nor U11893 (N_11893,N_10711,N_10729);
nor U11894 (N_11894,N_10767,N_10334);
nand U11895 (N_11895,N_10942,N_10895);
xnor U11896 (N_11896,N_10543,N_10391);
nand U11897 (N_11897,N_10230,N_10778);
nor U11898 (N_11898,N_10454,N_10214);
and U11899 (N_11899,N_10706,N_10582);
or U11900 (N_11900,N_10380,N_10713);
xnor U11901 (N_11901,N_10429,N_10556);
nand U11902 (N_11902,N_10272,N_10845);
xor U11903 (N_11903,N_10641,N_10450);
and U11904 (N_11904,N_10295,N_10843);
xnor U11905 (N_11905,N_10531,N_10022);
or U11906 (N_11906,N_10395,N_10813);
or U11907 (N_11907,N_10369,N_10118);
xor U11908 (N_11908,N_10812,N_10420);
or U11909 (N_11909,N_10174,N_10486);
nor U11910 (N_11910,N_10719,N_10642);
xor U11911 (N_11911,N_10462,N_10946);
nor U11912 (N_11912,N_10070,N_10851);
nor U11913 (N_11913,N_10313,N_10473);
nand U11914 (N_11914,N_10977,N_10155);
and U11915 (N_11915,N_10951,N_10777);
nor U11916 (N_11916,N_10657,N_10836);
or U11917 (N_11917,N_10457,N_10810);
nor U11918 (N_11918,N_10501,N_10392);
nand U11919 (N_11919,N_10098,N_10498);
and U11920 (N_11920,N_10802,N_10936);
nand U11921 (N_11921,N_10247,N_10755);
or U11922 (N_11922,N_10854,N_10269);
or U11923 (N_11923,N_10955,N_10367);
and U11924 (N_11924,N_10212,N_10650);
and U11925 (N_11925,N_10820,N_10647);
nor U11926 (N_11926,N_10124,N_10225);
xor U11927 (N_11927,N_10053,N_10617);
nand U11928 (N_11928,N_10054,N_10303);
nor U11929 (N_11929,N_10122,N_10348);
nand U11930 (N_11930,N_10709,N_10500);
nand U11931 (N_11931,N_10677,N_10761);
or U11932 (N_11932,N_10098,N_10257);
or U11933 (N_11933,N_10944,N_10967);
or U11934 (N_11934,N_10335,N_10471);
and U11935 (N_11935,N_10189,N_10098);
nand U11936 (N_11936,N_10706,N_10395);
or U11937 (N_11937,N_10756,N_10128);
nor U11938 (N_11938,N_10163,N_10581);
nand U11939 (N_11939,N_10476,N_10450);
and U11940 (N_11940,N_10594,N_10622);
nand U11941 (N_11941,N_10381,N_10585);
and U11942 (N_11942,N_10537,N_10448);
or U11943 (N_11943,N_10944,N_10494);
nor U11944 (N_11944,N_10110,N_10669);
and U11945 (N_11945,N_10330,N_10337);
nor U11946 (N_11946,N_10321,N_10388);
or U11947 (N_11947,N_10830,N_10886);
nand U11948 (N_11948,N_10267,N_10574);
nand U11949 (N_11949,N_10767,N_10949);
xor U11950 (N_11950,N_10928,N_10579);
nand U11951 (N_11951,N_10318,N_10321);
nand U11952 (N_11952,N_10539,N_10985);
nor U11953 (N_11953,N_10469,N_10877);
and U11954 (N_11954,N_10248,N_10102);
or U11955 (N_11955,N_10807,N_10624);
nand U11956 (N_11956,N_10094,N_10337);
and U11957 (N_11957,N_10588,N_10124);
and U11958 (N_11958,N_10417,N_10248);
nand U11959 (N_11959,N_10705,N_10989);
nor U11960 (N_11960,N_10947,N_10861);
and U11961 (N_11961,N_10451,N_10361);
xor U11962 (N_11962,N_10051,N_10947);
nor U11963 (N_11963,N_10642,N_10943);
nand U11964 (N_11964,N_10320,N_10784);
nor U11965 (N_11965,N_10625,N_10638);
nor U11966 (N_11966,N_10954,N_10037);
nand U11967 (N_11967,N_10417,N_10498);
xnor U11968 (N_11968,N_10384,N_10715);
or U11969 (N_11969,N_10196,N_10514);
nor U11970 (N_11970,N_10468,N_10698);
and U11971 (N_11971,N_10130,N_10069);
nand U11972 (N_11972,N_10369,N_10105);
nor U11973 (N_11973,N_10586,N_10164);
xor U11974 (N_11974,N_10112,N_10868);
nor U11975 (N_11975,N_10230,N_10709);
nand U11976 (N_11976,N_10913,N_10577);
nor U11977 (N_11977,N_10444,N_10247);
nand U11978 (N_11978,N_10918,N_10583);
or U11979 (N_11979,N_10225,N_10950);
nor U11980 (N_11980,N_10983,N_10699);
nor U11981 (N_11981,N_10958,N_10555);
xnor U11982 (N_11982,N_10516,N_10827);
nor U11983 (N_11983,N_10507,N_10757);
nand U11984 (N_11984,N_10754,N_10930);
xor U11985 (N_11985,N_10197,N_10911);
or U11986 (N_11986,N_10187,N_10835);
xnor U11987 (N_11987,N_10325,N_10493);
or U11988 (N_11988,N_10045,N_10177);
and U11989 (N_11989,N_10229,N_10692);
xor U11990 (N_11990,N_10291,N_10432);
and U11991 (N_11991,N_10089,N_10487);
and U11992 (N_11992,N_10901,N_10410);
and U11993 (N_11993,N_10037,N_10412);
nand U11994 (N_11994,N_10718,N_10568);
and U11995 (N_11995,N_10412,N_10128);
or U11996 (N_11996,N_10467,N_10411);
xnor U11997 (N_11997,N_10636,N_10168);
and U11998 (N_11998,N_10614,N_10669);
nor U11999 (N_11999,N_10848,N_10753);
xor U12000 (N_12000,N_11390,N_11137);
and U12001 (N_12001,N_11914,N_11686);
xnor U12002 (N_12002,N_11095,N_11804);
nor U12003 (N_12003,N_11967,N_11813);
and U12004 (N_12004,N_11668,N_11036);
nand U12005 (N_12005,N_11171,N_11466);
or U12006 (N_12006,N_11208,N_11975);
and U12007 (N_12007,N_11381,N_11379);
xnor U12008 (N_12008,N_11159,N_11770);
nor U12009 (N_12009,N_11020,N_11559);
nor U12010 (N_12010,N_11446,N_11657);
nand U12011 (N_12011,N_11439,N_11653);
or U12012 (N_12012,N_11553,N_11160);
xnor U12013 (N_12013,N_11806,N_11364);
and U12014 (N_12014,N_11085,N_11516);
or U12015 (N_12015,N_11180,N_11628);
nor U12016 (N_12016,N_11512,N_11838);
and U12017 (N_12017,N_11972,N_11795);
xnor U12018 (N_12018,N_11651,N_11754);
or U12019 (N_12019,N_11099,N_11848);
nor U12020 (N_12020,N_11461,N_11735);
nand U12021 (N_12021,N_11859,N_11501);
xnor U12022 (N_12022,N_11755,N_11699);
nand U12023 (N_12023,N_11278,N_11384);
or U12024 (N_12024,N_11345,N_11410);
xnor U12025 (N_12025,N_11986,N_11822);
or U12026 (N_12026,N_11059,N_11084);
nand U12027 (N_12027,N_11122,N_11569);
nand U12028 (N_12028,N_11323,N_11295);
xor U12029 (N_12029,N_11376,N_11109);
nor U12030 (N_12030,N_11332,N_11832);
or U12031 (N_12031,N_11337,N_11005);
and U12032 (N_12032,N_11163,N_11850);
nand U12033 (N_12033,N_11945,N_11821);
nor U12034 (N_12034,N_11719,N_11488);
and U12035 (N_12035,N_11871,N_11080);
xnor U12036 (N_12036,N_11522,N_11387);
and U12037 (N_12037,N_11851,N_11389);
and U12038 (N_12038,N_11016,N_11878);
or U12039 (N_12039,N_11973,N_11294);
nand U12040 (N_12040,N_11175,N_11117);
xnor U12041 (N_12041,N_11333,N_11862);
and U12042 (N_12042,N_11460,N_11268);
xor U12043 (N_12043,N_11775,N_11010);
or U12044 (N_12044,N_11713,N_11803);
and U12045 (N_12045,N_11716,N_11105);
and U12046 (N_12046,N_11664,N_11618);
xnor U12047 (N_12047,N_11107,N_11328);
nor U12048 (N_12048,N_11207,N_11074);
and U12049 (N_12049,N_11251,N_11982);
xor U12050 (N_12050,N_11825,N_11591);
or U12051 (N_12051,N_11079,N_11856);
or U12052 (N_12052,N_11827,N_11070);
and U12053 (N_12053,N_11032,N_11585);
nand U12054 (N_12054,N_11378,N_11284);
nand U12055 (N_12055,N_11923,N_11638);
nand U12056 (N_12056,N_11527,N_11318);
nor U12057 (N_12057,N_11508,N_11181);
nor U12058 (N_12058,N_11613,N_11210);
nor U12059 (N_12059,N_11089,N_11015);
nand U12060 (N_12060,N_11214,N_11977);
xnor U12061 (N_12061,N_11458,N_11550);
nand U12062 (N_12062,N_11455,N_11584);
or U12063 (N_12063,N_11991,N_11437);
xor U12064 (N_12064,N_11740,N_11952);
or U12065 (N_12065,N_11313,N_11001);
and U12066 (N_12066,N_11994,N_11477);
nor U12067 (N_12067,N_11843,N_11216);
nor U12068 (N_12068,N_11906,N_11700);
nor U12069 (N_12069,N_11561,N_11348);
and U12070 (N_12070,N_11291,N_11336);
and U12071 (N_12071,N_11281,N_11218);
nor U12072 (N_12072,N_11111,N_11257);
and U12073 (N_12073,N_11691,N_11764);
nand U12074 (N_12074,N_11509,N_11314);
or U12075 (N_12075,N_11583,N_11480);
and U12076 (N_12076,N_11063,N_11282);
or U12077 (N_12077,N_11671,N_11274);
and U12078 (N_12078,N_11834,N_11593);
or U12079 (N_12079,N_11418,N_11252);
xnor U12080 (N_12080,N_11510,N_11647);
nor U12081 (N_12081,N_11129,N_11103);
nor U12082 (N_12082,N_11718,N_11534);
nor U12083 (N_12083,N_11457,N_11845);
nor U12084 (N_12084,N_11641,N_11202);
or U12085 (N_12085,N_11570,N_11762);
and U12086 (N_12086,N_11022,N_11260);
xor U12087 (N_12087,N_11000,N_11658);
nand U12088 (N_12088,N_11443,N_11685);
and U12089 (N_12089,N_11748,N_11721);
nand U12090 (N_12090,N_11701,N_11689);
and U12091 (N_12091,N_11785,N_11893);
and U12092 (N_12092,N_11168,N_11717);
or U12093 (N_12093,N_11830,N_11956);
or U12094 (N_12094,N_11520,N_11909);
or U12095 (N_12095,N_11223,N_11092);
nor U12096 (N_12096,N_11027,N_11662);
xnor U12097 (N_12097,N_11007,N_11736);
nor U12098 (N_12098,N_11088,N_11616);
and U12099 (N_12099,N_11247,N_11575);
nand U12100 (N_12100,N_11130,N_11529);
xnor U12101 (N_12101,N_11212,N_11245);
or U12102 (N_12102,N_11363,N_11953);
or U12103 (N_12103,N_11886,N_11263);
or U12104 (N_12104,N_11265,N_11548);
nor U12105 (N_12105,N_11943,N_11530);
and U12106 (N_12106,N_11732,N_11523);
or U12107 (N_12107,N_11044,N_11841);
nand U12108 (N_12108,N_11349,N_11746);
or U12109 (N_12109,N_11517,N_11928);
xor U12110 (N_12110,N_11401,N_11026);
xnor U12111 (N_12111,N_11629,N_11555);
xor U12112 (N_12112,N_11852,N_11327);
and U12113 (N_12113,N_11744,N_11004);
nor U12114 (N_12114,N_11441,N_11743);
nor U12115 (N_12115,N_11579,N_11558);
or U12116 (N_12116,N_11675,N_11126);
and U12117 (N_12117,N_11377,N_11478);
or U12118 (N_12118,N_11464,N_11149);
nor U12119 (N_12119,N_11091,N_11786);
nand U12120 (N_12120,N_11935,N_11391);
and U12121 (N_12121,N_11541,N_11087);
or U12122 (N_12122,N_11759,N_11229);
nand U12123 (N_12123,N_11823,N_11898);
xnor U12124 (N_12124,N_11793,N_11836);
nand U12125 (N_12125,N_11152,N_11304);
and U12126 (N_12126,N_11649,N_11614);
xor U12127 (N_12127,N_11602,N_11609);
xor U12128 (N_12128,N_11076,N_11404);
xnor U12129 (N_12129,N_11896,N_11521);
xnor U12130 (N_12130,N_11166,N_11722);
and U12131 (N_12131,N_11046,N_11842);
nand U12132 (N_12132,N_11577,N_11114);
nor U12133 (N_12133,N_11456,N_11903);
nor U12134 (N_12134,N_11796,N_11101);
nor U12135 (N_12135,N_11473,N_11969);
or U12136 (N_12136,N_11885,N_11269);
nand U12137 (N_12137,N_11761,N_11853);
nand U12138 (N_12138,N_11778,N_11492);
xnor U12139 (N_12139,N_11985,N_11409);
nand U12140 (N_12140,N_11623,N_11396);
xor U12141 (N_12141,N_11965,N_11217);
or U12142 (N_12142,N_11835,N_11715);
and U12143 (N_12143,N_11067,N_11366);
nand U12144 (N_12144,N_11680,N_11470);
or U12145 (N_12145,N_11147,N_11193);
nor U12146 (N_12146,N_11753,N_11589);
nor U12147 (N_12147,N_11383,N_11050);
and U12148 (N_12148,N_11727,N_11188);
nor U12149 (N_12149,N_11014,N_11312);
or U12150 (N_12150,N_11317,N_11739);
xor U12151 (N_12151,N_11465,N_11599);
xor U12152 (N_12152,N_11695,N_11201);
nor U12153 (N_12153,N_11902,N_11655);
nand U12154 (N_12154,N_11343,N_11479);
and U12155 (N_12155,N_11447,N_11055);
or U12156 (N_12156,N_11272,N_11980);
xor U12157 (N_12157,N_11497,N_11119);
nor U12158 (N_12158,N_11400,N_11385);
nand U12159 (N_12159,N_11146,N_11824);
and U12160 (N_12160,N_11531,N_11243);
xnor U12161 (N_12161,N_11372,N_11543);
or U12162 (N_12162,N_11249,N_11929);
xor U12163 (N_12163,N_11681,N_11904);
nor U12164 (N_12164,N_11678,N_11254);
and U12165 (N_12165,N_11308,N_11426);
nand U12166 (N_12166,N_11043,N_11434);
nor U12167 (N_12167,N_11264,N_11725);
or U12168 (N_12168,N_11078,N_11205);
xor U12169 (N_12169,N_11692,N_11820);
xor U12170 (N_12170,N_11406,N_11781);
nand U12171 (N_12171,N_11472,N_11276);
or U12172 (N_12172,N_11791,N_11932);
xnor U12173 (N_12173,N_11397,N_11917);
nor U12174 (N_12174,N_11978,N_11515);
and U12175 (N_12175,N_11809,N_11169);
xor U12176 (N_12176,N_11773,N_11302);
or U12177 (N_12177,N_11948,N_11897);
xnor U12178 (N_12178,N_11086,N_11155);
and U12179 (N_12179,N_11135,N_11224);
or U12180 (N_12180,N_11448,N_11936);
or U12181 (N_12181,N_11197,N_11780);
or U12182 (N_12182,N_11857,N_11937);
and U12183 (N_12183,N_11233,N_11697);
nor U12184 (N_12184,N_11419,N_11560);
and U12185 (N_12185,N_11427,N_11631);
xnor U12186 (N_12186,N_11047,N_11394);
xnor U12187 (N_12187,N_11525,N_11557);
and U12188 (N_12188,N_11676,N_11944);
xor U12189 (N_12189,N_11632,N_11963);
nor U12190 (N_12190,N_11374,N_11993);
and U12191 (N_12191,N_11979,N_11301);
or U12192 (N_12192,N_11187,N_11453);
or U12193 (N_12193,N_11483,N_11590);
nor U12194 (N_12194,N_11061,N_11330);
nor U12195 (N_12195,N_11369,N_11942);
nand U12196 (N_12196,N_11325,N_11872);
xnor U12197 (N_12197,N_11742,N_11910);
xor U12198 (N_12198,N_11062,N_11905);
or U12199 (N_12199,N_11090,N_11927);
nor U12200 (N_12200,N_11572,N_11424);
or U12201 (N_12201,N_11661,N_11745);
xnor U12202 (N_12202,N_11826,N_11604);
and U12203 (N_12203,N_11574,N_11037);
and U12204 (N_12204,N_11578,N_11918);
or U12205 (N_12205,N_11733,N_11194);
nor U12206 (N_12206,N_11056,N_11006);
nand U12207 (N_12207,N_11771,N_11633);
nor U12208 (N_12208,N_11064,N_11949);
nor U12209 (N_12209,N_11462,N_11749);
xor U12210 (N_12210,N_11630,N_11815);
xor U12211 (N_12211,N_11113,N_11913);
nand U12212 (N_12212,N_11452,N_11476);
nand U12213 (N_12213,N_11941,N_11648);
nor U12214 (N_12214,N_11542,N_11758);
xor U12215 (N_12215,N_11884,N_11173);
or U12216 (N_12216,N_11615,N_11141);
nand U12217 (N_12217,N_11075,N_11204);
nor U12218 (N_12218,N_11601,N_11860);
nor U12219 (N_12219,N_11164,N_11428);
and U12220 (N_12220,N_11329,N_11679);
nor U12221 (N_12221,N_11189,N_11990);
nor U12222 (N_12222,N_11592,N_11066);
xor U12223 (N_12223,N_11507,N_11262);
or U12224 (N_12224,N_11855,N_11696);
xnor U12225 (N_12225,N_11386,N_11782);
nor U12226 (N_12226,N_11854,N_11463);
xnor U12227 (N_12227,N_11354,N_11726);
xnor U12228 (N_12228,N_11964,N_11071);
nand U12229 (N_12229,N_11494,N_11068);
nor U12230 (N_12230,N_11720,N_11586);
nand U12231 (N_12231,N_11132,N_11467);
or U12232 (N_12232,N_11203,N_11874);
xor U12233 (N_12233,N_11535,N_11118);
or U12234 (N_12234,N_11545,N_11013);
or U12235 (N_12235,N_11106,N_11421);
xnor U12236 (N_12236,N_11232,N_11236);
or U12237 (N_12237,N_11162,N_11959);
and U12238 (N_12238,N_11607,N_11285);
xnor U12239 (N_12239,N_11837,N_11346);
nand U12240 (N_12240,N_11420,N_11347);
xor U12241 (N_12241,N_11481,N_11298);
or U12242 (N_12242,N_11290,N_11563);
xnor U12243 (N_12243,N_11619,N_11528);
or U12244 (N_12244,N_11270,N_11792);
nand U12245 (N_12245,N_11581,N_11392);
or U12246 (N_12246,N_11435,N_11768);
xor U12247 (N_12247,N_11922,N_11663);
and U12248 (N_12248,N_11908,N_11220);
xnor U12249 (N_12249,N_11213,N_11030);
nor U12250 (N_12250,N_11505,N_11966);
nor U12251 (N_12251,N_11450,N_11684);
nor U12252 (N_12252,N_11708,N_11240);
nor U12253 (N_12253,N_11565,N_11309);
and U12254 (N_12254,N_11847,N_11142);
and U12255 (N_12255,N_11094,N_11417);
nor U12256 (N_12256,N_11587,N_11774);
or U12257 (N_12257,N_11829,N_11306);
nor U12258 (N_12258,N_11777,N_11765);
and U12259 (N_12259,N_11919,N_11981);
or U12260 (N_12260,N_11984,N_11297);
nand U12261 (N_12261,N_11414,N_11810);
nand U12262 (N_12262,N_11635,N_11081);
nor U12263 (N_12263,N_11538,N_11611);
and U12264 (N_12264,N_11248,N_11595);
or U12265 (N_12265,N_11698,N_11682);
or U12266 (N_12266,N_11367,N_11656);
or U12267 (N_12267,N_11858,N_11865);
nand U12268 (N_12268,N_11588,N_11797);
nor U12269 (N_12269,N_11195,N_11704);
or U12270 (N_12270,N_11665,N_11341);
xor U12271 (N_12271,N_11983,N_11199);
nand U12272 (N_12272,N_11031,N_11814);
xor U12273 (N_12273,N_11582,N_11408);
nand U12274 (N_12274,N_11659,N_11234);
or U12275 (N_12275,N_11546,N_11003);
nand U12276 (N_12276,N_11933,N_11703);
and U12277 (N_12277,N_11636,N_11807);
xor U12278 (N_12278,N_11018,N_11594);
nand U12279 (N_12279,N_11912,N_11499);
or U12280 (N_12280,N_11960,N_11108);
nor U12281 (N_12281,N_11468,N_11359);
nor U12282 (N_12282,N_11802,N_11562);
nor U12283 (N_12283,N_11183,N_11799);
xnor U12284 (N_12284,N_11888,N_11112);
and U12285 (N_12285,N_11620,N_11474);
and U12286 (N_12286,N_11110,N_11009);
nand U12287 (N_12287,N_11861,N_11186);
xor U12288 (N_12288,N_11019,N_11416);
xor U12289 (N_12289,N_11380,N_11567);
and U12290 (N_12290,N_11393,N_11485);
xor U12291 (N_12291,N_11403,N_11866);
or U12292 (N_12292,N_11280,N_11023);
xor U12293 (N_12293,N_11688,N_11549);
nand U12294 (N_12294,N_11051,N_11104);
xor U12295 (N_12295,N_11957,N_11215);
xor U12296 (N_12296,N_11976,N_11669);
or U12297 (N_12297,N_11828,N_11503);
nand U12298 (N_12298,N_11028,N_11170);
or U12299 (N_12299,N_11812,N_11643);
nor U12300 (N_12300,N_11605,N_11911);
nor U12301 (N_12301,N_11987,N_11017);
nand U12302 (N_12302,N_11864,N_11490);
nor U12303 (N_12303,N_11789,N_11433);
nor U12304 (N_12304,N_11571,N_11355);
nor U12305 (N_12305,N_11098,N_11891);
or U12306 (N_12306,N_11767,N_11877);
xor U12307 (N_12307,N_11120,N_11894);
nor U12308 (N_12308,N_11954,N_11365);
nand U12309 (N_12309,N_11939,N_11266);
nor U12310 (N_12310,N_11576,N_11706);
nand U12311 (N_12311,N_11375,N_11011);
and U12312 (N_12312,N_11951,N_11921);
or U12313 (N_12313,N_11737,N_11645);
nor U12314 (N_12314,N_11564,N_11311);
and U12315 (N_12315,N_11707,N_11580);
nor U12316 (N_12316,N_11506,N_11801);
nor U12317 (N_12317,N_11596,N_11840);
nor U12318 (N_12318,N_11116,N_11261);
or U12319 (N_12319,N_11486,N_11892);
and U12320 (N_12320,N_11222,N_11045);
nand U12321 (N_12321,N_11161,N_11926);
and U12322 (N_12322,N_11321,N_11998);
nor U12323 (N_12323,N_11626,N_11039);
and U12324 (N_12324,N_11551,N_11352);
or U12325 (N_12325,N_11382,N_11250);
or U12326 (N_12326,N_11711,N_11253);
nor U12327 (N_12327,N_11724,N_11185);
nor U12328 (N_12328,N_11683,N_11598);
nand U12329 (N_12329,N_11934,N_11140);
and U12330 (N_12330,N_11869,N_11846);
xor U12331 (N_12331,N_11670,N_11831);
or U12332 (N_12332,N_11178,N_11154);
or U12333 (N_12333,N_11674,N_11407);
or U12334 (N_12334,N_11412,N_11514);
nand U12335 (N_12335,N_11144,N_11138);
and U12336 (N_12336,N_11415,N_11573);
nor U12337 (N_12337,N_11438,N_11242);
nor U12338 (N_12338,N_11459,N_11370);
and U12339 (N_12339,N_11167,N_11504);
nor U12340 (N_12340,N_11766,N_11996);
and U12341 (N_12341,N_11226,N_11617);
xnor U12342 (N_12342,N_11054,N_11052);
and U12343 (N_12343,N_11289,N_11907);
or U12344 (N_12344,N_11277,N_11184);
nand U12345 (N_12345,N_11729,N_11231);
and U12346 (N_12346,N_11191,N_11060);
nand U12347 (N_12347,N_11500,N_11511);
xor U12348 (N_12348,N_11296,N_11305);
nor U12349 (N_12349,N_11950,N_11388);
nor U12350 (N_12350,N_11879,N_11300);
and U12351 (N_12351,N_11444,N_11058);
nand U12352 (N_12352,N_11053,N_11145);
xnor U12353 (N_12353,N_11876,N_11411);
and U12354 (N_12354,N_11361,N_11057);
nor U12355 (N_12355,N_11273,N_11818);
xor U12356 (N_12356,N_11687,N_11946);
and U12357 (N_12357,N_11293,N_11962);
and U12358 (N_12358,N_11165,N_11238);
and U12359 (N_12359,N_11241,N_11422);
nor U12360 (N_12360,N_11041,N_11035);
nor U12361 (N_12361,N_11873,N_11315);
nor U12362 (N_12362,N_11326,N_11431);
nor U12363 (N_12363,N_11350,N_11134);
xnor U12364 (N_12364,N_11258,N_11065);
or U12365 (N_12365,N_11819,N_11395);
nor U12366 (N_12366,N_11093,N_11083);
or U12367 (N_12367,N_11900,N_11432);
xor U12368 (N_12368,N_11714,N_11730);
nand U12369 (N_12369,N_11554,N_11772);
nor U12370 (N_12370,N_11320,N_11029);
nand U12371 (N_12371,N_11221,N_11608);
nor U12372 (N_12372,N_11817,N_11469);
and U12373 (N_12373,N_11808,N_11600);
and U12374 (N_12374,N_11547,N_11622);
and U12375 (N_12375,N_11287,N_11398);
xnor U12376 (N_12376,N_11798,N_11310);
nand U12377 (N_12377,N_11324,N_11292);
or U12378 (N_12378,N_11693,N_11524);
or U12379 (N_12379,N_11637,N_11271);
nor U12380 (N_12380,N_11568,N_11513);
or U12381 (N_12381,N_11491,N_11881);
or U12382 (N_12382,N_11756,N_11179);
xnor U12383 (N_12383,N_11901,N_11425);
xor U12384 (N_12384,N_11360,N_11034);
or U12385 (N_12385,N_11652,N_11989);
xnor U12386 (N_12386,N_11709,N_11750);
or U12387 (N_12387,N_11518,N_11961);
nand U12388 (N_12388,N_11021,N_11237);
xor U12389 (N_12389,N_11331,N_11533);
nand U12390 (N_12390,N_11915,N_11784);
or U12391 (N_12391,N_11536,N_11747);
nand U12392 (N_12392,N_11153,N_11157);
nor U12393 (N_12393,N_11702,N_11495);
nand U12394 (N_12394,N_11454,N_11351);
and U12395 (N_12395,N_11621,N_11800);
nor U12396 (N_12396,N_11307,N_11471);
or U12397 (N_12397,N_11493,N_11625);
xnor U12398 (N_12398,N_11899,N_11940);
nor U12399 (N_12399,N_11958,N_11342);
xnor U12400 (N_12400,N_11779,N_11040);
nand U12401 (N_12401,N_11597,N_11069);
nand U12402 (N_12402,N_11805,N_11225);
nand U12403 (N_12403,N_11368,N_11883);
or U12404 (N_12404,N_11256,N_11206);
nor U12405 (N_12405,N_11870,N_11445);
xnor U12406 (N_12406,N_11868,N_11102);
and U12407 (N_12407,N_11760,N_11423);
and U12408 (N_12408,N_11151,N_11672);
nor U12409 (N_12409,N_11228,N_11358);
nor U12410 (N_12410,N_11988,N_11219);
nor U12411 (N_12411,N_11440,N_11413);
and U12412 (N_12412,N_11344,N_11539);
and U12413 (N_12413,N_11211,N_11123);
or U12414 (N_12414,N_11124,N_11710);
xnor U12415 (N_12415,N_11496,N_11924);
nand U12416 (N_12416,N_11882,N_11133);
xor U12417 (N_12417,N_11666,N_11190);
xnor U12418 (N_12418,N_11811,N_11487);
xor U12419 (N_12419,N_11610,N_11938);
nor U12420 (N_12420,N_11025,N_11660);
nand U12421 (N_12421,N_11498,N_11705);
and U12422 (N_12422,N_11603,N_11259);
and U12423 (N_12423,N_11849,N_11402);
nand U12424 (N_12424,N_11286,N_11667);
nor U12425 (N_12425,N_11136,N_11042);
nor U12426 (N_12426,N_11442,N_11844);
nand U12427 (N_12427,N_11783,N_11970);
nand U12428 (N_12428,N_11148,N_11920);
and U12429 (N_12429,N_11024,N_11997);
xnor U12430 (N_12430,N_11731,N_11757);
nor U12431 (N_12431,N_11640,N_11209);
and U12432 (N_12432,N_11451,N_11319);
nor U12433 (N_12433,N_11356,N_11839);
nand U12434 (N_12434,N_11752,N_11172);
xnor U12435 (N_12435,N_11339,N_11198);
nor U12436 (N_12436,N_11650,N_11788);
nand U12437 (N_12437,N_11794,N_11880);
xnor U12438 (N_12438,N_11176,N_11096);
xnor U12439 (N_12439,N_11115,N_11673);
and U12440 (N_12440,N_11244,N_11992);
nor U12441 (N_12441,N_11048,N_11303);
or U12442 (N_12442,N_11646,N_11947);
xnor U12443 (N_12443,N_11863,N_11227);
and U12444 (N_12444,N_11239,N_11357);
or U12445 (N_12445,N_11279,N_11728);
nand U12446 (N_12446,N_11156,N_11787);
or U12447 (N_12447,N_11235,N_11429);
or U12448 (N_12448,N_11288,N_11131);
and U12449 (N_12449,N_11230,N_11275);
or U12450 (N_12450,N_11532,N_11995);
nand U12451 (N_12451,N_11887,N_11299);
and U12452 (N_12452,N_11012,N_11627);
nand U12453 (N_12453,N_11246,N_11931);
and U12454 (N_12454,N_11544,N_11738);
or U12455 (N_12455,N_11335,N_11556);
nor U12456 (N_12456,N_11540,N_11519);
nor U12457 (N_12457,N_11482,N_11449);
nand U12458 (N_12458,N_11316,N_11200);
nor U12459 (N_12459,N_11362,N_11008);
and U12460 (N_12460,N_11033,N_11971);
or U12461 (N_12461,N_11125,N_11537);
and U12462 (N_12462,N_11875,N_11723);
xnor U12463 (N_12463,N_11642,N_11955);
nand U12464 (N_12464,N_11430,N_11267);
nand U12465 (N_12465,N_11049,N_11405);
or U12466 (N_12466,N_11867,N_11639);
nor U12467 (N_12467,N_11097,N_11127);
nand U12468 (N_12468,N_11174,N_11916);
xor U12469 (N_12469,N_11930,N_11566);
nand U12470 (N_12470,N_11889,N_11751);
and U12471 (N_12471,N_11073,N_11371);
nand U12472 (N_12472,N_11353,N_11999);
or U12473 (N_12473,N_11741,N_11816);
nor U12474 (N_12474,N_11139,N_11340);
or U12475 (N_12475,N_11968,N_11082);
nand U12476 (N_12476,N_11255,N_11002);
xor U12477 (N_12477,N_11143,N_11038);
xor U12478 (N_12478,N_11077,N_11192);
and U12479 (N_12479,N_11634,N_11196);
or U12480 (N_12480,N_11654,N_11690);
or U12481 (N_12481,N_11763,N_11769);
or U12482 (N_12482,N_11833,N_11150);
xnor U12483 (N_12483,N_11100,N_11890);
or U12484 (N_12484,N_11399,N_11322);
or U12485 (N_12485,N_11734,N_11121);
and U12486 (N_12486,N_11182,N_11895);
and U12487 (N_12487,N_11502,N_11489);
or U12488 (N_12488,N_11925,N_11974);
and U12489 (N_12489,N_11776,N_11158);
xnor U12490 (N_12490,N_11484,N_11177);
or U12491 (N_12491,N_11334,N_11526);
or U12492 (N_12492,N_11475,N_11373);
and U12493 (N_12493,N_11128,N_11790);
and U12494 (N_12494,N_11624,N_11072);
or U12495 (N_12495,N_11677,N_11712);
or U12496 (N_12496,N_11436,N_11338);
or U12497 (N_12497,N_11644,N_11283);
and U12498 (N_12498,N_11552,N_11694);
nor U12499 (N_12499,N_11606,N_11612);
nand U12500 (N_12500,N_11335,N_11238);
xor U12501 (N_12501,N_11269,N_11574);
xor U12502 (N_12502,N_11793,N_11012);
nand U12503 (N_12503,N_11449,N_11540);
xor U12504 (N_12504,N_11824,N_11406);
nand U12505 (N_12505,N_11268,N_11696);
or U12506 (N_12506,N_11847,N_11018);
xnor U12507 (N_12507,N_11065,N_11286);
nor U12508 (N_12508,N_11935,N_11162);
xor U12509 (N_12509,N_11224,N_11736);
nor U12510 (N_12510,N_11845,N_11848);
xnor U12511 (N_12511,N_11669,N_11363);
nor U12512 (N_12512,N_11551,N_11298);
nand U12513 (N_12513,N_11505,N_11074);
and U12514 (N_12514,N_11527,N_11759);
xnor U12515 (N_12515,N_11664,N_11205);
xor U12516 (N_12516,N_11252,N_11493);
and U12517 (N_12517,N_11003,N_11941);
nor U12518 (N_12518,N_11095,N_11880);
nand U12519 (N_12519,N_11927,N_11891);
or U12520 (N_12520,N_11635,N_11036);
and U12521 (N_12521,N_11817,N_11316);
xnor U12522 (N_12522,N_11748,N_11799);
nor U12523 (N_12523,N_11442,N_11400);
nand U12524 (N_12524,N_11702,N_11575);
or U12525 (N_12525,N_11304,N_11145);
nand U12526 (N_12526,N_11392,N_11364);
and U12527 (N_12527,N_11682,N_11236);
nor U12528 (N_12528,N_11081,N_11110);
and U12529 (N_12529,N_11277,N_11489);
and U12530 (N_12530,N_11305,N_11298);
xor U12531 (N_12531,N_11763,N_11395);
nor U12532 (N_12532,N_11843,N_11433);
or U12533 (N_12533,N_11202,N_11865);
or U12534 (N_12534,N_11319,N_11763);
and U12535 (N_12535,N_11564,N_11108);
or U12536 (N_12536,N_11566,N_11436);
nor U12537 (N_12537,N_11752,N_11356);
xor U12538 (N_12538,N_11448,N_11895);
nand U12539 (N_12539,N_11275,N_11856);
or U12540 (N_12540,N_11370,N_11388);
xnor U12541 (N_12541,N_11365,N_11448);
or U12542 (N_12542,N_11152,N_11908);
and U12543 (N_12543,N_11422,N_11504);
xnor U12544 (N_12544,N_11546,N_11043);
and U12545 (N_12545,N_11647,N_11931);
or U12546 (N_12546,N_11985,N_11610);
xnor U12547 (N_12547,N_11856,N_11585);
xor U12548 (N_12548,N_11278,N_11335);
and U12549 (N_12549,N_11007,N_11866);
nand U12550 (N_12550,N_11958,N_11465);
and U12551 (N_12551,N_11168,N_11671);
or U12552 (N_12552,N_11213,N_11915);
xnor U12553 (N_12553,N_11767,N_11467);
or U12554 (N_12554,N_11087,N_11519);
xnor U12555 (N_12555,N_11678,N_11527);
and U12556 (N_12556,N_11927,N_11416);
nand U12557 (N_12557,N_11856,N_11938);
nor U12558 (N_12558,N_11766,N_11482);
or U12559 (N_12559,N_11396,N_11946);
xnor U12560 (N_12560,N_11874,N_11724);
nand U12561 (N_12561,N_11946,N_11635);
xor U12562 (N_12562,N_11293,N_11374);
and U12563 (N_12563,N_11206,N_11508);
nor U12564 (N_12564,N_11367,N_11574);
nor U12565 (N_12565,N_11375,N_11135);
nor U12566 (N_12566,N_11771,N_11497);
or U12567 (N_12567,N_11169,N_11801);
xnor U12568 (N_12568,N_11051,N_11639);
nor U12569 (N_12569,N_11509,N_11939);
nor U12570 (N_12570,N_11705,N_11954);
nand U12571 (N_12571,N_11250,N_11360);
nand U12572 (N_12572,N_11056,N_11325);
nand U12573 (N_12573,N_11866,N_11897);
and U12574 (N_12574,N_11936,N_11265);
nand U12575 (N_12575,N_11366,N_11448);
nor U12576 (N_12576,N_11026,N_11239);
nand U12577 (N_12577,N_11822,N_11337);
and U12578 (N_12578,N_11002,N_11992);
nand U12579 (N_12579,N_11933,N_11334);
xnor U12580 (N_12580,N_11382,N_11054);
and U12581 (N_12581,N_11741,N_11119);
nand U12582 (N_12582,N_11008,N_11013);
nand U12583 (N_12583,N_11553,N_11597);
xnor U12584 (N_12584,N_11744,N_11067);
and U12585 (N_12585,N_11614,N_11793);
nand U12586 (N_12586,N_11547,N_11802);
or U12587 (N_12587,N_11194,N_11651);
or U12588 (N_12588,N_11020,N_11557);
xor U12589 (N_12589,N_11294,N_11708);
or U12590 (N_12590,N_11633,N_11736);
and U12591 (N_12591,N_11431,N_11624);
xor U12592 (N_12592,N_11620,N_11383);
or U12593 (N_12593,N_11682,N_11056);
and U12594 (N_12594,N_11207,N_11539);
or U12595 (N_12595,N_11513,N_11791);
and U12596 (N_12596,N_11711,N_11736);
nand U12597 (N_12597,N_11469,N_11951);
xnor U12598 (N_12598,N_11975,N_11178);
xnor U12599 (N_12599,N_11985,N_11665);
nor U12600 (N_12600,N_11457,N_11967);
or U12601 (N_12601,N_11175,N_11072);
nand U12602 (N_12602,N_11172,N_11486);
or U12603 (N_12603,N_11983,N_11514);
and U12604 (N_12604,N_11688,N_11042);
nor U12605 (N_12605,N_11967,N_11381);
and U12606 (N_12606,N_11987,N_11638);
nor U12607 (N_12607,N_11997,N_11497);
nand U12608 (N_12608,N_11261,N_11792);
or U12609 (N_12609,N_11180,N_11328);
nor U12610 (N_12610,N_11011,N_11129);
and U12611 (N_12611,N_11226,N_11718);
and U12612 (N_12612,N_11650,N_11137);
nand U12613 (N_12613,N_11592,N_11882);
nor U12614 (N_12614,N_11913,N_11530);
nor U12615 (N_12615,N_11079,N_11246);
and U12616 (N_12616,N_11458,N_11217);
nand U12617 (N_12617,N_11784,N_11091);
xnor U12618 (N_12618,N_11310,N_11042);
or U12619 (N_12619,N_11564,N_11768);
nor U12620 (N_12620,N_11064,N_11952);
xnor U12621 (N_12621,N_11491,N_11985);
xor U12622 (N_12622,N_11111,N_11535);
xnor U12623 (N_12623,N_11657,N_11236);
nor U12624 (N_12624,N_11364,N_11560);
nand U12625 (N_12625,N_11962,N_11255);
nor U12626 (N_12626,N_11018,N_11933);
or U12627 (N_12627,N_11414,N_11625);
nor U12628 (N_12628,N_11267,N_11287);
nor U12629 (N_12629,N_11804,N_11143);
nand U12630 (N_12630,N_11230,N_11137);
nor U12631 (N_12631,N_11646,N_11834);
or U12632 (N_12632,N_11026,N_11257);
nor U12633 (N_12633,N_11000,N_11845);
or U12634 (N_12634,N_11243,N_11311);
xor U12635 (N_12635,N_11380,N_11365);
xnor U12636 (N_12636,N_11950,N_11375);
and U12637 (N_12637,N_11555,N_11294);
nor U12638 (N_12638,N_11036,N_11991);
or U12639 (N_12639,N_11760,N_11172);
nand U12640 (N_12640,N_11327,N_11506);
xor U12641 (N_12641,N_11382,N_11538);
and U12642 (N_12642,N_11859,N_11568);
nand U12643 (N_12643,N_11061,N_11258);
nand U12644 (N_12644,N_11758,N_11358);
nand U12645 (N_12645,N_11372,N_11143);
or U12646 (N_12646,N_11818,N_11401);
and U12647 (N_12647,N_11871,N_11018);
nor U12648 (N_12648,N_11868,N_11455);
or U12649 (N_12649,N_11626,N_11765);
or U12650 (N_12650,N_11464,N_11033);
nor U12651 (N_12651,N_11884,N_11180);
nand U12652 (N_12652,N_11867,N_11378);
xnor U12653 (N_12653,N_11447,N_11026);
or U12654 (N_12654,N_11711,N_11062);
or U12655 (N_12655,N_11645,N_11326);
and U12656 (N_12656,N_11177,N_11504);
and U12657 (N_12657,N_11079,N_11210);
and U12658 (N_12658,N_11680,N_11216);
or U12659 (N_12659,N_11948,N_11630);
nand U12660 (N_12660,N_11479,N_11622);
and U12661 (N_12661,N_11045,N_11400);
nand U12662 (N_12662,N_11667,N_11679);
or U12663 (N_12663,N_11741,N_11617);
nand U12664 (N_12664,N_11240,N_11522);
nor U12665 (N_12665,N_11902,N_11127);
xnor U12666 (N_12666,N_11183,N_11390);
or U12667 (N_12667,N_11737,N_11959);
nor U12668 (N_12668,N_11781,N_11914);
and U12669 (N_12669,N_11223,N_11435);
or U12670 (N_12670,N_11019,N_11661);
and U12671 (N_12671,N_11882,N_11136);
and U12672 (N_12672,N_11539,N_11013);
nor U12673 (N_12673,N_11245,N_11782);
or U12674 (N_12674,N_11924,N_11747);
or U12675 (N_12675,N_11379,N_11273);
nor U12676 (N_12676,N_11779,N_11369);
and U12677 (N_12677,N_11247,N_11406);
or U12678 (N_12678,N_11368,N_11129);
and U12679 (N_12679,N_11785,N_11890);
nor U12680 (N_12680,N_11006,N_11231);
xnor U12681 (N_12681,N_11250,N_11570);
nand U12682 (N_12682,N_11352,N_11805);
or U12683 (N_12683,N_11504,N_11238);
or U12684 (N_12684,N_11228,N_11445);
xnor U12685 (N_12685,N_11447,N_11110);
xor U12686 (N_12686,N_11487,N_11386);
and U12687 (N_12687,N_11234,N_11501);
nor U12688 (N_12688,N_11414,N_11529);
nor U12689 (N_12689,N_11958,N_11679);
xor U12690 (N_12690,N_11162,N_11408);
nand U12691 (N_12691,N_11506,N_11770);
nor U12692 (N_12692,N_11741,N_11079);
and U12693 (N_12693,N_11614,N_11602);
nand U12694 (N_12694,N_11547,N_11935);
nor U12695 (N_12695,N_11667,N_11959);
or U12696 (N_12696,N_11803,N_11362);
and U12697 (N_12697,N_11470,N_11026);
or U12698 (N_12698,N_11287,N_11260);
and U12699 (N_12699,N_11079,N_11721);
nor U12700 (N_12700,N_11979,N_11019);
nand U12701 (N_12701,N_11612,N_11624);
and U12702 (N_12702,N_11733,N_11822);
xor U12703 (N_12703,N_11419,N_11926);
or U12704 (N_12704,N_11865,N_11724);
or U12705 (N_12705,N_11268,N_11143);
nand U12706 (N_12706,N_11988,N_11463);
and U12707 (N_12707,N_11524,N_11828);
xor U12708 (N_12708,N_11739,N_11774);
or U12709 (N_12709,N_11538,N_11549);
nor U12710 (N_12710,N_11780,N_11102);
or U12711 (N_12711,N_11252,N_11877);
xnor U12712 (N_12712,N_11548,N_11244);
or U12713 (N_12713,N_11681,N_11026);
xnor U12714 (N_12714,N_11911,N_11264);
xnor U12715 (N_12715,N_11165,N_11872);
xnor U12716 (N_12716,N_11969,N_11377);
xnor U12717 (N_12717,N_11901,N_11482);
xnor U12718 (N_12718,N_11943,N_11736);
and U12719 (N_12719,N_11236,N_11922);
xor U12720 (N_12720,N_11521,N_11227);
and U12721 (N_12721,N_11902,N_11697);
nand U12722 (N_12722,N_11999,N_11649);
nand U12723 (N_12723,N_11904,N_11212);
xor U12724 (N_12724,N_11250,N_11747);
nand U12725 (N_12725,N_11171,N_11443);
or U12726 (N_12726,N_11719,N_11034);
and U12727 (N_12727,N_11823,N_11841);
xnor U12728 (N_12728,N_11349,N_11101);
or U12729 (N_12729,N_11825,N_11278);
nor U12730 (N_12730,N_11203,N_11826);
nand U12731 (N_12731,N_11210,N_11111);
nand U12732 (N_12732,N_11064,N_11698);
or U12733 (N_12733,N_11862,N_11201);
nor U12734 (N_12734,N_11906,N_11145);
nor U12735 (N_12735,N_11701,N_11681);
and U12736 (N_12736,N_11994,N_11404);
xor U12737 (N_12737,N_11666,N_11761);
nor U12738 (N_12738,N_11763,N_11627);
and U12739 (N_12739,N_11163,N_11795);
xor U12740 (N_12740,N_11279,N_11379);
xor U12741 (N_12741,N_11314,N_11076);
xnor U12742 (N_12742,N_11970,N_11887);
nand U12743 (N_12743,N_11808,N_11217);
or U12744 (N_12744,N_11481,N_11833);
nor U12745 (N_12745,N_11486,N_11130);
nor U12746 (N_12746,N_11658,N_11352);
xor U12747 (N_12747,N_11520,N_11820);
or U12748 (N_12748,N_11987,N_11320);
nand U12749 (N_12749,N_11621,N_11864);
nor U12750 (N_12750,N_11928,N_11831);
xnor U12751 (N_12751,N_11584,N_11401);
or U12752 (N_12752,N_11048,N_11820);
nand U12753 (N_12753,N_11999,N_11675);
xnor U12754 (N_12754,N_11421,N_11166);
or U12755 (N_12755,N_11147,N_11162);
or U12756 (N_12756,N_11018,N_11129);
xnor U12757 (N_12757,N_11457,N_11444);
and U12758 (N_12758,N_11367,N_11290);
nand U12759 (N_12759,N_11253,N_11602);
nor U12760 (N_12760,N_11102,N_11715);
nor U12761 (N_12761,N_11273,N_11816);
xor U12762 (N_12762,N_11057,N_11639);
nor U12763 (N_12763,N_11697,N_11696);
and U12764 (N_12764,N_11303,N_11564);
and U12765 (N_12765,N_11256,N_11985);
or U12766 (N_12766,N_11070,N_11326);
and U12767 (N_12767,N_11081,N_11305);
or U12768 (N_12768,N_11578,N_11673);
or U12769 (N_12769,N_11744,N_11778);
xor U12770 (N_12770,N_11241,N_11627);
or U12771 (N_12771,N_11475,N_11633);
or U12772 (N_12772,N_11907,N_11243);
or U12773 (N_12773,N_11711,N_11356);
or U12774 (N_12774,N_11177,N_11077);
or U12775 (N_12775,N_11895,N_11775);
xnor U12776 (N_12776,N_11374,N_11913);
nand U12777 (N_12777,N_11127,N_11546);
nand U12778 (N_12778,N_11334,N_11755);
and U12779 (N_12779,N_11187,N_11849);
xor U12780 (N_12780,N_11234,N_11908);
and U12781 (N_12781,N_11995,N_11813);
and U12782 (N_12782,N_11561,N_11450);
and U12783 (N_12783,N_11011,N_11948);
nor U12784 (N_12784,N_11896,N_11412);
and U12785 (N_12785,N_11869,N_11463);
and U12786 (N_12786,N_11658,N_11589);
or U12787 (N_12787,N_11811,N_11481);
and U12788 (N_12788,N_11387,N_11487);
nor U12789 (N_12789,N_11609,N_11381);
and U12790 (N_12790,N_11277,N_11764);
xnor U12791 (N_12791,N_11236,N_11824);
nand U12792 (N_12792,N_11053,N_11499);
and U12793 (N_12793,N_11683,N_11678);
xor U12794 (N_12794,N_11436,N_11660);
xor U12795 (N_12795,N_11193,N_11226);
xnor U12796 (N_12796,N_11297,N_11959);
or U12797 (N_12797,N_11268,N_11580);
nor U12798 (N_12798,N_11635,N_11017);
and U12799 (N_12799,N_11099,N_11263);
and U12800 (N_12800,N_11627,N_11229);
or U12801 (N_12801,N_11665,N_11697);
nor U12802 (N_12802,N_11325,N_11033);
or U12803 (N_12803,N_11137,N_11298);
and U12804 (N_12804,N_11823,N_11872);
and U12805 (N_12805,N_11454,N_11202);
xor U12806 (N_12806,N_11607,N_11716);
xor U12807 (N_12807,N_11386,N_11018);
xnor U12808 (N_12808,N_11931,N_11157);
nand U12809 (N_12809,N_11434,N_11054);
nand U12810 (N_12810,N_11443,N_11675);
nand U12811 (N_12811,N_11943,N_11458);
xor U12812 (N_12812,N_11457,N_11689);
nand U12813 (N_12813,N_11272,N_11083);
xnor U12814 (N_12814,N_11717,N_11863);
and U12815 (N_12815,N_11411,N_11221);
or U12816 (N_12816,N_11463,N_11850);
nor U12817 (N_12817,N_11738,N_11083);
nand U12818 (N_12818,N_11543,N_11666);
or U12819 (N_12819,N_11355,N_11795);
nand U12820 (N_12820,N_11865,N_11824);
xnor U12821 (N_12821,N_11675,N_11484);
xor U12822 (N_12822,N_11208,N_11288);
xnor U12823 (N_12823,N_11982,N_11564);
nor U12824 (N_12824,N_11392,N_11913);
xnor U12825 (N_12825,N_11715,N_11421);
xnor U12826 (N_12826,N_11964,N_11317);
xor U12827 (N_12827,N_11929,N_11231);
and U12828 (N_12828,N_11476,N_11569);
xor U12829 (N_12829,N_11462,N_11265);
or U12830 (N_12830,N_11251,N_11035);
nor U12831 (N_12831,N_11304,N_11762);
or U12832 (N_12832,N_11767,N_11248);
and U12833 (N_12833,N_11149,N_11360);
nor U12834 (N_12834,N_11213,N_11782);
and U12835 (N_12835,N_11867,N_11908);
or U12836 (N_12836,N_11583,N_11940);
nor U12837 (N_12837,N_11712,N_11364);
nor U12838 (N_12838,N_11280,N_11514);
and U12839 (N_12839,N_11795,N_11892);
nand U12840 (N_12840,N_11831,N_11832);
and U12841 (N_12841,N_11546,N_11614);
nor U12842 (N_12842,N_11672,N_11045);
nand U12843 (N_12843,N_11922,N_11696);
and U12844 (N_12844,N_11359,N_11442);
or U12845 (N_12845,N_11798,N_11260);
nand U12846 (N_12846,N_11423,N_11345);
nand U12847 (N_12847,N_11460,N_11987);
nand U12848 (N_12848,N_11938,N_11984);
xnor U12849 (N_12849,N_11640,N_11024);
or U12850 (N_12850,N_11861,N_11364);
nand U12851 (N_12851,N_11040,N_11848);
and U12852 (N_12852,N_11644,N_11849);
nor U12853 (N_12853,N_11236,N_11087);
or U12854 (N_12854,N_11916,N_11122);
or U12855 (N_12855,N_11783,N_11875);
nor U12856 (N_12856,N_11024,N_11378);
and U12857 (N_12857,N_11178,N_11397);
xnor U12858 (N_12858,N_11267,N_11199);
nor U12859 (N_12859,N_11299,N_11715);
and U12860 (N_12860,N_11380,N_11416);
and U12861 (N_12861,N_11358,N_11248);
xor U12862 (N_12862,N_11382,N_11536);
nor U12863 (N_12863,N_11514,N_11576);
xor U12864 (N_12864,N_11028,N_11648);
and U12865 (N_12865,N_11083,N_11516);
xor U12866 (N_12866,N_11625,N_11801);
and U12867 (N_12867,N_11040,N_11555);
nor U12868 (N_12868,N_11376,N_11341);
or U12869 (N_12869,N_11272,N_11275);
or U12870 (N_12870,N_11724,N_11659);
xnor U12871 (N_12871,N_11614,N_11376);
and U12872 (N_12872,N_11131,N_11304);
xnor U12873 (N_12873,N_11753,N_11344);
and U12874 (N_12874,N_11843,N_11373);
nor U12875 (N_12875,N_11306,N_11251);
xor U12876 (N_12876,N_11755,N_11492);
nor U12877 (N_12877,N_11989,N_11719);
nand U12878 (N_12878,N_11341,N_11732);
or U12879 (N_12879,N_11768,N_11618);
and U12880 (N_12880,N_11174,N_11342);
nand U12881 (N_12881,N_11678,N_11192);
xor U12882 (N_12882,N_11478,N_11120);
and U12883 (N_12883,N_11097,N_11542);
or U12884 (N_12884,N_11439,N_11382);
nand U12885 (N_12885,N_11099,N_11347);
xnor U12886 (N_12886,N_11219,N_11850);
and U12887 (N_12887,N_11322,N_11943);
nand U12888 (N_12888,N_11913,N_11160);
or U12889 (N_12889,N_11898,N_11535);
xor U12890 (N_12890,N_11683,N_11010);
nor U12891 (N_12891,N_11664,N_11581);
xnor U12892 (N_12892,N_11641,N_11672);
nand U12893 (N_12893,N_11483,N_11831);
and U12894 (N_12894,N_11145,N_11590);
xnor U12895 (N_12895,N_11812,N_11702);
nand U12896 (N_12896,N_11647,N_11477);
xor U12897 (N_12897,N_11230,N_11884);
nand U12898 (N_12898,N_11773,N_11354);
xor U12899 (N_12899,N_11333,N_11091);
xnor U12900 (N_12900,N_11619,N_11577);
nand U12901 (N_12901,N_11987,N_11857);
and U12902 (N_12902,N_11952,N_11010);
nor U12903 (N_12903,N_11802,N_11529);
or U12904 (N_12904,N_11466,N_11751);
or U12905 (N_12905,N_11005,N_11925);
xnor U12906 (N_12906,N_11540,N_11538);
or U12907 (N_12907,N_11237,N_11521);
xor U12908 (N_12908,N_11928,N_11575);
nor U12909 (N_12909,N_11631,N_11784);
and U12910 (N_12910,N_11322,N_11842);
nand U12911 (N_12911,N_11573,N_11563);
and U12912 (N_12912,N_11639,N_11238);
nand U12913 (N_12913,N_11856,N_11894);
or U12914 (N_12914,N_11211,N_11935);
and U12915 (N_12915,N_11973,N_11227);
xnor U12916 (N_12916,N_11607,N_11621);
xor U12917 (N_12917,N_11795,N_11174);
or U12918 (N_12918,N_11968,N_11431);
xnor U12919 (N_12919,N_11650,N_11328);
nand U12920 (N_12920,N_11986,N_11526);
nand U12921 (N_12921,N_11953,N_11104);
nor U12922 (N_12922,N_11148,N_11176);
nor U12923 (N_12923,N_11884,N_11812);
and U12924 (N_12924,N_11624,N_11820);
nand U12925 (N_12925,N_11791,N_11149);
nor U12926 (N_12926,N_11230,N_11219);
and U12927 (N_12927,N_11462,N_11057);
or U12928 (N_12928,N_11862,N_11317);
xor U12929 (N_12929,N_11588,N_11379);
and U12930 (N_12930,N_11058,N_11600);
nor U12931 (N_12931,N_11018,N_11575);
xor U12932 (N_12932,N_11705,N_11119);
or U12933 (N_12933,N_11550,N_11320);
nand U12934 (N_12934,N_11096,N_11908);
nand U12935 (N_12935,N_11336,N_11129);
or U12936 (N_12936,N_11793,N_11942);
xor U12937 (N_12937,N_11344,N_11435);
xor U12938 (N_12938,N_11107,N_11694);
and U12939 (N_12939,N_11040,N_11292);
or U12940 (N_12940,N_11692,N_11009);
nand U12941 (N_12941,N_11347,N_11452);
xor U12942 (N_12942,N_11035,N_11535);
nor U12943 (N_12943,N_11836,N_11189);
or U12944 (N_12944,N_11680,N_11138);
xor U12945 (N_12945,N_11475,N_11160);
nand U12946 (N_12946,N_11426,N_11535);
nor U12947 (N_12947,N_11588,N_11989);
or U12948 (N_12948,N_11830,N_11128);
xor U12949 (N_12949,N_11878,N_11659);
xor U12950 (N_12950,N_11925,N_11825);
and U12951 (N_12951,N_11593,N_11976);
nor U12952 (N_12952,N_11098,N_11128);
xor U12953 (N_12953,N_11900,N_11753);
or U12954 (N_12954,N_11678,N_11769);
nor U12955 (N_12955,N_11592,N_11327);
nand U12956 (N_12956,N_11511,N_11815);
xor U12957 (N_12957,N_11081,N_11976);
nand U12958 (N_12958,N_11556,N_11884);
and U12959 (N_12959,N_11780,N_11728);
and U12960 (N_12960,N_11842,N_11348);
xnor U12961 (N_12961,N_11220,N_11098);
and U12962 (N_12962,N_11222,N_11385);
nand U12963 (N_12963,N_11222,N_11204);
or U12964 (N_12964,N_11811,N_11137);
and U12965 (N_12965,N_11935,N_11306);
nand U12966 (N_12966,N_11641,N_11515);
xnor U12967 (N_12967,N_11023,N_11828);
nand U12968 (N_12968,N_11677,N_11929);
xor U12969 (N_12969,N_11416,N_11297);
or U12970 (N_12970,N_11620,N_11531);
or U12971 (N_12971,N_11503,N_11653);
xor U12972 (N_12972,N_11107,N_11515);
and U12973 (N_12973,N_11126,N_11555);
xnor U12974 (N_12974,N_11629,N_11817);
and U12975 (N_12975,N_11653,N_11933);
and U12976 (N_12976,N_11457,N_11199);
xor U12977 (N_12977,N_11919,N_11943);
or U12978 (N_12978,N_11640,N_11406);
and U12979 (N_12979,N_11216,N_11713);
nor U12980 (N_12980,N_11371,N_11993);
nor U12981 (N_12981,N_11948,N_11109);
or U12982 (N_12982,N_11062,N_11813);
xor U12983 (N_12983,N_11800,N_11017);
or U12984 (N_12984,N_11252,N_11737);
and U12985 (N_12985,N_11575,N_11633);
xnor U12986 (N_12986,N_11190,N_11623);
and U12987 (N_12987,N_11993,N_11282);
or U12988 (N_12988,N_11162,N_11785);
and U12989 (N_12989,N_11757,N_11890);
nor U12990 (N_12990,N_11792,N_11374);
xnor U12991 (N_12991,N_11329,N_11785);
or U12992 (N_12992,N_11538,N_11428);
or U12993 (N_12993,N_11379,N_11865);
nor U12994 (N_12994,N_11156,N_11453);
nor U12995 (N_12995,N_11276,N_11381);
nand U12996 (N_12996,N_11203,N_11822);
and U12997 (N_12997,N_11037,N_11179);
nand U12998 (N_12998,N_11307,N_11503);
and U12999 (N_12999,N_11356,N_11080);
xnor U13000 (N_13000,N_12666,N_12253);
and U13001 (N_13001,N_12409,N_12298);
nand U13002 (N_13002,N_12630,N_12206);
nand U13003 (N_13003,N_12896,N_12668);
or U13004 (N_13004,N_12034,N_12921);
nand U13005 (N_13005,N_12315,N_12820);
and U13006 (N_13006,N_12613,N_12130);
nor U13007 (N_13007,N_12371,N_12712);
nor U13008 (N_13008,N_12767,N_12801);
nand U13009 (N_13009,N_12335,N_12098);
and U13010 (N_13010,N_12734,N_12363);
and U13011 (N_13011,N_12405,N_12947);
nand U13012 (N_13012,N_12512,N_12148);
or U13013 (N_13013,N_12653,N_12854);
or U13014 (N_13014,N_12431,N_12636);
nor U13015 (N_13015,N_12380,N_12511);
nand U13016 (N_13016,N_12264,N_12863);
or U13017 (N_13017,N_12418,N_12879);
nor U13018 (N_13018,N_12463,N_12458);
nor U13019 (N_13019,N_12196,N_12460);
or U13020 (N_13020,N_12743,N_12012);
and U13021 (N_13021,N_12741,N_12086);
nand U13022 (N_13022,N_12422,N_12145);
or U13023 (N_13023,N_12607,N_12089);
nand U13024 (N_13024,N_12269,N_12758);
xor U13025 (N_13025,N_12878,N_12679);
nand U13026 (N_13026,N_12830,N_12410);
and U13027 (N_13027,N_12326,N_12153);
xor U13028 (N_13028,N_12141,N_12402);
nand U13029 (N_13029,N_12891,N_12680);
nand U13030 (N_13030,N_12053,N_12260);
or U13031 (N_13031,N_12194,N_12969);
and U13032 (N_13032,N_12276,N_12800);
nor U13033 (N_13033,N_12869,N_12008);
nor U13034 (N_13034,N_12439,N_12814);
nor U13035 (N_13035,N_12441,N_12728);
or U13036 (N_13036,N_12336,N_12781);
nor U13037 (N_13037,N_12654,N_12585);
xnor U13038 (N_13038,N_12088,N_12268);
nor U13039 (N_13039,N_12274,N_12270);
or U13040 (N_13040,N_12513,N_12765);
and U13041 (N_13041,N_12818,N_12306);
xnor U13042 (N_13042,N_12462,N_12442);
nor U13043 (N_13043,N_12261,N_12573);
nand U13044 (N_13044,N_12722,N_12533);
xor U13045 (N_13045,N_12045,N_12877);
nor U13046 (N_13046,N_12964,N_12074);
nor U13047 (N_13047,N_12783,N_12397);
nor U13048 (N_13048,N_12273,N_12614);
or U13049 (N_13049,N_12282,N_12903);
nand U13050 (N_13050,N_12381,N_12184);
nand U13051 (N_13051,N_12127,N_12251);
nor U13052 (N_13052,N_12024,N_12707);
xnor U13053 (N_13053,N_12425,N_12938);
nor U13054 (N_13054,N_12929,N_12774);
xnor U13055 (N_13055,N_12207,N_12976);
xnor U13056 (N_13056,N_12019,N_12702);
xnor U13057 (N_13057,N_12242,N_12255);
or U13058 (N_13058,N_12448,N_12889);
nor U13059 (N_13059,N_12182,N_12404);
nor U13060 (N_13060,N_12093,N_12732);
or U13061 (N_13061,N_12189,N_12091);
xnor U13062 (N_13062,N_12939,N_12620);
nand U13063 (N_13063,N_12514,N_12050);
xnor U13064 (N_13064,N_12882,N_12014);
or U13065 (N_13065,N_12487,N_12786);
nand U13066 (N_13066,N_12884,N_12279);
and U13067 (N_13067,N_12539,N_12049);
xor U13068 (N_13068,N_12331,N_12694);
xnor U13069 (N_13069,N_12673,N_12945);
or U13070 (N_13070,N_12561,N_12224);
xor U13071 (N_13071,N_12423,N_12684);
nand U13072 (N_13072,N_12575,N_12633);
xor U13073 (N_13073,N_12243,N_12726);
xnor U13074 (N_13074,N_12919,N_12044);
xnor U13075 (N_13075,N_12432,N_12411);
or U13076 (N_13076,N_12280,N_12337);
nand U13077 (N_13077,N_12526,N_12004);
xor U13078 (N_13078,N_12187,N_12105);
nor U13079 (N_13079,N_12011,N_12435);
xnor U13080 (N_13080,N_12565,N_12340);
xnor U13081 (N_13081,N_12623,N_12547);
or U13082 (N_13082,N_12698,N_12374);
nor U13083 (N_13083,N_12087,N_12924);
or U13084 (N_13084,N_12991,N_12813);
or U13085 (N_13085,N_12061,N_12406);
nor U13086 (N_13086,N_12385,N_12659);
nand U13087 (N_13087,N_12731,N_12876);
or U13088 (N_13088,N_12793,N_12847);
xor U13089 (N_13089,N_12020,N_12824);
nor U13090 (N_13090,N_12318,N_12930);
nor U13091 (N_13091,N_12199,N_12389);
or U13092 (N_13092,N_12447,N_12332);
and U13093 (N_13093,N_12475,N_12853);
xnor U13094 (N_13094,N_12424,N_12366);
and U13095 (N_13095,N_12073,N_12150);
nand U13096 (N_13096,N_12103,N_12700);
nand U13097 (N_13097,N_12809,N_12957);
or U13098 (N_13098,N_12713,N_12277);
nand U13099 (N_13099,N_12505,N_12845);
xnor U13100 (N_13100,N_12772,N_12911);
nor U13101 (N_13101,N_12035,N_12655);
xor U13102 (N_13102,N_12022,N_12506);
and U13103 (N_13103,N_12382,N_12092);
xor U13104 (N_13104,N_12197,N_12499);
nand U13105 (N_13105,N_12346,N_12616);
xnor U13106 (N_13106,N_12691,N_12085);
and U13107 (N_13107,N_12443,N_12535);
and U13108 (N_13108,N_12980,N_12163);
and U13109 (N_13109,N_12844,N_12619);
nand U13110 (N_13110,N_12730,N_12683);
nor U13111 (N_13111,N_12392,N_12135);
nor U13112 (N_13112,N_12601,N_12874);
nand U13113 (N_13113,N_12245,N_12909);
and U13114 (N_13114,N_12586,N_12241);
nor U13115 (N_13115,N_12151,N_12168);
xnor U13116 (N_13116,N_12681,N_12204);
xnor U13117 (N_13117,N_12622,N_12927);
and U13118 (N_13118,N_12605,N_12572);
xor U13119 (N_13119,N_12489,N_12912);
xnor U13120 (N_13120,N_12519,N_12894);
nand U13121 (N_13121,N_12795,N_12946);
xnor U13122 (N_13122,N_12500,N_12275);
xnor U13123 (N_13123,N_12288,N_12704);
nand U13124 (N_13124,N_12674,N_12333);
and U13125 (N_13125,N_12648,N_12828);
nand U13126 (N_13126,N_12379,N_12716);
or U13127 (N_13127,N_12583,N_12940);
nor U13128 (N_13128,N_12450,N_12110);
or U13129 (N_13129,N_12477,N_12757);
or U13130 (N_13130,N_12117,N_12481);
or U13131 (N_13131,N_12016,N_12313);
nor U13132 (N_13132,N_12030,N_12624);
xnor U13133 (N_13133,N_12688,N_12143);
and U13134 (N_13134,N_12358,N_12023);
nand U13135 (N_13135,N_12100,N_12183);
or U13136 (N_13136,N_12949,N_12522);
and U13137 (N_13137,N_12762,N_12827);
nor U13138 (N_13138,N_12436,N_12651);
or U13139 (N_13139,N_12888,N_12075);
and U13140 (N_13140,N_12538,N_12835);
nand U13141 (N_13141,N_12562,N_12094);
and U13142 (N_13142,N_12026,N_12661);
nor U13143 (N_13143,N_12871,N_12552);
or U13144 (N_13144,N_12308,N_12796);
nand U13145 (N_13145,N_12761,N_12071);
and U13146 (N_13146,N_12805,N_12490);
and U13147 (N_13147,N_12574,N_12042);
or U13148 (N_13148,N_12584,N_12753);
and U13149 (N_13149,N_12373,N_12319);
and U13150 (N_13150,N_12887,N_12198);
nor U13151 (N_13151,N_12192,N_12311);
xor U13152 (N_13152,N_12995,N_12589);
nor U13153 (N_13153,N_12330,N_12480);
or U13154 (N_13154,N_12498,N_12556);
nand U13155 (N_13155,N_12587,N_12367);
nor U13156 (N_13156,N_12900,N_12735);
nor U13157 (N_13157,N_12915,N_12532);
and U13158 (N_13158,N_12777,N_12027);
and U13159 (N_13159,N_12039,N_12545);
xor U13160 (N_13160,N_12858,N_12440);
and U13161 (N_13161,N_12317,N_12898);
and U13162 (N_13162,N_12842,N_12375);
nor U13163 (N_13163,N_12802,N_12662);
or U13164 (N_13164,N_12862,N_12948);
nor U13165 (N_13165,N_12213,N_12908);
nand U13166 (N_13166,N_12467,N_12686);
or U13167 (N_13167,N_12338,N_12438);
nand U13168 (N_13168,N_12567,N_12256);
nor U13169 (N_13169,N_12803,N_12396);
or U13170 (N_13170,N_12483,N_12115);
or U13171 (N_13171,N_12162,N_12119);
nand U13172 (N_13172,N_12365,N_12598);
nor U13173 (N_13173,N_12631,N_12059);
nand U13174 (N_13174,N_12357,N_12983);
nand U13175 (N_13175,N_12880,N_12300);
xnor U13176 (N_13176,N_12111,N_12857);
nand U13177 (N_13177,N_12920,N_12928);
nand U13178 (N_13178,N_12839,N_12452);
or U13179 (N_13179,N_12142,N_12356);
nand U13180 (N_13180,N_12953,N_12961);
nand U13181 (N_13181,N_12473,N_12872);
xnor U13182 (N_13182,N_12109,N_12246);
nand U13183 (N_13183,N_12797,N_12923);
or U13184 (N_13184,N_12459,N_12064);
nand U13185 (N_13185,N_12750,N_12247);
or U13186 (N_13186,N_12017,N_12540);
nor U13187 (N_13187,N_12848,N_12348);
xnor U13188 (N_13188,N_12811,N_12551);
or U13189 (N_13189,N_12591,N_12124);
xnor U13190 (N_13190,N_12203,N_12951);
nor U13191 (N_13191,N_12868,N_12593);
xnor U13192 (N_13192,N_12350,N_12295);
and U13193 (N_13193,N_12342,N_12705);
nor U13194 (N_13194,N_12324,N_12541);
xor U13195 (N_13195,N_12553,N_12998);
or U13196 (N_13196,N_12901,N_12077);
or U13197 (N_13197,N_12977,N_12979);
nor U13198 (N_13198,N_12696,N_12852);
nor U13199 (N_13199,N_12208,N_12592);
or U13200 (N_13200,N_12334,N_12474);
xnor U13201 (N_13201,N_12046,N_12984);
and U13202 (N_13202,N_12353,N_12417);
or U13203 (N_13203,N_12286,N_12377);
and U13204 (N_13204,N_12082,N_12076);
nand U13205 (N_13205,N_12225,N_12727);
or U13206 (N_13206,N_12174,N_12725);
nand U13207 (N_13207,N_12149,N_12158);
nand U13208 (N_13208,N_12263,N_12861);
nand U13209 (N_13209,N_12955,N_12383);
or U13210 (N_13210,N_12209,N_12554);
nand U13211 (N_13211,N_12217,N_12544);
nor U13212 (N_13212,N_12733,N_12769);
or U13213 (N_13213,N_12952,N_12740);
nand U13214 (N_13214,N_12906,N_12904);
xor U13215 (N_13215,N_12658,N_12237);
nor U13216 (N_13216,N_12576,N_12465);
and U13217 (N_13217,N_12936,N_12766);
nor U13218 (N_13218,N_12195,N_12159);
nand U13219 (N_13219,N_12122,N_12695);
nand U13220 (N_13220,N_12052,N_12309);
xnor U13221 (N_13221,N_12492,N_12006);
xnor U13222 (N_13222,N_12644,N_12515);
and U13223 (N_13223,N_12671,N_12285);
xor U13224 (N_13224,N_12981,N_12025);
and U13225 (N_13225,N_12007,N_12388);
nand U13226 (N_13226,N_12621,N_12628);
or U13227 (N_13227,N_12883,N_12287);
or U13228 (N_13228,N_12643,N_12962);
nand U13229 (N_13229,N_12387,N_12864);
xnor U13230 (N_13230,N_12033,N_12775);
and U13231 (N_13231,N_12294,N_12354);
nand U13232 (N_13232,N_12170,N_12232);
nand U13233 (N_13233,N_12823,N_12067);
or U13234 (N_13234,N_12164,N_12079);
and U13235 (N_13235,N_12746,N_12994);
nand U13236 (N_13236,N_12993,N_12663);
xor U13237 (N_13237,N_12488,N_12254);
and U13238 (N_13238,N_12495,N_12136);
xor U13239 (N_13239,N_12084,N_12875);
or U13240 (N_13240,N_12560,N_12770);
and U13241 (N_13241,N_12973,N_12051);
or U13242 (N_13242,N_12491,N_12013);
nor U13243 (N_13243,N_12118,N_12239);
or U13244 (N_13244,N_12714,N_12699);
nand U13245 (N_13245,N_12937,N_12219);
xor U13246 (N_13246,N_12637,N_12398);
nor U13247 (N_13247,N_12469,N_12099);
nand U13248 (N_13248,N_12860,N_12126);
xnor U13249 (N_13249,N_12468,N_12031);
nor U13250 (N_13250,N_12910,N_12461);
or U13251 (N_13251,N_12407,N_12559);
or U13252 (N_13252,N_12555,N_12886);
xnor U13253 (N_13253,N_12185,N_12116);
or U13254 (N_13254,N_12010,N_12779);
or U13255 (N_13255,N_12617,N_12221);
xnor U13256 (N_13256,N_12133,N_12597);
nor U13257 (N_13257,N_12101,N_12790);
and U13258 (N_13258,N_12036,N_12018);
nor U13259 (N_13259,N_12866,N_12784);
nand U13260 (N_13260,N_12521,N_12687);
xnor U13261 (N_13261,N_12179,N_12152);
or U13262 (N_13262,N_12466,N_12629);
xor U13263 (N_13263,N_12055,N_12132);
nand U13264 (N_13264,N_12240,N_12789);
and U13265 (N_13265,N_12451,N_12646);
or U13266 (N_13266,N_12171,N_12855);
nor U13267 (N_13267,N_12478,N_12359);
or U13268 (N_13268,N_12181,N_12129);
and U13269 (N_13269,N_12453,N_12138);
nor U13270 (N_13270,N_12250,N_12314);
xor U13271 (N_13271,N_12502,N_12302);
nand U13272 (N_13272,N_12167,N_12230);
nand U13273 (N_13273,N_12278,N_12248);
and U13274 (N_13274,N_12697,N_12665);
nor U13275 (N_13275,N_12083,N_12914);
xor U13276 (N_13276,N_12283,N_12768);
nor U13277 (N_13277,N_12773,N_12916);
or U13278 (N_13278,N_12721,N_12566);
nor U13279 (N_13279,N_12625,N_12815);
and U13280 (N_13280,N_12220,N_12744);
and U13281 (N_13281,N_12627,N_12634);
and U13282 (N_13282,N_12485,N_12216);
and U13283 (N_13283,N_12941,N_12106);
or U13284 (N_13284,N_12120,N_12798);
or U13285 (N_13285,N_12710,N_12907);
xnor U13286 (N_13286,N_12021,N_12497);
xnor U13287 (N_13287,N_12229,N_12228);
or U13288 (N_13288,N_12390,N_12484);
and U13289 (N_13289,N_12708,N_12832);
nor U13290 (N_13290,N_12403,N_12751);
xor U13291 (N_13291,N_12218,N_12144);
nand U13292 (N_13292,N_12426,N_12943);
and U13293 (N_13293,N_12657,N_12368);
xnor U13294 (N_13294,N_12062,N_12542);
nand U13295 (N_13295,N_12266,N_12987);
and U13296 (N_13296,N_12530,N_12345);
or U13297 (N_13297,N_12291,N_12549);
nor U13298 (N_13298,N_12156,N_12177);
xnor U13299 (N_13299,N_12428,N_12180);
xnor U13300 (N_13300,N_12518,N_12455);
and U13301 (N_13301,N_12808,N_12227);
or U13302 (N_13302,N_12233,N_12434);
or U13303 (N_13303,N_12290,N_12978);
nand U13304 (N_13304,N_12186,N_12244);
or U13305 (N_13305,N_12437,N_12967);
and U13306 (N_13306,N_12899,N_12343);
xor U13307 (N_13307,N_12711,N_12057);
and U13308 (N_13308,N_12486,N_12926);
nor U13309 (N_13309,N_12078,N_12040);
nand U13310 (N_13310,N_12931,N_12446);
and U13311 (N_13311,N_12009,N_12265);
xor U13312 (N_13312,N_12370,N_12416);
nand U13313 (N_13313,N_12905,N_12701);
or U13314 (N_13314,N_12344,N_12493);
or U13315 (N_13315,N_12176,N_12529);
nand U13316 (N_13316,N_12304,N_12558);
nand U13317 (N_13317,N_12165,N_12670);
xnor U13318 (N_13318,N_12037,N_12272);
nor U13319 (N_13319,N_12161,N_12822);
or U13320 (N_13320,N_12960,N_12408);
or U13321 (N_13321,N_12231,N_12550);
nor U13322 (N_13322,N_12043,N_12667);
and U13323 (N_13323,N_12054,N_12913);
nor U13324 (N_13324,N_12881,N_12582);
or U13325 (N_13325,N_12546,N_12996);
nor U13326 (N_13326,N_12525,N_12739);
and U13327 (N_13327,N_12341,N_12096);
nor U13328 (N_13328,N_12072,N_12131);
xor U13329 (N_13329,N_12234,N_12785);
nor U13330 (N_13330,N_12169,N_12956);
or U13331 (N_13331,N_12709,N_12193);
and U13332 (N_13332,N_12807,N_12137);
and U13333 (N_13333,N_12850,N_12672);
nor U13334 (N_13334,N_12301,N_12361);
and U13335 (N_13335,N_12415,N_12048);
xor U13336 (N_13336,N_12258,N_12412);
xor U13337 (N_13337,N_12201,N_12959);
nand U13338 (N_13338,N_12639,N_12003);
xnor U13339 (N_13339,N_12420,N_12190);
nand U13340 (N_13340,N_12327,N_12376);
and U13341 (N_13341,N_12147,N_12501);
nor U13342 (N_13342,N_12950,N_12972);
xnor U13343 (N_13343,N_12935,N_12594);
or U13344 (N_13344,N_12840,N_12577);
or U13345 (N_13345,N_12843,N_12482);
or U13346 (N_13346,N_12305,N_12178);
or U13347 (N_13347,N_12384,N_12588);
and U13348 (N_13348,N_12296,N_12760);
nor U13349 (N_13349,N_12610,N_12215);
nand U13350 (N_13350,N_12323,N_12873);
nor U13351 (N_13351,N_12347,N_12222);
and U13352 (N_13352,N_12838,N_12271);
nor U13353 (N_13353,N_12214,N_12974);
or U13354 (N_13354,N_12738,N_12609);
and U13355 (N_13355,N_12211,N_12826);
nand U13356 (N_13356,N_12472,N_12108);
or U13357 (N_13357,N_12471,N_12596);
nor U13358 (N_13358,N_12351,N_12917);
or U13359 (N_13359,N_12836,N_12259);
nor U13360 (N_13360,N_12649,N_12524);
xnor U13361 (N_13361,N_12401,N_12504);
nand U13362 (N_13362,N_12509,N_12479);
and U13363 (N_13363,N_12812,N_12395);
or U13364 (N_13364,N_12157,N_12780);
xor U13365 (N_13365,N_12339,N_12191);
xor U13366 (N_13366,N_12029,N_12693);
nor U13367 (N_13367,N_12128,N_12413);
or U13368 (N_13368,N_12841,N_12692);
xnor U13369 (N_13369,N_12971,N_12364);
or U13370 (N_13370,N_12837,N_12536);
and U13371 (N_13371,N_12641,N_12429);
or U13372 (N_13372,N_12252,N_12355);
or U13373 (N_13373,N_12281,N_12669);
and U13374 (N_13374,N_12989,N_12717);
xor U13375 (N_13375,N_12457,N_12284);
xnor U13376 (N_13376,N_12508,N_12675);
xnor U13377 (N_13377,N_12070,N_12548);
nor U13378 (N_13378,N_12001,N_12262);
or U13379 (N_13379,N_12867,N_12104);
or U13380 (N_13380,N_12819,N_12564);
or U13381 (N_13381,N_12745,N_12997);
xnor U13382 (N_13382,N_12325,N_12982);
nand U13383 (N_13383,N_12985,N_12421);
nor U13384 (N_13384,N_12494,N_12792);
xnor U13385 (N_13385,N_12000,N_12267);
or U13386 (N_13386,N_12257,N_12752);
xor U13387 (N_13387,N_12321,N_12534);
nand U13388 (N_13388,N_12865,N_12897);
xor U13389 (N_13389,N_12788,N_12656);
nor U13390 (N_13390,N_12032,N_12932);
nor U13391 (N_13391,N_12747,N_12297);
nor U13392 (N_13392,N_12729,N_12706);
xnor U13393 (N_13393,N_12097,N_12427);
and U13394 (N_13394,N_12754,N_12322);
and U13395 (N_13395,N_12102,N_12372);
nand U13396 (N_13396,N_12581,N_12470);
nand U13397 (N_13397,N_12015,N_12703);
and U13398 (N_13398,N_12080,N_12892);
nand U13399 (N_13399,N_12527,N_12954);
xnor U13400 (N_13400,N_12238,N_12557);
or U13401 (N_13401,N_12890,N_12794);
and U13402 (N_13402,N_12604,N_12058);
xor U13403 (N_13403,N_12507,N_12289);
xnor U13404 (N_13404,N_12816,N_12378);
or U13405 (N_13405,N_12090,N_12893);
and U13406 (N_13406,N_12293,N_12825);
xor U13407 (N_13407,N_12362,N_12329);
and U13408 (N_13408,N_12642,N_12715);
or U13409 (N_13409,N_12352,N_12925);
xor U13410 (N_13410,N_12066,N_12678);
nor U13411 (N_13411,N_12172,N_12791);
nor U13412 (N_13412,N_12677,N_12310);
and U13413 (N_13413,N_12303,N_12724);
xnor U13414 (N_13414,N_12782,N_12123);
or U13415 (N_13415,N_12134,N_12571);
or U13416 (N_13416,N_12810,N_12933);
nor U13417 (N_13417,N_12517,N_12114);
nand U13418 (N_13418,N_12113,N_12682);
or U13419 (N_13419,N_12771,N_12069);
nand U13420 (N_13420,N_12520,N_12849);
nand U13421 (N_13421,N_12543,N_12503);
nor U13422 (N_13422,N_12223,N_12175);
nand U13423 (N_13423,N_12394,N_12060);
or U13424 (N_13424,N_12449,N_12831);
or U13425 (N_13425,N_12320,N_12047);
nor U13426 (N_13426,N_12249,N_12676);
and U13427 (N_13427,N_12859,N_12817);
nor U13428 (N_13428,N_12764,N_12778);
xnor U13429 (N_13429,N_12121,N_12205);
nor U13430 (N_13430,N_12200,N_12834);
and U13431 (N_13431,N_12107,N_12360);
and U13432 (N_13432,N_12599,N_12737);
and U13433 (N_13433,N_12723,N_12063);
or U13434 (N_13434,N_12393,N_12292);
xnor U13435 (N_13435,N_12081,N_12755);
and U13436 (N_13436,N_12433,N_12068);
xnor U13437 (N_13437,N_12464,N_12608);
and U13438 (N_13438,N_12125,N_12414);
nand U13439 (N_13439,N_12603,N_12400);
nor U13440 (N_13440,N_12719,N_12895);
or U13441 (N_13441,N_12650,N_12002);
or U13442 (N_13442,N_12166,N_12690);
or U13443 (N_13443,N_12992,N_12602);
or U13444 (N_13444,N_12988,N_12885);
nand U13445 (N_13445,N_12570,N_12618);
xnor U13446 (N_13446,N_12160,N_12568);
nand U13447 (N_13447,N_12445,N_12612);
nor U13448 (N_13448,N_12173,N_12226);
xnor U13449 (N_13449,N_12038,N_12188);
or U13450 (N_13450,N_12776,N_12647);
nand U13451 (N_13451,N_12578,N_12510);
and U13452 (N_13452,N_12563,N_12399);
or U13453 (N_13453,N_12028,N_12833);
and U13454 (N_13454,N_12312,N_12328);
nand U13455 (N_13455,N_12922,N_12146);
nand U13456 (N_13456,N_12632,N_12645);
nor U13457 (N_13457,N_12870,N_12299);
nand U13458 (N_13458,N_12748,N_12419);
or U13459 (N_13459,N_12689,N_12369);
xor U13460 (N_13460,N_12391,N_12851);
nand U13461 (N_13461,N_12531,N_12155);
and U13462 (N_13462,N_12056,N_12759);
and U13463 (N_13463,N_12965,N_12804);
and U13464 (N_13464,N_12806,N_12970);
and U13465 (N_13465,N_12718,N_12999);
and U13466 (N_13466,N_12918,N_12430);
nand U13467 (N_13467,N_12615,N_12756);
and U13468 (N_13468,N_12944,N_12966);
nand U13469 (N_13469,N_12685,N_12990);
or U13470 (N_13470,N_12986,N_12537);
or U13471 (N_13471,N_12902,N_12821);
nand U13472 (N_13472,N_12580,N_12742);
nor U13473 (N_13473,N_12664,N_12112);
and U13474 (N_13474,N_12934,N_12476);
or U13475 (N_13475,N_12005,N_12942);
xor U13476 (N_13476,N_12963,N_12523);
nand U13477 (N_13477,N_12958,N_12202);
xnor U13478 (N_13478,N_12846,N_12606);
or U13479 (N_13479,N_12095,N_12626);
and U13480 (N_13480,N_12611,N_12856);
and U13481 (N_13481,N_12579,N_12635);
nand U13482 (N_13482,N_12139,N_12496);
or U13483 (N_13483,N_12787,N_12154);
nor U13484 (N_13484,N_12652,N_12975);
nand U13485 (N_13485,N_12516,N_12799);
nand U13486 (N_13486,N_12968,N_12307);
xor U13487 (N_13487,N_12316,N_12528);
or U13488 (N_13488,N_12600,N_12736);
and U13489 (N_13489,N_12386,N_12454);
xnor U13490 (N_13490,N_12212,N_12660);
and U13491 (N_13491,N_12210,N_12720);
xnor U13492 (N_13492,N_12829,N_12236);
or U13493 (N_13493,N_12349,N_12065);
and U13494 (N_13494,N_12763,N_12590);
and U13495 (N_13495,N_12569,N_12640);
nand U13496 (N_13496,N_12595,N_12456);
nor U13497 (N_13497,N_12638,N_12140);
xor U13498 (N_13498,N_12235,N_12444);
and U13499 (N_13499,N_12041,N_12749);
and U13500 (N_13500,N_12199,N_12594);
xor U13501 (N_13501,N_12951,N_12150);
xor U13502 (N_13502,N_12330,N_12656);
nand U13503 (N_13503,N_12100,N_12624);
xnor U13504 (N_13504,N_12029,N_12347);
xor U13505 (N_13505,N_12814,N_12753);
or U13506 (N_13506,N_12204,N_12457);
nor U13507 (N_13507,N_12048,N_12849);
xor U13508 (N_13508,N_12411,N_12274);
nand U13509 (N_13509,N_12844,N_12446);
nor U13510 (N_13510,N_12321,N_12429);
nor U13511 (N_13511,N_12061,N_12792);
nand U13512 (N_13512,N_12971,N_12451);
and U13513 (N_13513,N_12950,N_12590);
or U13514 (N_13514,N_12735,N_12248);
nand U13515 (N_13515,N_12845,N_12673);
nand U13516 (N_13516,N_12071,N_12927);
or U13517 (N_13517,N_12759,N_12027);
nor U13518 (N_13518,N_12806,N_12928);
nand U13519 (N_13519,N_12375,N_12970);
nor U13520 (N_13520,N_12391,N_12491);
nor U13521 (N_13521,N_12709,N_12499);
or U13522 (N_13522,N_12858,N_12295);
or U13523 (N_13523,N_12140,N_12461);
or U13524 (N_13524,N_12465,N_12615);
xor U13525 (N_13525,N_12439,N_12001);
and U13526 (N_13526,N_12436,N_12342);
nand U13527 (N_13527,N_12955,N_12919);
nand U13528 (N_13528,N_12169,N_12801);
nand U13529 (N_13529,N_12617,N_12190);
xor U13530 (N_13530,N_12640,N_12979);
and U13531 (N_13531,N_12420,N_12526);
nand U13532 (N_13532,N_12675,N_12800);
and U13533 (N_13533,N_12882,N_12917);
nor U13534 (N_13534,N_12079,N_12300);
and U13535 (N_13535,N_12010,N_12194);
or U13536 (N_13536,N_12129,N_12169);
xor U13537 (N_13537,N_12773,N_12570);
and U13538 (N_13538,N_12883,N_12125);
nand U13539 (N_13539,N_12390,N_12618);
nor U13540 (N_13540,N_12988,N_12435);
and U13541 (N_13541,N_12180,N_12945);
nand U13542 (N_13542,N_12534,N_12994);
nor U13543 (N_13543,N_12013,N_12159);
or U13544 (N_13544,N_12009,N_12196);
and U13545 (N_13545,N_12660,N_12658);
nor U13546 (N_13546,N_12116,N_12640);
nor U13547 (N_13547,N_12481,N_12631);
nor U13548 (N_13548,N_12209,N_12806);
and U13549 (N_13549,N_12772,N_12483);
and U13550 (N_13550,N_12913,N_12257);
nor U13551 (N_13551,N_12468,N_12854);
xnor U13552 (N_13552,N_12543,N_12662);
nor U13553 (N_13553,N_12089,N_12605);
or U13554 (N_13554,N_12167,N_12664);
and U13555 (N_13555,N_12654,N_12510);
nor U13556 (N_13556,N_12454,N_12790);
or U13557 (N_13557,N_12601,N_12115);
nor U13558 (N_13558,N_12815,N_12480);
or U13559 (N_13559,N_12846,N_12015);
nor U13560 (N_13560,N_12282,N_12751);
and U13561 (N_13561,N_12020,N_12533);
nand U13562 (N_13562,N_12120,N_12227);
and U13563 (N_13563,N_12115,N_12487);
or U13564 (N_13564,N_12991,N_12014);
and U13565 (N_13565,N_12173,N_12627);
nor U13566 (N_13566,N_12786,N_12676);
nand U13567 (N_13567,N_12196,N_12289);
xor U13568 (N_13568,N_12237,N_12536);
or U13569 (N_13569,N_12273,N_12524);
nand U13570 (N_13570,N_12723,N_12091);
xnor U13571 (N_13571,N_12629,N_12194);
or U13572 (N_13572,N_12754,N_12829);
nor U13573 (N_13573,N_12941,N_12276);
or U13574 (N_13574,N_12965,N_12679);
xnor U13575 (N_13575,N_12836,N_12494);
nor U13576 (N_13576,N_12857,N_12759);
and U13577 (N_13577,N_12770,N_12789);
nand U13578 (N_13578,N_12678,N_12203);
nor U13579 (N_13579,N_12400,N_12525);
or U13580 (N_13580,N_12581,N_12830);
and U13581 (N_13581,N_12811,N_12979);
nor U13582 (N_13582,N_12480,N_12257);
nand U13583 (N_13583,N_12502,N_12344);
or U13584 (N_13584,N_12926,N_12814);
xnor U13585 (N_13585,N_12304,N_12901);
xnor U13586 (N_13586,N_12020,N_12469);
nor U13587 (N_13587,N_12889,N_12751);
or U13588 (N_13588,N_12264,N_12038);
xor U13589 (N_13589,N_12140,N_12363);
nand U13590 (N_13590,N_12651,N_12393);
and U13591 (N_13591,N_12289,N_12629);
nand U13592 (N_13592,N_12438,N_12250);
or U13593 (N_13593,N_12031,N_12289);
nand U13594 (N_13594,N_12432,N_12302);
xor U13595 (N_13595,N_12457,N_12987);
xor U13596 (N_13596,N_12256,N_12999);
or U13597 (N_13597,N_12377,N_12078);
or U13598 (N_13598,N_12081,N_12877);
and U13599 (N_13599,N_12006,N_12708);
nand U13600 (N_13600,N_12206,N_12785);
nor U13601 (N_13601,N_12344,N_12066);
nand U13602 (N_13602,N_12238,N_12023);
nand U13603 (N_13603,N_12085,N_12546);
or U13604 (N_13604,N_12664,N_12121);
nor U13605 (N_13605,N_12843,N_12370);
xnor U13606 (N_13606,N_12954,N_12714);
xnor U13607 (N_13607,N_12910,N_12798);
xor U13608 (N_13608,N_12758,N_12747);
and U13609 (N_13609,N_12041,N_12150);
nor U13610 (N_13610,N_12761,N_12105);
xor U13611 (N_13611,N_12267,N_12792);
nand U13612 (N_13612,N_12472,N_12771);
nand U13613 (N_13613,N_12317,N_12158);
and U13614 (N_13614,N_12692,N_12906);
xor U13615 (N_13615,N_12740,N_12311);
nor U13616 (N_13616,N_12780,N_12132);
or U13617 (N_13617,N_12117,N_12261);
and U13618 (N_13618,N_12892,N_12765);
and U13619 (N_13619,N_12266,N_12260);
xnor U13620 (N_13620,N_12755,N_12896);
and U13621 (N_13621,N_12469,N_12450);
and U13622 (N_13622,N_12003,N_12344);
xor U13623 (N_13623,N_12842,N_12143);
and U13624 (N_13624,N_12973,N_12467);
and U13625 (N_13625,N_12661,N_12616);
nor U13626 (N_13626,N_12221,N_12514);
nand U13627 (N_13627,N_12550,N_12431);
and U13628 (N_13628,N_12315,N_12190);
nand U13629 (N_13629,N_12767,N_12038);
and U13630 (N_13630,N_12325,N_12682);
nand U13631 (N_13631,N_12724,N_12258);
and U13632 (N_13632,N_12421,N_12333);
nand U13633 (N_13633,N_12162,N_12100);
nor U13634 (N_13634,N_12289,N_12135);
and U13635 (N_13635,N_12697,N_12293);
or U13636 (N_13636,N_12934,N_12173);
nor U13637 (N_13637,N_12541,N_12576);
nor U13638 (N_13638,N_12209,N_12856);
nand U13639 (N_13639,N_12254,N_12640);
or U13640 (N_13640,N_12248,N_12942);
and U13641 (N_13641,N_12227,N_12637);
nand U13642 (N_13642,N_12569,N_12247);
or U13643 (N_13643,N_12904,N_12179);
xor U13644 (N_13644,N_12407,N_12202);
xor U13645 (N_13645,N_12815,N_12367);
and U13646 (N_13646,N_12442,N_12895);
nand U13647 (N_13647,N_12291,N_12568);
and U13648 (N_13648,N_12926,N_12608);
xnor U13649 (N_13649,N_12670,N_12696);
xnor U13650 (N_13650,N_12205,N_12134);
xnor U13651 (N_13651,N_12196,N_12710);
xor U13652 (N_13652,N_12746,N_12073);
or U13653 (N_13653,N_12473,N_12754);
nor U13654 (N_13654,N_12600,N_12997);
and U13655 (N_13655,N_12173,N_12736);
and U13656 (N_13656,N_12806,N_12666);
or U13657 (N_13657,N_12903,N_12305);
nor U13658 (N_13658,N_12421,N_12332);
or U13659 (N_13659,N_12497,N_12009);
or U13660 (N_13660,N_12868,N_12104);
and U13661 (N_13661,N_12817,N_12684);
and U13662 (N_13662,N_12257,N_12262);
xnor U13663 (N_13663,N_12925,N_12904);
or U13664 (N_13664,N_12402,N_12521);
xnor U13665 (N_13665,N_12819,N_12726);
or U13666 (N_13666,N_12405,N_12195);
nor U13667 (N_13667,N_12753,N_12785);
nand U13668 (N_13668,N_12407,N_12996);
nand U13669 (N_13669,N_12642,N_12760);
nand U13670 (N_13670,N_12149,N_12957);
nor U13671 (N_13671,N_12695,N_12762);
and U13672 (N_13672,N_12192,N_12486);
and U13673 (N_13673,N_12199,N_12146);
xor U13674 (N_13674,N_12569,N_12567);
nand U13675 (N_13675,N_12450,N_12250);
xnor U13676 (N_13676,N_12424,N_12568);
or U13677 (N_13677,N_12913,N_12270);
and U13678 (N_13678,N_12875,N_12800);
nor U13679 (N_13679,N_12557,N_12045);
or U13680 (N_13680,N_12474,N_12073);
or U13681 (N_13681,N_12001,N_12011);
and U13682 (N_13682,N_12014,N_12046);
nor U13683 (N_13683,N_12225,N_12541);
or U13684 (N_13684,N_12440,N_12618);
or U13685 (N_13685,N_12479,N_12854);
and U13686 (N_13686,N_12343,N_12361);
xnor U13687 (N_13687,N_12666,N_12547);
nor U13688 (N_13688,N_12128,N_12755);
and U13689 (N_13689,N_12291,N_12674);
and U13690 (N_13690,N_12962,N_12405);
or U13691 (N_13691,N_12401,N_12306);
xor U13692 (N_13692,N_12339,N_12941);
xnor U13693 (N_13693,N_12945,N_12938);
nand U13694 (N_13694,N_12559,N_12080);
or U13695 (N_13695,N_12822,N_12766);
xor U13696 (N_13696,N_12563,N_12199);
xnor U13697 (N_13697,N_12222,N_12525);
or U13698 (N_13698,N_12864,N_12220);
nand U13699 (N_13699,N_12433,N_12604);
or U13700 (N_13700,N_12752,N_12657);
nor U13701 (N_13701,N_12226,N_12731);
and U13702 (N_13702,N_12350,N_12110);
and U13703 (N_13703,N_12999,N_12022);
nand U13704 (N_13704,N_12566,N_12638);
and U13705 (N_13705,N_12238,N_12921);
and U13706 (N_13706,N_12418,N_12586);
and U13707 (N_13707,N_12896,N_12740);
or U13708 (N_13708,N_12326,N_12785);
and U13709 (N_13709,N_12216,N_12651);
nor U13710 (N_13710,N_12416,N_12018);
or U13711 (N_13711,N_12806,N_12938);
nand U13712 (N_13712,N_12486,N_12373);
nand U13713 (N_13713,N_12130,N_12761);
nand U13714 (N_13714,N_12509,N_12863);
nor U13715 (N_13715,N_12698,N_12715);
nor U13716 (N_13716,N_12934,N_12500);
nand U13717 (N_13717,N_12482,N_12593);
and U13718 (N_13718,N_12303,N_12131);
nand U13719 (N_13719,N_12772,N_12344);
nand U13720 (N_13720,N_12747,N_12613);
and U13721 (N_13721,N_12171,N_12688);
or U13722 (N_13722,N_12417,N_12917);
and U13723 (N_13723,N_12603,N_12781);
or U13724 (N_13724,N_12869,N_12726);
nand U13725 (N_13725,N_12464,N_12336);
nor U13726 (N_13726,N_12548,N_12487);
nand U13727 (N_13727,N_12004,N_12275);
nor U13728 (N_13728,N_12462,N_12845);
xor U13729 (N_13729,N_12465,N_12717);
nor U13730 (N_13730,N_12056,N_12211);
nor U13731 (N_13731,N_12808,N_12903);
xor U13732 (N_13732,N_12654,N_12847);
or U13733 (N_13733,N_12798,N_12079);
or U13734 (N_13734,N_12476,N_12421);
and U13735 (N_13735,N_12662,N_12329);
nor U13736 (N_13736,N_12444,N_12425);
nand U13737 (N_13737,N_12244,N_12694);
and U13738 (N_13738,N_12147,N_12244);
or U13739 (N_13739,N_12995,N_12325);
xnor U13740 (N_13740,N_12251,N_12528);
nand U13741 (N_13741,N_12555,N_12584);
xor U13742 (N_13742,N_12753,N_12036);
and U13743 (N_13743,N_12997,N_12022);
or U13744 (N_13744,N_12582,N_12437);
or U13745 (N_13745,N_12492,N_12294);
xor U13746 (N_13746,N_12278,N_12679);
nor U13747 (N_13747,N_12775,N_12039);
nand U13748 (N_13748,N_12860,N_12601);
nor U13749 (N_13749,N_12139,N_12135);
xnor U13750 (N_13750,N_12812,N_12940);
and U13751 (N_13751,N_12017,N_12067);
xnor U13752 (N_13752,N_12161,N_12071);
xnor U13753 (N_13753,N_12117,N_12015);
and U13754 (N_13754,N_12752,N_12061);
nand U13755 (N_13755,N_12716,N_12609);
or U13756 (N_13756,N_12880,N_12353);
and U13757 (N_13757,N_12575,N_12296);
and U13758 (N_13758,N_12473,N_12155);
nand U13759 (N_13759,N_12537,N_12677);
nand U13760 (N_13760,N_12920,N_12222);
xor U13761 (N_13761,N_12549,N_12476);
nor U13762 (N_13762,N_12871,N_12777);
xnor U13763 (N_13763,N_12102,N_12064);
nor U13764 (N_13764,N_12733,N_12310);
nand U13765 (N_13765,N_12150,N_12871);
and U13766 (N_13766,N_12072,N_12508);
nand U13767 (N_13767,N_12614,N_12933);
nor U13768 (N_13768,N_12965,N_12375);
and U13769 (N_13769,N_12375,N_12610);
nor U13770 (N_13770,N_12662,N_12205);
nand U13771 (N_13771,N_12495,N_12655);
and U13772 (N_13772,N_12469,N_12758);
or U13773 (N_13773,N_12960,N_12804);
nor U13774 (N_13774,N_12996,N_12911);
xor U13775 (N_13775,N_12562,N_12398);
nor U13776 (N_13776,N_12880,N_12121);
xor U13777 (N_13777,N_12374,N_12459);
nor U13778 (N_13778,N_12746,N_12144);
or U13779 (N_13779,N_12181,N_12228);
nor U13780 (N_13780,N_12119,N_12301);
xor U13781 (N_13781,N_12632,N_12876);
nor U13782 (N_13782,N_12419,N_12131);
and U13783 (N_13783,N_12561,N_12896);
nor U13784 (N_13784,N_12404,N_12841);
xor U13785 (N_13785,N_12179,N_12166);
nand U13786 (N_13786,N_12935,N_12390);
xnor U13787 (N_13787,N_12923,N_12855);
or U13788 (N_13788,N_12435,N_12935);
or U13789 (N_13789,N_12059,N_12376);
nand U13790 (N_13790,N_12614,N_12574);
and U13791 (N_13791,N_12573,N_12592);
xnor U13792 (N_13792,N_12685,N_12616);
and U13793 (N_13793,N_12677,N_12416);
nand U13794 (N_13794,N_12206,N_12751);
nand U13795 (N_13795,N_12705,N_12350);
xor U13796 (N_13796,N_12229,N_12182);
or U13797 (N_13797,N_12299,N_12173);
xnor U13798 (N_13798,N_12067,N_12846);
xnor U13799 (N_13799,N_12386,N_12671);
nand U13800 (N_13800,N_12791,N_12779);
nor U13801 (N_13801,N_12018,N_12207);
nand U13802 (N_13802,N_12261,N_12536);
nor U13803 (N_13803,N_12213,N_12080);
and U13804 (N_13804,N_12112,N_12282);
and U13805 (N_13805,N_12515,N_12512);
or U13806 (N_13806,N_12644,N_12940);
xor U13807 (N_13807,N_12267,N_12761);
nand U13808 (N_13808,N_12757,N_12986);
nand U13809 (N_13809,N_12421,N_12779);
nand U13810 (N_13810,N_12373,N_12776);
xnor U13811 (N_13811,N_12831,N_12415);
nor U13812 (N_13812,N_12069,N_12994);
nand U13813 (N_13813,N_12180,N_12327);
and U13814 (N_13814,N_12219,N_12406);
nor U13815 (N_13815,N_12273,N_12605);
nor U13816 (N_13816,N_12788,N_12793);
nor U13817 (N_13817,N_12052,N_12034);
nor U13818 (N_13818,N_12993,N_12776);
nand U13819 (N_13819,N_12847,N_12668);
and U13820 (N_13820,N_12395,N_12290);
or U13821 (N_13821,N_12562,N_12908);
nand U13822 (N_13822,N_12907,N_12100);
or U13823 (N_13823,N_12710,N_12439);
nor U13824 (N_13824,N_12389,N_12912);
xnor U13825 (N_13825,N_12836,N_12179);
xnor U13826 (N_13826,N_12010,N_12253);
or U13827 (N_13827,N_12999,N_12869);
and U13828 (N_13828,N_12019,N_12798);
nand U13829 (N_13829,N_12380,N_12538);
nor U13830 (N_13830,N_12199,N_12251);
nand U13831 (N_13831,N_12553,N_12340);
xnor U13832 (N_13832,N_12542,N_12808);
and U13833 (N_13833,N_12556,N_12362);
and U13834 (N_13834,N_12262,N_12943);
and U13835 (N_13835,N_12279,N_12145);
nand U13836 (N_13836,N_12286,N_12285);
and U13837 (N_13837,N_12953,N_12280);
or U13838 (N_13838,N_12729,N_12383);
xor U13839 (N_13839,N_12805,N_12150);
nand U13840 (N_13840,N_12562,N_12414);
nor U13841 (N_13841,N_12139,N_12495);
nor U13842 (N_13842,N_12239,N_12587);
nand U13843 (N_13843,N_12177,N_12049);
xnor U13844 (N_13844,N_12217,N_12252);
xor U13845 (N_13845,N_12081,N_12808);
and U13846 (N_13846,N_12144,N_12455);
and U13847 (N_13847,N_12714,N_12509);
nor U13848 (N_13848,N_12522,N_12008);
and U13849 (N_13849,N_12273,N_12745);
and U13850 (N_13850,N_12082,N_12166);
and U13851 (N_13851,N_12389,N_12384);
nand U13852 (N_13852,N_12167,N_12520);
xnor U13853 (N_13853,N_12409,N_12583);
nor U13854 (N_13854,N_12079,N_12086);
or U13855 (N_13855,N_12311,N_12993);
and U13856 (N_13856,N_12642,N_12538);
xnor U13857 (N_13857,N_12552,N_12050);
and U13858 (N_13858,N_12954,N_12268);
or U13859 (N_13859,N_12082,N_12384);
nand U13860 (N_13860,N_12003,N_12931);
or U13861 (N_13861,N_12581,N_12481);
nor U13862 (N_13862,N_12205,N_12708);
nand U13863 (N_13863,N_12939,N_12565);
xor U13864 (N_13864,N_12698,N_12471);
nand U13865 (N_13865,N_12017,N_12259);
nand U13866 (N_13866,N_12095,N_12340);
nand U13867 (N_13867,N_12759,N_12350);
nand U13868 (N_13868,N_12948,N_12034);
and U13869 (N_13869,N_12020,N_12953);
or U13870 (N_13870,N_12518,N_12220);
nor U13871 (N_13871,N_12319,N_12416);
nor U13872 (N_13872,N_12858,N_12016);
xor U13873 (N_13873,N_12851,N_12184);
or U13874 (N_13874,N_12243,N_12935);
nor U13875 (N_13875,N_12656,N_12687);
or U13876 (N_13876,N_12775,N_12958);
nand U13877 (N_13877,N_12349,N_12072);
and U13878 (N_13878,N_12965,N_12584);
nor U13879 (N_13879,N_12299,N_12655);
or U13880 (N_13880,N_12709,N_12991);
nand U13881 (N_13881,N_12384,N_12995);
xnor U13882 (N_13882,N_12496,N_12797);
and U13883 (N_13883,N_12578,N_12269);
or U13884 (N_13884,N_12239,N_12443);
xor U13885 (N_13885,N_12525,N_12461);
nor U13886 (N_13886,N_12478,N_12527);
nand U13887 (N_13887,N_12233,N_12829);
or U13888 (N_13888,N_12979,N_12231);
nand U13889 (N_13889,N_12414,N_12485);
nand U13890 (N_13890,N_12391,N_12600);
and U13891 (N_13891,N_12932,N_12514);
or U13892 (N_13892,N_12264,N_12201);
nor U13893 (N_13893,N_12967,N_12599);
and U13894 (N_13894,N_12051,N_12913);
nor U13895 (N_13895,N_12711,N_12811);
nand U13896 (N_13896,N_12987,N_12130);
nor U13897 (N_13897,N_12425,N_12103);
nand U13898 (N_13898,N_12131,N_12329);
xor U13899 (N_13899,N_12699,N_12760);
and U13900 (N_13900,N_12521,N_12029);
or U13901 (N_13901,N_12768,N_12267);
and U13902 (N_13902,N_12367,N_12305);
nand U13903 (N_13903,N_12554,N_12832);
nand U13904 (N_13904,N_12941,N_12440);
nor U13905 (N_13905,N_12983,N_12852);
nor U13906 (N_13906,N_12832,N_12349);
nor U13907 (N_13907,N_12594,N_12785);
nor U13908 (N_13908,N_12534,N_12256);
and U13909 (N_13909,N_12869,N_12815);
xor U13910 (N_13910,N_12634,N_12819);
xor U13911 (N_13911,N_12284,N_12817);
and U13912 (N_13912,N_12855,N_12030);
xnor U13913 (N_13913,N_12732,N_12898);
and U13914 (N_13914,N_12227,N_12837);
or U13915 (N_13915,N_12319,N_12642);
or U13916 (N_13916,N_12601,N_12513);
nand U13917 (N_13917,N_12538,N_12065);
nor U13918 (N_13918,N_12422,N_12165);
and U13919 (N_13919,N_12126,N_12899);
nand U13920 (N_13920,N_12459,N_12104);
and U13921 (N_13921,N_12719,N_12372);
nand U13922 (N_13922,N_12666,N_12187);
nand U13923 (N_13923,N_12553,N_12500);
nor U13924 (N_13924,N_12605,N_12760);
nor U13925 (N_13925,N_12715,N_12079);
xnor U13926 (N_13926,N_12659,N_12870);
nor U13927 (N_13927,N_12156,N_12908);
nor U13928 (N_13928,N_12725,N_12675);
xor U13929 (N_13929,N_12710,N_12289);
xor U13930 (N_13930,N_12207,N_12569);
and U13931 (N_13931,N_12326,N_12770);
xnor U13932 (N_13932,N_12650,N_12043);
nand U13933 (N_13933,N_12314,N_12319);
xor U13934 (N_13934,N_12123,N_12651);
xnor U13935 (N_13935,N_12180,N_12504);
and U13936 (N_13936,N_12925,N_12236);
nor U13937 (N_13937,N_12937,N_12295);
and U13938 (N_13938,N_12915,N_12334);
nor U13939 (N_13939,N_12984,N_12989);
nand U13940 (N_13940,N_12939,N_12539);
xnor U13941 (N_13941,N_12209,N_12492);
or U13942 (N_13942,N_12797,N_12104);
nand U13943 (N_13943,N_12504,N_12646);
or U13944 (N_13944,N_12673,N_12583);
or U13945 (N_13945,N_12949,N_12801);
xnor U13946 (N_13946,N_12431,N_12985);
xnor U13947 (N_13947,N_12262,N_12648);
xor U13948 (N_13948,N_12125,N_12010);
xor U13949 (N_13949,N_12002,N_12458);
or U13950 (N_13950,N_12760,N_12728);
and U13951 (N_13951,N_12268,N_12017);
nor U13952 (N_13952,N_12045,N_12979);
nor U13953 (N_13953,N_12423,N_12765);
xor U13954 (N_13954,N_12195,N_12704);
or U13955 (N_13955,N_12666,N_12532);
and U13956 (N_13956,N_12838,N_12127);
and U13957 (N_13957,N_12939,N_12644);
nand U13958 (N_13958,N_12434,N_12155);
nor U13959 (N_13959,N_12538,N_12029);
nand U13960 (N_13960,N_12439,N_12905);
or U13961 (N_13961,N_12809,N_12303);
or U13962 (N_13962,N_12882,N_12814);
or U13963 (N_13963,N_12651,N_12323);
nand U13964 (N_13964,N_12443,N_12595);
and U13965 (N_13965,N_12179,N_12312);
or U13966 (N_13966,N_12561,N_12860);
or U13967 (N_13967,N_12774,N_12338);
nor U13968 (N_13968,N_12209,N_12883);
or U13969 (N_13969,N_12670,N_12277);
xnor U13970 (N_13970,N_12637,N_12221);
nand U13971 (N_13971,N_12607,N_12192);
nor U13972 (N_13972,N_12124,N_12680);
xor U13973 (N_13973,N_12440,N_12759);
nand U13974 (N_13974,N_12406,N_12466);
xor U13975 (N_13975,N_12583,N_12825);
nor U13976 (N_13976,N_12698,N_12371);
xnor U13977 (N_13977,N_12555,N_12086);
nand U13978 (N_13978,N_12299,N_12555);
nor U13979 (N_13979,N_12926,N_12031);
or U13980 (N_13980,N_12368,N_12890);
and U13981 (N_13981,N_12660,N_12861);
and U13982 (N_13982,N_12820,N_12894);
nand U13983 (N_13983,N_12721,N_12958);
xnor U13984 (N_13984,N_12981,N_12922);
nand U13985 (N_13985,N_12719,N_12869);
or U13986 (N_13986,N_12954,N_12931);
or U13987 (N_13987,N_12995,N_12474);
nor U13988 (N_13988,N_12012,N_12402);
nor U13989 (N_13989,N_12772,N_12937);
and U13990 (N_13990,N_12909,N_12381);
nand U13991 (N_13991,N_12237,N_12755);
or U13992 (N_13992,N_12292,N_12512);
or U13993 (N_13993,N_12465,N_12977);
nor U13994 (N_13994,N_12239,N_12058);
and U13995 (N_13995,N_12873,N_12293);
xnor U13996 (N_13996,N_12171,N_12974);
xor U13997 (N_13997,N_12061,N_12833);
or U13998 (N_13998,N_12139,N_12383);
nor U13999 (N_13999,N_12974,N_12154);
nand U14000 (N_14000,N_13489,N_13618);
nor U14001 (N_14001,N_13832,N_13148);
nand U14002 (N_14002,N_13919,N_13781);
and U14003 (N_14003,N_13518,N_13596);
nor U14004 (N_14004,N_13927,N_13532);
nor U14005 (N_14005,N_13437,N_13225);
nor U14006 (N_14006,N_13341,N_13971);
nand U14007 (N_14007,N_13878,N_13805);
xor U14008 (N_14008,N_13821,N_13775);
or U14009 (N_14009,N_13553,N_13807);
xor U14010 (N_14010,N_13755,N_13824);
xor U14011 (N_14011,N_13817,N_13865);
nor U14012 (N_14012,N_13229,N_13051);
xnor U14013 (N_14013,N_13132,N_13086);
nand U14014 (N_14014,N_13862,N_13870);
or U14015 (N_14015,N_13448,N_13970);
xor U14016 (N_14016,N_13520,N_13257);
nor U14017 (N_14017,N_13439,N_13203);
and U14018 (N_14018,N_13026,N_13994);
nor U14019 (N_14019,N_13679,N_13839);
xor U14020 (N_14020,N_13285,N_13370);
nand U14021 (N_14021,N_13393,N_13101);
or U14022 (N_14022,N_13571,N_13277);
nand U14023 (N_14023,N_13294,N_13055);
nor U14024 (N_14024,N_13222,N_13117);
nand U14025 (N_14025,N_13706,N_13872);
nor U14026 (N_14026,N_13302,N_13897);
and U14027 (N_14027,N_13417,N_13295);
xnor U14028 (N_14028,N_13627,N_13435);
nand U14029 (N_14029,N_13179,N_13178);
nand U14030 (N_14030,N_13834,N_13092);
or U14031 (N_14031,N_13748,N_13703);
or U14032 (N_14032,N_13044,N_13979);
and U14033 (N_14033,N_13153,N_13105);
nor U14034 (N_14034,N_13264,N_13884);
and U14035 (N_14035,N_13660,N_13898);
or U14036 (N_14036,N_13053,N_13737);
xnor U14037 (N_14037,N_13646,N_13658);
or U14038 (N_14038,N_13586,N_13918);
and U14039 (N_14039,N_13033,N_13461);
xor U14040 (N_14040,N_13736,N_13836);
xnor U14041 (N_14041,N_13759,N_13367);
and U14042 (N_14042,N_13364,N_13621);
nand U14043 (N_14043,N_13497,N_13459);
nor U14044 (N_14044,N_13454,N_13280);
nor U14045 (N_14045,N_13546,N_13920);
nand U14046 (N_14046,N_13882,N_13813);
xnor U14047 (N_14047,N_13510,N_13485);
nor U14048 (N_14048,N_13482,N_13268);
nor U14049 (N_14049,N_13355,N_13296);
and U14050 (N_14050,N_13320,N_13058);
xnor U14051 (N_14051,N_13360,N_13182);
or U14052 (N_14052,N_13931,N_13456);
and U14053 (N_14053,N_13568,N_13964);
and U14054 (N_14054,N_13036,N_13321);
or U14055 (N_14055,N_13120,N_13893);
xor U14056 (N_14056,N_13168,N_13123);
nand U14057 (N_14057,N_13035,N_13198);
xnor U14058 (N_14058,N_13030,N_13413);
and U14059 (N_14059,N_13206,N_13625);
nor U14060 (N_14060,N_13386,N_13316);
and U14061 (N_14061,N_13709,N_13351);
nor U14062 (N_14062,N_13371,N_13157);
or U14063 (N_14063,N_13756,N_13921);
or U14064 (N_14064,N_13833,N_13039);
and U14065 (N_14065,N_13125,N_13126);
nor U14066 (N_14066,N_13438,N_13056);
nor U14067 (N_14067,N_13721,N_13276);
nor U14068 (N_14068,N_13040,N_13134);
and U14069 (N_14069,N_13619,N_13152);
and U14070 (N_14070,N_13701,N_13659);
or U14071 (N_14071,N_13888,N_13477);
and U14072 (N_14072,N_13547,N_13585);
nor U14073 (N_14073,N_13233,N_13366);
nand U14074 (N_14074,N_13905,N_13318);
and U14075 (N_14075,N_13488,N_13758);
xor U14076 (N_14076,N_13790,N_13702);
xor U14077 (N_14077,N_13800,N_13672);
nor U14078 (N_14078,N_13440,N_13717);
xnor U14079 (N_14079,N_13550,N_13972);
or U14080 (N_14080,N_13106,N_13292);
nand U14081 (N_14081,N_13667,N_13904);
nand U14082 (N_14082,N_13473,N_13326);
nand U14083 (N_14083,N_13691,N_13981);
or U14084 (N_14084,N_13275,N_13772);
nor U14085 (N_14085,N_13365,N_13543);
nand U14086 (N_14086,N_13825,N_13572);
and U14087 (N_14087,N_13840,N_13259);
xor U14088 (N_14088,N_13648,N_13782);
nand U14089 (N_14089,N_13034,N_13287);
xnor U14090 (N_14090,N_13348,N_13591);
xor U14091 (N_14091,N_13804,N_13031);
nand U14092 (N_14092,N_13284,N_13094);
xnor U14093 (N_14093,N_13216,N_13629);
or U14094 (N_14094,N_13845,N_13345);
and U14095 (N_14095,N_13029,N_13687);
xnor U14096 (N_14096,N_13849,N_13688);
nand U14097 (N_14097,N_13556,N_13457);
or U14098 (N_14098,N_13997,N_13963);
or U14099 (N_14099,N_13502,N_13795);
nand U14100 (N_14100,N_13171,N_13697);
and U14101 (N_14101,N_13463,N_13262);
nand U14102 (N_14102,N_13575,N_13899);
and U14103 (N_14103,N_13140,N_13911);
or U14104 (N_14104,N_13490,N_13147);
nor U14105 (N_14105,N_13181,N_13993);
nor U14106 (N_14106,N_13323,N_13549);
nor U14107 (N_14107,N_13398,N_13496);
and U14108 (N_14108,N_13559,N_13760);
or U14109 (N_14109,N_13347,N_13065);
or U14110 (N_14110,N_13534,N_13923);
or U14111 (N_14111,N_13630,N_13339);
nor U14112 (N_14112,N_13633,N_13976);
nand U14113 (N_14113,N_13769,N_13666);
or U14114 (N_14114,N_13680,N_13192);
xor U14115 (N_14115,N_13467,N_13723);
and U14116 (N_14116,N_13372,N_13357);
nor U14117 (N_14117,N_13169,N_13661);
nand U14118 (N_14118,N_13059,N_13214);
nor U14119 (N_14119,N_13244,N_13221);
nor U14120 (N_14120,N_13005,N_13910);
nor U14121 (N_14121,N_13241,N_13530);
and U14122 (N_14122,N_13838,N_13067);
xnor U14123 (N_14123,N_13319,N_13279);
nor U14124 (N_14124,N_13451,N_13852);
nand U14125 (N_14125,N_13460,N_13445);
and U14126 (N_14126,N_13606,N_13803);
nand U14127 (N_14127,N_13443,N_13242);
and U14128 (N_14128,N_13462,N_13476);
or U14129 (N_14129,N_13024,N_13087);
and U14130 (N_14130,N_13552,N_13853);
or U14131 (N_14131,N_13074,N_13137);
and U14132 (N_14132,N_13388,N_13327);
and U14133 (N_14133,N_13391,N_13639);
nand U14134 (N_14134,N_13762,N_13004);
or U14135 (N_14135,N_13990,N_13806);
and U14136 (N_14136,N_13215,N_13917);
nand U14137 (N_14137,N_13542,N_13789);
or U14138 (N_14138,N_13733,N_13317);
xor U14139 (N_14139,N_13195,N_13421);
and U14140 (N_14140,N_13708,N_13934);
nand U14141 (N_14141,N_13566,N_13631);
and U14142 (N_14142,N_13634,N_13042);
nor U14143 (N_14143,N_13522,N_13097);
or U14144 (N_14144,N_13871,N_13114);
nand U14145 (N_14145,N_13232,N_13499);
or U14146 (N_14146,N_13901,N_13382);
or U14147 (N_14147,N_13263,N_13239);
or U14148 (N_14148,N_13980,N_13777);
xor U14149 (N_14149,N_13635,N_13186);
nand U14150 (N_14150,N_13731,N_13397);
or U14151 (N_14151,N_13307,N_13512);
or U14152 (N_14152,N_13113,N_13465);
nor U14153 (N_14153,N_13765,N_13955);
nand U14154 (N_14154,N_13309,N_13098);
or U14155 (N_14155,N_13342,N_13643);
and U14156 (N_14156,N_13330,N_13536);
xor U14157 (N_14157,N_13442,N_13669);
or U14158 (N_14158,N_13681,N_13592);
and U14159 (N_14159,N_13541,N_13404);
nand U14160 (N_14160,N_13551,N_13902);
nor U14161 (N_14161,N_13304,N_13109);
nand U14162 (N_14162,N_13662,N_13859);
nor U14163 (N_14163,N_13656,N_13582);
and U14164 (N_14164,N_13025,N_13607);
nor U14165 (N_14165,N_13715,N_13017);
and U14166 (N_14166,N_13686,N_13692);
nand U14167 (N_14167,N_13811,N_13243);
nand U14168 (N_14168,N_13819,N_13190);
and U14169 (N_14169,N_13091,N_13315);
xnor U14170 (N_14170,N_13245,N_13486);
xnor U14171 (N_14171,N_13332,N_13632);
xnor U14172 (N_14172,N_13193,N_13450);
or U14173 (N_14173,N_13752,N_13900);
nand U14174 (N_14174,N_13914,N_13150);
nand U14175 (N_14175,N_13487,N_13930);
and U14176 (N_14176,N_13954,N_13768);
nor U14177 (N_14177,N_13481,N_13107);
nor U14178 (N_14178,N_13174,N_13533);
nand U14179 (N_14179,N_13828,N_13857);
nor U14180 (N_14180,N_13061,N_13118);
nor U14181 (N_14181,N_13589,N_13308);
nor U14182 (N_14182,N_13776,N_13141);
nand U14183 (N_14183,N_13331,N_13563);
or U14184 (N_14184,N_13949,N_13475);
xnor U14185 (N_14185,N_13281,N_13016);
and U14186 (N_14186,N_13472,N_13139);
and U14187 (N_14187,N_13410,N_13427);
or U14188 (N_14188,N_13735,N_13945);
xor U14189 (N_14189,N_13373,N_13299);
nor U14190 (N_14190,N_13389,N_13506);
xor U14191 (N_14191,N_13060,N_13887);
and U14192 (N_14192,N_13324,N_13773);
nand U14193 (N_14193,N_13835,N_13915);
and U14194 (N_14194,N_13100,N_13064);
or U14195 (N_14195,N_13217,N_13256);
nor U14196 (N_14196,N_13414,N_13802);
xor U14197 (N_14197,N_13238,N_13711);
and U14198 (N_14198,N_13785,N_13652);
xnor U14199 (N_14199,N_13780,N_13753);
nor U14200 (N_14200,N_13283,N_13492);
or U14201 (N_14201,N_13668,N_13479);
or U14202 (N_14202,N_13260,N_13778);
or U14203 (N_14203,N_13224,N_13858);
nand U14204 (N_14204,N_13088,N_13713);
nor U14205 (N_14205,N_13602,N_13986);
xor U14206 (N_14206,N_13555,N_13188);
nor U14207 (N_14207,N_13503,N_13941);
and U14208 (N_14208,N_13590,N_13998);
or U14209 (N_14209,N_13588,N_13164);
nand U14210 (N_14210,N_13535,N_13526);
nand U14211 (N_14211,N_13982,N_13185);
nor U14212 (N_14212,N_13663,N_13809);
or U14213 (N_14213,N_13237,N_13749);
nand U14214 (N_14214,N_13167,N_13199);
and U14215 (N_14215,N_13474,N_13218);
nor U14216 (N_14216,N_13724,N_13129);
nand U14217 (N_14217,N_13890,N_13583);
xor U14218 (N_14218,N_13396,N_13407);
nor U14219 (N_14219,N_13261,N_13162);
or U14220 (N_14220,N_13430,N_13622);
or U14221 (N_14221,N_13343,N_13049);
nand U14222 (N_14222,N_13289,N_13842);
nand U14223 (N_14223,N_13306,N_13310);
nor U14224 (N_14224,N_13075,N_13494);
nor U14225 (N_14225,N_13202,N_13464);
or U14226 (N_14226,N_13201,N_13587);
and U14227 (N_14227,N_13411,N_13651);
nor U14228 (N_14228,N_13368,N_13952);
nand U14229 (N_14229,N_13999,N_13846);
xnor U14230 (N_14230,N_13626,N_13558);
nand U14231 (N_14231,N_13767,N_13598);
or U14232 (N_14232,N_13693,N_13291);
xor U14233 (N_14233,N_13400,N_13957);
or U14234 (N_14234,N_13154,N_13507);
nand U14235 (N_14235,N_13014,N_13788);
or U14236 (N_14236,N_13615,N_13340);
nor U14237 (N_14237,N_13314,N_13160);
or U14238 (N_14238,N_13246,N_13557);
nand U14239 (N_14239,N_13251,N_13424);
nor U14240 (N_14240,N_13358,N_13070);
xnor U14241 (N_14241,N_13678,N_13922);
xnor U14242 (N_14242,N_13151,N_13664);
xnor U14243 (N_14243,N_13783,N_13798);
or U14244 (N_14244,N_13740,N_13929);
xor U14245 (N_14245,N_13468,N_13328);
nand U14246 (N_14246,N_13333,N_13995);
and U14247 (N_14247,N_13223,N_13066);
nor U14248 (N_14248,N_13637,N_13676);
nor U14249 (N_14249,N_13418,N_13799);
or U14250 (N_14250,N_13714,N_13210);
nor U14251 (N_14251,N_13511,N_13581);
xor U14252 (N_14252,N_13916,N_13329);
and U14253 (N_14253,N_13002,N_13127);
nand U14254 (N_14254,N_13903,N_13027);
and U14255 (N_14255,N_13992,N_13612);
and U14256 (N_14256,N_13829,N_13376);
nor U14257 (N_14257,N_13390,N_13948);
and U14258 (N_14258,N_13613,N_13211);
or U14259 (N_14259,N_13471,N_13936);
xnor U14260 (N_14260,N_13278,N_13718);
or U14261 (N_14261,N_13253,N_13081);
nand U14262 (N_14262,N_13861,N_13077);
xor U14263 (N_14263,N_13774,N_13924);
nand U14264 (N_14264,N_13197,N_13975);
xor U14265 (N_14265,N_13548,N_13796);
nor U14266 (N_14266,N_13416,N_13823);
nor U14267 (N_14267,N_13599,N_13848);
nor U14268 (N_14268,N_13739,N_13394);
or U14269 (N_14269,N_13521,N_13335);
xnor U14270 (N_14270,N_13009,N_13868);
and U14271 (N_14271,N_13111,N_13022);
or U14272 (N_14272,N_13729,N_13951);
nor U14273 (N_14273,N_13983,N_13742);
and U14274 (N_14274,N_13699,N_13399);
nor U14275 (N_14275,N_13766,N_13433);
nor U14276 (N_14276,N_13529,N_13851);
and U14277 (N_14277,N_13793,N_13973);
xnor U14278 (N_14278,N_13205,N_13158);
nand U14279 (N_14279,N_13191,N_13977);
nor U14280 (N_14280,N_13079,N_13072);
nor U14281 (N_14281,N_13093,N_13144);
and U14282 (N_14282,N_13712,N_13392);
or U14283 (N_14283,N_13562,N_13353);
and U14284 (N_14284,N_13743,N_13677);
and U14285 (N_14285,N_13584,N_13083);
nand U14286 (N_14286,N_13670,N_13683);
nand U14287 (N_14287,N_13883,N_13565);
or U14288 (N_14288,N_13354,N_13933);
and U14289 (N_14289,N_13786,N_13705);
nand U14290 (N_14290,N_13272,N_13213);
and U14291 (N_14291,N_13968,N_13466);
nor U14292 (N_14292,N_13322,N_13441);
xor U14293 (N_14293,N_13010,N_13363);
nand U14294 (N_14294,N_13401,N_13844);
and U14295 (N_14295,N_13513,N_13818);
nor U14296 (N_14296,N_13493,N_13704);
nand U14297 (N_14297,N_13038,N_13913);
or U14298 (N_14298,N_13946,N_13112);
nor U14299 (N_14299,N_13978,N_13636);
nand U14300 (N_14300,N_13956,N_13876);
xnor U14301 (N_14301,N_13644,N_13751);
or U14302 (N_14302,N_13344,N_13674);
xor U14303 (N_14303,N_13909,N_13425);
or U14304 (N_14304,N_13727,N_13003);
nand U14305 (N_14305,N_13537,N_13642);
xnor U14306 (N_14306,N_13236,N_13624);
nor U14307 (N_14307,N_13048,N_13671);
xnor U14308 (N_14308,N_13734,N_13082);
and U14309 (N_14309,N_13008,N_13124);
nor U14310 (N_14310,N_13227,N_13231);
and U14311 (N_14311,N_13271,N_13987);
or U14312 (N_14312,N_13928,N_13935);
or U14313 (N_14313,N_13645,N_13561);
nor U14314 (N_14314,N_13050,N_13614);
nand U14315 (N_14315,N_13267,N_13886);
xor U14316 (N_14316,N_13896,N_13128);
xor U14317 (N_14317,N_13000,N_13073);
or U14318 (N_14318,N_13593,N_13657);
or U14319 (N_14319,N_13089,N_13047);
nor U14320 (N_14320,N_13710,N_13429);
nor U14321 (N_14321,N_13207,N_13447);
and U14322 (N_14322,N_13528,N_13006);
xor U14323 (N_14323,N_13062,N_13515);
or U14324 (N_14324,N_13266,N_13177);
nand U14325 (N_14325,N_13453,N_13426);
and U14326 (N_14326,N_13122,N_13673);
xnor U14327 (N_14327,N_13784,N_13078);
or U14328 (N_14328,N_13495,N_13569);
and U14329 (N_14329,N_13754,N_13801);
and U14330 (N_14330,N_13880,N_13133);
and U14331 (N_14331,N_13716,N_13046);
and U14332 (N_14332,N_13538,N_13791);
nor U14333 (N_14333,N_13170,N_13020);
or U14334 (N_14334,N_13325,N_13436);
or U14335 (N_14335,N_13269,N_13084);
or U14336 (N_14336,N_13184,N_13045);
nand U14337 (N_14337,N_13362,N_13043);
xnor U14338 (N_14338,N_13578,N_13406);
xnor U14339 (N_14339,N_13240,N_13069);
and U14340 (N_14340,N_13402,N_13722);
nand U14341 (N_14341,N_13810,N_13194);
or U14342 (N_14342,N_13469,N_13820);
and U14343 (N_14343,N_13480,N_13385);
nor U14344 (N_14344,N_13580,N_13369);
xor U14345 (N_14345,N_13301,N_13270);
and U14346 (N_14346,N_13690,N_13096);
nor U14347 (N_14347,N_13564,N_13432);
and U14348 (N_14348,N_13290,N_13252);
or U14349 (N_14349,N_13808,N_13455);
nor U14350 (N_14350,N_13505,N_13054);
nor U14351 (N_14351,N_13166,N_13962);
xnor U14352 (N_14352,N_13063,N_13514);
xor U14353 (N_14353,N_13080,N_13208);
and U14354 (N_14354,N_13012,N_13491);
nand U14355 (N_14355,N_13349,N_13119);
or U14356 (N_14356,N_13604,N_13187);
or U14357 (N_14357,N_13867,N_13746);
nor U14358 (N_14358,N_13570,N_13816);
and U14359 (N_14359,N_13508,N_13961);
xor U14360 (N_14360,N_13273,N_13444);
xor U14361 (N_14361,N_13356,N_13408);
nand U14362 (N_14362,N_13984,N_13189);
and U14363 (N_14363,N_13866,N_13745);
or U14364 (N_14364,N_13605,N_13761);
nor U14365 (N_14365,N_13787,N_13594);
xnor U14366 (N_14366,N_13940,N_13311);
or U14367 (N_14367,N_13350,N_13452);
xnor U14368 (N_14368,N_13682,N_13741);
nand U14369 (N_14369,N_13212,N_13869);
xor U14370 (N_14370,N_13675,N_13361);
nor U14371 (N_14371,N_13937,N_13312);
or U14372 (N_14372,N_13959,N_13966);
and U14373 (N_14373,N_13611,N_13540);
and U14374 (N_14374,N_13830,N_13303);
xnor U14375 (N_14375,N_13110,N_13728);
xor U14376 (N_14376,N_13085,N_13374);
nor U14377 (N_14377,N_13274,N_13149);
nand U14378 (N_14378,N_13359,N_13384);
or U14379 (N_14379,N_13943,N_13653);
and U14380 (N_14380,N_13763,N_13601);
xnor U14381 (N_14381,N_13131,N_13875);
xor U14382 (N_14382,N_13792,N_13831);
xnor U14383 (N_14383,N_13172,N_13856);
or U14384 (N_14384,N_13932,N_13595);
xnor U14385 (N_14385,N_13747,N_13235);
xor U14386 (N_14386,N_13864,N_13879);
xor U14387 (N_14387,N_13509,N_13300);
or U14388 (N_14388,N_13874,N_13527);
or U14389 (N_14389,N_13104,N_13379);
and U14390 (N_14390,N_13814,N_13597);
nor U14391 (N_14391,N_13220,N_13422);
nor U14392 (N_14392,N_13484,N_13173);
xnor U14393 (N_14393,N_13011,N_13628);
nor U14394 (N_14394,N_13052,N_13609);
and U14395 (N_14395,N_13608,N_13163);
nand U14396 (N_14396,N_13574,N_13947);
nand U14397 (N_14397,N_13873,N_13337);
and U14398 (N_14398,N_13116,N_13617);
nand U14399 (N_14399,N_13577,N_13576);
and U14400 (N_14400,N_13375,N_13944);
xor U14401 (N_14401,N_13684,N_13383);
xnor U14402 (N_14402,N_13130,N_13544);
xor U14403 (N_14403,N_13090,N_13431);
or U14404 (N_14404,N_13906,N_13458);
and U14405 (N_14405,N_13286,N_13726);
nand U14406 (N_14406,N_13738,N_13881);
nand U14407 (N_14407,N_13560,N_13007);
and U14408 (N_14408,N_13183,N_13750);
nand U14409 (N_14409,N_13732,N_13265);
or U14410 (N_14410,N_13524,N_13019);
or U14411 (N_14411,N_13689,N_13757);
or U14412 (N_14412,N_13837,N_13950);
nand U14413 (N_14413,N_13381,N_13665);
nand U14414 (N_14414,N_13305,N_13988);
xor U14415 (N_14415,N_13143,N_13942);
and U14416 (N_14416,N_13135,N_13640);
nor U14417 (N_14417,N_13145,N_13121);
xor U14418 (N_14418,N_13478,N_13226);
nor U14419 (N_14419,N_13771,N_13412);
or U14420 (N_14420,N_13654,N_13209);
or U14421 (N_14421,N_13891,N_13200);
xor U14422 (N_14422,N_13960,N_13338);
nor U14423 (N_14423,N_13623,N_13554);
and U14424 (N_14424,N_13420,N_13037);
or U14425 (N_14425,N_13403,N_13099);
and U14426 (N_14426,N_13523,N_13254);
xnor U14427 (N_14427,N_13969,N_13539);
nor U14428 (N_14428,N_13965,N_13610);
and U14429 (N_14429,N_13655,N_13707);
nand U14430 (N_14430,N_13519,N_13579);
nand U14431 (N_14431,N_13854,N_13926);
and U14432 (N_14432,N_13641,N_13255);
xnor U14433 (N_14433,N_13288,N_13377);
and U14434 (N_14434,N_13531,N_13146);
or U14435 (N_14435,N_13649,N_13647);
xnor U14436 (N_14436,N_13638,N_13395);
xnor U14437 (N_14437,N_13352,N_13068);
nand U14438 (N_14438,N_13908,N_13219);
nor U14439 (N_14439,N_13504,N_13812);
and U14440 (N_14440,N_13380,N_13567);
or U14441 (N_14441,N_13293,N_13863);
nand U14442 (N_14442,N_13415,N_13603);
and U14443 (N_14443,N_13938,N_13015);
nand U14444 (N_14444,N_13071,N_13847);
xor U14445 (N_14445,N_13161,N_13387);
xor U14446 (N_14446,N_13449,N_13860);
and U14447 (N_14447,N_13958,N_13939);
xor U14448 (N_14448,N_13248,N_13405);
nor U14449 (N_14449,N_13855,N_13907);
xor U14450 (N_14450,N_13138,N_13770);
or U14451 (N_14451,N_13719,N_13041);
nor U14452 (N_14452,N_13013,N_13779);
nand U14453 (N_14453,N_13889,N_13498);
nand U14454 (N_14454,N_13953,N_13698);
xnor U14455 (N_14455,N_13346,N_13925);
nor U14456 (N_14456,N_13985,N_13912);
xnor U14457 (N_14457,N_13827,N_13843);
and U14458 (N_14458,N_13234,N_13685);
or U14459 (N_14459,N_13165,N_13794);
nor U14460 (N_14460,N_13028,N_13516);
nor U14461 (N_14461,N_13620,N_13103);
nand U14462 (N_14462,N_13517,N_13470);
and U14463 (N_14463,N_13298,N_13996);
xor U14464 (N_14464,N_13730,N_13650);
and U14465 (N_14465,N_13336,N_13989);
or U14466 (N_14466,N_13032,N_13545);
and U14467 (N_14467,N_13700,N_13378);
and U14468 (N_14468,N_13720,N_13196);
nand U14469 (N_14469,N_13744,N_13822);
nand U14470 (N_14470,N_13419,N_13204);
or U14471 (N_14471,N_13616,N_13115);
nor U14472 (N_14472,N_13500,N_13695);
xor U14473 (N_14473,N_13282,N_13483);
or U14474 (N_14474,N_13018,N_13076);
nor U14475 (N_14475,N_13155,N_13892);
xnor U14476 (N_14476,N_13423,N_13230);
xor U14477 (N_14477,N_13102,N_13815);
nor U14478 (N_14478,N_13967,N_13885);
nor U14479 (N_14479,N_13991,N_13694);
nand U14480 (N_14480,N_13764,N_13156);
and U14481 (N_14481,N_13095,N_13850);
nor U14482 (N_14482,N_13446,N_13434);
and U14483 (N_14483,N_13247,N_13826);
nand U14484 (N_14484,N_13409,N_13428);
nor U14485 (N_14485,N_13057,N_13313);
and U14486 (N_14486,N_13877,N_13142);
nand U14487 (N_14487,N_13258,N_13175);
xnor U14488 (N_14488,N_13108,N_13297);
or U14489 (N_14489,N_13573,N_13974);
and U14490 (N_14490,N_13136,N_13250);
xor U14491 (N_14491,N_13249,N_13600);
nand U14492 (N_14492,N_13021,N_13334);
nand U14493 (N_14493,N_13895,N_13894);
xnor U14494 (N_14494,N_13725,N_13696);
and U14495 (N_14495,N_13841,N_13797);
nand U14496 (N_14496,N_13159,N_13180);
and U14497 (N_14497,N_13176,N_13001);
xor U14498 (N_14498,N_13228,N_13023);
or U14499 (N_14499,N_13501,N_13525);
and U14500 (N_14500,N_13105,N_13389);
xor U14501 (N_14501,N_13138,N_13702);
or U14502 (N_14502,N_13181,N_13322);
or U14503 (N_14503,N_13881,N_13882);
and U14504 (N_14504,N_13464,N_13367);
nor U14505 (N_14505,N_13680,N_13187);
and U14506 (N_14506,N_13820,N_13594);
and U14507 (N_14507,N_13517,N_13424);
and U14508 (N_14508,N_13286,N_13624);
or U14509 (N_14509,N_13138,N_13928);
or U14510 (N_14510,N_13398,N_13521);
or U14511 (N_14511,N_13752,N_13368);
and U14512 (N_14512,N_13401,N_13686);
xor U14513 (N_14513,N_13561,N_13063);
and U14514 (N_14514,N_13422,N_13084);
nor U14515 (N_14515,N_13936,N_13636);
and U14516 (N_14516,N_13491,N_13826);
xnor U14517 (N_14517,N_13610,N_13269);
and U14518 (N_14518,N_13729,N_13807);
nand U14519 (N_14519,N_13967,N_13174);
and U14520 (N_14520,N_13407,N_13228);
xnor U14521 (N_14521,N_13864,N_13138);
nand U14522 (N_14522,N_13723,N_13680);
or U14523 (N_14523,N_13243,N_13082);
and U14524 (N_14524,N_13935,N_13070);
and U14525 (N_14525,N_13958,N_13697);
nor U14526 (N_14526,N_13586,N_13636);
xor U14527 (N_14527,N_13321,N_13207);
xor U14528 (N_14528,N_13292,N_13376);
and U14529 (N_14529,N_13520,N_13177);
xor U14530 (N_14530,N_13593,N_13200);
xnor U14531 (N_14531,N_13146,N_13399);
nor U14532 (N_14532,N_13897,N_13256);
nand U14533 (N_14533,N_13328,N_13205);
nor U14534 (N_14534,N_13481,N_13613);
xnor U14535 (N_14535,N_13032,N_13433);
xor U14536 (N_14536,N_13226,N_13939);
nand U14537 (N_14537,N_13436,N_13539);
nor U14538 (N_14538,N_13399,N_13578);
or U14539 (N_14539,N_13963,N_13415);
nand U14540 (N_14540,N_13541,N_13998);
xnor U14541 (N_14541,N_13383,N_13087);
nor U14542 (N_14542,N_13617,N_13923);
nand U14543 (N_14543,N_13987,N_13246);
xor U14544 (N_14544,N_13597,N_13716);
and U14545 (N_14545,N_13872,N_13259);
or U14546 (N_14546,N_13527,N_13546);
and U14547 (N_14547,N_13152,N_13371);
nor U14548 (N_14548,N_13163,N_13700);
or U14549 (N_14549,N_13588,N_13667);
nor U14550 (N_14550,N_13573,N_13150);
or U14551 (N_14551,N_13441,N_13507);
nand U14552 (N_14552,N_13489,N_13445);
xnor U14553 (N_14553,N_13956,N_13200);
nand U14554 (N_14554,N_13619,N_13963);
nand U14555 (N_14555,N_13699,N_13547);
xnor U14556 (N_14556,N_13215,N_13291);
nand U14557 (N_14557,N_13316,N_13352);
or U14558 (N_14558,N_13318,N_13598);
and U14559 (N_14559,N_13926,N_13697);
nor U14560 (N_14560,N_13721,N_13874);
xnor U14561 (N_14561,N_13383,N_13926);
and U14562 (N_14562,N_13744,N_13497);
and U14563 (N_14563,N_13884,N_13044);
nand U14564 (N_14564,N_13270,N_13920);
nand U14565 (N_14565,N_13724,N_13396);
xor U14566 (N_14566,N_13953,N_13516);
and U14567 (N_14567,N_13242,N_13001);
and U14568 (N_14568,N_13662,N_13652);
nor U14569 (N_14569,N_13623,N_13920);
and U14570 (N_14570,N_13719,N_13219);
and U14571 (N_14571,N_13522,N_13171);
xnor U14572 (N_14572,N_13961,N_13440);
or U14573 (N_14573,N_13628,N_13248);
xnor U14574 (N_14574,N_13045,N_13585);
nand U14575 (N_14575,N_13770,N_13003);
xor U14576 (N_14576,N_13994,N_13301);
nor U14577 (N_14577,N_13065,N_13715);
nand U14578 (N_14578,N_13339,N_13694);
nor U14579 (N_14579,N_13604,N_13292);
or U14580 (N_14580,N_13737,N_13374);
nor U14581 (N_14581,N_13318,N_13132);
nor U14582 (N_14582,N_13819,N_13053);
or U14583 (N_14583,N_13141,N_13129);
or U14584 (N_14584,N_13057,N_13067);
nor U14585 (N_14585,N_13828,N_13060);
xnor U14586 (N_14586,N_13655,N_13962);
and U14587 (N_14587,N_13601,N_13232);
nor U14588 (N_14588,N_13906,N_13375);
nand U14589 (N_14589,N_13595,N_13135);
and U14590 (N_14590,N_13246,N_13732);
nand U14591 (N_14591,N_13918,N_13616);
or U14592 (N_14592,N_13978,N_13621);
xor U14593 (N_14593,N_13893,N_13815);
xnor U14594 (N_14594,N_13442,N_13476);
or U14595 (N_14595,N_13772,N_13513);
nand U14596 (N_14596,N_13601,N_13270);
or U14597 (N_14597,N_13657,N_13568);
and U14598 (N_14598,N_13669,N_13436);
nor U14599 (N_14599,N_13068,N_13198);
nor U14600 (N_14600,N_13578,N_13334);
and U14601 (N_14601,N_13914,N_13298);
and U14602 (N_14602,N_13089,N_13618);
and U14603 (N_14603,N_13820,N_13356);
nand U14604 (N_14604,N_13455,N_13766);
nor U14605 (N_14605,N_13404,N_13432);
nor U14606 (N_14606,N_13894,N_13418);
or U14607 (N_14607,N_13373,N_13921);
xnor U14608 (N_14608,N_13330,N_13875);
or U14609 (N_14609,N_13866,N_13705);
or U14610 (N_14610,N_13590,N_13925);
nand U14611 (N_14611,N_13928,N_13298);
nor U14612 (N_14612,N_13917,N_13606);
or U14613 (N_14613,N_13098,N_13958);
or U14614 (N_14614,N_13375,N_13655);
and U14615 (N_14615,N_13512,N_13362);
or U14616 (N_14616,N_13401,N_13309);
nand U14617 (N_14617,N_13294,N_13223);
nor U14618 (N_14618,N_13510,N_13138);
xnor U14619 (N_14619,N_13878,N_13728);
and U14620 (N_14620,N_13679,N_13217);
nor U14621 (N_14621,N_13914,N_13390);
nor U14622 (N_14622,N_13807,N_13455);
nor U14623 (N_14623,N_13609,N_13687);
and U14624 (N_14624,N_13039,N_13047);
and U14625 (N_14625,N_13491,N_13180);
and U14626 (N_14626,N_13193,N_13847);
nor U14627 (N_14627,N_13383,N_13592);
xnor U14628 (N_14628,N_13566,N_13192);
nand U14629 (N_14629,N_13237,N_13352);
nand U14630 (N_14630,N_13021,N_13104);
or U14631 (N_14631,N_13179,N_13253);
xnor U14632 (N_14632,N_13640,N_13317);
or U14633 (N_14633,N_13602,N_13591);
nand U14634 (N_14634,N_13329,N_13751);
nand U14635 (N_14635,N_13613,N_13203);
xor U14636 (N_14636,N_13842,N_13407);
nor U14637 (N_14637,N_13321,N_13857);
xor U14638 (N_14638,N_13850,N_13933);
and U14639 (N_14639,N_13431,N_13660);
xor U14640 (N_14640,N_13467,N_13279);
or U14641 (N_14641,N_13389,N_13541);
xor U14642 (N_14642,N_13407,N_13212);
xor U14643 (N_14643,N_13073,N_13616);
or U14644 (N_14644,N_13184,N_13464);
and U14645 (N_14645,N_13403,N_13515);
nand U14646 (N_14646,N_13921,N_13197);
xnor U14647 (N_14647,N_13114,N_13368);
nand U14648 (N_14648,N_13102,N_13588);
and U14649 (N_14649,N_13079,N_13425);
or U14650 (N_14650,N_13228,N_13768);
nor U14651 (N_14651,N_13165,N_13379);
nor U14652 (N_14652,N_13323,N_13180);
nor U14653 (N_14653,N_13695,N_13807);
and U14654 (N_14654,N_13829,N_13355);
and U14655 (N_14655,N_13914,N_13477);
or U14656 (N_14656,N_13369,N_13051);
nand U14657 (N_14657,N_13736,N_13848);
nand U14658 (N_14658,N_13980,N_13672);
nor U14659 (N_14659,N_13711,N_13676);
and U14660 (N_14660,N_13742,N_13327);
or U14661 (N_14661,N_13428,N_13834);
xnor U14662 (N_14662,N_13082,N_13112);
and U14663 (N_14663,N_13034,N_13602);
and U14664 (N_14664,N_13227,N_13368);
and U14665 (N_14665,N_13507,N_13468);
and U14666 (N_14666,N_13301,N_13057);
or U14667 (N_14667,N_13578,N_13281);
or U14668 (N_14668,N_13838,N_13362);
and U14669 (N_14669,N_13891,N_13430);
nor U14670 (N_14670,N_13935,N_13415);
nand U14671 (N_14671,N_13932,N_13157);
or U14672 (N_14672,N_13244,N_13322);
and U14673 (N_14673,N_13283,N_13864);
nand U14674 (N_14674,N_13357,N_13860);
nand U14675 (N_14675,N_13945,N_13412);
nor U14676 (N_14676,N_13898,N_13140);
and U14677 (N_14677,N_13587,N_13352);
and U14678 (N_14678,N_13728,N_13941);
nor U14679 (N_14679,N_13658,N_13746);
or U14680 (N_14680,N_13227,N_13203);
nor U14681 (N_14681,N_13787,N_13694);
nand U14682 (N_14682,N_13286,N_13937);
or U14683 (N_14683,N_13007,N_13162);
xnor U14684 (N_14684,N_13731,N_13437);
and U14685 (N_14685,N_13208,N_13985);
and U14686 (N_14686,N_13374,N_13659);
and U14687 (N_14687,N_13404,N_13878);
or U14688 (N_14688,N_13423,N_13817);
nor U14689 (N_14689,N_13909,N_13740);
or U14690 (N_14690,N_13457,N_13845);
or U14691 (N_14691,N_13955,N_13050);
xor U14692 (N_14692,N_13984,N_13490);
nor U14693 (N_14693,N_13075,N_13905);
and U14694 (N_14694,N_13132,N_13085);
and U14695 (N_14695,N_13843,N_13571);
nand U14696 (N_14696,N_13496,N_13421);
nand U14697 (N_14697,N_13962,N_13691);
nand U14698 (N_14698,N_13633,N_13403);
nand U14699 (N_14699,N_13826,N_13392);
nand U14700 (N_14700,N_13336,N_13283);
or U14701 (N_14701,N_13414,N_13322);
or U14702 (N_14702,N_13802,N_13957);
xnor U14703 (N_14703,N_13447,N_13846);
and U14704 (N_14704,N_13907,N_13587);
and U14705 (N_14705,N_13230,N_13029);
and U14706 (N_14706,N_13287,N_13329);
or U14707 (N_14707,N_13364,N_13146);
nor U14708 (N_14708,N_13533,N_13652);
or U14709 (N_14709,N_13072,N_13452);
or U14710 (N_14710,N_13593,N_13865);
xor U14711 (N_14711,N_13459,N_13396);
nor U14712 (N_14712,N_13961,N_13697);
xor U14713 (N_14713,N_13267,N_13246);
and U14714 (N_14714,N_13723,N_13803);
or U14715 (N_14715,N_13720,N_13009);
nand U14716 (N_14716,N_13238,N_13183);
nor U14717 (N_14717,N_13425,N_13046);
xnor U14718 (N_14718,N_13095,N_13027);
xor U14719 (N_14719,N_13406,N_13089);
xnor U14720 (N_14720,N_13502,N_13547);
or U14721 (N_14721,N_13658,N_13010);
or U14722 (N_14722,N_13431,N_13592);
and U14723 (N_14723,N_13063,N_13338);
or U14724 (N_14724,N_13572,N_13287);
nand U14725 (N_14725,N_13443,N_13782);
or U14726 (N_14726,N_13069,N_13732);
and U14727 (N_14727,N_13743,N_13820);
nand U14728 (N_14728,N_13656,N_13154);
nand U14729 (N_14729,N_13944,N_13460);
or U14730 (N_14730,N_13691,N_13643);
or U14731 (N_14731,N_13939,N_13073);
xnor U14732 (N_14732,N_13188,N_13853);
nor U14733 (N_14733,N_13854,N_13935);
or U14734 (N_14734,N_13916,N_13353);
and U14735 (N_14735,N_13405,N_13945);
or U14736 (N_14736,N_13633,N_13380);
xor U14737 (N_14737,N_13189,N_13464);
nand U14738 (N_14738,N_13695,N_13499);
nand U14739 (N_14739,N_13137,N_13296);
and U14740 (N_14740,N_13562,N_13839);
xnor U14741 (N_14741,N_13007,N_13333);
or U14742 (N_14742,N_13028,N_13857);
nand U14743 (N_14743,N_13462,N_13944);
and U14744 (N_14744,N_13580,N_13730);
nor U14745 (N_14745,N_13651,N_13058);
nor U14746 (N_14746,N_13875,N_13230);
nor U14747 (N_14747,N_13260,N_13465);
nor U14748 (N_14748,N_13808,N_13025);
and U14749 (N_14749,N_13773,N_13818);
nor U14750 (N_14750,N_13898,N_13589);
and U14751 (N_14751,N_13517,N_13768);
and U14752 (N_14752,N_13642,N_13425);
nor U14753 (N_14753,N_13175,N_13662);
nor U14754 (N_14754,N_13906,N_13014);
xnor U14755 (N_14755,N_13553,N_13323);
xnor U14756 (N_14756,N_13948,N_13675);
or U14757 (N_14757,N_13534,N_13420);
and U14758 (N_14758,N_13231,N_13947);
or U14759 (N_14759,N_13827,N_13672);
and U14760 (N_14760,N_13847,N_13999);
and U14761 (N_14761,N_13750,N_13995);
or U14762 (N_14762,N_13034,N_13980);
nand U14763 (N_14763,N_13095,N_13422);
nand U14764 (N_14764,N_13216,N_13768);
or U14765 (N_14765,N_13140,N_13940);
or U14766 (N_14766,N_13259,N_13877);
or U14767 (N_14767,N_13236,N_13834);
xnor U14768 (N_14768,N_13106,N_13299);
nor U14769 (N_14769,N_13977,N_13180);
nand U14770 (N_14770,N_13488,N_13985);
xnor U14771 (N_14771,N_13709,N_13716);
and U14772 (N_14772,N_13135,N_13869);
or U14773 (N_14773,N_13931,N_13277);
nor U14774 (N_14774,N_13805,N_13027);
nand U14775 (N_14775,N_13358,N_13588);
nand U14776 (N_14776,N_13456,N_13950);
nor U14777 (N_14777,N_13251,N_13887);
or U14778 (N_14778,N_13314,N_13357);
nand U14779 (N_14779,N_13911,N_13450);
xnor U14780 (N_14780,N_13892,N_13791);
or U14781 (N_14781,N_13412,N_13185);
nand U14782 (N_14782,N_13386,N_13793);
xnor U14783 (N_14783,N_13273,N_13703);
or U14784 (N_14784,N_13448,N_13499);
nand U14785 (N_14785,N_13053,N_13440);
or U14786 (N_14786,N_13744,N_13902);
xnor U14787 (N_14787,N_13931,N_13748);
nor U14788 (N_14788,N_13052,N_13106);
nand U14789 (N_14789,N_13351,N_13751);
and U14790 (N_14790,N_13453,N_13770);
or U14791 (N_14791,N_13664,N_13671);
nand U14792 (N_14792,N_13497,N_13191);
and U14793 (N_14793,N_13531,N_13310);
nor U14794 (N_14794,N_13420,N_13549);
xnor U14795 (N_14795,N_13493,N_13498);
or U14796 (N_14796,N_13612,N_13959);
xor U14797 (N_14797,N_13209,N_13347);
xor U14798 (N_14798,N_13665,N_13166);
nand U14799 (N_14799,N_13795,N_13824);
nand U14800 (N_14800,N_13543,N_13875);
and U14801 (N_14801,N_13589,N_13333);
and U14802 (N_14802,N_13843,N_13355);
xnor U14803 (N_14803,N_13984,N_13548);
and U14804 (N_14804,N_13214,N_13179);
and U14805 (N_14805,N_13312,N_13977);
and U14806 (N_14806,N_13602,N_13951);
nand U14807 (N_14807,N_13501,N_13664);
or U14808 (N_14808,N_13276,N_13426);
and U14809 (N_14809,N_13875,N_13318);
nand U14810 (N_14810,N_13376,N_13999);
nor U14811 (N_14811,N_13042,N_13445);
nor U14812 (N_14812,N_13482,N_13950);
and U14813 (N_14813,N_13249,N_13930);
or U14814 (N_14814,N_13119,N_13804);
or U14815 (N_14815,N_13824,N_13431);
or U14816 (N_14816,N_13604,N_13917);
nor U14817 (N_14817,N_13235,N_13653);
xor U14818 (N_14818,N_13698,N_13226);
nand U14819 (N_14819,N_13726,N_13029);
or U14820 (N_14820,N_13102,N_13854);
xor U14821 (N_14821,N_13004,N_13363);
or U14822 (N_14822,N_13565,N_13129);
xnor U14823 (N_14823,N_13810,N_13185);
and U14824 (N_14824,N_13662,N_13939);
and U14825 (N_14825,N_13275,N_13851);
nor U14826 (N_14826,N_13335,N_13037);
and U14827 (N_14827,N_13077,N_13493);
xnor U14828 (N_14828,N_13041,N_13477);
or U14829 (N_14829,N_13074,N_13959);
xnor U14830 (N_14830,N_13286,N_13969);
nor U14831 (N_14831,N_13891,N_13504);
and U14832 (N_14832,N_13067,N_13082);
nor U14833 (N_14833,N_13840,N_13982);
nand U14834 (N_14834,N_13799,N_13020);
and U14835 (N_14835,N_13172,N_13267);
nand U14836 (N_14836,N_13734,N_13883);
and U14837 (N_14837,N_13230,N_13401);
nand U14838 (N_14838,N_13031,N_13537);
nor U14839 (N_14839,N_13312,N_13328);
nor U14840 (N_14840,N_13227,N_13189);
and U14841 (N_14841,N_13405,N_13300);
xnor U14842 (N_14842,N_13898,N_13011);
or U14843 (N_14843,N_13109,N_13045);
nor U14844 (N_14844,N_13131,N_13929);
or U14845 (N_14845,N_13473,N_13688);
xor U14846 (N_14846,N_13421,N_13320);
xor U14847 (N_14847,N_13768,N_13904);
nand U14848 (N_14848,N_13094,N_13731);
nand U14849 (N_14849,N_13252,N_13191);
nand U14850 (N_14850,N_13701,N_13138);
nor U14851 (N_14851,N_13644,N_13052);
nand U14852 (N_14852,N_13513,N_13567);
nor U14853 (N_14853,N_13519,N_13127);
and U14854 (N_14854,N_13249,N_13354);
xor U14855 (N_14855,N_13004,N_13014);
and U14856 (N_14856,N_13589,N_13293);
nand U14857 (N_14857,N_13059,N_13718);
or U14858 (N_14858,N_13689,N_13215);
nor U14859 (N_14859,N_13682,N_13559);
nor U14860 (N_14860,N_13585,N_13129);
nand U14861 (N_14861,N_13331,N_13156);
xor U14862 (N_14862,N_13861,N_13169);
and U14863 (N_14863,N_13930,N_13713);
xor U14864 (N_14864,N_13802,N_13164);
and U14865 (N_14865,N_13377,N_13640);
or U14866 (N_14866,N_13698,N_13665);
nand U14867 (N_14867,N_13563,N_13628);
nor U14868 (N_14868,N_13229,N_13697);
or U14869 (N_14869,N_13486,N_13710);
or U14870 (N_14870,N_13587,N_13664);
and U14871 (N_14871,N_13630,N_13928);
or U14872 (N_14872,N_13414,N_13776);
nand U14873 (N_14873,N_13664,N_13456);
nor U14874 (N_14874,N_13598,N_13799);
nand U14875 (N_14875,N_13514,N_13874);
nand U14876 (N_14876,N_13379,N_13193);
or U14877 (N_14877,N_13192,N_13143);
nand U14878 (N_14878,N_13647,N_13924);
and U14879 (N_14879,N_13314,N_13952);
and U14880 (N_14880,N_13843,N_13254);
xor U14881 (N_14881,N_13732,N_13200);
xor U14882 (N_14882,N_13305,N_13297);
and U14883 (N_14883,N_13592,N_13336);
xnor U14884 (N_14884,N_13812,N_13259);
nor U14885 (N_14885,N_13402,N_13453);
or U14886 (N_14886,N_13900,N_13552);
and U14887 (N_14887,N_13169,N_13305);
xnor U14888 (N_14888,N_13622,N_13257);
nor U14889 (N_14889,N_13865,N_13690);
nand U14890 (N_14890,N_13876,N_13357);
or U14891 (N_14891,N_13803,N_13490);
nand U14892 (N_14892,N_13327,N_13434);
nor U14893 (N_14893,N_13281,N_13032);
and U14894 (N_14894,N_13402,N_13187);
xor U14895 (N_14895,N_13650,N_13814);
nand U14896 (N_14896,N_13729,N_13249);
nor U14897 (N_14897,N_13978,N_13279);
nand U14898 (N_14898,N_13799,N_13858);
xnor U14899 (N_14899,N_13312,N_13025);
xor U14900 (N_14900,N_13141,N_13086);
nor U14901 (N_14901,N_13707,N_13791);
nand U14902 (N_14902,N_13081,N_13285);
nor U14903 (N_14903,N_13657,N_13222);
xor U14904 (N_14904,N_13079,N_13594);
or U14905 (N_14905,N_13990,N_13465);
nor U14906 (N_14906,N_13832,N_13595);
or U14907 (N_14907,N_13893,N_13472);
nand U14908 (N_14908,N_13468,N_13630);
nand U14909 (N_14909,N_13188,N_13527);
xor U14910 (N_14910,N_13730,N_13214);
and U14911 (N_14911,N_13508,N_13414);
xor U14912 (N_14912,N_13142,N_13884);
or U14913 (N_14913,N_13294,N_13631);
xor U14914 (N_14914,N_13669,N_13756);
nand U14915 (N_14915,N_13817,N_13658);
and U14916 (N_14916,N_13765,N_13510);
xnor U14917 (N_14917,N_13046,N_13861);
and U14918 (N_14918,N_13437,N_13439);
and U14919 (N_14919,N_13929,N_13335);
and U14920 (N_14920,N_13323,N_13471);
xnor U14921 (N_14921,N_13677,N_13511);
nand U14922 (N_14922,N_13367,N_13042);
and U14923 (N_14923,N_13470,N_13889);
or U14924 (N_14924,N_13399,N_13986);
or U14925 (N_14925,N_13654,N_13784);
or U14926 (N_14926,N_13186,N_13924);
xor U14927 (N_14927,N_13679,N_13051);
and U14928 (N_14928,N_13735,N_13764);
nor U14929 (N_14929,N_13978,N_13451);
nor U14930 (N_14930,N_13645,N_13991);
nand U14931 (N_14931,N_13260,N_13163);
nor U14932 (N_14932,N_13479,N_13270);
and U14933 (N_14933,N_13013,N_13458);
nand U14934 (N_14934,N_13899,N_13409);
and U14935 (N_14935,N_13334,N_13587);
and U14936 (N_14936,N_13661,N_13939);
or U14937 (N_14937,N_13314,N_13900);
nand U14938 (N_14938,N_13267,N_13382);
nand U14939 (N_14939,N_13863,N_13832);
xor U14940 (N_14940,N_13444,N_13718);
or U14941 (N_14941,N_13847,N_13454);
and U14942 (N_14942,N_13824,N_13455);
xnor U14943 (N_14943,N_13749,N_13442);
nor U14944 (N_14944,N_13621,N_13049);
or U14945 (N_14945,N_13863,N_13606);
or U14946 (N_14946,N_13207,N_13459);
nand U14947 (N_14947,N_13504,N_13697);
and U14948 (N_14948,N_13164,N_13957);
or U14949 (N_14949,N_13734,N_13610);
nor U14950 (N_14950,N_13294,N_13893);
and U14951 (N_14951,N_13774,N_13186);
nand U14952 (N_14952,N_13916,N_13717);
and U14953 (N_14953,N_13210,N_13049);
xnor U14954 (N_14954,N_13118,N_13583);
and U14955 (N_14955,N_13776,N_13816);
nand U14956 (N_14956,N_13319,N_13820);
nor U14957 (N_14957,N_13309,N_13120);
or U14958 (N_14958,N_13123,N_13899);
or U14959 (N_14959,N_13728,N_13211);
and U14960 (N_14960,N_13780,N_13855);
xnor U14961 (N_14961,N_13300,N_13590);
or U14962 (N_14962,N_13333,N_13489);
xnor U14963 (N_14963,N_13709,N_13614);
nor U14964 (N_14964,N_13100,N_13400);
xnor U14965 (N_14965,N_13256,N_13812);
nand U14966 (N_14966,N_13816,N_13942);
and U14967 (N_14967,N_13984,N_13999);
nand U14968 (N_14968,N_13935,N_13909);
nand U14969 (N_14969,N_13601,N_13864);
or U14970 (N_14970,N_13158,N_13147);
and U14971 (N_14971,N_13167,N_13349);
nand U14972 (N_14972,N_13769,N_13619);
and U14973 (N_14973,N_13705,N_13163);
and U14974 (N_14974,N_13027,N_13655);
nand U14975 (N_14975,N_13741,N_13610);
or U14976 (N_14976,N_13170,N_13302);
and U14977 (N_14977,N_13308,N_13932);
nand U14978 (N_14978,N_13445,N_13747);
xor U14979 (N_14979,N_13785,N_13079);
xor U14980 (N_14980,N_13102,N_13409);
xor U14981 (N_14981,N_13879,N_13008);
and U14982 (N_14982,N_13097,N_13982);
nor U14983 (N_14983,N_13907,N_13174);
xnor U14984 (N_14984,N_13763,N_13543);
nor U14985 (N_14985,N_13284,N_13212);
or U14986 (N_14986,N_13290,N_13440);
xnor U14987 (N_14987,N_13403,N_13772);
and U14988 (N_14988,N_13178,N_13650);
nor U14989 (N_14989,N_13685,N_13107);
and U14990 (N_14990,N_13504,N_13860);
xor U14991 (N_14991,N_13048,N_13325);
xor U14992 (N_14992,N_13929,N_13738);
nor U14993 (N_14993,N_13137,N_13547);
xor U14994 (N_14994,N_13043,N_13220);
or U14995 (N_14995,N_13868,N_13670);
nand U14996 (N_14996,N_13103,N_13789);
nand U14997 (N_14997,N_13735,N_13253);
and U14998 (N_14998,N_13478,N_13969);
or U14999 (N_14999,N_13226,N_13232);
and U15000 (N_15000,N_14698,N_14554);
nand U15001 (N_15001,N_14732,N_14865);
xor U15002 (N_15002,N_14248,N_14617);
and U15003 (N_15003,N_14590,N_14498);
and U15004 (N_15004,N_14052,N_14273);
and U15005 (N_15005,N_14810,N_14583);
and U15006 (N_15006,N_14020,N_14943);
and U15007 (N_15007,N_14392,N_14568);
or U15008 (N_15008,N_14644,N_14992);
nand U15009 (N_15009,N_14356,N_14038);
and U15010 (N_15010,N_14632,N_14671);
and U15011 (N_15011,N_14885,N_14205);
nor U15012 (N_15012,N_14308,N_14315);
or U15013 (N_15013,N_14913,N_14677);
and U15014 (N_15014,N_14218,N_14477);
or U15015 (N_15015,N_14789,N_14040);
or U15016 (N_15016,N_14719,N_14480);
or U15017 (N_15017,N_14488,N_14512);
or U15018 (N_15018,N_14202,N_14853);
and U15019 (N_15019,N_14075,N_14999);
and U15020 (N_15020,N_14118,N_14405);
nand U15021 (N_15021,N_14960,N_14263);
or U15022 (N_15022,N_14080,N_14550);
nor U15023 (N_15023,N_14884,N_14760);
or U15024 (N_15024,N_14807,N_14949);
nor U15025 (N_15025,N_14422,N_14186);
nand U15026 (N_15026,N_14267,N_14069);
xor U15027 (N_15027,N_14328,N_14923);
xor U15028 (N_15028,N_14428,N_14362);
or U15029 (N_15029,N_14514,N_14784);
nand U15030 (N_15030,N_14723,N_14805);
nor U15031 (N_15031,N_14402,N_14822);
nand U15032 (N_15032,N_14003,N_14433);
and U15033 (N_15033,N_14228,N_14821);
and U15034 (N_15034,N_14570,N_14011);
and U15035 (N_15035,N_14833,N_14114);
or U15036 (N_15036,N_14601,N_14458);
xor U15037 (N_15037,N_14142,N_14256);
or U15038 (N_15038,N_14781,N_14758);
nand U15039 (N_15039,N_14503,N_14301);
nor U15040 (N_15040,N_14354,N_14643);
nand U15041 (N_15041,N_14928,N_14337);
nor U15042 (N_15042,N_14975,N_14146);
or U15043 (N_15043,N_14450,N_14072);
and U15044 (N_15044,N_14286,N_14318);
xor U15045 (N_15045,N_14430,N_14795);
nor U15046 (N_15046,N_14538,N_14193);
or U15047 (N_15047,N_14857,N_14324);
and U15048 (N_15048,N_14360,N_14639);
xnor U15049 (N_15049,N_14084,N_14908);
nor U15050 (N_15050,N_14579,N_14887);
and U15051 (N_15051,N_14692,N_14086);
or U15052 (N_15052,N_14194,N_14492);
and U15053 (N_15053,N_14123,N_14007);
xnor U15054 (N_15054,N_14203,N_14872);
and U15055 (N_15055,N_14525,N_14546);
nand U15056 (N_15056,N_14591,N_14325);
or U15057 (N_15057,N_14729,N_14759);
nand U15058 (N_15058,N_14598,N_14547);
or U15059 (N_15059,N_14945,N_14612);
or U15060 (N_15060,N_14953,N_14956);
or U15061 (N_15061,N_14342,N_14957);
and U15062 (N_15062,N_14024,N_14100);
nor U15063 (N_15063,N_14766,N_14183);
or U15064 (N_15064,N_14469,N_14066);
and U15065 (N_15065,N_14264,N_14606);
or U15066 (N_15066,N_14721,N_14169);
or U15067 (N_15067,N_14965,N_14855);
and U15068 (N_15068,N_14646,N_14605);
xor U15069 (N_15069,N_14834,N_14168);
nand U15070 (N_15070,N_14609,N_14633);
nand U15071 (N_15071,N_14571,N_14708);
nor U15072 (N_15072,N_14389,N_14743);
or U15073 (N_15073,N_14312,N_14128);
nand U15074 (N_15074,N_14474,N_14587);
or U15075 (N_15075,N_14777,N_14504);
and U15076 (N_15076,N_14010,N_14476);
and U15077 (N_15077,N_14836,N_14030);
nand U15078 (N_15078,N_14636,N_14297);
nor U15079 (N_15079,N_14303,N_14115);
nand U15080 (N_15080,N_14838,N_14152);
or U15081 (N_15081,N_14008,N_14877);
xor U15082 (N_15082,N_14326,N_14154);
and U15083 (N_15083,N_14544,N_14515);
xnor U15084 (N_15084,N_14377,N_14062);
or U15085 (N_15085,N_14645,N_14306);
or U15086 (N_15086,N_14958,N_14158);
nor U15087 (N_15087,N_14627,N_14156);
or U15088 (N_15088,N_14981,N_14418);
xor U15089 (N_15089,N_14811,N_14473);
nand U15090 (N_15090,N_14533,N_14816);
and U15091 (N_15091,N_14915,N_14406);
xnor U15092 (N_15092,N_14738,N_14762);
xor U15093 (N_15093,N_14924,N_14260);
nand U15094 (N_15094,N_14638,N_14272);
nor U15095 (N_15095,N_14025,N_14597);
nor U15096 (N_15096,N_14883,N_14988);
nand U15097 (N_15097,N_14974,N_14148);
nor U15098 (N_15098,N_14283,N_14447);
xnor U15099 (N_15099,N_14284,N_14268);
nor U15100 (N_15100,N_14888,N_14001);
and U15101 (N_15101,N_14790,N_14112);
or U15102 (N_15102,N_14680,N_14387);
nor U15103 (N_15103,N_14959,N_14728);
xnor U15104 (N_15104,N_14175,N_14464);
and U15105 (N_15105,N_14942,N_14061);
xor U15106 (N_15106,N_14954,N_14352);
or U15107 (N_15107,N_14179,N_14341);
nand U15108 (N_15108,N_14806,N_14220);
nand U15109 (N_15109,N_14564,N_14290);
xnor U15110 (N_15110,N_14056,N_14427);
or U15111 (N_15111,N_14879,N_14407);
or U15112 (N_15112,N_14487,N_14714);
nor U15113 (N_15113,N_14497,N_14215);
and U15114 (N_15114,N_14232,N_14028);
or U15115 (N_15115,N_14794,N_14217);
nand U15116 (N_15116,N_14854,N_14425);
nand U15117 (N_15117,N_14894,N_14471);
nand U15118 (N_15118,N_14358,N_14771);
and U15119 (N_15119,N_14350,N_14511);
nand U15120 (N_15120,N_14819,N_14847);
nand U15121 (N_15121,N_14505,N_14578);
and U15122 (N_15122,N_14964,N_14426);
nor U15123 (N_15123,N_14886,N_14088);
xor U15124 (N_15124,N_14882,N_14907);
nor U15125 (N_15125,N_14850,N_14249);
nor U15126 (N_15126,N_14460,N_14357);
nor U15127 (N_15127,N_14394,N_14033);
nor U15128 (N_15128,N_14371,N_14468);
nor U15129 (N_15129,N_14799,N_14167);
and U15130 (N_15130,N_14305,N_14434);
and U15131 (N_15131,N_14933,N_14300);
and U15132 (N_15132,N_14802,N_14779);
xor U15133 (N_15133,N_14935,N_14594);
nand U15134 (N_15134,N_14071,N_14094);
and U15135 (N_15135,N_14764,N_14919);
nand U15136 (N_15136,N_14237,N_14610);
xnor U15137 (N_15137,N_14529,N_14153);
nor U15138 (N_15138,N_14369,N_14439);
or U15139 (N_15139,N_14979,N_14615);
xnor U15140 (N_15140,N_14563,N_14769);
or U15141 (N_15141,N_14496,N_14410);
nand U15142 (N_15142,N_14087,N_14629);
nor U15143 (N_15143,N_14293,N_14348);
or U15144 (N_15144,N_14296,N_14330);
and U15145 (N_15145,N_14673,N_14077);
or U15146 (N_15146,N_14095,N_14310);
nor U15147 (N_15147,N_14800,N_14791);
nand U15148 (N_15148,N_14448,N_14274);
nor U15149 (N_15149,N_14495,N_14876);
nor U15150 (N_15150,N_14182,N_14345);
nor U15151 (N_15151,N_14262,N_14682);
nand U15152 (N_15152,N_14436,N_14659);
nor U15153 (N_15153,N_14285,N_14572);
and U15154 (N_15154,N_14212,N_14842);
and U15155 (N_15155,N_14768,N_14299);
and U15156 (N_15156,N_14889,N_14927);
and U15157 (N_15157,N_14607,N_14839);
nand U15158 (N_15158,N_14619,N_14720);
nor U15159 (N_15159,N_14171,N_14419);
or U15160 (N_15160,N_14699,N_14366);
nand U15161 (N_15161,N_14437,N_14491);
or U15162 (N_15162,N_14574,N_14302);
nor U15163 (N_15163,N_14722,N_14778);
and U15164 (N_15164,N_14107,N_14870);
and U15165 (N_15165,N_14524,N_14133);
and U15166 (N_15166,N_14431,N_14294);
nand U15167 (N_15167,N_14081,N_14320);
or U15168 (N_15168,N_14670,N_14143);
and U15169 (N_15169,N_14047,N_14014);
nor U15170 (N_15170,N_14841,N_14986);
xnor U15171 (N_15171,N_14364,N_14197);
and U15172 (N_15172,N_14519,N_14552);
nand U15173 (N_15173,N_14036,N_14104);
and U15174 (N_15174,N_14400,N_14798);
xnor U15175 (N_15175,N_14950,N_14322);
nor U15176 (N_15176,N_14507,N_14185);
xor U15177 (N_15177,N_14292,N_14832);
or U15178 (N_15178,N_14741,N_14067);
or U15179 (N_15179,N_14740,N_14313);
nand U15180 (N_15180,N_14097,N_14749);
nand U15181 (N_15181,N_14211,N_14716);
and U15182 (N_15182,N_14948,N_14204);
xnor U15183 (N_15183,N_14901,N_14125);
and U15184 (N_15184,N_14868,N_14737);
xnor U15185 (N_15185,N_14730,N_14650);
and U15186 (N_15186,N_14751,N_14560);
or U15187 (N_15187,N_14027,N_14170);
nand U15188 (N_15188,N_14291,N_14098);
or U15189 (N_15189,N_14208,N_14706);
and U15190 (N_15190,N_14139,N_14969);
and U15191 (N_15191,N_14481,N_14184);
and U15192 (N_15192,N_14614,N_14365);
nand U15193 (N_15193,N_14690,N_14165);
xor U15194 (N_15194,N_14982,N_14166);
nand U15195 (N_15195,N_14178,N_14825);
nand U15196 (N_15196,N_14526,N_14412);
nor U15197 (N_15197,N_14648,N_14335);
or U15198 (N_15198,N_14089,N_14952);
or U15199 (N_15199,N_14135,N_14903);
xor U15200 (N_15200,N_14508,N_14846);
or U15201 (N_15201,N_14177,N_14029);
nand U15202 (N_15202,N_14382,N_14788);
or U15203 (N_15203,N_14881,N_14987);
or U15204 (N_15204,N_14454,N_14852);
xor U15205 (N_15205,N_14219,N_14984);
nand U15206 (N_15206,N_14622,N_14667);
or U15207 (N_15207,N_14102,N_14830);
and U15208 (N_15208,N_14336,N_14864);
and U15209 (N_15209,N_14332,N_14835);
nand U15210 (N_15210,N_14349,N_14596);
xor U15211 (N_15211,N_14711,N_14809);
nor U15212 (N_15212,N_14748,N_14843);
and U15213 (N_15213,N_14936,N_14654);
and U15214 (N_15214,N_14528,N_14628);
and U15215 (N_15215,N_14656,N_14672);
xor U15216 (N_15216,N_14813,N_14998);
and U15217 (N_15217,N_14727,N_14941);
nand U15218 (N_15218,N_14517,N_14259);
and U15219 (N_15219,N_14584,N_14490);
and U15220 (N_15220,N_14224,N_14686);
nor U15221 (N_15221,N_14559,N_14993);
nor U15222 (N_15222,N_14398,N_14994);
nand U15223 (N_15223,N_14049,N_14931);
nand U15224 (N_15224,N_14467,N_14851);
nor U15225 (N_15225,N_14192,N_14314);
nor U15226 (N_15226,N_14386,N_14618);
or U15227 (N_15227,N_14149,N_14113);
nor U15228 (N_15228,N_14420,N_14076);
nor U15229 (N_15229,N_14150,N_14017);
xnor U15230 (N_15230,N_14586,N_14929);
xnor U15231 (N_15231,N_14421,N_14122);
or U15232 (N_15232,N_14316,N_14724);
or U15233 (N_15233,N_14311,N_14642);
or U15234 (N_15234,N_14347,N_14739);
nand U15235 (N_15235,N_14926,N_14675);
or U15236 (N_15236,N_14461,N_14449);
nand U15237 (N_15237,N_14108,N_14577);
xnor U15238 (N_15238,N_14199,N_14531);
nand U15239 (N_15239,N_14668,N_14018);
and U15240 (N_15240,N_14712,N_14361);
or U15241 (N_15241,N_14780,N_14718);
or U15242 (N_15242,N_14890,N_14472);
nand U15243 (N_15243,N_14190,N_14101);
nand U15244 (N_15244,N_14270,N_14961);
or U15245 (N_15245,N_14390,N_14506);
nor U15246 (N_15246,N_14625,N_14092);
nand U15247 (N_15247,N_14438,N_14042);
and U15248 (N_15248,N_14022,N_14000);
nand U15249 (N_15249,N_14276,N_14207);
nor U15250 (N_15250,N_14717,N_14174);
xor U15251 (N_15251,N_14824,N_14026);
nor U15252 (N_15252,N_14770,N_14991);
xor U15253 (N_15253,N_14374,N_14611);
xor U15254 (N_15254,N_14580,N_14944);
and U15255 (N_15255,N_14837,N_14653);
nand U15256 (N_15256,N_14378,N_14391);
xnor U15257 (N_15257,N_14823,N_14288);
nor U15258 (N_15258,N_14683,N_14188);
and U15259 (N_15259,N_14106,N_14917);
and U15260 (N_15260,N_14130,N_14539);
nor U15261 (N_15261,N_14602,N_14209);
nand U15262 (N_15262,N_14589,N_14340);
and U15263 (N_15263,N_14695,N_14678);
nor U15264 (N_15264,N_14814,N_14637);
and U15265 (N_15265,N_14869,N_14446);
and U15266 (N_15266,N_14747,N_14765);
nand U15267 (N_15267,N_14657,N_14085);
xnor U15268 (N_15268,N_14750,N_14697);
and U15269 (N_15269,N_14016,N_14962);
xor U15270 (N_15270,N_14616,N_14878);
and U15271 (N_15271,N_14973,N_14367);
and U15272 (N_15272,N_14375,N_14767);
nor U15273 (N_15273,N_14109,N_14415);
nand U15274 (N_15274,N_14408,N_14527);
nand U15275 (N_15275,N_14327,N_14479);
and U15276 (N_15276,N_14261,N_14754);
or U15277 (N_15277,N_14746,N_14756);
or U15278 (N_15278,N_14275,N_14015);
xor U15279 (N_15279,N_14796,N_14561);
or U15280 (N_15280,N_14989,N_14745);
nor U15281 (N_15281,N_14862,N_14626);
xor U15282 (N_15282,N_14424,N_14702);
or U15283 (N_15283,N_14532,N_14588);
and U15284 (N_15284,N_14021,N_14689);
nor U15285 (N_15285,N_14909,N_14280);
xor U15286 (N_15286,N_14551,N_14793);
xnor U15287 (N_15287,N_14782,N_14801);
xor U15288 (N_15288,N_14082,N_14399);
nor U15289 (N_15289,N_14726,N_14457);
or U15290 (N_15290,N_14828,N_14681);
nor U15291 (N_15291,N_14817,N_14455);
nor U15292 (N_15292,N_14501,N_14581);
or U15293 (N_15293,N_14053,N_14921);
and U15294 (N_15294,N_14701,N_14110);
xor U15295 (N_15295,N_14009,N_14569);
nor U15296 (N_15296,N_14573,N_14196);
nor U15297 (N_15297,N_14829,N_14006);
xor U15298 (N_15298,N_14388,N_14858);
xor U15299 (N_15299,N_14640,N_14844);
and U15300 (N_15300,N_14966,N_14096);
nand U15301 (N_15301,N_14200,N_14592);
and U15302 (N_15302,N_14787,N_14246);
nand U15303 (N_15303,N_14860,N_14485);
nand U15304 (N_15304,N_14126,N_14383);
or U15305 (N_15305,N_14411,N_14304);
and U15306 (N_15306,N_14381,N_14057);
and U15307 (N_15307,N_14258,N_14013);
nor U15308 (N_15308,N_14380,N_14910);
or U15309 (N_15309,N_14353,N_14213);
nand U15310 (N_15310,N_14269,N_14867);
or U15311 (N_15311,N_14666,N_14379);
nand U15312 (N_15312,N_14694,N_14932);
and U15313 (N_15313,N_14500,N_14906);
and U15314 (N_15314,N_14334,N_14997);
or U15315 (N_15315,N_14278,N_14757);
and U15316 (N_15316,N_14499,N_14543);
nor U15317 (N_15317,N_14774,N_14621);
or U15318 (N_15318,N_14189,N_14555);
and U15319 (N_15319,N_14651,N_14920);
xor U15320 (N_15320,N_14938,N_14922);
nor U15321 (N_15321,N_14631,N_14660);
and U15322 (N_15322,N_14875,N_14105);
nor U15323 (N_15323,N_14039,N_14652);
xor U15324 (N_15324,N_14250,N_14818);
xor U15325 (N_15325,N_14676,N_14783);
or U15326 (N_15326,N_14873,N_14159);
xnor U15327 (N_15327,N_14240,N_14265);
xor U15328 (N_15328,N_14462,N_14603);
xnor U15329 (N_15329,N_14404,N_14140);
and U15330 (N_15330,N_14566,N_14043);
or U15331 (N_15331,N_14247,N_14535);
nor U15332 (N_15332,N_14227,N_14074);
nand U15333 (N_15333,N_14339,N_14343);
or U15334 (N_15334,N_14634,N_14079);
and U15335 (N_15335,N_14073,N_14704);
xor U15336 (N_15336,N_14160,N_14441);
nor U15337 (N_15337,N_14871,N_14731);
or U15338 (N_15338,N_14236,N_14911);
nor U15339 (N_15339,N_14214,N_14620);
nor U15340 (N_15340,N_14946,N_14482);
xnor U15341 (N_15341,N_14849,N_14661);
and U15342 (N_15342,N_14662,N_14895);
or U15343 (N_15343,N_14376,N_14968);
or U15344 (N_15344,N_14161,N_14164);
and U15345 (N_15345,N_14147,N_14937);
or U15346 (N_15346,N_14172,N_14393);
nand U15347 (N_15347,N_14144,N_14252);
xor U15348 (N_15348,N_14060,N_14930);
nor U15349 (N_15349,N_14912,N_14051);
nand U15350 (N_15350,N_14736,N_14363);
xnor U15351 (N_15351,N_14565,N_14241);
or U15352 (N_15352,N_14282,N_14733);
and U15353 (N_15353,N_14201,N_14647);
nand U15354 (N_15354,N_14516,N_14127);
or U15355 (N_15355,N_14744,N_14298);
xnor U15356 (N_15356,N_14576,N_14831);
or U15357 (N_15357,N_14845,N_14486);
nor U15358 (N_15358,N_14173,N_14198);
nor U15359 (N_15359,N_14874,N_14058);
nor U15360 (N_15360,N_14116,N_14509);
and U15361 (N_15361,N_14715,N_14048);
or U15362 (N_15362,N_14983,N_14608);
xnor U15363 (N_15363,N_14710,N_14230);
or U15364 (N_15364,N_14827,N_14245);
nand U15365 (N_15365,N_14502,N_14233);
xnor U15366 (N_15366,N_14368,N_14990);
or U15367 (N_15367,N_14483,N_14373);
nand U15368 (N_15368,N_14521,N_14808);
nor U15369 (N_15369,N_14812,N_14331);
and U15370 (N_15370,N_14763,N_14775);
and U15371 (N_15371,N_14856,N_14068);
xnor U15372 (N_15372,N_14333,N_14880);
and U15373 (N_15373,N_14896,N_14649);
and U15374 (N_15374,N_14493,N_14664);
xnor U15375 (N_15375,N_14254,N_14557);
xor U15376 (N_15376,N_14395,N_14141);
nand U15377 (N_15377,N_14687,N_14899);
xor U15378 (N_15378,N_14900,N_14396);
nand U15379 (N_15379,N_14226,N_14065);
nand U15380 (N_15380,N_14513,N_14279);
and U15381 (N_15381,N_14289,N_14815);
nor U15382 (N_15382,N_14083,N_14225);
nor U15383 (N_15383,N_14035,N_14002);
and U15384 (N_15384,N_14103,N_14707);
or U15385 (N_15385,N_14070,N_14776);
xnor U15386 (N_15386,N_14967,N_14195);
and U15387 (N_15387,N_14534,N_14826);
or U15388 (N_15388,N_14019,N_14124);
xnor U15389 (N_15389,N_14914,N_14893);
xor U15390 (N_15390,N_14281,N_14222);
xor U15391 (N_15391,N_14444,N_14307);
and U15392 (N_15392,N_14585,N_14239);
nor U15393 (N_15393,N_14537,N_14703);
nor U15394 (N_15394,N_14093,N_14925);
nor U15395 (N_15395,N_14545,N_14466);
or U15396 (N_15396,N_14445,N_14734);
nand U15397 (N_15397,N_14669,N_14266);
or U15398 (N_15398,N_14005,N_14530);
and U15399 (N_15399,N_14157,N_14897);
nand U15400 (N_15400,N_14820,N_14613);
and U15401 (N_15401,N_14655,N_14786);
nor U15402 (N_15402,N_14548,N_14995);
nor U15403 (N_15403,N_14976,N_14663);
nor U15404 (N_15404,N_14696,N_14055);
xor U15405 (N_15405,N_14023,N_14041);
xnor U15406 (N_15406,N_14091,N_14034);
xor U15407 (N_15407,N_14414,N_14134);
and U15408 (N_15408,N_14359,N_14323);
xnor U15409 (N_15409,N_14059,N_14977);
nand U15410 (N_15410,N_14489,N_14216);
nor U15411 (N_15411,N_14947,N_14432);
xor U15412 (N_15412,N_14321,N_14658);
nor U15413 (N_15413,N_14129,N_14234);
xnor U15414 (N_15414,N_14145,N_14012);
nor U15415 (N_15415,N_14980,N_14451);
or U15416 (N_15416,N_14484,N_14223);
nand U15417 (N_15417,N_14440,N_14423);
or U15418 (N_15418,N_14955,N_14562);
and U15419 (N_15419,N_14709,N_14970);
nand U15420 (N_15420,N_14044,N_14329);
or U15421 (N_15421,N_14522,N_14772);
or U15422 (N_15422,N_14892,N_14078);
xor U15423 (N_15423,N_14693,N_14401);
nand U15424 (N_15424,N_14181,N_14478);
nor U15425 (N_15425,N_14685,N_14317);
and U15426 (N_15426,N_14295,N_14996);
xnor U15427 (N_15427,N_14155,N_14804);
nor U15428 (N_15428,N_14409,N_14630);
xor U15429 (N_15429,N_14684,N_14385);
or U15430 (N_15430,N_14972,N_14985);
or U15431 (N_15431,N_14384,N_14163);
and U15432 (N_15432,N_14861,N_14567);
xor U15433 (N_15433,N_14742,N_14674);
xor U15434 (N_15434,N_14037,N_14131);
nand U15435 (N_15435,N_14735,N_14898);
or U15436 (N_15436,N_14797,N_14251);
or U15437 (N_15437,N_14064,N_14099);
xnor U15438 (N_15438,N_14176,N_14575);
and U15439 (N_15439,N_14238,N_14866);
nor U15440 (N_15440,N_14494,N_14713);
nor U15441 (N_15441,N_14475,N_14465);
nand U15442 (N_15442,N_14940,N_14624);
or U15443 (N_15443,N_14523,N_14046);
xnor U15444 (N_15444,N_14417,N_14755);
nor U15445 (N_15445,N_14257,N_14863);
and U15446 (N_15446,N_14370,N_14518);
nor U15447 (N_15447,N_14679,N_14120);
nand U15448 (N_15448,N_14542,N_14429);
nand U15449 (N_15449,N_14397,N_14346);
or U15450 (N_15450,N_14792,N_14229);
xor U15451 (N_15451,N_14403,N_14848);
nor U15452 (N_15452,N_14137,N_14582);
and U15453 (N_15453,N_14191,N_14136);
nor U15454 (N_15454,N_14221,N_14971);
and U15455 (N_15455,N_14623,N_14604);
xor U15456 (N_15456,N_14761,N_14558);
nand U15457 (N_15457,N_14442,N_14705);
nor U15458 (N_15458,N_14600,N_14470);
or U15459 (N_15459,N_14891,N_14978);
and U15460 (N_15460,N_14700,N_14840);
nand U15461 (N_15461,N_14355,N_14725);
xor U15462 (N_15462,N_14688,N_14413);
or U15463 (N_15463,N_14032,N_14916);
nor U15464 (N_15464,N_14351,N_14255);
xnor U15465 (N_15465,N_14242,N_14435);
or U15466 (N_15466,N_14753,N_14031);
nor U15467 (N_15467,N_14271,N_14540);
xor U15468 (N_15468,N_14372,N_14595);
and U15469 (N_15469,N_14556,N_14963);
and U15470 (N_15470,N_14162,N_14132);
or U15471 (N_15471,N_14338,N_14090);
or U15472 (N_15472,N_14045,N_14541);
nand U15473 (N_15473,N_14138,N_14416);
nand U15474 (N_15474,N_14459,N_14117);
or U15475 (N_15475,N_14244,N_14918);
and U15476 (N_15476,N_14453,N_14859);
or U15477 (N_15477,N_14277,N_14180);
nor U15478 (N_15478,N_14536,N_14773);
nor U15479 (N_15479,N_14635,N_14243);
or U15480 (N_15480,N_14054,N_14443);
and U15481 (N_15481,N_14553,N_14905);
nand U15482 (N_15482,N_14231,N_14951);
nand U15483 (N_15483,N_14111,N_14665);
and U15484 (N_15484,N_14641,N_14119);
nor U15485 (N_15485,N_14210,N_14463);
nor U15486 (N_15486,N_14549,N_14785);
or U15487 (N_15487,N_14691,N_14235);
nor U15488 (N_15488,N_14452,N_14063);
or U15489 (N_15489,N_14344,N_14510);
or U15490 (N_15490,N_14599,N_14151);
xor U15491 (N_15491,N_14287,N_14752);
nor U15492 (N_15492,N_14803,N_14309);
and U15493 (N_15493,N_14456,N_14187);
xnor U15494 (N_15494,N_14004,N_14050);
nand U15495 (N_15495,N_14319,N_14902);
or U15496 (N_15496,N_14593,N_14253);
and U15497 (N_15497,N_14206,N_14939);
and U15498 (N_15498,N_14934,N_14904);
and U15499 (N_15499,N_14520,N_14121);
and U15500 (N_15500,N_14534,N_14850);
nand U15501 (N_15501,N_14268,N_14718);
or U15502 (N_15502,N_14632,N_14766);
and U15503 (N_15503,N_14557,N_14253);
xor U15504 (N_15504,N_14645,N_14696);
xor U15505 (N_15505,N_14742,N_14691);
nand U15506 (N_15506,N_14074,N_14546);
xnor U15507 (N_15507,N_14685,N_14365);
xor U15508 (N_15508,N_14496,N_14559);
xor U15509 (N_15509,N_14579,N_14125);
nand U15510 (N_15510,N_14613,N_14346);
nand U15511 (N_15511,N_14927,N_14759);
xnor U15512 (N_15512,N_14940,N_14390);
xnor U15513 (N_15513,N_14787,N_14955);
nor U15514 (N_15514,N_14347,N_14773);
and U15515 (N_15515,N_14078,N_14839);
and U15516 (N_15516,N_14904,N_14754);
nor U15517 (N_15517,N_14032,N_14373);
nor U15518 (N_15518,N_14581,N_14798);
nand U15519 (N_15519,N_14915,N_14921);
nor U15520 (N_15520,N_14868,N_14887);
and U15521 (N_15521,N_14564,N_14971);
nand U15522 (N_15522,N_14522,N_14982);
xnor U15523 (N_15523,N_14224,N_14896);
or U15524 (N_15524,N_14142,N_14247);
or U15525 (N_15525,N_14455,N_14934);
or U15526 (N_15526,N_14411,N_14662);
xor U15527 (N_15527,N_14591,N_14304);
nor U15528 (N_15528,N_14148,N_14104);
and U15529 (N_15529,N_14603,N_14312);
nor U15530 (N_15530,N_14845,N_14900);
and U15531 (N_15531,N_14812,N_14039);
and U15532 (N_15532,N_14380,N_14641);
or U15533 (N_15533,N_14555,N_14121);
and U15534 (N_15534,N_14997,N_14390);
nor U15535 (N_15535,N_14556,N_14454);
nor U15536 (N_15536,N_14802,N_14016);
xor U15537 (N_15537,N_14905,N_14504);
xor U15538 (N_15538,N_14625,N_14112);
and U15539 (N_15539,N_14422,N_14263);
xor U15540 (N_15540,N_14960,N_14403);
xnor U15541 (N_15541,N_14340,N_14348);
nor U15542 (N_15542,N_14761,N_14708);
or U15543 (N_15543,N_14418,N_14874);
xnor U15544 (N_15544,N_14297,N_14878);
or U15545 (N_15545,N_14612,N_14277);
xnor U15546 (N_15546,N_14466,N_14862);
or U15547 (N_15547,N_14764,N_14902);
and U15548 (N_15548,N_14096,N_14694);
or U15549 (N_15549,N_14605,N_14743);
nor U15550 (N_15550,N_14364,N_14898);
xor U15551 (N_15551,N_14352,N_14841);
and U15552 (N_15552,N_14491,N_14326);
nor U15553 (N_15553,N_14197,N_14340);
xor U15554 (N_15554,N_14138,N_14047);
nor U15555 (N_15555,N_14108,N_14586);
nand U15556 (N_15556,N_14075,N_14984);
nand U15557 (N_15557,N_14524,N_14281);
xnor U15558 (N_15558,N_14482,N_14650);
nand U15559 (N_15559,N_14735,N_14003);
xnor U15560 (N_15560,N_14754,N_14017);
xnor U15561 (N_15561,N_14406,N_14685);
xor U15562 (N_15562,N_14209,N_14868);
and U15563 (N_15563,N_14234,N_14339);
nor U15564 (N_15564,N_14322,N_14173);
nand U15565 (N_15565,N_14486,N_14193);
nor U15566 (N_15566,N_14575,N_14219);
nand U15567 (N_15567,N_14244,N_14106);
or U15568 (N_15568,N_14259,N_14187);
or U15569 (N_15569,N_14514,N_14376);
and U15570 (N_15570,N_14634,N_14619);
and U15571 (N_15571,N_14948,N_14962);
and U15572 (N_15572,N_14621,N_14932);
and U15573 (N_15573,N_14651,N_14807);
or U15574 (N_15574,N_14262,N_14155);
nand U15575 (N_15575,N_14071,N_14933);
nor U15576 (N_15576,N_14873,N_14557);
nor U15577 (N_15577,N_14013,N_14012);
and U15578 (N_15578,N_14920,N_14474);
and U15579 (N_15579,N_14141,N_14883);
nor U15580 (N_15580,N_14785,N_14682);
or U15581 (N_15581,N_14017,N_14265);
and U15582 (N_15582,N_14132,N_14006);
xnor U15583 (N_15583,N_14713,N_14177);
nand U15584 (N_15584,N_14885,N_14636);
or U15585 (N_15585,N_14012,N_14204);
xor U15586 (N_15586,N_14993,N_14994);
and U15587 (N_15587,N_14145,N_14362);
nand U15588 (N_15588,N_14091,N_14108);
xor U15589 (N_15589,N_14262,N_14686);
and U15590 (N_15590,N_14443,N_14575);
or U15591 (N_15591,N_14841,N_14253);
and U15592 (N_15592,N_14747,N_14188);
nor U15593 (N_15593,N_14086,N_14365);
xor U15594 (N_15594,N_14053,N_14234);
and U15595 (N_15595,N_14744,N_14979);
and U15596 (N_15596,N_14043,N_14345);
xnor U15597 (N_15597,N_14878,N_14562);
xnor U15598 (N_15598,N_14279,N_14646);
and U15599 (N_15599,N_14895,N_14717);
or U15600 (N_15600,N_14178,N_14218);
xnor U15601 (N_15601,N_14687,N_14976);
xnor U15602 (N_15602,N_14301,N_14866);
xor U15603 (N_15603,N_14803,N_14011);
nor U15604 (N_15604,N_14431,N_14922);
nor U15605 (N_15605,N_14655,N_14170);
or U15606 (N_15606,N_14175,N_14966);
nor U15607 (N_15607,N_14611,N_14830);
xor U15608 (N_15608,N_14210,N_14318);
or U15609 (N_15609,N_14206,N_14848);
or U15610 (N_15610,N_14728,N_14895);
nand U15611 (N_15611,N_14749,N_14959);
and U15612 (N_15612,N_14219,N_14669);
nand U15613 (N_15613,N_14178,N_14705);
and U15614 (N_15614,N_14484,N_14737);
nand U15615 (N_15615,N_14945,N_14338);
and U15616 (N_15616,N_14277,N_14144);
or U15617 (N_15617,N_14179,N_14140);
and U15618 (N_15618,N_14638,N_14476);
and U15619 (N_15619,N_14187,N_14423);
nand U15620 (N_15620,N_14533,N_14564);
xor U15621 (N_15621,N_14990,N_14227);
nor U15622 (N_15622,N_14987,N_14904);
nand U15623 (N_15623,N_14252,N_14834);
or U15624 (N_15624,N_14166,N_14323);
xor U15625 (N_15625,N_14149,N_14865);
or U15626 (N_15626,N_14141,N_14029);
or U15627 (N_15627,N_14065,N_14975);
or U15628 (N_15628,N_14618,N_14244);
or U15629 (N_15629,N_14111,N_14459);
or U15630 (N_15630,N_14646,N_14162);
and U15631 (N_15631,N_14025,N_14370);
nor U15632 (N_15632,N_14798,N_14056);
nand U15633 (N_15633,N_14903,N_14727);
and U15634 (N_15634,N_14954,N_14722);
nor U15635 (N_15635,N_14522,N_14269);
xor U15636 (N_15636,N_14677,N_14393);
or U15637 (N_15637,N_14841,N_14030);
and U15638 (N_15638,N_14640,N_14794);
xor U15639 (N_15639,N_14617,N_14302);
and U15640 (N_15640,N_14178,N_14985);
or U15641 (N_15641,N_14436,N_14686);
nand U15642 (N_15642,N_14232,N_14476);
nor U15643 (N_15643,N_14736,N_14129);
nand U15644 (N_15644,N_14822,N_14081);
nor U15645 (N_15645,N_14552,N_14415);
and U15646 (N_15646,N_14128,N_14872);
and U15647 (N_15647,N_14962,N_14283);
xnor U15648 (N_15648,N_14336,N_14428);
and U15649 (N_15649,N_14097,N_14214);
xor U15650 (N_15650,N_14783,N_14374);
and U15651 (N_15651,N_14874,N_14557);
xor U15652 (N_15652,N_14948,N_14840);
nand U15653 (N_15653,N_14352,N_14547);
nor U15654 (N_15654,N_14711,N_14956);
nand U15655 (N_15655,N_14094,N_14275);
nand U15656 (N_15656,N_14367,N_14085);
or U15657 (N_15657,N_14006,N_14470);
and U15658 (N_15658,N_14130,N_14483);
nor U15659 (N_15659,N_14616,N_14060);
xor U15660 (N_15660,N_14729,N_14544);
or U15661 (N_15661,N_14251,N_14435);
xnor U15662 (N_15662,N_14762,N_14160);
and U15663 (N_15663,N_14663,N_14458);
nand U15664 (N_15664,N_14551,N_14948);
or U15665 (N_15665,N_14137,N_14208);
nand U15666 (N_15666,N_14967,N_14647);
nand U15667 (N_15667,N_14167,N_14755);
xnor U15668 (N_15668,N_14333,N_14432);
nand U15669 (N_15669,N_14757,N_14460);
and U15670 (N_15670,N_14454,N_14847);
or U15671 (N_15671,N_14260,N_14607);
nand U15672 (N_15672,N_14553,N_14386);
and U15673 (N_15673,N_14680,N_14114);
or U15674 (N_15674,N_14879,N_14919);
xnor U15675 (N_15675,N_14437,N_14178);
nor U15676 (N_15676,N_14720,N_14166);
xnor U15677 (N_15677,N_14330,N_14119);
and U15678 (N_15678,N_14347,N_14641);
or U15679 (N_15679,N_14041,N_14438);
nor U15680 (N_15680,N_14975,N_14358);
xor U15681 (N_15681,N_14656,N_14991);
nor U15682 (N_15682,N_14294,N_14016);
nor U15683 (N_15683,N_14390,N_14134);
nor U15684 (N_15684,N_14691,N_14655);
xor U15685 (N_15685,N_14577,N_14583);
nand U15686 (N_15686,N_14576,N_14881);
xor U15687 (N_15687,N_14571,N_14025);
nor U15688 (N_15688,N_14959,N_14487);
nand U15689 (N_15689,N_14895,N_14328);
or U15690 (N_15690,N_14398,N_14852);
and U15691 (N_15691,N_14930,N_14728);
or U15692 (N_15692,N_14507,N_14134);
nand U15693 (N_15693,N_14776,N_14527);
nand U15694 (N_15694,N_14495,N_14928);
and U15695 (N_15695,N_14162,N_14969);
xnor U15696 (N_15696,N_14320,N_14512);
nor U15697 (N_15697,N_14157,N_14035);
and U15698 (N_15698,N_14534,N_14351);
nor U15699 (N_15699,N_14568,N_14618);
nand U15700 (N_15700,N_14177,N_14193);
nand U15701 (N_15701,N_14084,N_14007);
xnor U15702 (N_15702,N_14098,N_14819);
nand U15703 (N_15703,N_14689,N_14655);
xnor U15704 (N_15704,N_14644,N_14039);
xnor U15705 (N_15705,N_14690,N_14888);
xnor U15706 (N_15706,N_14942,N_14012);
nor U15707 (N_15707,N_14583,N_14069);
nand U15708 (N_15708,N_14080,N_14665);
xor U15709 (N_15709,N_14596,N_14634);
and U15710 (N_15710,N_14488,N_14260);
nor U15711 (N_15711,N_14017,N_14437);
nor U15712 (N_15712,N_14705,N_14847);
and U15713 (N_15713,N_14920,N_14069);
and U15714 (N_15714,N_14656,N_14715);
nor U15715 (N_15715,N_14791,N_14520);
xor U15716 (N_15716,N_14543,N_14748);
nor U15717 (N_15717,N_14681,N_14899);
and U15718 (N_15718,N_14158,N_14468);
nor U15719 (N_15719,N_14120,N_14979);
xor U15720 (N_15720,N_14739,N_14354);
nand U15721 (N_15721,N_14833,N_14536);
xor U15722 (N_15722,N_14132,N_14351);
and U15723 (N_15723,N_14760,N_14967);
nor U15724 (N_15724,N_14919,N_14306);
nor U15725 (N_15725,N_14527,N_14710);
nand U15726 (N_15726,N_14455,N_14561);
xor U15727 (N_15727,N_14391,N_14263);
nor U15728 (N_15728,N_14909,N_14331);
xnor U15729 (N_15729,N_14522,N_14571);
xor U15730 (N_15730,N_14543,N_14980);
xor U15731 (N_15731,N_14907,N_14795);
and U15732 (N_15732,N_14783,N_14768);
or U15733 (N_15733,N_14069,N_14092);
nand U15734 (N_15734,N_14092,N_14117);
or U15735 (N_15735,N_14681,N_14243);
nor U15736 (N_15736,N_14576,N_14656);
nor U15737 (N_15737,N_14856,N_14298);
or U15738 (N_15738,N_14556,N_14337);
and U15739 (N_15739,N_14455,N_14848);
nand U15740 (N_15740,N_14033,N_14268);
nor U15741 (N_15741,N_14067,N_14633);
and U15742 (N_15742,N_14261,N_14594);
or U15743 (N_15743,N_14810,N_14228);
nor U15744 (N_15744,N_14850,N_14109);
nor U15745 (N_15745,N_14905,N_14358);
nand U15746 (N_15746,N_14499,N_14079);
and U15747 (N_15747,N_14611,N_14650);
and U15748 (N_15748,N_14177,N_14000);
nand U15749 (N_15749,N_14774,N_14758);
xnor U15750 (N_15750,N_14141,N_14133);
nand U15751 (N_15751,N_14146,N_14044);
nand U15752 (N_15752,N_14583,N_14710);
xnor U15753 (N_15753,N_14659,N_14393);
nand U15754 (N_15754,N_14434,N_14639);
nor U15755 (N_15755,N_14745,N_14568);
nor U15756 (N_15756,N_14763,N_14849);
and U15757 (N_15757,N_14673,N_14307);
nand U15758 (N_15758,N_14746,N_14972);
nand U15759 (N_15759,N_14193,N_14995);
nor U15760 (N_15760,N_14187,N_14010);
and U15761 (N_15761,N_14200,N_14453);
xor U15762 (N_15762,N_14518,N_14440);
or U15763 (N_15763,N_14406,N_14042);
nand U15764 (N_15764,N_14212,N_14296);
or U15765 (N_15765,N_14949,N_14074);
nor U15766 (N_15766,N_14585,N_14183);
or U15767 (N_15767,N_14131,N_14331);
nand U15768 (N_15768,N_14505,N_14966);
or U15769 (N_15769,N_14797,N_14131);
and U15770 (N_15770,N_14670,N_14892);
nor U15771 (N_15771,N_14238,N_14007);
xor U15772 (N_15772,N_14339,N_14657);
xor U15773 (N_15773,N_14381,N_14665);
nand U15774 (N_15774,N_14188,N_14360);
nand U15775 (N_15775,N_14348,N_14875);
nor U15776 (N_15776,N_14221,N_14550);
nand U15777 (N_15777,N_14887,N_14307);
and U15778 (N_15778,N_14154,N_14740);
xnor U15779 (N_15779,N_14668,N_14901);
and U15780 (N_15780,N_14716,N_14142);
xor U15781 (N_15781,N_14020,N_14616);
or U15782 (N_15782,N_14431,N_14982);
or U15783 (N_15783,N_14235,N_14383);
nand U15784 (N_15784,N_14739,N_14392);
nand U15785 (N_15785,N_14452,N_14931);
or U15786 (N_15786,N_14875,N_14627);
xnor U15787 (N_15787,N_14460,N_14751);
nand U15788 (N_15788,N_14134,N_14696);
nor U15789 (N_15789,N_14263,N_14232);
or U15790 (N_15790,N_14508,N_14230);
nand U15791 (N_15791,N_14204,N_14197);
or U15792 (N_15792,N_14538,N_14986);
or U15793 (N_15793,N_14503,N_14892);
nand U15794 (N_15794,N_14217,N_14915);
or U15795 (N_15795,N_14557,N_14915);
and U15796 (N_15796,N_14461,N_14035);
nand U15797 (N_15797,N_14864,N_14815);
and U15798 (N_15798,N_14152,N_14057);
nor U15799 (N_15799,N_14360,N_14516);
or U15800 (N_15800,N_14253,N_14877);
xnor U15801 (N_15801,N_14998,N_14560);
and U15802 (N_15802,N_14594,N_14659);
and U15803 (N_15803,N_14277,N_14319);
or U15804 (N_15804,N_14716,N_14891);
and U15805 (N_15805,N_14189,N_14116);
and U15806 (N_15806,N_14891,N_14416);
xnor U15807 (N_15807,N_14322,N_14986);
xnor U15808 (N_15808,N_14370,N_14716);
or U15809 (N_15809,N_14681,N_14096);
or U15810 (N_15810,N_14683,N_14153);
xnor U15811 (N_15811,N_14762,N_14221);
xnor U15812 (N_15812,N_14958,N_14402);
or U15813 (N_15813,N_14256,N_14908);
nand U15814 (N_15814,N_14895,N_14770);
and U15815 (N_15815,N_14341,N_14147);
or U15816 (N_15816,N_14549,N_14459);
or U15817 (N_15817,N_14682,N_14719);
nand U15818 (N_15818,N_14395,N_14253);
or U15819 (N_15819,N_14610,N_14687);
xnor U15820 (N_15820,N_14435,N_14179);
and U15821 (N_15821,N_14739,N_14365);
nor U15822 (N_15822,N_14582,N_14638);
nor U15823 (N_15823,N_14394,N_14854);
nor U15824 (N_15824,N_14339,N_14590);
or U15825 (N_15825,N_14072,N_14524);
and U15826 (N_15826,N_14290,N_14286);
and U15827 (N_15827,N_14848,N_14801);
nand U15828 (N_15828,N_14142,N_14096);
nor U15829 (N_15829,N_14437,N_14103);
and U15830 (N_15830,N_14033,N_14204);
nand U15831 (N_15831,N_14270,N_14283);
or U15832 (N_15832,N_14147,N_14939);
nor U15833 (N_15833,N_14366,N_14210);
nand U15834 (N_15834,N_14286,N_14837);
or U15835 (N_15835,N_14581,N_14063);
xnor U15836 (N_15836,N_14120,N_14068);
nor U15837 (N_15837,N_14789,N_14690);
nor U15838 (N_15838,N_14827,N_14850);
nand U15839 (N_15839,N_14762,N_14697);
xor U15840 (N_15840,N_14647,N_14430);
or U15841 (N_15841,N_14416,N_14676);
nand U15842 (N_15842,N_14343,N_14454);
xnor U15843 (N_15843,N_14122,N_14533);
and U15844 (N_15844,N_14970,N_14071);
nand U15845 (N_15845,N_14789,N_14357);
and U15846 (N_15846,N_14882,N_14672);
xnor U15847 (N_15847,N_14989,N_14774);
and U15848 (N_15848,N_14606,N_14652);
nand U15849 (N_15849,N_14781,N_14453);
xor U15850 (N_15850,N_14275,N_14626);
nand U15851 (N_15851,N_14954,N_14140);
or U15852 (N_15852,N_14722,N_14236);
nand U15853 (N_15853,N_14468,N_14070);
xor U15854 (N_15854,N_14511,N_14486);
and U15855 (N_15855,N_14559,N_14439);
xnor U15856 (N_15856,N_14516,N_14314);
nand U15857 (N_15857,N_14369,N_14194);
nor U15858 (N_15858,N_14567,N_14267);
and U15859 (N_15859,N_14202,N_14483);
nor U15860 (N_15860,N_14143,N_14446);
and U15861 (N_15861,N_14600,N_14554);
nand U15862 (N_15862,N_14009,N_14072);
xor U15863 (N_15863,N_14938,N_14083);
nor U15864 (N_15864,N_14520,N_14242);
xor U15865 (N_15865,N_14177,N_14033);
nand U15866 (N_15866,N_14318,N_14224);
or U15867 (N_15867,N_14768,N_14467);
xnor U15868 (N_15868,N_14308,N_14300);
or U15869 (N_15869,N_14433,N_14742);
and U15870 (N_15870,N_14030,N_14784);
nor U15871 (N_15871,N_14517,N_14140);
nor U15872 (N_15872,N_14440,N_14510);
nand U15873 (N_15873,N_14668,N_14748);
nor U15874 (N_15874,N_14699,N_14260);
and U15875 (N_15875,N_14301,N_14752);
nor U15876 (N_15876,N_14477,N_14279);
nor U15877 (N_15877,N_14751,N_14973);
and U15878 (N_15878,N_14876,N_14720);
nand U15879 (N_15879,N_14120,N_14970);
and U15880 (N_15880,N_14410,N_14487);
nand U15881 (N_15881,N_14292,N_14319);
and U15882 (N_15882,N_14561,N_14881);
nand U15883 (N_15883,N_14493,N_14007);
xor U15884 (N_15884,N_14017,N_14926);
or U15885 (N_15885,N_14453,N_14323);
xnor U15886 (N_15886,N_14538,N_14975);
nor U15887 (N_15887,N_14045,N_14703);
xor U15888 (N_15888,N_14356,N_14554);
and U15889 (N_15889,N_14097,N_14195);
and U15890 (N_15890,N_14544,N_14113);
nand U15891 (N_15891,N_14894,N_14991);
nor U15892 (N_15892,N_14138,N_14483);
and U15893 (N_15893,N_14966,N_14370);
nand U15894 (N_15894,N_14906,N_14967);
xor U15895 (N_15895,N_14981,N_14830);
or U15896 (N_15896,N_14389,N_14594);
xnor U15897 (N_15897,N_14472,N_14700);
nand U15898 (N_15898,N_14172,N_14957);
nand U15899 (N_15899,N_14238,N_14851);
or U15900 (N_15900,N_14477,N_14979);
or U15901 (N_15901,N_14330,N_14238);
and U15902 (N_15902,N_14383,N_14148);
nand U15903 (N_15903,N_14253,N_14807);
nor U15904 (N_15904,N_14356,N_14182);
nor U15905 (N_15905,N_14088,N_14010);
xnor U15906 (N_15906,N_14009,N_14639);
nor U15907 (N_15907,N_14215,N_14514);
nand U15908 (N_15908,N_14104,N_14493);
xor U15909 (N_15909,N_14152,N_14785);
and U15910 (N_15910,N_14252,N_14707);
and U15911 (N_15911,N_14490,N_14538);
and U15912 (N_15912,N_14270,N_14089);
or U15913 (N_15913,N_14009,N_14408);
xor U15914 (N_15914,N_14688,N_14588);
or U15915 (N_15915,N_14128,N_14863);
or U15916 (N_15916,N_14119,N_14691);
or U15917 (N_15917,N_14383,N_14845);
nor U15918 (N_15918,N_14989,N_14474);
nand U15919 (N_15919,N_14967,N_14489);
nand U15920 (N_15920,N_14683,N_14780);
or U15921 (N_15921,N_14685,N_14258);
nor U15922 (N_15922,N_14954,N_14148);
nand U15923 (N_15923,N_14392,N_14526);
and U15924 (N_15924,N_14106,N_14549);
nor U15925 (N_15925,N_14933,N_14336);
nand U15926 (N_15926,N_14007,N_14337);
xor U15927 (N_15927,N_14163,N_14893);
xnor U15928 (N_15928,N_14393,N_14524);
nand U15929 (N_15929,N_14938,N_14679);
and U15930 (N_15930,N_14905,N_14791);
nor U15931 (N_15931,N_14582,N_14773);
xor U15932 (N_15932,N_14241,N_14165);
or U15933 (N_15933,N_14917,N_14286);
and U15934 (N_15934,N_14790,N_14189);
xor U15935 (N_15935,N_14468,N_14928);
xnor U15936 (N_15936,N_14328,N_14441);
nor U15937 (N_15937,N_14004,N_14443);
xor U15938 (N_15938,N_14727,N_14728);
nor U15939 (N_15939,N_14952,N_14950);
or U15940 (N_15940,N_14464,N_14614);
nand U15941 (N_15941,N_14140,N_14655);
or U15942 (N_15942,N_14366,N_14926);
xor U15943 (N_15943,N_14833,N_14829);
and U15944 (N_15944,N_14497,N_14384);
xnor U15945 (N_15945,N_14782,N_14848);
xnor U15946 (N_15946,N_14201,N_14896);
nor U15947 (N_15947,N_14339,N_14291);
xnor U15948 (N_15948,N_14632,N_14738);
and U15949 (N_15949,N_14930,N_14358);
nand U15950 (N_15950,N_14675,N_14486);
nor U15951 (N_15951,N_14816,N_14216);
nand U15952 (N_15952,N_14410,N_14092);
nor U15953 (N_15953,N_14892,N_14442);
nand U15954 (N_15954,N_14652,N_14692);
and U15955 (N_15955,N_14849,N_14370);
xnor U15956 (N_15956,N_14381,N_14223);
xnor U15957 (N_15957,N_14088,N_14707);
and U15958 (N_15958,N_14290,N_14954);
and U15959 (N_15959,N_14038,N_14061);
or U15960 (N_15960,N_14731,N_14350);
nor U15961 (N_15961,N_14140,N_14903);
nor U15962 (N_15962,N_14747,N_14165);
nor U15963 (N_15963,N_14509,N_14254);
nor U15964 (N_15964,N_14589,N_14056);
or U15965 (N_15965,N_14193,N_14468);
xor U15966 (N_15966,N_14290,N_14652);
nand U15967 (N_15967,N_14909,N_14335);
nand U15968 (N_15968,N_14743,N_14869);
nand U15969 (N_15969,N_14694,N_14547);
nor U15970 (N_15970,N_14403,N_14345);
xor U15971 (N_15971,N_14308,N_14195);
xor U15972 (N_15972,N_14282,N_14542);
xnor U15973 (N_15973,N_14721,N_14042);
xor U15974 (N_15974,N_14714,N_14102);
or U15975 (N_15975,N_14009,N_14530);
nor U15976 (N_15976,N_14800,N_14164);
xnor U15977 (N_15977,N_14229,N_14615);
xnor U15978 (N_15978,N_14558,N_14363);
and U15979 (N_15979,N_14727,N_14009);
nor U15980 (N_15980,N_14412,N_14596);
nand U15981 (N_15981,N_14210,N_14792);
or U15982 (N_15982,N_14873,N_14001);
and U15983 (N_15983,N_14991,N_14943);
and U15984 (N_15984,N_14538,N_14243);
and U15985 (N_15985,N_14193,N_14254);
nand U15986 (N_15986,N_14743,N_14346);
nand U15987 (N_15987,N_14476,N_14570);
nand U15988 (N_15988,N_14093,N_14018);
or U15989 (N_15989,N_14314,N_14076);
xor U15990 (N_15990,N_14520,N_14685);
nor U15991 (N_15991,N_14076,N_14921);
nand U15992 (N_15992,N_14472,N_14452);
and U15993 (N_15993,N_14183,N_14972);
xnor U15994 (N_15994,N_14780,N_14112);
or U15995 (N_15995,N_14064,N_14306);
and U15996 (N_15996,N_14937,N_14562);
and U15997 (N_15997,N_14369,N_14927);
nor U15998 (N_15998,N_14796,N_14456);
and U15999 (N_15999,N_14787,N_14210);
xor U16000 (N_16000,N_15172,N_15888);
or U16001 (N_16001,N_15929,N_15443);
xnor U16002 (N_16002,N_15072,N_15787);
and U16003 (N_16003,N_15703,N_15613);
xor U16004 (N_16004,N_15115,N_15418);
nand U16005 (N_16005,N_15351,N_15565);
and U16006 (N_16006,N_15191,N_15931);
xor U16007 (N_16007,N_15981,N_15283);
nor U16008 (N_16008,N_15642,N_15951);
and U16009 (N_16009,N_15815,N_15405);
nand U16010 (N_16010,N_15227,N_15907);
or U16011 (N_16011,N_15204,N_15450);
nor U16012 (N_16012,N_15140,N_15767);
nand U16013 (N_16013,N_15363,N_15459);
nand U16014 (N_16014,N_15282,N_15202);
and U16015 (N_16015,N_15148,N_15725);
nor U16016 (N_16016,N_15924,N_15686);
xnor U16017 (N_16017,N_15223,N_15723);
nand U16018 (N_16018,N_15315,N_15597);
or U16019 (N_16019,N_15238,N_15831);
or U16020 (N_16020,N_15491,N_15999);
xor U16021 (N_16021,N_15112,N_15380);
and U16022 (N_16022,N_15068,N_15819);
xnor U16023 (N_16023,N_15991,N_15231);
or U16024 (N_16024,N_15938,N_15063);
nand U16025 (N_16025,N_15579,N_15937);
xor U16026 (N_16026,N_15697,N_15113);
or U16027 (N_16027,N_15719,N_15590);
and U16028 (N_16028,N_15521,N_15838);
xor U16029 (N_16029,N_15034,N_15196);
and U16030 (N_16030,N_15249,N_15095);
xnor U16031 (N_16031,N_15587,N_15771);
nand U16032 (N_16032,N_15673,N_15812);
and U16033 (N_16033,N_15147,N_15466);
nor U16034 (N_16034,N_15876,N_15846);
nand U16035 (N_16035,N_15904,N_15626);
xor U16036 (N_16036,N_15615,N_15797);
xor U16037 (N_16037,N_15500,N_15326);
and U16038 (N_16038,N_15990,N_15738);
xor U16039 (N_16039,N_15395,N_15736);
nor U16040 (N_16040,N_15858,N_15588);
and U16041 (N_16041,N_15292,N_15730);
xnor U16042 (N_16042,N_15643,N_15414);
and U16043 (N_16043,N_15277,N_15535);
or U16044 (N_16044,N_15605,N_15765);
and U16045 (N_16045,N_15547,N_15941);
and U16046 (N_16046,N_15811,N_15229);
nor U16047 (N_16047,N_15375,N_15413);
nor U16048 (N_16048,N_15632,N_15721);
nor U16049 (N_16049,N_15988,N_15728);
or U16050 (N_16050,N_15260,N_15267);
or U16051 (N_16051,N_15825,N_15653);
nand U16052 (N_16052,N_15428,N_15665);
or U16053 (N_16053,N_15659,N_15798);
and U16054 (N_16054,N_15671,N_15756);
nor U16055 (N_16055,N_15293,N_15766);
xor U16056 (N_16056,N_15483,N_15928);
nor U16057 (N_16057,N_15463,N_15799);
and U16058 (N_16058,N_15207,N_15830);
or U16059 (N_16059,N_15433,N_15410);
xor U16060 (N_16060,N_15821,N_15108);
nor U16061 (N_16061,N_15447,N_15442);
or U16062 (N_16062,N_15000,N_15852);
nand U16063 (N_16063,N_15402,N_15173);
xor U16064 (N_16064,N_15814,N_15120);
or U16065 (N_16065,N_15305,N_15685);
nand U16066 (N_16066,N_15142,N_15822);
xor U16067 (N_16067,N_15906,N_15083);
xor U16068 (N_16068,N_15166,N_15054);
xor U16069 (N_16069,N_15057,N_15015);
and U16070 (N_16070,N_15397,N_15412);
nand U16071 (N_16071,N_15183,N_15064);
or U16072 (N_16072,N_15448,N_15704);
nor U16073 (N_16073,N_15969,N_15808);
or U16074 (N_16074,N_15340,N_15435);
xor U16075 (N_16075,N_15079,N_15194);
nor U16076 (N_16076,N_15549,N_15836);
xnor U16077 (N_16077,N_15584,N_15657);
and U16078 (N_16078,N_15827,N_15263);
or U16079 (N_16079,N_15205,N_15037);
xnor U16080 (N_16080,N_15854,N_15520);
or U16081 (N_16081,N_15461,N_15592);
or U16082 (N_16082,N_15634,N_15201);
nor U16083 (N_16083,N_15700,N_15984);
xor U16084 (N_16084,N_15155,N_15917);
xnor U16085 (N_16085,N_15041,N_15832);
and U16086 (N_16086,N_15385,N_15135);
xnor U16087 (N_16087,N_15608,N_15646);
nor U16088 (N_16088,N_15705,N_15633);
xnor U16089 (N_16089,N_15164,N_15768);
nor U16090 (N_16090,N_15694,N_15962);
or U16091 (N_16091,N_15058,N_15562);
and U16092 (N_16092,N_15949,N_15366);
nand U16093 (N_16093,N_15022,N_15559);
and U16094 (N_16094,N_15474,N_15291);
nand U16095 (N_16095,N_15880,N_15921);
xnor U16096 (N_16096,N_15722,N_15099);
xnor U16097 (N_16097,N_15488,N_15735);
or U16098 (N_16098,N_15352,N_15525);
nand U16099 (N_16099,N_15137,N_15593);
nand U16100 (N_16100,N_15645,N_15975);
or U16101 (N_16101,N_15048,N_15689);
nand U16102 (N_16102,N_15098,N_15104);
nand U16103 (N_16103,N_15075,N_15629);
and U16104 (N_16104,N_15555,N_15641);
nand U16105 (N_16105,N_15720,N_15499);
nor U16106 (N_16106,N_15586,N_15308);
or U16107 (N_16107,N_15698,N_15986);
or U16108 (N_16108,N_15853,N_15900);
xor U16109 (N_16109,N_15234,N_15253);
nand U16110 (N_16110,N_15387,N_15367);
xor U16111 (N_16111,N_15203,N_15976);
nor U16112 (N_16112,N_15709,N_15649);
or U16113 (N_16113,N_15193,N_15237);
nor U16114 (N_16114,N_15136,N_15561);
xor U16115 (N_16115,N_15651,N_15493);
or U16116 (N_16116,N_15464,N_15431);
and U16117 (N_16117,N_15751,N_15716);
nand U16118 (N_16118,N_15742,N_15603);
or U16119 (N_16119,N_15407,N_15256);
or U16120 (N_16120,N_15262,N_15779);
xor U16121 (N_16121,N_15954,N_15701);
and U16122 (N_16122,N_15328,N_15492);
and U16123 (N_16123,N_15837,N_15732);
xnor U16124 (N_16124,N_15222,N_15484);
nand U16125 (N_16125,N_15743,N_15866);
nor U16126 (N_16126,N_15364,N_15179);
nand U16127 (N_16127,N_15446,N_15420);
or U16128 (N_16128,N_15266,N_15995);
xor U16129 (N_16129,N_15760,N_15080);
and U16130 (N_16130,N_15871,N_15254);
and U16131 (N_16131,N_15206,N_15043);
nor U16132 (N_16132,N_15211,N_15131);
nand U16133 (N_16133,N_15505,N_15388);
or U16134 (N_16134,N_15383,N_15033);
or U16135 (N_16135,N_15576,N_15750);
xnor U16136 (N_16136,N_15895,N_15512);
nor U16137 (N_16137,N_15806,N_15479);
or U16138 (N_16138,N_15497,N_15539);
nand U16139 (N_16139,N_15882,N_15478);
nor U16140 (N_16140,N_15240,N_15910);
nand U16141 (N_16141,N_15920,N_15905);
xor U16142 (N_16142,N_15176,N_15485);
xnor U16143 (N_16143,N_15517,N_15486);
xor U16144 (N_16144,N_15423,N_15655);
nand U16145 (N_16145,N_15225,N_15745);
nor U16146 (N_16146,N_15272,N_15153);
nor U16147 (N_16147,N_15636,N_15506);
nor U16148 (N_16148,N_15144,N_15898);
xnor U16149 (N_16149,N_15313,N_15213);
or U16150 (N_16150,N_15609,N_15758);
or U16151 (N_16151,N_15785,N_15356);
or U16152 (N_16152,N_15312,N_15596);
and U16153 (N_16153,N_15169,N_15740);
nor U16154 (N_16154,N_15754,N_15824);
nand U16155 (N_16155,N_15016,N_15829);
or U16156 (N_16156,N_15394,N_15541);
and U16157 (N_16157,N_15945,N_15175);
nand U16158 (N_16158,N_15580,N_15970);
nand U16159 (N_16159,N_15612,N_15417);
or U16160 (N_16160,N_15384,N_15794);
xor U16161 (N_16161,N_15971,N_15059);
nor U16162 (N_16162,N_15027,N_15557);
and U16163 (N_16163,N_15069,N_15350);
and U16164 (N_16164,N_15803,N_15001);
and U16165 (N_16165,N_15040,N_15449);
nor U16166 (N_16166,N_15729,N_15759);
or U16167 (N_16167,N_15828,N_15601);
nand U16168 (N_16168,N_15585,N_15875);
or U16169 (N_16169,N_15322,N_15044);
or U16170 (N_16170,N_15560,N_15024);
or U16171 (N_16171,N_15070,N_15973);
or U16172 (N_16172,N_15713,N_15092);
nor U16173 (N_16173,N_15323,N_15595);
or U16174 (N_16174,N_15977,N_15556);
and U16175 (N_16175,N_15167,N_15473);
nor U16176 (N_16176,N_15007,N_15067);
nand U16177 (N_16177,N_15424,N_15494);
or U16178 (N_16178,N_15869,N_15021);
xnor U16179 (N_16179,N_15490,N_15020);
nand U16180 (N_16180,N_15285,N_15933);
or U16181 (N_16181,N_15273,N_15763);
nand U16182 (N_16182,N_15564,N_15019);
or U16183 (N_16183,N_15538,N_15747);
or U16184 (N_16184,N_15246,N_15823);
or U16185 (N_16185,N_15269,N_15746);
and U16186 (N_16186,N_15582,N_15036);
or U16187 (N_16187,N_15950,N_15879);
or U16188 (N_16188,N_15839,N_15014);
or U16189 (N_16189,N_15679,N_15923);
or U16190 (N_16190,N_15245,N_15084);
and U16191 (N_16191,N_15338,N_15537);
xor U16192 (N_16192,N_15124,N_15476);
xor U16193 (N_16193,N_15878,N_15724);
or U16194 (N_16194,N_15681,N_15631);
nand U16195 (N_16195,N_15526,N_15310);
and U16196 (N_16196,N_15727,N_15856);
nand U16197 (N_16197,N_15158,N_15678);
xor U16198 (N_16198,N_15082,N_15668);
and U16199 (N_16199,N_15516,N_15749);
and U16200 (N_16200,N_15816,N_15863);
nor U16201 (N_16201,N_15451,N_15487);
nor U16202 (N_16202,N_15542,N_15130);
xor U16203 (N_16203,N_15445,N_15126);
and U16204 (N_16204,N_15826,N_15699);
and U16205 (N_16205,N_15983,N_15029);
xor U16206 (N_16206,N_15004,N_15091);
or U16207 (N_16207,N_15648,N_15170);
and U16208 (N_16208,N_15536,N_15706);
nand U16209 (N_16209,N_15873,N_15925);
nor U16210 (N_16210,N_15242,N_15687);
nor U16211 (N_16211,N_15885,N_15307);
and U16212 (N_16212,N_15591,N_15770);
or U16213 (N_16213,N_15477,N_15421);
nor U16214 (N_16214,N_15133,N_15711);
xor U16215 (N_16215,N_15119,N_15660);
nor U16216 (N_16216,N_15100,N_15437);
xor U16217 (N_16217,N_15683,N_15300);
nor U16218 (N_16218,N_15287,N_15049);
nor U16219 (N_16219,N_15411,N_15061);
or U16220 (N_16220,N_15845,N_15677);
or U16221 (N_16221,N_15042,N_15047);
nor U16222 (N_16222,N_15009,N_15475);
and U16223 (N_16223,N_15343,N_15220);
xnor U16224 (N_16224,N_15553,N_15141);
or U16225 (N_16225,N_15399,N_15422);
nand U16226 (N_16226,N_15532,N_15214);
nor U16227 (N_16227,N_15200,N_15919);
or U16228 (N_16228,N_15224,N_15509);
nand U16229 (N_16229,N_15341,N_15997);
and U16230 (N_16230,N_15345,N_15122);
and U16231 (N_16231,N_15165,N_15748);
and U16232 (N_16232,N_15622,N_15502);
or U16233 (N_16233,N_15623,N_15355);
xnor U16234 (N_16234,N_15480,N_15056);
nand U16235 (N_16235,N_15843,N_15501);
nand U16236 (N_16236,N_15780,N_15400);
and U16237 (N_16237,N_15334,N_15031);
xnor U16238 (N_16238,N_15777,N_15666);
or U16239 (N_16239,N_15149,N_15373);
or U16240 (N_16240,N_15216,N_15081);
and U16241 (N_16241,N_15255,N_15469);
and U16242 (N_16242,N_15299,N_15775);
nand U16243 (N_16243,N_15909,N_15809);
xnor U16244 (N_16244,N_15504,N_15614);
nor U16245 (N_16245,N_15918,N_15154);
xor U16246 (N_16246,N_15050,N_15381);
and U16247 (N_16247,N_15891,N_15163);
xnor U16248 (N_16248,N_15415,N_15864);
xnor U16249 (N_16249,N_15602,N_15911);
and U16250 (N_16250,N_15624,N_15670);
nor U16251 (N_16251,N_15090,N_15489);
nor U16252 (N_16252,N_15529,N_15996);
nand U16253 (N_16253,N_15077,N_15693);
nor U16254 (N_16254,N_15181,N_15757);
and U16255 (N_16255,N_15319,N_15270);
xnor U16256 (N_16256,N_15708,N_15248);
xor U16257 (N_16257,N_15610,N_15177);
nor U16258 (N_16258,N_15017,N_15524);
nand U16259 (N_16259,N_15638,N_15055);
xor U16260 (N_16260,N_15637,N_15859);
nor U16261 (N_16261,N_15128,N_15661);
and U16262 (N_16262,N_15134,N_15008);
and U16263 (N_16263,N_15235,N_15114);
nor U16264 (N_16264,N_15051,N_15625);
nor U16265 (N_16265,N_15250,N_15994);
nor U16266 (N_16266,N_15886,N_15406);
or U16267 (N_16267,N_15023,N_15534);
and U16268 (N_16268,N_15573,N_15288);
nand U16269 (N_16269,N_15718,N_15676);
nor U16270 (N_16270,N_15271,N_15965);
or U16271 (N_16271,N_15887,N_15786);
or U16272 (N_16272,N_15953,N_15993);
nor U16273 (N_16273,N_15842,N_15574);
and U16274 (N_16274,N_15012,N_15890);
xor U16275 (N_16275,N_15046,N_15662);
and U16276 (N_16276,N_15978,N_15003);
xnor U16277 (N_16277,N_15302,N_15457);
or U16278 (N_16278,N_15324,N_15386);
or U16279 (N_16279,N_15374,N_15416);
nand U16280 (N_16280,N_15569,N_15578);
or U16281 (N_16281,N_15784,N_15835);
or U16282 (N_16282,N_15789,N_15184);
nand U16283 (N_16283,N_15316,N_15377);
or U16284 (N_16284,N_15604,N_15752);
nor U16285 (N_16285,N_15434,N_15296);
nand U16286 (N_16286,N_15208,N_15301);
xnor U16287 (N_16287,N_15939,N_15030);
nand U16288 (N_16288,N_15178,N_15116);
nor U16289 (N_16289,N_15371,N_15897);
xnor U16290 (N_16290,N_15289,N_15998);
and U16291 (N_16291,N_15782,N_15519);
xnor U16292 (N_16292,N_15279,N_15465);
nor U16293 (N_16293,N_15792,N_15074);
nand U16294 (N_16294,N_15966,N_15714);
xor U16295 (N_16295,N_15947,N_15396);
and U16296 (N_16296,N_15621,N_15598);
nor U16297 (N_16297,N_15453,N_15514);
and U16298 (N_16298,N_15548,N_15664);
xnor U16299 (N_16299,N_15157,N_15106);
or U16300 (N_16300,N_15810,N_15353);
xnor U16301 (N_16301,N_15073,N_15159);
and U16302 (N_16302,N_15168,N_15382);
nor U16303 (N_16303,N_15276,N_15393);
and U16304 (N_16304,N_15795,N_15972);
xor U16305 (N_16305,N_15989,N_15652);
xnor U16306 (N_16306,N_15861,N_15259);
and U16307 (N_16307,N_15425,N_15817);
or U16308 (N_16308,N_15550,N_15849);
nor U16309 (N_16309,N_15791,N_15118);
and U16310 (N_16310,N_15675,N_15755);
and U16311 (N_16311,N_15132,N_15093);
or U16312 (N_16312,N_15545,N_15065);
or U16313 (N_16313,N_15577,N_15712);
or U16314 (N_16314,N_15640,N_15498);
nand U16315 (N_16315,N_15589,N_15028);
and U16316 (N_16316,N_15635,N_15688);
nand U16317 (N_16317,N_15802,N_15894);
nand U16318 (N_16318,N_15117,N_15889);
and U16319 (N_16319,N_15575,N_15109);
nor U16320 (N_16320,N_15199,N_15855);
nor U16321 (N_16321,N_15913,N_15357);
xor U16322 (N_16322,N_15527,N_15195);
or U16323 (N_16323,N_15268,N_15533);
xor U16324 (N_16324,N_15097,N_15121);
nor U16325 (N_16325,N_15303,N_15339);
or U16326 (N_16326,N_15959,N_15197);
nand U16327 (N_16327,N_15228,N_15820);
nand U16328 (N_16328,N_15600,N_15311);
xor U16329 (N_16329,N_15684,N_15731);
and U16330 (N_16330,N_15335,N_15974);
or U16331 (N_16331,N_15964,N_15346);
nor U16332 (N_16332,N_15439,N_15628);
xnor U16333 (N_16333,N_15129,N_15967);
xnor U16334 (N_16334,N_15005,N_15275);
nand U16335 (N_16335,N_15523,N_15510);
nand U16336 (N_16336,N_15813,N_15680);
nor U16337 (N_16337,N_15101,N_15060);
nor U16338 (N_16338,N_15252,N_15801);
or U16339 (N_16339,N_15543,N_15111);
nor U16340 (N_16340,N_15644,N_15881);
xnor U16341 (N_16341,N_15247,N_15985);
and U16342 (N_16342,N_15281,N_15123);
xnor U16343 (N_16343,N_15314,N_15327);
xor U16344 (N_16344,N_15125,N_15552);
or U16345 (N_16345,N_15934,N_15554);
or U16346 (N_16346,N_15682,N_15800);
or U16347 (N_16347,N_15440,N_15233);
xor U16348 (N_16348,N_15215,N_15943);
and U16349 (N_16349,N_15026,N_15304);
nand U16350 (N_16350,N_15696,N_15715);
nand U16351 (N_16351,N_15370,N_15778);
nor U16352 (N_16352,N_15658,N_15330);
and U16353 (N_16353,N_15734,N_15209);
nor U16354 (N_16354,N_15518,N_15567);
and U16355 (N_16355,N_15805,N_15744);
nand U16356 (N_16356,N_15348,N_15409);
nand U16357 (N_16357,N_15025,N_15896);
nand U16358 (N_16358,N_15221,N_15035);
or U16359 (N_16359,N_15432,N_15515);
nand U16360 (N_16360,N_15217,N_15607);
or U16361 (N_16361,N_15188,N_15702);
nor U16362 (N_16362,N_15558,N_15438);
xor U16363 (N_16363,N_15261,N_15764);
xnor U16364 (N_16364,N_15926,N_15606);
and U16365 (N_16365,N_15963,N_15583);
nor U16366 (N_16366,N_15707,N_15337);
nor U16367 (N_16367,N_15306,N_15690);
xor U16368 (N_16368,N_15390,N_15062);
or U16369 (N_16369,N_15455,N_15982);
nor U16370 (N_16370,N_15290,N_15672);
and U16371 (N_16371,N_15860,N_15189);
nor U16372 (N_16372,N_15987,N_15695);
nor U16373 (N_16373,N_15544,N_15865);
and U16374 (N_16374,N_15344,N_15944);
xnor U16375 (N_16375,N_15392,N_15317);
xor U16376 (N_16376,N_15495,N_15156);
nor U16377 (N_16377,N_15472,N_15710);
and U16378 (N_16378,N_15088,N_15236);
nor U16379 (N_16379,N_15389,N_15232);
and U16380 (N_16380,N_15460,N_15572);
nor U16381 (N_16381,N_15329,N_15654);
or U16382 (N_16382,N_15807,N_15226);
and U16383 (N_16383,N_15733,N_15462);
nor U16384 (N_16384,N_15912,N_15620);
and U16385 (N_16385,N_15468,N_15663);
and U16386 (N_16386,N_15427,N_15467);
xor U16387 (N_16387,N_15833,N_15511);
and U16388 (N_16388,N_15650,N_15528);
nand U16389 (N_16389,N_15737,N_15139);
or U16390 (N_16390,N_15094,N_15360);
or U16391 (N_16391,N_15630,N_15401);
and U16392 (N_16392,N_15066,N_15076);
xnor U16393 (N_16393,N_15530,N_15930);
or U16394 (N_16394,N_15834,N_15772);
xnor U16395 (N_16395,N_15325,N_15470);
or U16396 (N_16396,N_15127,N_15368);
xnor U16397 (N_16397,N_15336,N_15096);
or U16398 (N_16398,N_15150,N_15298);
or U16399 (N_16399,N_15230,N_15739);
and U16400 (N_16400,N_15619,N_15187);
xnor U16401 (N_16401,N_15883,N_15916);
and U16402 (N_16402,N_15085,N_15927);
nor U16403 (N_16403,N_15741,N_15874);
nor U16404 (N_16404,N_15948,N_15570);
xnor U16405 (N_16405,N_15185,N_15089);
xnor U16406 (N_16406,N_15251,N_15294);
and U16407 (N_16407,N_15376,N_15192);
nor U16408 (N_16408,N_15320,N_15145);
nand U16409 (N_16409,N_15243,N_15404);
nand U16410 (N_16410,N_15331,N_15171);
and U16411 (N_16411,N_15430,N_15956);
xor U16412 (N_16412,N_15110,N_15773);
or U16413 (N_16413,N_15398,N_15297);
xnor U16414 (N_16414,N_15753,N_15274);
xnor U16415 (N_16415,N_15979,N_15471);
or U16416 (N_16416,N_15551,N_15482);
nor U16417 (N_16417,N_15496,N_15295);
nand U16418 (N_16418,N_15162,N_15940);
and U16419 (N_16419,N_15952,N_15342);
nand U16420 (N_16420,N_15508,N_15361);
xor U16421 (N_16421,N_15309,N_15265);
nor U16422 (N_16422,N_15408,N_15152);
and U16423 (N_16423,N_15102,N_15513);
nand U16424 (N_16424,N_15992,N_15656);
and U16425 (N_16425,N_15796,N_15053);
nand U16426 (N_16426,N_15507,N_15667);
xor U16427 (N_16427,N_15793,N_15781);
and U16428 (N_16428,N_15958,N_15006);
or U16429 (N_16429,N_15627,N_15540);
xnor U16430 (N_16430,N_15844,N_15378);
nor U16431 (N_16431,N_15901,N_15870);
and U16432 (N_16432,N_15071,N_15946);
nand U16433 (N_16433,N_15426,N_15674);
nand U16434 (N_16434,N_15321,N_15481);
nand U16435 (N_16435,N_15349,N_15138);
or U16436 (N_16436,N_15045,N_15914);
nand U16437 (N_16437,N_15531,N_15354);
or U16438 (N_16438,N_15892,N_15454);
or U16439 (N_16439,N_15761,N_15618);
nand U16440 (N_16440,N_15258,N_15862);
nor U16441 (N_16441,N_15444,N_15280);
or U16442 (N_16442,N_15818,N_15563);
nor U16443 (N_16443,N_15616,N_15241);
or U16444 (N_16444,N_15010,N_15932);
and U16445 (N_16445,N_15286,N_15955);
nand U16446 (N_16446,N_15915,N_15333);
and U16447 (N_16447,N_15935,N_15086);
nand U16448 (N_16448,N_15039,N_15669);
nand U16449 (N_16449,N_15571,N_15284);
xnor U16450 (N_16450,N_15639,N_15219);
nor U16451 (N_16451,N_15899,N_15790);
xor U16452 (N_16452,N_15372,N_15968);
and U16453 (N_16453,N_15503,N_15143);
nand U16454 (N_16454,N_15936,N_15332);
xor U16455 (N_16455,N_15180,N_15867);
or U16456 (N_16456,N_15002,N_15419);
and U16457 (N_16457,N_15018,N_15052);
nand U16458 (N_16458,N_15452,N_15429);
and U16459 (N_16459,N_15013,N_15960);
xnor U16460 (N_16460,N_15957,N_15851);
or U16461 (N_16461,N_15961,N_15847);
xor U16462 (N_16462,N_15762,N_15617);
nor U16463 (N_16463,N_15776,N_15868);
or U16464 (N_16464,N_15198,N_15726);
nand U16465 (N_16465,N_15391,N_15257);
xor U16466 (N_16466,N_15884,N_15032);
xnor U16467 (N_16467,N_15038,N_15893);
nand U16468 (N_16468,N_15212,N_15369);
nand U16469 (N_16469,N_15872,N_15087);
or U16470 (N_16470,N_15647,N_15788);
nand U16471 (N_16471,N_15318,N_15078);
or U16472 (N_16472,N_15186,N_15161);
nand U16473 (N_16473,N_15458,N_15902);
nand U16474 (N_16474,N_15611,N_15599);
or U16475 (N_16475,N_15903,N_15568);
and U16476 (N_16476,N_15804,N_15174);
and U16477 (N_16477,N_15848,N_15908);
nor U16478 (N_16478,N_15011,N_15359);
nand U16479 (N_16479,N_15840,N_15436);
nand U16480 (N_16480,N_15210,N_15151);
xor U16481 (N_16481,N_15522,N_15456);
nor U16482 (N_16482,N_15850,N_15717);
xor U16483 (N_16483,N_15105,N_15365);
nor U16484 (N_16484,N_15691,N_15769);
xor U16485 (N_16485,N_15783,N_15857);
xnor U16486 (N_16486,N_15218,N_15239);
xor U16487 (N_16487,N_15362,N_15877);
xnor U16488 (N_16488,N_15146,N_15103);
xnor U16489 (N_16489,N_15347,N_15566);
or U16490 (N_16490,N_15581,N_15244);
nand U16491 (N_16491,N_15190,N_15594);
xnor U16492 (N_16492,N_15692,N_15182);
nand U16493 (N_16493,N_15278,N_15379);
nand U16494 (N_16494,N_15942,N_15980);
or U16495 (N_16495,N_15841,N_15922);
and U16496 (N_16496,N_15264,N_15403);
nor U16497 (N_16497,N_15160,N_15107);
xor U16498 (N_16498,N_15358,N_15546);
xor U16499 (N_16499,N_15774,N_15441);
and U16500 (N_16500,N_15835,N_15497);
and U16501 (N_16501,N_15132,N_15283);
xor U16502 (N_16502,N_15953,N_15326);
xnor U16503 (N_16503,N_15971,N_15922);
nand U16504 (N_16504,N_15142,N_15769);
nor U16505 (N_16505,N_15128,N_15180);
or U16506 (N_16506,N_15023,N_15609);
nand U16507 (N_16507,N_15158,N_15255);
xnor U16508 (N_16508,N_15993,N_15688);
or U16509 (N_16509,N_15818,N_15835);
xor U16510 (N_16510,N_15069,N_15398);
nor U16511 (N_16511,N_15310,N_15596);
and U16512 (N_16512,N_15279,N_15325);
nor U16513 (N_16513,N_15485,N_15338);
and U16514 (N_16514,N_15348,N_15959);
and U16515 (N_16515,N_15615,N_15155);
xnor U16516 (N_16516,N_15598,N_15602);
nand U16517 (N_16517,N_15522,N_15194);
xor U16518 (N_16518,N_15296,N_15074);
xor U16519 (N_16519,N_15793,N_15526);
nand U16520 (N_16520,N_15220,N_15671);
nor U16521 (N_16521,N_15921,N_15320);
xor U16522 (N_16522,N_15237,N_15078);
nand U16523 (N_16523,N_15747,N_15392);
and U16524 (N_16524,N_15474,N_15567);
nand U16525 (N_16525,N_15409,N_15589);
nand U16526 (N_16526,N_15855,N_15016);
nand U16527 (N_16527,N_15891,N_15792);
nand U16528 (N_16528,N_15524,N_15372);
nand U16529 (N_16529,N_15006,N_15765);
nand U16530 (N_16530,N_15684,N_15970);
and U16531 (N_16531,N_15050,N_15198);
nor U16532 (N_16532,N_15055,N_15695);
and U16533 (N_16533,N_15797,N_15543);
and U16534 (N_16534,N_15218,N_15151);
and U16535 (N_16535,N_15408,N_15318);
nor U16536 (N_16536,N_15180,N_15327);
nor U16537 (N_16537,N_15618,N_15853);
xor U16538 (N_16538,N_15975,N_15059);
xor U16539 (N_16539,N_15412,N_15185);
nor U16540 (N_16540,N_15012,N_15886);
or U16541 (N_16541,N_15403,N_15299);
xor U16542 (N_16542,N_15109,N_15063);
xor U16543 (N_16543,N_15043,N_15713);
nor U16544 (N_16544,N_15083,N_15848);
nor U16545 (N_16545,N_15901,N_15178);
nand U16546 (N_16546,N_15119,N_15465);
xor U16547 (N_16547,N_15895,N_15127);
nand U16548 (N_16548,N_15921,N_15019);
and U16549 (N_16549,N_15974,N_15388);
nor U16550 (N_16550,N_15477,N_15819);
xnor U16551 (N_16551,N_15299,N_15506);
and U16552 (N_16552,N_15598,N_15639);
xnor U16553 (N_16553,N_15974,N_15924);
nand U16554 (N_16554,N_15147,N_15597);
nor U16555 (N_16555,N_15257,N_15685);
nor U16556 (N_16556,N_15368,N_15409);
and U16557 (N_16557,N_15235,N_15312);
xor U16558 (N_16558,N_15440,N_15699);
nand U16559 (N_16559,N_15859,N_15068);
nor U16560 (N_16560,N_15260,N_15549);
or U16561 (N_16561,N_15629,N_15058);
nand U16562 (N_16562,N_15017,N_15749);
nand U16563 (N_16563,N_15339,N_15649);
nor U16564 (N_16564,N_15888,N_15691);
xor U16565 (N_16565,N_15616,N_15251);
and U16566 (N_16566,N_15130,N_15809);
and U16567 (N_16567,N_15115,N_15882);
or U16568 (N_16568,N_15171,N_15525);
nand U16569 (N_16569,N_15975,N_15101);
nand U16570 (N_16570,N_15064,N_15652);
nand U16571 (N_16571,N_15212,N_15620);
nand U16572 (N_16572,N_15211,N_15767);
or U16573 (N_16573,N_15927,N_15207);
xor U16574 (N_16574,N_15970,N_15108);
xnor U16575 (N_16575,N_15530,N_15818);
and U16576 (N_16576,N_15410,N_15091);
nand U16577 (N_16577,N_15287,N_15568);
nand U16578 (N_16578,N_15971,N_15612);
nor U16579 (N_16579,N_15941,N_15533);
xor U16580 (N_16580,N_15710,N_15041);
or U16581 (N_16581,N_15837,N_15769);
nor U16582 (N_16582,N_15251,N_15611);
nor U16583 (N_16583,N_15858,N_15078);
xnor U16584 (N_16584,N_15561,N_15962);
nor U16585 (N_16585,N_15908,N_15734);
and U16586 (N_16586,N_15807,N_15421);
nand U16587 (N_16587,N_15036,N_15318);
xor U16588 (N_16588,N_15005,N_15539);
and U16589 (N_16589,N_15438,N_15998);
or U16590 (N_16590,N_15828,N_15637);
nand U16591 (N_16591,N_15405,N_15669);
xor U16592 (N_16592,N_15369,N_15021);
or U16593 (N_16593,N_15459,N_15105);
xor U16594 (N_16594,N_15437,N_15897);
nand U16595 (N_16595,N_15689,N_15697);
and U16596 (N_16596,N_15099,N_15955);
xnor U16597 (N_16597,N_15200,N_15428);
nor U16598 (N_16598,N_15939,N_15754);
and U16599 (N_16599,N_15606,N_15030);
xor U16600 (N_16600,N_15342,N_15788);
nand U16601 (N_16601,N_15146,N_15479);
and U16602 (N_16602,N_15191,N_15915);
xnor U16603 (N_16603,N_15891,N_15295);
nor U16604 (N_16604,N_15291,N_15420);
or U16605 (N_16605,N_15757,N_15516);
or U16606 (N_16606,N_15837,N_15824);
nand U16607 (N_16607,N_15539,N_15764);
xnor U16608 (N_16608,N_15120,N_15723);
nand U16609 (N_16609,N_15613,N_15296);
xor U16610 (N_16610,N_15528,N_15553);
nor U16611 (N_16611,N_15267,N_15378);
or U16612 (N_16612,N_15852,N_15404);
nand U16613 (N_16613,N_15378,N_15285);
xor U16614 (N_16614,N_15431,N_15806);
or U16615 (N_16615,N_15602,N_15005);
nand U16616 (N_16616,N_15008,N_15224);
or U16617 (N_16617,N_15007,N_15507);
nor U16618 (N_16618,N_15297,N_15953);
and U16619 (N_16619,N_15705,N_15156);
nand U16620 (N_16620,N_15987,N_15781);
nor U16621 (N_16621,N_15689,N_15993);
xnor U16622 (N_16622,N_15642,N_15325);
nand U16623 (N_16623,N_15186,N_15824);
and U16624 (N_16624,N_15143,N_15607);
and U16625 (N_16625,N_15798,N_15914);
nand U16626 (N_16626,N_15838,N_15087);
nand U16627 (N_16627,N_15307,N_15284);
nand U16628 (N_16628,N_15014,N_15654);
and U16629 (N_16629,N_15900,N_15730);
and U16630 (N_16630,N_15110,N_15419);
or U16631 (N_16631,N_15496,N_15119);
nand U16632 (N_16632,N_15684,N_15323);
or U16633 (N_16633,N_15137,N_15624);
and U16634 (N_16634,N_15297,N_15904);
nand U16635 (N_16635,N_15536,N_15910);
xnor U16636 (N_16636,N_15740,N_15277);
nand U16637 (N_16637,N_15242,N_15954);
nor U16638 (N_16638,N_15127,N_15944);
or U16639 (N_16639,N_15243,N_15528);
and U16640 (N_16640,N_15447,N_15586);
nor U16641 (N_16641,N_15171,N_15944);
and U16642 (N_16642,N_15639,N_15201);
xor U16643 (N_16643,N_15575,N_15681);
and U16644 (N_16644,N_15916,N_15717);
nor U16645 (N_16645,N_15541,N_15832);
nor U16646 (N_16646,N_15649,N_15812);
nand U16647 (N_16647,N_15427,N_15517);
or U16648 (N_16648,N_15900,N_15308);
xor U16649 (N_16649,N_15810,N_15609);
nor U16650 (N_16650,N_15748,N_15185);
and U16651 (N_16651,N_15563,N_15617);
and U16652 (N_16652,N_15185,N_15538);
or U16653 (N_16653,N_15952,N_15377);
nand U16654 (N_16654,N_15098,N_15807);
or U16655 (N_16655,N_15017,N_15515);
xor U16656 (N_16656,N_15306,N_15114);
and U16657 (N_16657,N_15540,N_15666);
nor U16658 (N_16658,N_15057,N_15085);
and U16659 (N_16659,N_15952,N_15103);
nor U16660 (N_16660,N_15030,N_15241);
and U16661 (N_16661,N_15112,N_15655);
xor U16662 (N_16662,N_15877,N_15586);
nor U16663 (N_16663,N_15959,N_15141);
or U16664 (N_16664,N_15469,N_15654);
and U16665 (N_16665,N_15934,N_15865);
nand U16666 (N_16666,N_15500,N_15414);
and U16667 (N_16667,N_15171,N_15027);
nor U16668 (N_16668,N_15751,N_15892);
nand U16669 (N_16669,N_15222,N_15172);
or U16670 (N_16670,N_15421,N_15531);
xnor U16671 (N_16671,N_15867,N_15881);
nor U16672 (N_16672,N_15314,N_15817);
nand U16673 (N_16673,N_15988,N_15552);
and U16674 (N_16674,N_15916,N_15722);
or U16675 (N_16675,N_15071,N_15036);
and U16676 (N_16676,N_15804,N_15949);
nand U16677 (N_16677,N_15036,N_15280);
nand U16678 (N_16678,N_15584,N_15799);
xnor U16679 (N_16679,N_15447,N_15802);
and U16680 (N_16680,N_15624,N_15079);
nor U16681 (N_16681,N_15636,N_15699);
xor U16682 (N_16682,N_15204,N_15750);
and U16683 (N_16683,N_15664,N_15913);
nand U16684 (N_16684,N_15081,N_15610);
or U16685 (N_16685,N_15161,N_15718);
or U16686 (N_16686,N_15395,N_15034);
xnor U16687 (N_16687,N_15295,N_15326);
xnor U16688 (N_16688,N_15511,N_15659);
or U16689 (N_16689,N_15669,N_15014);
or U16690 (N_16690,N_15048,N_15955);
or U16691 (N_16691,N_15293,N_15369);
and U16692 (N_16692,N_15685,N_15669);
nand U16693 (N_16693,N_15879,N_15645);
nor U16694 (N_16694,N_15762,N_15508);
nor U16695 (N_16695,N_15111,N_15785);
or U16696 (N_16696,N_15731,N_15259);
or U16697 (N_16697,N_15433,N_15362);
xor U16698 (N_16698,N_15460,N_15301);
and U16699 (N_16699,N_15509,N_15003);
xor U16700 (N_16700,N_15976,N_15853);
nand U16701 (N_16701,N_15531,N_15527);
or U16702 (N_16702,N_15542,N_15724);
xor U16703 (N_16703,N_15142,N_15459);
xnor U16704 (N_16704,N_15443,N_15264);
nor U16705 (N_16705,N_15150,N_15587);
or U16706 (N_16706,N_15763,N_15233);
xor U16707 (N_16707,N_15115,N_15378);
xnor U16708 (N_16708,N_15704,N_15954);
nand U16709 (N_16709,N_15896,N_15850);
and U16710 (N_16710,N_15977,N_15149);
or U16711 (N_16711,N_15193,N_15617);
nand U16712 (N_16712,N_15522,N_15694);
or U16713 (N_16713,N_15934,N_15659);
xor U16714 (N_16714,N_15058,N_15999);
nand U16715 (N_16715,N_15731,N_15434);
nor U16716 (N_16716,N_15073,N_15442);
and U16717 (N_16717,N_15164,N_15736);
nor U16718 (N_16718,N_15182,N_15406);
and U16719 (N_16719,N_15419,N_15130);
and U16720 (N_16720,N_15839,N_15862);
xnor U16721 (N_16721,N_15918,N_15377);
and U16722 (N_16722,N_15699,N_15530);
xor U16723 (N_16723,N_15725,N_15151);
and U16724 (N_16724,N_15143,N_15810);
nand U16725 (N_16725,N_15560,N_15702);
or U16726 (N_16726,N_15119,N_15208);
nor U16727 (N_16727,N_15556,N_15837);
nand U16728 (N_16728,N_15411,N_15304);
xor U16729 (N_16729,N_15052,N_15499);
nor U16730 (N_16730,N_15830,N_15065);
and U16731 (N_16731,N_15463,N_15923);
nor U16732 (N_16732,N_15624,N_15648);
nand U16733 (N_16733,N_15574,N_15248);
xnor U16734 (N_16734,N_15946,N_15701);
nor U16735 (N_16735,N_15459,N_15037);
xor U16736 (N_16736,N_15119,N_15329);
and U16737 (N_16737,N_15361,N_15206);
nor U16738 (N_16738,N_15896,N_15432);
nand U16739 (N_16739,N_15726,N_15912);
or U16740 (N_16740,N_15008,N_15768);
and U16741 (N_16741,N_15457,N_15205);
and U16742 (N_16742,N_15158,N_15212);
and U16743 (N_16743,N_15196,N_15302);
and U16744 (N_16744,N_15425,N_15726);
nand U16745 (N_16745,N_15754,N_15217);
nand U16746 (N_16746,N_15054,N_15155);
and U16747 (N_16747,N_15393,N_15953);
xnor U16748 (N_16748,N_15500,N_15083);
nand U16749 (N_16749,N_15734,N_15732);
xnor U16750 (N_16750,N_15006,N_15963);
nor U16751 (N_16751,N_15543,N_15441);
nor U16752 (N_16752,N_15824,N_15010);
nand U16753 (N_16753,N_15578,N_15089);
nand U16754 (N_16754,N_15373,N_15848);
or U16755 (N_16755,N_15386,N_15775);
and U16756 (N_16756,N_15001,N_15034);
or U16757 (N_16757,N_15062,N_15040);
and U16758 (N_16758,N_15270,N_15067);
and U16759 (N_16759,N_15997,N_15059);
nand U16760 (N_16760,N_15496,N_15854);
or U16761 (N_16761,N_15066,N_15314);
and U16762 (N_16762,N_15407,N_15952);
and U16763 (N_16763,N_15258,N_15383);
nor U16764 (N_16764,N_15632,N_15031);
nor U16765 (N_16765,N_15341,N_15303);
nand U16766 (N_16766,N_15826,N_15391);
or U16767 (N_16767,N_15667,N_15668);
and U16768 (N_16768,N_15754,N_15979);
nor U16769 (N_16769,N_15427,N_15598);
and U16770 (N_16770,N_15192,N_15464);
nand U16771 (N_16771,N_15038,N_15848);
nor U16772 (N_16772,N_15726,N_15528);
and U16773 (N_16773,N_15255,N_15394);
xnor U16774 (N_16774,N_15490,N_15099);
nor U16775 (N_16775,N_15823,N_15736);
nand U16776 (N_16776,N_15141,N_15552);
nand U16777 (N_16777,N_15620,N_15794);
or U16778 (N_16778,N_15741,N_15911);
xnor U16779 (N_16779,N_15775,N_15536);
or U16780 (N_16780,N_15559,N_15119);
xnor U16781 (N_16781,N_15482,N_15733);
or U16782 (N_16782,N_15840,N_15620);
nor U16783 (N_16783,N_15713,N_15446);
xnor U16784 (N_16784,N_15477,N_15856);
and U16785 (N_16785,N_15212,N_15130);
nand U16786 (N_16786,N_15550,N_15507);
nand U16787 (N_16787,N_15224,N_15585);
nand U16788 (N_16788,N_15472,N_15891);
nor U16789 (N_16789,N_15183,N_15585);
xnor U16790 (N_16790,N_15771,N_15937);
or U16791 (N_16791,N_15591,N_15204);
xor U16792 (N_16792,N_15390,N_15536);
xnor U16793 (N_16793,N_15680,N_15625);
nor U16794 (N_16794,N_15297,N_15377);
xnor U16795 (N_16795,N_15261,N_15832);
xor U16796 (N_16796,N_15996,N_15249);
xor U16797 (N_16797,N_15145,N_15472);
or U16798 (N_16798,N_15045,N_15583);
nand U16799 (N_16799,N_15115,N_15862);
nor U16800 (N_16800,N_15576,N_15634);
or U16801 (N_16801,N_15802,N_15329);
nor U16802 (N_16802,N_15596,N_15867);
or U16803 (N_16803,N_15910,N_15592);
xor U16804 (N_16804,N_15965,N_15605);
and U16805 (N_16805,N_15434,N_15076);
xnor U16806 (N_16806,N_15660,N_15246);
and U16807 (N_16807,N_15055,N_15256);
and U16808 (N_16808,N_15825,N_15826);
nor U16809 (N_16809,N_15007,N_15578);
or U16810 (N_16810,N_15012,N_15590);
and U16811 (N_16811,N_15357,N_15076);
xor U16812 (N_16812,N_15691,N_15879);
or U16813 (N_16813,N_15784,N_15144);
and U16814 (N_16814,N_15404,N_15763);
or U16815 (N_16815,N_15981,N_15685);
and U16816 (N_16816,N_15504,N_15202);
nand U16817 (N_16817,N_15985,N_15329);
or U16818 (N_16818,N_15037,N_15125);
nor U16819 (N_16819,N_15400,N_15137);
nand U16820 (N_16820,N_15338,N_15105);
and U16821 (N_16821,N_15760,N_15923);
nor U16822 (N_16822,N_15531,N_15235);
and U16823 (N_16823,N_15324,N_15507);
nand U16824 (N_16824,N_15019,N_15244);
and U16825 (N_16825,N_15515,N_15706);
xnor U16826 (N_16826,N_15642,N_15009);
nor U16827 (N_16827,N_15052,N_15728);
and U16828 (N_16828,N_15282,N_15733);
and U16829 (N_16829,N_15379,N_15666);
nor U16830 (N_16830,N_15743,N_15281);
nor U16831 (N_16831,N_15428,N_15676);
and U16832 (N_16832,N_15335,N_15311);
nor U16833 (N_16833,N_15755,N_15312);
nand U16834 (N_16834,N_15737,N_15418);
nand U16835 (N_16835,N_15246,N_15365);
nor U16836 (N_16836,N_15224,N_15658);
or U16837 (N_16837,N_15012,N_15478);
or U16838 (N_16838,N_15736,N_15364);
or U16839 (N_16839,N_15612,N_15137);
or U16840 (N_16840,N_15327,N_15541);
or U16841 (N_16841,N_15613,N_15530);
or U16842 (N_16842,N_15575,N_15088);
or U16843 (N_16843,N_15073,N_15826);
and U16844 (N_16844,N_15962,N_15481);
nor U16845 (N_16845,N_15489,N_15065);
and U16846 (N_16846,N_15460,N_15296);
nor U16847 (N_16847,N_15129,N_15931);
nand U16848 (N_16848,N_15969,N_15619);
xnor U16849 (N_16849,N_15674,N_15390);
or U16850 (N_16850,N_15845,N_15319);
xor U16851 (N_16851,N_15888,N_15423);
and U16852 (N_16852,N_15283,N_15223);
and U16853 (N_16853,N_15805,N_15168);
and U16854 (N_16854,N_15741,N_15669);
nand U16855 (N_16855,N_15982,N_15285);
nor U16856 (N_16856,N_15761,N_15573);
xor U16857 (N_16857,N_15851,N_15778);
xnor U16858 (N_16858,N_15016,N_15306);
xnor U16859 (N_16859,N_15411,N_15557);
nand U16860 (N_16860,N_15732,N_15295);
nor U16861 (N_16861,N_15477,N_15487);
nor U16862 (N_16862,N_15192,N_15037);
or U16863 (N_16863,N_15097,N_15346);
nand U16864 (N_16864,N_15156,N_15889);
nand U16865 (N_16865,N_15268,N_15455);
nor U16866 (N_16866,N_15604,N_15395);
or U16867 (N_16867,N_15140,N_15172);
xor U16868 (N_16868,N_15279,N_15170);
or U16869 (N_16869,N_15542,N_15653);
xor U16870 (N_16870,N_15027,N_15301);
or U16871 (N_16871,N_15033,N_15336);
or U16872 (N_16872,N_15644,N_15195);
and U16873 (N_16873,N_15048,N_15248);
or U16874 (N_16874,N_15674,N_15223);
xor U16875 (N_16875,N_15003,N_15683);
or U16876 (N_16876,N_15555,N_15324);
nor U16877 (N_16877,N_15885,N_15084);
nor U16878 (N_16878,N_15350,N_15227);
and U16879 (N_16879,N_15451,N_15143);
xnor U16880 (N_16880,N_15574,N_15715);
and U16881 (N_16881,N_15336,N_15928);
or U16882 (N_16882,N_15948,N_15466);
and U16883 (N_16883,N_15606,N_15482);
nor U16884 (N_16884,N_15918,N_15072);
or U16885 (N_16885,N_15274,N_15446);
nor U16886 (N_16886,N_15647,N_15485);
or U16887 (N_16887,N_15523,N_15765);
nand U16888 (N_16888,N_15190,N_15927);
nand U16889 (N_16889,N_15949,N_15788);
or U16890 (N_16890,N_15767,N_15019);
nor U16891 (N_16891,N_15848,N_15546);
nand U16892 (N_16892,N_15110,N_15691);
or U16893 (N_16893,N_15305,N_15509);
xnor U16894 (N_16894,N_15221,N_15761);
nor U16895 (N_16895,N_15956,N_15543);
or U16896 (N_16896,N_15189,N_15534);
or U16897 (N_16897,N_15331,N_15731);
nor U16898 (N_16898,N_15482,N_15320);
xor U16899 (N_16899,N_15400,N_15447);
and U16900 (N_16900,N_15512,N_15701);
nand U16901 (N_16901,N_15692,N_15407);
and U16902 (N_16902,N_15082,N_15208);
nor U16903 (N_16903,N_15616,N_15652);
and U16904 (N_16904,N_15026,N_15832);
and U16905 (N_16905,N_15200,N_15112);
or U16906 (N_16906,N_15203,N_15624);
nor U16907 (N_16907,N_15303,N_15028);
and U16908 (N_16908,N_15418,N_15525);
and U16909 (N_16909,N_15934,N_15211);
xnor U16910 (N_16910,N_15793,N_15957);
nor U16911 (N_16911,N_15195,N_15849);
or U16912 (N_16912,N_15266,N_15542);
or U16913 (N_16913,N_15567,N_15139);
or U16914 (N_16914,N_15152,N_15077);
and U16915 (N_16915,N_15523,N_15239);
xor U16916 (N_16916,N_15958,N_15433);
xnor U16917 (N_16917,N_15360,N_15586);
or U16918 (N_16918,N_15469,N_15548);
nor U16919 (N_16919,N_15707,N_15571);
nand U16920 (N_16920,N_15185,N_15741);
or U16921 (N_16921,N_15855,N_15868);
xnor U16922 (N_16922,N_15656,N_15477);
nand U16923 (N_16923,N_15102,N_15314);
nand U16924 (N_16924,N_15754,N_15074);
nand U16925 (N_16925,N_15332,N_15559);
nor U16926 (N_16926,N_15483,N_15517);
nand U16927 (N_16927,N_15037,N_15154);
and U16928 (N_16928,N_15697,N_15621);
nor U16929 (N_16929,N_15397,N_15864);
nor U16930 (N_16930,N_15679,N_15129);
and U16931 (N_16931,N_15964,N_15149);
or U16932 (N_16932,N_15981,N_15187);
nor U16933 (N_16933,N_15046,N_15448);
or U16934 (N_16934,N_15288,N_15033);
nor U16935 (N_16935,N_15659,N_15701);
nand U16936 (N_16936,N_15527,N_15283);
nor U16937 (N_16937,N_15471,N_15085);
and U16938 (N_16938,N_15867,N_15990);
and U16939 (N_16939,N_15494,N_15389);
or U16940 (N_16940,N_15629,N_15868);
nand U16941 (N_16941,N_15446,N_15543);
and U16942 (N_16942,N_15257,N_15618);
xor U16943 (N_16943,N_15082,N_15423);
nand U16944 (N_16944,N_15924,N_15381);
nor U16945 (N_16945,N_15866,N_15268);
nand U16946 (N_16946,N_15193,N_15619);
or U16947 (N_16947,N_15673,N_15640);
xnor U16948 (N_16948,N_15520,N_15535);
and U16949 (N_16949,N_15882,N_15858);
nand U16950 (N_16950,N_15293,N_15332);
nor U16951 (N_16951,N_15848,N_15610);
or U16952 (N_16952,N_15597,N_15027);
xor U16953 (N_16953,N_15866,N_15393);
and U16954 (N_16954,N_15034,N_15218);
or U16955 (N_16955,N_15208,N_15057);
nand U16956 (N_16956,N_15307,N_15040);
xor U16957 (N_16957,N_15897,N_15011);
nor U16958 (N_16958,N_15565,N_15601);
nand U16959 (N_16959,N_15285,N_15842);
and U16960 (N_16960,N_15762,N_15751);
nor U16961 (N_16961,N_15512,N_15400);
and U16962 (N_16962,N_15374,N_15631);
nand U16963 (N_16963,N_15533,N_15403);
nor U16964 (N_16964,N_15547,N_15892);
or U16965 (N_16965,N_15300,N_15697);
or U16966 (N_16966,N_15198,N_15151);
nor U16967 (N_16967,N_15324,N_15079);
and U16968 (N_16968,N_15161,N_15501);
nand U16969 (N_16969,N_15459,N_15234);
or U16970 (N_16970,N_15770,N_15099);
nand U16971 (N_16971,N_15462,N_15198);
nor U16972 (N_16972,N_15901,N_15225);
and U16973 (N_16973,N_15832,N_15126);
nand U16974 (N_16974,N_15048,N_15729);
xor U16975 (N_16975,N_15153,N_15387);
and U16976 (N_16976,N_15472,N_15901);
nor U16977 (N_16977,N_15637,N_15278);
nand U16978 (N_16978,N_15966,N_15366);
nand U16979 (N_16979,N_15227,N_15856);
nand U16980 (N_16980,N_15671,N_15120);
nor U16981 (N_16981,N_15986,N_15069);
and U16982 (N_16982,N_15364,N_15049);
nand U16983 (N_16983,N_15240,N_15934);
or U16984 (N_16984,N_15846,N_15230);
and U16985 (N_16985,N_15938,N_15285);
nor U16986 (N_16986,N_15907,N_15067);
or U16987 (N_16987,N_15286,N_15869);
nor U16988 (N_16988,N_15742,N_15211);
xnor U16989 (N_16989,N_15094,N_15386);
xnor U16990 (N_16990,N_15695,N_15785);
xnor U16991 (N_16991,N_15742,N_15192);
xor U16992 (N_16992,N_15975,N_15795);
or U16993 (N_16993,N_15530,N_15431);
xnor U16994 (N_16994,N_15375,N_15884);
or U16995 (N_16995,N_15324,N_15660);
nand U16996 (N_16996,N_15974,N_15991);
nor U16997 (N_16997,N_15038,N_15674);
and U16998 (N_16998,N_15019,N_15359);
or U16999 (N_16999,N_15448,N_15973);
nor U17000 (N_17000,N_16908,N_16819);
nand U17001 (N_17001,N_16031,N_16496);
nor U17002 (N_17002,N_16915,N_16884);
nor U17003 (N_17003,N_16696,N_16733);
nor U17004 (N_17004,N_16038,N_16864);
or U17005 (N_17005,N_16875,N_16162);
and U17006 (N_17006,N_16593,N_16928);
nand U17007 (N_17007,N_16887,N_16486);
and U17008 (N_17008,N_16353,N_16188);
or U17009 (N_17009,N_16872,N_16158);
nor U17010 (N_17010,N_16754,N_16848);
xnor U17011 (N_17011,N_16983,N_16902);
nor U17012 (N_17012,N_16351,N_16451);
nor U17013 (N_17013,N_16361,N_16005);
nor U17014 (N_17014,N_16044,N_16316);
or U17015 (N_17015,N_16524,N_16610);
nor U17016 (N_17016,N_16366,N_16438);
nand U17017 (N_17017,N_16342,N_16512);
and U17018 (N_17018,N_16133,N_16258);
or U17019 (N_17019,N_16203,N_16926);
nor U17020 (N_17020,N_16103,N_16963);
nand U17021 (N_17021,N_16781,N_16552);
or U17022 (N_17022,N_16629,N_16426);
and U17023 (N_17023,N_16738,N_16533);
xor U17024 (N_17024,N_16084,N_16731);
and U17025 (N_17025,N_16171,N_16198);
or U17026 (N_17026,N_16125,N_16013);
nor U17027 (N_17027,N_16907,N_16692);
or U17028 (N_17028,N_16228,N_16276);
xor U17029 (N_17029,N_16183,N_16235);
nand U17030 (N_17030,N_16446,N_16889);
nor U17031 (N_17031,N_16626,N_16530);
nor U17032 (N_17032,N_16097,N_16663);
and U17033 (N_17033,N_16018,N_16197);
xor U17034 (N_17034,N_16566,N_16893);
or U17035 (N_17035,N_16580,N_16355);
and U17036 (N_17036,N_16615,N_16665);
or U17037 (N_17037,N_16664,N_16861);
nand U17038 (N_17038,N_16204,N_16271);
or U17039 (N_17039,N_16888,N_16348);
xnor U17040 (N_17040,N_16151,N_16093);
or U17041 (N_17041,N_16064,N_16740);
xor U17042 (N_17042,N_16784,N_16466);
nand U17043 (N_17043,N_16360,N_16009);
or U17044 (N_17044,N_16489,N_16949);
xnor U17045 (N_17045,N_16409,N_16955);
nor U17046 (N_17046,N_16972,N_16840);
nor U17047 (N_17047,N_16106,N_16225);
or U17048 (N_17048,N_16761,N_16930);
nor U17049 (N_17049,N_16620,N_16985);
nor U17050 (N_17050,N_16283,N_16645);
nor U17051 (N_17051,N_16898,N_16567);
or U17052 (N_17052,N_16801,N_16677);
nand U17053 (N_17053,N_16913,N_16500);
nor U17054 (N_17054,N_16613,N_16901);
and U17055 (N_17055,N_16790,N_16384);
nand U17056 (N_17056,N_16541,N_16497);
and U17057 (N_17057,N_16614,N_16783);
and U17058 (N_17058,N_16518,N_16722);
xnor U17059 (N_17059,N_16660,N_16027);
nor U17060 (N_17060,N_16358,N_16558);
nor U17061 (N_17061,N_16286,N_16473);
nand U17062 (N_17062,N_16788,N_16357);
or U17063 (N_17063,N_16549,N_16433);
or U17064 (N_17064,N_16394,N_16818);
or U17065 (N_17065,N_16595,N_16229);
nand U17066 (N_17066,N_16914,N_16135);
nand U17067 (N_17067,N_16362,N_16751);
xnor U17068 (N_17068,N_16467,N_16363);
xor U17069 (N_17069,N_16508,N_16432);
nor U17070 (N_17070,N_16092,N_16445);
xor U17071 (N_17071,N_16643,N_16220);
or U17072 (N_17072,N_16634,N_16756);
nor U17073 (N_17073,N_16759,N_16159);
xnor U17074 (N_17074,N_16318,N_16107);
or U17075 (N_17075,N_16123,N_16155);
nand U17076 (N_17076,N_16701,N_16846);
and U17077 (N_17077,N_16042,N_16002);
xor U17078 (N_17078,N_16623,N_16544);
xnor U17079 (N_17079,N_16332,N_16628);
xnor U17080 (N_17080,N_16839,N_16128);
and U17081 (N_17081,N_16873,N_16215);
and U17082 (N_17082,N_16718,N_16705);
or U17083 (N_17083,N_16310,N_16447);
nand U17084 (N_17084,N_16837,N_16014);
xor U17085 (N_17085,N_16841,N_16509);
or U17086 (N_17086,N_16369,N_16545);
nand U17087 (N_17087,N_16116,N_16279);
xnor U17088 (N_17088,N_16862,N_16134);
nor U17089 (N_17089,N_16689,N_16410);
or U17090 (N_17090,N_16959,N_16216);
xnor U17091 (N_17091,N_16789,N_16295);
and U17092 (N_17092,N_16737,N_16618);
xor U17093 (N_17093,N_16745,N_16205);
nor U17094 (N_17094,N_16559,N_16821);
xor U17095 (N_17095,N_16883,N_16562);
nor U17096 (N_17096,N_16870,N_16658);
and U17097 (N_17097,N_16556,N_16146);
nand U17098 (N_17098,N_16047,N_16523);
nand U17099 (N_17099,N_16016,N_16569);
xor U17100 (N_17100,N_16234,N_16494);
xor U17101 (N_17101,N_16655,N_16023);
and U17102 (N_17102,N_16323,N_16944);
nand U17103 (N_17103,N_16961,N_16498);
and U17104 (N_17104,N_16108,N_16417);
and U17105 (N_17105,N_16505,N_16603);
xnor U17106 (N_17106,N_16314,N_16322);
nor U17107 (N_17107,N_16670,N_16101);
nor U17108 (N_17108,N_16163,N_16194);
and U17109 (N_17109,N_16117,N_16504);
nand U17110 (N_17110,N_16189,N_16397);
or U17111 (N_17111,N_16966,N_16997);
or U17112 (N_17112,N_16390,N_16906);
nand U17113 (N_17113,N_16817,N_16709);
xnor U17114 (N_17114,N_16441,N_16806);
nand U17115 (N_17115,N_16828,N_16695);
xnor U17116 (N_17116,N_16430,N_16130);
xnor U17117 (N_17117,N_16999,N_16049);
or U17118 (N_17118,N_16771,N_16777);
or U17119 (N_17119,N_16086,N_16024);
and U17120 (N_17120,N_16510,N_16034);
xor U17121 (N_17121,N_16903,N_16578);
or U17122 (N_17122,N_16482,N_16631);
or U17123 (N_17123,N_16551,N_16379);
and U17124 (N_17124,N_16401,N_16844);
and U17125 (N_17125,N_16589,N_16778);
nor U17126 (N_17126,N_16074,N_16109);
nand U17127 (N_17127,N_16293,N_16674);
nand U17128 (N_17128,N_16392,N_16240);
or U17129 (N_17129,N_16126,N_16327);
nand U17130 (N_17130,N_16406,N_16691);
nor U17131 (N_17131,N_16483,N_16706);
nand U17132 (N_17132,N_16909,N_16829);
nor U17133 (N_17133,N_16968,N_16742);
nand U17134 (N_17134,N_16780,N_16324);
or U17135 (N_17135,N_16904,N_16847);
or U17136 (N_17136,N_16054,N_16880);
xnor U17137 (N_17137,N_16448,N_16572);
nor U17138 (N_17138,N_16176,N_16824);
xor U17139 (N_17139,N_16585,N_16476);
and U17140 (N_17140,N_16395,N_16127);
nand U17141 (N_17141,N_16199,N_16779);
and U17142 (N_17142,N_16251,N_16319);
and U17143 (N_17143,N_16553,N_16536);
and U17144 (N_17144,N_16732,N_16259);
xnor U17145 (N_17145,N_16577,N_16192);
xor U17146 (N_17146,N_16265,N_16682);
and U17147 (N_17147,N_16814,N_16184);
nor U17148 (N_17148,N_16548,N_16795);
or U17149 (N_17149,N_16687,N_16803);
and U17150 (N_17150,N_16538,N_16953);
nor U17151 (N_17151,N_16081,N_16244);
or U17152 (N_17152,N_16343,N_16166);
and U17153 (N_17153,N_16517,N_16281);
nand U17154 (N_17154,N_16052,N_16377);
and U17155 (N_17155,N_16746,N_16338);
or U17156 (N_17156,N_16137,N_16493);
or U17157 (N_17157,N_16206,N_16799);
or U17158 (N_17158,N_16213,N_16651);
or U17159 (N_17159,N_16440,N_16762);
nor U17160 (N_17160,N_16036,N_16161);
nor U17161 (N_17161,N_16753,N_16833);
nand U17162 (N_17162,N_16444,N_16333);
nor U17163 (N_17163,N_16980,N_16245);
nor U17164 (N_17164,N_16879,N_16029);
xor U17165 (N_17165,N_16969,N_16532);
and U17166 (N_17166,N_16543,N_16481);
or U17167 (N_17167,N_16724,N_16954);
or U17168 (N_17168,N_16150,N_16739);
or U17169 (N_17169,N_16752,N_16082);
or U17170 (N_17170,N_16601,N_16942);
nand U17171 (N_17171,N_16380,N_16998);
and U17172 (N_17172,N_16630,N_16303);
xor U17173 (N_17173,N_16878,N_16227);
or U17174 (N_17174,N_16877,N_16698);
or U17175 (N_17175,N_16186,N_16419);
nand U17176 (N_17176,N_16748,N_16675);
xnor U17177 (N_17177,N_16713,N_16490);
nor U17178 (N_17178,N_16055,N_16897);
or U17179 (N_17179,N_16404,N_16564);
nand U17180 (N_17180,N_16237,N_16527);
nand U17181 (N_17181,N_16495,N_16511);
nand U17182 (N_17182,N_16113,N_16573);
nand U17183 (N_17183,N_16267,N_16871);
nand U17184 (N_17184,N_16347,N_16398);
xor U17185 (N_17185,N_16991,N_16937);
xnor U17186 (N_17186,N_16326,N_16480);
xnor U17187 (N_17187,N_16212,N_16669);
xor U17188 (N_17188,N_16934,N_16423);
nand U17189 (N_17189,N_16179,N_16951);
and U17190 (N_17190,N_16852,N_16672);
or U17191 (N_17191,N_16019,N_16911);
or U17192 (N_17192,N_16025,N_16656);
xnor U17193 (N_17193,N_16869,N_16078);
xnor U17194 (N_17194,N_16071,N_16411);
or U17195 (N_17195,N_16947,N_16020);
nand U17196 (N_17196,N_16579,N_16305);
or U17197 (N_17197,N_16121,N_16758);
xor U17198 (N_17198,N_16571,N_16767);
xor U17199 (N_17199,N_16400,N_16866);
or U17200 (N_17200,N_16238,N_16885);
xor U17201 (N_17201,N_16102,N_16975);
xnor U17202 (N_17202,N_16646,N_16375);
and U17203 (N_17203,N_16637,N_16749);
nor U17204 (N_17204,N_16300,N_16503);
or U17205 (N_17205,N_16600,N_16320);
xor U17206 (N_17206,N_16030,N_16041);
and U17207 (N_17207,N_16546,N_16252);
or U17208 (N_17208,N_16407,N_16261);
nor U17209 (N_17209,N_16588,N_16219);
and U17210 (N_17210,N_16098,N_16491);
and U17211 (N_17211,N_16960,N_16141);
and U17212 (N_17212,N_16597,N_16325);
or U17213 (N_17213,N_16195,N_16772);
nand U17214 (N_17214,N_16170,N_16138);
xor U17215 (N_17215,N_16568,N_16900);
nand U17216 (N_17216,N_16297,N_16415);
or U17217 (N_17217,N_16680,N_16831);
xor U17218 (N_17218,N_16574,N_16590);
xor U17219 (N_17219,N_16033,N_16273);
nor U17220 (N_17220,N_16609,N_16515);
and U17221 (N_17221,N_16987,N_16091);
or U17222 (N_17222,N_16442,N_16557);
or U17223 (N_17223,N_16439,N_16717);
xnor U17224 (N_17224,N_16714,N_16173);
and U17225 (N_17225,N_16269,N_16797);
and U17226 (N_17226,N_16344,N_16886);
xnor U17227 (N_17227,N_16399,N_16932);
and U17228 (N_17228,N_16927,N_16461);
nor U17229 (N_17229,N_16272,N_16858);
or U17230 (N_17230,N_16266,N_16214);
or U17231 (N_17231,N_16187,N_16825);
xor U17232 (N_17232,N_16067,N_16422);
or U17233 (N_17233,N_16863,N_16096);
or U17234 (N_17234,N_16690,N_16529);
nor U17235 (N_17235,N_16891,N_16456);
xor U17236 (N_17236,N_16586,N_16012);
xor U17237 (N_17237,N_16925,N_16037);
xor U17238 (N_17238,N_16736,N_16154);
nand U17239 (N_17239,N_16140,N_16584);
xor U17240 (N_17240,N_16750,N_16337);
nor U17241 (N_17241,N_16607,N_16153);
or U17242 (N_17242,N_16662,N_16611);
nor U17243 (N_17243,N_16475,N_16519);
nor U17244 (N_17244,N_16434,N_16356);
nor U17245 (N_17245,N_16413,N_16167);
or U17246 (N_17246,N_16899,N_16405);
nand U17247 (N_17247,N_16554,N_16633);
xor U17248 (N_17248,N_16624,N_16436);
or U17249 (N_17249,N_16382,N_16367);
nor U17250 (N_17250,N_16652,N_16522);
or U17251 (N_17251,N_16421,N_16056);
xor U17252 (N_17252,N_16474,N_16791);
nand U17253 (N_17253,N_16068,N_16807);
xor U17254 (N_17254,N_16851,N_16144);
and U17255 (N_17255,N_16874,N_16370);
nand U17256 (N_17256,N_16372,N_16956);
nand U17257 (N_17257,N_16804,N_16542);
xnor U17258 (N_17258,N_16798,N_16472);
nand U17259 (N_17259,N_16428,N_16022);
nor U17260 (N_17260,N_16565,N_16301);
or U17261 (N_17261,N_16936,N_16231);
and U17262 (N_17262,N_16015,N_16371);
xor U17263 (N_17263,N_16119,N_16485);
or U17264 (N_17264,N_16262,N_16946);
nor U17265 (N_17265,N_16492,N_16711);
nand U17266 (N_17266,N_16180,N_16335);
nand U17267 (N_17267,N_16260,N_16006);
and U17268 (N_17268,N_16003,N_16191);
or U17269 (N_17269,N_16792,N_16311);
nor U17270 (N_17270,N_16115,N_16182);
and U17271 (N_17271,N_16350,N_16149);
nor U17272 (N_17272,N_16986,N_16604);
nor U17273 (N_17273,N_16264,N_16061);
and U17274 (N_17274,N_16349,N_16994);
and U17275 (N_17275,N_16051,N_16704);
nand U17276 (N_17276,N_16805,N_16834);
and U17277 (N_17277,N_16378,N_16827);
or U17278 (N_17278,N_16217,N_16919);
nor U17279 (N_17279,N_16059,N_16592);
or U17280 (N_17280,N_16977,N_16118);
nand U17281 (N_17281,N_16339,N_16521);
or U17282 (N_17282,N_16826,N_16550);
or U17283 (N_17283,N_16881,N_16948);
or U17284 (N_17284,N_16010,N_16274);
nand U17285 (N_17285,N_16331,N_16035);
nand U17286 (N_17286,N_16796,N_16707);
nor U17287 (N_17287,N_16243,N_16328);
and U17288 (N_17288,N_16688,N_16679);
nor U17289 (N_17289,N_16666,N_16894);
xor U17290 (N_17290,N_16905,N_16974);
nand U17291 (N_17291,N_16516,N_16028);
and U17292 (N_17292,N_16450,N_16254);
nor U17293 (N_17293,N_16471,N_16703);
nor U17294 (N_17294,N_16278,N_16226);
nand U17295 (N_17295,N_16224,N_16683);
and U17296 (N_17296,N_16810,N_16315);
and U17297 (N_17297,N_16685,N_16636);
or U17298 (N_17298,N_16202,N_16429);
and U17299 (N_17299,N_16210,N_16768);
nand U17300 (N_17300,N_16488,N_16032);
nand U17301 (N_17301,N_16285,N_16336);
and U17302 (N_17302,N_16385,N_16001);
nor U17303 (N_17303,N_16236,N_16459);
or U17304 (N_17304,N_16329,N_16793);
nor U17305 (N_17305,N_16304,N_16287);
or U17306 (N_17306,N_16060,N_16594);
nor U17307 (N_17307,N_16587,N_16280);
xor U17308 (N_17308,N_16063,N_16599);
nand U17309 (N_17309,N_16616,N_16513);
nand U17310 (N_17310,N_16843,N_16352);
xnor U17311 (N_17311,N_16867,N_16723);
nand U17312 (N_17312,N_16995,N_16648);
nand U17313 (N_17313,N_16935,N_16321);
xor U17314 (N_17314,N_16940,N_16290);
or U17315 (N_17315,N_16653,N_16976);
nor U17316 (N_17316,N_16555,N_16386);
nor U17317 (N_17317,N_16835,N_16921);
and U17318 (N_17318,N_16850,N_16922);
nand U17319 (N_17319,N_16437,N_16952);
nand U17320 (N_17320,N_16988,N_16563);
nand U17321 (N_17321,N_16085,N_16561);
xor U17322 (N_17322,N_16933,N_16642);
and U17323 (N_17323,N_16916,N_16465);
and U17324 (N_17324,N_16143,N_16598);
and U17325 (N_17325,N_16918,N_16431);
or U17326 (N_17326,N_16857,N_16910);
xnor U17327 (N_17327,N_16292,N_16105);
and U17328 (N_17328,N_16070,N_16782);
nor U17329 (N_17329,N_16537,N_16077);
nand U17330 (N_17330,N_16499,N_16172);
or U17331 (N_17331,N_16979,N_16619);
nand U17332 (N_17332,N_16268,N_16712);
and U17333 (N_17333,N_16196,N_16147);
and U17334 (N_17334,N_16139,N_16640);
and U17335 (N_17335,N_16958,N_16345);
xor U17336 (N_17336,N_16697,N_16945);
nand U17337 (N_17337,N_16816,N_16414);
and U17338 (N_17338,N_16452,N_16207);
nand U17339 (N_17339,N_16288,N_16506);
or U17340 (N_17340,N_16160,N_16865);
nand U17341 (N_17341,N_16800,N_16168);
and U17342 (N_17342,N_16809,N_16741);
or U17343 (N_17343,N_16306,N_16298);
xnor U17344 (N_17344,N_16247,N_16787);
nor U17345 (N_17345,N_16760,N_16747);
nor U17346 (N_17346,N_16811,N_16755);
nand U17347 (N_17347,N_16175,N_16514);
nand U17348 (N_17348,N_16868,N_16836);
or U17349 (N_17349,N_16993,N_16686);
or U17350 (N_17350,N_16221,N_16403);
xnor U17351 (N_17351,N_16608,N_16313);
xnor U17352 (N_17352,N_16291,N_16560);
or U17353 (N_17353,N_16941,N_16849);
xor U17354 (N_17354,N_16725,N_16896);
xor U17355 (N_17355,N_16764,N_16726);
nor U17356 (N_17356,N_16769,N_16455);
nand U17357 (N_17357,N_16094,N_16309);
xnor U17358 (N_17358,N_16981,N_16334);
and U17359 (N_17359,N_16647,N_16045);
and U17360 (N_17360,N_16469,N_16046);
xor U17361 (N_17361,N_16470,N_16062);
nand U17362 (N_17362,N_16924,N_16808);
or U17363 (N_17363,N_16853,N_16222);
and U17364 (N_17364,N_16520,N_16164);
nor U17365 (N_17365,N_16729,N_16124);
nor U17366 (N_17366,N_16962,N_16088);
xnor U17367 (N_17367,N_16699,N_16007);
nor U17368 (N_17368,N_16275,N_16131);
xnor U17369 (N_17369,N_16057,N_16364);
nor U17370 (N_17370,N_16970,N_16462);
or U17371 (N_17371,N_16678,N_16122);
nor U17372 (N_17372,N_16635,N_16708);
and U17373 (N_17373,N_16048,N_16190);
and U17374 (N_17374,N_16720,N_16408);
nand U17375 (N_17375,N_16734,N_16876);
xnor U17376 (N_17376,N_16823,N_16458);
nor U17377 (N_17377,N_16912,N_16487);
or U17378 (N_17378,N_16694,N_16359);
nor U17379 (N_17379,N_16786,N_16354);
or U17380 (N_17380,N_16069,N_16043);
xnor U17381 (N_17381,N_16744,N_16090);
xnor U17382 (N_17382,N_16632,N_16671);
xnor U17383 (N_17383,N_16727,N_16743);
or U17384 (N_17384,N_16710,N_16178);
or U17385 (N_17385,N_16895,N_16021);
nand U17386 (N_17386,N_16622,N_16528);
xnor U17387 (N_17387,N_16457,N_16242);
and U17388 (N_17388,N_16299,N_16453);
nor U17389 (N_17389,N_16539,N_16185);
and U17390 (N_17390,N_16661,N_16484);
xnor U17391 (N_17391,N_16340,N_16501);
xor U17392 (N_17392,N_16100,N_16882);
or U17393 (N_17393,N_16776,N_16250);
and U17394 (N_17394,N_16855,N_16802);
or U17395 (N_17395,N_16770,N_16065);
nand U17396 (N_17396,N_16388,N_16302);
xor U17397 (N_17397,N_16284,N_16965);
or U17398 (N_17398,N_16463,N_16950);
xnor U17399 (N_17399,N_16263,N_16531);
nand U17400 (N_17400,N_16230,N_16617);
or U17401 (N_17401,N_16464,N_16104);
xor U17402 (N_17402,N_16169,N_16087);
nor U17403 (N_17403,N_16971,N_16152);
nor U17404 (N_17404,N_16420,N_16076);
or U17405 (N_17405,N_16815,N_16612);
nor U17406 (N_17406,N_16606,N_16923);
nand U17407 (N_17407,N_16424,N_16765);
nor U17408 (N_17408,N_16794,N_16766);
nand U17409 (N_17409,N_16477,N_16289);
xnor U17410 (N_17410,N_16418,N_16657);
xnor U17411 (N_17411,N_16992,N_16650);
nor U17412 (N_17412,N_16050,N_16540);
nand U17413 (N_17413,N_16412,N_16943);
or U17414 (N_17414,N_16854,N_16040);
xor U17415 (N_17415,N_16095,N_16373);
or U17416 (N_17416,N_16639,N_16621);
nand U17417 (N_17417,N_16075,N_16365);
or U17418 (N_17418,N_16211,N_16547);
and U17419 (N_17419,N_16389,N_16233);
nand U17420 (N_17420,N_16860,N_16201);
xnor U17421 (N_17421,N_16938,N_16427);
or U17422 (N_17422,N_16066,N_16017);
and U17423 (N_17423,N_16193,N_16468);
and U17424 (N_17424,N_16341,N_16200);
nand U17425 (N_17425,N_16393,N_16253);
nor U17426 (N_17426,N_16218,N_16845);
or U17427 (N_17427,N_16110,N_16004);
or U17428 (N_17428,N_16376,N_16120);
and U17429 (N_17429,N_16581,N_16330);
or U17430 (N_17430,N_16443,N_16813);
nor U17431 (N_17431,N_16676,N_16307);
xnor U17432 (N_17432,N_16625,N_16693);
or U17433 (N_17433,N_16246,N_16239);
xor U17434 (N_17434,N_16856,N_16931);
nand U17435 (N_17435,N_16757,N_16255);
nor U17436 (N_17436,N_16990,N_16282);
nor U17437 (N_17437,N_16832,N_16728);
and U17438 (N_17438,N_16730,N_16502);
and U17439 (N_17439,N_16602,N_16920);
and U17440 (N_17440,N_16039,N_16374);
and U17441 (N_17441,N_16079,N_16241);
and U17442 (N_17442,N_16830,N_16576);
or U17443 (N_17443,N_16702,N_16526);
or U17444 (N_17444,N_16312,N_16391);
or U17445 (N_17445,N_16719,N_16774);
nand U17446 (N_17446,N_16454,N_16008);
xnor U17447 (N_17447,N_16989,N_16425);
nand U17448 (N_17448,N_16317,N_16684);
or U17449 (N_17449,N_16649,N_16416);
nor U17450 (N_17450,N_16248,N_16478);
nor U17451 (N_17451,N_16525,N_16256);
xor U17452 (N_17452,N_16381,N_16089);
nor U17453 (N_17453,N_16982,N_16929);
or U17454 (N_17454,N_16591,N_16296);
nand U17455 (N_17455,N_16308,N_16644);
and U17456 (N_17456,N_16681,N_16114);
nor U17457 (N_17457,N_16083,N_16939);
nand U17458 (N_17458,N_16072,N_16099);
nand U17459 (N_17459,N_16967,N_16638);
and U17460 (N_17460,N_16402,N_16249);
and U17461 (N_17461,N_16181,N_16346);
nand U17462 (N_17462,N_16583,N_16859);
and U17463 (N_17463,N_16842,N_16964);
or U17464 (N_17464,N_16368,N_16396);
nor U17465 (N_17465,N_16735,N_16890);
xnor U17466 (N_17466,N_16812,N_16984);
xnor U17467 (N_17467,N_16148,N_16387);
and U17468 (N_17468,N_16142,N_16177);
nor U17469 (N_17469,N_16570,N_16270);
or U17470 (N_17470,N_16080,N_16917);
nand U17471 (N_17471,N_16973,N_16145);
or U17472 (N_17472,N_16822,N_16763);
or U17473 (N_17473,N_16449,N_16654);
nand U17474 (N_17474,N_16715,N_16785);
and U17475 (N_17475,N_16535,N_16575);
nor U17476 (N_17476,N_16775,N_16129);
nor U17477 (N_17477,N_16058,N_16165);
or U17478 (N_17478,N_16460,N_16820);
nor U17479 (N_17479,N_16605,N_16136);
or U17480 (N_17480,N_16174,N_16208);
and U17481 (N_17481,N_16507,N_16957);
xnor U17482 (N_17482,N_16000,N_16667);
and U17483 (N_17483,N_16659,N_16383);
nor U17484 (N_17484,N_16534,N_16157);
nor U17485 (N_17485,N_16978,N_16892);
nand U17486 (N_17486,N_16700,N_16627);
nand U17487 (N_17487,N_16277,N_16721);
xor U17488 (N_17488,N_16294,N_16223);
or U17489 (N_17489,N_16668,N_16011);
nand U17490 (N_17490,N_16026,N_16132);
and U17491 (N_17491,N_16773,N_16112);
xnor U17492 (N_17492,N_16996,N_16257);
nand U17493 (N_17493,N_16156,N_16673);
or U17494 (N_17494,N_16073,N_16111);
and U17495 (N_17495,N_16838,N_16232);
xor U17496 (N_17496,N_16716,N_16435);
or U17497 (N_17497,N_16479,N_16582);
and U17498 (N_17498,N_16641,N_16209);
nor U17499 (N_17499,N_16053,N_16596);
or U17500 (N_17500,N_16516,N_16961);
xnor U17501 (N_17501,N_16161,N_16552);
and U17502 (N_17502,N_16641,N_16325);
nor U17503 (N_17503,N_16539,N_16689);
nor U17504 (N_17504,N_16385,N_16412);
nand U17505 (N_17505,N_16007,N_16166);
xnor U17506 (N_17506,N_16487,N_16921);
nor U17507 (N_17507,N_16788,N_16557);
and U17508 (N_17508,N_16048,N_16366);
or U17509 (N_17509,N_16587,N_16832);
and U17510 (N_17510,N_16144,N_16640);
nor U17511 (N_17511,N_16099,N_16344);
nand U17512 (N_17512,N_16538,N_16352);
nor U17513 (N_17513,N_16512,N_16033);
and U17514 (N_17514,N_16158,N_16129);
nor U17515 (N_17515,N_16449,N_16268);
nand U17516 (N_17516,N_16785,N_16350);
or U17517 (N_17517,N_16516,N_16080);
nor U17518 (N_17518,N_16225,N_16904);
or U17519 (N_17519,N_16589,N_16748);
xor U17520 (N_17520,N_16937,N_16645);
and U17521 (N_17521,N_16433,N_16550);
and U17522 (N_17522,N_16528,N_16890);
xnor U17523 (N_17523,N_16223,N_16867);
nor U17524 (N_17524,N_16070,N_16589);
nand U17525 (N_17525,N_16573,N_16175);
and U17526 (N_17526,N_16131,N_16881);
or U17527 (N_17527,N_16421,N_16169);
or U17528 (N_17528,N_16056,N_16235);
or U17529 (N_17529,N_16181,N_16740);
nor U17530 (N_17530,N_16447,N_16521);
and U17531 (N_17531,N_16041,N_16114);
xor U17532 (N_17532,N_16290,N_16690);
and U17533 (N_17533,N_16472,N_16949);
nor U17534 (N_17534,N_16471,N_16140);
xnor U17535 (N_17535,N_16613,N_16633);
or U17536 (N_17536,N_16649,N_16803);
and U17537 (N_17537,N_16931,N_16726);
and U17538 (N_17538,N_16749,N_16325);
nand U17539 (N_17539,N_16768,N_16247);
nor U17540 (N_17540,N_16538,N_16690);
xor U17541 (N_17541,N_16340,N_16306);
xor U17542 (N_17542,N_16295,N_16866);
and U17543 (N_17543,N_16037,N_16789);
or U17544 (N_17544,N_16780,N_16692);
or U17545 (N_17545,N_16909,N_16606);
nor U17546 (N_17546,N_16574,N_16811);
or U17547 (N_17547,N_16999,N_16247);
nand U17548 (N_17548,N_16050,N_16617);
and U17549 (N_17549,N_16919,N_16608);
nand U17550 (N_17550,N_16816,N_16064);
nor U17551 (N_17551,N_16650,N_16391);
xnor U17552 (N_17552,N_16525,N_16296);
nor U17553 (N_17553,N_16768,N_16925);
or U17554 (N_17554,N_16587,N_16013);
or U17555 (N_17555,N_16577,N_16415);
nor U17556 (N_17556,N_16097,N_16149);
nor U17557 (N_17557,N_16462,N_16327);
nand U17558 (N_17558,N_16196,N_16999);
xnor U17559 (N_17559,N_16443,N_16835);
and U17560 (N_17560,N_16996,N_16954);
and U17561 (N_17561,N_16958,N_16523);
or U17562 (N_17562,N_16156,N_16441);
xor U17563 (N_17563,N_16519,N_16912);
and U17564 (N_17564,N_16023,N_16657);
and U17565 (N_17565,N_16400,N_16274);
or U17566 (N_17566,N_16909,N_16921);
xor U17567 (N_17567,N_16590,N_16990);
and U17568 (N_17568,N_16072,N_16205);
xnor U17569 (N_17569,N_16601,N_16573);
xnor U17570 (N_17570,N_16525,N_16329);
or U17571 (N_17571,N_16886,N_16722);
and U17572 (N_17572,N_16778,N_16816);
nand U17573 (N_17573,N_16800,N_16668);
and U17574 (N_17574,N_16137,N_16427);
and U17575 (N_17575,N_16437,N_16286);
xor U17576 (N_17576,N_16909,N_16381);
or U17577 (N_17577,N_16580,N_16613);
xnor U17578 (N_17578,N_16565,N_16472);
xor U17579 (N_17579,N_16803,N_16439);
xor U17580 (N_17580,N_16683,N_16230);
nor U17581 (N_17581,N_16843,N_16164);
nand U17582 (N_17582,N_16502,N_16659);
nor U17583 (N_17583,N_16932,N_16014);
and U17584 (N_17584,N_16118,N_16924);
or U17585 (N_17585,N_16515,N_16412);
and U17586 (N_17586,N_16074,N_16652);
or U17587 (N_17587,N_16176,N_16136);
nand U17588 (N_17588,N_16913,N_16296);
xor U17589 (N_17589,N_16715,N_16070);
nor U17590 (N_17590,N_16369,N_16494);
nand U17591 (N_17591,N_16320,N_16120);
or U17592 (N_17592,N_16466,N_16276);
nor U17593 (N_17593,N_16190,N_16107);
nand U17594 (N_17594,N_16885,N_16511);
xor U17595 (N_17595,N_16269,N_16732);
xor U17596 (N_17596,N_16133,N_16641);
nand U17597 (N_17597,N_16567,N_16592);
xor U17598 (N_17598,N_16782,N_16405);
nor U17599 (N_17599,N_16062,N_16781);
nand U17600 (N_17600,N_16409,N_16166);
nor U17601 (N_17601,N_16747,N_16624);
nor U17602 (N_17602,N_16304,N_16960);
nor U17603 (N_17603,N_16443,N_16028);
nor U17604 (N_17604,N_16611,N_16506);
nor U17605 (N_17605,N_16855,N_16709);
and U17606 (N_17606,N_16512,N_16589);
and U17607 (N_17607,N_16335,N_16260);
or U17608 (N_17608,N_16080,N_16567);
nor U17609 (N_17609,N_16113,N_16630);
nor U17610 (N_17610,N_16003,N_16359);
and U17611 (N_17611,N_16075,N_16731);
xnor U17612 (N_17612,N_16157,N_16866);
and U17613 (N_17613,N_16986,N_16844);
nor U17614 (N_17614,N_16137,N_16731);
nor U17615 (N_17615,N_16678,N_16358);
or U17616 (N_17616,N_16635,N_16491);
or U17617 (N_17617,N_16424,N_16222);
nor U17618 (N_17618,N_16982,N_16758);
or U17619 (N_17619,N_16565,N_16416);
xnor U17620 (N_17620,N_16778,N_16649);
xnor U17621 (N_17621,N_16125,N_16681);
and U17622 (N_17622,N_16326,N_16672);
and U17623 (N_17623,N_16827,N_16794);
nor U17624 (N_17624,N_16949,N_16662);
or U17625 (N_17625,N_16965,N_16829);
and U17626 (N_17626,N_16269,N_16063);
nand U17627 (N_17627,N_16525,N_16369);
nor U17628 (N_17628,N_16531,N_16749);
and U17629 (N_17629,N_16474,N_16552);
nor U17630 (N_17630,N_16933,N_16445);
nor U17631 (N_17631,N_16099,N_16870);
or U17632 (N_17632,N_16834,N_16105);
or U17633 (N_17633,N_16462,N_16457);
nand U17634 (N_17634,N_16290,N_16644);
xnor U17635 (N_17635,N_16834,N_16134);
or U17636 (N_17636,N_16835,N_16673);
nand U17637 (N_17637,N_16077,N_16003);
nor U17638 (N_17638,N_16720,N_16341);
xnor U17639 (N_17639,N_16495,N_16659);
and U17640 (N_17640,N_16158,N_16505);
or U17641 (N_17641,N_16791,N_16531);
or U17642 (N_17642,N_16734,N_16297);
or U17643 (N_17643,N_16734,N_16293);
and U17644 (N_17644,N_16819,N_16874);
or U17645 (N_17645,N_16988,N_16938);
xnor U17646 (N_17646,N_16741,N_16885);
and U17647 (N_17647,N_16481,N_16718);
nand U17648 (N_17648,N_16666,N_16681);
or U17649 (N_17649,N_16843,N_16409);
and U17650 (N_17650,N_16683,N_16685);
nand U17651 (N_17651,N_16428,N_16113);
nor U17652 (N_17652,N_16140,N_16067);
nor U17653 (N_17653,N_16371,N_16755);
nand U17654 (N_17654,N_16430,N_16036);
or U17655 (N_17655,N_16056,N_16685);
nor U17656 (N_17656,N_16541,N_16668);
and U17657 (N_17657,N_16456,N_16194);
nand U17658 (N_17658,N_16028,N_16577);
xor U17659 (N_17659,N_16573,N_16900);
nor U17660 (N_17660,N_16449,N_16734);
or U17661 (N_17661,N_16677,N_16384);
or U17662 (N_17662,N_16547,N_16745);
and U17663 (N_17663,N_16878,N_16720);
or U17664 (N_17664,N_16998,N_16052);
nor U17665 (N_17665,N_16468,N_16449);
or U17666 (N_17666,N_16250,N_16113);
nand U17667 (N_17667,N_16729,N_16463);
and U17668 (N_17668,N_16323,N_16059);
nor U17669 (N_17669,N_16477,N_16914);
or U17670 (N_17670,N_16724,N_16231);
xor U17671 (N_17671,N_16045,N_16185);
and U17672 (N_17672,N_16459,N_16646);
nor U17673 (N_17673,N_16622,N_16539);
and U17674 (N_17674,N_16416,N_16580);
nor U17675 (N_17675,N_16886,N_16887);
nand U17676 (N_17676,N_16436,N_16853);
and U17677 (N_17677,N_16704,N_16585);
xnor U17678 (N_17678,N_16184,N_16322);
or U17679 (N_17679,N_16931,N_16014);
xor U17680 (N_17680,N_16524,N_16092);
nand U17681 (N_17681,N_16422,N_16808);
and U17682 (N_17682,N_16674,N_16436);
xor U17683 (N_17683,N_16956,N_16183);
or U17684 (N_17684,N_16741,N_16323);
nor U17685 (N_17685,N_16047,N_16808);
or U17686 (N_17686,N_16995,N_16326);
nand U17687 (N_17687,N_16881,N_16577);
or U17688 (N_17688,N_16473,N_16677);
nand U17689 (N_17689,N_16479,N_16383);
xnor U17690 (N_17690,N_16664,N_16883);
xor U17691 (N_17691,N_16776,N_16455);
xor U17692 (N_17692,N_16392,N_16108);
nor U17693 (N_17693,N_16788,N_16174);
nand U17694 (N_17694,N_16450,N_16083);
and U17695 (N_17695,N_16601,N_16250);
xnor U17696 (N_17696,N_16474,N_16470);
xor U17697 (N_17697,N_16843,N_16694);
xnor U17698 (N_17698,N_16098,N_16604);
or U17699 (N_17699,N_16676,N_16570);
nand U17700 (N_17700,N_16439,N_16284);
xor U17701 (N_17701,N_16172,N_16453);
or U17702 (N_17702,N_16260,N_16060);
nor U17703 (N_17703,N_16056,N_16191);
nor U17704 (N_17704,N_16810,N_16983);
nand U17705 (N_17705,N_16908,N_16548);
nand U17706 (N_17706,N_16311,N_16919);
nor U17707 (N_17707,N_16236,N_16802);
nor U17708 (N_17708,N_16371,N_16082);
nor U17709 (N_17709,N_16514,N_16709);
nand U17710 (N_17710,N_16917,N_16732);
nor U17711 (N_17711,N_16467,N_16061);
nand U17712 (N_17712,N_16232,N_16654);
nor U17713 (N_17713,N_16059,N_16614);
xor U17714 (N_17714,N_16010,N_16128);
or U17715 (N_17715,N_16171,N_16652);
and U17716 (N_17716,N_16377,N_16087);
or U17717 (N_17717,N_16095,N_16618);
nor U17718 (N_17718,N_16334,N_16426);
nand U17719 (N_17719,N_16775,N_16079);
nor U17720 (N_17720,N_16980,N_16218);
nand U17721 (N_17721,N_16045,N_16449);
and U17722 (N_17722,N_16315,N_16796);
nand U17723 (N_17723,N_16105,N_16652);
or U17724 (N_17724,N_16158,N_16524);
nand U17725 (N_17725,N_16873,N_16244);
or U17726 (N_17726,N_16259,N_16938);
xnor U17727 (N_17727,N_16031,N_16460);
nand U17728 (N_17728,N_16397,N_16854);
nor U17729 (N_17729,N_16653,N_16172);
nand U17730 (N_17730,N_16790,N_16584);
or U17731 (N_17731,N_16854,N_16121);
and U17732 (N_17732,N_16887,N_16161);
or U17733 (N_17733,N_16337,N_16673);
nor U17734 (N_17734,N_16062,N_16101);
or U17735 (N_17735,N_16007,N_16553);
nand U17736 (N_17736,N_16226,N_16049);
and U17737 (N_17737,N_16736,N_16517);
xnor U17738 (N_17738,N_16454,N_16341);
nand U17739 (N_17739,N_16480,N_16577);
or U17740 (N_17740,N_16136,N_16166);
nand U17741 (N_17741,N_16140,N_16073);
or U17742 (N_17742,N_16108,N_16123);
or U17743 (N_17743,N_16939,N_16493);
nor U17744 (N_17744,N_16093,N_16822);
xor U17745 (N_17745,N_16098,N_16216);
or U17746 (N_17746,N_16885,N_16850);
xor U17747 (N_17747,N_16287,N_16526);
nor U17748 (N_17748,N_16542,N_16455);
or U17749 (N_17749,N_16935,N_16211);
or U17750 (N_17750,N_16845,N_16102);
xnor U17751 (N_17751,N_16389,N_16011);
or U17752 (N_17752,N_16372,N_16334);
nor U17753 (N_17753,N_16173,N_16947);
nand U17754 (N_17754,N_16366,N_16281);
nor U17755 (N_17755,N_16055,N_16526);
nor U17756 (N_17756,N_16737,N_16821);
xnor U17757 (N_17757,N_16339,N_16585);
or U17758 (N_17758,N_16466,N_16129);
or U17759 (N_17759,N_16410,N_16303);
xnor U17760 (N_17760,N_16374,N_16583);
xnor U17761 (N_17761,N_16998,N_16242);
nor U17762 (N_17762,N_16205,N_16774);
xor U17763 (N_17763,N_16664,N_16089);
nor U17764 (N_17764,N_16310,N_16131);
xnor U17765 (N_17765,N_16605,N_16870);
and U17766 (N_17766,N_16289,N_16147);
or U17767 (N_17767,N_16389,N_16400);
xnor U17768 (N_17768,N_16122,N_16121);
xor U17769 (N_17769,N_16423,N_16854);
nand U17770 (N_17770,N_16890,N_16539);
and U17771 (N_17771,N_16951,N_16196);
nand U17772 (N_17772,N_16517,N_16477);
nor U17773 (N_17773,N_16247,N_16244);
xnor U17774 (N_17774,N_16674,N_16152);
and U17775 (N_17775,N_16306,N_16056);
or U17776 (N_17776,N_16057,N_16618);
xor U17777 (N_17777,N_16076,N_16840);
nor U17778 (N_17778,N_16779,N_16992);
nor U17779 (N_17779,N_16728,N_16577);
nor U17780 (N_17780,N_16731,N_16539);
xor U17781 (N_17781,N_16112,N_16144);
nand U17782 (N_17782,N_16770,N_16492);
nor U17783 (N_17783,N_16452,N_16530);
nor U17784 (N_17784,N_16664,N_16003);
or U17785 (N_17785,N_16836,N_16733);
nand U17786 (N_17786,N_16709,N_16006);
nand U17787 (N_17787,N_16860,N_16578);
or U17788 (N_17788,N_16070,N_16265);
and U17789 (N_17789,N_16339,N_16537);
nor U17790 (N_17790,N_16853,N_16830);
xnor U17791 (N_17791,N_16054,N_16222);
and U17792 (N_17792,N_16132,N_16156);
xnor U17793 (N_17793,N_16338,N_16193);
xnor U17794 (N_17794,N_16959,N_16644);
and U17795 (N_17795,N_16390,N_16104);
xor U17796 (N_17796,N_16245,N_16420);
nor U17797 (N_17797,N_16741,N_16921);
or U17798 (N_17798,N_16339,N_16482);
nor U17799 (N_17799,N_16367,N_16544);
and U17800 (N_17800,N_16794,N_16785);
xnor U17801 (N_17801,N_16012,N_16360);
nor U17802 (N_17802,N_16392,N_16347);
or U17803 (N_17803,N_16751,N_16898);
nor U17804 (N_17804,N_16345,N_16587);
and U17805 (N_17805,N_16982,N_16526);
or U17806 (N_17806,N_16828,N_16760);
xor U17807 (N_17807,N_16095,N_16123);
xor U17808 (N_17808,N_16050,N_16041);
xnor U17809 (N_17809,N_16062,N_16087);
xnor U17810 (N_17810,N_16045,N_16377);
and U17811 (N_17811,N_16761,N_16515);
or U17812 (N_17812,N_16145,N_16801);
and U17813 (N_17813,N_16847,N_16744);
nor U17814 (N_17814,N_16717,N_16871);
nor U17815 (N_17815,N_16492,N_16478);
or U17816 (N_17816,N_16760,N_16867);
and U17817 (N_17817,N_16283,N_16672);
or U17818 (N_17818,N_16795,N_16881);
nor U17819 (N_17819,N_16076,N_16035);
xor U17820 (N_17820,N_16722,N_16418);
nand U17821 (N_17821,N_16527,N_16954);
nand U17822 (N_17822,N_16991,N_16611);
nand U17823 (N_17823,N_16293,N_16653);
and U17824 (N_17824,N_16732,N_16308);
xor U17825 (N_17825,N_16803,N_16079);
xor U17826 (N_17826,N_16795,N_16056);
nor U17827 (N_17827,N_16703,N_16747);
and U17828 (N_17828,N_16171,N_16426);
nor U17829 (N_17829,N_16731,N_16793);
nor U17830 (N_17830,N_16584,N_16883);
nor U17831 (N_17831,N_16862,N_16704);
xnor U17832 (N_17832,N_16753,N_16141);
nor U17833 (N_17833,N_16074,N_16320);
nor U17834 (N_17834,N_16346,N_16495);
and U17835 (N_17835,N_16210,N_16767);
and U17836 (N_17836,N_16021,N_16501);
xnor U17837 (N_17837,N_16093,N_16944);
xnor U17838 (N_17838,N_16054,N_16665);
and U17839 (N_17839,N_16385,N_16364);
xnor U17840 (N_17840,N_16868,N_16686);
nor U17841 (N_17841,N_16769,N_16737);
and U17842 (N_17842,N_16626,N_16028);
and U17843 (N_17843,N_16446,N_16357);
xnor U17844 (N_17844,N_16302,N_16164);
nand U17845 (N_17845,N_16223,N_16172);
xor U17846 (N_17846,N_16216,N_16286);
xor U17847 (N_17847,N_16523,N_16083);
or U17848 (N_17848,N_16532,N_16771);
nand U17849 (N_17849,N_16363,N_16063);
nand U17850 (N_17850,N_16147,N_16047);
and U17851 (N_17851,N_16287,N_16256);
nor U17852 (N_17852,N_16406,N_16610);
and U17853 (N_17853,N_16186,N_16684);
nand U17854 (N_17854,N_16094,N_16574);
nor U17855 (N_17855,N_16702,N_16850);
or U17856 (N_17856,N_16765,N_16923);
or U17857 (N_17857,N_16887,N_16570);
xnor U17858 (N_17858,N_16518,N_16508);
or U17859 (N_17859,N_16629,N_16484);
nand U17860 (N_17860,N_16453,N_16966);
nor U17861 (N_17861,N_16188,N_16505);
or U17862 (N_17862,N_16450,N_16801);
and U17863 (N_17863,N_16741,N_16028);
and U17864 (N_17864,N_16508,N_16215);
or U17865 (N_17865,N_16722,N_16918);
nand U17866 (N_17866,N_16835,N_16666);
and U17867 (N_17867,N_16145,N_16074);
and U17868 (N_17868,N_16242,N_16930);
nor U17869 (N_17869,N_16055,N_16337);
xnor U17870 (N_17870,N_16965,N_16503);
xnor U17871 (N_17871,N_16905,N_16078);
and U17872 (N_17872,N_16719,N_16857);
nand U17873 (N_17873,N_16919,N_16482);
and U17874 (N_17874,N_16725,N_16349);
xor U17875 (N_17875,N_16812,N_16349);
nor U17876 (N_17876,N_16484,N_16532);
nor U17877 (N_17877,N_16551,N_16149);
xnor U17878 (N_17878,N_16242,N_16944);
nor U17879 (N_17879,N_16784,N_16959);
xnor U17880 (N_17880,N_16801,N_16623);
nand U17881 (N_17881,N_16081,N_16114);
nand U17882 (N_17882,N_16646,N_16751);
xnor U17883 (N_17883,N_16701,N_16840);
nor U17884 (N_17884,N_16888,N_16734);
or U17885 (N_17885,N_16151,N_16122);
nand U17886 (N_17886,N_16970,N_16998);
nor U17887 (N_17887,N_16039,N_16126);
or U17888 (N_17888,N_16462,N_16261);
nand U17889 (N_17889,N_16742,N_16393);
nor U17890 (N_17890,N_16192,N_16962);
or U17891 (N_17891,N_16891,N_16489);
nand U17892 (N_17892,N_16408,N_16233);
nand U17893 (N_17893,N_16527,N_16434);
nor U17894 (N_17894,N_16477,N_16606);
nor U17895 (N_17895,N_16493,N_16397);
and U17896 (N_17896,N_16172,N_16369);
xnor U17897 (N_17897,N_16646,N_16638);
nand U17898 (N_17898,N_16932,N_16885);
and U17899 (N_17899,N_16263,N_16128);
and U17900 (N_17900,N_16696,N_16548);
and U17901 (N_17901,N_16949,N_16753);
nor U17902 (N_17902,N_16536,N_16256);
and U17903 (N_17903,N_16435,N_16597);
and U17904 (N_17904,N_16159,N_16571);
or U17905 (N_17905,N_16369,N_16002);
and U17906 (N_17906,N_16853,N_16021);
nand U17907 (N_17907,N_16153,N_16436);
nand U17908 (N_17908,N_16781,N_16150);
xor U17909 (N_17909,N_16817,N_16855);
and U17910 (N_17910,N_16719,N_16229);
or U17911 (N_17911,N_16431,N_16970);
nor U17912 (N_17912,N_16089,N_16561);
xor U17913 (N_17913,N_16041,N_16010);
and U17914 (N_17914,N_16948,N_16027);
and U17915 (N_17915,N_16291,N_16182);
nand U17916 (N_17916,N_16636,N_16643);
xor U17917 (N_17917,N_16395,N_16879);
xor U17918 (N_17918,N_16336,N_16018);
xnor U17919 (N_17919,N_16624,N_16883);
nand U17920 (N_17920,N_16481,N_16727);
xor U17921 (N_17921,N_16014,N_16475);
nand U17922 (N_17922,N_16215,N_16511);
or U17923 (N_17923,N_16202,N_16845);
nand U17924 (N_17924,N_16073,N_16158);
nand U17925 (N_17925,N_16956,N_16192);
or U17926 (N_17926,N_16423,N_16467);
or U17927 (N_17927,N_16852,N_16091);
or U17928 (N_17928,N_16849,N_16852);
nand U17929 (N_17929,N_16819,N_16688);
nor U17930 (N_17930,N_16133,N_16889);
nand U17931 (N_17931,N_16281,N_16668);
nand U17932 (N_17932,N_16385,N_16129);
nor U17933 (N_17933,N_16722,N_16768);
nand U17934 (N_17934,N_16197,N_16232);
nor U17935 (N_17935,N_16259,N_16693);
and U17936 (N_17936,N_16167,N_16992);
nand U17937 (N_17937,N_16489,N_16613);
and U17938 (N_17938,N_16529,N_16626);
or U17939 (N_17939,N_16312,N_16505);
and U17940 (N_17940,N_16256,N_16358);
and U17941 (N_17941,N_16895,N_16647);
nand U17942 (N_17942,N_16087,N_16343);
nand U17943 (N_17943,N_16225,N_16785);
xor U17944 (N_17944,N_16270,N_16463);
xnor U17945 (N_17945,N_16796,N_16961);
and U17946 (N_17946,N_16465,N_16463);
nor U17947 (N_17947,N_16565,N_16561);
nand U17948 (N_17948,N_16067,N_16473);
nand U17949 (N_17949,N_16058,N_16112);
nor U17950 (N_17950,N_16652,N_16476);
xor U17951 (N_17951,N_16200,N_16141);
nor U17952 (N_17952,N_16606,N_16586);
nand U17953 (N_17953,N_16406,N_16460);
nand U17954 (N_17954,N_16890,N_16700);
and U17955 (N_17955,N_16926,N_16270);
nor U17956 (N_17956,N_16613,N_16904);
nor U17957 (N_17957,N_16211,N_16561);
xor U17958 (N_17958,N_16938,N_16142);
and U17959 (N_17959,N_16353,N_16605);
xnor U17960 (N_17960,N_16026,N_16554);
and U17961 (N_17961,N_16454,N_16771);
xor U17962 (N_17962,N_16090,N_16231);
nand U17963 (N_17963,N_16359,N_16642);
or U17964 (N_17964,N_16136,N_16467);
nand U17965 (N_17965,N_16833,N_16146);
and U17966 (N_17966,N_16009,N_16664);
nor U17967 (N_17967,N_16550,N_16539);
nand U17968 (N_17968,N_16613,N_16247);
and U17969 (N_17969,N_16499,N_16264);
nand U17970 (N_17970,N_16485,N_16773);
xnor U17971 (N_17971,N_16507,N_16293);
xnor U17972 (N_17972,N_16735,N_16507);
nor U17973 (N_17973,N_16328,N_16347);
xnor U17974 (N_17974,N_16826,N_16505);
and U17975 (N_17975,N_16941,N_16505);
or U17976 (N_17976,N_16225,N_16128);
and U17977 (N_17977,N_16870,N_16391);
or U17978 (N_17978,N_16841,N_16476);
nand U17979 (N_17979,N_16270,N_16302);
nor U17980 (N_17980,N_16475,N_16169);
and U17981 (N_17981,N_16741,N_16183);
xor U17982 (N_17982,N_16723,N_16817);
and U17983 (N_17983,N_16549,N_16974);
or U17984 (N_17984,N_16642,N_16134);
xor U17985 (N_17985,N_16843,N_16788);
xnor U17986 (N_17986,N_16033,N_16667);
xor U17987 (N_17987,N_16632,N_16137);
or U17988 (N_17988,N_16527,N_16548);
nor U17989 (N_17989,N_16315,N_16871);
nand U17990 (N_17990,N_16574,N_16779);
or U17991 (N_17991,N_16312,N_16752);
or U17992 (N_17992,N_16821,N_16921);
or U17993 (N_17993,N_16818,N_16910);
nand U17994 (N_17994,N_16255,N_16054);
nand U17995 (N_17995,N_16988,N_16005);
nand U17996 (N_17996,N_16223,N_16059);
and U17997 (N_17997,N_16226,N_16785);
nor U17998 (N_17998,N_16984,N_16866);
nor U17999 (N_17999,N_16529,N_16480);
and U18000 (N_18000,N_17164,N_17882);
xnor U18001 (N_18001,N_17498,N_17246);
nor U18002 (N_18002,N_17703,N_17033);
nand U18003 (N_18003,N_17960,N_17530);
xnor U18004 (N_18004,N_17435,N_17817);
nor U18005 (N_18005,N_17282,N_17311);
and U18006 (N_18006,N_17627,N_17385);
xor U18007 (N_18007,N_17630,N_17854);
and U18008 (N_18008,N_17716,N_17302);
xnor U18009 (N_18009,N_17834,N_17429);
nor U18010 (N_18010,N_17256,N_17196);
and U18011 (N_18011,N_17513,N_17649);
and U18012 (N_18012,N_17329,N_17014);
xor U18013 (N_18013,N_17933,N_17170);
and U18014 (N_18014,N_17792,N_17327);
nor U18015 (N_18015,N_17326,N_17022);
or U18016 (N_18016,N_17724,N_17713);
or U18017 (N_18017,N_17147,N_17367);
nand U18018 (N_18018,N_17184,N_17454);
nand U18019 (N_18019,N_17228,N_17337);
xnor U18020 (N_18020,N_17797,N_17643);
xor U18021 (N_18021,N_17511,N_17440);
nor U18022 (N_18022,N_17269,N_17897);
or U18023 (N_18023,N_17614,N_17119);
nand U18024 (N_18024,N_17777,N_17274);
or U18025 (N_18025,N_17330,N_17050);
nor U18026 (N_18026,N_17814,N_17027);
xnor U18027 (N_18027,N_17870,N_17958);
nor U18028 (N_18028,N_17839,N_17827);
nand U18029 (N_18029,N_17430,N_17217);
nor U18030 (N_18030,N_17881,N_17035);
or U18031 (N_18031,N_17542,N_17500);
and U18032 (N_18032,N_17657,N_17725);
nor U18033 (N_18033,N_17205,N_17998);
nor U18034 (N_18034,N_17158,N_17846);
nor U18035 (N_18035,N_17481,N_17504);
and U18036 (N_18036,N_17991,N_17512);
xnor U18037 (N_18037,N_17115,N_17539);
nor U18038 (N_18038,N_17732,N_17128);
and U18039 (N_18039,N_17038,N_17366);
xor U18040 (N_18040,N_17772,N_17324);
xor U18041 (N_18041,N_17284,N_17123);
xnor U18042 (N_18042,N_17719,N_17080);
nand U18043 (N_18043,N_17737,N_17702);
xor U18044 (N_18044,N_17253,N_17532);
nor U18045 (N_18045,N_17825,N_17893);
nand U18046 (N_18046,N_17585,N_17801);
or U18047 (N_18047,N_17616,N_17306);
or U18048 (N_18048,N_17784,N_17473);
and U18049 (N_18049,N_17736,N_17851);
xnor U18050 (N_18050,N_17235,N_17578);
and U18051 (N_18051,N_17470,N_17364);
and U18052 (N_18052,N_17178,N_17304);
nand U18053 (N_18053,N_17360,N_17187);
nand U18054 (N_18054,N_17541,N_17706);
nor U18055 (N_18055,N_17670,N_17740);
or U18056 (N_18056,N_17632,N_17489);
or U18057 (N_18057,N_17661,N_17995);
nand U18058 (N_18058,N_17894,N_17179);
nand U18059 (N_18059,N_17445,N_17727);
xor U18060 (N_18060,N_17949,N_17798);
and U18061 (N_18061,N_17533,N_17638);
or U18062 (N_18062,N_17457,N_17303);
or U18063 (N_18063,N_17656,N_17193);
nand U18064 (N_18064,N_17767,N_17804);
and U18065 (N_18065,N_17689,N_17260);
nand U18066 (N_18066,N_17186,N_17721);
nor U18067 (N_18067,N_17211,N_17848);
nand U18068 (N_18068,N_17712,N_17058);
xnor U18069 (N_18069,N_17754,N_17416);
and U18070 (N_18070,N_17667,N_17734);
and U18071 (N_18071,N_17644,N_17259);
or U18072 (N_18072,N_17354,N_17421);
xnor U18073 (N_18073,N_17771,N_17499);
nand U18074 (N_18074,N_17990,N_17313);
or U18075 (N_18075,N_17864,N_17983);
and U18076 (N_18076,N_17060,N_17456);
xnor U18077 (N_18077,N_17546,N_17538);
or U18078 (N_18078,N_17688,N_17907);
nand U18079 (N_18079,N_17493,N_17800);
or U18080 (N_18080,N_17595,N_17908);
xnor U18081 (N_18081,N_17185,N_17034);
nand U18082 (N_18082,N_17382,N_17258);
xor U18083 (N_18083,N_17224,N_17475);
xnor U18084 (N_18084,N_17929,N_17947);
or U18085 (N_18085,N_17890,N_17066);
nand U18086 (N_18086,N_17016,N_17073);
or U18087 (N_18087,N_17902,N_17793);
nor U18088 (N_18088,N_17357,N_17815);
and U18089 (N_18089,N_17888,N_17519);
and U18090 (N_18090,N_17979,N_17130);
nand U18091 (N_18091,N_17895,N_17932);
xor U18092 (N_18092,N_17984,N_17601);
and U18093 (N_18093,N_17915,N_17999);
nor U18094 (N_18094,N_17353,N_17321);
xnor U18095 (N_18095,N_17494,N_17889);
nand U18096 (N_18096,N_17629,N_17399);
xnor U18097 (N_18097,N_17172,N_17218);
or U18098 (N_18098,N_17446,N_17537);
nor U18099 (N_18099,N_17203,N_17666);
and U18100 (N_18100,N_17510,N_17559);
and U18101 (N_18101,N_17518,N_17459);
or U18102 (N_18102,N_17183,N_17091);
or U18103 (N_18103,N_17904,N_17124);
xnor U18104 (N_18104,N_17816,N_17396);
and U18105 (N_18105,N_17220,N_17845);
or U18106 (N_18106,N_17820,N_17344);
nand U18107 (N_18107,N_17129,N_17913);
xor U18108 (N_18108,N_17738,N_17605);
nor U18109 (N_18109,N_17450,N_17189);
nand U18110 (N_18110,N_17790,N_17230);
or U18111 (N_18111,N_17005,N_17608);
nor U18112 (N_18112,N_17660,N_17223);
xnor U18113 (N_18113,N_17868,N_17215);
or U18114 (N_18114,N_17380,N_17955);
nor U18115 (N_18115,N_17965,N_17098);
xnor U18116 (N_18116,N_17505,N_17583);
nand U18117 (N_18117,N_17783,N_17628);
nor U18118 (N_18118,N_17349,N_17507);
nor U18119 (N_18119,N_17535,N_17462);
nor U18120 (N_18120,N_17696,N_17351);
xor U18121 (N_18121,N_17658,N_17819);
and U18122 (N_18122,N_17867,N_17837);
and U18123 (N_18123,N_17049,N_17503);
and U18124 (N_18124,N_17836,N_17233);
nand U18125 (N_18125,N_17097,N_17569);
or U18126 (N_18126,N_17557,N_17144);
nand U18127 (N_18127,N_17502,N_17176);
nand U18128 (N_18128,N_17662,N_17461);
nor U18129 (N_18129,N_17191,N_17392);
nor U18130 (N_18130,N_17645,N_17150);
or U18131 (N_18131,N_17755,N_17331);
and U18132 (N_18132,N_17579,N_17883);
xor U18133 (N_18133,N_17765,N_17099);
nand U18134 (N_18134,N_17674,N_17808);
or U18135 (N_18135,N_17297,N_17722);
or U18136 (N_18136,N_17101,N_17928);
nand U18137 (N_18137,N_17015,N_17387);
or U18138 (N_18138,N_17280,N_17698);
or U18139 (N_18139,N_17003,N_17561);
and U18140 (N_18140,N_17672,N_17198);
nand U18141 (N_18141,N_17690,N_17679);
xnor U18142 (N_18142,N_17480,N_17781);
or U18143 (N_18143,N_17789,N_17972);
and U18144 (N_18144,N_17550,N_17173);
xnor U18145 (N_18145,N_17395,N_17718);
nand U18146 (N_18146,N_17753,N_17594);
nor U18147 (N_18147,N_17394,N_17611);
or U18148 (N_18148,N_17342,N_17948);
or U18149 (N_18149,N_17403,N_17156);
nor U18150 (N_18150,N_17476,N_17121);
nand U18151 (N_18151,N_17132,N_17835);
nand U18152 (N_18152,N_17365,N_17917);
xnor U18153 (N_18153,N_17285,N_17602);
xor U18154 (N_18154,N_17522,N_17149);
xor U18155 (N_18155,N_17409,N_17886);
xnor U18156 (N_18156,N_17333,N_17386);
or U18157 (N_18157,N_17523,N_17940);
xnor U18158 (N_18158,N_17756,N_17796);
and U18159 (N_18159,N_17350,N_17934);
and U18160 (N_18160,N_17226,N_17201);
nand U18161 (N_18161,N_17245,N_17930);
and U18162 (N_18162,N_17731,N_17267);
nand U18163 (N_18163,N_17566,N_17390);
or U18164 (N_18164,N_17707,N_17131);
xnor U18165 (N_18165,N_17992,N_17479);
nand U18166 (N_18166,N_17251,N_17885);
and U18167 (N_18167,N_17104,N_17053);
and U18168 (N_18168,N_17458,N_17239);
nor U18169 (N_18169,N_17813,N_17216);
or U18170 (N_18170,N_17401,N_17869);
nor U18171 (N_18171,N_17584,N_17163);
or U18172 (N_18172,N_17126,N_17412);
and U18173 (N_18173,N_17199,N_17597);
nor U18174 (N_18174,N_17708,N_17574);
nand U18175 (N_18175,N_17957,N_17914);
nand U18176 (N_18176,N_17213,N_17593);
xnor U18177 (N_18177,N_17142,N_17775);
xnor U18178 (N_18178,N_17424,N_17271);
and U18179 (N_18179,N_17279,N_17116);
nor U18180 (N_18180,N_17317,N_17202);
nor U18181 (N_18181,N_17155,N_17439);
xnor U18182 (N_18182,N_17204,N_17410);
xnor U18183 (N_18183,N_17174,N_17840);
xnor U18184 (N_18184,N_17105,N_17041);
xnor U18185 (N_18185,N_17741,N_17653);
nand U18186 (N_18186,N_17175,N_17810);
or U18187 (N_18187,N_17023,N_17582);
nor U18188 (N_18188,N_17953,N_17857);
nor U18189 (N_18189,N_17094,N_17369);
xnor U18190 (N_18190,N_17111,N_17451);
nand U18191 (N_18191,N_17229,N_17418);
nor U18192 (N_18192,N_17361,N_17540);
nor U18193 (N_18193,N_17009,N_17381);
xor U18194 (N_18194,N_17844,N_17137);
nor U18195 (N_18195,N_17562,N_17341);
xnor U18196 (N_18196,N_17340,N_17580);
nand U18197 (N_18197,N_17257,N_17545);
xor U18198 (N_18198,N_17905,N_17596);
or U18199 (N_18199,N_17044,N_17560);
nor U18200 (N_18200,N_17521,N_17927);
xnor U18201 (N_18201,N_17607,N_17310);
nand U18202 (N_18202,N_17296,N_17809);
nor U18203 (N_18203,N_17109,N_17946);
and U18204 (N_18204,N_17609,N_17770);
or U18205 (N_18205,N_17008,N_17799);
or U18206 (N_18206,N_17743,N_17400);
nand U18207 (N_18207,N_17024,N_17414);
xor U18208 (N_18208,N_17241,N_17676);
and U18209 (N_18209,N_17705,N_17923);
and U18210 (N_18210,N_17768,N_17633);
xor U18211 (N_18211,N_17752,N_17135);
or U18212 (N_18212,N_17020,N_17025);
nor U18213 (N_18213,N_17478,N_17264);
or U18214 (N_18214,N_17046,N_17549);
xnor U18215 (N_18215,N_17081,N_17273);
nor U18216 (N_18216,N_17452,N_17134);
nor U18217 (N_18217,N_17878,N_17455);
xor U18218 (N_18218,N_17085,N_17962);
nor U18219 (N_18219,N_17648,N_17346);
nand U18220 (N_18220,N_17860,N_17862);
and U18221 (N_18221,N_17056,N_17637);
nand U18222 (N_18222,N_17944,N_17336);
or U18223 (N_18223,N_17778,N_17898);
or U18224 (N_18224,N_17723,N_17673);
or U18225 (N_18225,N_17055,N_17288);
xor U18226 (N_18226,N_17751,N_17477);
or U18227 (N_18227,N_17420,N_17573);
nand U18228 (N_18228,N_17240,N_17106);
nor U18229 (N_18229,N_17717,N_17000);
nor U18230 (N_18230,N_17236,N_17291);
xor U18231 (N_18231,N_17833,N_17818);
or U18232 (N_18232,N_17286,N_17266);
nor U18233 (N_18233,N_17745,N_17697);
xnor U18234 (N_18234,N_17831,N_17695);
and U18235 (N_18235,N_17626,N_17048);
nand U18236 (N_18236,N_17334,N_17262);
and U18237 (N_18237,N_17806,N_17681);
and U18238 (N_18238,N_17275,N_17467);
nand U18239 (N_18239,N_17181,N_17423);
nand U18240 (N_18240,N_17875,N_17576);
nand U18241 (N_18241,N_17987,N_17985);
and U18242 (N_18242,N_17971,N_17376);
and U18243 (N_18243,N_17293,N_17428);
xnor U18244 (N_18244,N_17515,N_17243);
nor U18245 (N_18245,N_17136,N_17460);
nor U18246 (N_18246,N_17847,N_17036);
or U18247 (N_18247,N_17299,N_17685);
nand U18248 (N_18248,N_17071,N_17100);
and U18249 (N_18249,N_17952,N_17794);
or U18250 (N_18250,N_17988,N_17853);
and U18251 (N_18251,N_17887,N_17042);
nand U18252 (N_18252,N_17120,N_17018);
or U18253 (N_18253,N_17852,N_17391);
xnor U18254 (N_18254,N_17077,N_17617);
xor U18255 (N_18255,N_17884,N_17069);
xor U18256 (N_18256,N_17182,N_17320);
nor U18257 (N_18257,N_17981,N_17973);
xor U18258 (N_18258,N_17664,N_17552);
xor U18259 (N_18259,N_17338,N_17675);
nor U18260 (N_18260,N_17861,N_17671);
and U18261 (N_18261,N_17209,N_17486);
nor U18262 (N_18262,N_17082,N_17701);
or U18263 (N_18263,N_17567,N_17910);
xnor U18264 (N_18264,N_17490,N_17222);
nor U18265 (N_18265,N_17974,N_17919);
xor U18266 (N_18266,N_17002,N_17612);
or U18267 (N_18267,N_17787,N_17484);
or U18268 (N_18268,N_17619,N_17556);
nor U18269 (N_18269,N_17406,N_17072);
and U18270 (N_18270,N_17849,N_17733);
nor U18271 (N_18271,N_17047,N_17766);
or U18272 (N_18272,N_17352,N_17654);
and U18273 (N_18273,N_17729,N_17699);
and U18274 (N_18274,N_17856,N_17146);
nand U18275 (N_18275,N_17465,N_17600);
nor U18276 (N_18276,N_17052,N_17501);
nor U18277 (N_18277,N_17265,N_17975);
nand U18278 (N_18278,N_17232,N_17323);
and U18279 (N_18279,N_17903,N_17029);
xnor U18280 (N_18280,N_17281,N_17892);
or U18281 (N_18281,N_17314,N_17832);
or U18282 (N_18282,N_17826,N_17374);
xor U18283 (N_18283,N_17355,N_17590);
nor U18284 (N_18284,N_17531,N_17305);
nand U18285 (N_18285,N_17263,N_17372);
and U18286 (N_18286,N_17599,N_17488);
nor U18287 (N_18287,N_17298,N_17307);
and U18288 (N_18288,N_17828,N_17166);
nand U18289 (N_18289,N_17431,N_17936);
and U18290 (N_18290,N_17037,N_17659);
and U18291 (N_18291,N_17709,N_17339);
and U18292 (N_18292,N_17970,N_17565);
nor U18293 (N_18293,N_17634,N_17362);
and U18294 (N_18294,N_17370,N_17017);
xor U18295 (N_18295,N_17436,N_17117);
and U18296 (N_18296,N_17212,N_17348);
nand U18297 (N_18297,N_17425,N_17891);
nand U18298 (N_18298,N_17192,N_17610);
and U18299 (N_18299,N_17980,N_17624);
and U18300 (N_18300,N_17102,N_17151);
nor U18301 (N_18301,N_17730,N_17141);
nand U18302 (N_18302,N_17750,N_17976);
xor U18303 (N_18303,N_17295,N_17270);
xnor U18304 (N_18304,N_17997,N_17841);
and U18305 (N_18305,N_17802,N_17742);
and U18306 (N_18306,N_17994,N_17700);
xor U18307 (N_18307,N_17227,N_17843);
and U18308 (N_18308,N_17921,N_17277);
nor U18309 (N_18309,N_17786,N_17631);
nand U18310 (N_18310,N_17438,N_17554);
nand U18311 (N_18311,N_17829,N_17208);
nor U18312 (N_18312,N_17922,N_17443);
xor U18313 (N_18313,N_17062,N_17735);
nand U18314 (N_18314,N_17879,N_17553);
and U18315 (N_18315,N_17858,N_17650);
nor U18316 (N_18316,N_17899,N_17300);
nand U18317 (N_18317,N_17509,N_17757);
nand U18318 (N_18318,N_17032,N_17093);
nand U18319 (N_18319,N_17063,N_17520);
or U18320 (N_18320,N_17328,N_17125);
nor U18321 (N_18321,N_17383,N_17168);
xor U18322 (N_18322,N_17639,N_17606);
or U18323 (N_18323,N_17118,N_17272);
or U18324 (N_18324,N_17603,N_17950);
or U18325 (N_18325,N_17095,N_17384);
and U18326 (N_18326,N_17951,N_17564);
nor U18327 (N_18327,N_17335,N_17761);
or U18328 (N_18328,N_17855,N_17678);
or U18329 (N_18329,N_17900,N_17096);
and U18330 (N_18330,N_17345,N_17823);
nand U18331 (N_18331,N_17647,N_17591);
xnor U18332 (N_18332,N_17363,N_17563);
nand U18333 (N_18333,N_17776,N_17551);
xor U18334 (N_18334,N_17524,N_17555);
or U18335 (N_18335,N_17916,N_17964);
nand U18336 (N_18336,N_17325,N_17165);
nor U18337 (N_18337,N_17043,N_17686);
nand U18338 (N_18338,N_17318,N_17728);
nor U18339 (N_18339,N_17061,N_17087);
nor U18340 (N_18340,N_17982,N_17157);
xnor U18341 (N_18341,N_17939,N_17108);
or U18342 (N_18342,N_17103,N_17693);
and U18343 (N_18343,N_17031,N_17759);
or U18344 (N_18344,N_17859,N_17373);
xor U18345 (N_18345,N_17824,N_17358);
xnor U18346 (N_18346,N_17961,N_17514);
or U18347 (N_18347,N_17219,N_17011);
nor U18348 (N_18348,N_17138,N_17159);
nand U18349 (N_18349,N_17937,N_17497);
or U18350 (N_18350,N_17059,N_17110);
xnor U18351 (N_18351,N_17194,N_17668);
and U18352 (N_18352,N_17237,N_17057);
nor U18353 (N_18353,N_17437,N_17162);
nand U18354 (N_18354,N_17726,N_17359);
xor U18355 (N_18355,N_17078,N_17665);
nor U18356 (N_18356,N_17850,N_17877);
and U18357 (N_18357,N_17575,N_17154);
and U18358 (N_18358,N_17838,N_17866);
nand U18359 (N_18359,N_17398,N_17986);
and U18360 (N_18360,N_17687,N_17788);
and U18361 (N_18361,N_17873,N_17920);
xor U18362 (N_18362,N_17356,N_17250);
nor U18363 (N_18363,N_17112,N_17803);
and U18364 (N_18364,N_17422,N_17758);
and U18365 (N_18365,N_17210,N_17943);
or U18366 (N_18366,N_17704,N_17516);
nand U18367 (N_18367,N_17415,N_17030);
and U18368 (N_18368,N_17487,N_17148);
and U18369 (N_18369,N_17180,N_17413);
nand U18370 (N_18370,N_17083,N_17558);
nor U18371 (N_18371,N_17064,N_17571);
xor U18372 (N_18372,N_17680,N_17931);
or U18373 (N_18373,N_17433,N_17397);
or U18374 (N_18374,N_17464,N_17427);
nor U18375 (N_18375,N_17089,N_17959);
or U18376 (N_18376,N_17065,N_17876);
nor U18377 (N_18377,N_17388,N_17641);
nor U18378 (N_18378,N_17577,N_17492);
nor U18379 (N_18379,N_17076,N_17684);
or U18380 (N_18380,N_17402,N_17769);
or U18381 (N_18381,N_17589,N_17942);
nand U18382 (N_18382,N_17710,N_17068);
or U18383 (N_18383,N_17744,N_17739);
nand U18384 (N_18384,N_17244,N_17993);
and U18385 (N_18385,N_17655,N_17663);
or U18386 (N_18386,N_17434,N_17874);
xnor U18387 (N_18387,N_17525,N_17248);
or U18388 (N_18388,N_17469,N_17088);
nor U18389 (N_18389,N_17954,N_17026);
nor U18390 (N_18390,N_17528,N_17622);
or U18391 (N_18391,N_17368,N_17544);
xor U18392 (N_18392,N_17587,N_17863);
nand U18393 (N_18393,N_17238,N_17911);
xor U18394 (N_18394,N_17805,N_17526);
and U18395 (N_18395,N_17004,N_17040);
and U18396 (N_18396,N_17651,N_17534);
and U18397 (N_18397,N_17268,N_17517);
nand U18398 (N_18398,N_17315,N_17200);
nand U18399 (N_18399,N_17652,N_17309);
nand U18400 (N_18400,N_17746,N_17592);
xnor U18401 (N_18401,N_17242,N_17720);
or U18402 (N_18402,N_17114,N_17586);
and U18403 (N_18403,N_17234,N_17570);
nand U18404 (N_18404,N_17070,N_17683);
nand U18405 (N_18405,N_17466,N_17225);
nand U18406 (N_18406,N_17871,N_17371);
nor U18407 (N_18407,N_17393,N_17086);
xor U18408 (N_18408,N_17762,N_17276);
nor U18409 (N_18409,N_17621,N_17956);
nor U18410 (N_18410,N_17912,N_17442);
and U18411 (N_18411,N_17084,N_17278);
xnor U18412 (N_18412,N_17812,N_17906);
and U18413 (N_18413,N_17308,N_17620);
xor U18414 (N_18414,N_17941,N_17945);
xor U18415 (N_18415,N_17231,N_17635);
xor U18416 (N_18416,N_17195,N_17019);
and U18417 (N_18417,N_17640,N_17214);
and U18418 (N_18418,N_17051,N_17795);
nand U18419 (N_18419,N_17791,N_17715);
xnor U18420 (N_18420,N_17347,N_17010);
nor U18421 (N_18421,N_17548,N_17773);
nand U18422 (N_18422,N_17901,N_17880);
nor U18423 (N_18423,N_17448,N_17143);
and U18424 (N_18424,N_17977,N_17935);
and U18425 (N_18425,N_17811,N_17604);
or U18426 (N_18426,N_17572,N_17377);
nand U18427 (N_18427,N_17247,N_17407);
xnor U18428 (N_18428,N_17312,N_17332);
nand U18429 (N_18429,N_17909,N_17483);
or U18430 (N_18430,N_17079,N_17006);
and U18431 (N_18431,N_17289,N_17007);
and U18432 (N_18432,N_17254,N_17821);
and U18433 (N_18433,N_17529,N_17188);
or U18434 (N_18434,N_17013,N_17714);
xnor U18435 (N_18435,N_17918,N_17426);
and U18436 (N_18436,N_17691,N_17054);
or U18437 (N_18437,N_17496,N_17568);
nor U18438 (N_18438,N_17598,N_17419);
xnor U18439 (N_18439,N_17379,N_17343);
nor U18440 (N_18440,N_17039,N_17692);
nand U18441 (N_18441,N_17764,N_17169);
nor U18442 (N_18442,N_17842,N_17167);
xnor U18443 (N_18443,N_17780,N_17506);
and U18444 (N_18444,N_17177,N_17012);
nor U18445 (N_18445,N_17581,N_17160);
or U18446 (N_18446,N_17292,N_17417);
and U18447 (N_18447,N_17411,N_17107);
xor U18448 (N_18448,N_17441,N_17319);
nand U18449 (N_18449,N_17969,N_17472);
nand U18450 (N_18450,N_17543,N_17028);
and U18451 (N_18451,N_17963,N_17140);
and U18452 (N_18452,N_17547,N_17067);
nor U18453 (N_18453,N_17133,N_17536);
and U18454 (N_18454,N_17779,N_17807);
nand U18455 (N_18455,N_17322,N_17782);
nor U18456 (N_18456,N_17045,N_17996);
nand U18457 (N_18457,N_17207,N_17113);
or U18458 (N_18458,N_17978,N_17968);
and U18459 (N_18459,N_17139,N_17763);
and U18460 (N_18460,N_17749,N_17527);
nand U18461 (N_18461,N_17444,N_17127);
xnor U18462 (N_18462,N_17316,N_17197);
xnor U18463 (N_18463,N_17774,N_17938);
xor U18464 (N_18464,N_17152,N_17485);
nand U18465 (N_18465,N_17283,N_17449);
or U18466 (N_18466,N_17508,N_17453);
xor U18467 (N_18467,N_17748,N_17122);
nor U18468 (N_18468,N_17001,N_17287);
and U18469 (N_18469,N_17491,N_17872);
and U18470 (N_18470,N_17588,N_17145);
xnor U18471 (N_18471,N_17636,N_17290);
nor U18472 (N_18472,N_17171,N_17694);
nor U18473 (N_18473,N_17405,N_17896);
nor U18474 (N_18474,N_17618,N_17925);
xor U18475 (N_18475,N_17711,N_17090);
nor U18476 (N_18476,N_17206,N_17967);
and U18477 (N_18477,N_17249,N_17646);
or U18478 (N_18478,N_17389,N_17074);
nand U18479 (N_18479,N_17625,N_17471);
xnor U18480 (N_18480,N_17682,N_17153);
nor U18481 (N_18481,N_17301,N_17482);
and U18482 (N_18482,N_17830,N_17408);
nor U18483 (N_18483,N_17785,N_17615);
xnor U18484 (N_18484,N_17190,N_17822);
and U18485 (N_18485,N_17432,N_17669);
and U18486 (N_18486,N_17642,N_17474);
nand U18487 (N_18487,N_17989,N_17252);
or U18488 (N_18488,N_17613,N_17294);
nand U18489 (N_18489,N_17092,N_17463);
nand U18490 (N_18490,N_17404,N_17378);
nand U18491 (N_18491,N_17747,N_17075);
and U18492 (N_18492,N_17447,N_17021);
nor U18493 (N_18493,N_17623,N_17926);
xnor U18494 (N_18494,N_17261,N_17865);
xnor U18495 (N_18495,N_17495,N_17255);
or U18496 (N_18496,N_17375,N_17966);
xor U18497 (N_18497,N_17468,N_17924);
or U18498 (N_18498,N_17161,N_17677);
nor U18499 (N_18499,N_17221,N_17760);
and U18500 (N_18500,N_17765,N_17885);
xor U18501 (N_18501,N_17565,N_17417);
nand U18502 (N_18502,N_17989,N_17728);
and U18503 (N_18503,N_17395,N_17010);
xor U18504 (N_18504,N_17528,N_17815);
or U18505 (N_18505,N_17132,N_17184);
nor U18506 (N_18506,N_17949,N_17269);
and U18507 (N_18507,N_17725,N_17860);
nor U18508 (N_18508,N_17135,N_17820);
and U18509 (N_18509,N_17647,N_17439);
and U18510 (N_18510,N_17815,N_17201);
and U18511 (N_18511,N_17456,N_17193);
nand U18512 (N_18512,N_17425,N_17607);
nor U18513 (N_18513,N_17963,N_17579);
and U18514 (N_18514,N_17355,N_17568);
or U18515 (N_18515,N_17731,N_17570);
xnor U18516 (N_18516,N_17584,N_17783);
nor U18517 (N_18517,N_17685,N_17067);
nand U18518 (N_18518,N_17962,N_17155);
nand U18519 (N_18519,N_17275,N_17089);
xnor U18520 (N_18520,N_17590,N_17252);
and U18521 (N_18521,N_17293,N_17477);
xor U18522 (N_18522,N_17230,N_17278);
xnor U18523 (N_18523,N_17724,N_17292);
and U18524 (N_18524,N_17241,N_17720);
nand U18525 (N_18525,N_17539,N_17850);
nor U18526 (N_18526,N_17249,N_17200);
nand U18527 (N_18527,N_17809,N_17796);
and U18528 (N_18528,N_17372,N_17721);
nand U18529 (N_18529,N_17346,N_17547);
nand U18530 (N_18530,N_17266,N_17260);
xor U18531 (N_18531,N_17992,N_17977);
or U18532 (N_18532,N_17550,N_17782);
and U18533 (N_18533,N_17261,N_17997);
and U18534 (N_18534,N_17619,N_17962);
xnor U18535 (N_18535,N_17730,N_17870);
or U18536 (N_18536,N_17259,N_17898);
xnor U18537 (N_18537,N_17373,N_17140);
or U18538 (N_18538,N_17590,N_17603);
nand U18539 (N_18539,N_17659,N_17579);
xnor U18540 (N_18540,N_17634,N_17701);
nand U18541 (N_18541,N_17194,N_17230);
xnor U18542 (N_18542,N_17155,N_17150);
nand U18543 (N_18543,N_17916,N_17097);
or U18544 (N_18544,N_17962,N_17575);
and U18545 (N_18545,N_17533,N_17632);
nor U18546 (N_18546,N_17789,N_17287);
xor U18547 (N_18547,N_17967,N_17467);
nor U18548 (N_18548,N_17619,N_17204);
nor U18549 (N_18549,N_17184,N_17482);
xnor U18550 (N_18550,N_17029,N_17947);
xor U18551 (N_18551,N_17880,N_17823);
nand U18552 (N_18552,N_17414,N_17023);
nand U18553 (N_18553,N_17998,N_17208);
nor U18554 (N_18554,N_17303,N_17993);
nand U18555 (N_18555,N_17381,N_17894);
or U18556 (N_18556,N_17535,N_17862);
nor U18557 (N_18557,N_17093,N_17703);
xor U18558 (N_18558,N_17059,N_17615);
or U18559 (N_18559,N_17756,N_17041);
nor U18560 (N_18560,N_17156,N_17172);
or U18561 (N_18561,N_17450,N_17166);
or U18562 (N_18562,N_17835,N_17725);
nand U18563 (N_18563,N_17055,N_17166);
and U18564 (N_18564,N_17756,N_17659);
nand U18565 (N_18565,N_17540,N_17800);
nor U18566 (N_18566,N_17315,N_17226);
and U18567 (N_18567,N_17179,N_17612);
or U18568 (N_18568,N_17898,N_17691);
nor U18569 (N_18569,N_17972,N_17403);
nor U18570 (N_18570,N_17030,N_17935);
and U18571 (N_18571,N_17357,N_17422);
or U18572 (N_18572,N_17878,N_17888);
and U18573 (N_18573,N_17981,N_17914);
nor U18574 (N_18574,N_17660,N_17089);
nand U18575 (N_18575,N_17218,N_17314);
nand U18576 (N_18576,N_17343,N_17509);
or U18577 (N_18577,N_17819,N_17037);
nor U18578 (N_18578,N_17223,N_17084);
and U18579 (N_18579,N_17199,N_17285);
nand U18580 (N_18580,N_17118,N_17446);
xor U18581 (N_18581,N_17424,N_17531);
and U18582 (N_18582,N_17018,N_17673);
xnor U18583 (N_18583,N_17232,N_17460);
nor U18584 (N_18584,N_17665,N_17568);
or U18585 (N_18585,N_17915,N_17956);
nor U18586 (N_18586,N_17156,N_17968);
nor U18587 (N_18587,N_17561,N_17660);
xnor U18588 (N_18588,N_17912,N_17092);
xor U18589 (N_18589,N_17573,N_17582);
nand U18590 (N_18590,N_17880,N_17211);
and U18591 (N_18591,N_17291,N_17409);
or U18592 (N_18592,N_17573,N_17718);
nand U18593 (N_18593,N_17908,N_17538);
and U18594 (N_18594,N_17414,N_17326);
xor U18595 (N_18595,N_17637,N_17341);
nor U18596 (N_18596,N_17987,N_17086);
or U18597 (N_18597,N_17964,N_17235);
and U18598 (N_18598,N_17664,N_17690);
nor U18599 (N_18599,N_17605,N_17093);
xnor U18600 (N_18600,N_17198,N_17035);
nand U18601 (N_18601,N_17310,N_17544);
and U18602 (N_18602,N_17044,N_17693);
nand U18603 (N_18603,N_17263,N_17934);
nand U18604 (N_18604,N_17271,N_17556);
and U18605 (N_18605,N_17057,N_17231);
nor U18606 (N_18606,N_17746,N_17694);
or U18607 (N_18607,N_17144,N_17544);
nand U18608 (N_18608,N_17470,N_17469);
nand U18609 (N_18609,N_17622,N_17828);
xor U18610 (N_18610,N_17792,N_17947);
nand U18611 (N_18611,N_17882,N_17657);
or U18612 (N_18612,N_17819,N_17681);
xor U18613 (N_18613,N_17774,N_17882);
xor U18614 (N_18614,N_17204,N_17544);
nand U18615 (N_18615,N_17964,N_17484);
and U18616 (N_18616,N_17356,N_17337);
nor U18617 (N_18617,N_17100,N_17740);
nand U18618 (N_18618,N_17800,N_17767);
nor U18619 (N_18619,N_17404,N_17670);
nor U18620 (N_18620,N_17602,N_17380);
and U18621 (N_18621,N_17279,N_17153);
nand U18622 (N_18622,N_17969,N_17149);
and U18623 (N_18623,N_17720,N_17635);
nand U18624 (N_18624,N_17054,N_17713);
nand U18625 (N_18625,N_17620,N_17127);
xnor U18626 (N_18626,N_17371,N_17159);
nor U18627 (N_18627,N_17995,N_17684);
and U18628 (N_18628,N_17561,N_17589);
nand U18629 (N_18629,N_17082,N_17003);
nor U18630 (N_18630,N_17963,N_17479);
or U18631 (N_18631,N_17380,N_17608);
or U18632 (N_18632,N_17614,N_17835);
nand U18633 (N_18633,N_17964,N_17741);
and U18634 (N_18634,N_17964,N_17006);
nor U18635 (N_18635,N_17800,N_17059);
nor U18636 (N_18636,N_17895,N_17935);
or U18637 (N_18637,N_17353,N_17535);
xnor U18638 (N_18638,N_17821,N_17269);
xor U18639 (N_18639,N_17822,N_17227);
xnor U18640 (N_18640,N_17100,N_17173);
xnor U18641 (N_18641,N_17229,N_17161);
nand U18642 (N_18642,N_17126,N_17026);
nand U18643 (N_18643,N_17177,N_17894);
xnor U18644 (N_18644,N_17032,N_17619);
nand U18645 (N_18645,N_17959,N_17572);
nand U18646 (N_18646,N_17996,N_17426);
xor U18647 (N_18647,N_17513,N_17905);
or U18648 (N_18648,N_17182,N_17594);
nand U18649 (N_18649,N_17266,N_17778);
nor U18650 (N_18650,N_17342,N_17789);
xnor U18651 (N_18651,N_17585,N_17368);
nand U18652 (N_18652,N_17730,N_17898);
and U18653 (N_18653,N_17705,N_17116);
or U18654 (N_18654,N_17523,N_17491);
or U18655 (N_18655,N_17612,N_17244);
xor U18656 (N_18656,N_17546,N_17779);
or U18657 (N_18657,N_17615,N_17619);
and U18658 (N_18658,N_17896,N_17175);
nor U18659 (N_18659,N_17254,N_17570);
xor U18660 (N_18660,N_17351,N_17695);
and U18661 (N_18661,N_17342,N_17561);
nor U18662 (N_18662,N_17784,N_17432);
nand U18663 (N_18663,N_17748,N_17520);
and U18664 (N_18664,N_17540,N_17024);
and U18665 (N_18665,N_17015,N_17602);
xor U18666 (N_18666,N_17248,N_17116);
and U18667 (N_18667,N_17016,N_17373);
nand U18668 (N_18668,N_17643,N_17166);
xnor U18669 (N_18669,N_17170,N_17905);
nand U18670 (N_18670,N_17894,N_17661);
nor U18671 (N_18671,N_17063,N_17625);
or U18672 (N_18672,N_17615,N_17140);
and U18673 (N_18673,N_17340,N_17533);
xnor U18674 (N_18674,N_17148,N_17051);
nand U18675 (N_18675,N_17766,N_17708);
and U18676 (N_18676,N_17974,N_17726);
xnor U18677 (N_18677,N_17896,N_17987);
xnor U18678 (N_18678,N_17858,N_17188);
nand U18679 (N_18679,N_17166,N_17817);
and U18680 (N_18680,N_17475,N_17953);
nand U18681 (N_18681,N_17626,N_17151);
nand U18682 (N_18682,N_17539,N_17170);
nand U18683 (N_18683,N_17358,N_17309);
nand U18684 (N_18684,N_17643,N_17507);
xor U18685 (N_18685,N_17481,N_17558);
nor U18686 (N_18686,N_17109,N_17939);
or U18687 (N_18687,N_17853,N_17112);
or U18688 (N_18688,N_17828,N_17178);
and U18689 (N_18689,N_17970,N_17126);
or U18690 (N_18690,N_17309,N_17141);
nand U18691 (N_18691,N_17671,N_17720);
or U18692 (N_18692,N_17687,N_17419);
or U18693 (N_18693,N_17687,N_17811);
nand U18694 (N_18694,N_17380,N_17993);
nand U18695 (N_18695,N_17261,N_17953);
nor U18696 (N_18696,N_17732,N_17397);
and U18697 (N_18697,N_17901,N_17258);
or U18698 (N_18698,N_17271,N_17891);
nor U18699 (N_18699,N_17702,N_17931);
xnor U18700 (N_18700,N_17041,N_17950);
and U18701 (N_18701,N_17618,N_17047);
nand U18702 (N_18702,N_17205,N_17789);
or U18703 (N_18703,N_17690,N_17108);
nor U18704 (N_18704,N_17170,N_17267);
or U18705 (N_18705,N_17278,N_17874);
and U18706 (N_18706,N_17480,N_17929);
nor U18707 (N_18707,N_17933,N_17173);
or U18708 (N_18708,N_17847,N_17151);
nand U18709 (N_18709,N_17204,N_17433);
or U18710 (N_18710,N_17431,N_17347);
and U18711 (N_18711,N_17023,N_17540);
or U18712 (N_18712,N_17786,N_17721);
or U18713 (N_18713,N_17081,N_17029);
and U18714 (N_18714,N_17280,N_17470);
or U18715 (N_18715,N_17816,N_17244);
nor U18716 (N_18716,N_17315,N_17594);
and U18717 (N_18717,N_17865,N_17615);
and U18718 (N_18718,N_17797,N_17554);
or U18719 (N_18719,N_17282,N_17497);
nor U18720 (N_18720,N_17766,N_17532);
nor U18721 (N_18721,N_17244,N_17766);
nor U18722 (N_18722,N_17372,N_17244);
nor U18723 (N_18723,N_17571,N_17617);
and U18724 (N_18724,N_17847,N_17731);
or U18725 (N_18725,N_17784,N_17754);
or U18726 (N_18726,N_17890,N_17811);
or U18727 (N_18727,N_17942,N_17112);
nor U18728 (N_18728,N_17917,N_17378);
or U18729 (N_18729,N_17197,N_17804);
or U18730 (N_18730,N_17241,N_17789);
xor U18731 (N_18731,N_17001,N_17568);
nor U18732 (N_18732,N_17655,N_17555);
or U18733 (N_18733,N_17904,N_17954);
and U18734 (N_18734,N_17206,N_17161);
and U18735 (N_18735,N_17882,N_17649);
nand U18736 (N_18736,N_17238,N_17777);
or U18737 (N_18737,N_17236,N_17244);
nand U18738 (N_18738,N_17378,N_17984);
nor U18739 (N_18739,N_17482,N_17171);
xnor U18740 (N_18740,N_17075,N_17308);
xnor U18741 (N_18741,N_17422,N_17237);
and U18742 (N_18742,N_17219,N_17203);
nor U18743 (N_18743,N_17366,N_17381);
and U18744 (N_18744,N_17200,N_17192);
and U18745 (N_18745,N_17472,N_17354);
and U18746 (N_18746,N_17104,N_17480);
nor U18747 (N_18747,N_17376,N_17270);
xnor U18748 (N_18748,N_17422,N_17875);
xor U18749 (N_18749,N_17737,N_17693);
or U18750 (N_18750,N_17398,N_17989);
xor U18751 (N_18751,N_17205,N_17216);
and U18752 (N_18752,N_17760,N_17101);
nand U18753 (N_18753,N_17288,N_17486);
xor U18754 (N_18754,N_17368,N_17450);
or U18755 (N_18755,N_17526,N_17731);
and U18756 (N_18756,N_17930,N_17879);
nand U18757 (N_18757,N_17819,N_17742);
nor U18758 (N_18758,N_17242,N_17093);
nand U18759 (N_18759,N_17883,N_17225);
nand U18760 (N_18760,N_17532,N_17457);
and U18761 (N_18761,N_17383,N_17018);
nor U18762 (N_18762,N_17559,N_17700);
nor U18763 (N_18763,N_17551,N_17399);
nand U18764 (N_18764,N_17495,N_17007);
and U18765 (N_18765,N_17121,N_17604);
nand U18766 (N_18766,N_17531,N_17333);
or U18767 (N_18767,N_17164,N_17873);
and U18768 (N_18768,N_17907,N_17092);
nand U18769 (N_18769,N_17589,N_17918);
xor U18770 (N_18770,N_17583,N_17661);
xor U18771 (N_18771,N_17036,N_17107);
and U18772 (N_18772,N_17370,N_17768);
and U18773 (N_18773,N_17804,N_17382);
xor U18774 (N_18774,N_17401,N_17539);
nor U18775 (N_18775,N_17720,N_17308);
xor U18776 (N_18776,N_17216,N_17525);
or U18777 (N_18777,N_17913,N_17200);
nand U18778 (N_18778,N_17691,N_17241);
and U18779 (N_18779,N_17135,N_17323);
nor U18780 (N_18780,N_17756,N_17656);
xor U18781 (N_18781,N_17990,N_17774);
nand U18782 (N_18782,N_17972,N_17240);
nor U18783 (N_18783,N_17110,N_17231);
and U18784 (N_18784,N_17122,N_17156);
nand U18785 (N_18785,N_17821,N_17952);
nor U18786 (N_18786,N_17981,N_17943);
nor U18787 (N_18787,N_17832,N_17779);
and U18788 (N_18788,N_17375,N_17891);
or U18789 (N_18789,N_17928,N_17750);
nand U18790 (N_18790,N_17504,N_17300);
nand U18791 (N_18791,N_17432,N_17894);
and U18792 (N_18792,N_17012,N_17596);
and U18793 (N_18793,N_17972,N_17740);
or U18794 (N_18794,N_17119,N_17846);
nand U18795 (N_18795,N_17535,N_17095);
and U18796 (N_18796,N_17217,N_17331);
nand U18797 (N_18797,N_17866,N_17967);
nor U18798 (N_18798,N_17502,N_17507);
xor U18799 (N_18799,N_17315,N_17244);
and U18800 (N_18800,N_17130,N_17539);
xnor U18801 (N_18801,N_17593,N_17914);
nor U18802 (N_18802,N_17966,N_17296);
or U18803 (N_18803,N_17515,N_17591);
and U18804 (N_18804,N_17038,N_17843);
xnor U18805 (N_18805,N_17110,N_17938);
nor U18806 (N_18806,N_17239,N_17784);
or U18807 (N_18807,N_17369,N_17515);
or U18808 (N_18808,N_17010,N_17239);
nand U18809 (N_18809,N_17707,N_17214);
or U18810 (N_18810,N_17797,N_17942);
or U18811 (N_18811,N_17462,N_17780);
or U18812 (N_18812,N_17251,N_17628);
and U18813 (N_18813,N_17949,N_17737);
nor U18814 (N_18814,N_17019,N_17753);
or U18815 (N_18815,N_17370,N_17262);
nand U18816 (N_18816,N_17616,N_17398);
xor U18817 (N_18817,N_17001,N_17749);
and U18818 (N_18818,N_17534,N_17742);
nor U18819 (N_18819,N_17144,N_17230);
and U18820 (N_18820,N_17676,N_17605);
xnor U18821 (N_18821,N_17745,N_17658);
or U18822 (N_18822,N_17456,N_17491);
nand U18823 (N_18823,N_17539,N_17018);
and U18824 (N_18824,N_17544,N_17912);
nand U18825 (N_18825,N_17209,N_17191);
or U18826 (N_18826,N_17355,N_17790);
and U18827 (N_18827,N_17057,N_17570);
or U18828 (N_18828,N_17281,N_17870);
and U18829 (N_18829,N_17202,N_17091);
xor U18830 (N_18830,N_17459,N_17363);
and U18831 (N_18831,N_17779,N_17078);
xnor U18832 (N_18832,N_17206,N_17663);
nor U18833 (N_18833,N_17181,N_17270);
or U18834 (N_18834,N_17298,N_17042);
and U18835 (N_18835,N_17077,N_17051);
and U18836 (N_18836,N_17953,N_17981);
xor U18837 (N_18837,N_17499,N_17564);
xor U18838 (N_18838,N_17306,N_17734);
or U18839 (N_18839,N_17970,N_17966);
nor U18840 (N_18840,N_17362,N_17959);
xnor U18841 (N_18841,N_17518,N_17541);
or U18842 (N_18842,N_17992,N_17801);
or U18843 (N_18843,N_17233,N_17187);
or U18844 (N_18844,N_17226,N_17502);
xnor U18845 (N_18845,N_17691,N_17336);
or U18846 (N_18846,N_17636,N_17344);
nand U18847 (N_18847,N_17276,N_17896);
nor U18848 (N_18848,N_17396,N_17238);
or U18849 (N_18849,N_17400,N_17753);
xnor U18850 (N_18850,N_17647,N_17885);
nand U18851 (N_18851,N_17307,N_17458);
nor U18852 (N_18852,N_17034,N_17981);
nand U18853 (N_18853,N_17340,N_17965);
nand U18854 (N_18854,N_17169,N_17930);
and U18855 (N_18855,N_17526,N_17540);
xor U18856 (N_18856,N_17837,N_17283);
xnor U18857 (N_18857,N_17851,N_17469);
xor U18858 (N_18858,N_17901,N_17976);
and U18859 (N_18859,N_17452,N_17596);
nor U18860 (N_18860,N_17048,N_17454);
xor U18861 (N_18861,N_17503,N_17322);
or U18862 (N_18862,N_17201,N_17191);
nand U18863 (N_18863,N_17805,N_17893);
nand U18864 (N_18864,N_17997,N_17885);
xor U18865 (N_18865,N_17217,N_17639);
and U18866 (N_18866,N_17092,N_17955);
or U18867 (N_18867,N_17342,N_17763);
and U18868 (N_18868,N_17578,N_17902);
and U18869 (N_18869,N_17401,N_17923);
nor U18870 (N_18870,N_17264,N_17387);
nor U18871 (N_18871,N_17974,N_17437);
xor U18872 (N_18872,N_17579,N_17113);
or U18873 (N_18873,N_17894,N_17163);
xnor U18874 (N_18874,N_17962,N_17040);
xnor U18875 (N_18875,N_17026,N_17297);
nand U18876 (N_18876,N_17586,N_17331);
or U18877 (N_18877,N_17757,N_17239);
and U18878 (N_18878,N_17258,N_17360);
nand U18879 (N_18879,N_17538,N_17831);
nand U18880 (N_18880,N_17512,N_17587);
and U18881 (N_18881,N_17459,N_17785);
nand U18882 (N_18882,N_17854,N_17157);
nor U18883 (N_18883,N_17610,N_17132);
and U18884 (N_18884,N_17592,N_17752);
xor U18885 (N_18885,N_17538,N_17877);
or U18886 (N_18886,N_17623,N_17807);
nand U18887 (N_18887,N_17451,N_17581);
or U18888 (N_18888,N_17766,N_17236);
and U18889 (N_18889,N_17428,N_17748);
nor U18890 (N_18890,N_17528,N_17821);
nor U18891 (N_18891,N_17462,N_17080);
or U18892 (N_18892,N_17977,N_17932);
xor U18893 (N_18893,N_17838,N_17622);
and U18894 (N_18894,N_17847,N_17031);
and U18895 (N_18895,N_17948,N_17658);
nor U18896 (N_18896,N_17498,N_17732);
and U18897 (N_18897,N_17934,N_17223);
and U18898 (N_18898,N_17237,N_17709);
and U18899 (N_18899,N_17380,N_17812);
nor U18900 (N_18900,N_17325,N_17007);
and U18901 (N_18901,N_17353,N_17614);
nor U18902 (N_18902,N_17263,N_17297);
nor U18903 (N_18903,N_17541,N_17627);
xnor U18904 (N_18904,N_17844,N_17302);
xor U18905 (N_18905,N_17405,N_17599);
nor U18906 (N_18906,N_17397,N_17828);
nor U18907 (N_18907,N_17517,N_17266);
xor U18908 (N_18908,N_17639,N_17293);
xnor U18909 (N_18909,N_17821,N_17343);
nor U18910 (N_18910,N_17999,N_17781);
xor U18911 (N_18911,N_17184,N_17092);
nor U18912 (N_18912,N_17393,N_17946);
nand U18913 (N_18913,N_17406,N_17278);
and U18914 (N_18914,N_17413,N_17965);
and U18915 (N_18915,N_17937,N_17266);
or U18916 (N_18916,N_17370,N_17743);
xnor U18917 (N_18917,N_17741,N_17012);
nand U18918 (N_18918,N_17896,N_17399);
nor U18919 (N_18919,N_17653,N_17052);
and U18920 (N_18920,N_17099,N_17077);
nand U18921 (N_18921,N_17180,N_17746);
nand U18922 (N_18922,N_17035,N_17820);
or U18923 (N_18923,N_17710,N_17393);
xnor U18924 (N_18924,N_17079,N_17228);
or U18925 (N_18925,N_17112,N_17438);
nand U18926 (N_18926,N_17670,N_17126);
nand U18927 (N_18927,N_17210,N_17474);
xor U18928 (N_18928,N_17770,N_17147);
or U18929 (N_18929,N_17748,N_17040);
and U18930 (N_18930,N_17637,N_17994);
xor U18931 (N_18931,N_17257,N_17408);
and U18932 (N_18932,N_17248,N_17849);
nand U18933 (N_18933,N_17842,N_17155);
nand U18934 (N_18934,N_17247,N_17228);
and U18935 (N_18935,N_17798,N_17731);
and U18936 (N_18936,N_17678,N_17747);
and U18937 (N_18937,N_17756,N_17545);
nor U18938 (N_18938,N_17626,N_17271);
and U18939 (N_18939,N_17531,N_17429);
or U18940 (N_18940,N_17759,N_17229);
and U18941 (N_18941,N_17105,N_17240);
xnor U18942 (N_18942,N_17194,N_17975);
and U18943 (N_18943,N_17394,N_17499);
nand U18944 (N_18944,N_17151,N_17150);
nor U18945 (N_18945,N_17279,N_17695);
nor U18946 (N_18946,N_17417,N_17683);
nor U18947 (N_18947,N_17229,N_17571);
nor U18948 (N_18948,N_17491,N_17344);
xor U18949 (N_18949,N_17768,N_17456);
xnor U18950 (N_18950,N_17798,N_17689);
xnor U18951 (N_18951,N_17462,N_17106);
or U18952 (N_18952,N_17876,N_17790);
nor U18953 (N_18953,N_17516,N_17361);
xor U18954 (N_18954,N_17321,N_17570);
nor U18955 (N_18955,N_17969,N_17945);
nor U18956 (N_18956,N_17981,N_17718);
nor U18957 (N_18957,N_17577,N_17276);
and U18958 (N_18958,N_17863,N_17784);
or U18959 (N_18959,N_17170,N_17435);
and U18960 (N_18960,N_17278,N_17043);
nand U18961 (N_18961,N_17086,N_17294);
and U18962 (N_18962,N_17499,N_17032);
or U18963 (N_18963,N_17688,N_17107);
and U18964 (N_18964,N_17383,N_17875);
xnor U18965 (N_18965,N_17855,N_17890);
xor U18966 (N_18966,N_17651,N_17596);
and U18967 (N_18967,N_17558,N_17957);
nand U18968 (N_18968,N_17848,N_17410);
nor U18969 (N_18969,N_17765,N_17909);
or U18970 (N_18970,N_17101,N_17293);
and U18971 (N_18971,N_17568,N_17873);
and U18972 (N_18972,N_17239,N_17507);
xnor U18973 (N_18973,N_17311,N_17148);
nor U18974 (N_18974,N_17474,N_17983);
or U18975 (N_18975,N_17058,N_17244);
and U18976 (N_18976,N_17222,N_17471);
xor U18977 (N_18977,N_17974,N_17997);
nor U18978 (N_18978,N_17490,N_17739);
xnor U18979 (N_18979,N_17123,N_17788);
xnor U18980 (N_18980,N_17675,N_17796);
nor U18981 (N_18981,N_17482,N_17784);
xor U18982 (N_18982,N_17848,N_17098);
and U18983 (N_18983,N_17246,N_17525);
nand U18984 (N_18984,N_17423,N_17799);
xnor U18985 (N_18985,N_17189,N_17467);
nand U18986 (N_18986,N_17812,N_17459);
nor U18987 (N_18987,N_17069,N_17880);
nor U18988 (N_18988,N_17718,N_17813);
xor U18989 (N_18989,N_17258,N_17136);
and U18990 (N_18990,N_17901,N_17599);
and U18991 (N_18991,N_17739,N_17986);
nor U18992 (N_18992,N_17275,N_17190);
nor U18993 (N_18993,N_17653,N_17177);
or U18994 (N_18994,N_17061,N_17145);
nand U18995 (N_18995,N_17944,N_17155);
nor U18996 (N_18996,N_17807,N_17133);
nand U18997 (N_18997,N_17522,N_17858);
nor U18998 (N_18998,N_17867,N_17495);
or U18999 (N_18999,N_17476,N_17258);
nand U19000 (N_19000,N_18919,N_18366);
nand U19001 (N_19001,N_18857,N_18827);
xor U19002 (N_19002,N_18218,N_18726);
nand U19003 (N_19003,N_18011,N_18182);
xor U19004 (N_19004,N_18341,N_18696);
or U19005 (N_19005,N_18718,N_18312);
and U19006 (N_19006,N_18727,N_18483);
xor U19007 (N_19007,N_18095,N_18323);
nand U19008 (N_19008,N_18743,N_18675);
and U19009 (N_19009,N_18789,N_18210);
nor U19010 (N_19010,N_18464,N_18353);
nand U19011 (N_19011,N_18206,N_18290);
nor U19012 (N_19012,N_18374,N_18269);
nor U19013 (N_19013,N_18546,N_18632);
or U19014 (N_19014,N_18503,N_18631);
and U19015 (N_19015,N_18902,N_18278);
or U19016 (N_19016,N_18669,N_18164);
xnor U19017 (N_19017,N_18895,N_18375);
xnor U19018 (N_19018,N_18547,N_18322);
nand U19019 (N_19019,N_18197,N_18015);
and U19020 (N_19020,N_18300,N_18404);
or U19021 (N_19021,N_18167,N_18746);
or U19022 (N_19022,N_18199,N_18814);
nand U19023 (N_19023,N_18180,N_18572);
xor U19024 (N_19024,N_18621,N_18087);
or U19025 (N_19025,N_18119,N_18472);
nand U19026 (N_19026,N_18660,N_18562);
or U19027 (N_19027,N_18338,N_18777);
xnor U19028 (N_19028,N_18220,N_18630);
or U19029 (N_19029,N_18122,N_18380);
xnor U19030 (N_19030,N_18608,N_18331);
xnor U19031 (N_19031,N_18448,N_18575);
and U19032 (N_19032,N_18779,N_18602);
nor U19033 (N_19033,N_18301,N_18420);
nor U19034 (N_19034,N_18767,N_18748);
and U19035 (N_19035,N_18279,N_18153);
and U19036 (N_19036,N_18392,N_18913);
and U19037 (N_19037,N_18930,N_18496);
or U19038 (N_19038,N_18633,N_18571);
nand U19039 (N_19039,N_18840,N_18057);
or U19040 (N_19040,N_18741,N_18401);
or U19041 (N_19041,N_18061,N_18173);
and U19042 (N_19042,N_18045,N_18983);
nor U19043 (N_19043,N_18558,N_18489);
nor U19044 (N_19044,N_18988,N_18155);
and U19045 (N_19045,N_18869,N_18202);
nand U19046 (N_19046,N_18710,N_18271);
nand U19047 (N_19047,N_18276,N_18280);
nor U19048 (N_19048,N_18358,N_18624);
and U19049 (N_19049,N_18993,N_18107);
nor U19050 (N_19050,N_18359,N_18788);
and U19051 (N_19051,N_18805,N_18591);
nor U19052 (N_19052,N_18021,N_18193);
and U19053 (N_19053,N_18260,N_18140);
nor U19054 (N_19054,N_18198,N_18294);
and U19055 (N_19055,N_18031,N_18683);
or U19056 (N_19056,N_18791,N_18931);
or U19057 (N_19057,N_18835,N_18717);
nor U19058 (N_19058,N_18085,N_18634);
xnor U19059 (N_19059,N_18352,N_18256);
and U19060 (N_19060,N_18311,N_18189);
xor U19061 (N_19061,N_18695,N_18399);
nor U19062 (N_19062,N_18272,N_18787);
nor U19063 (N_19063,N_18798,N_18561);
or U19064 (N_19064,N_18918,N_18247);
xnor U19065 (N_19065,N_18491,N_18243);
or U19066 (N_19066,N_18022,N_18810);
or U19067 (N_19067,N_18690,N_18679);
or U19068 (N_19068,N_18775,N_18136);
nor U19069 (N_19069,N_18953,N_18487);
and U19070 (N_19070,N_18668,N_18349);
or U19071 (N_19071,N_18543,N_18288);
xor U19072 (N_19072,N_18772,N_18151);
and U19073 (N_19073,N_18365,N_18172);
or U19074 (N_19074,N_18860,N_18117);
and U19075 (N_19075,N_18799,N_18568);
and U19076 (N_19076,N_18043,N_18008);
nand U19077 (N_19077,N_18653,N_18815);
xor U19078 (N_19078,N_18019,N_18490);
nor U19079 (N_19079,N_18262,N_18523);
xor U19080 (N_19080,N_18701,N_18509);
nand U19081 (N_19081,N_18177,N_18030);
or U19082 (N_19082,N_18549,N_18601);
and U19083 (N_19083,N_18314,N_18285);
nand U19084 (N_19084,N_18398,N_18332);
or U19085 (N_19085,N_18208,N_18303);
nand U19086 (N_19086,N_18744,N_18065);
xor U19087 (N_19087,N_18124,N_18093);
xnor U19088 (N_19088,N_18098,N_18733);
or U19089 (N_19089,N_18101,N_18966);
and U19090 (N_19090,N_18094,N_18284);
and U19091 (N_19091,N_18148,N_18475);
xor U19092 (N_19092,N_18364,N_18405);
or U19093 (N_19093,N_18765,N_18152);
nand U19094 (N_19094,N_18028,N_18510);
and U19095 (N_19095,N_18872,N_18935);
xor U19096 (N_19096,N_18335,N_18035);
nor U19097 (N_19097,N_18986,N_18644);
xnor U19098 (N_19098,N_18051,N_18379);
nand U19099 (N_19099,N_18736,N_18059);
or U19100 (N_19100,N_18427,N_18821);
nand U19101 (N_19101,N_18006,N_18126);
and U19102 (N_19102,N_18830,N_18563);
and U19103 (N_19103,N_18014,N_18474);
and U19104 (N_19104,N_18424,N_18909);
or U19105 (N_19105,N_18944,N_18952);
or U19106 (N_19106,N_18688,N_18064);
nand U19107 (N_19107,N_18992,N_18072);
nand U19108 (N_19108,N_18654,N_18264);
nand U19109 (N_19109,N_18881,N_18397);
nor U19110 (N_19110,N_18773,N_18851);
or U19111 (N_19111,N_18071,N_18443);
xnor U19112 (N_19112,N_18003,N_18484);
xnor U19113 (N_19113,N_18305,N_18808);
or U19114 (N_19114,N_18975,N_18212);
or U19115 (N_19115,N_18712,N_18223);
xor U19116 (N_19116,N_18069,N_18998);
nand U19117 (N_19117,N_18730,N_18048);
nor U19118 (N_19118,N_18425,N_18382);
xnor U19119 (N_19119,N_18393,N_18056);
nand U19120 (N_19120,N_18747,N_18135);
and U19121 (N_19121,N_18402,N_18336);
and U19122 (N_19122,N_18261,N_18482);
and U19123 (N_19123,N_18343,N_18987);
or U19124 (N_19124,N_18234,N_18979);
or U19125 (N_19125,N_18948,N_18273);
nand U19126 (N_19126,N_18797,N_18333);
nor U19127 (N_19127,N_18978,N_18384);
xor U19128 (N_19128,N_18159,N_18831);
or U19129 (N_19129,N_18565,N_18586);
nor U19130 (N_19130,N_18694,N_18873);
nor U19131 (N_19131,N_18502,N_18409);
nand U19132 (N_19132,N_18004,N_18096);
nand U19133 (N_19133,N_18242,N_18149);
nand U19134 (N_19134,N_18850,N_18699);
nor U19135 (N_19135,N_18629,N_18722);
nor U19136 (N_19136,N_18592,N_18689);
nor U19137 (N_19137,N_18617,N_18583);
nand U19138 (N_19138,N_18837,N_18790);
nand U19139 (N_19139,N_18698,N_18046);
xnor U19140 (N_19140,N_18974,N_18756);
xor U19141 (N_19141,N_18897,N_18680);
xor U19142 (N_19142,N_18517,N_18664);
nand U19143 (N_19143,N_18326,N_18864);
xnor U19144 (N_19144,N_18761,N_18406);
nor U19145 (N_19145,N_18597,N_18967);
and U19146 (N_19146,N_18697,N_18954);
or U19147 (N_19147,N_18950,N_18934);
xor U19148 (N_19148,N_18169,N_18268);
and U19149 (N_19149,N_18745,N_18876);
nand U19150 (N_19150,N_18859,N_18686);
and U19151 (N_19151,N_18054,N_18800);
nor U19152 (N_19152,N_18070,N_18351);
and U19153 (N_19153,N_18267,N_18762);
xnor U19154 (N_19154,N_18481,N_18076);
or U19155 (N_19155,N_18113,N_18504);
or U19156 (N_19156,N_18163,N_18663);
nor U19157 (N_19157,N_18754,N_18002);
or U19158 (N_19158,N_18385,N_18099);
or U19159 (N_19159,N_18838,N_18829);
or U19160 (N_19160,N_18582,N_18204);
or U19161 (N_19161,N_18622,N_18053);
or U19162 (N_19162,N_18104,N_18457);
nor U19163 (N_19163,N_18520,N_18593);
or U19164 (N_19164,N_18982,N_18783);
nand U19165 (N_19165,N_18228,N_18714);
or U19166 (N_19166,N_18647,N_18346);
or U19167 (N_19167,N_18729,N_18728);
xnor U19168 (N_19168,N_18885,N_18186);
xnor U19169 (N_19169,N_18758,N_18009);
or U19170 (N_19170,N_18190,N_18903);
and U19171 (N_19171,N_18479,N_18657);
nand U19172 (N_19172,N_18996,N_18058);
nor U19173 (N_19173,N_18465,N_18700);
and U19174 (N_19174,N_18020,N_18943);
or U19175 (N_19175,N_18068,N_18893);
or U19176 (N_19176,N_18626,N_18347);
or U19177 (N_19177,N_18802,N_18554);
and U19178 (N_19178,N_18555,N_18038);
or U19179 (N_19179,N_18154,N_18102);
or U19180 (N_19180,N_18032,N_18492);
or U19181 (N_19181,N_18682,N_18445);
and U19182 (N_19182,N_18957,N_18413);
nor U19183 (N_19183,N_18759,N_18047);
and U19184 (N_19184,N_18086,N_18209);
xnor U19185 (N_19185,N_18388,N_18125);
nor U19186 (N_19186,N_18920,N_18486);
and U19187 (N_19187,N_18693,N_18073);
nor U19188 (N_19188,N_18620,N_18970);
xor U19189 (N_19189,N_18883,N_18027);
and U19190 (N_19190,N_18213,N_18557);
or U19191 (N_19191,N_18141,N_18131);
and U19192 (N_19192,N_18577,N_18360);
nor U19193 (N_19193,N_18587,N_18116);
and U19194 (N_19194,N_18369,N_18599);
xor U19195 (N_19195,N_18725,N_18853);
nor U19196 (N_19196,N_18991,N_18812);
xor U19197 (N_19197,N_18016,N_18412);
xnor U19198 (N_19198,N_18438,N_18614);
or U19199 (N_19199,N_18877,N_18940);
or U19200 (N_19200,N_18144,N_18778);
xor U19201 (N_19201,N_18636,N_18724);
nor U19202 (N_19202,N_18478,N_18844);
or U19203 (N_19203,N_18786,N_18833);
and U19204 (N_19204,N_18033,N_18329);
nand U19205 (N_19205,N_18922,N_18738);
or U19206 (N_19206,N_18249,N_18550);
or U19207 (N_19207,N_18569,N_18961);
or U19208 (N_19208,N_18176,N_18801);
nor U19209 (N_19209,N_18171,N_18731);
xor U19210 (N_19210,N_18477,N_18536);
nand U19211 (N_19211,N_18292,N_18973);
xnor U19212 (N_19212,N_18884,N_18556);
xnor U19213 (N_19213,N_18062,N_18133);
nor U19214 (N_19214,N_18342,N_18936);
nand U19215 (N_19215,N_18255,N_18795);
nand U19216 (N_19216,N_18813,N_18981);
nand U19217 (N_19217,N_18063,N_18105);
nor U19218 (N_19218,N_18834,N_18676);
nand U19219 (N_19219,N_18236,N_18941);
nor U19220 (N_19220,N_18115,N_18960);
nand U19221 (N_19221,N_18755,N_18611);
xnor U19222 (N_19222,N_18766,N_18108);
nand U19223 (N_19223,N_18473,N_18867);
nor U19224 (N_19224,N_18499,N_18408);
nor U19225 (N_19225,N_18244,N_18146);
and U19226 (N_19226,N_18692,N_18422);
and U19227 (N_19227,N_18447,N_18764);
nor U19228 (N_19228,N_18110,N_18560);
xnor U19229 (N_19229,N_18576,N_18304);
xor U19230 (N_19230,N_18715,N_18354);
nor U19231 (N_19231,N_18836,N_18887);
nand U19232 (N_19232,N_18559,N_18917);
nand U19233 (N_19233,N_18911,N_18532);
or U19234 (N_19234,N_18650,N_18013);
or U19235 (N_19235,N_18250,N_18513);
nor U19236 (N_19236,N_18946,N_18299);
and U19237 (N_19237,N_18367,N_18429);
xnor U19238 (N_19238,N_18528,N_18187);
and U19239 (N_19239,N_18892,N_18763);
xnor U19240 (N_19240,N_18395,N_18589);
nand U19241 (N_19241,N_18253,N_18955);
or U19242 (N_19242,N_18678,N_18460);
nor U19243 (N_19243,N_18120,N_18564);
and U19244 (N_19244,N_18515,N_18407);
and U19245 (N_19245,N_18390,N_18471);
or U19246 (N_19246,N_18861,N_18753);
nand U19247 (N_19247,N_18822,N_18868);
xnor U19248 (N_19248,N_18286,N_18453);
nand U19249 (N_19249,N_18307,N_18495);
nor U19250 (N_19250,N_18709,N_18656);
nand U19251 (N_19251,N_18348,N_18467);
and U19252 (N_19252,N_18325,N_18672);
xnor U19253 (N_19253,N_18450,N_18605);
xnor U19254 (N_19254,N_18681,N_18588);
or U19255 (N_19255,N_18316,N_18646);
or U19256 (N_19256,N_18277,N_18452);
nor U19257 (N_19257,N_18553,N_18449);
xnor U19258 (N_19258,N_18968,N_18820);
or U19259 (N_19259,N_18103,N_18241);
and U19260 (N_19260,N_18426,N_18328);
nand U19261 (N_19261,N_18649,N_18114);
nand U19262 (N_19262,N_18055,N_18990);
nand U19263 (N_19263,N_18781,N_18995);
or U19264 (N_19264,N_18324,N_18356);
and U19265 (N_19265,N_18188,N_18081);
or U19266 (N_19266,N_18079,N_18078);
nand U19267 (N_19267,N_18886,N_18924);
xnor U19268 (N_19268,N_18904,N_18196);
or U19269 (N_19269,N_18265,N_18372);
nand U19270 (N_19270,N_18907,N_18889);
or U19271 (N_19271,N_18371,N_18052);
or U19272 (N_19272,N_18616,N_18123);
nand U19273 (N_19273,N_18252,N_18421);
nand U19274 (N_19274,N_18642,N_18809);
or U19275 (N_19275,N_18819,N_18157);
or U19276 (N_19276,N_18293,N_18824);
nand U19277 (N_19277,N_18742,N_18514);
nor U19278 (N_19278,N_18932,N_18283);
xnor U19279 (N_19279,N_18604,N_18428);
xor U19280 (N_19280,N_18468,N_18227);
xor U19281 (N_19281,N_18685,N_18165);
or U19282 (N_19282,N_18965,N_18898);
nor U19283 (N_19283,N_18084,N_18309);
nor U19284 (N_19284,N_18274,N_18923);
xor U19285 (N_19285,N_18240,N_18900);
nor U19286 (N_19286,N_18410,N_18839);
and U19287 (N_19287,N_18376,N_18574);
and U19288 (N_19288,N_18205,N_18702);
and U19289 (N_19289,N_18541,N_18036);
or U19290 (N_19290,N_18044,N_18050);
nor U19291 (N_19291,N_18615,N_18089);
xnor U19292 (N_19292,N_18512,N_18083);
or U19293 (N_19293,N_18842,N_18221);
nand U19294 (N_19294,N_18908,N_18925);
nand U19295 (N_19295,N_18436,N_18355);
and U19296 (N_19296,N_18544,N_18259);
xnor U19297 (N_19297,N_18871,N_18566);
or U19298 (N_19298,N_18750,N_18785);
nand U19299 (N_19299,N_18161,N_18999);
or U19300 (N_19300,N_18581,N_18201);
or U19301 (N_19301,N_18012,N_18000);
and U19302 (N_19302,N_18217,N_18958);
or U19303 (N_19303,N_18458,N_18927);
and U19304 (N_19304,N_18846,N_18191);
or U19305 (N_19305,N_18807,N_18915);
and U19306 (N_19306,N_18378,N_18929);
or U19307 (N_19307,N_18441,N_18381);
xnor U19308 (N_19308,N_18508,N_18570);
nor U19309 (N_19309,N_18875,N_18854);
and U19310 (N_19310,N_18075,N_18803);
or U19311 (N_19311,N_18832,N_18112);
nand U19312 (N_19312,N_18841,N_18901);
and U19313 (N_19313,N_18878,N_18295);
or U19314 (N_19314,N_18818,N_18655);
or U19315 (N_19315,N_18129,N_18207);
nand U19316 (N_19316,N_18315,N_18529);
nor U19317 (N_19317,N_18670,N_18239);
nor U19318 (N_19318,N_18118,N_18548);
nand U19319 (N_19319,N_18383,N_18005);
or U19320 (N_19320,N_18039,N_18708);
or U19321 (N_19321,N_18363,N_18147);
xor U19322 (N_19322,N_18488,N_18308);
and U19323 (N_19323,N_18962,N_18567);
nand U19324 (N_19324,N_18029,N_18551);
nand U19325 (N_19325,N_18432,N_18266);
xnor U19326 (N_19326,N_18185,N_18752);
xor U19327 (N_19327,N_18297,N_18034);
xnor U19328 (N_19328,N_18370,N_18691);
nor U19329 (N_19329,N_18825,N_18435);
nor U19330 (N_19330,N_18454,N_18879);
nor U19331 (N_19331,N_18880,N_18628);
nor U19332 (N_19332,N_18639,N_18142);
xnor U19333 (N_19333,N_18769,N_18721);
nand U19334 (N_19334,N_18519,N_18439);
nor U19335 (N_19335,N_18442,N_18640);
nor U19336 (N_19336,N_18178,N_18313);
nor U19337 (N_19337,N_18001,N_18989);
nand U19338 (N_19338,N_18462,N_18320);
or U19339 (N_19339,N_18774,N_18446);
and U19340 (N_19340,N_18673,N_18501);
or U19341 (N_19341,N_18362,N_18156);
or U19342 (N_19342,N_18806,N_18166);
xnor U19343 (N_19343,N_18826,N_18476);
nor U19344 (N_19344,N_18852,N_18132);
xnor U19345 (N_19345,N_18912,N_18216);
or U19346 (N_19346,N_18828,N_18684);
xnor U19347 (N_19347,N_18430,N_18947);
and U19348 (N_19348,N_18150,N_18662);
and U19349 (N_19349,N_18985,N_18776);
or U19350 (N_19350,N_18074,N_18984);
xor U19351 (N_19351,N_18711,N_18192);
nor U19352 (N_19352,N_18100,N_18179);
xor U19353 (N_19353,N_18905,N_18470);
xnor U19354 (N_19354,N_18246,N_18600);
xor U19355 (N_19355,N_18796,N_18933);
xnor U19356 (N_19356,N_18373,N_18749);
nor U19357 (N_19357,N_18494,N_18254);
nand U19358 (N_19358,N_18067,N_18232);
nor U19359 (N_19359,N_18926,N_18637);
nor U19360 (N_19360,N_18431,N_18534);
nand U19361 (N_19361,N_18230,N_18782);
or U19362 (N_19362,N_18317,N_18461);
and U19363 (N_19363,N_18263,N_18394);
or U19364 (N_19364,N_18545,N_18040);
nand U19365 (N_19365,N_18651,N_18882);
or U19366 (N_19366,N_18526,N_18584);
nor U19367 (N_19367,N_18865,N_18235);
or U19368 (N_19368,N_18097,N_18816);
and U19369 (N_19369,N_18906,N_18951);
and U19370 (N_19370,N_18321,N_18848);
nor U19371 (N_19371,N_18456,N_18914);
and U19372 (N_19372,N_18258,N_18768);
and U19373 (N_19373,N_18870,N_18862);
and U19374 (N_19374,N_18419,N_18891);
or U19375 (N_19375,N_18652,N_18007);
nor U19376 (N_19376,N_18181,N_18527);
or U19377 (N_19377,N_18916,N_18275);
and U19378 (N_19378,N_18677,N_18257);
or U19379 (N_19379,N_18340,N_18337);
nand U19380 (N_19380,N_18018,N_18770);
and U19381 (N_19381,N_18368,N_18585);
nor U19382 (N_19382,N_18183,N_18713);
or U19383 (N_19383,N_18158,N_18506);
or U19384 (N_19384,N_18847,N_18010);
or U19385 (N_19385,N_18200,N_18145);
xnor U19386 (N_19386,N_18345,N_18080);
or U19387 (N_19387,N_18792,N_18418);
and U19388 (N_19388,N_18455,N_18480);
nor U19389 (N_19389,N_18469,N_18451);
and U19390 (N_19390,N_18623,N_18938);
and U19391 (N_19391,N_18739,N_18433);
nor U19392 (N_19392,N_18175,N_18434);
xnor U19393 (N_19393,N_18823,N_18899);
xor U19394 (N_19394,N_18088,N_18703);
nand U19395 (N_19395,N_18327,N_18521);
xor U19396 (N_19396,N_18737,N_18863);
or U19397 (N_19397,N_18440,N_18524);
or U19398 (N_19398,N_18910,N_18598);
nor U19399 (N_19399,N_18849,N_18289);
and U19400 (N_19400,N_18516,N_18195);
nor U19401 (N_19401,N_18139,N_18194);
xnor U19402 (N_19402,N_18606,N_18302);
nand U19403 (N_19403,N_18665,N_18498);
and U19404 (N_19404,N_18972,N_18444);
and U19405 (N_19405,N_18077,N_18666);
nor U19406 (N_19406,N_18607,N_18511);
xor U19407 (N_19407,N_18416,N_18411);
nor U19408 (N_19408,N_18248,N_18595);
or U19409 (N_19409,N_18287,N_18757);
or U19410 (N_19410,N_18579,N_18310);
and U19411 (N_19411,N_18856,N_18414);
nand U19412 (N_19412,N_18613,N_18705);
and U19413 (N_19413,N_18091,N_18533);
or U19414 (N_19414,N_18760,N_18270);
nor U19415 (N_19415,N_18535,N_18997);
xnor U19416 (N_19416,N_18659,N_18518);
and U19417 (N_19417,N_18794,N_18531);
and U19418 (N_19418,N_18386,N_18580);
xnor U19419 (N_19419,N_18638,N_18603);
and U19420 (N_19420,N_18224,N_18658);
nor U19421 (N_19421,N_18130,N_18716);
and U19422 (N_19422,N_18890,N_18609);
nor U19423 (N_19423,N_18921,N_18066);
and U19424 (N_19424,N_18811,N_18391);
nor U19425 (N_19425,N_18400,N_18214);
nor U19426 (N_19426,N_18160,N_18466);
xnor U19427 (N_19427,N_18578,N_18222);
nand U19428 (N_19428,N_18417,N_18229);
and U19429 (N_19429,N_18596,N_18121);
nor U19430 (N_19430,N_18537,N_18625);
and U19431 (N_19431,N_18771,N_18497);
and U19432 (N_19432,N_18437,N_18874);
and U19433 (N_19433,N_18784,N_18855);
nor U19434 (N_19434,N_18706,N_18858);
nand U19435 (N_19435,N_18971,N_18361);
nor U19436 (N_19436,N_18648,N_18318);
nand U19437 (N_19437,N_18894,N_18994);
nor U19438 (N_19438,N_18845,N_18866);
and U19439 (N_19439,N_18319,N_18538);
xor U19440 (N_19440,N_18671,N_18026);
and U19441 (N_19441,N_18357,N_18162);
nor U19442 (N_19442,N_18463,N_18704);
xor U19443 (N_19443,N_18415,N_18111);
and U19444 (N_19444,N_18023,N_18281);
nand U19445 (N_19445,N_18896,N_18339);
nand U19446 (N_19446,N_18233,N_18674);
nand U19447 (N_19447,N_18540,N_18720);
xnor U19448 (N_19448,N_18049,N_18377);
nand U19449 (N_19449,N_18937,N_18522);
or U19450 (N_19450,N_18667,N_18344);
and U19451 (N_19451,N_18949,N_18751);
or U19452 (N_19452,N_18928,N_18612);
nor U19453 (N_19453,N_18459,N_18500);
nor U19454 (N_19454,N_18530,N_18219);
nand U19455 (N_19455,N_18942,N_18888);
xor U19456 (N_19456,N_18184,N_18389);
nor U19457 (N_19457,N_18025,N_18485);
and U19458 (N_19458,N_18168,N_18939);
nand U19459 (N_19459,N_18817,N_18734);
and U19460 (N_19460,N_18945,N_18618);
and U19461 (N_19461,N_18641,N_18134);
nor U19462 (N_19462,N_18017,N_18963);
and U19463 (N_19463,N_18396,N_18170);
xor U19464 (N_19464,N_18610,N_18956);
or U19465 (N_19465,N_18143,N_18505);
nand U19466 (N_19466,N_18330,N_18843);
xnor U19467 (N_19467,N_18296,N_18215);
or U19468 (N_19468,N_18635,N_18306);
or U19469 (N_19469,N_18707,N_18423);
and U19470 (N_19470,N_18282,N_18226);
nor U19471 (N_19471,N_18291,N_18387);
xnor U19472 (N_19472,N_18174,N_18037);
and U19473 (N_19473,N_18251,N_18334);
xor U19474 (N_19474,N_18128,N_18127);
xor U19475 (N_19475,N_18542,N_18060);
and U19476 (N_19476,N_18959,N_18661);
xnor U19477 (N_19477,N_18627,N_18507);
and U19478 (N_19478,N_18719,N_18024);
and U19479 (N_19479,N_18594,N_18793);
xor U19480 (N_19480,N_18735,N_18041);
nor U19481 (N_19481,N_18964,N_18298);
nor U19482 (N_19482,N_18619,N_18245);
nand U19483 (N_19483,N_18977,N_18138);
nor U19484 (N_19484,N_18109,N_18238);
or U19485 (N_19485,N_18573,N_18082);
or U19486 (N_19486,N_18552,N_18780);
nor U19487 (N_19487,N_18723,N_18645);
nor U19488 (N_19488,N_18092,N_18350);
and U19489 (N_19489,N_18643,N_18137);
and U19490 (N_19490,N_18804,N_18590);
nand U19491 (N_19491,N_18969,N_18732);
and U19492 (N_19492,N_18980,N_18493);
xnor U19493 (N_19493,N_18403,N_18090);
nand U19494 (N_19494,N_18203,N_18225);
nand U19495 (N_19495,N_18106,N_18211);
nand U19496 (N_19496,N_18687,N_18740);
xor U19497 (N_19497,N_18042,N_18525);
xor U19498 (N_19498,N_18539,N_18231);
or U19499 (N_19499,N_18237,N_18976);
xor U19500 (N_19500,N_18893,N_18581);
and U19501 (N_19501,N_18854,N_18786);
xnor U19502 (N_19502,N_18783,N_18908);
nand U19503 (N_19503,N_18293,N_18018);
and U19504 (N_19504,N_18379,N_18754);
or U19505 (N_19505,N_18967,N_18413);
nand U19506 (N_19506,N_18865,N_18556);
xnor U19507 (N_19507,N_18967,N_18067);
nand U19508 (N_19508,N_18622,N_18377);
and U19509 (N_19509,N_18736,N_18804);
or U19510 (N_19510,N_18031,N_18941);
nor U19511 (N_19511,N_18754,N_18523);
nor U19512 (N_19512,N_18001,N_18287);
nand U19513 (N_19513,N_18003,N_18792);
nand U19514 (N_19514,N_18093,N_18996);
xnor U19515 (N_19515,N_18508,N_18706);
or U19516 (N_19516,N_18191,N_18708);
nor U19517 (N_19517,N_18967,N_18821);
nand U19518 (N_19518,N_18727,N_18722);
or U19519 (N_19519,N_18061,N_18456);
nor U19520 (N_19520,N_18980,N_18003);
and U19521 (N_19521,N_18681,N_18668);
nor U19522 (N_19522,N_18070,N_18085);
or U19523 (N_19523,N_18184,N_18073);
nor U19524 (N_19524,N_18074,N_18385);
nor U19525 (N_19525,N_18898,N_18267);
xnor U19526 (N_19526,N_18767,N_18316);
nand U19527 (N_19527,N_18114,N_18934);
xor U19528 (N_19528,N_18802,N_18507);
and U19529 (N_19529,N_18063,N_18033);
nand U19530 (N_19530,N_18174,N_18530);
nor U19531 (N_19531,N_18159,N_18152);
nor U19532 (N_19532,N_18315,N_18450);
xor U19533 (N_19533,N_18097,N_18215);
or U19534 (N_19534,N_18477,N_18143);
nor U19535 (N_19535,N_18614,N_18264);
or U19536 (N_19536,N_18233,N_18185);
and U19537 (N_19537,N_18405,N_18302);
xor U19538 (N_19538,N_18250,N_18632);
xnor U19539 (N_19539,N_18361,N_18143);
nand U19540 (N_19540,N_18261,N_18685);
and U19541 (N_19541,N_18218,N_18903);
xor U19542 (N_19542,N_18540,N_18241);
and U19543 (N_19543,N_18333,N_18653);
nand U19544 (N_19544,N_18775,N_18930);
nand U19545 (N_19545,N_18051,N_18030);
xnor U19546 (N_19546,N_18813,N_18561);
or U19547 (N_19547,N_18451,N_18258);
xnor U19548 (N_19548,N_18966,N_18571);
nor U19549 (N_19549,N_18295,N_18243);
nor U19550 (N_19550,N_18874,N_18404);
or U19551 (N_19551,N_18285,N_18599);
or U19552 (N_19552,N_18206,N_18365);
nand U19553 (N_19553,N_18717,N_18599);
and U19554 (N_19554,N_18596,N_18867);
xnor U19555 (N_19555,N_18413,N_18631);
or U19556 (N_19556,N_18807,N_18350);
xor U19557 (N_19557,N_18974,N_18385);
xnor U19558 (N_19558,N_18055,N_18798);
xnor U19559 (N_19559,N_18789,N_18066);
or U19560 (N_19560,N_18300,N_18095);
and U19561 (N_19561,N_18304,N_18499);
nand U19562 (N_19562,N_18599,N_18669);
nor U19563 (N_19563,N_18627,N_18372);
nand U19564 (N_19564,N_18486,N_18913);
nand U19565 (N_19565,N_18136,N_18934);
or U19566 (N_19566,N_18980,N_18767);
nand U19567 (N_19567,N_18920,N_18038);
and U19568 (N_19568,N_18859,N_18702);
or U19569 (N_19569,N_18694,N_18889);
nor U19570 (N_19570,N_18718,N_18005);
and U19571 (N_19571,N_18075,N_18878);
nor U19572 (N_19572,N_18540,N_18576);
nand U19573 (N_19573,N_18632,N_18462);
xnor U19574 (N_19574,N_18486,N_18260);
xnor U19575 (N_19575,N_18893,N_18597);
and U19576 (N_19576,N_18371,N_18623);
and U19577 (N_19577,N_18070,N_18778);
or U19578 (N_19578,N_18690,N_18066);
xor U19579 (N_19579,N_18149,N_18441);
and U19580 (N_19580,N_18568,N_18293);
xor U19581 (N_19581,N_18361,N_18038);
nand U19582 (N_19582,N_18444,N_18996);
nand U19583 (N_19583,N_18280,N_18839);
nor U19584 (N_19584,N_18855,N_18386);
xnor U19585 (N_19585,N_18386,N_18017);
nand U19586 (N_19586,N_18873,N_18470);
nand U19587 (N_19587,N_18374,N_18991);
nand U19588 (N_19588,N_18170,N_18859);
and U19589 (N_19589,N_18122,N_18978);
or U19590 (N_19590,N_18530,N_18813);
xor U19591 (N_19591,N_18407,N_18687);
or U19592 (N_19592,N_18484,N_18648);
nor U19593 (N_19593,N_18813,N_18760);
and U19594 (N_19594,N_18228,N_18846);
nand U19595 (N_19595,N_18453,N_18441);
nor U19596 (N_19596,N_18886,N_18083);
or U19597 (N_19597,N_18065,N_18494);
xor U19598 (N_19598,N_18151,N_18276);
nor U19599 (N_19599,N_18845,N_18150);
nand U19600 (N_19600,N_18979,N_18943);
and U19601 (N_19601,N_18731,N_18588);
xnor U19602 (N_19602,N_18673,N_18942);
or U19603 (N_19603,N_18924,N_18001);
nand U19604 (N_19604,N_18214,N_18859);
nand U19605 (N_19605,N_18629,N_18688);
and U19606 (N_19606,N_18910,N_18666);
or U19607 (N_19607,N_18965,N_18838);
nand U19608 (N_19608,N_18967,N_18692);
and U19609 (N_19609,N_18604,N_18182);
nor U19610 (N_19610,N_18515,N_18634);
nor U19611 (N_19611,N_18555,N_18321);
nand U19612 (N_19612,N_18198,N_18943);
and U19613 (N_19613,N_18144,N_18837);
nor U19614 (N_19614,N_18524,N_18442);
and U19615 (N_19615,N_18530,N_18762);
xnor U19616 (N_19616,N_18290,N_18147);
nand U19617 (N_19617,N_18980,N_18532);
and U19618 (N_19618,N_18346,N_18278);
xor U19619 (N_19619,N_18694,N_18020);
xor U19620 (N_19620,N_18038,N_18189);
xor U19621 (N_19621,N_18482,N_18072);
nand U19622 (N_19622,N_18935,N_18551);
xor U19623 (N_19623,N_18275,N_18402);
nand U19624 (N_19624,N_18072,N_18562);
or U19625 (N_19625,N_18447,N_18689);
xor U19626 (N_19626,N_18460,N_18005);
nand U19627 (N_19627,N_18980,N_18471);
nand U19628 (N_19628,N_18492,N_18788);
or U19629 (N_19629,N_18182,N_18334);
nand U19630 (N_19630,N_18654,N_18802);
nor U19631 (N_19631,N_18862,N_18049);
xor U19632 (N_19632,N_18421,N_18051);
and U19633 (N_19633,N_18001,N_18629);
and U19634 (N_19634,N_18310,N_18961);
nand U19635 (N_19635,N_18057,N_18567);
xnor U19636 (N_19636,N_18380,N_18771);
nand U19637 (N_19637,N_18050,N_18532);
and U19638 (N_19638,N_18207,N_18218);
or U19639 (N_19639,N_18705,N_18496);
or U19640 (N_19640,N_18143,N_18479);
nand U19641 (N_19641,N_18249,N_18818);
xnor U19642 (N_19642,N_18479,N_18737);
nor U19643 (N_19643,N_18238,N_18042);
nor U19644 (N_19644,N_18372,N_18695);
and U19645 (N_19645,N_18876,N_18600);
xor U19646 (N_19646,N_18680,N_18641);
and U19647 (N_19647,N_18376,N_18745);
nand U19648 (N_19648,N_18060,N_18136);
nand U19649 (N_19649,N_18646,N_18175);
or U19650 (N_19650,N_18906,N_18202);
and U19651 (N_19651,N_18793,N_18308);
xor U19652 (N_19652,N_18653,N_18747);
and U19653 (N_19653,N_18908,N_18920);
nor U19654 (N_19654,N_18261,N_18993);
or U19655 (N_19655,N_18084,N_18645);
and U19656 (N_19656,N_18986,N_18882);
nand U19657 (N_19657,N_18101,N_18193);
or U19658 (N_19658,N_18031,N_18462);
nand U19659 (N_19659,N_18251,N_18657);
nand U19660 (N_19660,N_18713,N_18393);
or U19661 (N_19661,N_18083,N_18013);
nand U19662 (N_19662,N_18783,N_18343);
or U19663 (N_19663,N_18595,N_18639);
and U19664 (N_19664,N_18818,N_18918);
nand U19665 (N_19665,N_18412,N_18474);
nand U19666 (N_19666,N_18040,N_18280);
or U19667 (N_19667,N_18949,N_18931);
nand U19668 (N_19668,N_18701,N_18054);
or U19669 (N_19669,N_18214,N_18675);
or U19670 (N_19670,N_18921,N_18498);
xnor U19671 (N_19671,N_18570,N_18150);
nand U19672 (N_19672,N_18914,N_18330);
or U19673 (N_19673,N_18916,N_18155);
xor U19674 (N_19674,N_18311,N_18019);
nand U19675 (N_19675,N_18343,N_18993);
or U19676 (N_19676,N_18368,N_18358);
xor U19677 (N_19677,N_18238,N_18529);
and U19678 (N_19678,N_18524,N_18749);
xor U19679 (N_19679,N_18399,N_18198);
nand U19680 (N_19680,N_18833,N_18138);
and U19681 (N_19681,N_18296,N_18632);
and U19682 (N_19682,N_18161,N_18462);
nand U19683 (N_19683,N_18099,N_18459);
or U19684 (N_19684,N_18073,N_18818);
xor U19685 (N_19685,N_18083,N_18854);
and U19686 (N_19686,N_18863,N_18349);
nand U19687 (N_19687,N_18552,N_18193);
and U19688 (N_19688,N_18476,N_18494);
or U19689 (N_19689,N_18320,N_18673);
xnor U19690 (N_19690,N_18495,N_18116);
xor U19691 (N_19691,N_18563,N_18557);
nand U19692 (N_19692,N_18330,N_18195);
nand U19693 (N_19693,N_18648,N_18461);
xnor U19694 (N_19694,N_18701,N_18385);
xnor U19695 (N_19695,N_18561,N_18480);
nand U19696 (N_19696,N_18839,N_18601);
nor U19697 (N_19697,N_18081,N_18722);
and U19698 (N_19698,N_18730,N_18843);
nand U19699 (N_19699,N_18900,N_18448);
xnor U19700 (N_19700,N_18191,N_18895);
and U19701 (N_19701,N_18026,N_18299);
or U19702 (N_19702,N_18440,N_18172);
xor U19703 (N_19703,N_18336,N_18373);
or U19704 (N_19704,N_18911,N_18971);
or U19705 (N_19705,N_18002,N_18631);
nand U19706 (N_19706,N_18902,N_18441);
xor U19707 (N_19707,N_18499,N_18780);
nand U19708 (N_19708,N_18837,N_18496);
or U19709 (N_19709,N_18814,N_18053);
or U19710 (N_19710,N_18441,N_18585);
nor U19711 (N_19711,N_18017,N_18795);
or U19712 (N_19712,N_18305,N_18352);
nand U19713 (N_19713,N_18210,N_18992);
xnor U19714 (N_19714,N_18912,N_18109);
or U19715 (N_19715,N_18017,N_18124);
or U19716 (N_19716,N_18768,N_18578);
and U19717 (N_19717,N_18110,N_18497);
or U19718 (N_19718,N_18296,N_18665);
nand U19719 (N_19719,N_18341,N_18144);
or U19720 (N_19720,N_18742,N_18771);
xor U19721 (N_19721,N_18074,N_18329);
and U19722 (N_19722,N_18247,N_18043);
and U19723 (N_19723,N_18114,N_18950);
nor U19724 (N_19724,N_18943,N_18258);
nand U19725 (N_19725,N_18893,N_18663);
xnor U19726 (N_19726,N_18107,N_18966);
and U19727 (N_19727,N_18472,N_18729);
or U19728 (N_19728,N_18801,N_18971);
nor U19729 (N_19729,N_18901,N_18830);
nor U19730 (N_19730,N_18096,N_18161);
nor U19731 (N_19731,N_18462,N_18472);
nand U19732 (N_19732,N_18649,N_18280);
xor U19733 (N_19733,N_18033,N_18224);
xnor U19734 (N_19734,N_18760,N_18594);
xnor U19735 (N_19735,N_18386,N_18069);
nor U19736 (N_19736,N_18437,N_18852);
xor U19737 (N_19737,N_18022,N_18000);
and U19738 (N_19738,N_18719,N_18744);
xnor U19739 (N_19739,N_18911,N_18156);
nand U19740 (N_19740,N_18837,N_18418);
or U19741 (N_19741,N_18345,N_18571);
nand U19742 (N_19742,N_18820,N_18683);
xnor U19743 (N_19743,N_18648,N_18025);
or U19744 (N_19744,N_18530,N_18514);
xor U19745 (N_19745,N_18438,N_18881);
and U19746 (N_19746,N_18106,N_18686);
xnor U19747 (N_19747,N_18570,N_18642);
xor U19748 (N_19748,N_18392,N_18852);
xnor U19749 (N_19749,N_18062,N_18993);
nor U19750 (N_19750,N_18357,N_18339);
or U19751 (N_19751,N_18648,N_18679);
and U19752 (N_19752,N_18649,N_18503);
nand U19753 (N_19753,N_18554,N_18516);
nor U19754 (N_19754,N_18559,N_18207);
or U19755 (N_19755,N_18449,N_18993);
nor U19756 (N_19756,N_18135,N_18890);
and U19757 (N_19757,N_18080,N_18731);
and U19758 (N_19758,N_18747,N_18873);
or U19759 (N_19759,N_18579,N_18764);
nor U19760 (N_19760,N_18022,N_18667);
xor U19761 (N_19761,N_18187,N_18445);
nor U19762 (N_19762,N_18152,N_18834);
xnor U19763 (N_19763,N_18911,N_18081);
xnor U19764 (N_19764,N_18224,N_18404);
xnor U19765 (N_19765,N_18444,N_18543);
xor U19766 (N_19766,N_18702,N_18951);
xnor U19767 (N_19767,N_18643,N_18605);
nor U19768 (N_19768,N_18925,N_18664);
or U19769 (N_19769,N_18144,N_18385);
nand U19770 (N_19770,N_18261,N_18131);
xor U19771 (N_19771,N_18345,N_18684);
nor U19772 (N_19772,N_18071,N_18511);
or U19773 (N_19773,N_18110,N_18676);
or U19774 (N_19774,N_18341,N_18009);
xor U19775 (N_19775,N_18784,N_18404);
or U19776 (N_19776,N_18872,N_18980);
nor U19777 (N_19777,N_18106,N_18822);
nor U19778 (N_19778,N_18484,N_18900);
nor U19779 (N_19779,N_18379,N_18308);
xnor U19780 (N_19780,N_18146,N_18500);
or U19781 (N_19781,N_18062,N_18309);
and U19782 (N_19782,N_18902,N_18388);
nand U19783 (N_19783,N_18790,N_18110);
and U19784 (N_19784,N_18462,N_18085);
nor U19785 (N_19785,N_18333,N_18839);
or U19786 (N_19786,N_18130,N_18628);
nand U19787 (N_19787,N_18173,N_18509);
nor U19788 (N_19788,N_18772,N_18146);
nor U19789 (N_19789,N_18057,N_18787);
xnor U19790 (N_19790,N_18239,N_18509);
xnor U19791 (N_19791,N_18310,N_18115);
or U19792 (N_19792,N_18584,N_18376);
xor U19793 (N_19793,N_18470,N_18948);
nand U19794 (N_19794,N_18560,N_18299);
xor U19795 (N_19795,N_18297,N_18987);
xnor U19796 (N_19796,N_18746,N_18675);
or U19797 (N_19797,N_18275,N_18209);
and U19798 (N_19798,N_18145,N_18616);
nand U19799 (N_19799,N_18529,N_18482);
or U19800 (N_19800,N_18236,N_18106);
or U19801 (N_19801,N_18304,N_18955);
nor U19802 (N_19802,N_18698,N_18651);
nand U19803 (N_19803,N_18865,N_18549);
xor U19804 (N_19804,N_18554,N_18903);
nand U19805 (N_19805,N_18167,N_18996);
or U19806 (N_19806,N_18506,N_18611);
xor U19807 (N_19807,N_18203,N_18007);
or U19808 (N_19808,N_18018,N_18619);
and U19809 (N_19809,N_18448,N_18870);
nand U19810 (N_19810,N_18731,N_18713);
nor U19811 (N_19811,N_18353,N_18390);
or U19812 (N_19812,N_18794,N_18844);
xnor U19813 (N_19813,N_18180,N_18649);
nand U19814 (N_19814,N_18320,N_18004);
xnor U19815 (N_19815,N_18293,N_18860);
nand U19816 (N_19816,N_18694,N_18684);
or U19817 (N_19817,N_18735,N_18495);
xor U19818 (N_19818,N_18690,N_18060);
and U19819 (N_19819,N_18764,N_18586);
xnor U19820 (N_19820,N_18003,N_18252);
nor U19821 (N_19821,N_18442,N_18387);
or U19822 (N_19822,N_18370,N_18348);
or U19823 (N_19823,N_18624,N_18310);
nand U19824 (N_19824,N_18707,N_18740);
and U19825 (N_19825,N_18033,N_18521);
or U19826 (N_19826,N_18746,N_18980);
or U19827 (N_19827,N_18869,N_18746);
or U19828 (N_19828,N_18185,N_18425);
xor U19829 (N_19829,N_18558,N_18569);
xor U19830 (N_19830,N_18196,N_18287);
nor U19831 (N_19831,N_18598,N_18941);
nor U19832 (N_19832,N_18094,N_18395);
nor U19833 (N_19833,N_18676,N_18120);
xnor U19834 (N_19834,N_18321,N_18157);
nor U19835 (N_19835,N_18188,N_18511);
nor U19836 (N_19836,N_18191,N_18370);
and U19837 (N_19837,N_18203,N_18346);
xor U19838 (N_19838,N_18788,N_18627);
nor U19839 (N_19839,N_18335,N_18829);
nor U19840 (N_19840,N_18791,N_18754);
nand U19841 (N_19841,N_18821,N_18045);
xnor U19842 (N_19842,N_18324,N_18453);
or U19843 (N_19843,N_18657,N_18318);
xnor U19844 (N_19844,N_18937,N_18409);
or U19845 (N_19845,N_18691,N_18561);
xor U19846 (N_19846,N_18163,N_18582);
xnor U19847 (N_19847,N_18820,N_18518);
and U19848 (N_19848,N_18802,N_18850);
and U19849 (N_19849,N_18700,N_18286);
nor U19850 (N_19850,N_18040,N_18881);
or U19851 (N_19851,N_18771,N_18412);
and U19852 (N_19852,N_18024,N_18678);
nand U19853 (N_19853,N_18025,N_18718);
or U19854 (N_19854,N_18682,N_18791);
and U19855 (N_19855,N_18265,N_18024);
nand U19856 (N_19856,N_18260,N_18027);
xor U19857 (N_19857,N_18794,N_18709);
nand U19858 (N_19858,N_18646,N_18438);
xor U19859 (N_19859,N_18218,N_18438);
or U19860 (N_19860,N_18699,N_18013);
and U19861 (N_19861,N_18719,N_18347);
or U19862 (N_19862,N_18924,N_18501);
xnor U19863 (N_19863,N_18012,N_18029);
nor U19864 (N_19864,N_18608,N_18664);
xnor U19865 (N_19865,N_18169,N_18931);
nand U19866 (N_19866,N_18117,N_18700);
nor U19867 (N_19867,N_18753,N_18724);
or U19868 (N_19868,N_18159,N_18123);
nor U19869 (N_19869,N_18111,N_18414);
or U19870 (N_19870,N_18616,N_18247);
nand U19871 (N_19871,N_18705,N_18462);
or U19872 (N_19872,N_18912,N_18775);
and U19873 (N_19873,N_18879,N_18745);
or U19874 (N_19874,N_18661,N_18608);
and U19875 (N_19875,N_18510,N_18630);
nand U19876 (N_19876,N_18704,N_18153);
nor U19877 (N_19877,N_18266,N_18782);
xnor U19878 (N_19878,N_18001,N_18600);
and U19879 (N_19879,N_18762,N_18667);
or U19880 (N_19880,N_18433,N_18996);
xnor U19881 (N_19881,N_18571,N_18719);
nand U19882 (N_19882,N_18316,N_18051);
or U19883 (N_19883,N_18967,N_18810);
and U19884 (N_19884,N_18694,N_18134);
xor U19885 (N_19885,N_18704,N_18833);
nor U19886 (N_19886,N_18181,N_18090);
nor U19887 (N_19887,N_18927,N_18948);
and U19888 (N_19888,N_18957,N_18288);
nand U19889 (N_19889,N_18688,N_18659);
xor U19890 (N_19890,N_18222,N_18298);
nor U19891 (N_19891,N_18643,N_18641);
xor U19892 (N_19892,N_18934,N_18517);
or U19893 (N_19893,N_18491,N_18753);
xor U19894 (N_19894,N_18654,N_18553);
xor U19895 (N_19895,N_18711,N_18597);
nand U19896 (N_19896,N_18723,N_18040);
nand U19897 (N_19897,N_18569,N_18857);
xor U19898 (N_19898,N_18009,N_18522);
nor U19899 (N_19899,N_18831,N_18692);
or U19900 (N_19900,N_18158,N_18260);
nand U19901 (N_19901,N_18167,N_18823);
xnor U19902 (N_19902,N_18523,N_18628);
nor U19903 (N_19903,N_18116,N_18108);
or U19904 (N_19904,N_18774,N_18666);
and U19905 (N_19905,N_18794,N_18920);
xnor U19906 (N_19906,N_18119,N_18670);
xor U19907 (N_19907,N_18561,N_18453);
xnor U19908 (N_19908,N_18781,N_18838);
xor U19909 (N_19909,N_18948,N_18488);
and U19910 (N_19910,N_18148,N_18533);
nand U19911 (N_19911,N_18990,N_18779);
nor U19912 (N_19912,N_18782,N_18361);
and U19913 (N_19913,N_18533,N_18052);
and U19914 (N_19914,N_18743,N_18547);
nor U19915 (N_19915,N_18701,N_18469);
or U19916 (N_19916,N_18131,N_18134);
and U19917 (N_19917,N_18652,N_18003);
or U19918 (N_19918,N_18618,N_18120);
and U19919 (N_19919,N_18494,N_18495);
xor U19920 (N_19920,N_18603,N_18852);
and U19921 (N_19921,N_18921,N_18231);
or U19922 (N_19922,N_18382,N_18573);
nand U19923 (N_19923,N_18381,N_18546);
nand U19924 (N_19924,N_18351,N_18879);
and U19925 (N_19925,N_18481,N_18099);
nand U19926 (N_19926,N_18582,N_18425);
nor U19927 (N_19927,N_18889,N_18888);
nor U19928 (N_19928,N_18042,N_18354);
nor U19929 (N_19929,N_18843,N_18932);
and U19930 (N_19930,N_18735,N_18275);
and U19931 (N_19931,N_18432,N_18762);
and U19932 (N_19932,N_18432,N_18368);
and U19933 (N_19933,N_18331,N_18070);
and U19934 (N_19934,N_18492,N_18435);
xnor U19935 (N_19935,N_18294,N_18826);
or U19936 (N_19936,N_18291,N_18305);
xnor U19937 (N_19937,N_18855,N_18545);
or U19938 (N_19938,N_18863,N_18668);
or U19939 (N_19939,N_18836,N_18419);
nand U19940 (N_19940,N_18246,N_18321);
nor U19941 (N_19941,N_18542,N_18032);
nand U19942 (N_19942,N_18385,N_18218);
nand U19943 (N_19943,N_18613,N_18519);
xor U19944 (N_19944,N_18082,N_18949);
or U19945 (N_19945,N_18287,N_18723);
nor U19946 (N_19946,N_18205,N_18437);
and U19947 (N_19947,N_18051,N_18001);
nand U19948 (N_19948,N_18895,N_18785);
or U19949 (N_19949,N_18116,N_18562);
and U19950 (N_19950,N_18560,N_18672);
or U19951 (N_19951,N_18336,N_18236);
xor U19952 (N_19952,N_18885,N_18151);
and U19953 (N_19953,N_18323,N_18843);
xor U19954 (N_19954,N_18665,N_18249);
nand U19955 (N_19955,N_18430,N_18183);
nand U19956 (N_19956,N_18900,N_18095);
nor U19957 (N_19957,N_18745,N_18203);
and U19958 (N_19958,N_18534,N_18420);
xnor U19959 (N_19959,N_18218,N_18817);
nand U19960 (N_19960,N_18232,N_18077);
xnor U19961 (N_19961,N_18821,N_18172);
or U19962 (N_19962,N_18317,N_18564);
xor U19963 (N_19963,N_18343,N_18928);
or U19964 (N_19964,N_18688,N_18121);
or U19965 (N_19965,N_18985,N_18680);
xnor U19966 (N_19966,N_18147,N_18701);
nand U19967 (N_19967,N_18017,N_18213);
nor U19968 (N_19968,N_18633,N_18902);
nor U19969 (N_19969,N_18559,N_18623);
nor U19970 (N_19970,N_18385,N_18528);
nor U19971 (N_19971,N_18252,N_18555);
and U19972 (N_19972,N_18668,N_18771);
xor U19973 (N_19973,N_18752,N_18139);
or U19974 (N_19974,N_18933,N_18342);
and U19975 (N_19975,N_18711,N_18991);
and U19976 (N_19976,N_18952,N_18321);
nor U19977 (N_19977,N_18451,N_18542);
nor U19978 (N_19978,N_18588,N_18679);
or U19979 (N_19979,N_18093,N_18477);
xnor U19980 (N_19980,N_18557,N_18040);
nand U19981 (N_19981,N_18242,N_18015);
nand U19982 (N_19982,N_18328,N_18521);
or U19983 (N_19983,N_18149,N_18384);
nor U19984 (N_19984,N_18342,N_18789);
xor U19985 (N_19985,N_18694,N_18602);
xnor U19986 (N_19986,N_18345,N_18001);
xnor U19987 (N_19987,N_18656,N_18274);
nor U19988 (N_19988,N_18662,N_18804);
or U19989 (N_19989,N_18260,N_18245);
nand U19990 (N_19990,N_18213,N_18295);
nor U19991 (N_19991,N_18145,N_18627);
nor U19992 (N_19992,N_18457,N_18139);
nand U19993 (N_19993,N_18720,N_18039);
and U19994 (N_19994,N_18409,N_18853);
and U19995 (N_19995,N_18878,N_18424);
nor U19996 (N_19996,N_18022,N_18391);
and U19997 (N_19997,N_18408,N_18304);
or U19998 (N_19998,N_18788,N_18930);
nand U19999 (N_19999,N_18871,N_18434);
and UO_0 (O_0,N_19834,N_19133);
or UO_1 (O_1,N_19424,N_19219);
nor UO_2 (O_2,N_19692,N_19950);
and UO_3 (O_3,N_19134,N_19736);
nor UO_4 (O_4,N_19232,N_19747);
or UO_5 (O_5,N_19877,N_19245);
and UO_6 (O_6,N_19029,N_19414);
or UO_7 (O_7,N_19577,N_19331);
xnor UO_8 (O_8,N_19495,N_19138);
nand UO_9 (O_9,N_19338,N_19938);
nand UO_10 (O_10,N_19843,N_19066);
nor UO_11 (O_11,N_19516,N_19943);
nand UO_12 (O_12,N_19361,N_19615);
nor UO_13 (O_13,N_19222,N_19044);
xnor UO_14 (O_14,N_19586,N_19140);
or UO_15 (O_15,N_19654,N_19201);
or UO_16 (O_16,N_19558,N_19087);
or UO_17 (O_17,N_19005,N_19343);
xnor UO_18 (O_18,N_19339,N_19885);
and UO_19 (O_19,N_19939,N_19024);
xnor UO_20 (O_20,N_19022,N_19532);
nand UO_21 (O_21,N_19537,N_19540);
or UO_22 (O_22,N_19327,N_19784);
and UO_23 (O_23,N_19047,N_19409);
or UO_24 (O_24,N_19709,N_19627);
or UO_25 (O_25,N_19124,N_19267);
and UO_26 (O_26,N_19909,N_19553);
and UO_27 (O_27,N_19274,N_19421);
xor UO_28 (O_28,N_19551,N_19153);
and UO_29 (O_29,N_19839,N_19651);
nand UO_30 (O_30,N_19836,N_19977);
nor UO_31 (O_31,N_19178,N_19999);
and UO_32 (O_32,N_19790,N_19247);
nor UO_33 (O_33,N_19521,N_19152);
nand UO_34 (O_34,N_19924,N_19063);
xnor UO_35 (O_35,N_19599,N_19486);
xor UO_36 (O_36,N_19815,N_19766);
and UO_37 (O_37,N_19082,N_19882);
nand UO_38 (O_38,N_19783,N_19927);
xor UO_39 (O_39,N_19813,N_19846);
or UO_40 (O_40,N_19502,N_19268);
nor UO_41 (O_41,N_19369,N_19099);
and UO_42 (O_42,N_19561,N_19590);
nor UO_43 (O_43,N_19919,N_19866);
or UO_44 (O_44,N_19230,N_19196);
nor UO_45 (O_45,N_19761,N_19275);
and UO_46 (O_46,N_19566,N_19605);
xnor UO_47 (O_47,N_19143,N_19818);
and UO_48 (O_48,N_19353,N_19391);
or UO_49 (O_49,N_19241,N_19979);
nand UO_50 (O_50,N_19775,N_19347);
nor UO_51 (O_51,N_19157,N_19655);
nand UO_52 (O_52,N_19904,N_19876);
nor UO_53 (O_53,N_19300,N_19425);
nand UO_54 (O_54,N_19127,N_19714);
or UO_55 (O_55,N_19811,N_19150);
xnor UO_56 (O_56,N_19541,N_19445);
or UO_57 (O_57,N_19437,N_19474);
and UO_58 (O_58,N_19442,N_19806);
or UO_59 (O_59,N_19522,N_19364);
and UO_60 (O_60,N_19996,N_19789);
nor UO_61 (O_61,N_19942,N_19740);
nor UO_62 (O_62,N_19148,N_19292);
xnor UO_63 (O_63,N_19609,N_19160);
xnor UO_64 (O_64,N_19632,N_19040);
or UO_65 (O_65,N_19955,N_19083);
nand UO_66 (O_66,N_19928,N_19895);
nand UO_67 (O_67,N_19491,N_19606);
nor UO_68 (O_68,N_19897,N_19908);
nand UO_69 (O_69,N_19929,N_19980);
and UO_70 (O_70,N_19049,N_19101);
nand UO_71 (O_71,N_19428,N_19475);
and UO_72 (O_72,N_19764,N_19753);
nor UO_73 (O_73,N_19595,N_19233);
or UO_74 (O_74,N_19849,N_19983);
or UO_75 (O_75,N_19628,N_19501);
or UO_76 (O_76,N_19518,N_19842);
nand UO_77 (O_77,N_19100,N_19989);
nor UO_78 (O_78,N_19700,N_19054);
or UO_79 (O_79,N_19611,N_19270);
xor UO_80 (O_80,N_19854,N_19337);
or UO_81 (O_81,N_19830,N_19868);
xor UO_82 (O_82,N_19010,N_19390);
or UO_83 (O_83,N_19976,N_19172);
nand UO_84 (O_84,N_19956,N_19888);
and UO_85 (O_85,N_19778,N_19450);
or UO_86 (O_86,N_19588,N_19793);
xor UO_87 (O_87,N_19372,N_19023);
nand UO_88 (O_88,N_19995,N_19525);
xnor UO_89 (O_89,N_19526,N_19720);
nor UO_90 (O_90,N_19696,N_19397);
and UO_91 (O_91,N_19462,N_19405);
or UO_92 (O_92,N_19771,N_19918);
xnor UO_93 (O_93,N_19803,N_19637);
and UO_94 (O_94,N_19021,N_19860);
and UO_95 (O_95,N_19772,N_19574);
nor UO_96 (O_96,N_19591,N_19972);
nor UO_97 (O_97,N_19017,N_19038);
nand UO_98 (O_98,N_19642,N_19310);
xnor UO_99 (O_99,N_19953,N_19587);
xnor UO_100 (O_100,N_19559,N_19964);
nand UO_101 (O_101,N_19848,N_19042);
nand UO_102 (O_102,N_19239,N_19332);
xor UO_103 (O_103,N_19886,N_19546);
or UO_104 (O_104,N_19136,N_19602);
nand UO_105 (O_105,N_19304,N_19785);
nor UO_106 (O_106,N_19795,N_19682);
or UO_107 (O_107,N_19097,N_19528);
or UO_108 (O_108,N_19028,N_19323);
xor UO_109 (O_109,N_19913,N_19780);
and UO_110 (O_110,N_19455,N_19672);
and UO_111 (O_111,N_19821,N_19648);
nand UO_112 (O_112,N_19542,N_19378);
nor UO_113 (O_113,N_19847,N_19725);
xor UO_114 (O_114,N_19175,N_19098);
or UO_115 (O_115,N_19809,N_19253);
and UO_116 (O_116,N_19858,N_19216);
nand UO_117 (O_117,N_19823,N_19721);
nand UO_118 (O_118,N_19570,N_19857);
xor UO_119 (O_119,N_19246,N_19679);
nand UO_120 (O_120,N_19717,N_19549);
xnor UO_121 (O_121,N_19156,N_19534);
and UO_122 (O_122,N_19004,N_19265);
nor UO_123 (O_123,N_19151,N_19906);
nand UO_124 (O_124,N_19604,N_19277);
xnor UO_125 (O_125,N_19724,N_19556);
nor UO_126 (O_126,N_19200,N_19204);
and UO_127 (O_127,N_19598,N_19110);
xnor UO_128 (O_128,N_19058,N_19808);
xor UO_129 (O_129,N_19872,N_19184);
nor UO_130 (O_130,N_19238,N_19743);
and UO_131 (O_131,N_19722,N_19217);
xnor UO_132 (O_132,N_19986,N_19105);
xor UO_133 (O_133,N_19734,N_19739);
nand UO_134 (O_134,N_19478,N_19535);
or UO_135 (O_135,N_19427,N_19601);
or UO_136 (O_136,N_19731,N_19746);
nor UO_137 (O_137,N_19658,N_19266);
and UO_138 (O_138,N_19170,N_19176);
or UO_139 (O_139,N_19417,N_19861);
nor UO_140 (O_140,N_19394,N_19431);
nor UO_141 (O_141,N_19827,N_19687);
or UO_142 (O_142,N_19992,N_19710);
xnor UO_143 (O_143,N_19420,N_19207);
nand UO_144 (O_144,N_19562,N_19223);
or UO_145 (O_145,N_19645,N_19481);
nand UO_146 (O_146,N_19752,N_19915);
nor UO_147 (O_147,N_19161,N_19096);
or UO_148 (O_148,N_19062,N_19723);
nor UO_149 (O_149,N_19027,N_19893);
nor UO_150 (O_150,N_19891,N_19622);
nand UO_151 (O_151,N_19666,N_19695);
nor UO_152 (O_152,N_19814,N_19254);
nor UO_153 (O_153,N_19545,N_19833);
or UO_154 (O_154,N_19012,N_19822);
or UO_155 (O_155,N_19874,N_19359);
xor UO_156 (O_156,N_19756,N_19884);
or UO_157 (O_157,N_19197,N_19335);
nand UO_158 (O_158,N_19608,N_19046);
nand UO_159 (O_159,N_19837,N_19146);
or UO_160 (O_160,N_19869,N_19325);
nor UO_161 (O_161,N_19064,N_19459);
nor UO_162 (O_162,N_19053,N_19504);
or UO_163 (O_163,N_19195,N_19289);
nor UO_164 (O_164,N_19086,N_19061);
or UO_165 (O_165,N_19212,N_19807);
xor UO_166 (O_166,N_19059,N_19631);
xor UO_167 (O_167,N_19191,N_19826);
nor UO_168 (O_168,N_19707,N_19515);
xnor UO_169 (O_169,N_19978,N_19494);
nand UO_170 (O_170,N_19520,N_19926);
nor UO_171 (O_171,N_19467,N_19930);
and UO_172 (O_172,N_19531,N_19711);
xor UO_173 (O_173,N_19003,N_19998);
xor UO_174 (O_174,N_19295,N_19352);
nand UO_175 (O_175,N_19900,N_19228);
nor UO_176 (O_176,N_19850,N_19031);
nand UO_177 (O_177,N_19356,N_19294);
nor UO_178 (O_178,N_19384,N_19430);
xnor UO_179 (O_179,N_19312,N_19748);
or UO_180 (O_180,N_19460,N_19508);
nor UO_181 (O_181,N_19342,N_19358);
xnor UO_182 (O_182,N_19712,N_19859);
xor UO_183 (O_183,N_19825,N_19831);
nor UO_184 (O_184,N_19092,N_19792);
nor UO_185 (O_185,N_19050,N_19411);
or UO_186 (O_186,N_19400,N_19444);
or UO_187 (O_187,N_19963,N_19781);
xnor UO_188 (O_188,N_19940,N_19701);
and UO_189 (O_189,N_19936,N_19804);
xor UO_190 (O_190,N_19603,N_19765);
or UO_191 (O_191,N_19910,N_19290);
nor UO_192 (O_192,N_19280,N_19681);
and UO_193 (O_193,N_19041,N_19640);
nand UO_194 (O_194,N_19382,N_19068);
nand UO_195 (O_195,N_19530,N_19434);
and UO_196 (O_196,N_19203,N_19669);
xor UO_197 (O_197,N_19510,N_19788);
xnor UO_198 (O_198,N_19987,N_19131);
and UO_199 (O_199,N_19320,N_19423);
or UO_200 (O_200,N_19738,N_19167);
nand UO_201 (O_201,N_19935,N_19705);
or UO_202 (O_202,N_19240,N_19898);
nor UO_203 (O_203,N_19311,N_19519);
and UO_204 (O_204,N_19536,N_19177);
nand UO_205 (O_205,N_19630,N_19768);
xor UO_206 (O_206,N_19621,N_19291);
nand UO_207 (O_207,N_19664,N_19000);
xnor UO_208 (O_208,N_19864,N_19227);
xnor UO_209 (O_209,N_19899,N_19596);
nand UO_210 (O_210,N_19773,N_19344);
nand UO_211 (O_211,N_19413,N_19180);
or UO_212 (O_212,N_19547,N_19517);
nand UO_213 (O_213,N_19305,N_19279);
xnor UO_214 (O_214,N_19506,N_19635);
or UO_215 (O_215,N_19284,N_19081);
and UO_216 (O_216,N_19346,N_19639);
or UO_217 (O_217,N_19137,N_19912);
nor UO_218 (O_218,N_19688,N_19169);
nand UO_219 (O_219,N_19727,N_19851);
and UO_220 (O_220,N_19438,N_19048);
xnor UO_221 (O_221,N_19514,N_19164);
nand UO_222 (O_222,N_19366,N_19398);
nand UO_223 (O_223,N_19213,N_19067);
nor UO_224 (O_224,N_19115,N_19961);
xnor UO_225 (O_225,N_19319,N_19190);
xor UO_226 (O_226,N_19260,N_19569);
or UO_227 (O_227,N_19816,N_19435);
xnor UO_228 (O_228,N_19759,N_19647);
nor UO_229 (O_229,N_19488,N_19659);
or UO_230 (O_230,N_19817,N_19917);
nand UO_231 (O_231,N_19464,N_19057);
xnor UO_232 (O_232,N_19243,N_19341);
and UO_233 (O_233,N_19447,N_19933);
xnor UO_234 (O_234,N_19149,N_19675);
nor UO_235 (O_235,N_19957,N_19568);
and UO_236 (O_236,N_19656,N_19357);
or UO_237 (O_237,N_19244,N_19796);
and UO_238 (O_238,N_19465,N_19168);
nand UO_239 (O_239,N_19463,N_19163);
nand UO_240 (O_240,N_19523,N_19729);
and UO_241 (O_241,N_19077,N_19008);
nor UO_242 (O_242,N_19030,N_19155);
and UO_243 (O_243,N_19680,N_19433);
nor UO_244 (O_244,N_19819,N_19745);
or UO_245 (O_245,N_19316,N_19457);
nor UO_246 (O_246,N_19626,N_19485);
and UO_247 (O_247,N_19043,N_19799);
xor UO_248 (O_248,N_19315,N_19862);
or UO_249 (O_249,N_19403,N_19879);
xor UO_250 (O_250,N_19194,N_19482);
nor UO_251 (O_251,N_19234,N_19966);
and UO_252 (O_252,N_19890,N_19144);
or UO_253 (O_253,N_19828,N_19511);
nand UO_254 (O_254,N_19370,N_19374);
xor UO_255 (O_255,N_19563,N_19162);
and UO_256 (O_256,N_19074,N_19544);
and UO_257 (O_257,N_19399,N_19301);
or UO_258 (O_258,N_19782,N_19840);
xnor UO_259 (O_259,N_19363,N_19173);
xnor UO_260 (O_260,N_19770,N_19103);
xnor UO_261 (O_261,N_19767,N_19691);
nand UO_262 (O_262,N_19250,N_19334);
nand UO_263 (O_263,N_19261,N_19011);
or UO_264 (O_264,N_19597,N_19797);
nand UO_265 (O_265,N_19122,N_19065);
nand UO_266 (O_266,N_19051,N_19135);
nor UO_267 (O_267,N_19503,N_19443);
nand UO_268 (O_268,N_19154,N_19252);
nand UO_269 (O_269,N_19584,N_19844);
or UO_270 (O_270,N_19496,N_19901);
and UO_271 (O_271,N_19873,N_19629);
or UO_272 (O_272,N_19962,N_19922);
and UO_273 (O_273,N_19618,N_19794);
nand UO_274 (O_274,N_19355,N_19832);
nor UO_275 (O_275,N_19580,N_19557);
xor UO_276 (O_276,N_19385,N_19288);
nor UO_277 (O_277,N_19193,N_19007);
xnor UO_278 (O_278,N_19393,N_19845);
xor UO_279 (O_279,N_19726,N_19129);
xnor UO_280 (O_280,N_19902,N_19209);
nand UO_281 (O_281,N_19299,N_19104);
or UO_282 (O_282,N_19205,N_19644);
nor UO_283 (O_283,N_19056,N_19760);
xor UO_284 (O_284,N_19708,N_19662);
xnor UO_285 (O_285,N_19026,N_19538);
nor UO_286 (O_286,N_19365,N_19881);
nand UO_287 (O_287,N_19446,N_19954);
or UO_288 (O_288,N_19617,N_19490);
xor UO_289 (O_289,N_19937,N_19282);
nor UO_290 (O_290,N_19932,N_19013);
nor UO_291 (O_291,N_19255,N_19718);
or UO_292 (O_292,N_19896,N_19777);
or UO_293 (O_293,N_19202,N_19527);
nor UO_294 (O_294,N_19550,N_19111);
or UO_295 (O_295,N_19235,N_19470);
xor UO_296 (O_296,N_19641,N_19947);
nand UO_297 (O_297,N_19293,N_19671);
nor UO_298 (O_298,N_19841,N_19383);
nand UO_299 (O_299,N_19226,N_19719);
and UO_300 (O_300,N_19322,N_19883);
and UO_301 (O_301,N_19123,N_19774);
nor UO_302 (O_302,N_19451,N_19985);
and UO_303 (O_303,N_19565,N_19091);
and UO_304 (O_304,N_19045,N_19313);
nor UO_305 (O_305,N_19875,N_19916);
nand UO_306 (O_306,N_19674,N_19218);
nand UO_307 (O_307,N_19458,N_19019);
xor UO_308 (O_308,N_19991,N_19307);
xor UO_309 (O_309,N_19117,N_19221);
nor UO_310 (O_310,N_19529,N_19921);
and UO_311 (O_311,N_19368,N_19614);
nand UO_312 (O_312,N_19259,N_19824);
nor UO_313 (O_313,N_19468,N_19564);
xor UO_314 (O_314,N_19441,N_19340);
nor UO_315 (O_315,N_19829,N_19970);
and UO_316 (O_316,N_19499,N_19646);
xor UO_317 (O_317,N_19380,N_19006);
and UO_318 (O_318,N_19974,N_19329);
xnor UO_319 (O_319,N_19256,N_19089);
nor UO_320 (O_320,N_19702,N_19052);
nand UO_321 (O_321,N_19419,N_19107);
and UO_322 (O_322,N_19395,N_19592);
and UO_323 (O_323,N_19032,N_19185);
xor UO_324 (O_324,N_19142,N_19229);
and UO_325 (O_325,N_19037,N_19552);
nand UO_326 (O_326,N_19479,N_19249);
or UO_327 (O_327,N_19112,N_19035);
and UO_328 (O_328,N_19704,N_19432);
xnor UO_329 (O_329,N_19483,N_19020);
xor UO_330 (O_330,N_19406,N_19934);
or UO_331 (O_331,N_19732,N_19330);
nand UO_332 (O_332,N_19415,N_19166);
nand UO_333 (O_333,N_19619,N_19471);
xor UO_334 (O_334,N_19994,N_19225);
nand UO_335 (O_335,N_19779,N_19524);
nor UO_336 (O_336,N_19199,N_19607);
nor UO_337 (O_337,N_19461,N_19348);
or UO_338 (O_338,N_19500,N_19578);
nand UO_339 (O_339,N_19871,N_19533);
nand UO_340 (O_340,N_19625,N_19147);
nor UO_341 (O_341,N_19762,N_19440);
nand UO_342 (O_342,N_19750,N_19703);
and UO_343 (O_343,N_19095,N_19685);
or UO_344 (O_344,N_19683,N_19220);
and UO_345 (O_345,N_19237,N_19663);
nor UO_346 (O_346,N_19981,N_19251);
nand UO_347 (O_347,N_19993,N_19211);
nor UO_348 (O_348,N_19351,N_19298);
and UO_349 (O_349,N_19278,N_19755);
and UO_350 (O_350,N_19080,N_19242);
nor UO_351 (O_351,N_19386,N_19758);
or UO_352 (O_352,N_19125,N_19333);
nor UO_353 (O_353,N_19119,N_19798);
xnor UO_354 (O_354,N_19033,N_19911);
and UO_355 (O_355,N_19667,N_19810);
or UO_356 (O_356,N_19623,N_19668);
xnor UO_357 (O_357,N_19009,N_19812);
or UO_358 (O_358,N_19257,N_19971);
xor UO_359 (O_359,N_19426,N_19113);
or UO_360 (O_360,N_19215,N_19960);
nand UO_361 (O_361,N_19984,N_19802);
nor UO_362 (O_362,N_19371,N_19036);
nand UO_363 (O_363,N_19643,N_19145);
and UO_364 (O_364,N_19948,N_19543);
or UO_365 (O_365,N_19636,N_19555);
and UO_366 (O_366,N_19324,N_19865);
or UO_367 (O_367,N_19585,N_19130);
nand UO_368 (O_368,N_19132,N_19676);
and UO_369 (O_369,N_19477,N_19071);
nor UO_370 (O_370,N_19072,N_19579);
and UO_371 (O_371,N_19408,N_19497);
nor UO_372 (O_372,N_19165,N_19039);
nand UO_373 (O_373,N_19326,N_19069);
and UO_374 (O_374,N_19716,N_19094);
or UO_375 (O_375,N_19264,N_19946);
nor UO_376 (O_376,N_19018,N_19554);
or UO_377 (O_377,N_19573,N_19404);
nor UO_378 (O_378,N_19863,N_19141);
xnor UO_379 (O_379,N_19713,N_19944);
xnor UO_380 (O_380,N_19387,N_19480);
nor UO_381 (O_381,N_19016,N_19751);
nor UO_382 (O_382,N_19410,N_19835);
or UO_383 (O_383,N_19572,N_19453);
nand UO_384 (O_384,N_19236,N_19073);
or UO_385 (O_385,N_19730,N_19263);
nor UO_386 (O_386,N_19345,N_19763);
or UO_387 (O_387,N_19997,N_19093);
nor UO_388 (O_388,N_19694,N_19078);
xnor UO_389 (O_389,N_19801,N_19187);
or UO_390 (O_390,N_19192,N_19594);
or UO_391 (O_391,N_19975,N_19466);
nand UO_392 (O_392,N_19174,N_19698);
nor UO_393 (O_393,N_19297,N_19287);
nor UO_394 (O_394,N_19476,N_19181);
nor UO_395 (O_395,N_19484,N_19412);
nand UO_396 (O_396,N_19638,N_19076);
and UO_397 (O_397,N_19706,N_19905);
nor UO_398 (O_398,N_19283,N_19958);
nor UO_399 (O_399,N_19684,N_19689);
nor UO_400 (O_400,N_19354,N_19120);
or UO_401 (O_401,N_19616,N_19969);
nand UO_402 (O_402,N_19452,N_19951);
xor UO_403 (O_403,N_19742,N_19472);
nor UO_404 (O_404,N_19448,N_19401);
nand UO_405 (O_405,N_19248,N_19931);
and UO_406 (O_406,N_19690,N_19853);
and UO_407 (O_407,N_19769,N_19660);
or UO_408 (O_408,N_19657,N_19610);
and UO_409 (O_409,N_19593,N_19649);
xor UO_410 (O_410,N_19894,N_19581);
and UO_411 (O_411,N_19273,N_19262);
or UO_412 (O_412,N_19673,N_19612);
and UO_413 (O_413,N_19852,N_19118);
nand UO_414 (O_414,N_19303,N_19487);
nor UO_415 (O_415,N_19941,N_19973);
nand UO_416 (O_416,N_19686,N_19376);
xnor UO_417 (O_417,N_19949,N_19429);
or UO_418 (O_418,N_19988,N_19085);
or UO_419 (O_419,N_19381,N_19377);
xor UO_420 (O_420,N_19188,N_19002);
xnor UO_421 (O_421,N_19678,N_19805);
and UO_422 (O_422,N_19820,N_19108);
and UO_423 (O_423,N_19634,N_19735);
nor UO_424 (O_424,N_19737,N_19088);
nand UO_425 (O_425,N_19661,N_19548);
or UO_426 (O_426,N_19126,N_19281);
and UO_427 (O_427,N_19296,N_19128);
or UO_428 (O_428,N_19416,N_19318);
xor UO_429 (O_429,N_19867,N_19513);
and UO_430 (O_430,N_19576,N_19286);
and UO_431 (O_431,N_19582,N_19920);
and UO_432 (O_432,N_19379,N_19328);
xor UO_433 (O_433,N_19952,N_19733);
nor UO_434 (O_434,N_19418,N_19914);
or UO_435 (O_435,N_19362,N_19102);
nand UO_436 (O_436,N_19258,N_19889);
or UO_437 (O_437,N_19741,N_19109);
or UO_438 (O_438,N_19407,N_19982);
or UO_439 (O_439,N_19907,N_19367);
nand UO_440 (O_440,N_19389,N_19454);
nand UO_441 (O_441,N_19090,N_19171);
or UO_442 (O_442,N_19186,N_19498);
xnor UO_443 (O_443,N_19493,N_19880);
and UO_444 (O_444,N_19276,N_19210);
xor UO_445 (O_445,N_19034,N_19079);
and UO_446 (O_446,N_19179,N_19600);
xnor UO_447 (O_447,N_19001,N_19015);
and UO_448 (O_448,N_19624,N_19728);
nor UO_449 (O_449,N_19159,N_19925);
nor UO_450 (O_450,N_19571,N_19903);
and UO_451 (O_451,N_19633,N_19014);
or UO_452 (O_452,N_19892,N_19776);
or UO_453 (O_453,N_19422,N_19838);
xor UO_454 (O_454,N_19613,N_19650);
nor UO_455 (O_455,N_19449,N_19314);
xnor UO_456 (O_456,N_19959,N_19182);
and UO_457 (O_457,N_19436,N_19306);
xnor UO_458 (O_458,N_19787,N_19302);
or UO_459 (O_459,N_19208,N_19388);
and UO_460 (O_460,N_19583,N_19317);
and UO_461 (O_461,N_19653,N_19715);
nor UO_462 (O_462,N_19060,N_19693);
and UO_463 (O_463,N_19749,N_19575);
or UO_464 (O_464,N_19652,N_19589);
and UO_465 (O_465,N_19923,N_19375);
and UO_466 (O_466,N_19670,N_19965);
nor UO_467 (O_467,N_19189,N_19336);
nor UO_468 (O_468,N_19665,N_19373);
nor UO_469 (O_469,N_19198,N_19855);
and UO_470 (O_470,N_19084,N_19114);
xor UO_471 (O_471,N_19439,N_19183);
or UO_472 (O_472,N_19505,N_19214);
and UO_473 (O_473,N_19512,N_19757);
nor UO_474 (O_474,N_19106,N_19744);
and UO_475 (O_475,N_19139,N_19677);
and UO_476 (O_476,N_19070,N_19360);
nor UO_477 (O_477,N_19887,N_19224);
xor UO_478 (O_478,N_19116,N_19990);
and UO_479 (O_479,N_19560,N_19870);
nand UO_480 (O_480,N_19945,N_19856);
or UO_481 (O_481,N_19699,N_19507);
or UO_482 (O_482,N_19055,N_19269);
nand UO_483 (O_483,N_19396,N_19509);
or UO_484 (O_484,N_19308,N_19349);
xnor UO_485 (O_485,N_19968,N_19272);
xnor UO_486 (O_486,N_19321,N_19800);
nor UO_487 (O_487,N_19878,N_19456);
xor UO_488 (O_488,N_19285,N_19489);
nor UO_489 (O_489,N_19158,N_19350);
and UO_490 (O_490,N_19469,N_19567);
and UO_491 (O_491,N_19492,N_19539);
nand UO_492 (O_492,N_19754,N_19271);
xor UO_493 (O_493,N_19791,N_19121);
or UO_494 (O_494,N_19206,N_19402);
and UO_495 (O_495,N_19967,N_19025);
xor UO_496 (O_496,N_19620,N_19309);
nand UO_497 (O_497,N_19392,N_19473);
nor UO_498 (O_498,N_19786,N_19697);
nand UO_499 (O_499,N_19231,N_19075);
nor UO_500 (O_500,N_19218,N_19575);
nor UO_501 (O_501,N_19216,N_19815);
and UO_502 (O_502,N_19602,N_19827);
and UO_503 (O_503,N_19501,N_19927);
or UO_504 (O_504,N_19270,N_19900);
or UO_505 (O_505,N_19814,N_19782);
and UO_506 (O_506,N_19068,N_19865);
or UO_507 (O_507,N_19084,N_19854);
or UO_508 (O_508,N_19635,N_19926);
xor UO_509 (O_509,N_19790,N_19258);
nor UO_510 (O_510,N_19626,N_19211);
and UO_511 (O_511,N_19801,N_19899);
or UO_512 (O_512,N_19942,N_19620);
nor UO_513 (O_513,N_19474,N_19750);
or UO_514 (O_514,N_19496,N_19914);
nand UO_515 (O_515,N_19270,N_19136);
nand UO_516 (O_516,N_19328,N_19770);
xnor UO_517 (O_517,N_19590,N_19762);
and UO_518 (O_518,N_19919,N_19258);
and UO_519 (O_519,N_19976,N_19767);
or UO_520 (O_520,N_19485,N_19975);
or UO_521 (O_521,N_19090,N_19878);
or UO_522 (O_522,N_19083,N_19754);
nor UO_523 (O_523,N_19129,N_19592);
nor UO_524 (O_524,N_19914,N_19145);
or UO_525 (O_525,N_19887,N_19277);
or UO_526 (O_526,N_19105,N_19055);
or UO_527 (O_527,N_19506,N_19156);
nand UO_528 (O_528,N_19459,N_19047);
and UO_529 (O_529,N_19985,N_19355);
nor UO_530 (O_530,N_19194,N_19854);
nor UO_531 (O_531,N_19399,N_19738);
nor UO_532 (O_532,N_19544,N_19331);
xnor UO_533 (O_533,N_19088,N_19820);
and UO_534 (O_534,N_19815,N_19721);
or UO_535 (O_535,N_19501,N_19281);
xnor UO_536 (O_536,N_19799,N_19059);
and UO_537 (O_537,N_19530,N_19674);
or UO_538 (O_538,N_19817,N_19313);
or UO_539 (O_539,N_19584,N_19085);
or UO_540 (O_540,N_19986,N_19229);
nand UO_541 (O_541,N_19925,N_19061);
xnor UO_542 (O_542,N_19217,N_19145);
nand UO_543 (O_543,N_19692,N_19467);
nor UO_544 (O_544,N_19529,N_19415);
or UO_545 (O_545,N_19280,N_19079);
xnor UO_546 (O_546,N_19211,N_19046);
or UO_547 (O_547,N_19547,N_19599);
nor UO_548 (O_548,N_19909,N_19609);
or UO_549 (O_549,N_19671,N_19689);
xnor UO_550 (O_550,N_19191,N_19326);
xor UO_551 (O_551,N_19183,N_19597);
nand UO_552 (O_552,N_19500,N_19524);
nand UO_553 (O_553,N_19564,N_19693);
nand UO_554 (O_554,N_19236,N_19994);
xor UO_555 (O_555,N_19701,N_19401);
nand UO_556 (O_556,N_19595,N_19454);
xnor UO_557 (O_557,N_19452,N_19366);
xor UO_558 (O_558,N_19197,N_19529);
xnor UO_559 (O_559,N_19477,N_19228);
and UO_560 (O_560,N_19638,N_19513);
or UO_561 (O_561,N_19035,N_19585);
and UO_562 (O_562,N_19104,N_19682);
nor UO_563 (O_563,N_19685,N_19828);
nor UO_564 (O_564,N_19141,N_19487);
xor UO_565 (O_565,N_19326,N_19849);
xnor UO_566 (O_566,N_19666,N_19797);
and UO_567 (O_567,N_19078,N_19901);
xnor UO_568 (O_568,N_19335,N_19326);
nor UO_569 (O_569,N_19645,N_19851);
and UO_570 (O_570,N_19758,N_19622);
and UO_571 (O_571,N_19698,N_19984);
xnor UO_572 (O_572,N_19883,N_19020);
or UO_573 (O_573,N_19780,N_19960);
xor UO_574 (O_574,N_19818,N_19188);
nand UO_575 (O_575,N_19020,N_19389);
or UO_576 (O_576,N_19028,N_19178);
or UO_577 (O_577,N_19303,N_19890);
and UO_578 (O_578,N_19872,N_19902);
nor UO_579 (O_579,N_19591,N_19687);
xor UO_580 (O_580,N_19110,N_19263);
xnor UO_581 (O_581,N_19029,N_19827);
xnor UO_582 (O_582,N_19151,N_19753);
and UO_583 (O_583,N_19886,N_19223);
or UO_584 (O_584,N_19117,N_19980);
and UO_585 (O_585,N_19766,N_19667);
nand UO_586 (O_586,N_19818,N_19042);
nor UO_587 (O_587,N_19101,N_19201);
nor UO_588 (O_588,N_19925,N_19132);
nand UO_589 (O_589,N_19823,N_19615);
and UO_590 (O_590,N_19854,N_19513);
nor UO_591 (O_591,N_19806,N_19579);
nor UO_592 (O_592,N_19456,N_19177);
nand UO_593 (O_593,N_19607,N_19525);
and UO_594 (O_594,N_19874,N_19234);
and UO_595 (O_595,N_19679,N_19981);
xnor UO_596 (O_596,N_19633,N_19048);
xor UO_597 (O_597,N_19142,N_19175);
or UO_598 (O_598,N_19291,N_19695);
or UO_599 (O_599,N_19427,N_19209);
xnor UO_600 (O_600,N_19690,N_19056);
nor UO_601 (O_601,N_19577,N_19976);
and UO_602 (O_602,N_19330,N_19578);
nor UO_603 (O_603,N_19419,N_19558);
nor UO_604 (O_604,N_19234,N_19242);
nor UO_605 (O_605,N_19493,N_19590);
nand UO_606 (O_606,N_19174,N_19259);
or UO_607 (O_607,N_19701,N_19680);
nor UO_608 (O_608,N_19608,N_19810);
nor UO_609 (O_609,N_19294,N_19012);
nand UO_610 (O_610,N_19846,N_19166);
nand UO_611 (O_611,N_19433,N_19388);
nand UO_612 (O_612,N_19058,N_19020);
and UO_613 (O_613,N_19438,N_19945);
and UO_614 (O_614,N_19726,N_19579);
or UO_615 (O_615,N_19797,N_19997);
xnor UO_616 (O_616,N_19128,N_19492);
or UO_617 (O_617,N_19279,N_19532);
and UO_618 (O_618,N_19164,N_19033);
xnor UO_619 (O_619,N_19857,N_19831);
or UO_620 (O_620,N_19209,N_19199);
nor UO_621 (O_621,N_19934,N_19151);
nand UO_622 (O_622,N_19932,N_19034);
nor UO_623 (O_623,N_19323,N_19265);
and UO_624 (O_624,N_19427,N_19978);
nand UO_625 (O_625,N_19409,N_19993);
and UO_626 (O_626,N_19318,N_19813);
or UO_627 (O_627,N_19236,N_19116);
xor UO_628 (O_628,N_19667,N_19741);
and UO_629 (O_629,N_19239,N_19147);
xnor UO_630 (O_630,N_19580,N_19573);
xor UO_631 (O_631,N_19883,N_19807);
xor UO_632 (O_632,N_19329,N_19633);
or UO_633 (O_633,N_19798,N_19141);
nand UO_634 (O_634,N_19607,N_19618);
xor UO_635 (O_635,N_19598,N_19045);
or UO_636 (O_636,N_19675,N_19220);
nor UO_637 (O_637,N_19782,N_19100);
and UO_638 (O_638,N_19933,N_19824);
nor UO_639 (O_639,N_19802,N_19025);
and UO_640 (O_640,N_19610,N_19120);
nand UO_641 (O_641,N_19397,N_19580);
nor UO_642 (O_642,N_19776,N_19167);
or UO_643 (O_643,N_19071,N_19846);
nor UO_644 (O_644,N_19194,N_19195);
nor UO_645 (O_645,N_19547,N_19780);
nand UO_646 (O_646,N_19954,N_19576);
and UO_647 (O_647,N_19336,N_19618);
and UO_648 (O_648,N_19604,N_19352);
nand UO_649 (O_649,N_19007,N_19577);
xor UO_650 (O_650,N_19241,N_19136);
and UO_651 (O_651,N_19871,N_19205);
and UO_652 (O_652,N_19761,N_19063);
xor UO_653 (O_653,N_19098,N_19847);
xnor UO_654 (O_654,N_19129,N_19529);
and UO_655 (O_655,N_19431,N_19311);
nand UO_656 (O_656,N_19765,N_19311);
nor UO_657 (O_657,N_19927,N_19017);
nor UO_658 (O_658,N_19220,N_19805);
nand UO_659 (O_659,N_19443,N_19804);
or UO_660 (O_660,N_19462,N_19861);
xor UO_661 (O_661,N_19577,N_19440);
or UO_662 (O_662,N_19473,N_19070);
nor UO_663 (O_663,N_19598,N_19530);
nand UO_664 (O_664,N_19265,N_19613);
nor UO_665 (O_665,N_19071,N_19448);
xnor UO_666 (O_666,N_19753,N_19236);
xor UO_667 (O_667,N_19659,N_19970);
and UO_668 (O_668,N_19815,N_19715);
xor UO_669 (O_669,N_19699,N_19878);
xor UO_670 (O_670,N_19458,N_19596);
nand UO_671 (O_671,N_19694,N_19045);
xnor UO_672 (O_672,N_19149,N_19478);
and UO_673 (O_673,N_19082,N_19068);
or UO_674 (O_674,N_19935,N_19936);
xnor UO_675 (O_675,N_19357,N_19705);
and UO_676 (O_676,N_19933,N_19912);
nor UO_677 (O_677,N_19779,N_19713);
and UO_678 (O_678,N_19581,N_19877);
nor UO_679 (O_679,N_19951,N_19208);
or UO_680 (O_680,N_19761,N_19752);
nor UO_681 (O_681,N_19951,N_19598);
and UO_682 (O_682,N_19859,N_19203);
or UO_683 (O_683,N_19192,N_19137);
xor UO_684 (O_684,N_19423,N_19430);
nor UO_685 (O_685,N_19964,N_19102);
xnor UO_686 (O_686,N_19181,N_19693);
and UO_687 (O_687,N_19744,N_19392);
nor UO_688 (O_688,N_19278,N_19118);
xor UO_689 (O_689,N_19065,N_19012);
or UO_690 (O_690,N_19465,N_19339);
and UO_691 (O_691,N_19423,N_19080);
xnor UO_692 (O_692,N_19166,N_19621);
nand UO_693 (O_693,N_19435,N_19748);
xor UO_694 (O_694,N_19993,N_19471);
nand UO_695 (O_695,N_19949,N_19102);
nand UO_696 (O_696,N_19476,N_19705);
or UO_697 (O_697,N_19602,N_19736);
xor UO_698 (O_698,N_19752,N_19083);
nand UO_699 (O_699,N_19882,N_19583);
or UO_700 (O_700,N_19544,N_19045);
and UO_701 (O_701,N_19392,N_19299);
and UO_702 (O_702,N_19398,N_19040);
xor UO_703 (O_703,N_19564,N_19645);
or UO_704 (O_704,N_19796,N_19038);
and UO_705 (O_705,N_19315,N_19219);
or UO_706 (O_706,N_19706,N_19710);
nor UO_707 (O_707,N_19545,N_19937);
nor UO_708 (O_708,N_19469,N_19962);
and UO_709 (O_709,N_19428,N_19650);
or UO_710 (O_710,N_19594,N_19643);
and UO_711 (O_711,N_19426,N_19475);
nand UO_712 (O_712,N_19696,N_19032);
or UO_713 (O_713,N_19374,N_19467);
and UO_714 (O_714,N_19816,N_19671);
and UO_715 (O_715,N_19139,N_19063);
and UO_716 (O_716,N_19665,N_19077);
or UO_717 (O_717,N_19965,N_19630);
nand UO_718 (O_718,N_19629,N_19388);
nand UO_719 (O_719,N_19008,N_19795);
xor UO_720 (O_720,N_19523,N_19077);
or UO_721 (O_721,N_19496,N_19053);
nand UO_722 (O_722,N_19830,N_19488);
xor UO_723 (O_723,N_19534,N_19678);
nand UO_724 (O_724,N_19213,N_19524);
and UO_725 (O_725,N_19292,N_19166);
xor UO_726 (O_726,N_19572,N_19694);
xnor UO_727 (O_727,N_19084,N_19530);
nor UO_728 (O_728,N_19237,N_19460);
nand UO_729 (O_729,N_19476,N_19112);
xor UO_730 (O_730,N_19146,N_19486);
xnor UO_731 (O_731,N_19693,N_19989);
xor UO_732 (O_732,N_19464,N_19888);
or UO_733 (O_733,N_19632,N_19548);
xor UO_734 (O_734,N_19954,N_19115);
and UO_735 (O_735,N_19686,N_19466);
and UO_736 (O_736,N_19277,N_19850);
and UO_737 (O_737,N_19444,N_19758);
and UO_738 (O_738,N_19430,N_19029);
xor UO_739 (O_739,N_19685,N_19714);
and UO_740 (O_740,N_19396,N_19680);
nand UO_741 (O_741,N_19525,N_19769);
or UO_742 (O_742,N_19444,N_19943);
xor UO_743 (O_743,N_19173,N_19343);
or UO_744 (O_744,N_19730,N_19662);
nand UO_745 (O_745,N_19578,N_19535);
nor UO_746 (O_746,N_19013,N_19743);
xnor UO_747 (O_747,N_19967,N_19112);
xnor UO_748 (O_748,N_19406,N_19842);
and UO_749 (O_749,N_19654,N_19623);
or UO_750 (O_750,N_19303,N_19720);
nor UO_751 (O_751,N_19450,N_19744);
nor UO_752 (O_752,N_19785,N_19673);
and UO_753 (O_753,N_19263,N_19184);
or UO_754 (O_754,N_19034,N_19737);
xor UO_755 (O_755,N_19690,N_19052);
nor UO_756 (O_756,N_19135,N_19780);
and UO_757 (O_757,N_19527,N_19561);
or UO_758 (O_758,N_19588,N_19872);
or UO_759 (O_759,N_19160,N_19177);
xnor UO_760 (O_760,N_19630,N_19862);
nor UO_761 (O_761,N_19042,N_19762);
nand UO_762 (O_762,N_19609,N_19137);
and UO_763 (O_763,N_19574,N_19646);
nor UO_764 (O_764,N_19553,N_19648);
xor UO_765 (O_765,N_19499,N_19239);
or UO_766 (O_766,N_19930,N_19704);
and UO_767 (O_767,N_19365,N_19354);
nand UO_768 (O_768,N_19029,N_19785);
nor UO_769 (O_769,N_19864,N_19792);
and UO_770 (O_770,N_19013,N_19320);
or UO_771 (O_771,N_19794,N_19029);
or UO_772 (O_772,N_19038,N_19496);
xor UO_773 (O_773,N_19977,N_19512);
nand UO_774 (O_774,N_19601,N_19207);
nand UO_775 (O_775,N_19568,N_19404);
xor UO_776 (O_776,N_19109,N_19512);
and UO_777 (O_777,N_19324,N_19185);
xor UO_778 (O_778,N_19387,N_19691);
nor UO_779 (O_779,N_19972,N_19738);
xnor UO_780 (O_780,N_19054,N_19193);
or UO_781 (O_781,N_19471,N_19378);
nor UO_782 (O_782,N_19788,N_19085);
xnor UO_783 (O_783,N_19447,N_19496);
and UO_784 (O_784,N_19510,N_19573);
nor UO_785 (O_785,N_19756,N_19470);
and UO_786 (O_786,N_19100,N_19317);
nor UO_787 (O_787,N_19890,N_19559);
xor UO_788 (O_788,N_19689,N_19233);
nand UO_789 (O_789,N_19208,N_19719);
xor UO_790 (O_790,N_19644,N_19523);
or UO_791 (O_791,N_19269,N_19864);
or UO_792 (O_792,N_19421,N_19972);
nand UO_793 (O_793,N_19927,N_19306);
nor UO_794 (O_794,N_19385,N_19560);
nand UO_795 (O_795,N_19997,N_19240);
nor UO_796 (O_796,N_19059,N_19774);
or UO_797 (O_797,N_19862,N_19865);
xnor UO_798 (O_798,N_19693,N_19732);
xnor UO_799 (O_799,N_19168,N_19924);
nor UO_800 (O_800,N_19585,N_19662);
or UO_801 (O_801,N_19949,N_19178);
or UO_802 (O_802,N_19418,N_19015);
nand UO_803 (O_803,N_19883,N_19931);
xor UO_804 (O_804,N_19898,N_19019);
nor UO_805 (O_805,N_19019,N_19136);
nor UO_806 (O_806,N_19967,N_19185);
or UO_807 (O_807,N_19892,N_19732);
xor UO_808 (O_808,N_19429,N_19039);
and UO_809 (O_809,N_19965,N_19019);
or UO_810 (O_810,N_19993,N_19026);
nor UO_811 (O_811,N_19000,N_19606);
nand UO_812 (O_812,N_19395,N_19927);
or UO_813 (O_813,N_19992,N_19942);
nor UO_814 (O_814,N_19773,N_19892);
or UO_815 (O_815,N_19280,N_19785);
and UO_816 (O_816,N_19148,N_19170);
nor UO_817 (O_817,N_19574,N_19363);
or UO_818 (O_818,N_19793,N_19224);
nand UO_819 (O_819,N_19328,N_19857);
xnor UO_820 (O_820,N_19714,N_19862);
nand UO_821 (O_821,N_19613,N_19771);
or UO_822 (O_822,N_19912,N_19000);
or UO_823 (O_823,N_19254,N_19288);
or UO_824 (O_824,N_19775,N_19271);
nand UO_825 (O_825,N_19297,N_19268);
and UO_826 (O_826,N_19026,N_19962);
or UO_827 (O_827,N_19879,N_19894);
xor UO_828 (O_828,N_19635,N_19486);
and UO_829 (O_829,N_19750,N_19162);
and UO_830 (O_830,N_19123,N_19801);
nor UO_831 (O_831,N_19695,N_19806);
nor UO_832 (O_832,N_19259,N_19231);
nor UO_833 (O_833,N_19827,N_19532);
and UO_834 (O_834,N_19552,N_19200);
xor UO_835 (O_835,N_19785,N_19054);
and UO_836 (O_836,N_19444,N_19967);
nand UO_837 (O_837,N_19472,N_19409);
xor UO_838 (O_838,N_19886,N_19521);
xor UO_839 (O_839,N_19918,N_19131);
and UO_840 (O_840,N_19503,N_19897);
xnor UO_841 (O_841,N_19981,N_19156);
nand UO_842 (O_842,N_19798,N_19890);
nor UO_843 (O_843,N_19615,N_19941);
nor UO_844 (O_844,N_19505,N_19788);
and UO_845 (O_845,N_19533,N_19430);
nor UO_846 (O_846,N_19610,N_19309);
and UO_847 (O_847,N_19373,N_19951);
xnor UO_848 (O_848,N_19800,N_19043);
or UO_849 (O_849,N_19497,N_19624);
nand UO_850 (O_850,N_19851,N_19036);
xor UO_851 (O_851,N_19406,N_19653);
nor UO_852 (O_852,N_19711,N_19422);
nand UO_853 (O_853,N_19249,N_19702);
nor UO_854 (O_854,N_19805,N_19299);
nand UO_855 (O_855,N_19118,N_19308);
nand UO_856 (O_856,N_19902,N_19082);
nand UO_857 (O_857,N_19060,N_19590);
or UO_858 (O_858,N_19354,N_19259);
or UO_859 (O_859,N_19289,N_19897);
xnor UO_860 (O_860,N_19062,N_19032);
nor UO_861 (O_861,N_19546,N_19452);
xnor UO_862 (O_862,N_19445,N_19134);
or UO_863 (O_863,N_19007,N_19518);
nand UO_864 (O_864,N_19421,N_19767);
nor UO_865 (O_865,N_19979,N_19328);
and UO_866 (O_866,N_19606,N_19670);
and UO_867 (O_867,N_19672,N_19562);
nor UO_868 (O_868,N_19914,N_19183);
nand UO_869 (O_869,N_19901,N_19192);
and UO_870 (O_870,N_19134,N_19128);
nor UO_871 (O_871,N_19850,N_19463);
nand UO_872 (O_872,N_19218,N_19637);
xnor UO_873 (O_873,N_19559,N_19821);
xor UO_874 (O_874,N_19856,N_19296);
nor UO_875 (O_875,N_19082,N_19694);
or UO_876 (O_876,N_19520,N_19972);
and UO_877 (O_877,N_19925,N_19409);
and UO_878 (O_878,N_19077,N_19618);
nor UO_879 (O_879,N_19313,N_19195);
and UO_880 (O_880,N_19188,N_19952);
nor UO_881 (O_881,N_19369,N_19176);
or UO_882 (O_882,N_19068,N_19086);
nor UO_883 (O_883,N_19614,N_19287);
nand UO_884 (O_884,N_19878,N_19697);
nor UO_885 (O_885,N_19122,N_19319);
nor UO_886 (O_886,N_19026,N_19371);
or UO_887 (O_887,N_19699,N_19541);
xnor UO_888 (O_888,N_19633,N_19712);
xnor UO_889 (O_889,N_19018,N_19850);
nand UO_890 (O_890,N_19841,N_19489);
and UO_891 (O_891,N_19977,N_19109);
and UO_892 (O_892,N_19330,N_19288);
or UO_893 (O_893,N_19528,N_19976);
or UO_894 (O_894,N_19324,N_19077);
xnor UO_895 (O_895,N_19508,N_19194);
xnor UO_896 (O_896,N_19373,N_19655);
nand UO_897 (O_897,N_19124,N_19995);
and UO_898 (O_898,N_19721,N_19276);
or UO_899 (O_899,N_19948,N_19351);
xor UO_900 (O_900,N_19162,N_19318);
xnor UO_901 (O_901,N_19293,N_19320);
nor UO_902 (O_902,N_19060,N_19709);
xnor UO_903 (O_903,N_19108,N_19441);
and UO_904 (O_904,N_19026,N_19075);
nand UO_905 (O_905,N_19672,N_19829);
nor UO_906 (O_906,N_19391,N_19687);
nor UO_907 (O_907,N_19075,N_19302);
nor UO_908 (O_908,N_19571,N_19164);
xnor UO_909 (O_909,N_19243,N_19765);
xnor UO_910 (O_910,N_19232,N_19400);
and UO_911 (O_911,N_19566,N_19493);
xnor UO_912 (O_912,N_19672,N_19742);
xor UO_913 (O_913,N_19295,N_19974);
nor UO_914 (O_914,N_19976,N_19364);
nand UO_915 (O_915,N_19698,N_19213);
nand UO_916 (O_916,N_19479,N_19905);
nand UO_917 (O_917,N_19780,N_19030);
nand UO_918 (O_918,N_19951,N_19715);
and UO_919 (O_919,N_19153,N_19277);
nor UO_920 (O_920,N_19599,N_19414);
nor UO_921 (O_921,N_19402,N_19368);
xnor UO_922 (O_922,N_19812,N_19745);
or UO_923 (O_923,N_19927,N_19670);
nand UO_924 (O_924,N_19740,N_19211);
and UO_925 (O_925,N_19078,N_19102);
and UO_926 (O_926,N_19774,N_19551);
nand UO_927 (O_927,N_19851,N_19629);
nand UO_928 (O_928,N_19600,N_19903);
and UO_929 (O_929,N_19034,N_19058);
xor UO_930 (O_930,N_19125,N_19535);
nand UO_931 (O_931,N_19117,N_19971);
or UO_932 (O_932,N_19998,N_19239);
nand UO_933 (O_933,N_19320,N_19861);
nand UO_934 (O_934,N_19419,N_19474);
nor UO_935 (O_935,N_19035,N_19276);
and UO_936 (O_936,N_19377,N_19151);
and UO_937 (O_937,N_19879,N_19952);
xor UO_938 (O_938,N_19056,N_19701);
nor UO_939 (O_939,N_19509,N_19953);
and UO_940 (O_940,N_19259,N_19329);
nor UO_941 (O_941,N_19933,N_19769);
and UO_942 (O_942,N_19946,N_19510);
and UO_943 (O_943,N_19319,N_19410);
xnor UO_944 (O_944,N_19618,N_19311);
nor UO_945 (O_945,N_19247,N_19527);
nand UO_946 (O_946,N_19280,N_19274);
nor UO_947 (O_947,N_19307,N_19487);
nand UO_948 (O_948,N_19637,N_19899);
nand UO_949 (O_949,N_19730,N_19424);
nand UO_950 (O_950,N_19194,N_19514);
xor UO_951 (O_951,N_19023,N_19985);
nand UO_952 (O_952,N_19476,N_19066);
and UO_953 (O_953,N_19268,N_19596);
nor UO_954 (O_954,N_19205,N_19791);
and UO_955 (O_955,N_19948,N_19571);
nor UO_956 (O_956,N_19820,N_19449);
xnor UO_957 (O_957,N_19715,N_19176);
xor UO_958 (O_958,N_19674,N_19200);
or UO_959 (O_959,N_19434,N_19979);
xnor UO_960 (O_960,N_19310,N_19382);
nor UO_961 (O_961,N_19074,N_19344);
and UO_962 (O_962,N_19529,N_19721);
or UO_963 (O_963,N_19515,N_19397);
nand UO_964 (O_964,N_19993,N_19449);
nor UO_965 (O_965,N_19520,N_19760);
xnor UO_966 (O_966,N_19813,N_19849);
xor UO_967 (O_967,N_19306,N_19844);
xnor UO_968 (O_968,N_19146,N_19616);
nor UO_969 (O_969,N_19114,N_19763);
nand UO_970 (O_970,N_19603,N_19370);
or UO_971 (O_971,N_19393,N_19627);
xnor UO_972 (O_972,N_19863,N_19388);
nor UO_973 (O_973,N_19155,N_19872);
and UO_974 (O_974,N_19456,N_19701);
or UO_975 (O_975,N_19400,N_19160);
xnor UO_976 (O_976,N_19610,N_19651);
nor UO_977 (O_977,N_19089,N_19930);
nand UO_978 (O_978,N_19034,N_19465);
nor UO_979 (O_979,N_19871,N_19451);
and UO_980 (O_980,N_19297,N_19159);
or UO_981 (O_981,N_19274,N_19886);
nor UO_982 (O_982,N_19684,N_19776);
and UO_983 (O_983,N_19669,N_19527);
and UO_984 (O_984,N_19841,N_19405);
and UO_985 (O_985,N_19347,N_19664);
xnor UO_986 (O_986,N_19119,N_19761);
xnor UO_987 (O_987,N_19404,N_19085);
xor UO_988 (O_988,N_19112,N_19251);
xor UO_989 (O_989,N_19510,N_19123);
or UO_990 (O_990,N_19952,N_19180);
nor UO_991 (O_991,N_19660,N_19280);
nor UO_992 (O_992,N_19449,N_19593);
nor UO_993 (O_993,N_19505,N_19344);
xor UO_994 (O_994,N_19357,N_19665);
and UO_995 (O_995,N_19332,N_19919);
xor UO_996 (O_996,N_19262,N_19039);
xor UO_997 (O_997,N_19942,N_19540);
or UO_998 (O_998,N_19739,N_19858);
xor UO_999 (O_999,N_19586,N_19299);
nand UO_1000 (O_1000,N_19839,N_19456);
nand UO_1001 (O_1001,N_19144,N_19656);
or UO_1002 (O_1002,N_19531,N_19277);
xnor UO_1003 (O_1003,N_19115,N_19782);
and UO_1004 (O_1004,N_19340,N_19707);
xnor UO_1005 (O_1005,N_19997,N_19911);
or UO_1006 (O_1006,N_19271,N_19065);
nor UO_1007 (O_1007,N_19530,N_19992);
xor UO_1008 (O_1008,N_19841,N_19676);
xor UO_1009 (O_1009,N_19618,N_19839);
nand UO_1010 (O_1010,N_19703,N_19172);
nor UO_1011 (O_1011,N_19550,N_19411);
or UO_1012 (O_1012,N_19475,N_19616);
nor UO_1013 (O_1013,N_19923,N_19830);
nand UO_1014 (O_1014,N_19103,N_19157);
nand UO_1015 (O_1015,N_19516,N_19251);
and UO_1016 (O_1016,N_19034,N_19100);
xor UO_1017 (O_1017,N_19329,N_19110);
nand UO_1018 (O_1018,N_19178,N_19005);
nand UO_1019 (O_1019,N_19374,N_19311);
nor UO_1020 (O_1020,N_19751,N_19696);
and UO_1021 (O_1021,N_19098,N_19759);
nor UO_1022 (O_1022,N_19124,N_19070);
nand UO_1023 (O_1023,N_19535,N_19371);
xnor UO_1024 (O_1024,N_19127,N_19934);
xor UO_1025 (O_1025,N_19715,N_19189);
and UO_1026 (O_1026,N_19276,N_19582);
nand UO_1027 (O_1027,N_19046,N_19104);
nor UO_1028 (O_1028,N_19574,N_19769);
nand UO_1029 (O_1029,N_19216,N_19096);
nor UO_1030 (O_1030,N_19220,N_19042);
xor UO_1031 (O_1031,N_19645,N_19751);
and UO_1032 (O_1032,N_19795,N_19429);
xnor UO_1033 (O_1033,N_19227,N_19544);
xor UO_1034 (O_1034,N_19131,N_19426);
xor UO_1035 (O_1035,N_19094,N_19180);
nor UO_1036 (O_1036,N_19828,N_19664);
xor UO_1037 (O_1037,N_19398,N_19881);
and UO_1038 (O_1038,N_19488,N_19374);
nand UO_1039 (O_1039,N_19461,N_19262);
or UO_1040 (O_1040,N_19587,N_19256);
nor UO_1041 (O_1041,N_19464,N_19288);
nor UO_1042 (O_1042,N_19721,N_19049);
and UO_1043 (O_1043,N_19447,N_19710);
and UO_1044 (O_1044,N_19658,N_19603);
nand UO_1045 (O_1045,N_19028,N_19805);
nor UO_1046 (O_1046,N_19515,N_19988);
nand UO_1047 (O_1047,N_19453,N_19380);
xor UO_1048 (O_1048,N_19696,N_19323);
and UO_1049 (O_1049,N_19590,N_19276);
nor UO_1050 (O_1050,N_19700,N_19991);
xnor UO_1051 (O_1051,N_19497,N_19613);
or UO_1052 (O_1052,N_19529,N_19466);
nand UO_1053 (O_1053,N_19455,N_19357);
and UO_1054 (O_1054,N_19008,N_19927);
and UO_1055 (O_1055,N_19762,N_19236);
xnor UO_1056 (O_1056,N_19064,N_19666);
xor UO_1057 (O_1057,N_19883,N_19645);
nor UO_1058 (O_1058,N_19920,N_19685);
and UO_1059 (O_1059,N_19792,N_19478);
nand UO_1060 (O_1060,N_19471,N_19294);
or UO_1061 (O_1061,N_19782,N_19324);
nand UO_1062 (O_1062,N_19594,N_19387);
nor UO_1063 (O_1063,N_19972,N_19061);
nand UO_1064 (O_1064,N_19434,N_19265);
or UO_1065 (O_1065,N_19437,N_19336);
and UO_1066 (O_1066,N_19237,N_19296);
xor UO_1067 (O_1067,N_19390,N_19234);
nor UO_1068 (O_1068,N_19083,N_19868);
xor UO_1069 (O_1069,N_19874,N_19250);
and UO_1070 (O_1070,N_19492,N_19573);
nor UO_1071 (O_1071,N_19147,N_19728);
nand UO_1072 (O_1072,N_19103,N_19499);
and UO_1073 (O_1073,N_19120,N_19897);
nand UO_1074 (O_1074,N_19418,N_19692);
xor UO_1075 (O_1075,N_19756,N_19691);
xnor UO_1076 (O_1076,N_19798,N_19183);
or UO_1077 (O_1077,N_19661,N_19007);
or UO_1078 (O_1078,N_19725,N_19276);
nor UO_1079 (O_1079,N_19146,N_19343);
nor UO_1080 (O_1080,N_19042,N_19776);
and UO_1081 (O_1081,N_19322,N_19134);
or UO_1082 (O_1082,N_19966,N_19474);
or UO_1083 (O_1083,N_19002,N_19107);
or UO_1084 (O_1084,N_19517,N_19179);
nand UO_1085 (O_1085,N_19816,N_19083);
and UO_1086 (O_1086,N_19783,N_19869);
and UO_1087 (O_1087,N_19971,N_19701);
nand UO_1088 (O_1088,N_19560,N_19447);
nand UO_1089 (O_1089,N_19598,N_19428);
and UO_1090 (O_1090,N_19315,N_19783);
or UO_1091 (O_1091,N_19204,N_19591);
or UO_1092 (O_1092,N_19637,N_19621);
or UO_1093 (O_1093,N_19123,N_19632);
xnor UO_1094 (O_1094,N_19018,N_19370);
nand UO_1095 (O_1095,N_19231,N_19277);
xnor UO_1096 (O_1096,N_19614,N_19168);
xnor UO_1097 (O_1097,N_19229,N_19440);
and UO_1098 (O_1098,N_19144,N_19451);
and UO_1099 (O_1099,N_19347,N_19093);
nand UO_1100 (O_1100,N_19111,N_19077);
and UO_1101 (O_1101,N_19599,N_19202);
or UO_1102 (O_1102,N_19823,N_19430);
xnor UO_1103 (O_1103,N_19232,N_19951);
or UO_1104 (O_1104,N_19346,N_19445);
nor UO_1105 (O_1105,N_19996,N_19870);
or UO_1106 (O_1106,N_19173,N_19212);
and UO_1107 (O_1107,N_19478,N_19249);
or UO_1108 (O_1108,N_19606,N_19525);
xor UO_1109 (O_1109,N_19866,N_19944);
nor UO_1110 (O_1110,N_19192,N_19904);
xor UO_1111 (O_1111,N_19872,N_19574);
or UO_1112 (O_1112,N_19620,N_19251);
nand UO_1113 (O_1113,N_19103,N_19584);
nand UO_1114 (O_1114,N_19669,N_19892);
or UO_1115 (O_1115,N_19957,N_19248);
nor UO_1116 (O_1116,N_19879,N_19834);
xor UO_1117 (O_1117,N_19783,N_19481);
xor UO_1118 (O_1118,N_19797,N_19831);
nor UO_1119 (O_1119,N_19875,N_19595);
nand UO_1120 (O_1120,N_19139,N_19509);
nor UO_1121 (O_1121,N_19999,N_19616);
nand UO_1122 (O_1122,N_19316,N_19658);
nand UO_1123 (O_1123,N_19178,N_19905);
or UO_1124 (O_1124,N_19103,N_19467);
nor UO_1125 (O_1125,N_19329,N_19744);
and UO_1126 (O_1126,N_19528,N_19014);
nand UO_1127 (O_1127,N_19918,N_19521);
or UO_1128 (O_1128,N_19208,N_19360);
or UO_1129 (O_1129,N_19949,N_19894);
and UO_1130 (O_1130,N_19959,N_19036);
and UO_1131 (O_1131,N_19073,N_19567);
or UO_1132 (O_1132,N_19524,N_19370);
or UO_1133 (O_1133,N_19618,N_19709);
nor UO_1134 (O_1134,N_19614,N_19753);
or UO_1135 (O_1135,N_19447,N_19149);
or UO_1136 (O_1136,N_19263,N_19083);
nand UO_1137 (O_1137,N_19387,N_19896);
xnor UO_1138 (O_1138,N_19397,N_19143);
nand UO_1139 (O_1139,N_19413,N_19487);
and UO_1140 (O_1140,N_19022,N_19297);
and UO_1141 (O_1141,N_19017,N_19751);
nor UO_1142 (O_1142,N_19853,N_19733);
and UO_1143 (O_1143,N_19550,N_19097);
xor UO_1144 (O_1144,N_19063,N_19809);
or UO_1145 (O_1145,N_19117,N_19047);
xnor UO_1146 (O_1146,N_19674,N_19900);
and UO_1147 (O_1147,N_19159,N_19944);
xor UO_1148 (O_1148,N_19057,N_19434);
or UO_1149 (O_1149,N_19020,N_19334);
nand UO_1150 (O_1150,N_19151,N_19550);
nand UO_1151 (O_1151,N_19942,N_19053);
or UO_1152 (O_1152,N_19147,N_19457);
nor UO_1153 (O_1153,N_19095,N_19031);
xor UO_1154 (O_1154,N_19208,N_19745);
xor UO_1155 (O_1155,N_19171,N_19616);
nor UO_1156 (O_1156,N_19310,N_19527);
nor UO_1157 (O_1157,N_19782,N_19049);
and UO_1158 (O_1158,N_19927,N_19997);
or UO_1159 (O_1159,N_19987,N_19773);
xor UO_1160 (O_1160,N_19001,N_19245);
or UO_1161 (O_1161,N_19983,N_19179);
nand UO_1162 (O_1162,N_19161,N_19460);
or UO_1163 (O_1163,N_19692,N_19024);
and UO_1164 (O_1164,N_19187,N_19611);
xor UO_1165 (O_1165,N_19240,N_19840);
and UO_1166 (O_1166,N_19664,N_19617);
xnor UO_1167 (O_1167,N_19002,N_19293);
and UO_1168 (O_1168,N_19566,N_19742);
xor UO_1169 (O_1169,N_19230,N_19491);
or UO_1170 (O_1170,N_19005,N_19582);
xnor UO_1171 (O_1171,N_19084,N_19500);
nand UO_1172 (O_1172,N_19608,N_19171);
nand UO_1173 (O_1173,N_19826,N_19927);
nor UO_1174 (O_1174,N_19345,N_19201);
and UO_1175 (O_1175,N_19131,N_19742);
and UO_1176 (O_1176,N_19132,N_19885);
or UO_1177 (O_1177,N_19662,N_19646);
xnor UO_1178 (O_1178,N_19585,N_19140);
nand UO_1179 (O_1179,N_19952,N_19334);
and UO_1180 (O_1180,N_19596,N_19674);
nor UO_1181 (O_1181,N_19870,N_19321);
nor UO_1182 (O_1182,N_19398,N_19401);
nor UO_1183 (O_1183,N_19547,N_19757);
or UO_1184 (O_1184,N_19998,N_19696);
and UO_1185 (O_1185,N_19929,N_19235);
or UO_1186 (O_1186,N_19252,N_19653);
and UO_1187 (O_1187,N_19969,N_19889);
xnor UO_1188 (O_1188,N_19850,N_19172);
xnor UO_1189 (O_1189,N_19134,N_19854);
nand UO_1190 (O_1190,N_19379,N_19183);
and UO_1191 (O_1191,N_19349,N_19125);
nor UO_1192 (O_1192,N_19591,N_19536);
and UO_1193 (O_1193,N_19014,N_19517);
nor UO_1194 (O_1194,N_19042,N_19991);
xnor UO_1195 (O_1195,N_19671,N_19271);
or UO_1196 (O_1196,N_19911,N_19387);
and UO_1197 (O_1197,N_19759,N_19745);
nand UO_1198 (O_1198,N_19373,N_19901);
nand UO_1199 (O_1199,N_19245,N_19920);
nand UO_1200 (O_1200,N_19819,N_19670);
nor UO_1201 (O_1201,N_19955,N_19569);
nor UO_1202 (O_1202,N_19302,N_19886);
or UO_1203 (O_1203,N_19133,N_19660);
nand UO_1204 (O_1204,N_19476,N_19683);
and UO_1205 (O_1205,N_19632,N_19030);
or UO_1206 (O_1206,N_19596,N_19350);
xor UO_1207 (O_1207,N_19438,N_19272);
nor UO_1208 (O_1208,N_19282,N_19004);
nor UO_1209 (O_1209,N_19286,N_19901);
xnor UO_1210 (O_1210,N_19278,N_19282);
xor UO_1211 (O_1211,N_19484,N_19388);
xnor UO_1212 (O_1212,N_19887,N_19026);
and UO_1213 (O_1213,N_19766,N_19012);
nand UO_1214 (O_1214,N_19069,N_19251);
nor UO_1215 (O_1215,N_19143,N_19814);
and UO_1216 (O_1216,N_19696,N_19777);
or UO_1217 (O_1217,N_19483,N_19911);
xnor UO_1218 (O_1218,N_19675,N_19215);
nand UO_1219 (O_1219,N_19087,N_19435);
or UO_1220 (O_1220,N_19977,N_19026);
xnor UO_1221 (O_1221,N_19686,N_19532);
xnor UO_1222 (O_1222,N_19564,N_19230);
and UO_1223 (O_1223,N_19140,N_19498);
nor UO_1224 (O_1224,N_19422,N_19529);
and UO_1225 (O_1225,N_19084,N_19216);
or UO_1226 (O_1226,N_19027,N_19464);
nand UO_1227 (O_1227,N_19017,N_19018);
nor UO_1228 (O_1228,N_19704,N_19418);
nand UO_1229 (O_1229,N_19723,N_19053);
nand UO_1230 (O_1230,N_19317,N_19223);
xor UO_1231 (O_1231,N_19510,N_19992);
xnor UO_1232 (O_1232,N_19598,N_19704);
and UO_1233 (O_1233,N_19328,N_19507);
nand UO_1234 (O_1234,N_19230,N_19519);
nor UO_1235 (O_1235,N_19924,N_19729);
xnor UO_1236 (O_1236,N_19478,N_19708);
xnor UO_1237 (O_1237,N_19791,N_19402);
or UO_1238 (O_1238,N_19184,N_19339);
xor UO_1239 (O_1239,N_19545,N_19676);
nand UO_1240 (O_1240,N_19562,N_19294);
xor UO_1241 (O_1241,N_19493,N_19093);
nor UO_1242 (O_1242,N_19043,N_19159);
nand UO_1243 (O_1243,N_19894,N_19168);
nor UO_1244 (O_1244,N_19536,N_19495);
nor UO_1245 (O_1245,N_19940,N_19290);
nand UO_1246 (O_1246,N_19814,N_19001);
nand UO_1247 (O_1247,N_19776,N_19429);
nor UO_1248 (O_1248,N_19605,N_19892);
and UO_1249 (O_1249,N_19647,N_19992);
and UO_1250 (O_1250,N_19884,N_19658);
and UO_1251 (O_1251,N_19338,N_19415);
xor UO_1252 (O_1252,N_19317,N_19797);
nor UO_1253 (O_1253,N_19488,N_19621);
and UO_1254 (O_1254,N_19418,N_19092);
or UO_1255 (O_1255,N_19170,N_19484);
xor UO_1256 (O_1256,N_19350,N_19009);
nand UO_1257 (O_1257,N_19662,N_19469);
or UO_1258 (O_1258,N_19034,N_19451);
nand UO_1259 (O_1259,N_19751,N_19018);
nor UO_1260 (O_1260,N_19323,N_19727);
nand UO_1261 (O_1261,N_19060,N_19990);
or UO_1262 (O_1262,N_19527,N_19064);
nand UO_1263 (O_1263,N_19506,N_19776);
or UO_1264 (O_1264,N_19876,N_19311);
nand UO_1265 (O_1265,N_19294,N_19339);
nand UO_1266 (O_1266,N_19483,N_19585);
nor UO_1267 (O_1267,N_19201,N_19061);
nor UO_1268 (O_1268,N_19409,N_19160);
and UO_1269 (O_1269,N_19800,N_19515);
or UO_1270 (O_1270,N_19998,N_19789);
xnor UO_1271 (O_1271,N_19140,N_19120);
and UO_1272 (O_1272,N_19276,N_19254);
and UO_1273 (O_1273,N_19292,N_19050);
nand UO_1274 (O_1274,N_19534,N_19103);
nand UO_1275 (O_1275,N_19902,N_19786);
nand UO_1276 (O_1276,N_19535,N_19191);
and UO_1277 (O_1277,N_19591,N_19981);
xor UO_1278 (O_1278,N_19143,N_19673);
and UO_1279 (O_1279,N_19881,N_19451);
xor UO_1280 (O_1280,N_19939,N_19550);
xnor UO_1281 (O_1281,N_19359,N_19497);
nand UO_1282 (O_1282,N_19733,N_19297);
nor UO_1283 (O_1283,N_19541,N_19907);
nor UO_1284 (O_1284,N_19718,N_19024);
nor UO_1285 (O_1285,N_19457,N_19710);
nand UO_1286 (O_1286,N_19640,N_19924);
nand UO_1287 (O_1287,N_19984,N_19467);
nor UO_1288 (O_1288,N_19880,N_19212);
nor UO_1289 (O_1289,N_19428,N_19299);
nor UO_1290 (O_1290,N_19331,N_19171);
nor UO_1291 (O_1291,N_19073,N_19556);
or UO_1292 (O_1292,N_19893,N_19333);
nand UO_1293 (O_1293,N_19587,N_19215);
or UO_1294 (O_1294,N_19996,N_19540);
nor UO_1295 (O_1295,N_19427,N_19697);
nand UO_1296 (O_1296,N_19485,N_19387);
nor UO_1297 (O_1297,N_19197,N_19850);
or UO_1298 (O_1298,N_19659,N_19020);
xor UO_1299 (O_1299,N_19904,N_19793);
xnor UO_1300 (O_1300,N_19725,N_19509);
nand UO_1301 (O_1301,N_19065,N_19253);
nand UO_1302 (O_1302,N_19137,N_19754);
nor UO_1303 (O_1303,N_19688,N_19306);
nor UO_1304 (O_1304,N_19815,N_19080);
or UO_1305 (O_1305,N_19178,N_19587);
xor UO_1306 (O_1306,N_19895,N_19975);
or UO_1307 (O_1307,N_19044,N_19182);
nor UO_1308 (O_1308,N_19821,N_19210);
nand UO_1309 (O_1309,N_19958,N_19254);
and UO_1310 (O_1310,N_19194,N_19969);
nand UO_1311 (O_1311,N_19768,N_19448);
and UO_1312 (O_1312,N_19317,N_19986);
or UO_1313 (O_1313,N_19741,N_19210);
and UO_1314 (O_1314,N_19741,N_19656);
nor UO_1315 (O_1315,N_19982,N_19397);
or UO_1316 (O_1316,N_19147,N_19219);
xor UO_1317 (O_1317,N_19041,N_19771);
and UO_1318 (O_1318,N_19266,N_19174);
or UO_1319 (O_1319,N_19801,N_19548);
and UO_1320 (O_1320,N_19127,N_19759);
xnor UO_1321 (O_1321,N_19631,N_19209);
and UO_1322 (O_1322,N_19995,N_19886);
xnor UO_1323 (O_1323,N_19106,N_19946);
and UO_1324 (O_1324,N_19206,N_19871);
nand UO_1325 (O_1325,N_19249,N_19688);
xor UO_1326 (O_1326,N_19544,N_19222);
xnor UO_1327 (O_1327,N_19336,N_19980);
xor UO_1328 (O_1328,N_19260,N_19255);
nand UO_1329 (O_1329,N_19043,N_19353);
nand UO_1330 (O_1330,N_19582,N_19483);
xor UO_1331 (O_1331,N_19868,N_19085);
or UO_1332 (O_1332,N_19193,N_19992);
or UO_1333 (O_1333,N_19105,N_19866);
nor UO_1334 (O_1334,N_19627,N_19095);
and UO_1335 (O_1335,N_19516,N_19842);
nor UO_1336 (O_1336,N_19705,N_19330);
or UO_1337 (O_1337,N_19141,N_19306);
nand UO_1338 (O_1338,N_19809,N_19596);
xnor UO_1339 (O_1339,N_19653,N_19195);
nor UO_1340 (O_1340,N_19658,N_19449);
nor UO_1341 (O_1341,N_19559,N_19873);
nor UO_1342 (O_1342,N_19384,N_19887);
and UO_1343 (O_1343,N_19024,N_19727);
xnor UO_1344 (O_1344,N_19449,N_19693);
or UO_1345 (O_1345,N_19171,N_19651);
xor UO_1346 (O_1346,N_19533,N_19339);
xnor UO_1347 (O_1347,N_19997,N_19138);
or UO_1348 (O_1348,N_19158,N_19201);
and UO_1349 (O_1349,N_19974,N_19819);
xor UO_1350 (O_1350,N_19034,N_19338);
nand UO_1351 (O_1351,N_19985,N_19782);
xnor UO_1352 (O_1352,N_19932,N_19716);
xnor UO_1353 (O_1353,N_19079,N_19678);
xor UO_1354 (O_1354,N_19473,N_19589);
xnor UO_1355 (O_1355,N_19812,N_19109);
or UO_1356 (O_1356,N_19303,N_19045);
nand UO_1357 (O_1357,N_19840,N_19276);
nor UO_1358 (O_1358,N_19987,N_19345);
nand UO_1359 (O_1359,N_19170,N_19763);
nor UO_1360 (O_1360,N_19972,N_19383);
nand UO_1361 (O_1361,N_19206,N_19650);
and UO_1362 (O_1362,N_19861,N_19823);
nor UO_1363 (O_1363,N_19683,N_19645);
xnor UO_1364 (O_1364,N_19499,N_19925);
xnor UO_1365 (O_1365,N_19355,N_19078);
or UO_1366 (O_1366,N_19247,N_19893);
and UO_1367 (O_1367,N_19662,N_19405);
nor UO_1368 (O_1368,N_19077,N_19772);
nand UO_1369 (O_1369,N_19518,N_19926);
xor UO_1370 (O_1370,N_19628,N_19065);
nand UO_1371 (O_1371,N_19540,N_19603);
nor UO_1372 (O_1372,N_19896,N_19345);
or UO_1373 (O_1373,N_19271,N_19406);
or UO_1374 (O_1374,N_19753,N_19564);
xnor UO_1375 (O_1375,N_19051,N_19077);
xor UO_1376 (O_1376,N_19674,N_19418);
nand UO_1377 (O_1377,N_19599,N_19653);
and UO_1378 (O_1378,N_19359,N_19349);
xor UO_1379 (O_1379,N_19728,N_19174);
or UO_1380 (O_1380,N_19165,N_19344);
or UO_1381 (O_1381,N_19301,N_19020);
nand UO_1382 (O_1382,N_19766,N_19127);
nor UO_1383 (O_1383,N_19254,N_19579);
xor UO_1384 (O_1384,N_19492,N_19144);
nor UO_1385 (O_1385,N_19959,N_19971);
nand UO_1386 (O_1386,N_19244,N_19901);
nor UO_1387 (O_1387,N_19427,N_19647);
nand UO_1388 (O_1388,N_19410,N_19314);
nand UO_1389 (O_1389,N_19960,N_19011);
nand UO_1390 (O_1390,N_19655,N_19494);
or UO_1391 (O_1391,N_19413,N_19285);
xor UO_1392 (O_1392,N_19744,N_19139);
nor UO_1393 (O_1393,N_19440,N_19797);
xnor UO_1394 (O_1394,N_19976,N_19930);
xor UO_1395 (O_1395,N_19504,N_19729);
nor UO_1396 (O_1396,N_19310,N_19541);
nand UO_1397 (O_1397,N_19954,N_19680);
nor UO_1398 (O_1398,N_19219,N_19068);
nor UO_1399 (O_1399,N_19904,N_19384);
or UO_1400 (O_1400,N_19272,N_19538);
nand UO_1401 (O_1401,N_19770,N_19842);
and UO_1402 (O_1402,N_19778,N_19973);
xnor UO_1403 (O_1403,N_19749,N_19507);
and UO_1404 (O_1404,N_19623,N_19903);
and UO_1405 (O_1405,N_19802,N_19755);
and UO_1406 (O_1406,N_19787,N_19325);
nor UO_1407 (O_1407,N_19666,N_19306);
xnor UO_1408 (O_1408,N_19372,N_19293);
or UO_1409 (O_1409,N_19414,N_19225);
nand UO_1410 (O_1410,N_19835,N_19239);
nand UO_1411 (O_1411,N_19560,N_19241);
or UO_1412 (O_1412,N_19054,N_19262);
nor UO_1413 (O_1413,N_19592,N_19833);
or UO_1414 (O_1414,N_19883,N_19070);
and UO_1415 (O_1415,N_19329,N_19833);
nand UO_1416 (O_1416,N_19476,N_19754);
nor UO_1417 (O_1417,N_19444,N_19897);
nor UO_1418 (O_1418,N_19547,N_19924);
and UO_1419 (O_1419,N_19855,N_19934);
or UO_1420 (O_1420,N_19486,N_19768);
xnor UO_1421 (O_1421,N_19731,N_19966);
xnor UO_1422 (O_1422,N_19372,N_19220);
xnor UO_1423 (O_1423,N_19111,N_19489);
xnor UO_1424 (O_1424,N_19030,N_19625);
and UO_1425 (O_1425,N_19440,N_19469);
or UO_1426 (O_1426,N_19514,N_19619);
xnor UO_1427 (O_1427,N_19652,N_19336);
nor UO_1428 (O_1428,N_19299,N_19913);
or UO_1429 (O_1429,N_19854,N_19382);
and UO_1430 (O_1430,N_19393,N_19949);
nand UO_1431 (O_1431,N_19548,N_19939);
and UO_1432 (O_1432,N_19016,N_19027);
or UO_1433 (O_1433,N_19698,N_19625);
nand UO_1434 (O_1434,N_19143,N_19782);
xnor UO_1435 (O_1435,N_19102,N_19413);
nand UO_1436 (O_1436,N_19432,N_19603);
and UO_1437 (O_1437,N_19655,N_19642);
and UO_1438 (O_1438,N_19554,N_19674);
xor UO_1439 (O_1439,N_19618,N_19404);
nor UO_1440 (O_1440,N_19986,N_19425);
nor UO_1441 (O_1441,N_19759,N_19291);
xor UO_1442 (O_1442,N_19837,N_19595);
nor UO_1443 (O_1443,N_19914,N_19587);
and UO_1444 (O_1444,N_19442,N_19595);
nor UO_1445 (O_1445,N_19108,N_19126);
xor UO_1446 (O_1446,N_19711,N_19397);
and UO_1447 (O_1447,N_19097,N_19382);
and UO_1448 (O_1448,N_19557,N_19366);
xor UO_1449 (O_1449,N_19065,N_19155);
nor UO_1450 (O_1450,N_19923,N_19904);
or UO_1451 (O_1451,N_19791,N_19542);
nor UO_1452 (O_1452,N_19828,N_19787);
or UO_1453 (O_1453,N_19062,N_19350);
nand UO_1454 (O_1454,N_19239,N_19982);
and UO_1455 (O_1455,N_19403,N_19418);
nor UO_1456 (O_1456,N_19081,N_19259);
and UO_1457 (O_1457,N_19498,N_19567);
nand UO_1458 (O_1458,N_19056,N_19171);
xor UO_1459 (O_1459,N_19272,N_19542);
xor UO_1460 (O_1460,N_19646,N_19323);
or UO_1461 (O_1461,N_19495,N_19466);
and UO_1462 (O_1462,N_19109,N_19247);
or UO_1463 (O_1463,N_19996,N_19927);
and UO_1464 (O_1464,N_19920,N_19182);
nand UO_1465 (O_1465,N_19190,N_19283);
nand UO_1466 (O_1466,N_19502,N_19352);
or UO_1467 (O_1467,N_19546,N_19700);
nand UO_1468 (O_1468,N_19181,N_19686);
nand UO_1469 (O_1469,N_19136,N_19782);
xor UO_1470 (O_1470,N_19028,N_19104);
nand UO_1471 (O_1471,N_19126,N_19711);
or UO_1472 (O_1472,N_19064,N_19604);
nand UO_1473 (O_1473,N_19465,N_19637);
and UO_1474 (O_1474,N_19716,N_19843);
nand UO_1475 (O_1475,N_19530,N_19148);
nor UO_1476 (O_1476,N_19146,N_19395);
xnor UO_1477 (O_1477,N_19545,N_19609);
or UO_1478 (O_1478,N_19974,N_19697);
and UO_1479 (O_1479,N_19403,N_19413);
nor UO_1480 (O_1480,N_19847,N_19321);
and UO_1481 (O_1481,N_19716,N_19232);
xnor UO_1482 (O_1482,N_19798,N_19598);
nor UO_1483 (O_1483,N_19089,N_19901);
xor UO_1484 (O_1484,N_19906,N_19725);
xnor UO_1485 (O_1485,N_19822,N_19588);
and UO_1486 (O_1486,N_19861,N_19373);
xor UO_1487 (O_1487,N_19178,N_19886);
nand UO_1488 (O_1488,N_19695,N_19003);
nand UO_1489 (O_1489,N_19939,N_19137);
xnor UO_1490 (O_1490,N_19140,N_19924);
and UO_1491 (O_1491,N_19514,N_19574);
and UO_1492 (O_1492,N_19010,N_19990);
nand UO_1493 (O_1493,N_19544,N_19020);
xor UO_1494 (O_1494,N_19419,N_19053);
nor UO_1495 (O_1495,N_19890,N_19654);
nor UO_1496 (O_1496,N_19510,N_19995);
or UO_1497 (O_1497,N_19748,N_19797);
xor UO_1498 (O_1498,N_19083,N_19038);
nor UO_1499 (O_1499,N_19557,N_19739);
nand UO_1500 (O_1500,N_19983,N_19702);
nor UO_1501 (O_1501,N_19811,N_19999);
and UO_1502 (O_1502,N_19108,N_19369);
or UO_1503 (O_1503,N_19242,N_19503);
or UO_1504 (O_1504,N_19118,N_19261);
nor UO_1505 (O_1505,N_19926,N_19369);
and UO_1506 (O_1506,N_19022,N_19466);
nor UO_1507 (O_1507,N_19744,N_19739);
nor UO_1508 (O_1508,N_19987,N_19780);
or UO_1509 (O_1509,N_19942,N_19180);
nor UO_1510 (O_1510,N_19954,N_19948);
nand UO_1511 (O_1511,N_19524,N_19693);
nand UO_1512 (O_1512,N_19101,N_19593);
nand UO_1513 (O_1513,N_19621,N_19306);
and UO_1514 (O_1514,N_19100,N_19917);
xor UO_1515 (O_1515,N_19666,N_19035);
or UO_1516 (O_1516,N_19218,N_19934);
or UO_1517 (O_1517,N_19800,N_19404);
xnor UO_1518 (O_1518,N_19332,N_19211);
and UO_1519 (O_1519,N_19324,N_19239);
or UO_1520 (O_1520,N_19760,N_19994);
and UO_1521 (O_1521,N_19964,N_19229);
nand UO_1522 (O_1522,N_19994,N_19880);
nor UO_1523 (O_1523,N_19029,N_19993);
xor UO_1524 (O_1524,N_19647,N_19918);
and UO_1525 (O_1525,N_19161,N_19860);
nor UO_1526 (O_1526,N_19818,N_19621);
nand UO_1527 (O_1527,N_19957,N_19684);
and UO_1528 (O_1528,N_19949,N_19977);
xor UO_1529 (O_1529,N_19889,N_19506);
nor UO_1530 (O_1530,N_19392,N_19633);
nor UO_1531 (O_1531,N_19128,N_19828);
xor UO_1532 (O_1532,N_19671,N_19388);
nand UO_1533 (O_1533,N_19077,N_19935);
xnor UO_1534 (O_1534,N_19654,N_19192);
or UO_1535 (O_1535,N_19719,N_19596);
and UO_1536 (O_1536,N_19464,N_19655);
xor UO_1537 (O_1537,N_19194,N_19576);
nand UO_1538 (O_1538,N_19741,N_19984);
or UO_1539 (O_1539,N_19608,N_19733);
nor UO_1540 (O_1540,N_19492,N_19012);
and UO_1541 (O_1541,N_19808,N_19128);
nor UO_1542 (O_1542,N_19960,N_19744);
nand UO_1543 (O_1543,N_19139,N_19783);
nand UO_1544 (O_1544,N_19508,N_19287);
nand UO_1545 (O_1545,N_19315,N_19110);
nor UO_1546 (O_1546,N_19452,N_19197);
xnor UO_1547 (O_1547,N_19538,N_19429);
xnor UO_1548 (O_1548,N_19015,N_19646);
xor UO_1549 (O_1549,N_19225,N_19216);
and UO_1550 (O_1550,N_19394,N_19496);
nand UO_1551 (O_1551,N_19068,N_19733);
xor UO_1552 (O_1552,N_19770,N_19505);
xor UO_1553 (O_1553,N_19593,N_19459);
and UO_1554 (O_1554,N_19237,N_19347);
or UO_1555 (O_1555,N_19934,N_19105);
nor UO_1556 (O_1556,N_19924,N_19859);
xor UO_1557 (O_1557,N_19620,N_19295);
or UO_1558 (O_1558,N_19791,N_19897);
nor UO_1559 (O_1559,N_19917,N_19421);
or UO_1560 (O_1560,N_19690,N_19477);
and UO_1561 (O_1561,N_19672,N_19348);
nand UO_1562 (O_1562,N_19373,N_19069);
xor UO_1563 (O_1563,N_19611,N_19102);
nor UO_1564 (O_1564,N_19741,N_19971);
or UO_1565 (O_1565,N_19618,N_19733);
nor UO_1566 (O_1566,N_19883,N_19213);
nand UO_1567 (O_1567,N_19147,N_19407);
nor UO_1568 (O_1568,N_19838,N_19653);
or UO_1569 (O_1569,N_19977,N_19787);
nand UO_1570 (O_1570,N_19640,N_19534);
xnor UO_1571 (O_1571,N_19231,N_19009);
nand UO_1572 (O_1572,N_19923,N_19238);
nand UO_1573 (O_1573,N_19755,N_19164);
nand UO_1574 (O_1574,N_19638,N_19061);
and UO_1575 (O_1575,N_19421,N_19636);
xnor UO_1576 (O_1576,N_19038,N_19397);
or UO_1577 (O_1577,N_19536,N_19094);
or UO_1578 (O_1578,N_19353,N_19261);
nor UO_1579 (O_1579,N_19445,N_19547);
nor UO_1580 (O_1580,N_19738,N_19177);
nand UO_1581 (O_1581,N_19198,N_19869);
or UO_1582 (O_1582,N_19103,N_19781);
xnor UO_1583 (O_1583,N_19610,N_19923);
nor UO_1584 (O_1584,N_19127,N_19158);
xor UO_1585 (O_1585,N_19307,N_19551);
nand UO_1586 (O_1586,N_19715,N_19416);
and UO_1587 (O_1587,N_19627,N_19400);
and UO_1588 (O_1588,N_19836,N_19097);
and UO_1589 (O_1589,N_19219,N_19074);
xor UO_1590 (O_1590,N_19691,N_19956);
nor UO_1591 (O_1591,N_19676,N_19287);
and UO_1592 (O_1592,N_19975,N_19305);
and UO_1593 (O_1593,N_19077,N_19204);
or UO_1594 (O_1594,N_19907,N_19182);
nor UO_1595 (O_1595,N_19699,N_19157);
nand UO_1596 (O_1596,N_19749,N_19690);
nor UO_1597 (O_1597,N_19697,N_19331);
nand UO_1598 (O_1598,N_19732,N_19713);
nand UO_1599 (O_1599,N_19096,N_19547);
nand UO_1600 (O_1600,N_19066,N_19783);
xor UO_1601 (O_1601,N_19215,N_19189);
and UO_1602 (O_1602,N_19266,N_19779);
nor UO_1603 (O_1603,N_19699,N_19735);
xor UO_1604 (O_1604,N_19165,N_19949);
nand UO_1605 (O_1605,N_19824,N_19967);
or UO_1606 (O_1606,N_19671,N_19469);
and UO_1607 (O_1607,N_19636,N_19546);
xor UO_1608 (O_1608,N_19607,N_19787);
or UO_1609 (O_1609,N_19184,N_19998);
nand UO_1610 (O_1610,N_19351,N_19716);
nor UO_1611 (O_1611,N_19851,N_19152);
or UO_1612 (O_1612,N_19241,N_19114);
nor UO_1613 (O_1613,N_19805,N_19561);
and UO_1614 (O_1614,N_19015,N_19707);
or UO_1615 (O_1615,N_19250,N_19855);
and UO_1616 (O_1616,N_19869,N_19549);
or UO_1617 (O_1617,N_19725,N_19642);
and UO_1618 (O_1618,N_19153,N_19089);
nor UO_1619 (O_1619,N_19691,N_19185);
or UO_1620 (O_1620,N_19506,N_19251);
xor UO_1621 (O_1621,N_19620,N_19416);
nor UO_1622 (O_1622,N_19643,N_19885);
nor UO_1623 (O_1623,N_19223,N_19778);
nor UO_1624 (O_1624,N_19743,N_19862);
or UO_1625 (O_1625,N_19868,N_19465);
nand UO_1626 (O_1626,N_19883,N_19643);
nand UO_1627 (O_1627,N_19089,N_19362);
xor UO_1628 (O_1628,N_19473,N_19214);
and UO_1629 (O_1629,N_19667,N_19395);
nand UO_1630 (O_1630,N_19460,N_19273);
nand UO_1631 (O_1631,N_19736,N_19144);
xor UO_1632 (O_1632,N_19024,N_19437);
and UO_1633 (O_1633,N_19312,N_19713);
nor UO_1634 (O_1634,N_19547,N_19286);
or UO_1635 (O_1635,N_19888,N_19264);
nor UO_1636 (O_1636,N_19848,N_19593);
nor UO_1637 (O_1637,N_19510,N_19768);
or UO_1638 (O_1638,N_19978,N_19742);
nor UO_1639 (O_1639,N_19150,N_19784);
or UO_1640 (O_1640,N_19735,N_19509);
and UO_1641 (O_1641,N_19296,N_19469);
and UO_1642 (O_1642,N_19515,N_19253);
xnor UO_1643 (O_1643,N_19111,N_19945);
or UO_1644 (O_1644,N_19600,N_19398);
and UO_1645 (O_1645,N_19371,N_19283);
xnor UO_1646 (O_1646,N_19004,N_19019);
nand UO_1647 (O_1647,N_19583,N_19741);
xnor UO_1648 (O_1648,N_19513,N_19999);
or UO_1649 (O_1649,N_19400,N_19624);
nand UO_1650 (O_1650,N_19545,N_19631);
nor UO_1651 (O_1651,N_19570,N_19821);
nand UO_1652 (O_1652,N_19426,N_19514);
or UO_1653 (O_1653,N_19709,N_19094);
xnor UO_1654 (O_1654,N_19485,N_19258);
nor UO_1655 (O_1655,N_19627,N_19911);
and UO_1656 (O_1656,N_19172,N_19525);
and UO_1657 (O_1657,N_19677,N_19132);
nor UO_1658 (O_1658,N_19532,N_19432);
nand UO_1659 (O_1659,N_19000,N_19717);
nand UO_1660 (O_1660,N_19821,N_19836);
nor UO_1661 (O_1661,N_19381,N_19730);
and UO_1662 (O_1662,N_19310,N_19126);
nand UO_1663 (O_1663,N_19928,N_19188);
xnor UO_1664 (O_1664,N_19460,N_19700);
and UO_1665 (O_1665,N_19682,N_19430);
and UO_1666 (O_1666,N_19152,N_19648);
nor UO_1667 (O_1667,N_19206,N_19792);
and UO_1668 (O_1668,N_19723,N_19507);
nand UO_1669 (O_1669,N_19319,N_19921);
nand UO_1670 (O_1670,N_19571,N_19161);
nor UO_1671 (O_1671,N_19160,N_19892);
nor UO_1672 (O_1672,N_19326,N_19846);
xor UO_1673 (O_1673,N_19928,N_19235);
xor UO_1674 (O_1674,N_19797,N_19901);
and UO_1675 (O_1675,N_19540,N_19107);
xor UO_1676 (O_1676,N_19086,N_19635);
and UO_1677 (O_1677,N_19863,N_19595);
and UO_1678 (O_1678,N_19671,N_19500);
or UO_1679 (O_1679,N_19273,N_19840);
and UO_1680 (O_1680,N_19241,N_19163);
xnor UO_1681 (O_1681,N_19478,N_19178);
xnor UO_1682 (O_1682,N_19322,N_19607);
nor UO_1683 (O_1683,N_19862,N_19087);
nor UO_1684 (O_1684,N_19664,N_19112);
xor UO_1685 (O_1685,N_19273,N_19928);
or UO_1686 (O_1686,N_19295,N_19187);
and UO_1687 (O_1687,N_19970,N_19190);
nand UO_1688 (O_1688,N_19259,N_19195);
and UO_1689 (O_1689,N_19911,N_19059);
nor UO_1690 (O_1690,N_19641,N_19603);
and UO_1691 (O_1691,N_19157,N_19292);
and UO_1692 (O_1692,N_19472,N_19844);
nor UO_1693 (O_1693,N_19725,N_19298);
or UO_1694 (O_1694,N_19210,N_19543);
nand UO_1695 (O_1695,N_19682,N_19470);
nand UO_1696 (O_1696,N_19437,N_19260);
nand UO_1697 (O_1697,N_19648,N_19763);
or UO_1698 (O_1698,N_19698,N_19795);
and UO_1699 (O_1699,N_19947,N_19103);
or UO_1700 (O_1700,N_19200,N_19162);
and UO_1701 (O_1701,N_19895,N_19747);
or UO_1702 (O_1702,N_19453,N_19197);
xor UO_1703 (O_1703,N_19312,N_19591);
xnor UO_1704 (O_1704,N_19060,N_19391);
xnor UO_1705 (O_1705,N_19175,N_19805);
and UO_1706 (O_1706,N_19457,N_19604);
xnor UO_1707 (O_1707,N_19938,N_19940);
and UO_1708 (O_1708,N_19117,N_19100);
and UO_1709 (O_1709,N_19484,N_19461);
xor UO_1710 (O_1710,N_19122,N_19204);
xnor UO_1711 (O_1711,N_19175,N_19768);
nand UO_1712 (O_1712,N_19863,N_19647);
nor UO_1713 (O_1713,N_19452,N_19635);
and UO_1714 (O_1714,N_19137,N_19989);
nand UO_1715 (O_1715,N_19606,N_19944);
xnor UO_1716 (O_1716,N_19476,N_19119);
nor UO_1717 (O_1717,N_19865,N_19187);
or UO_1718 (O_1718,N_19019,N_19682);
and UO_1719 (O_1719,N_19860,N_19697);
nor UO_1720 (O_1720,N_19537,N_19846);
xnor UO_1721 (O_1721,N_19551,N_19563);
and UO_1722 (O_1722,N_19538,N_19325);
or UO_1723 (O_1723,N_19953,N_19667);
and UO_1724 (O_1724,N_19250,N_19079);
nor UO_1725 (O_1725,N_19972,N_19829);
nor UO_1726 (O_1726,N_19616,N_19785);
and UO_1727 (O_1727,N_19992,N_19038);
nand UO_1728 (O_1728,N_19016,N_19896);
and UO_1729 (O_1729,N_19823,N_19189);
nand UO_1730 (O_1730,N_19079,N_19440);
or UO_1731 (O_1731,N_19216,N_19511);
xor UO_1732 (O_1732,N_19574,N_19324);
xor UO_1733 (O_1733,N_19207,N_19951);
nor UO_1734 (O_1734,N_19940,N_19089);
nand UO_1735 (O_1735,N_19862,N_19285);
nand UO_1736 (O_1736,N_19512,N_19592);
nor UO_1737 (O_1737,N_19721,N_19898);
xnor UO_1738 (O_1738,N_19452,N_19530);
xnor UO_1739 (O_1739,N_19190,N_19100);
xnor UO_1740 (O_1740,N_19079,N_19477);
xnor UO_1741 (O_1741,N_19541,N_19385);
and UO_1742 (O_1742,N_19331,N_19839);
xor UO_1743 (O_1743,N_19108,N_19580);
or UO_1744 (O_1744,N_19214,N_19563);
and UO_1745 (O_1745,N_19712,N_19563);
and UO_1746 (O_1746,N_19819,N_19244);
nand UO_1747 (O_1747,N_19795,N_19543);
xor UO_1748 (O_1748,N_19288,N_19655);
nor UO_1749 (O_1749,N_19906,N_19025);
xor UO_1750 (O_1750,N_19917,N_19399);
nor UO_1751 (O_1751,N_19588,N_19278);
or UO_1752 (O_1752,N_19467,N_19595);
xor UO_1753 (O_1753,N_19958,N_19055);
xnor UO_1754 (O_1754,N_19346,N_19884);
or UO_1755 (O_1755,N_19388,N_19335);
xnor UO_1756 (O_1756,N_19635,N_19433);
and UO_1757 (O_1757,N_19105,N_19874);
nand UO_1758 (O_1758,N_19832,N_19039);
xor UO_1759 (O_1759,N_19575,N_19986);
xor UO_1760 (O_1760,N_19042,N_19184);
nand UO_1761 (O_1761,N_19144,N_19939);
xor UO_1762 (O_1762,N_19361,N_19427);
nor UO_1763 (O_1763,N_19028,N_19232);
nand UO_1764 (O_1764,N_19494,N_19614);
or UO_1765 (O_1765,N_19641,N_19563);
xor UO_1766 (O_1766,N_19405,N_19941);
nor UO_1767 (O_1767,N_19923,N_19347);
or UO_1768 (O_1768,N_19629,N_19485);
or UO_1769 (O_1769,N_19227,N_19599);
xnor UO_1770 (O_1770,N_19476,N_19573);
and UO_1771 (O_1771,N_19252,N_19408);
and UO_1772 (O_1772,N_19934,N_19356);
xor UO_1773 (O_1773,N_19367,N_19252);
nor UO_1774 (O_1774,N_19139,N_19958);
and UO_1775 (O_1775,N_19909,N_19209);
xor UO_1776 (O_1776,N_19944,N_19568);
and UO_1777 (O_1777,N_19740,N_19342);
or UO_1778 (O_1778,N_19691,N_19612);
or UO_1779 (O_1779,N_19299,N_19848);
xnor UO_1780 (O_1780,N_19607,N_19838);
nand UO_1781 (O_1781,N_19029,N_19690);
and UO_1782 (O_1782,N_19627,N_19963);
and UO_1783 (O_1783,N_19632,N_19759);
and UO_1784 (O_1784,N_19856,N_19537);
nor UO_1785 (O_1785,N_19561,N_19456);
and UO_1786 (O_1786,N_19062,N_19236);
nor UO_1787 (O_1787,N_19679,N_19824);
nor UO_1788 (O_1788,N_19003,N_19081);
xor UO_1789 (O_1789,N_19559,N_19986);
and UO_1790 (O_1790,N_19891,N_19090);
nor UO_1791 (O_1791,N_19133,N_19309);
and UO_1792 (O_1792,N_19236,N_19398);
and UO_1793 (O_1793,N_19488,N_19516);
or UO_1794 (O_1794,N_19861,N_19673);
nand UO_1795 (O_1795,N_19613,N_19162);
or UO_1796 (O_1796,N_19600,N_19681);
nor UO_1797 (O_1797,N_19058,N_19195);
nor UO_1798 (O_1798,N_19166,N_19221);
nor UO_1799 (O_1799,N_19023,N_19069);
and UO_1800 (O_1800,N_19090,N_19516);
and UO_1801 (O_1801,N_19798,N_19380);
and UO_1802 (O_1802,N_19330,N_19706);
xor UO_1803 (O_1803,N_19761,N_19645);
xnor UO_1804 (O_1804,N_19469,N_19900);
nand UO_1805 (O_1805,N_19360,N_19950);
nand UO_1806 (O_1806,N_19938,N_19955);
xor UO_1807 (O_1807,N_19323,N_19006);
and UO_1808 (O_1808,N_19609,N_19746);
xor UO_1809 (O_1809,N_19339,N_19695);
nor UO_1810 (O_1810,N_19617,N_19619);
nor UO_1811 (O_1811,N_19940,N_19230);
and UO_1812 (O_1812,N_19020,N_19792);
nor UO_1813 (O_1813,N_19092,N_19685);
or UO_1814 (O_1814,N_19347,N_19048);
or UO_1815 (O_1815,N_19930,N_19155);
nor UO_1816 (O_1816,N_19295,N_19921);
nor UO_1817 (O_1817,N_19080,N_19627);
and UO_1818 (O_1818,N_19765,N_19308);
xnor UO_1819 (O_1819,N_19403,N_19598);
nor UO_1820 (O_1820,N_19665,N_19849);
or UO_1821 (O_1821,N_19438,N_19646);
or UO_1822 (O_1822,N_19810,N_19067);
and UO_1823 (O_1823,N_19297,N_19725);
nand UO_1824 (O_1824,N_19130,N_19461);
nor UO_1825 (O_1825,N_19092,N_19766);
and UO_1826 (O_1826,N_19446,N_19905);
and UO_1827 (O_1827,N_19318,N_19354);
xor UO_1828 (O_1828,N_19327,N_19729);
nand UO_1829 (O_1829,N_19542,N_19240);
nor UO_1830 (O_1830,N_19866,N_19140);
or UO_1831 (O_1831,N_19236,N_19488);
or UO_1832 (O_1832,N_19281,N_19828);
and UO_1833 (O_1833,N_19050,N_19206);
nor UO_1834 (O_1834,N_19990,N_19063);
nand UO_1835 (O_1835,N_19886,N_19643);
and UO_1836 (O_1836,N_19728,N_19996);
xor UO_1837 (O_1837,N_19848,N_19039);
or UO_1838 (O_1838,N_19205,N_19557);
nand UO_1839 (O_1839,N_19266,N_19906);
xnor UO_1840 (O_1840,N_19513,N_19922);
and UO_1841 (O_1841,N_19726,N_19303);
nand UO_1842 (O_1842,N_19830,N_19890);
and UO_1843 (O_1843,N_19912,N_19388);
nor UO_1844 (O_1844,N_19544,N_19352);
or UO_1845 (O_1845,N_19343,N_19207);
or UO_1846 (O_1846,N_19794,N_19096);
nor UO_1847 (O_1847,N_19749,N_19394);
and UO_1848 (O_1848,N_19863,N_19913);
xor UO_1849 (O_1849,N_19258,N_19891);
and UO_1850 (O_1850,N_19620,N_19045);
and UO_1851 (O_1851,N_19018,N_19298);
nor UO_1852 (O_1852,N_19611,N_19141);
nand UO_1853 (O_1853,N_19554,N_19072);
nand UO_1854 (O_1854,N_19510,N_19791);
nand UO_1855 (O_1855,N_19328,N_19808);
and UO_1856 (O_1856,N_19821,N_19368);
nand UO_1857 (O_1857,N_19303,N_19043);
xnor UO_1858 (O_1858,N_19807,N_19160);
nand UO_1859 (O_1859,N_19811,N_19473);
nand UO_1860 (O_1860,N_19876,N_19835);
nand UO_1861 (O_1861,N_19819,N_19765);
nor UO_1862 (O_1862,N_19517,N_19654);
xor UO_1863 (O_1863,N_19259,N_19998);
nand UO_1864 (O_1864,N_19966,N_19211);
and UO_1865 (O_1865,N_19849,N_19396);
nor UO_1866 (O_1866,N_19619,N_19054);
nor UO_1867 (O_1867,N_19014,N_19213);
xor UO_1868 (O_1868,N_19584,N_19674);
xor UO_1869 (O_1869,N_19960,N_19905);
nand UO_1870 (O_1870,N_19606,N_19078);
nand UO_1871 (O_1871,N_19039,N_19491);
or UO_1872 (O_1872,N_19366,N_19233);
xor UO_1873 (O_1873,N_19105,N_19550);
nor UO_1874 (O_1874,N_19105,N_19292);
and UO_1875 (O_1875,N_19800,N_19985);
and UO_1876 (O_1876,N_19951,N_19404);
nor UO_1877 (O_1877,N_19176,N_19287);
and UO_1878 (O_1878,N_19625,N_19582);
nand UO_1879 (O_1879,N_19953,N_19312);
xnor UO_1880 (O_1880,N_19402,N_19704);
nor UO_1881 (O_1881,N_19552,N_19164);
or UO_1882 (O_1882,N_19466,N_19342);
nor UO_1883 (O_1883,N_19720,N_19759);
nand UO_1884 (O_1884,N_19058,N_19600);
or UO_1885 (O_1885,N_19559,N_19693);
xnor UO_1886 (O_1886,N_19563,N_19857);
or UO_1887 (O_1887,N_19862,N_19531);
nand UO_1888 (O_1888,N_19706,N_19337);
or UO_1889 (O_1889,N_19127,N_19568);
xnor UO_1890 (O_1890,N_19602,N_19609);
and UO_1891 (O_1891,N_19080,N_19022);
nor UO_1892 (O_1892,N_19566,N_19725);
and UO_1893 (O_1893,N_19874,N_19304);
or UO_1894 (O_1894,N_19704,N_19708);
or UO_1895 (O_1895,N_19477,N_19647);
or UO_1896 (O_1896,N_19825,N_19887);
or UO_1897 (O_1897,N_19650,N_19583);
nor UO_1898 (O_1898,N_19359,N_19533);
and UO_1899 (O_1899,N_19399,N_19273);
xor UO_1900 (O_1900,N_19423,N_19579);
xnor UO_1901 (O_1901,N_19899,N_19147);
or UO_1902 (O_1902,N_19325,N_19252);
xor UO_1903 (O_1903,N_19348,N_19395);
nor UO_1904 (O_1904,N_19213,N_19467);
or UO_1905 (O_1905,N_19550,N_19648);
xnor UO_1906 (O_1906,N_19994,N_19474);
xor UO_1907 (O_1907,N_19889,N_19992);
xor UO_1908 (O_1908,N_19628,N_19206);
or UO_1909 (O_1909,N_19581,N_19870);
nor UO_1910 (O_1910,N_19557,N_19562);
nand UO_1911 (O_1911,N_19320,N_19802);
or UO_1912 (O_1912,N_19658,N_19043);
xor UO_1913 (O_1913,N_19314,N_19405);
xnor UO_1914 (O_1914,N_19400,N_19185);
nand UO_1915 (O_1915,N_19977,N_19324);
or UO_1916 (O_1916,N_19165,N_19994);
and UO_1917 (O_1917,N_19814,N_19728);
nor UO_1918 (O_1918,N_19857,N_19214);
and UO_1919 (O_1919,N_19328,N_19362);
xor UO_1920 (O_1920,N_19170,N_19215);
nand UO_1921 (O_1921,N_19613,N_19749);
and UO_1922 (O_1922,N_19312,N_19934);
xnor UO_1923 (O_1923,N_19011,N_19822);
and UO_1924 (O_1924,N_19594,N_19399);
xor UO_1925 (O_1925,N_19380,N_19623);
nand UO_1926 (O_1926,N_19209,N_19481);
and UO_1927 (O_1927,N_19356,N_19840);
nor UO_1928 (O_1928,N_19810,N_19839);
xor UO_1929 (O_1929,N_19755,N_19136);
nand UO_1930 (O_1930,N_19239,N_19526);
nand UO_1931 (O_1931,N_19147,N_19259);
xor UO_1932 (O_1932,N_19695,N_19081);
or UO_1933 (O_1933,N_19597,N_19484);
nand UO_1934 (O_1934,N_19176,N_19604);
nand UO_1935 (O_1935,N_19079,N_19646);
xnor UO_1936 (O_1936,N_19922,N_19135);
or UO_1937 (O_1937,N_19843,N_19148);
xor UO_1938 (O_1938,N_19950,N_19371);
nor UO_1939 (O_1939,N_19158,N_19562);
nor UO_1940 (O_1940,N_19165,N_19147);
xnor UO_1941 (O_1941,N_19063,N_19541);
nand UO_1942 (O_1942,N_19033,N_19247);
and UO_1943 (O_1943,N_19556,N_19999);
and UO_1944 (O_1944,N_19128,N_19165);
and UO_1945 (O_1945,N_19428,N_19028);
nor UO_1946 (O_1946,N_19105,N_19044);
or UO_1947 (O_1947,N_19881,N_19448);
xnor UO_1948 (O_1948,N_19015,N_19422);
nor UO_1949 (O_1949,N_19861,N_19930);
nand UO_1950 (O_1950,N_19936,N_19077);
xnor UO_1951 (O_1951,N_19347,N_19354);
and UO_1952 (O_1952,N_19832,N_19536);
nand UO_1953 (O_1953,N_19507,N_19440);
nand UO_1954 (O_1954,N_19490,N_19652);
and UO_1955 (O_1955,N_19344,N_19462);
nor UO_1956 (O_1956,N_19787,N_19628);
xor UO_1957 (O_1957,N_19200,N_19509);
or UO_1958 (O_1958,N_19669,N_19398);
nand UO_1959 (O_1959,N_19846,N_19228);
xor UO_1960 (O_1960,N_19153,N_19051);
and UO_1961 (O_1961,N_19627,N_19059);
nor UO_1962 (O_1962,N_19829,N_19605);
nand UO_1963 (O_1963,N_19943,N_19980);
or UO_1964 (O_1964,N_19465,N_19069);
or UO_1965 (O_1965,N_19973,N_19969);
xor UO_1966 (O_1966,N_19177,N_19657);
nand UO_1967 (O_1967,N_19507,N_19233);
and UO_1968 (O_1968,N_19446,N_19268);
or UO_1969 (O_1969,N_19175,N_19437);
or UO_1970 (O_1970,N_19712,N_19940);
and UO_1971 (O_1971,N_19614,N_19183);
and UO_1972 (O_1972,N_19774,N_19360);
or UO_1973 (O_1973,N_19739,N_19159);
nand UO_1974 (O_1974,N_19126,N_19003);
or UO_1975 (O_1975,N_19361,N_19348);
and UO_1976 (O_1976,N_19179,N_19479);
or UO_1977 (O_1977,N_19324,N_19102);
nand UO_1978 (O_1978,N_19670,N_19884);
or UO_1979 (O_1979,N_19282,N_19030);
nor UO_1980 (O_1980,N_19693,N_19321);
and UO_1981 (O_1981,N_19555,N_19753);
and UO_1982 (O_1982,N_19819,N_19281);
and UO_1983 (O_1983,N_19743,N_19703);
nand UO_1984 (O_1984,N_19393,N_19989);
nand UO_1985 (O_1985,N_19274,N_19900);
and UO_1986 (O_1986,N_19832,N_19651);
nor UO_1987 (O_1987,N_19918,N_19428);
xnor UO_1988 (O_1988,N_19554,N_19858);
and UO_1989 (O_1989,N_19718,N_19250);
nor UO_1990 (O_1990,N_19640,N_19007);
or UO_1991 (O_1991,N_19207,N_19444);
xnor UO_1992 (O_1992,N_19953,N_19278);
nor UO_1993 (O_1993,N_19342,N_19079);
or UO_1994 (O_1994,N_19913,N_19724);
xnor UO_1995 (O_1995,N_19193,N_19328);
nand UO_1996 (O_1996,N_19550,N_19107);
or UO_1997 (O_1997,N_19106,N_19033);
nand UO_1998 (O_1998,N_19718,N_19069);
nand UO_1999 (O_1999,N_19917,N_19190);
xor UO_2000 (O_2000,N_19914,N_19549);
xor UO_2001 (O_2001,N_19272,N_19626);
or UO_2002 (O_2002,N_19798,N_19375);
nand UO_2003 (O_2003,N_19462,N_19446);
xor UO_2004 (O_2004,N_19381,N_19200);
nor UO_2005 (O_2005,N_19873,N_19622);
nor UO_2006 (O_2006,N_19048,N_19351);
nor UO_2007 (O_2007,N_19943,N_19626);
xnor UO_2008 (O_2008,N_19892,N_19252);
nor UO_2009 (O_2009,N_19272,N_19380);
or UO_2010 (O_2010,N_19580,N_19843);
nand UO_2011 (O_2011,N_19744,N_19824);
nand UO_2012 (O_2012,N_19647,N_19262);
xnor UO_2013 (O_2013,N_19719,N_19482);
and UO_2014 (O_2014,N_19082,N_19995);
and UO_2015 (O_2015,N_19259,N_19709);
or UO_2016 (O_2016,N_19170,N_19298);
xor UO_2017 (O_2017,N_19891,N_19492);
and UO_2018 (O_2018,N_19897,N_19453);
nor UO_2019 (O_2019,N_19265,N_19043);
nand UO_2020 (O_2020,N_19895,N_19399);
nand UO_2021 (O_2021,N_19659,N_19253);
xor UO_2022 (O_2022,N_19330,N_19807);
nor UO_2023 (O_2023,N_19635,N_19814);
and UO_2024 (O_2024,N_19359,N_19776);
and UO_2025 (O_2025,N_19727,N_19805);
and UO_2026 (O_2026,N_19424,N_19483);
nand UO_2027 (O_2027,N_19241,N_19301);
nand UO_2028 (O_2028,N_19392,N_19060);
or UO_2029 (O_2029,N_19298,N_19364);
xnor UO_2030 (O_2030,N_19995,N_19935);
or UO_2031 (O_2031,N_19419,N_19750);
and UO_2032 (O_2032,N_19756,N_19839);
or UO_2033 (O_2033,N_19450,N_19196);
nor UO_2034 (O_2034,N_19702,N_19664);
and UO_2035 (O_2035,N_19563,N_19872);
nor UO_2036 (O_2036,N_19228,N_19643);
and UO_2037 (O_2037,N_19563,N_19494);
nor UO_2038 (O_2038,N_19475,N_19522);
or UO_2039 (O_2039,N_19450,N_19116);
nor UO_2040 (O_2040,N_19600,N_19607);
xor UO_2041 (O_2041,N_19258,N_19713);
and UO_2042 (O_2042,N_19198,N_19388);
xor UO_2043 (O_2043,N_19089,N_19312);
and UO_2044 (O_2044,N_19707,N_19690);
or UO_2045 (O_2045,N_19455,N_19318);
nor UO_2046 (O_2046,N_19166,N_19856);
nand UO_2047 (O_2047,N_19999,N_19699);
and UO_2048 (O_2048,N_19596,N_19795);
nor UO_2049 (O_2049,N_19209,N_19246);
and UO_2050 (O_2050,N_19254,N_19795);
and UO_2051 (O_2051,N_19441,N_19705);
xor UO_2052 (O_2052,N_19099,N_19260);
nand UO_2053 (O_2053,N_19943,N_19212);
and UO_2054 (O_2054,N_19082,N_19035);
nand UO_2055 (O_2055,N_19607,N_19927);
nand UO_2056 (O_2056,N_19252,N_19793);
nor UO_2057 (O_2057,N_19224,N_19088);
xnor UO_2058 (O_2058,N_19194,N_19357);
nand UO_2059 (O_2059,N_19278,N_19745);
nor UO_2060 (O_2060,N_19301,N_19765);
xor UO_2061 (O_2061,N_19450,N_19491);
nand UO_2062 (O_2062,N_19883,N_19015);
xnor UO_2063 (O_2063,N_19053,N_19275);
or UO_2064 (O_2064,N_19554,N_19865);
nand UO_2065 (O_2065,N_19042,N_19453);
nand UO_2066 (O_2066,N_19331,N_19164);
nor UO_2067 (O_2067,N_19406,N_19459);
nor UO_2068 (O_2068,N_19620,N_19474);
nor UO_2069 (O_2069,N_19218,N_19930);
xor UO_2070 (O_2070,N_19383,N_19471);
nor UO_2071 (O_2071,N_19253,N_19725);
and UO_2072 (O_2072,N_19300,N_19144);
xnor UO_2073 (O_2073,N_19593,N_19224);
and UO_2074 (O_2074,N_19386,N_19751);
nor UO_2075 (O_2075,N_19263,N_19851);
and UO_2076 (O_2076,N_19507,N_19293);
or UO_2077 (O_2077,N_19356,N_19982);
nand UO_2078 (O_2078,N_19217,N_19672);
nor UO_2079 (O_2079,N_19447,N_19482);
nor UO_2080 (O_2080,N_19647,N_19930);
nor UO_2081 (O_2081,N_19546,N_19439);
xor UO_2082 (O_2082,N_19428,N_19990);
nor UO_2083 (O_2083,N_19800,N_19088);
or UO_2084 (O_2084,N_19984,N_19601);
and UO_2085 (O_2085,N_19939,N_19553);
xnor UO_2086 (O_2086,N_19299,N_19846);
nor UO_2087 (O_2087,N_19573,N_19417);
xnor UO_2088 (O_2088,N_19924,N_19857);
and UO_2089 (O_2089,N_19513,N_19301);
xnor UO_2090 (O_2090,N_19209,N_19619);
and UO_2091 (O_2091,N_19651,N_19563);
xnor UO_2092 (O_2092,N_19641,N_19217);
nor UO_2093 (O_2093,N_19318,N_19585);
nor UO_2094 (O_2094,N_19070,N_19077);
nand UO_2095 (O_2095,N_19124,N_19395);
and UO_2096 (O_2096,N_19961,N_19983);
xor UO_2097 (O_2097,N_19111,N_19063);
nor UO_2098 (O_2098,N_19346,N_19197);
xnor UO_2099 (O_2099,N_19445,N_19616);
xor UO_2100 (O_2100,N_19774,N_19844);
or UO_2101 (O_2101,N_19513,N_19086);
or UO_2102 (O_2102,N_19312,N_19377);
nand UO_2103 (O_2103,N_19585,N_19099);
or UO_2104 (O_2104,N_19053,N_19953);
xor UO_2105 (O_2105,N_19219,N_19844);
xnor UO_2106 (O_2106,N_19351,N_19737);
or UO_2107 (O_2107,N_19472,N_19277);
or UO_2108 (O_2108,N_19640,N_19318);
and UO_2109 (O_2109,N_19960,N_19969);
and UO_2110 (O_2110,N_19192,N_19916);
nand UO_2111 (O_2111,N_19882,N_19091);
and UO_2112 (O_2112,N_19652,N_19133);
nor UO_2113 (O_2113,N_19160,N_19486);
or UO_2114 (O_2114,N_19743,N_19335);
nor UO_2115 (O_2115,N_19944,N_19141);
nand UO_2116 (O_2116,N_19038,N_19280);
nor UO_2117 (O_2117,N_19466,N_19347);
nor UO_2118 (O_2118,N_19084,N_19222);
nor UO_2119 (O_2119,N_19257,N_19194);
nand UO_2120 (O_2120,N_19388,N_19104);
nand UO_2121 (O_2121,N_19010,N_19193);
xnor UO_2122 (O_2122,N_19480,N_19640);
nand UO_2123 (O_2123,N_19284,N_19765);
nor UO_2124 (O_2124,N_19968,N_19548);
or UO_2125 (O_2125,N_19123,N_19982);
or UO_2126 (O_2126,N_19538,N_19409);
xnor UO_2127 (O_2127,N_19951,N_19056);
xnor UO_2128 (O_2128,N_19857,N_19677);
xnor UO_2129 (O_2129,N_19805,N_19839);
and UO_2130 (O_2130,N_19990,N_19624);
nor UO_2131 (O_2131,N_19927,N_19773);
and UO_2132 (O_2132,N_19361,N_19476);
nand UO_2133 (O_2133,N_19482,N_19262);
nor UO_2134 (O_2134,N_19014,N_19794);
nand UO_2135 (O_2135,N_19877,N_19307);
and UO_2136 (O_2136,N_19660,N_19128);
or UO_2137 (O_2137,N_19259,N_19675);
nor UO_2138 (O_2138,N_19808,N_19633);
xor UO_2139 (O_2139,N_19731,N_19159);
nor UO_2140 (O_2140,N_19167,N_19791);
nor UO_2141 (O_2141,N_19102,N_19122);
and UO_2142 (O_2142,N_19300,N_19959);
nand UO_2143 (O_2143,N_19095,N_19696);
or UO_2144 (O_2144,N_19123,N_19515);
and UO_2145 (O_2145,N_19657,N_19631);
xnor UO_2146 (O_2146,N_19499,N_19878);
and UO_2147 (O_2147,N_19748,N_19266);
nor UO_2148 (O_2148,N_19934,N_19671);
nor UO_2149 (O_2149,N_19966,N_19674);
xnor UO_2150 (O_2150,N_19668,N_19497);
nand UO_2151 (O_2151,N_19806,N_19001);
and UO_2152 (O_2152,N_19549,N_19365);
xnor UO_2153 (O_2153,N_19459,N_19360);
nand UO_2154 (O_2154,N_19286,N_19824);
or UO_2155 (O_2155,N_19670,N_19057);
or UO_2156 (O_2156,N_19208,N_19465);
and UO_2157 (O_2157,N_19058,N_19984);
nor UO_2158 (O_2158,N_19734,N_19804);
xor UO_2159 (O_2159,N_19308,N_19335);
xnor UO_2160 (O_2160,N_19175,N_19020);
nand UO_2161 (O_2161,N_19462,N_19142);
and UO_2162 (O_2162,N_19577,N_19401);
nor UO_2163 (O_2163,N_19526,N_19993);
or UO_2164 (O_2164,N_19474,N_19195);
xor UO_2165 (O_2165,N_19824,N_19518);
nor UO_2166 (O_2166,N_19803,N_19535);
xor UO_2167 (O_2167,N_19278,N_19615);
nor UO_2168 (O_2168,N_19378,N_19137);
nor UO_2169 (O_2169,N_19040,N_19286);
or UO_2170 (O_2170,N_19947,N_19811);
or UO_2171 (O_2171,N_19039,N_19306);
and UO_2172 (O_2172,N_19153,N_19685);
and UO_2173 (O_2173,N_19957,N_19147);
and UO_2174 (O_2174,N_19114,N_19989);
and UO_2175 (O_2175,N_19856,N_19282);
and UO_2176 (O_2176,N_19543,N_19824);
and UO_2177 (O_2177,N_19661,N_19514);
nor UO_2178 (O_2178,N_19671,N_19491);
xnor UO_2179 (O_2179,N_19122,N_19703);
and UO_2180 (O_2180,N_19028,N_19572);
xnor UO_2181 (O_2181,N_19218,N_19300);
xor UO_2182 (O_2182,N_19925,N_19299);
and UO_2183 (O_2183,N_19216,N_19542);
nor UO_2184 (O_2184,N_19973,N_19695);
nand UO_2185 (O_2185,N_19525,N_19429);
xor UO_2186 (O_2186,N_19085,N_19364);
and UO_2187 (O_2187,N_19348,N_19266);
nand UO_2188 (O_2188,N_19281,N_19413);
xnor UO_2189 (O_2189,N_19578,N_19390);
xnor UO_2190 (O_2190,N_19434,N_19437);
and UO_2191 (O_2191,N_19628,N_19783);
xnor UO_2192 (O_2192,N_19061,N_19905);
and UO_2193 (O_2193,N_19121,N_19869);
nor UO_2194 (O_2194,N_19064,N_19327);
nand UO_2195 (O_2195,N_19961,N_19448);
nand UO_2196 (O_2196,N_19211,N_19829);
or UO_2197 (O_2197,N_19021,N_19847);
and UO_2198 (O_2198,N_19232,N_19629);
nor UO_2199 (O_2199,N_19457,N_19606);
and UO_2200 (O_2200,N_19338,N_19726);
nand UO_2201 (O_2201,N_19516,N_19384);
nor UO_2202 (O_2202,N_19020,N_19350);
xnor UO_2203 (O_2203,N_19732,N_19830);
nand UO_2204 (O_2204,N_19315,N_19816);
and UO_2205 (O_2205,N_19360,N_19926);
nand UO_2206 (O_2206,N_19093,N_19526);
nand UO_2207 (O_2207,N_19656,N_19972);
and UO_2208 (O_2208,N_19471,N_19185);
nor UO_2209 (O_2209,N_19584,N_19266);
nand UO_2210 (O_2210,N_19893,N_19214);
nor UO_2211 (O_2211,N_19715,N_19583);
or UO_2212 (O_2212,N_19069,N_19715);
and UO_2213 (O_2213,N_19491,N_19150);
nand UO_2214 (O_2214,N_19616,N_19585);
xor UO_2215 (O_2215,N_19106,N_19863);
nor UO_2216 (O_2216,N_19950,N_19384);
nor UO_2217 (O_2217,N_19731,N_19382);
or UO_2218 (O_2218,N_19404,N_19355);
or UO_2219 (O_2219,N_19401,N_19688);
nand UO_2220 (O_2220,N_19361,N_19277);
nor UO_2221 (O_2221,N_19204,N_19822);
or UO_2222 (O_2222,N_19347,N_19590);
nand UO_2223 (O_2223,N_19133,N_19433);
nor UO_2224 (O_2224,N_19825,N_19550);
and UO_2225 (O_2225,N_19835,N_19684);
xor UO_2226 (O_2226,N_19526,N_19078);
nor UO_2227 (O_2227,N_19434,N_19331);
nor UO_2228 (O_2228,N_19130,N_19577);
or UO_2229 (O_2229,N_19825,N_19054);
nand UO_2230 (O_2230,N_19960,N_19490);
nand UO_2231 (O_2231,N_19496,N_19468);
or UO_2232 (O_2232,N_19615,N_19126);
and UO_2233 (O_2233,N_19505,N_19162);
nor UO_2234 (O_2234,N_19606,N_19779);
or UO_2235 (O_2235,N_19341,N_19332);
nand UO_2236 (O_2236,N_19697,N_19602);
or UO_2237 (O_2237,N_19204,N_19823);
nor UO_2238 (O_2238,N_19533,N_19717);
nor UO_2239 (O_2239,N_19692,N_19272);
xor UO_2240 (O_2240,N_19764,N_19093);
or UO_2241 (O_2241,N_19428,N_19364);
nand UO_2242 (O_2242,N_19385,N_19301);
nor UO_2243 (O_2243,N_19238,N_19741);
or UO_2244 (O_2244,N_19597,N_19665);
xnor UO_2245 (O_2245,N_19024,N_19886);
xor UO_2246 (O_2246,N_19647,N_19629);
nor UO_2247 (O_2247,N_19962,N_19898);
nor UO_2248 (O_2248,N_19570,N_19491);
nor UO_2249 (O_2249,N_19529,N_19578);
xor UO_2250 (O_2250,N_19632,N_19719);
and UO_2251 (O_2251,N_19264,N_19899);
or UO_2252 (O_2252,N_19257,N_19634);
or UO_2253 (O_2253,N_19876,N_19438);
nor UO_2254 (O_2254,N_19637,N_19208);
nand UO_2255 (O_2255,N_19258,N_19848);
and UO_2256 (O_2256,N_19073,N_19048);
nand UO_2257 (O_2257,N_19957,N_19004);
and UO_2258 (O_2258,N_19731,N_19248);
and UO_2259 (O_2259,N_19021,N_19347);
or UO_2260 (O_2260,N_19916,N_19364);
xnor UO_2261 (O_2261,N_19209,N_19161);
nand UO_2262 (O_2262,N_19835,N_19152);
xnor UO_2263 (O_2263,N_19510,N_19215);
or UO_2264 (O_2264,N_19659,N_19820);
or UO_2265 (O_2265,N_19605,N_19153);
nor UO_2266 (O_2266,N_19848,N_19511);
nor UO_2267 (O_2267,N_19529,N_19713);
and UO_2268 (O_2268,N_19701,N_19343);
nand UO_2269 (O_2269,N_19562,N_19645);
and UO_2270 (O_2270,N_19981,N_19429);
and UO_2271 (O_2271,N_19809,N_19239);
or UO_2272 (O_2272,N_19041,N_19930);
and UO_2273 (O_2273,N_19599,N_19570);
xor UO_2274 (O_2274,N_19120,N_19673);
nand UO_2275 (O_2275,N_19256,N_19808);
nor UO_2276 (O_2276,N_19617,N_19864);
nor UO_2277 (O_2277,N_19713,N_19283);
nand UO_2278 (O_2278,N_19892,N_19762);
nor UO_2279 (O_2279,N_19229,N_19923);
xor UO_2280 (O_2280,N_19010,N_19360);
and UO_2281 (O_2281,N_19029,N_19652);
or UO_2282 (O_2282,N_19397,N_19573);
nand UO_2283 (O_2283,N_19955,N_19618);
or UO_2284 (O_2284,N_19908,N_19939);
and UO_2285 (O_2285,N_19161,N_19494);
nand UO_2286 (O_2286,N_19629,N_19208);
nand UO_2287 (O_2287,N_19242,N_19244);
nor UO_2288 (O_2288,N_19950,N_19601);
nor UO_2289 (O_2289,N_19733,N_19541);
and UO_2290 (O_2290,N_19400,N_19915);
or UO_2291 (O_2291,N_19671,N_19416);
and UO_2292 (O_2292,N_19147,N_19911);
nand UO_2293 (O_2293,N_19898,N_19308);
nand UO_2294 (O_2294,N_19148,N_19219);
xnor UO_2295 (O_2295,N_19697,N_19128);
or UO_2296 (O_2296,N_19105,N_19009);
and UO_2297 (O_2297,N_19692,N_19499);
nor UO_2298 (O_2298,N_19492,N_19754);
and UO_2299 (O_2299,N_19525,N_19164);
xor UO_2300 (O_2300,N_19108,N_19579);
or UO_2301 (O_2301,N_19659,N_19353);
or UO_2302 (O_2302,N_19585,N_19655);
xor UO_2303 (O_2303,N_19230,N_19359);
xnor UO_2304 (O_2304,N_19184,N_19143);
nand UO_2305 (O_2305,N_19439,N_19564);
xnor UO_2306 (O_2306,N_19820,N_19786);
and UO_2307 (O_2307,N_19331,N_19322);
xnor UO_2308 (O_2308,N_19234,N_19590);
and UO_2309 (O_2309,N_19171,N_19812);
and UO_2310 (O_2310,N_19297,N_19895);
and UO_2311 (O_2311,N_19985,N_19276);
or UO_2312 (O_2312,N_19598,N_19218);
xor UO_2313 (O_2313,N_19166,N_19384);
nor UO_2314 (O_2314,N_19063,N_19978);
or UO_2315 (O_2315,N_19761,N_19220);
or UO_2316 (O_2316,N_19428,N_19779);
or UO_2317 (O_2317,N_19263,N_19969);
nor UO_2318 (O_2318,N_19330,N_19871);
nor UO_2319 (O_2319,N_19148,N_19660);
or UO_2320 (O_2320,N_19744,N_19836);
nand UO_2321 (O_2321,N_19866,N_19475);
or UO_2322 (O_2322,N_19767,N_19086);
nand UO_2323 (O_2323,N_19484,N_19824);
nand UO_2324 (O_2324,N_19267,N_19770);
nand UO_2325 (O_2325,N_19811,N_19621);
xor UO_2326 (O_2326,N_19115,N_19626);
and UO_2327 (O_2327,N_19279,N_19567);
and UO_2328 (O_2328,N_19775,N_19992);
nor UO_2329 (O_2329,N_19953,N_19708);
nor UO_2330 (O_2330,N_19362,N_19726);
or UO_2331 (O_2331,N_19304,N_19193);
nor UO_2332 (O_2332,N_19935,N_19454);
or UO_2333 (O_2333,N_19718,N_19412);
xor UO_2334 (O_2334,N_19068,N_19010);
or UO_2335 (O_2335,N_19314,N_19096);
xor UO_2336 (O_2336,N_19160,N_19614);
or UO_2337 (O_2337,N_19161,N_19572);
and UO_2338 (O_2338,N_19674,N_19724);
or UO_2339 (O_2339,N_19877,N_19647);
nor UO_2340 (O_2340,N_19039,N_19890);
or UO_2341 (O_2341,N_19063,N_19138);
and UO_2342 (O_2342,N_19131,N_19578);
xnor UO_2343 (O_2343,N_19974,N_19707);
or UO_2344 (O_2344,N_19974,N_19942);
or UO_2345 (O_2345,N_19952,N_19291);
nand UO_2346 (O_2346,N_19756,N_19496);
or UO_2347 (O_2347,N_19648,N_19119);
nor UO_2348 (O_2348,N_19501,N_19014);
or UO_2349 (O_2349,N_19547,N_19600);
nor UO_2350 (O_2350,N_19720,N_19379);
nor UO_2351 (O_2351,N_19170,N_19212);
and UO_2352 (O_2352,N_19438,N_19203);
nand UO_2353 (O_2353,N_19424,N_19217);
nand UO_2354 (O_2354,N_19977,N_19161);
or UO_2355 (O_2355,N_19041,N_19372);
nor UO_2356 (O_2356,N_19978,N_19389);
or UO_2357 (O_2357,N_19273,N_19293);
or UO_2358 (O_2358,N_19088,N_19924);
or UO_2359 (O_2359,N_19313,N_19720);
xnor UO_2360 (O_2360,N_19544,N_19683);
nand UO_2361 (O_2361,N_19207,N_19942);
or UO_2362 (O_2362,N_19359,N_19627);
nor UO_2363 (O_2363,N_19445,N_19308);
nand UO_2364 (O_2364,N_19044,N_19361);
and UO_2365 (O_2365,N_19943,N_19051);
and UO_2366 (O_2366,N_19513,N_19976);
nand UO_2367 (O_2367,N_19316,N_19088);
and UO_2368 (O_2368,N_19488,N_19784);
or UO_2369 (O_2369,N_19841,N_19507);
or UO_2370 (O_2370,N_19589,N_19492);
and UO_2371 (O_2371,N_19237,N_19018);
xnor UO_2372 (O_2372,N_19227,N_19488);
and UO_2373 (O_2373,N_19135,N_19513);
and UO_2374 (O_2374,N_19726,N_19317);
or UO_2375 (O_2375,N_19058,N_19652);
or UO_2376 (O_2376,N_19647,N_19652);
xor UO_2377 (O_2377,N_19895,N_19723);
xnor UO_2378 (O_2378,N_19492,N_19632);
nor UO_2379 (O_2379,N_19039,N_19924);
nor UO_2380 (O_2380,N_19152,N_19547);
or UO_2381 (O_2381,N_19057,N_19906);
and UO_2382 (O_2382,N_19111,N_19364);
and UO_2383 (O_2383,N_19732,N_19523);
and UO_2384 (O_2384,N_19676,N_19931);
nor UO_2385 (O_2385,N_19483,N_19370);
nand UO_2386 (O_2386,N_19128,N_19687);
or UO_2387 (O_2387,N_19513,N_19523);
nor UO_2388 (O_2388,N_19808,N_19157);
and UO_2389 (O_2389,N_19918,N_19606);
and UO_2390 (O_2390,N_19095,N_19939);
and UO_2391 (O_2391,N_19326,N_19034);
nand UO_2392 (O_2392,N_19825,N_19812);
xor UO_2393 (O_2393,N_19574,N_19849);
xor UO_2394 (O_2394,N_19445,N_19029);
and UO_2395 (O_2395,N_19567,N_19813);
nor UO_2396 (O_2396,N_19365,N_19455);
and UO_2397 (O_2397,N_19998,N_19915);
and UO_2398 (O_2398,N_19987,N_19336);
or UO_2399 (O_2399,N_19884,N_19623);
nor UO_2400 (O_2400,N_19144,N_19208);
xnor UO_2401 (O_2401,N_19321,N_19825);
and UO_2402 (O_2402,N_19215,N_19987);
nand UO_2403 (O_2403,N_19391,N_19329);
nor UO_2404 (O_2404,N_19921,N_19066);
and UO_2405 (O_2405,N_19829,N_19710);
and UO_2406 (O_2406,N_19112,N_19741);
nor UO_2407 (O_2407,N_19965,N_19345);
and UO_2408 (O_2408,N_19135,N_19321);
nand UO_2409 (O_2409,N_19013,N_19292);
and UO_2410 (O_2410,N_19882,N_19619);
nand UO_2411 (O_2411,N_19688,N_19729);
and UO_2412 (O_2412,N_19776,N_19129);
and UO_2413 (O_2413,N_19935,N_19716);
or UO_2414 (O_2414,N_19714,N_19323);
nor UO_2415 (O_2415,N_19926,N_19457);
and UO_2416 (O_2416,N_19038,N_19056);
nor UO_2417 (O_2417,N_19034,N_19558);
and UO_2418 (O_2418,N_19270,N_19862);
or UO_2419 (O_2419,N_19500,N_19042);
xor UO_2420 (O_2420,N_19692,N_19559);
xor UO_2421 (O_2421,N_19099,N_19346);
nor UO_2422 (O_2422,N_19060,N_19463);
nor UO_2423 (O_2423,N_19504,N_19045);
nor UO_2424 (O_2424,N_19070,N_19080);
and UO_2425 (O_2425,N_19806,N_19238);
and UO_2426 (O_2426,N_19502,N_19714);
nor UO_2427 (O_2427,N_19615,N_19425);
and UO_2428 (O_2428,N_19638,N_19288);
or UO_2429 (O_2429,N_19261,N_19953);
nand UO_2430 (O_2430,N_19002,N_19702);
nor UO_2431 (O_2431,N_19777,N_19926);
xnor UO_2432 (O_2432,N_19136,N_19738);
nand UO_2433 (O_2433,N_19021,N_19998);
or UO_2434 (O_2434,N_19361,N_19788);
nor UO_2435 (O_2435,N_19241,N_19215);
xnor UO_2436 (O_2436,N_19136,N_19815);
xor UO_2437 (O_2437,N_19888,N_19004);
or UO_2438 (O_2438,N_19518,N_19860);
xor UO_2439 (O_2439,N_19097,N_19502);
and UO_2440 (O_2440,N_19759,N_19047);
or UO_2441 (O_2441,N_19018,N_19144);
xor UO_2442 (O_2442,N_19656,N_19096);
xnor UO_2443 (O_2443,N_19026,N_19936);
and UO_2444 (O_2444,N_19629,N_19660);
xnor UO_2445 (O_2445,N_19285,N_19719);
or UO_2446 (O_2446,N_19378,N_19143);
nand UO_2447 (O_2447,N_19888,N_19741);
and UO_2448 (O_2448,N_19602,N_19358);
xnor UO_2449 (O_2449,N_19269,N_19519);
and UO_2450 (O_2450,N_19995,N_19105);
and UO_2451 (O_2451,N_19455,N_19668);
or UO_2452 (O_2452,N_19255,N_19829);
xnor UO_2453 (O_2453,N_19251,N_19784);
and UO_2454 (O_2454,N_19804,N_19546);
nor UO_2455 (O_2455,N_19642,N_19156);
xor UO_2456 (O_2456,N_19768,N_19549);
nor UO_2457 (O_2457,N_19055,N_19266);
nor UO_2458 (O_2458,N_19165,N_19914);
xnor UO_2459 (O_2459,N_19465,N_19765);
and UO_2460 (O_2460,N_19532,N_19429);
xnor UO_2461 (O_2461,N_19069,N_19091);
nand UO_2462 (O_2462,N_19016,N_19580);
and UO_2463 (O_2463,N_19845,N_19893);
and UO_2464 (O_2464,N_19568,N_19075);
nand UO_2465 (O_2465,N_19664,N_19837);
nor UO_2466 (O_2466,N_19876,N_19541);
or UO_2467 (O_2467,N_19577,N_19672);
nand UO_2468 (O_2468,N_19933,N_19953);
nor UO_2469 (O_2469,N_19195,N_19832);
and UO_2470 (O_2470,N_19982,N_19778);
nand UO_2471 (O_2471,N_19303,N_19865);
nor UO_2472 (O_2472,N_19228,N_19510);
nand UO_2473 (O_2473,N_19032,N_19544);
and UO_2474 (O_2474,N_19674,N_19094);
and UO_2475 (O_2475,N_19358,N_19208);
nand UO_2476 (O_2476,N_19199,N_19065);
or UO_2477 (O_2477,N_19170,N_19187);
nand UO_2478 (O_2478,N_19375,N_19400);
xnor UO_2479 (O_2479,N_19502,N_19908);
nor UO_2480 (O_2480,N_19914,N_19052);
xnor UO_2481 (O_2481,N_19658,N_19878);
or UO_2482 (O_2482,N_19771,N_19901);
nand UO_2483 (O_2483,N_19790,N_19382);
xnor UO_2484 (O_2484,N_19326,N_19741);
nand UO_2485 (O_2485,N_19203,N_19824);
xor UO_2486 (O_2486,N_19614,N_19418);
or UO_2487 (O_2487,N_19023,N_19212);
and UO_2488 (O_2488,N_19149,N_19888);
nand UO_2489 (O_2489,N_19824,N_19246);
nor UO_2490 (O_2490,N_19125,N_19292);
xor UO_2491 (O_2491,N_19397,N_19000);
and UO_2492 (O_2492,N_19663,N_19695);
xnor UO_2493 (O_2493,N_19537,N_19574);
xnor UO_2494 (O_2494,N_19329,N_19959);
or UO_2495 (O_2495,N_19329,N_19468);
xnor UO_2496 (O_2496,N_19394,N_19545);
nor UO_2497 (O_2497,N_19688,N_19991);
nor UO_2498 (O_2498,N_19279,N_19266);
nor UO_2499 (O_2499,N_19118,N_19052);
endmodule