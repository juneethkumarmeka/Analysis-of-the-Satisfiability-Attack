module basic_750_5000_1000_10_levels_1xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_301,In_544);
nand U1 (N_1,In_456,In_741);
or U2 (N_2,In_263,In_360);
nand U3 (N_3,In_629,In_672);
nand U4 (N_4,In_114,In_26);
nand U5 (N_5,In_261,In_661);
nand U6 (N_6,In_275,In_347);
nand U7 (N_7,In_366,In_432);
nand U8 (N_8,In_281,In_521);
or U9 (N_9,In_229,In_706);
or U10 (N_10,In_720,In_119);
and U11 (N_11,In_253,In_108);
nor U12 (N_12,In_440,In_523);
nor U13 (N_13,In_107,In_652);
or U14 (N_14,In_566,In_536);
and U15 (N_15,In_718,In_127);
and U16 (N_16,In_608,In_173);
and U17 (N_17,In_356,In_278);
or U18 (N_18,In_526,In_635);
and U19 (N_19,In_51,In_495);
nand U20 (N_20,In_726,In_65);
and U21 (N_21,In_244,In_176);
nor U22 (N_22,In_262,In_300);
nor U23 (N_23,In_742,In_739);
or U24 (N_24,In_654,In_567);
nor U25 (N_25,In_601,In_381);
or U26 (N_26,In_509,In_397);
or U27 (N_27,In_141,In_585);
and U28 (N_28,In_591,In_78);
and U29 (N_29,In_604,In_731);
or U30 (N_30,In_136,In_451);
or U31 (N_31,In_371,In_27);
nand U32 (N_32,In_687,In_401);
or U33 (N_33,In_427,In_286);
nor U34 (N_34,In_285,In_236);
or U35 (N_35,In_148,In_677);
nor U36 (N_36,In_363,In_660);
nor U37 (N_37,In_387,In_396);
nor U38 (N_38,In_35,In_369);
or U39 (N_39,In_250,In_69);
nand U40 (N_40,In_355,In_237);
and U41 (N_41,In_210,In_727);
nor U42 (N_42,In_129,In_159);
nor U43 (N_43,In_606,In_496);
nor U44 (N_44,In_53,In_499);
nand U45 (N_45,In_10,In_180);
nand U46 (N_46,In_191,In_149);
or U47 (N_47,In_106,In_354);
nor U48 (N_48,In_510,In_703);
nor U49 (N_49,In_577,In_242);
or U50 (N_50,In_166,In_623);
and U51 (N_51,In_374,In_597);
nand U52 (N_52,In_227,In_241);
and U53 (N_53,In_575,In_543);
nand U54 (N_54,In_336,In_418);
or U55 (N_55,In_505,In_125);
nand U56 (N_56,In_16,In_143);
nor U57 (N_57,In_452,In_330);
and U58 (N_58,In_444,In_639);
and U59 (N_59,In_458,In_232);
nand U60 (N_60,In_368,In_52);
nand U61 (N_61,In_18,In_67);
and U62 (N_62,In_200,In_137);
nand U63 (N_63,In_316,In_193);
or U64 (N_64,In_408,In_490);
nor U65 (N_65,In_247,In_353);
or U66 (N_66,In_676,In_359);
and U67 (N_67,In_269,In_192);
or U68 (N_68,In_344,In_625);
or U69 (N_69,In_728,In_744);
and U70 (N_70,In_76,In_416);
and U71 (N_71,In_637,In_423);
or U72 (N_72,In_383,In_178);
and U73 (N_73,In_649,In_158);
and U74 (N_74,In_134,In_667);
or U75 (N_75,In_556,In_626);
and U76 (N_76,In_583,In_25);
and U77 (N_77,In_708,In_573);
nor U78 (N_78,In_209,In_102);
nor U79 (N_79,In_712,In_633);
and U80 (N_80,In_645,In_346);
or U81 (N_81,In_19,In_562);
nor U82 (N_82,In_404,In_364);
nor U83 (N_83,In_607,In_235);
or U84 (N_84,In_707,In_735);
or U85 (N_85,In_584,In_75);
and U86 (N_86,In_553,In_375);
or U87 (N_87,In_502,In_61);
nand U88 (N_88,In_373,In_335);
nand U89 (N_89,In_181,In_698);
nor U90 (N_90,In_699,In_124);
or U91 (N_91,In_714,In_14);
or U92 (N_92,In_477,In_647);
and U93 (N_93,In_59,In_489);
and U94 (N_94,In_399,In_678);
nand U95 (N_95,In_504,In_131);
nor U96 (N_96,In_329,In_17);
nor U97 (N_97,In_132,In_559);
nand U98 (N_98,In_56,In_341);
and U99 (N_99,In_185,In_391);
or U100 (N_100,In_196,In_308);
and U101 (N_101,In_436,In_737);
and U102 (N_102,In_221,In_450);
or U103 (N_103,In_81,In_128);
nor U104 (N_104,In_289,In_77);
nor U105 (N_105,In_540,In_86);
and U106 (N_106,In_212,In_282);
or U107 (N_107,In_722,In_94);
nor U108 (N_108,In_385,In_31);
nand U109 (N_109,In_267,In_471);
nor U110 (N_110,In_587,In_251);
or U111 (N_111,In_651,In_157);
or U112 (N_112,In_670,In_88);
nor U113 (N_113,In_484,In_139);
and U114 (N_114,In_411,In_152);
nor U115 (N_115,In_4,In_29);
and U116 (N_116,In_497,In_135);
nor U117 (N_117,In_246,In_457);
nor U118 (N_118,In_474,In_34);
nor U119 (N_119,In_243,In_463);
nand U120 (N_120,In_288,In_231);
nand U121 (N_121,In_90,In_63);
and U122 (N_122,In_631,In_186);
and U123 (N_123,In_723,In_725);
or U124 (N_124,In_47,In_596);
nand U125 (N_125,In_207,In_367);
and U126 (N_126,In_311,In_564);
xor U127 (N_127,In_546,In_324);
nand U128 (N_128,In_475,In_254);
nand U129 (N_129,In_425,In_203);
nand U130 (N_130,In_362,In_320);
nor U131 (N_131,In_732,In_719);
or U132 (N_132,In_303,In_716);
nor U133 (N_133,In_618,In_350);
or U134 (N_134,In_721,In_296);
and U135 (N_135,In_379,In_555);
nor U136 (N_136,In_694,In_361);
nor U137 (N_137,In_20,In_454);
nor U138 (N_138,In_524,In_542);
nand U139 (N_139,In_511,In_669);
nand U140 (N_140,In_169,In_684);
nand U141 (N_141,In_150,In_225);
nor U142 (N_142,In_24,In_380);
and U143 (N_143,In_713,In_331);
nand U144 (N_144,In_648,In_195);
or U145 (N_145,In_249,In_462);
and U146 (N_146,In_748,In_117);
nand U147 (N_147,In_613,In_478);
or U148 (N_148,In_23,In_747);
nor U149 (N_149,In_163,In_689);
or U150 (N_150,In_120,In_211);
and U151 (N_151,In_668,In_274);
nand U152 (N_152,In_322,In_7);
nor U153 (N_153,In_206,In_460);
or U154 (N_154,In_421,In_435);
and U155 (N_155,In_527,In_268);
or U156 (N_156,In_258,In_663);
and U157 (N_157,In_617,In_1);
nor U158 (N_158,In_146,In_415);
nor U159 (N_159,In_307,In_315);
or U160 (N_160,In_15,In_118);
and U161 (N_161,In_147,In_409);
nor U162 (N_162,In_299,In_32);
nand U163 (N_163,In_54,In_257);
or U164 (N_164,In_529,In_172);
and U165 (N_165,In_434,In_548);
xor U166 (N_166,In_321,In_179);
nand U167 (N_167,In_58,In_390);
nor U168 (N_168,In_85,In_482);
or U169 (N_169,In_73,In_87);
nand U170 (N_170,In_184,In_252);
and U171 (N_171,In_101,In_394);
and U172 (N_172,In_691,In_441);
nor U173 (N_173,In_62,In_522);
nor U174 (N_174,In_170,In_205);
or U175 (N_175,In_80,In_255);
or U176 (N_176,In_386,In_2);
nand U177 (N_177,In_305,In_182);
and U178 (N_178,In_337,In_638);
nand U179 (N_179,In_519,In_64);
or U180 (N_180,In_420,In_412);
and U181 (N_181,In_264,In_154);
or U182 (N_182,In_541,In_686);
nand U183 (N_183,In_658,In_557);
or U184 (N_184,In_574,In_283);
and U185 (N_185,In_402,In_582);
nor U186 (N_186,In_6,In_612);
nand U187 (N_187,In_525,In_217);
nand U188 (N_188,In_164,In_60);
xnor U189 (N_189,In_641,In_160);
and U190 (N_190,In_579,In_410);
or U191 (N_191,In_292,In_593);
or U192 (N_192,In_702,In_318);
and U193 (N_193,In_46,In_438);
and U194 (N_194,In_666,In_594);
nor U195 (N_195,In_675,In_501);
and U196 (N_196,In_483,In_422);
and U197 (N_197,In_219,In_551);
nor U198 (N_198,In_498,In_204);
nor U199 (N_199,In_99,In_21);
nor U200 (N_200,In_578,In_561);
and U201 (N_201,In_50,In_419);
nand U202 (N_202,In_378,In_220);
or U203 (N_203,In_109,In_630);
or U204 (N_204,In_642,In_188);
and U205 (N_205,In_0,In_514);
and U206 (N_206,In_270,In_222);
nor U207 (N_207,In_603,In_294);
and U208 (N_208,In_469,In_620);
nand U209 (N_209,In_605,In_167);
and U210 (N_210,In_38,In_37);
and U211 (N_211,In_377,In_116);
nand U212 (N_212,In_576,In_290);
and U213 (N_213,In_323,In_485);
or U214 (N_214,In_66,In_395);
nand U215 (N_215,In_734,In_388);
and U216 (N_216,In_238,In_121);
nand U217 (N_217,In_466,In_437);
xor U218 (N_218,In_333,In_453);
nor U219 (N_219,In_168,In_89);
nand U220 (N_220,In_230,In_715);
or U221 (N_221,In_39,In_11);
or U222 (N_222,In_738,In_428);
nand U223 (N_223,In_545,In_468);
nand U224 (N_224,In_405,In_650);
nor U225 (N_225,In_424,In_293);
or U226 (N_226,In_486,In_534);
and U227 (N_227,In_479,In_443);
nor U228 (N_228,In_112,In_692);
and U229 (N_229,In_417,In_161);
or U230 (N_230,In_705,In_36);
or U231 (N_231,In_240,In_539);
nor U232 (N_232,In_44,In_165);
nand U233 (N_233,In_621,In_328);
or U234 (N_234,In_600,In_228);
and U235 (N_235,In_201,In_535);
or U236 (N_236,In_190,In_174);
nor U237 (N_237,In_162,In_685);
or U238 (N_238,In_277,In_538);
nor U239 (N_239,In_234,In_736);
or U240 (N_240,In_683,In_515);
nand U241 (N_241,In_358,In_665);
nand U242 (N_242,In_448,In_98);
and U243 (N_243,In_517,In_488);
and U244 (N_244,In_640,In_537);
nand U245 (N_245,In_740,In_572);
or U246 (N_246,In_403,In_704);
and U247 (N_247,In_455,In_215);
nor U248 (N_248,In_558,In_8);
or U249 (N_249,In_273,In_487);
or U250 (N_250,In_9,In_327);
or U251 (N_251,In_97,In_140);
nand U252 (N_252,In_194,In_309);
nand U253 (N_253,In_145,In_233);
or U254 (N_254,In_142,In_110);
or U255 (N_255,In_352,In_426);
and U256 (N_256,In_619,In_295);
and U257 (N_257,In_695,In_508);
nor U258 (N_258,In_357,In_96);
nor U259 (N_259,In_133,In_690);
nor U260 (N_260,In_198,In_334);
nor U261 (N_261,In_653,In_503);
and U262 (N_262,In_376,In_338);
or U263 (N_263,In_343,In_512);
nor U264 (N_264,In_400,In_459);
nor U265 (N_265,In_155,In_68);
or U266 (N_266,In_272,In_319);
nand U267 (N_267,In_616,In_465);
nor U268 (N_268,In_610,In_298);
and U269 (N_269,In_644,In_664);
nand U270 (N_270,In_563,In_105);
nand U271 (N_271,In_595,In_446);
nand U272 (N_272,In_100,In_467);
or U273 (N_273,In_122,In_287);
or U274 (N_274,In_680,In_554);
or U275 (N_275,In_144,In_589);
nand U276 (N_276,In_22,In_40);
nor U277 (N_277,In_547,In_79);
nand U278 (N_278,In_472,In_276);
nor U279 (N_279,In_393,In_332);
nor U280 (N_280,In_349,In_592);
or U281 (N_281,In_549,In_673);
or U282 (N_282,In_614,In_156);
and U283 (N_283,In_491,In_746);
nor U284 (N_284,In_565,In_431);
or U285 (N_285,In_183,In_43);
nor U286 (N_286,In_473,In_588);
nor U287 (N_287,In_113,In_216);
and U288 (N_288,In_3,In_516);
nand U289 (N_289,In_724,In_126);
or U290 (N_290,In_239,In_560);
nand U291 (N_291,In_681,In_72);
or U292 (N_292,In_636,In_743);
nand U293 (N_293,In_384,In_370);
nor U294 (N_294,In_55,In_213);
nor U295 (N_295,In_84,In_115);
nand U296 (N_296,In_581,In_710);
nor U297 (N_297,In_33,In_571);
nand U298 (N_298,In_314,In_260);
nand U299 (N_299,In_317,In_730);
or U300 (N_300,In_226,In_745);
or U301 (N_301,In_749,In_123);
nor U302 (N_302,In_701,In_95);
nor U303 (N_303,In_634,In_284);
nor U304 (N_304,In_82,In_655);
nor U305 (N_305,In_500,In_13);
nor U306 (N_306,In_439,In_414);
nand U307 (N_307,In_30,In_580);
nor U308 (N_308,In_104,In_461);
or U309 (N_309,In_494,In_83);
nand U310 (N_310,In_513,In_530);
nand U311 (N_311,In_93,In_70);
nand U312 (N_312,In_177,In_313);
nor U313 (N_313,In_492,In_709);
nand U314 (N_314,In_507,In_12);
or U315 (N_315,In_442,In_696);
nor U316 (N_316,In_248,In_493);
or U317 (N_317,In_602,In_326);
nor U318 (N_318,In_189,In_632);
nor U319 (N_319,In_297,In_175);
or U320 (N_320,In_339,In_306);
and U321 (N_321,In_615,In_611);
or U322 (N_322,In_91,In_656);
and U323 (N_323,In_48,In_506);
nand U324 (N_324,In_348,In_449);
and U325 (N_325,In_711,In_624);
or U326 (N_326,In_340,In_671);
nand U327 (N_327,In_717,In_700);
nand U328 (N_328,In_533,In_41);
nor U329 (N_329,In_280,In_71);
and U330 (N_330,In_697,In_345);
or U331 (N_331,In_659,In_187);
nand U332 (N_332,In_291,In_429);
and U333 (N_333,In_679,In_568);
nand U334 (N_334,In_407,In_218);
and U335 (N_335,In_528,In_325);
or U336 (N_336,In_627,In_476);
or U337 (N_337,In_413,In_481);
nand U338 (N_338,In_733,In_312);
nor U339 (N_339,In_49,In_74);
or U340 (N_340,In_271,In_406);
and U341 (N_341,In_365,In_202);
and U342 (N_342,In_130,In_256);
and U343 (N_343,In_430,In_279);
or U344 (N_344,In_433,In_266);
and U345 (N_345,In_138,In_197);
nand U346 (N_346,In_57,In_304);
or U347 (N_347,In_214,In_398);
nor U348 (N_348,In_342,In_447);
and U349 (N_349,In_445,In_171);
nand U350 (N_350,In_729,In_92);
and U351 (N_351,In_351,In_464);
nand U352 (N_352,In_392,In_657);
nand U353 (N_353,In_28,In_372);
or U354 (N_354,In_693,In_310);
or U355 (N_355,In_532,In_245);
and U356 (N_356,In_674,In_688);
or U357 (N_357,In_5,In_151);
or U358 (N_358,In_382,In_682);
or U359 (N_359,In_111,In_531);
and U360 (N_360,In_598,In_153);
nor U361 (N_361,In_42,In_622);
and U362 (N_362,In_662,In_45);
and U363 (N_363,In_552,In_646);
nand U364 (N_364,In_518,In_599);
or U365 (N_365,In_569,In_103);
nor U366 (N_366,In_550,In_223);
nor U367 (N_367,In_480,In_609);
and U368 (N_368,In_470,In_259);
or U369 (N_369,In_520,In_389);
or U370 (N_370,In_628,In_265);
or U371 (N_371,In_199,In_570);
or U372 (N_372,In_586,In_590);
nand U373 (N_373,In_224,In_208);
nand U374 (N_374,In_643,In_302);
or U375 (N_375,In_379,In_338);
or U376 (N_376,In_1,In_631);
nor U377 (N_377,In_65,In_43);
and U378 (N_378,In_219,In_444);
or U379 (N_379,In_568,In_282);
and U380 (N_380,In_591,In_272);
and U381 (N_381,In_481,In_668);
or U382 (N_382,In_613,In_575);
nor U383 (N_383,In_726,In_584);
nor U384 (N_384,In_631,In_651);
nor U385 (N_385,In_264,In_28);
nand U386 (N_386,In_270,In_17);
or U387 (N_387,In_381,In_75);
nor U388 (N_388,In_204,In_620);
nor U389 (N_389,In_695,In_341);
and U390 (N_390,In_23,In_228);
or U391 (N_391,In_238,In_537);
or U392 (N_392,In_448,In_146);
nand U393 (N_393,In_187,In_113);
or U394 (N_394,In_180,In_238);
nor U395 (N_395,In_16,In_472);
nor U396 (N_396,In_154,In_340);
and U397 (N_397,In_737,In_42);
nand U398 (N_398,In_554,In_74);
nand U399 (N_399,In_377,In_304);
or U400 (N_400,In_592,In_689);
or U401 (N_401,In_611,In_162);
and U402 (N_402,In_699,In_515);
nand U403 (N_403,In_202,In_669);
nor U404 (N_404,In_573,In_55);
nor U405 (N_405,In_504,In_222);
nor U406 (N_406,In_538,In_711);
and U407 (N_407,In_29,In_188);
or U408 (N_408,In_637,In_512);
nand U409 (N_409,In_433,In_85);
and U410 (N_410,In_437,In_717);
or U411 (N_411,In_202,In_738);
and U412 (N_412,In_360,In_256);
nor U413 (N_413,In_232,In_514);
xor U414 (N_414,In_632,In_215);
or U415 (N_415,In_474,In_273);
nor U416 (N_416,In_552,In_370);
or U417 (N_417,In_325,In_203);
nand U418 (N_418,In_152,In_283);
nor U419 (N_419,In_145,In_326);
nand U420 (N_420,In_249,In_48);
or U421 (N_421,In_424,In_56);
and U422 (N_422,In_385,In_114);
nor U423 (N_423,In_428,In_739);
or U424 (N_424,In_462,In_476);
nand U425 (N_425,In_340,In_582);
nand U426 (N_426,In_436,In_152);
nor U427 (N_427,In_538,In_653);
nor U428 (N_428,In_474,In_2);
and U429 (N_429,In_637,In_316);
nor U430 (N_430,In_729,In_149);
nor U431 (N_431,In_591,In_714);
nand U432 (N_432,In_102,In_46);
and U433 (N_433,In_157,In_460);
nand U434 (N_434,In_452,In_26);
nand U435 (N_435,In_628,In_303);
and U436 (N_436,In_250,In_371);
nor U437 (N_437,In_275,In_400);
or U438 (N_438,In_491,In_105);
nand U439 (N_439,In_64,In_521);
and U440 (N_440,In_109,In_261);
nor U441 (N_441,In_448,In_211);
nand U442 (N_442,In_358,In_568);
and U443 (N_443,In_388,In_314);
nor U444 (N_444,In_446,In_159);
nor U445 (N_445,In_236,In_731);
xor U446 (N_446,In_381,In_632);
nand U447 (N_447,In_541,In_385);
xnor U448 (N_448,In_336,In_98);
or U449 (N_449,In_651,In_315);
nor U450 (N_450,In_234,In_542);
and U451 (N_451,In_35,In_203);
nor U452 (N_452,In_206,In_101);
and U453 (N_453,In_357,In_84);
nand U454 (N_454,In_620,In_180);
and U455 (N_455,In_160,In_192);
and U456 (N_456,In_39,In_457);
nor U457 (N_457,In_113,In_582);
and U458 (N_458,In_260,In_215);
nor U459 (N_459,In_326,In_514);
or U460 (N_460,In_637,In_87);
and U461 (N_461,In_278,In_395);
and U462 (N_462,In_418,In_68);
and U463 (N_463,In_624,In_177);
or U464 (N_464,In_318,In_292);
nor U465 (N_465,In_574,In_35);
nor U466 (N_466,In_612,In_153);
or U467 (N_467,In_733,In_617);
nor U468 (N_468,In_586,In_644);
nor U469 (N_469,In_203,In_629);
nand U470 (N_470,In_451,In_662);
nand U471 (N_471,In_445,In_367);
nor U472 (N_472,In_47,In_484);
and U473 (N_473,In_18,In_373);
nor U474 (N_474,In_557,In_573);
or U475 (N_475,In_325,In_360);
nand U476 (N_476,In_6,In_445);
nand U477 (N_477,In_691,In_186);
nand U478 (N_478,In_144,In_665);
or U479 (N_479,In_527,In_629);
and U480 (N_480,In_710,In_4);
and U481 (N_481,In_629,In_666);
and U482 (N_482,In_477,In_636);
and U483 (N_483,In_462,In_253);
and U484 (N_484,In_4,In_1);
nand U485 (N_485,In_593,In_482);
and U486 (N_486,In_355,In_41);
nand U487 (N_487,In_500,In_656);
nand U488 (N_488,In_258,In_714);
nand U489 (N_489,In_338,In_585);
nor U490 (N_490,In_220,In_152);
nand U491 (N_491,In_376,In_593);
nand U492 (N_492,In_129,In_462);
nand U493 (N_493,In_703,In_220);
and U494 (N_494,In_619,In_134);
and U495 (N_495,In_613,In_711);
nor U496 (N_496,In_261,In_486);
or U497 (N_497,In_365,In_145);
and U498 (N_498,In_609,In_562);
and U499 (N_499,In_18,In_599);
or U500 (N_500,N_408,N_428);
and U501 (N_501,N_491,N_136);
nand U502 (N_502,N_38,N_268);
nand U503 (N_503,N_169,N_272);
nand U504 (N_504,N_165,N_267);
nand U505 (N_505,N_24,N_190);
nand U506 (N_506,N_243,N_79);
nand U507 (N_507,N_45,N_201);
nand U508 (N_508,N_343,N_295);
nor U509 (N_509,N_19,N_4);
or U510 (N_510,N_188,N_320);
or U511 (N_511,N_83,N_13);
nand U512 (N_512,N_328,N_393);
nor U513 (N_513,N_202,N_396);
or U514 (N_514,N_126,N_447);
nor U515 (N_515,N_325,N_60);
and U516 (N_516,N_367,N_218);
or U517 (N_517,N_234,N_253);
nor U518 (N_518,N_392,N_99);
nand U519 (N_519,N_239,N_336);
or U520 (N_520,N_465,N_266);
and U521 (N_521,N_6,N_462);
or U522 (N_522,N_59,N_249);
or U523 (N_523,N_379,N_170);
xnor U524 (N_524,N_252,N_35);
and U525 (N_525,N_488,N_296);
nor U526 (N_526,N_362,N_457);
nor U527 (N_527,N_432,N_85);
and U528 (N_528,N_459,N_208);
or U529 (N_529,N_193,N_482);
or U530 (N_530,N_317,N_134);
nand U531 (N_531,N_414,N_105);
and U532 (N_532,N_300,N_191);
nand U533 (N_533,N_387,N_36);
and U534 (N_534,N_271,N_65);
nand U535 (N_535,N_196,N_365);
and U536 (N_536,N_384,N_9);
or U537 (N_537,N_235,N_141);
nand U538 (N_538,N_102,N_291);
nor U539 (N_539,N_437,N_489);
nand U540 (N_540,N_331,N_70);
nand U541 (N_541,N_486,N_94);
nor U542 (N_542,N_119,N_163);
or U543 (N_543,N_440,N_12);
nand U544 (N_544,N_419,N_460);
and U545 (N_545,N_430,N_363);
nand U546 (N_546,N_138,N_400);
nor U547 (N_547,N_114,N_356);
and U548 (N_548,N_237,N_499);
nand U549 (N_549,N_158,N_251);
nand U550 (N_550,N_27,N_472);
nor U551 (N_551,N_55,N_391);
or U552 (N_552,N_127,N_276);
and U553 (N_553,N_52,N_452);
and U554 (N_554,N_51,N_497);
or U555 (N_555,N_405,N_468);
or U556 (N_556,N_28,N_474);
and U557 (N_557,N_184,N_471);
nand U558 (N_558,N_418,N_33);
nor U559 (N_559,N_179,N_464);
nor U560 (N_560,N_205,N_197);
or U561 (N_561,N_410,N_42);
nand U562 (N_562,N_398,N_492);
or U563 (N_563,N_444,N_135);
and U564 (N_564,N_376,N_153);
or U565 (N_565,N_370,N_92);
nand U566 (N_566,N_228,N_72);
or U567 (N_567,N_340,N_454);
nor U568 (N_568,N_290,N_349);
and U569 (N_569,N_137,N_441);
and U570 (N_570,N_443,N_394);
nor U571 (N_571,N_490,N_411);
or U572 (N_572,N_409,N_233);
or U573 (N_573,N_181,N_48);
and U574 (N_574,N_200,N_95);
nand U575 (N_575,N_15,N_285);
nor U576 (N_576,N_373,N_86);
and U577 (N_577,N_351,N_421);
or U578 (N_578,N_260,N_395);
nor U579 (N_579,N_309,N_159);
or U580 (N_580,N_401,N_467);
and U581 (N_581,N_46,N_355);
and U582 (N_582,N_292,N_280);
nor U583 (N_583,N_265,N_226);
and U584 (N_584,N_319,N_299);
and U585 (N_585,N_195,N_417);
nand U586 (N_586,N_483,N_90);
and U587 (N_587,N_18,N_415);
and U588 (N_588,N_154,N_286);
nor U589 (N_589,N_186,N_133);
nand U590 (N_590,N_298,N_223);
nor U591 (N_591,N_240,N_63);
nor U592 (N_592,N_487,N_87);
nor U593 (N_593,N_183,N_287);
nand U594 (N_594,N_366,N_54);
and U595 (N_595,N_470,N_232);
nor U596 (N_596,N_278,N_446);
or U597 (N_597,N_273,N_323);
and U598 (N_598,N_423,N_167);
and U599 (N_599,N_270,N_162);
or U600 (N_600,N_26,N_56);
or U601 (N_601,N_20,N_361);
or U602 (N_602,N_43,N_106);
and U603 (N_603,N_213,N_485);
and U604 (N_604,N_88,N_407);
nor U605 (N_605,N_142,N_120);
nand U606 (N_606,N_216,N_147);
nor U607 (N_607,N_314,N_310);
nor U608 (N_608,N_157,N_144);
and U609 (N_609,N_8,N_279);
and U610 (N_610,N_269,N_368);
and U611 (N_611,N_112,N_413);
nor U612 (N_612,N_123,N_412);
nand U613 (N_613,N_178,N_227);
nand U614 (N_614,N_283,N_466);
nand U615 (N_615,N_306,N_282);
nand U616 (N_616,N_455,N_185);
nand U617 (N_617,N_161,N_212);
or U618 (N_618,N_281,N_44);
or U619 (N_619,N_143,N_182);
nor U620 (N_620,N_477,N_353);
or U621 (N_621,N_74,N_22);
nand U622 (N_622,N_149,N_187);
nand U623 (N_623,N_372,N_25);
nor U624 (N_624,N_124,N_168);
or U625 (N_625,N_91,N_1);
nand U626 (N_626,N_128,N_364);
or U627 (N_627,N_380,N_493);
nand U628 (N_628,N_288,N_176);
nand U629 (N_629,N_302,N_98);
nand U630 (N_630,N_21,N_132);
and U631 (N_631,N_498,N_57);
nand U632 (N_632,N_342,N_93);
nor U633 (N_633,N_229,N_255);
nor U634 (N_634,N_66,N_164);
and U635 (N_635,N_438,N_104);
or U636 (N_636,N_352,N_427);
and U637 (N_637,N_264,N_82);
and U638 (N_638,N_348,N_5);
nor U639 (N_639,N_62,N_210);
nor U640 (N_640,N_236,N_53);
and U641 (N_641,N_76,N_425);
nand U642 (N_642,N_111,N_301);
nor U643 (N_643,N_166,N_326);
nand U644 (N_644,N_479,N_0);
or U645 (N_645,N_113,N_47);
and U646 (N_646,N_382,N_58);
and U647 (N_647,N_224,N_424);
or U648 (N_648,N_426,N_110);
or U649 (N_649,N_334,N_209);
or U650 (N_650,N_277,N_221);
xnor U651 (N_651,N_304,N_263);
and U652 (N_652,N_450,N_434);
nor U653 (N_653,N_318,N_381);
or U654 (N_654,N_84,N_118);
and U655 (N_655,N_247,N_345);
or U656 (N_656,N_152,N_145);
nand U657 (N_657,N_222,N_330);
and U658 (N_658,N_174,N_431);
or U659 (N_659,N_242,N_344);
or U660 (N_660,N_435,N_89);
nand U661 (N_661,N_420,N_338);
and U662 (N_662,N_49,N_108);
nor U663 (N_663,N_378,N_246);
and U664 (N_664,N_61,N_496);
nor U665 (N_665,N_199,N_316);
nand U666 (N_666,N_347,N_214);
or U667 (N_667,N_449,N_274);
nor U668 (N_668,N_406,N_37);
nor U669 (N_669,N_256,N_121);
nor U670 (N_670,N_100,N_359);
or U671 (N_671,N_203,N_71);
nand U672 (N_672,N_473,N_11);
nand U673 (N_673,N_175,N_386);
or U674 (N_674,N_129,N_475);
or U675 (N_675,N_458,N_225);
nand U676 (N_676,N_397,N_335);
and U677 (N_677,N_375,N_369);
nor U678 (N_678,N_189,N_231);
and U679 (N_679,N_383,N_109);
and U680 (N_680,N_146,N_481);
nand U681 (N_681,N_115,N_321);
nor U682 (N_682,N_461,N_377);
or U683 (N_683,N_103,N_2);
nor U684 (N_684,N_358,N_3);
or U685 (N_685,N_422,N_484);
or U686 (N_686,N_238,N_206);
and U687 (N_687,N_250,N_254);
or U688 (N_688,N_245,N_139);
and U689 (N_689,N_150,N_262);
nand U690 (N_690,N_305,N_148);
or U691 (N_691,N_220,N_404);
and U692 (N_692,N_346,N_360);
or U693 (N_693,N_204,N_389);
or U694 (N_694,N_31,N_211);
xnor U695 (N_695,N_442,N_297);
nand U696 (N_696,N_327,N_34);
nor U697 (N_697,N_308,N_32);
nor U698 (N_698,N_101,N_313);
or U699 (N_699,N_478,N_69);
nor U700 (N_700,N_303,N_388);
nand U701 (N_701,N_171,N_116);
or U702 (N_702,N_311,N_429);
xor U703 (N_703,N_456,N_219);
nand U704 (N_704,N_402,N_131);
nand U705 (N_705,N_289,N_259);
or U706 (N_706,N_230,N_333);
nor U707 (N_707,N_173,N_436);
nor U708 (N_708,N_30,N_341);
or U709 (N_709,N_324,N_374);
nor U710 (N_710,N_453,N_155);
and U711 (N_711,N_17,N_39);
nor U712 (N_712,N_337,N_198);
and U713 (N_713,N_294,N_399);
nand U714 (N_714,N_160,N_385);
and U715 (N_715,N_117,N_322);
nand U716 (N_716,N_469,N_64);
or U717 (N_717,N_258,N_29);
and U718 (N_718,N_107,N_332);
and U719 (N_719,N_329,N_494);
nor U720 (N_720,N_307,N_194);
or U721 (N_721,N_80,N_284);
and U722 (N_722,N_207,N_14);
and U723 (N_723,N_275,N_81);
and U724 (N_724,N_75,N_172);
nand U725 (N_725,N_257,N_215);
nor U726 (N_726,N_217,N_96);
xor U727 (N_727,N_241,N_315);
or U728 (N_728,N_403,N_180);
nor U729 (N_729,N_50,N_41);
nand U730 (N_730,N_151,N_244);
nor U731 (N_731,N_67,N_312);
or U732 (N_732,N_495,N_480);
and U733 (N_733,N_354,N_439);
or U734 (N_734,N_357,N_476);
and U735 (N_735,N_10,N_23);
or U736 (N_736,N_416,N_156);
and U737 (N_737,N_40,N_463);
nand U738 (N_738,N_140,N_77);
and U739 (N_739,N_122,N_451);
and U740 (N_740,N_248,N_293);
and U741 (N_741,N_390,N_371);
nor U742 (N_742,N_339,N_445);
nand U743 (N_743,N_177,N_192);
nand U744 (N_744,N_125,N_448);
nor U745 (N_745,N_97,N_7);
nor U746 (N_746,N_261,N_130);
and U747 (N_747,N_68,N_16);
or U748 (N_748,N_73,N_350);
nand U749 (N_749,N_433,N_78);
and U750 (N_750,N_243,N_404);
nor U751 (N_751,N_473,N_88);
nor U752 (N_752,N_138,N_60);
nand U753 (N_753,N_265,N_416);
nor U754 (N_754,N_8,N_305);
and U755 (N_755,N_425,N_105);
or U756 (N_756,N_441,N_196);
nand U757 (N_757,N_492,N_438);
nand U758 (N_758,N_456,N_205);
nor U759 (N_759,N_92,N_1);
and U760 (N_760,N_265,N_256);
and U761 (N_761,N_48,N_262);
nand U762 (N_762,N_376,N_138);
and U763 (N_763,N_62,N_355);
nor U764 (N_764,N_284,N_398);
or U765 (N_765,N_337,N_203);
nor U766 (N_766,N_89,N_206);
nor U767 (N_767,N_347,N_228);
and U768 (N_768,N_177,N_471);
or U769 (N_769,N_183,N_483);
nand U770 (N_770,N_327,N_241);
nand U771 (N_771,N_203,N_316);
and U772 (N_772,N_55,N_191);
or U773 (N_773,N_309,N_223);
nor U774 (N_774,N_25,N_277);
nand U775 (N_775,N_64,N_372);
nor U776 (N_776,N_103,N_309);
and U777 (N_777,N_408,N_107);
nor U778 (N_778,N_307,N_249);
nand U779 (N_779,N_277,N_28);
and U780 (N_780,N_446,N_181);
or U781 (N_781,N_360,N_320);
or U782 (N_782,N_499,N_433);
nand U783 (N_783,N_453,N_50);
and U784 (N_784,N_360,N_397);
or U785 (N_785,N_437,N_440);
nor U786 (N_786,N_479,N_440);
or U787 (N_787,N_20,N_245);
and U788 (N_788,N_171,N_70);
nor U789 (N_789,N_443,N_94);
and U790 (N_790,N_272,N_424);
nand U791 (N_791,N_128,N_296);
and U792 (N_792,N_435,N_360);
nor U793 (N_793,N_52,N_144);
nor U794 (N_794,N_407,N_344);
nand U795 (N_795,N_111,N_125);
and U796 (N_796,N_131,N_167);
nor U797 (N_797,N_12,N_91);
or U798 (N_798,N_287,N_294);
nor U799 (N_799,N_493,N_452);
and U800 (N_800,N_250,N_466);
nor U801 (N_801,N_15,N_410);
nor U802 (N_802,N_101,N_235);
and U803 (N_803,N_82,N_381);
nand U804 (N_804,N_135,N_204);
nand U805 (N_805,N_443,N_134);
nor U806 (N_806,N_479,N_450);
nand U807 (N_807,N_204,N_111);
nor U808 (N_808,N_421,N_62);
or U809 (N_809,N_450,N_427);
nand U810 (N_810,N_65,N_290);
nor U811 (N_811,N_115,N_28);
or U812 (N_812,N_440,N_434);
nor U813 (N_813,N_469,N_407);
nor U814 (N_814,N_466,N_19);
nor U815 (N_815,N_56,N_470);
nand U816 (N_816,N_358,N_430);
or U817 (N_817,N_88,N_12);
nand U818 (N_818,N_252,N_213);
or U819 (N_819,N_120,N_119);
nand U820 (N_820,N_6,N_360);
nor U821 (N_821,N_215,N_252);
nor U822 (N_822,N_439,N_430);
nor U823 (N_823,N_339,N_1);
or U824 (N_824,N_486,N_480);
nand U825 (N_825,N_336,N_112);
nand U826 (N_826,N_110,N_470);
nand U827 (N_827,N_41,N_24);
nand U828 (N_828,N_414,N_18);
nor U829 (N_829,N_51,N_60);
and U830 (N_830,N_150,N_256);
or U831 (N_831,N_403,N_215);
and U832 (N_832,N_274,N_22);
nand U833 (N_833,N_62,N_180);
and U834 (N_834,N_317,N_251);
nor U835 (N_835,N_497,N_79);
or U836 (N_836,N_125,N_127);
nand U837 (N_837,N_281,N_389);
and U838 (N_838,N_112,N_427);
nand U839 (N_839,N_116,N_408);
and U840 (N_840,N_34,N_317);
nand U841 (N_841,N_181,N_397);
or U842 (N_842,N_355,N_13);
nor U843 (N_843,N_312,N_350);
nand U844 (N_844,N_100,N_95);
nand U845 (N_845,N_194,N_40);
nand U846 (N_846,N_46,N_220);
or U847 (N_847,N_59,N_13);
and U848 (N_848,N_256,N_294);
nand U849 (N_849,N_196,N_26);
nand U850 (N_850,N_200,N_476);
nor U851 (N_851,N_344,N_299);
nor U852 (N_852,N_137,N_214);
and U853 (N_853,N_313,N_71);
and U854 (N_854,N_333,N_46);
xor U855 (N_855,N_398,N_399);
and U856 (N_856,N_348,N_230);
and U857 (N_857,N_245,N_241);
and U858 (N_858,N_117,N_164);
or U859 (N_859,N_242,N_431);
nand U860 (N_860,N_389,N_373);
and U861 (N_861,N_395,N_1);
nor U862 (N_862,N_281,N_403);
nand U863 (N_863,N_397,N_457);
or U864 (N_864,N_178,N_258);
nand U865 (N_865,N_469,N_483);
or U866 (N_866,N_230,N_360);
nand U867 (N_867,N_240,N_2);
nand U868 (N_868,N_403,N_102);
and U869 (N_869,N_344,N_479);
or U870 (N_870,N_319,N_64);
and U871 (N_871,N_309,N_289);
and U872 (N_872,N_55,N_44);
nor U873 (N_873,N_350,N_409);
nor U874 (N_874,N_65,N_50);
nor U875 (N_875,N_323,N_425);
and U876 (N_876,N_132,N_201);
nand U877 (N_877,N_497,N_126);
and U878 (N_878,N_498,N_107);
and U879 (N_879,N_246,N_118);
and U880 (N_880,N_213,N_447);
and U881 (N_881,N_435,N_158);
or U882 (N_882,N_494,N_320);
nor U883 (N_883,N_299,N_433);
and U884 (N_884,N_108,N_281);
or U885 (N_885,N_490,N_37);
or U886 (N_886,N_239,N_92);
nand U887 (N_887,N_213,N_101);
and U888 (N_888,N_165,N_122);
and U889 (N_889,N_27,N_22);
nand U890 (N_890,N_333,N_362);
nor U891 (N_891,N_145,N_1);
and U892 (N_892,N_196,N_112);
nand U893 (N_893,N_283,N_485);
or U894 (N_894,N_121,N_312);
nor U895 (N_895,N_310,N_438);
or U896 (N_896,N_194,N_140);
nand U897 (N_897,N_395,N_267);
or U898 (N_898,N_196,N_141);
or U899 (N_899,N_133,N_75);
nor U900 (N_900,N_483,N_103);
nand U901 (N_901,N_30,N_34);
or U902 (N_902,N_422,N_254);
nand U903 (N_903,N_120,N_327);
or U904 (N_904,N_51,N_271);
and U905 (N_905,N_110,N_53);
nor U906 (N_906,N_240,N_279);
and U907 (N_907,N_61,N_264);
nor U908 (N_908,N_427,N_301);
and U909 (N_909,N_113,N_353);
nand U910 (N_910,N_370,N_88);
nand U911 (N_911,N_1,N_369);
nor U912 (N_912,N_175,N_485);
or U913 (N_913,N_248,N_257);
and U914 (N_914,N_476,N_70);
nor U915 (N_915,N_52,N_217);
and U916 (N_916,N_214,N_405);
and U917 (N_917,N_105,N_447);
nand U918 (N_918,N_322,N_309);
and U919 (N_919,N_425,N_118);
and U920 (N_920,N_463,N_72);
and U921 (N_921,N_84,N_433);
nand U922 (N_922,N_286,N_379);
and U923 (N_923,N_485,N_189);
nor U924 (N_924,N_115,N_338);
nand U925 (N_925,N_390,N_93);
nor U926 (N_926,N_352,N_385);
or U927 (N_927,N_329,N_214);
or U928 (N_928,N_457,N_315);
and U929 (N_929,N_201,N_245);
nand U930 (N_930,N_70,N_124);
and U931 (N_931,N_23,N_415);
or U932 (N_932,N_287,N_444);
nand U933 (N_933,N_232,N_300);
and U934 (N_934,N_354,N_395);
or U935 (N_935,N_176,N_52);
and U936 (N_936,N_484,N_10);
or U937 (N_937,N_406,N_42);
or U938 (N_938,N_358,N_433);
nand U939 (N_939,N_56,N_44);
nand U940 (N_940,N_280,N_120);
nand U941 (N_941,N_195,N_496);
nor U942 (N_942,N_1,N_0);
nor U943 (N_943,N_278,N_361);
nor U944 (N_944,N_326,N_126);
nor U945 (N_945,N_1,N_335);
nor U946 (N_946,N_449,N_331);
xnor U947 (N_947,N_468,N_223);
or U948 (N_948,N_176,N_187);
nand U949 (N_949,N_145,N_440);
nand U950 (N_950,N_493,N_488);
nand U951 (N_951,N_471,N_383);
nand U952 (N_952,N_125,N_245);
or U953 (N_953,N_44,N_352);
or U954 (N_954,N_414,N_296);
or U955 (N_955,N_104,N_358);
nand U956 (N_956,N_318,N_452);
nor U957 (N_957,N_113,N_389);
nand U958 (N_958,N_386,N_302);
or U959 (N_959,N_443,N_423);
nor U960 (N_960,N_53,N_184);
nor U961 (N_961,N_125,N_479);
or U962 (N_962,N_168,N_91);
and U963 (N_963,N_293,N_388);
nand U964 (N_964,N_21,N_311);
and U965 (N_965,N_174,N_22);
or U966 (N_966,N_319,N_397);
nor U967 (N_967,N_125,N_50);
or U968 (N_968,N_285,N_89);
or U969 (N_969,N_176,N_260);
nand U970 (N_970,N_350,N_297);
nand U971 (N_971,N_145,N_449);
nand U972 (N_972,N_218,N_447);
nand U973 (N_973,N_333,N_385);
or U974 (N_974,N_3,N_74);
or U975 (N_975,N_120,N_351);
or U976 (N_976,N_125,N_268);
nand U977 (N_977,N_496,N_248);
nor U978 (N_978,N_214,N_432);
or U979 (N_979,N_311,N_209);
or U980 (N_980,N_287,N_277);
and U981 (N_981,N_75,N_238);
and U982 (N_982,N_233,N_102);
or U983 (N_983,N_304,N_61);
or U984 (N_984,N_205,N_344);
and U985 (N_985,N_68,N_234);
nor U986 (N_986,N_225,N_134);
nor U987 (N_987,N_309,N_449);
or U988 (N_988,N_156,N_129);
nor U989 (N_989,N_215,N_448);
or U990 (N_990,N_406,N_405);
or U991 (N_991,N_400,N_31);
nand U992 (N_992,N_268,N_102);
nand U993 (N_993,N_6,N_50);
nor U994 (N_994,N_367,N_126);
nand U995 (N_995,N_493,N_52);
nand U996 (N_996,N_324,N_385);
or U997 (N_997,N_276,N_389);
nand U998 (N_998,N_142,N_131);
and U999 (N_999,N_353,N_279);
and U1000 (N_1000,N_620,N_956);
or U1001 (N_1001,N_646,N_778);
nor U1002 (N_1002,N_599,N_842);
nor U1003 (N_1003,N_906,N_914);
nand U1004 (N_1004,N_882,N_843);
nor U1005 (N_1005,N_580,N_537);
nand U1006 (N_1006,N_686,N_762);
nand U1007 (N_1007,N_558,N_845);
or U1008 (N_1008,N_589,N_952);
xnor U1009 (N_1009,N_688,N_783);
or U1010 (N_1010,N_868,N_780);
nand U1011 (N_1011,N_940,N_689);
nor U1012 (N_1012,N_941,N_901);
and U1013 (N_1013,N_761,N_534);
and U1014 (N_1014,N_732,N_650);
or U1015 (N_1015,N_706,N_598);
nand U1016 (N_1016,N_705,N_877);
or U1017 (N_1017,N_814,N_570);
or U1018 (N_1018,N_567,N_789);
nor U1019 (N_1019,N_514,N_810);
nor U1020 (N_1020,N_861,N_645);
nand U1021 (N_1021,N_724,N_918);
or U1022 (N_1022,N_700,N_575);
nand U1023 (N_1023,N_963,N_747);
and U1024 (N_1024,N_709,N_798);
nor U1025 (N_1025,N_719,N_727);
nand U1026 (N_1026,N_880,N_750);
nor U1027 (N_1027,N_870,N_751);
and U1028 (N_1028,N_643,N_684);
nor U1029 (N_1029,N_640,N_964);
or U1030 (N_1030,N_765,N_586);
nor U1031 (N_1031,N_653,N_536);
and U1032 (N_1032,N_916,N_636);
or U1033 (N_1033,N_779,N_618);
or U1034 (N_1034,N_505,N_708);
or U1035 (N_1035,N_835,N_950);
or U1036 (N_1036,N_746,N_651);
nor U1037 (N_1037,N_829,N_990);
nor U1038 (N_1038,N_844,N_869);
nand U1039 (N_1039,N_714,N_960);
and U1040 (N_1040,N_953,N_803);
nand U1041 (N_1041,N_891,N_676);
nand U1042 (N_1042,N_763,N_788);
and U1043 (N_1043,N_951,N_931);
nand U1044 (N_1044,N_735,N_879);
and U1045 (N_1045,N_961,N_923);
and U1046 (N_1046,N_697,N_625);
or U1047 (N_1047,N_508,N_629);
or U1048 (N_1048,N_532,N_617);
and U1049 (N_1049,N_926,N_871);
and U1050 (N_1050,N_603,N_939);
or U1051 (N_1051,N_673,N_557);
and U1052 (N_1052,N_704,N_601);
nand U1053 (N_1053,N_602,N_989);
nand U1054 (N_1054,N_973,N_683);
nor U1055 (N_1055,N_635,N_933);
nand U1056 (N_1056,N_693,N_986);
and U1057 (N_1057,N_826,N_595);
nand U1058 (N_1058,N_720,N_573);
nor U1059 (N_1059,N_512,N_822);
or U1060 (N_1060,N_893,N_981);
or U1061 (N_1061,N_616,N_920);
nand U1062 (N_1062,N_942,N_972);
nand U1063 (N_1063,N_959,N_991);
nand U1064 (N_1064,N_787,N_875);
nor U1065 (N_1065,N_540,N_998);
nor U1066 (N_1066,N_506,N_526);
and U1067 (N_1067,N_548,N_626);
or U1068 (N_1068,N_800,N_630);
and U1069 (N_1069,N_621,N_654);
or U1070 (N_1070,N_610,N_976);
or U1071 (N_1071,N_738,N_828);
nor U1072 (N_1072,N_507,N_663);
nand U1073 (N_1073,N_628,N_695);
or U1074 (N_1074,N_587,N_816);
nor U1075 (N_1075,N_503,N_521);
and U1076 (N_1076,N_772,N_921);
nand U1077 (N_1077,N_564,N_569);
nand U1078 (N_1078,N_841,N_757);
nor U1079 (N_1079,N_716,N_588);
and U1080 (N_1080,N_611,N_519);
or U1081 (N_1081,N_895,N_988);
and U1082 (N_1082,N_802,N_922);
nand U1083 (N_1083,N_502,N_755);
and U1084 (N_1084,N_824,N_734);
nor U1085 (N_1085,N_815,N_773);
nor U1086 (N_1086,N_583,N_677);
or U1087 (N_1087,N_739,N_899);
and U1088 (N_1088,N_694,N_766);
nor U1089 (N_1089,N_666,N_885);
nand U1090 (N_1090,N_623,N_550);
or U1091 (N_1091,N_698,N_909);
or U1092 (N_1092,N_662,N_832);
or U1093 (N_1093,N_883,N_966);
and U1094 (N_1094,N_999,N_947);
and U1095 (N_1095,N_552,N_597);
or U1096 (N_1096,N_513,N_632);
nand U1097 (N_1097,N_996,N_690);
nor U1098 (N_1098,N_896,N_937);
nor U1099 (N_1099,N_574,N_744);
and U1100 (N_1100,N_878,N_886);
xnor U1101 (N_1101,N_791,N_553);
nor U1102 (N_1102,N_604,N_555);
xnor U1103 (N_1103,N_556,N_627);
or U1104 (N_1104,N_819,N_992);
nor U1105 (N_1105,N_712,N_946);
or U1106 (N_1106,N_656,N_551);
nand U1107 (N_1107,N_849,N_796);
nand U1108 (N_1108,N_865,N_591);
or U1109 (N_1109,N_915,N_969);
or U1110 (N_1110,N_671,N_544);
nand U1111 (N_1111,N_723,N_807);
and U1112 (N_1112,N_982,N_702);
nor U1113 (N_1113,N_609,N_754);
and U1114 (N_1114,N_774,N_888);
nand U1115 (N_1115,N_812,N_794);
nor U1116 (N_1116,N_582,N_954);
and U1117 (N_1117,N_511,N_839);
nor U1118 (N_1118,N_710,N_864);
and U1119 (N_1119,N_561,N_510);
nand U1120 (N_1120,N_782,N_758);
and U1121 (N_1121,N_631,N_934);
or U1122 (N_1122,N_854,N_806);
nor U1123 (N_1123,N_644,N_993);
nor U1124 (N_1124,N_957,N_935);
and U1125 (N_1125,N_545,N_622);
and U1126 (N_1126,N_892,N_848);
nand U1127 (N_1127,N_890,N_911);
nand U1128 (N_1128,N_995,N_793);
nor U1129 (N_1129,N_905,N_681);
nor U1130 (N_1130,N_549,N_516);
and U1131 (N_1131,N_527,N_847);
nand U1132 (N_1132,N_680,N_563);
and U1133 (N_1133,N_730,N_771);
nor U1134 (N_1134,N_786,N_838);
or U1135 (N_1135,N_713,N_860);
nor U1136 (N_1136,N_980,N_777);
and U1137 (N_1137,N_874,N_731);
and U1138 (N_1138,N_594,N_547);
and U1139 (N_1139,N_531,N_674);
or U1140 (N_1140,N_560,N_924);
nor U1141 (N_1141,N_785,N_997);
nor U1142 (N_1142,N_571,N_975);
and U1143 (N_1143,N_767,N_903);
and U1144 (N_1144,N_678,N_929);
and U1145 (N_1145,N_970,N_585);
or U1146 (N_1146,N_633,N_559);
and U1147 (N_1147,N_614,N_692);
and U1148 (N_1148,N_944,N_866);
nand U1149 (N_1149,N_703,N_760);
nor U1150 (N_1150,N_639,N_978);
nand U1151 (N_1151,N_523,N_768);
nor U1152 (N_1152,N_661,N_820);
nand U1153 (N_1153,N_596,N_930);
and U1154 (N_1154,N_742,N_679);
nor U1155 (N_1155,N_962,N_813);
nor U1156 (N_1156,N_696,N_568);
nor U1157 (N_1157,N_517,N_634);
nor U1158 (N_1158,N_823,N_817);
and U1159 (N_1159,N_799,N_538);
nand U1160 (N_1160,N_675,N_665);
xnor U1161 (N_1161,N_949,N_830);
nor U1162 (N_1162,N_863,N_669);
nor U1163 (N_1163,N_971,N_753);
nor U1164 (N_1164,N_528,N_943);
or U1165 (N_1165,N_509,N_932);
and U1166 (N_1166,N_658,N_974);
nor U1167 (N_1167,N_566,N_737);
nor U1168 (N_1168,N_851,N_858);
and U1169 (N_1169,N_721,N_852);
nand U1170 (N_1170,N_764,N_748);
or U1171 (N_1171,N_638,N_667);
nand U1172 (N_1172,N_715,N_590);
nor U1173 (N_1173,N_577,N_904);
nor U1174 (N_1174,N_801,N_752);
or U1175 (N_1175,N_659,N_958);
and U1176 (N_1176,N_725,N_792);
and U1177 (N_1177,N_862,N_805);
or U1178 (N_1178,N_908,N_907);
nand U1179 (N_1179,N_652,N_985);
and U1180 (N_1180,N_670,N_607);
and U1181 (N_1181,N_539,N_592);
and U1182 (N_1182,N_500,N_619);
nand U1183 (N_1183,N_711,N_707);
or U1184 (N_1184,N_718,N_685);
nor U1185 (N_1185,N_655,N_615);
nor U1186 (N_1186,N_776,N_736);
nor U1187 (N_1187,N_529,N_600);
or U1188 (N_1188,N_872,N_859);
nor U1189 (N_1189,N_613,N_795);
and U1190 (N_1190,N_672,N_525);
or U1191 (N_1191,N_897,N_910);
nor U1192 (N_1192,N_664,N_554);
and U1193 (N_1193,N_827,N_562);
nand U1194 (N_1194,N_894,N_927);
or U1195 (N_1195,N_804,N_699);
nor U1196 (N_1196,N_902,N_546);
and U1197 (N_1197,N_649,N_837);
or U1198 (N_1198,N_756,N_876);
nor U1199 (N_1199,N_809,N_781);
nand U1200 (N_1200,N_936,N_543);
or U1201 (N_1201,N_825,N_642);
or U1202 (N_1202,N_740,N_965);
or U1203 (N_1203,N_840,N_979);
nor U1204 (N_1204,N_749,N_745);
or U1205 (N_1205,N_504,N_660);
nor U1206 (N_1206,N_846,N_743);
and U1207 (N_1207,N_983,N_624);
nor U1208 (N_1208,N_717,N_881);
and U1209 (N_1209,N_769,N_612);
or U1210 (N_1210,N_968,N_797);
or U1211 (N_1211,N_542,N_917);
nor U1212 (N_1212,N_790,N_898);
and U1213 (N_1213,N_593,N_701);
or U1214 (N_1214,N_576,N_818);
nor U1215 (N_1215,N_775,N_955);
and U1216 (N_1216,N_967,N_853);
and U1217 (N_1217,N_722,N_833);
or U1218 (N_1218,N_821,N_524);
nor U1219 (N_1219,N_856,N_729);
and U1220 (N_1220,N_668,N_733);
nor U1221 (N_1221,N_984,N_579);
nand U1222 (N_1222,N_873,N_647);
and U1223 (N_1223,N_533,N_831);
and U1224 (N_1224,N_522,N_948);
nor U1225 (N_1225,N_784,N_515);
nor U1226 (N_1226,N_605,N_884);
nor U1227 (N_1227,N_726,N_572);
nand U1228 (N_1228,N_518,N_945);
nand U1229 (N_1229,N_867,N_687);
or U1230 (N_1230,N_691,N_541);
nor U1231 (N_1231,N_900,N_520);
nor U1232 (N_1232,N_855,N_584);
or U1233 (N_1233,N_928,N_657);
nor U1234 (N_1234,N_501,N_581);
xnor U1235 (N_1235,N_977,N_925);
and U1236 (N_1236,N_850,N_811);
nand U1237 (N_1237,N_913,N_530);
nor U1238 (N_1238,N_578,N_565);
or U1239 (N_1239,N_641,N_987);
or U1240 (N_1240,N_608,N_912);
nand U1241 (N_1241,N_728,N_938);
nand U1242 (N_1242,N_741,N_648);
or U1243 (N_1243,N_836,N_759);
and U1244 (N_1244,N_637,N_887);
nor U1245 (N_1245,N_857,N_919);
nor U1246 (N_1246,N_889,N_808);
nand U1247 (N_1247,N_606,N_994);
or U1248 (N_1248,N_770,N_535);
or U1249 (N_1249,N_682,N_834);
and U1250 (N_1250,N_585,N_785);
nor U1251 (N_1251,N_507,N_703);
nand U1252 (N_1252,N_932,N_635);
or U1253 (N_1253,N_546,N_699);
and U1254 (N_1254,N_526,N_697);
and U1255 (N_1255,N_519,N_749);
or U1256 (N_1256,N_589,N_696);
or U1257 (N_1257,N_574,N_564);
nor U1258 (N_1258,N_825,N_643);
nor U1259 (N_1259,N_755,N_848);
or U1260 (N_1260,N_504,N_853);
nand U1261 (N_1261,N_547,N_706);
nor U1262 (N_1262,N_863,N_937);
and U1263 (N_1263,N_863,N_699);
or U1264 (N_1264,N_916,N_898);
nand U1265 (N_1265,N_731,N_724);
and U1266 (N_1266,N_788,N_799);
nand U1267 (N_1267,N_740,N_684);
and U1268 (N_1268,N_747,N_893);
nor U1269 (N_1269,N_876,N_845);
nor U1270 (N_1270,N_578,N_829);
xor U1271 (N_1271,N_510,N_922);
or U1272 (N_1272,N_608,N_713);
nand U1273 (N_1273,N_667,N_878);
or U1274 (N_1274,N_914,N_625);
and U1275 (N_1275,N_761,N_914);
nand U1276 (N_1276,N_963,N_560);
and U1277 (N_1277,N_632,N_668);
and U1278 (N_1278,N_999,N_603);
nor U1279 (N_1279,N_927,N_615);
nor U1280 (N_1280,N_913,N_715);
nand U1281 (N_1281,N_586,N_624);
or U1282 (N_1282,N_993,N_976);
and U1283 (N_1283,N_920,N_600);
and U1284 (N_1284,N_763,N_724);
or U1285 (N_1285,N_962,N_765);
or U1286 (N_1286,N_546,N_586);
or U1287 (N_1287,N_682,N_642);
nor U1288 (N_1288,N_589,N_505);
nand U1289 (N_1289,N_500,N_947);
nand U1290 (N_1290,N_684,N_934);
or U1291 (N_1291,N_819,N_849);
nand U1292 (N_1292,N_763,N_866);
nand U1293 (N_1293,N_525,N_567);
nor U1294 (N_1294,N_800,N_566);
or U1295 (N_1295,N_689,N_612);
or U1296 (N_1296,N_943,N_630);
and U1297 (N_1297,N_932,N_707);
nor U1298 (N_1298,N_724,N_751);
and U1299 (N_1299,N_574,N_954);
or U1300 (N_1300,N_533,N_906);
or U1301 (N_1301,N_813,N_740);
or U1302 (N_1302,N_872,N_966);
or U1303 (N_1303,N_542,N_898);
or U1304 (N_1304,N_557,N_627);
nor U1305 (N_1305,N_846,N_773);
or U1306 (N_1306,N_629,N_691);
and U1307 (N_1307,N_910,N_501);
nand U1308 (N_1308,N_643,N_821);
and U1309 (N_1309,N_599,N_844);
and U1310 (N_1310,N_951,N_658);
and U1311 (N_1311,N_992,N_750);
nor U1312 (N_1312,N_660,N_944);
nand U1313 (N_1313,N_534,N_850);
nand U1314 (N_1314,N_895,N_765);
nand U1315 (N_1315,N_577,N_608);
and U1316 (N_1316,N_907,N_507);
and U1317 (N_1317,N_707,N_721);
nor U1318 (N_1318,N_625,N_750);
or U1319 (N_1319,N_664,N_772);
nor U1320 (N_1320,N_894,N_998);
nor U1321 (N_1321,N_566,N_927);
nand U1322 (N_1322,N_527,N_771);
and U1323 (N_1323,N_889,N_513);
xor U1324 (N_1324,N_519,N_717);
xnor U1325 (N_1325,N_898,N_921);
nand U1326 (N_1326,N_794,N_819);
nor U1327 (N_1327,N_532,N_950);
and U1328 (N_1328,N_684,N_998);
and U1329 (N_1329,N_792,N_631);
or U1330 (N_1330,N_681,N_980);
nand U1331 (N_1331,N_971,N_584);
or U1332 (N_1332,N_870,N_810);
nor U1333 (N_1333,N_724,N_639);
and U1334 (N_1334,N_677,N_551);
nand U1335 (N_1335,N_716,N_875);
nor U1336 (N_1336,N_891,N_964);
or U1337 (N_1337,N_808,N_798);
or U1338 (N_1338,N_640,N_748);
or U1339 (N_1339,N_583,N_540);
nand U1340 (N_1340,N_986,N_933);
xor U1341 (N_1341,N_962,N_894);
nor U1342 (N_1342,N_926,N_574);
and U1343 (N_1343,N_732,N_791);
or U1344 (N_1344,N_596,N_955);
or U1345 (N_1345,N_817,N_740);
or U1346 (N_1346,N_947,N_564);
or U1347 (N_1347,N_531,N_763);
nand U1348 (N_1348,N_636,N_577);
and U1349 (N_1349,N_796,N_741);
or U1350 (N_1350,N_591,N_608);
nand U1351 (N_1351,N_937,N_875);
or U1352 (N_1352,N_649,N_846);
nor U1353 (N_1353,N_751,N_814);
and U1354 (N_1354,N_567,N_971);
nor U1355 (N_1355,N_679,N_788);
nor U1356 (N_1356,N_722,N_605);
and U1357 (N_1357,N_629,N_663);
or U1358 (N_1358,N_746,N_682);
and U1359 (N_1359,N_694,N_569);
nor U1360 (N_1360,N_527,N_583);
nand U1361 (N_1361,N_519,N_637);
nor U1362 (N_1362,N_752,N_552);
or U1363 (N_1363,N_591,N_899);
and U1364 (N_1364,N_618,N_765);
nand U1365 (N_1365,N_611,N_830);
and U1366 (N_1366,N_843,N_508);
and U1367 (N_1367,N_776,N_666);
nand U1368 (N_1368,N_702,N_950);
nand U1369 (N_1369,N_623,N_942);
or U1370 (N_1370,N_753,N_696);
nand U1371 (N_1371,N_825,N_650);
nand U1372 (N_1372,N_675,N_521);
nor U1373 (N_1373,N_908,N_603);
and U1374 (N_1374,N_936,N_520);
nand U1375 (N_1375,N_656,N_696);
nand U1376 (N_1376,N_926,N_633);
nor U1377 (N_1377,N_561,N_618);
nand U1378 (N_1378,N_934,N_909);
or U1379 (N_1379,N_824,N_947);
nor U1380 (N_1380,N_840,N_927);
or U1381 (N_1381,N_871,N_644);
nor U1382 (N_1382,N_812,N_826);
nand U1383 (N_1383,N_773,N_601);
and U1384 (N_1384,N_545,N_521);
or U1385 (N_1385,N_736,N_886);
and U1386 (N_1386,N_824,N_669);
nand U1387 (N_1387,N_919,N_805);
nand U1388 (N_1388,N_752,N_874);
nand U1389 (N_1389,N_999,N_607);
nor U1390 (N_1390,N_834,N_753);
and U1391 (N_1391,N_721,N_928);
nand U1392 (N_1392,N_959,N_870);
and U1393 (N_1393,N_519,N_553);
and U1394 (N_1394,N_973,N_717);
nor U1395 (N_1395,N_688,N_994);
or U1396 (N_1396,N_800,N_720);
nand U1397 (N_1397,N_786,N_797);
nor U1398 (N_1398,N_890,N_713);
nand U1399 (N_1399,N_783,N_801);
nand U1400 (N_1400,N_690,N_536);
nor U1401 (N_1401,N_560,N_758);
xnor U1402 (N_1402,N_516,N_906);
nand U1403 (N_1403,N_678,N_654);
nand U1404 (N_1404,N_951,N_542);
or U1405 (N_1405,N_943,N_764);
and U1406 (N_1406,N_596,N_997);
nor U1407 (N_1407,N_705,N_675);
nor U1408 (N_1408,N_504,N_536);
or U1409 (N_1409,N_921,N_731);
nor U1410 (N_1410,N_810,N_943);
nand U1411 (N_1411,N_795,N_500);
nor U1412 (N_1412,N_951,N_879);
or U1413 (N_1413,N_950,N_934);
nor U1414 (N_1414,N_980,N_646);
and U1415 (N_1415,N_610,N_846);
nand U1416 (N_1416,N_651,N_557);
nand U1417 (N_1417,N_910,N_587);
or U1418 (N_1418,N_527,N_948);
nor U1419 (N_1419,N_877,N_522);
or U1420 (N_1420,N_718,N_646);
or U1421 (N_1421,N_813,N_769);
nand U1422 (N_1422,N_662,N_672);
nand U1423 (N_1423,N_918,N_748);
nand U1424 (N_1424,N_908,N_549);
or U1425 (N_1425,N_537,N_841);
or U1426 (N_1426,N_673,N_730);
nor U1427 (N_1427,N_596,N_809);
and U1428 (N_1428,N_681,N_850);
nand U1429 (N_1429,N_554,N_546);
and U1430 (N_1430,N_848,N_995);
nor U1431 (N_1431,N_847,N_844);
or U1432 (N_1432,N_795,N_972);
nand U1433 (N_1433,N_917,N_886);
or U1434 (N_1434,N_859,N_961);
nand U1435 (N_1435,N_510,N_955);
nand U1436 (N_1436,N_602,N_956);
nand U1437 (N_1437,N_923,N_938);
nor U1438 (N_1438,N_594,N_809);
or U1439 (N_1439,N_581,N_552);
nand U1440 (N_1440,N_990,N_717);
nor U1441 (N_1441,N_805,N_777);
and U1442 (N_1442,N_918,N_591);
or U1443 (N_1443,N_866,N_546);
or U1444 (N_1444,N_539,N_826);
nand U1445 (N_1445,N_691,N_537);
and U1446 (N_1446,N_908,N_671);
and U1447 (N_1447,N_668,N_660);
or U1448 (N_1448,N_932,N_688);
or U1449 (N_1449,N_881,N_937);
or U1450 (N_1450,N_847,N_683);
nand U1451 (N_1451,N_849,N_675);
nor U1452 (N_1452,N_977,N_911);
and U1453 (N_1453,N_746,N_706);
nor U1454 (N_1454,N_774,N_739);
nor U1455 (N_1455,N_586,N_895);
and U1456 (N_1456,N_517,N_564);
and U1457 (N_1457,N_723,N_733);
or U1458 (N_1458,N_865,N_927);
and U1459 (N_1459,N_997,N_865);
and U1460 (N_1460,N_976,N_546);
nor U1461 (N_1461,N_879,N_854);
and U1462 (N_1462,N_728,N_790);
and U1463 (N_1463,N_990,N_780);
nor U1464 (N_1464,N_976,N_632);
nand U1465 (N_1465,N_915,N_678);
and U1466 (N_1466,N_877,N_699);
or U1467 (N_1467,N_603,N_580);
or U1468 (N_1468,N_606,N_603);
or U1469 (N_1469,N_958,N_558);
nand U1470 (N_1470,N_883,N_928);
nor U1471 (N_1471,N_615,N_686);
or U1472 (N_1472,N_992,N_963);
and U1473 (N_1473,N_738,N_585);
and U1474 (N_1474,N_816,N_714);
nand U1475 (N_1475,N_939,N_891);
or U1476 (N_1476,N_607,N_869);
and U1477 (N_1477,N_845,N_578);
nand U1478 (N_1478,N_946,N_719);
nand U1479 (N_1479,N_574,N_678);
or U1480 (N_1480,N_886,N_704);
xor U1481 (N_1481,N_602,N_798);
nor U1482 (N_1482,N_600,N_661);
and U1483 (N_1483,N_617,N_569);
nor U1484 (N_1484,N_559,N_924);
and U1485 (N_1485,N_948,N_818);
or U1486 (N_1486,N_694,N_993);
or U1487 (N_1487,N_533,N_862);
xnor U1488 (N_1488,N_996,N_976);
nand U1489 (N_1489,N_830,N_605);
nor U1490 (N_1490,N_606,N_951);
nor U1491 (N_1491,N_647,N_587);
nand U1492 (N_1492,N_816,N_931);
or U1493 (N_1493,N_748,N_907);
xnor U1494 (N_1494,N_508,N_597);
nor U1495 (N_1495,N_943,N_745);
and U1496 (N_1496,N_756,N_564);
nor U1497 (N_1497,N_502,N_711);
or U1498 (N_1498,N_887,N_583);
and U1499 (N_1499,N_892,N_517);
nor U1500 (N_1500,N_1412,N_1378);
and U1501 (N_1501,N_1381,N_1213);
nor U1502 (N_1502,N_1462,N_1064);
and U1503 (N_1503,N_1382,N_1401);
nand U1504 (N_1504,N_1302,N_1206);
and U1505 (N_1505,N_1435,N_1455);
nor U1506 (N_1506,N_1334,N_1394);
nand U1507 (N_1507,N_1148,N_1010);
nor U1508 (N_1508,N_1432,N_1078);
or U1509 (N_1509,N_1489,N_1017);
and U1510 (N_1510,N_1217,N_1095);
or U1511 (N_1511,N_1289,N_1236);
or U1512 (N_1512,N_1147,N_1199);
and U1513 (N_1513,N_1397,N_1102);
and U1514 (N_1514,N_1362,N_1109);
nor U1515 (N_1515,N_1439,N_1121);
nand U1516 (N_1516,N_1088,N_1143);
or U1517 (N_1517,N_1417,N_1452);
or U1518 (N_1518,N_1306,N_1360);
and U1519 (N_1519,N_1049,N_1080);
nand U1520 (N_1520,N_1288,N_1136);
or U1521 (N_1521,N_1185,N_1387);
nand U1522 (N_1522,N_1267,N_1426);
or U1523 (N_1523,N_1234,N_1416);
nand U1524 (N_1524,N_1320,N_1488);
nand U1525 (N_1525,N_1056,N_1492);
or U1526 (N_1526,N_1420,N_1443);
or U1527 (N_1527,N_1449,N_1232);
nor U1528 (N_1528,N_1498,N_1166);
and U1529 (N_1529,N_1072,N_1176);
nor U1530 (N_1530,N_1235,N_1347);
and U1531 (N_1531,N_1231,N_1371);
and U1532 (N_1532,N_1421,N_1009);
and U1533 (N_1533,N_1007,N_1035);
and U1534 (N_1534,N_1290,N_1004);
nand U1535 (N_1535,N_1434,N_1295);
nand U1536 (N_1536,N_1238,N_1367);
or U1537 (N_1537,N_1250,N_1260);
nand U1538 (N_1538,N_1301,N_1027);
and U1539 (N_1539,N_1459,N_1285);
or U1540 (N_1540,N_1011,N_1319);
or U1541 (N_1541,N_1144,N_1385);
nor U1542 (N_1542,N_1042,N_1214);
nor U1543 (N_1543,N_1477,N_1113);
nor U1544 (N_1544,N_1265,N_1115);
nand U1545 (N_1545,N_1089,N_1456);
or U1546 (N_1546,N_1356,N_1475);
nor U1547 (N_1547,N_1384,N_1057);
or U1548 (N_1548,N_1066,N_1479);
and U1549 (N_1549,N_1329,N_1076);
nand U1550 (N_1550,N_1087,N_1023);
or U1551 (N_1551,N_1406,N_1457);
or U1552 (N_1552,N_1278,N_1326);
xnor U1553 (N_1553,N_1139,N_1386);
nor U1554 (N_1554,N_1225,N_1468);
or U1555 (N_1555,N_1469,N_1200);
nor U1556 (N_1556,N_1157,N_1149);
nand U1557 (N_1557,N_1476,N_1338);
nand U1558 (N_1558,N_1203,N_1237);
nand U1559 (N_1559,N_1103,N_1252);
and U1560 (N_1560,N_1163,N_1445);
or U1561 (N_1561,N_1423,N_1305);
and U1562 (N_1562,N_1204,N_1105);
or U1563 (N_1563,N_1414,N_1090);
nor U1564 (N_1564,N_1341,N_1496);
nor U1565 (N_1565,N_1248,N_1352);
or U1566 (N_1566,N_1344,N_1211);
nand U1567 (N_1567,N_1363,N_1467);
nand U1568 (N_1568,N_1133,N_1466);
and U1569 (N_1569,N_1030,N_1240);
nand U1570 (N_1570,N_1458,N_1291);
nor U1571 (N_1571,N_1223,N_1330);
or U1572 (N_1572,N_1368,N_1107);
nand U1573 (N_1573,N_1298,N_1034);
nand U1574 (N_1574,N_1059,N_1471);
nor U1575 (N_1575,N_1297,N_1257);
and U1576 (N_1576,N_1465,N_1051);
nand U1577 (N_1577,N_1001,N_1138);
and U1578 (N_1578,N_1392,N_1114);
or U1579 (N_1579,N_1012,N_1081);
nor U1580 (N_1580,N_1120,N_1020);
nand U1581 (N_1581,N_1170,N_1348);
or U1582 (N_1582,N_1155,N_1047);
nand U1583 (N_1583,N_1125,N_1003);
or U1584 (N_1584,N_1304,N_1427);
or U1585 (N_1585,N_1415,N_1242);
and U1586 (N_1586,N_1039,N_1050);
or U1587 (N_1587,N_1379,N_1013);
or U1588 (N_1588,N_1069,N_1116);
or U1589 (N_1589,N_1182,N_1097);
and U1590 (N_1590,N_1438,N_1118);
xor U1591 (N_1591,N_1111,N_1393);
and U1592 (N_1592,N_1303,N_1311);
and U1593 (N_1593,N_1454,N_1318);
nand U1594 (N_1594,N_1032,N_1487);
and U1595 (N_1595,N_1159,N_1130);
nand U1596 (N_1596,N_1191,N_1346);
nor U1597 (N_1597,N_1171,N_1422);
or U1598 (N_1598,N_1000,N_1212);
and U1599 (N_1599,N_1349,N_1292);
xor U1600 (N_1600,N_1307,N_1046);
or U1601 (N_1601,N_1286,N_1486);
or U1602 (N_1602,N_1036,N_1135);
or U1603 (N_1603,N_1315,N_1294);
nand U1604 (N_1604,N_1282,N_1313);
or U1605 (N_1605,N_1150,N_1075);
nand U1606 (N_1606,N_1332,N_1437);
nand U1607 (N_1607,N_1372,N_1016);
nor U1608 (N_1608,N_1430,N_1140);
nand U1609 (N_1609,N_1272,N_1428);
and U1610 (N_1610,N_1424,N_1491);
or U1611 (N_1611,N_1029,N_1048);
or U1612 (N_1612,N_1308,N_1331);
or U1613 (N_1613,N_1209,N_1085);
nand U1614 (N_1614,N_1403,N_1126);
and U1615 (N_1615,N_1407,N_1178);
and U1616 (N_1616,N_1061,N_1141);
nor U1617 (N_1617,N_1196,N_1478);
nor U1618 (N_1618,N_1262,N_1131);
nor U1619 (N_1619,N_1339,N_1377);
or U1620 (N_1620,N_1092,N_1220);
or U1621 (N_1621,N_1296,N_1222);
nor U1622 (N_1622,N_1345,N_1499);
and U1623 (N_1623,N_1173,N_1192);
and U1624 (N_1624,N_1253,N_1172);
nor U1625 (N_1625,N_1084,N_1184);
or U1626 (N_1626,N_1255,N_1482);
or U1627 (N_1627,N_1207,N_1431);
or U1628 (N_1628,N_1383,N_1463);
nor U1629 (N_1629,N_1104,N_1152);
nand U1630 (N_1630,N_1151,N_1227);
and U1631 (N_1631,N_1497,N_1336);
and U1632 (N_1632,N_1472,N_1380);
nand U1633 (N_1633,N_1040,N_1083);
and U1634 (N_1634,N_1256,N_1146);
or U1635 (N_1635,N_1074,N_1280);
nand U1636 (N_1636,N_1015,N_1405);
nand U1637 (N_1637,N_1054,N_1321);
or U1638 (N_1638,N_1183,N_1395);
nor U1639 (N_1639,N_1440,N_1300);
or U1640 (N_1640,N_1110,N_1094);
nor U1641 (N_1641,N_1293,N_1413);
and U1642 (N_1642,N_1369,N_1484);
nor U1643 (N_1643,N_1275,N_1241);
nand U1644 (N_1644,N_1408,N_1419);
nand U1645 (N_1645,N_1038,N_1274);
and U1646 (N_1646,N_1441,N_1358);
and U1647 (N_1647,N_1019,N_1106);
nand U1648 (N_1648,N_1194,N_1216);
nor U1649 (N_1649,N_1266,N_1355);
nor U1650 (N_1650,N_1108,N_1327);
nand U1651 (N_1651,N_1366,N_1096);
or U1652 (N_1652,N_1495,N_1208);
or U1653 (N_1653,N_1022,N_1021);
or U1654 (N_1654,N_1228,N_1180);
and U1655 (N_1655,N_1376,N_1276);
or U1656 (N_1656,N_1134,N_1205);
nand U1657 (N_1657,N_1229,N_1335);
nand U1658 (N_1658,N_1317,N_1370);
or U1659 (N_1659,N_1063,N_1142);
and U1660 (N_1660,N_1071,N_1145);
or U1661 (N_1661,N_1156,N_1247);
nor U1662 (N_1662,N_1337,N_1091);
nor U1663 (N_1663,N_1243,N_1068);
and U1664 (N_1664,N_1364,N_1357);
or U1665 (N_1665,N_1198,N_1167);
or U1666 (N_1666,N_1480,N_1398);
and U1667 (N_1667,N_1444,N_1093);
and U1668 (N_1668,N_1351,N_1060);
or U1669 (N_1669,N_1005,N_1375);
or U1670 (N_1670,N_1448,N_1045);
nor U1671 (N_1671,N_1284,N_1129);
nor U1672 (N_1672,N_1239,N_1224);
nor U1673 (N_1673,N_1154,N_1450);
nand U1674 (N_1674,N_1174,N_1188);
nand U1675 (N_1675,N_1100,N_1098);
and U1676 (N_1676,N_1067,N_1165);
or U1677 (N_1677,N_1436,N_1244);
nor U1678 (N_1678,N_1388,N_1195);
nor U1679 (N_1679,N_1254,N_1418);
nor U1680 (N_1680,N_1202,N_1189);
and U1681 (N_1681,N_1197,N_1123);
nor U1682 (N_1682,N_1014,N_1446);
or U1683 (N_1683,N_1354,N_1079);
nand U1684 (N_1684,N_1041,N_1353);
or U1685 (N_1685,N_1055,N_1324);
and U1686 (N_1686,N_1132,N_1028);
or U1687 (N_1687,N_1481,N_1323);
or U1688 (N_1688,N_1391,N_1077);
or U1689 (N_1689,N_1442,N_1230);
or U1690 (N_1690,N_1164,N_1246);
and U1691 (N_1691,N_1187,N_1026);
or U1692 (N_1692,N_1429,N_1474);
nand U1693 (N_1693,N_1433,N_1396);
nor U1694 (N_1694,N_1470,N_1117);
or U1695 (N_1695,N_1158,N_1374);
nand U1696 (N_1696,N_1400,N_1264);
nand U1697 (N_1697,N_1124,N_1287);
or U1698 (N_1698,N_1404,N_1086);
nand U1699 (N_1699,N_1314,N_1177);
nor U1700 (N_1700,N_1390,N_1219);
or U1701 (N_1701,N_1490,N_1112);
or U1702 (N_1702,N_1277,N_1322);
nor U1703 (N_1703,N_1190,N_1312);
nand U1704 (N_1704,N_1210,N_1411);
nor U1705 (N_1705,N_1161,N_1218);
and U1706 (N_1706,N_1122,N_1160);
or U1707 (N_1707,N_1447,N_1044);
nand U1708 (N_1708,N_1031,N_1065);
and U1709 (N_1709,N_1245,N_1451);
nor U1710 (N_1710,N_1485,N_1261);
nand U1711 (N_1711,N_1179,N_1299);
nand U1712 (N_1712,N_1181,N_1309);
and U1713 (N_1713,N_1410,N_1328);
nand U1714 (N_1714,N_1283,N_1453);
nand U1715 (N_1715,N_1073,N_1062);
or U1716 (N_1716,N_1006,N_1251);
nor U1717 (N_1717,N_1037,N_1258);
nor U1718 (N_1718,N_1402,N_1226);
nor U1719 (N_1719,N_1101,N_1186);
nor U1720 (N_1720,N_1070,N_1221);
nor U1721 (N_1721,N_1270,N_1193);
nor U1722 (N_1722,N_1233,N_1153);
nand U1723 (N_1723,N_1002,N_1461);
and U1724 (N_1724,N_1024,N_1316);
nor U1725 (N_1725,N_1494,N_1052);
nor U1726 (N_1726,N_1249,N_1119);
or U1727 (N_1727,N_1373,N_1215);
and U1728 (N_1728,N_1271,N_1058);
nand U1729 (N_1729,N_1361,N_1082);
or U1730 (N_1730,N_1043,N_1268);
and U1731 (N_1731,N_1162,N_1128);
nor U1732 (N_1732,N_1263,N_1342);
nor U1733 (N_1733,N_1025,N_1273);
and U1734 (N_1734,N_1269,N_1493);
or U1735 (N_1735,N_1008,N_1175);
xor U1736 (N_1736,N_1389,N_1483);
nor U1737 (N_1737,N_1359,N_1343);
and U1738 (N_1738,N_1127,N_1365);
nor U1739 (N_1739,N_1137,N_1099);
or U1740 (N_1740,N_1279,N_1399);
nor U1741 (N_1741,N_1473,N_1350);
and U1742 (N_1742,N_1409,N_1259);
or U1743 (N_1743,N_1425,N_1464);
and U1744 (N_1744,N_1333,N_1201);
or U1745 (N_1745,N_1281,N_1053);
and U1746 (N_1746,N_1168,N_1169);
nand U1747 (N_1747,N_1325,N_1460);
and U1748 (N_1748,N_1310,N_1340);
nor U1749 (N_1749,N_1018,N_1033);
or U1750 (N_1750,N_1356,N_1256);
and U1751 (N_1751,N_1499,N_1313);
or U1752 (N_1752,N_1183,N_1257);
nor U1753 (N_1753,N_1206,N_1452);
nand U1754 (N_1754,N_1294,N_1012);
nand U1755 (N_1755,N_1052,N_1247);
or U1756 (N_1756,N_1361,N_1384);
nor U1757 (N_1757,N_1419,N_1273);
or U1758 (N_1758,N_1288,N_1494);
or U1759 (N_1759,N_1258,N_1351);
or U1760 (N_1760,N_1346,N_1467);
nand U1761 (N_1761,N_1010,N_1396);
nand U1762 (N_1762,N_1004,N_1331);
and U1763 (N_1763,N_1407,N_1447);
and U1764 (N_1764,N_1103,N_1174);
nor U1765 (N_1765,N_1124,N_1420);
nand U1766 (N_1766,N_1163,N_1223);
or U1767 (N_1767,N_1378,N_1246);
nor U1768 (N_1768,N_1486,N_1340);
or U1769 (N_1769,N_1277,N_1483);
or U1770 (N_1770,N_1397,N_1138);
or U1771 (N_1771,N_1433,N_1209);
or U1772 (N_1772,N_1411,N_1134);
nor U1773 (N_1773,N_1163,N_1307);
and U1774 (N_1774,N_1012,N_1425);
or U1775 (N_1775,N_1080,N_1175);
or U1776 (N_1776,N_1145,N_1093);
nand U1777 (N_1777,N_1345,N_1218);
xor U1778 (N_1778,N_1229,N_1371);
nand U1779 (N_1779,N_1457,N_1211);
or U1780 (N_1780,N_1008,N_1251);
nor U1781 (N_1781,N_1368,N_1062);
nor U1782 (N_1782,N_1007,N_1096);
nand U1783 (N_1783,N_1231,N_1254);
or U1784 (N_1784,N_1049,N_1469);
nor U1785 (N_1785,N_1221,N_1010);
or U1786 (N_1786,N_1169,N_1475);
or U1787 (N_1787,N_1407,N_1309);
and U1788 (N_1788,N_1006,N_1402);
and U1789 (N_1789,N_1352,N_1264);
nor U1790 (N_1790,N_1252,N_1048);
nand U1791 (N_1791,N_1410,N_1448);
and U1792 (N_1792,N_1392,N_1145);
nor U1793 (N_1793,N_1008,N_1091);
nand U1794 (N_1794,N_1009,N_1186);
or U1795 (N_1795,N_1380,N_1190);
and U1796 (N_1796,N_1217,N_1379);
nor U1797 (N_1797,N_1425,N_1266);
nor U1798 (N_1798,N_1033,N_1113);
or U1799 (N_1799,N_1104,N_1250);
or U1800 (N_1800,N_1245,N_1158);
and U1801 (N_1801,N_1024,N_1391);
and U1802 (N_1802,N_1463,N_1451);
nand U1803 (N_1803,N_1341,N_1357);
nand U1804 (N_1804,N_1146,N_1306);
nand U1805 (N_1805,N_1070,N_1031);
nor U1806 (N_1806,N_1175,N_1384);
and U1807 (N_1807,N_1393,N_1031);
nand U1808 (N_1808,N_1199,N_1419);
or U1809 (N_1809,N_1482,N_1245);
and U1810 (N_1810,N_1256,N_1147);
or U1811 (N_1811,N_1377,N_1197);
and U1812 (N_1812,N_1444,N_1395);
nand U1813 (N_1813,N_1386,N_1295);
nand U1814 (N_1814,N_1344,N_1092);
nand U1815 (N_1815,N_1219,N_1409);
or U1816 (N_1816,N_1360,N_1224);
nand U1817 (N_1817,N_1356,N_1010);
nor U1818 (N_1818,N_1045,N_1302);
and U1819 (N_1819,N_1102,N_1433);
and U1820 (N_1820,N_1118,N_1072);
and U1821 (N_1821,N_1324,N_1108);
and U1822 (N_1822,N_1183,N_1036);
and U1823 (N_1823,N_1448,N_1260);
and U1824 (N_1824,N_1058,N_1330);
and U1825 (N_1825,N_1131,N_1239);
or U1826 (N_1826,N_1377,N_1391);
nand U1827 (N_1827,N_1199,N_1146);
nor U1828 (N_1828,N_1466,N_1489);
and U1829 (N_1829,N_1280,N_1432);
nor U1830 (N_1830,N_1371,N_1011);
nand U1831 (N_1831,N_1088,N_1322);
or U1832 (N_1832,N_1162,N_1330);
nand U1833 (N_1833,N_1469,N_1454);
nand U1834 (N_1834,N_1029,N_1469);
nand U1835 (N_1835,N_1415,N_1089);
and U1836 (N_1836,N_1215,N_1263);
nand U1837 (N_1837,N_1203,N_1193);
nand U1838 (N_1838,N_1118,N_1021);
nand U1839 (N_1839,N_1472,N_1237);
nand U1840 (N_1840,N_1016,N_1318);
or U1841 (N_1841,N_1049,N_1240);
and U1842 (N_1842,N_1429,N_1445);
and U1843 (N_1843,N_1452,N_1054);
and U1844 (N_1844,N_1340,N_1394);
or U1845 (N_1845,N_1162,N_1485);
nor U1846 (N_1846,N_1395,N_1130);
nand U1847 (N_1847,N_1399,N_1354);
nor U1848 (N_1848,N_1134,N_1227);
nand U1849 (N_1849,N_1252,N_1105);
nand U1850 (N_1850,N_1235,N_1292);
nor U1851 (N_1851,N_1124,N_1315);
nand U1852 (N_1852,N_1352,N_1014);
nor U1853 (N_1853,N_1183,N_1350);
or U1854 (N_1854,N_1298,N_1374);
nor U1855 (N_1855,N_1105,N_1406);
and U1856 (N_1856,N_1271,N_1221);
or U1857 (N_1857,N_1388,N_1358);
and U1858 (N_1858,N_1443,N_1322);
nor U1859 (N_1859,N_1252,N_1416);
or U1860 (N_1860,N_1470,N_1270);
and U1861 (N_1861,N_1300,N_1247);
or U1862 (N_1862,N_1228,N_1115);
and U1863 (N_1863,N_1261,N_1149);
or U1864 (N_1864,N_1393,N_1387);
or U1865 (N_1865,N_1300,N_1090);
or U1866 (N_1866,N_1353,N_1083);
or U1867 (N_1867,N_1332,N_1141);
nor U1868 (N_1868,N_1353,N_1423);
nor U1869 (N_1869,N_1295,N_1276);
and U1870 (N_1870,N_1172,N_1376);
or U1871 (N_1871,N_1251,N_1028);
and U1872 (N_1872,N_1483,N_1027);
nand U1873 (N_1873,N_1218,N_1048);
nand U1874 (N_1874,N_1367,N_1123);
nor U1875 (N_1875,N_1193,N_1021);
nor U1876 (N_1876,N_1181,N_1149);
nor U1877 (N_1877,N_1253,N_1489);
nand U1878 (N_1878,N_1172,N_1325);
nand U1879 (N_1879,N_1204,N_1296);
nor U1880 (N_1880,N_1453,N_1155);
nor U1881 (N_1881,N_1159,N_1107);
or U1882 (N_1882,N_1175,N_1004);
nor U1883 (N_1883,N_1431,N_1392);
or U1884 (N_1884,N_1293,N_1088);
nor U1885 (N_1885,N_1496,N_1377);
nand U1886 (N_1886,N_1031,N_1133);
and U1887 (N_1887,N_1160,N_1305);
or U1888 (N_1888,N_1059,N_1034);
and U1889 (N_1889,N_1336,N_1434);
nor U1890 (N_1890,N_1153,N_1156);
nand U1891 (N_1891,N_1470,N_1223);
and U1892 (N_1892,N_1418,N_1429);
or U1893 (N_1893,N_1411,N_1385);
and U1894 (N_1894,N_1435,N_1198);
nand U1895 (N_1895,N_1277,N_1224);
and U1896 (N_1896,N_1205,N_1080);
nand U1897 (N_1897,N_1060,N_1391);
nor U1898 (N_1898,N_1115,N_1057);
nand U1899 (N_1899,N_1229,N_1025);
and U1900 (N_1900,N_1441,N_1053);
nand U1901 (N_1901,N_1104,N_1436);
and U1902 (N_1902,N_1243,N_1082);
or U1903 (N_1903,N_1215,N_1350);
and U1904 (N_1904,N_1285,N_1208);
nand U1905 (N_1905,N_1120,N_1372);
nor U1906 (N_1906,N_1106,N_1174);
or U1907 (N_1907,N_1376,N_1409);
nand U1908 (N_1908,N_1036,N_1439);
or U1909 (N_1909,N_1134,N_1224);
or U1910 (N_1910,N_1469,N_1023);
nor U1911 (N_1911,N_1261,N_1315);
nor U1912 (N_1912,N_1049,N_1105);
or U1913 (N_1913,N_1325,N_1047);
and U1914 (N_1914,N_1083,N_1486);
xor U1915 (N_1915,N_1415,N_1401);
nor U1916 (N_1916,N_1330,N_1294);
nor U1917 (N_1917,N_1449,N_1057);
nor U1918 (N_1918,N_1257,N_1326);
nor U1919 (N_1919,N_1476,N_1027);
or U1920 (N_1920,N_1130,N_1156);
and U1921 (N_1921,N_1131,N_1463);
and U1922 (N_1922,N_1345,N_1242);
or U1923 (N_1923,N_1493,N_1435);
nand U1924 (N_1924,N_1269,N_1385);
or U1925 (N_1925,N_1021,N_1366);
nor U1926 (N_1926,N_1398,N_1157);
and U1927 (N_1927,N_1454,N_1358);
nor U1928 (N_1928,N_1290,N_1391);
and U1929 (N_1929,N_1125,N_1276);
or U1930 (N_1930,N_1383,N_1477);
and U1931 (N_1931,N_1461,N_1114);
and U1932 (N_1932,N_1293,N_1042);
or U1933 (N_1933,N_1356,N_1268);
and U1934 (N_1934,N_1265,N_1068);
nand U1935 (N_1935,N_1087,N_1460);
and U1936 (N_1936,N_1433,N_1361);
nand U1937 (N_1937,N_1307,N_1498);
nand U1938 (N_1938,N_1144,N_1072);
nand U1939 (N_1939,N_1021,N_1148);
or U1940 (N_1940,N_1410,N_1336);
nor U1941 (N_1941,N_1424,N_1293);
nor U1942 (N_1942,N_1270,N_1063);
or U1943 (N_1943,N_1028,N_1156);
or U1944 (N_1944,N_1475,N_1466);
nor U1945 (N_1945,N_1464,N_1183);
or U1946 (N_1946,N_1458,N_1372);
nor U1947 (N_1947,N_1295,N_1047);
or U1948 (N_1948,N_1469,N_1342);
or U1949 (N_1949,N_1385,N_1251);
or U1950 (N_1950,N_1187,N_1299);
or U1951 (N_1951,N_1158,N_1038);
nand U1952 (N_1952,N_1469,N_1199);
and U1953 (N_1953,N_1176,N_1180);
or U1954 (N_1954,N_1240,N_1115);
nor U1955 (N_1955,N_1244,N_1423);
and U1956 (N_1956,N_1244,N_1419);
and U1957 (N_1957,N_1124,N_1173);
or U1958 (N_1958,N_1162,N_1149);
and U1959 (N_1959,N_1060,N_1256);
nor U1960 (N_1960,N_1014,N_1202);
nor U1961 (N_1961,N_1473,N_1310);
and U1962 (N_1962,N_1477,N_1425);
nand U1963 (N_1963,N_1258,N_1141);
or U1964 (N_1964,N_1480,N_1466);
nor U1965 (N_1965,N_1118,N_1133);
nand U1966 (N_1966,N_1318,N_1167);
nor U1967 (N_1967,N_1244,N_1228);
nor U1968 (N_1968,N_1132,N_1182);
and U1969 (N_1969,N_1294,N_1049);
xnor U1970 (N_1970,N_1127,N_1010);
nor U1971 (N_1971,N_1420,N_1492);
nand U1972 (N_1972,N_1494,N_1089);
nor U1973 (N_1973,N_1133,N_1298);
xnor U1974 (N_1974,N_1246,N_1074);
nand U1975 (N_1975,N_1201,N_1024);
or U1976 (N_1976,N_1230,N_1182);
nand U1977 (N_1977,N_1486,N_1029);
nor U1978 (N_1978,N_1354,N_1476);
or U1979 (N_1979,N_1487,N_1249);
nand U1980 (N_1980,N_1428,N_1212);
or U1981 (N_1981,N_1311,N_1421);
nor U1982 (N_1982,N_1392,N_1419);
nand U1983 (N_1983,N_1060,N_1196);
or U1984 (N_1984,N_1438,N_1286);
and U1985 (N_1985,N_1352,N_1156);
nand U1986 (N_1986,N_1204,N_1403);
and U1987 (N_1987,N_1003,N_1292);
or U1988 (N_1988,N_1442,N_1330);
or U1989 (N_1989,N_1471,N_1203);
nand U1990 (N_1990,N_1452,N_1408);
or U1991 (N_1991,N_1391,N_1269);
nand U1992 (N_1992,N_1227,N_1156);
or U1993 (N_1993,N_1460,N_1178);
nand U1994 (N_1994,N_1229,N_1285);
or U1995 (N_1995,N_1062,N_1473);
nand U1996 (N_1996,N_1165,N_1474);
nor U1997 (N_1997,N_1469,N_1292);
or U1998 (N_1998,N_1392,N_1300);
nand U1999 (N_1999,N_1466,N_1212);
nor U2000 (N_2000,N_1552,N_1935);
xor U2001 (N_2001,N_1752,N_1586);
nor U2002 (N_2002,N_1634,N_1529);
nor U2003 (N_2003,N_1949,N_1670);
and U2004 (N_2004,N_1735,N_1561);
nor U2005 (N_2005,N_1628,N_1553);
or U2006 (N_2006,N_1546,N_1532);
nor U2007 (N_2007,N_1703,N_1873);
nand U2008 (N_2008,N_1655,N_1896);
and U2009 (N_2009,N_1901,N_1798);
nand U2010 (N_2010,N_1765,N_1698);
nor U2011 (N_2011,N_1519,N_1769);
and U2012 (N_2012,N_1506,N_1936);
nand U2013 (N_2013,N_1893,N_1815);
and U2014 (N_2014,N_1740,N_1800);
nor U2015 (N_2015,N_1932,N_1562);
and U2016 (N_2016,N_1930,N_1504);
and U2017 (N_2017,N_1599,N_1693);
and U2018 (N_2018,N_1672,N_1907);
nor U2019 (N_2019,N_1734,N_1678);
nand U2020 (N_2020,N_1874,N_1831);
nand U2021 (N_2021,N_1807,N_1975);
nand U2022 (N_2022,N_1967,N_1977);
and U2023 (N_2023,N_1652,N_1514);
and U2024 (N_2024,N_1875,N_1702);
nor U2025 (N_2025,N_1609,N_1738);
nor U2026 (N_2026,N_1550,N_1577);
nand U2027 (N_2027,N_1741,N_1952);
nand U2028 (N_2028,N_1786,N_1733);
and U2029 (N_2029,N_1699,N_1757);
nor U2030 (N_2030,N_1887,N_1598);
or U2031 (N_2031,N_1794,N_1864);
nand U2032 (N_2032,N_1938,N_1964);
or U2033 (N_2033,N_1826,N_1872);
nor U2034 (N_2034,N_1857,N_1665);
nor U2035 (N_2035,N_1660,N_1802);
nor U2036 (N_2036,N_1859,N_1908);
or U2037 (N_2037,N_1770,N_1641);
nand U2038 (N_2038,N_1521,N_1870);
nor U2039 (N_2039,N_1775,N_1920);
and U2040 (N_2040,N_1843,N_1902);
xnor U2041 (N_2041,N_1886,N_1994);
or U2042 (N_2042,N_1643,N_1718);
or U2043 (N_2043,N_1829,N_1990);
and U2044 (N_2044,N_1973,N_1675);
or U2045 (N_2045,N_1996,N_1695);
and U2046 (N_2046,N_1814,N_1663);
nor U2047 (N_2047,N_1540,N_1501);
nand U2048 (N_2048,N_1968,N_1632);
and U2049 (N_2049,N_1995,N_1659);
nand U2050 (N_2050,N_1544,N_1604);
nand U2051 (N_2051,N_1500,N_1690);
nand U2052 (N_2052,N_1674,N_1725);
nand U2053 (N_2053,N_1890,N_1899);
and U2054 (N_2054,N_1985,N_1945);
or U2055 (N_2055,N_1841,N_1957);
and U2056 (N_2056,N_1636,N_1897);
and U2057 (N_2057,N_1573,N_1779);
nor U2058 (N_2058,N_1683,N_1568);
nand U2059 (N_2059,N_1768,N_1993);
nand U2060 (N_2060,N_1680,N_1524);
nor U2061 (N_2061,N_1796,N_1523);
nor U2062 (N_2062,N_1502,N_1543);
nand U2063 (N_2063,N_1580,N_1830);
or U2064 (N_2064,N_1928,N_1513);
and U2065 (N_2065,N_1922,N_1608);
or U2066 (N_2066,N_1869,N_1816);
and U2067 (N_2067,N_1943,N_1720);
nor U2068 (N_2068,N_1845,N_1927);
nand U2069 (N_2069,N_1823,N_1732);
and U2070 (N_2070,N_1867,N_1960);
nand U2071 (N_2071,N_1595,N_1700);
and U2072 (N_2072,N_1792,N_1664);
and U2073 (N_2073,N_1976,N_1910);
nand U2074 (N_2074,N_1806,N_1578);
nor U2075 (N_2075,N_1619,N_1926);
or U2076 (N_2076,N_1620,N_1705);
nand U2077 (N_2077,N_1607,N_1605);
nor U2078 (N_2078,N_1853,N_1567);
nor U2079 (N_2079,N_1797,N_1530);
and U2080 (N_2080,N_1582,N_1635);
nor U2081 (N_2081,N_1687,N_1533);
nand U2082 (N_2082,N_1751,N_1618);
nor U2083 (N_2083,N_1746,N_1673);
xor U2084 (N_2084,N_1888,N_1731);
and U2085 (N_2085,N_1756,N_1842);
and U2086 (N_2086,N_1617,N_1820);
nor U2087 (N_2087,N_1653,N_1648);
and U2088 (N_2088,N_1835,N_1689);
nand U2089 (N_2089,N_1566,N_1959);
or U2090 (N_2090,N_1951,N_1772);
or U2091 (N_2091,N_1676,N_1801);
and U2092 (N_2092,N_1851,N_1894);
and U2093 (N_2093,N_1970,N_1818);
nor U2094 (N_2094,N_1627,N_1696);
and U2095 (N_2095,N_1505,N_1759);
nand U2096 (N_2096,N_1724,N_1592);
nor U2097 (N_2097,N_1889,N_1679);
or U2098 (N_2098,N_1623,N_1863);
or U2099 (N_2099,N_1817,N_1526);
nand U2100 (N_2100,N_1531,N_1900);
and U2101 (N_2101,N_1858,N_1677);
nand U2102 (N_2102,N_1574,N_1760);
nand U2103 (N_2103,N_1591,N_1744);
and U2104 (N_2104,N_1511,N_1795);
nor U2105 (N_2105,N_1962,N_1947);
xor U2106 (N_2106,N_1564,N_1658);
nor U2107 (N_2107,N_1998,N_1639);
nor U2108 (N_2108,N_1737,N_1966);
nor U2109 (N_2109,N_1766,N_1833);
or U2110 (N_2110,N_1522,N_1827);
nand U2111 (N_2111,N_1742,N_1767);
nand U2112 (N_2112,N_1915,N_1517);
or U2113 (N_2113,N_1810,N_1545);
and U2114 (N_2114,N_1783,N_1958);
or U2115 (N_2115,N_1644,N_1668);
nand U2116 (N_2116,N_1861,N_1850);
nor U2117 (N_2117,N_1777,N_1905);
nor U2118 (N_2118,N_1822,N_1761);
or U2119 (N_2119,N_1697,N_1560);
or U2120 (N_2120,N_1771,N_1593);
nor U2121 (N_2121,N_1836,N_1981);
nand U2122 (N_2122,N_1860,N_1538);
nand U2123 (N_2123,N_1581,N_1891);
nand U2124 (N_2124,N_1588,N_1610);
and U2125 (N_2125,N_1855,N_1931);
nand U2126 (N_2126,N_1535,N_1862);
and U2127 (N_2127,N_1624,N_1616);
nand U2128 (N_2128,N_1934,N_1984);
and U2129 (N_2129,N_1789,N_1584);
nand U2130 (N_2130,N_1594,N_1730);
nand U2131 (N_2131,N_1667,N_1585);
and U2132 (N_2132,N_1787,N_1963);
nand U2133 (N_2133,N_1914,N_1986);
nor U2134 (N_2134,N_1704,N_1763);
nand U2135 (N_2135,N_1969,N_1729);
nor U2136 (N_2136,N_1856,N_1534);
nor U2137 (N_2137,N_1603,N_1681);
or U2138 (N_2138,N_1716,N_1811);
or U2139 (N_2139,N_1812,N_1754);
nor U2140 (N_2140,N_1551,N_1509);
and U2141 (N_2141,N_1903,N_1512);
nor U2142 (N_2142,N_1837,N_1528);
and U2143 (N_2143,N_1909,N_1991);
nand U2144 (N_2144,N_1953,N_1656);
and U2145 (N_2145,N_1971,N_1999);
nor U2146 (N_2146,N_1865,N_1898);
nor U2147 (N_2147,N_1834,N_1736);
nor U2148 (N_2148,N_1884,N_1694);
nand U2149 (N_2149,N_1590,N_1640);
and U2150 (N_2150,N_1904,N_1715);
or U2151 (N_2151,N_1558,N_1917);
or U2152 (N_2152,N_1684,N_1948);
or U2153 (N_2153,N_1625,N_1753);
and U2154 (N_2154,N_1642,N_1633);
and U2155 (N_2155,N_1921,N_1848);
or U2156 (N_2156,N_1682,N_1638);
nand U2157 (N_2157,N_1776,N_1548);
or U2158 (N_2158,N_1589,N_1979);
nor U2159 (N_2159,N_1537,N_1885);
and U2160 (N_2160,N_1880,N_1507);
and U2161 (N_2161,N_1651,N_1989);
nor U2162 (N_2162,N_1596,N_1838);
nand U2163 (N_2163,N_1944,N_1774);
nand U2164 (N_2164,N_1879,N_1645);
nand U2165 (N_2165,N_1780,N_1709);
and U2166 (N_2166,N_1924,N_1637);
or U2167 (N_2167,N_1671,N_1799);
and U2168 (N_2168,N_1726,N_1954);
and U2169 (N_2169,N_1883,N_1516);
nor U2170 (N_2170,N_1912,N_1868);
nor U2171 (N_2171,N_1743,N_1758);
nor U2172 (N_2172,N_1613,N_1685);
nor U2173 (N_2173,N_1692,N_1961);
and U2174 (N_2174,N_1650,N_1727);
and U2175 (N_2175,N_1950,N_1583);
and U2176 (N_2176,N_1518,N_1929);
and U2177 (N_2177,N_1937,N_1892);
and U2178 (N_2178,N_1847,N_1657);
xnor U2179 (N_2179,N_1755,N_1541);
nand U2180 (N_2180,N_1821,N_1956);
and U2181 (N_2181,N_1721,N_1527);
nor U2182 (N_2182,N_1587,N_1747);
or U2183 (N_2183,N_1974,N_1819);
or U2184 (N_2184,N_1579,N_1788);
nor U2185 (N_2185,N_1626,N_1723);
nand U2186 (N_2186,N_1773,N_1785);
nor U2187 (N_2187,N_1600,N_1946);
nor U2188 (N_2188,N_1749,N_1824);
or U2189 (N_2189,N_1630,N_1666);
nand U2190 (N_2190,N_1876,N_1849);
nand U2191 (N_2191,N_1701,N_1520);
and U2192 (N_2192,N_1622,N_1554);
or U2193 (N_2193,N_1881,N_1846);
or U2194 (N_2194,N_1791,N_1559);
nor U2195 (N_2195,N_1717,N_1722);
nor U2196 (N_2196,N_1965,N_1556);
and U2197 (N_2197,N_1911,N_1955);
or U2198 (N_2198,N_1933,N_1631);
and U2199 (N_2199,N_1525,N_1571);
nand U2200 (N_2200,N_1597,N_1539);
and U2201 (N_2201,N_1918,N_1606);
and U2202 (N_2202,N_1621,N_1601);
and U2203 (N_2203,N_1508,N_1569);
and U2204 (N_2204,N_1750,N_1882);
nor U2205 (N_2205,N_1708,N_1503);
nand U2206 (N_2206,N_1828,N_1808);
or U2207 (N_2207,N_1778,N_1913);
nor U2208 (N_2208,N_1549,N_1992);
or U2209 (N_2209,N_1661,N_1793);
and U2210 (N_2210,N_1565,N_1510);
nand U2211 (N_2211,N_1547,N_1987);
nand U2212 (N_2212,N_1536,N_1982);
or U2213 (N_2213,N_1919,N_1940);
or U2214 (N_2214,N_1844,N_1781);
and U2215 (N_2215,N_1614,N_1941);
and U2216 (N_2216,N_1906,N_1745);
nand U2217 (N_2217,N_1612,N_1978);
or U2218 (N_2218,N_1572,N_1782);
nor U2219 (N_2219,N_1854,N_1719);
nand U2220 (N_2220,N_1710,N_1706);
nand U2221 (N_2221,N_1877,N_1784);
nor U2222 (N_2222,N_1647,N_1654);
and U2223 (N_2223,N_1691,N_1602);
or U2224 (N_2224,N_1714,N_1840);
nand U2225 (N_2225,N_1712,N_1804);
nor U2226 (N_2226,N_1669,N_1515);
or U2227 (N_2227,N_1866,N_1871);
or U2228 (N_2228,N_1813,N_1762);
nor U2229 (N_2229,N_1942,N_1895);
and U2230 (N_2230,N_1542,N_1925);
or U2231 (N_2231,N_1832,N_1611);
and U2232 (N_2232,N_1649,N_1615);
nand U2233 (N_2233,N_1764,N_1576);
and U2234 (N_2234,N_1980,N_1988);
or U2235 (N_2235,N_1688,N_1852);
nand U2236 (N_2236,N_1646,N_1629);
and U2237 (N_2237,N_1916,N_1563);
nand U2238 (N_2238,N_1805,N_1575);
or U2239 (N_2239,N_1983,N_1809);
nand U2240 (N_2240,N_1790,N_1825);
or U2241 (N_2241,N_1803,N_1662);
nor U2242 (N_2242,N_1713,N_1923);
or U2243 (N_2243,N_1570,N_1748);
nand U2244 (N_2244,N_1555,N_1972);
xnor U2245 (N_2245,N_1839,N_1939);
nor U2246 (N_2246,N_1997,N_1728);
nor U2247 (N_2247,N_1711,N_1686);
and U2248 (N_2248,N_1707,N_1739);
and U2249 (N_2249,N_1878,N_1557);
nor U2250 (N_2250,N_1579,N_1527);
and U2251 (N_2251,N_1523,N_1871);
nor U2252 (N_2252,N_1653,N_1981);
or U2253 (N_2253,N_1619,N_1617);
nand U2254 (N_2254,N_1915,N_1900);
nor U2255 (N_2255,N_1911,N_1763);
nor U2256 (N_2256,N_1651,N_1964);
nand U2257 (N_2257,N_1723,N_1530);
xnor U2258 (N_2258,N_1819,N_1808);
and U2259 (N_2259,N_1565,N_1549);
or U2260 (N_2260,N_1601,N_1757);
nand U2261 (N_2261,N_1779,N_1987);
and U2262 (N_2262,N_1981,N_1505);
or U2263 (N_2263,N_1518,N_1528);
nand U2264 (N_2264,N_1907,N_1584);
nand U2265 (N_2265,N_1512,N_1613);
or U2266 (N_2266,N_1973,N_1678);
and U2267 (N_2267,N_1514,N_1562);
and U2268 (N_2268,N_1930,N_1799);
and U2269 (N_2269,N_1868,N_1598);
or U2270 (N_2270,N_1658,N_1671);
or U2271 (N_2271,N_1677,N_1944);
and U2272 (N_2272,N_1980,N_1994);
nand U2273 (N_2273,N_1988,N_1892);
and U2274 (N_2274,N_1941,N_1944);
or U2275 (N_2275,N_1719,N_1956);
and U2276 (N_2276,N_1699,N_1548);
nand U2277 (N_2277,N_1783,N_1776);
or U2278 (N_2278,N_1669,N_1797);
and U2279 (N_2279,N_1872,N_1833);
and U2280 (N_2280,N_1716,N_1605);
nand U2281 (N_2281,N_1754,N_1894);
nor U2282 (N_2282,N_1565,N_1822);
nor U2283 (N_2283,N_1797,N_1666);
nand U2284 (N_2284,N_1673,N_1886);
nor U2285 (N_2285,N_1548,N_1771);
and U2286 (N_2286,N_1500,N_1753);
nor U2287 (N_2287,N_1793,N_1550);
or U2288 (N_2288,N_1717,N_1654);
nand U2289 (N_2289,N_1688,N_1538);
and U2290 (N_2290,N_1526,N_1527);
nor U2291 (N_2291,N_1642,N_1680);
or U2292 (N_2292,N_1998,N_1800);
and U2293 (N_2293,N_1997,N_1673);
and U2294 (N_2294,N_1789,N_1853);
nand U2295 (N_2295,N_1734,N_1870);
nand U2296 (N_2296,N_1677,N_1900);
or U2297 (N_2297,N_1596,N_1964);
or U2298 (N_2298,N_1593,N_1803);
and U2299 (N_2299,N_1677,N_1803);
nor U2300 (N_2300,N_1773,N_1813);
and U2301 (N_2301,N_1774,N_1694);
or U2302 (N_2302,N_1648,N_1900);
nor U2303 (N_2303,N_1877,N_1969);
nand U2304 (N_2304,N_1662,N_1538);
or U2305 (N_2305,N_1683,N_1679);
nor U2306 (N_2306,N_1657,N_1526);
nor U2307 (N_2307,N_1615,N_1956);
nand U2308 (N_2308,N_1747,N_1505);
and U2309 (N_2309,N_1754,N_1503);
or U2310 (N_2310,N_1873,N_1622);
nor U2311 (N_2311,N_1580,N_1670);
nand U2312 (N_2312,N_1631,N_1889);
or U2313 (N_2313,N_1918,N_1592);
nand U2314 (N_2314,N_1944,N_1878);
and U2315 (N_2315,N_1664,N_1745);
nor U2316 (N_2316,N_1525,N_1823);
nand U2317 (N_2317,N_1613,N_1902);
nand U2318 (N_2318,N_1875,N_1893);
nand U2319 (N_2319,N_1954,N_1581);
and U2320 (N_2320,N_1931,N_1787);
and U2321 (N_2321,N_1873,N_1530);
or U2322 (N_2322,N_1515,N_1966);
nand U2323 (N_2323,N_1957,N_1504);
and U2324 (N_2324,N_1592,N_1991);
and U2325 (N_2325,N_1777,N_1625);
nand U2326 (N_2326,N_1687,N_1755);
or U2327 (N_2327,N_1864,N_1703);
nand U2328 (N_2328,N_1578,N_1957);
nor U2329 (N_2329,N_1906,N_1549);
nor U2330 (N_2330,N_1510,N_1711);
nand U2331 (N_2331,N_1774,N_1541);
or U2332 (N_2332,N_1838,N_1689);
nand U2333 (N_2333,N_1551,N_1999);
nor U2334 (N_2334,N_1944,N_1751);
nor U2335 (N_2335,N_1574,N_1643);
and U2336 (N_2336,N_1802,N_1866);
or U2337 (N_2337,N_1561,N_1529);
nand U2338 (N_2338,N_1563,N_1972);
nand U2339 (N_2339,N_1716,N_1756);
and U2340 (N_2340,N_1650,N_1897);
and U2341 (N_2341,N_1541,N_1942);
nor U2342 (N_2342,N_1942,N_1576);
nand U2343 (N_2343,N_1916,N_1527);
nor U2344 (N_2344,N_1684,N_1607);
nand U2345 (N_2345,N_1920,N_1854);
nor U2346 (N_2346,N_1831,N_1815);
nor U2347 (N_2347,N_1686,N_1611);
nand U2348 (N_2348,N_1690,N_1651);
nor U2349 (N_2349,N_1911,N_1904);
and U2350 (N_2350,N_1933,N_1594);
nand U2351 (N_2351,N_1590,N_1683);
or U2352 (N_2352,N_1961,N_1820);
or U2353 (N_2353,N_1735,N_1673);
and U2354 (N_2354,N_1684,N_1763);
xnor U2355 (N_2355,N_1895,N_1735);
and U2356 (N_2356,N_1890,N_1733);
and U2357 (N_2357,N_1847,N_1605);
nand U2358 (N_2358,N_1526,N_1549);
and U2359 (N_2359,N_1564,N_1898);
nand U2360 (N_2360,N_1551,N_1766);
and U2361 (N_2361,N_1698,N_1813);
nor U2362 (N_2362,N_1885,N_1857);
nand U2363 (N_2363,N_1990,N_1649);
nand U2364 (N_2364,N_1524,N_1717);
or U2365 (N_2365,N_1716,N_1552);
nor U2366 (N_2366,N_1506,N_1617);
nand U2367 (N_2367,N_1725,N_1515);
and U2368 (N_2368,N_1692,N_1777);
nand U2369 (N_2369,N_1671,N_1535);
nand U2370 (N_2370,N_1619,N_1596);
nand U2371 (N_2371,N_1605,N_1512);
or U2372 (N_2372,N_1691,N_1770);
or U2373 (N_2373,N_1545,N_1598);
or U2374 (N_2374,N_1802,N_1776);
or U2375 (N_2375,N_1769,N_1871);
and U2376 (N_2376,N_1630,N_1844);
and U2377 (N_2377,N_1694,N_1868);
and U2378 (N_2378,N_1663,N_1589);
and U2379 (N_2379,N_1602,N_1827);
nor U2380 (N_2380,N_1774,N_1941);
nand U2381 (N_2381,N_1601,N_1835);
nand U2382 (N_2382,N_1636,N_1933);
nand U2383 (N_2383,N_1736,N_1580);
nand U2384 (N_2384,N_1597,N_1763);
nand U2385 (N_2385,N_1852,N_1733);
nor U2386 (N_2386,N_1700,N_1764);
and U2387 (N_2387,N_1656,N_1639);
or U2388 (N_2388,N_1829,N_1547);
nand U2389 (N_2389,N_1746,N_1610);
nand U2390 (N_2390,N_1694,N_1568);
nor U2391 (N_2391,N_1859,N_1722);
nor U2392 (N_2392,N_1588,N_1593);
nand U2393 (N_2393,N_1513,N_1617);
and U2394 (N_2394,N_1630,N_1745);
nand U2395 (N_2395,N_1599,N_1935);
xor U2396 (N_2396,N_1623,N_1605);
or U2397 (N_2397,N_1746,N_1762);
and U2398 (N_2398,N_1584,N_1619);
or U2399 (N_2399,N_1619,N_1542);
nand U2400 (N_2400,N_1727,N_1973);
nand U2401 (N_2401,N_1779,N_1606);
and U2402 (N_2402,N_1674,N_1788);
or U2403 (N_2403,N_1658,N_1684);
and U2404 (N_2404,N_1730,N_1760);
or U2405 (N_2405,N_1697,N_1859);
nand U2406 (N_2406,N_1755,N_1882);
nor U2407 (N_2407,N_1591,N_1776);
or U2408 (N_2408,N_1738,N_1783);
nand U2409 (N_2409,N_1520,N_1899);
nand U2410 (N_2410,N_1762,N_1754);
nand U2411 (N_2411,N_1751,N_1899);
or U2412 (N_2412,N_1680,N_1603);
and U2413 (N_2413,N_1793,N_1778);
and U2414 (N_2414,N_1591,N_1706);
nor U2415 (N_2415,N_1854,N_1900);
nor U2416 (N_2416,N_1572,N_1902);
nor U2417 (N_2417,N_1500,N_1577);
and U2418 (N_2418,N_1970,N_1914);
nor U2419 (N_2419,N_1949,N_1545);
nor U2420 (N_2420,N_1908,N_1874);
or U2421 (N_2421,N_1548,N_1592);
or U2422 (N_2422,N_1523,N_1914);
or U2423 (N_2423,N_1674,N_1845);
and U2424 (N_2424,N_1880,N_1679);
nand U2425 (N_2425,N_1747,N_1995);
and U2426 (N_2426,N_1704,N_1531);
or U2427 (N_2427,N_1714,N_1979);
or U2428 (N_2428,N_1631,N_1635);
and U2429 (N_2429,N_1701,N_1645);
or U2430 (N_2430,N_1670,N_1874);
and U2431 (N_2431,N_1797,N_1623);
or U2432 (N_2432,N_1859,N_1961);
or U2433 (N_2433,N_1553,N_1536);
or U2434 (N_2434,N_1991,N_1519);
and U2435 (N_2435,N_1836,N_1690);
nor U2436 (N_2436,N_1715,N_1709);
or U2437 (N_2437,N_1526,N_1923);
nand U2438 (N_2438,N_1573,N_1758);
and U2439 (N_2439,N_1949,N_1555);
nor U2440 (N_2440,N_1886,N_1753);
and U2441 (N_2441,N_1837,N_1818);
nor U2442 (N_2442,N_1959,N_1913);
or U2443 (N_2443,N_1940,N_1731);
and U2444 (N_2444,N_1904,N_1648);
and U2445 (N_2445,N_1818,N_1699);
and U2446 (N_2446,N_1792,N_1744);
and U2447 (N_2447,N_1643,N_1952);
nand U2448 (N_2448,N_1689,N_1526);
nor U2449 (N_2449,N_1825,N_1788);
nand U2450 (N_2450,N_1911,N_1908);
nand U2451 (N_2451,N_1903,N_1682);
nand U2452 (N_2452,N_1577,N_1839);
nand U2453 (N_2453,N_1982,N_1695);
and U2454 (N_2454,N_1955,N_1889);
and U2455 (N_2455,N_1560,N_1679);
nand U2456 (N_2456,N_1957,N_1691);
or U2457 (N_2457,N_1851,N_1668);
and U2458 (N_2458,N_1655,N_1588);
and U2459 (N_2459,N_1950,N_1503);
nand U2460 (N_2460,N_1769,N_1654);
and U2461 (N_2461,N_1540,N_1613);
nand U2462 (N_2462,N_1871,N_1553);
and U2463 (N_2463,N_1501,N_1949);
nand U2464 (N_2464,N_1641,N_1696);
nand U2465 (N_2465,N_1846,N_1933);
and U2466 (N_2466,N_1538,N_1531);
nor U2467 (N_2467,N_1511,N_1669);
nor U2468 (N_2468,N_1677,N_1767);
nor U2469 (N_2469,N_1933,N_1881);
nand U2470 (N_2470,N_1614,N_1509);
and U2471 (N_2471,N_1948,N_1710);
and U2472 (N_2472,N_1909,N_1630);
nor U2473 (N_2473,N_1604,N_1694);
nand U2474 (N_2474,N_1645,N_1536);
or U2475 (N_2475,N_1975,N_1542);
nand U2476 (N_2476,N_1537,N_1993);
nor U2477 (N_2477,N_1810,N_1566);
nand U2478 (N_2478,N_1506,N_1912);
nor U2479 (N_2479,N_1889,N_1526);
nand U2480 (N_2480,N_1856,N_1517);
and U2481 (N_2481,N_1670,N_1893);
and U2482 (N_2482,N_1654,N_1547);
or U2483 (N_2483,N_1808,N_1549);
and U2484 (N_2484,N_1866,N_1570);
and U2485 (N_2485,N_1506,N_1630);
nor U2486 (N_2486,N_1703,N_1796);
or U2487 (N_2487,N_1661,N_1579);
or U2488 (N_2488,N_1803,N_1833);
nand U2489 (N_2489,N_1690,N_1758);
and U2490 (N_2490,N_1600,N_1848);
or U2491 (N_2491,N_1876,N_1976);
nand U2492 (N_2492,N_1695,N_1652);
nand U2493 (N_2493,N_1614,N_1765);
nor U2494 (N_2494,N_1789,N_1683);
and U2495 (N_2495,N_1780,N_1915);
nor U2496 (N_2496,N_1620,N_1699);
and U2497 (N_2497,N_1769,N_1859);
and U2498 (N_2498,N_1592,N_1721);
or U2499 (N_2499,N_1698,N_1816);
or U2500 (N_2500,N_2385,N_2284);
and U2501 (N_2501,N_2414,N_2452);
and U2502 (N_2502,N_2336,N_2410);
nor U2503 (N_2503,N_2474,N_2369);
nand U2504 (N_2504,N_2015,N_2224);
and U2505 (N_2505,N_2008,N_2364);
or U2506 (N_2506,N_2132,N_2363);
or U2507 (N_2507,N_2466,N_2416);
nor U2508 (N_2508,N_2136,N_2139);
nand U2509 (N_2509,N_2433,N_2087);
nand U2510 (N_2510,N_2333,N_2248);
nand U2511 (N_2511,N_2066,N_2275);
or U2512 (N_2512,N_2358,N_2243);
and U2513 (N_2513,N_2396,N_2258);
and U2514 (N_2514,N_2187,N_2431);
or U2515 (N_2515,N_2437,N_2272);
or U2516 (N_2516,N_2372,N_2023);
nand U2517 (N_2517,N_2189,N_2121);
or U2518 (N_2518,N_2122,N_2293);
and U2519 (N_2519,N_2260,N_2482);
or U2520 (N_2520,N_2063,N_2062);
and U2521 (N_2521,N_2150,N_2216);
or U2522 (N_2522,N_2083,N_2427);
xnor U2523 (N_2523,N_2283,N_2404);
and U2524 (N_2524,N_2445,N_2027);
nor U2525 (N_2525,N_2418,N_2072);
nor U2526 (N_2526,N_2315,N_2355);
and U2527 (N_2527,N_2463,N_2135);
and U2528 (N_2528,N_2003,N_2183);
nand U2529 (N_2529,N_2324,N_2126);
and U2530 (N_2530,N_2245,N_2370);
or U2531 (N_2531,N_2421,N_2185);
and U2532 (N_2532,N_2460,N_2097);
and U2533 (N_2533,N_2093,N_2158);
nand U2534 (N_2534,N_2326,N_2345);
xnor U2535 (N_2535,N_2018,N_2312);
nand U2536 (N_2536,N_2049,N_2422);
or U2537 (N_2537,N_2367,N_2264);
nand U2538 (N_2538,N_2115,N_2134);
or U2539 (N_2539,N_2222,N_2489);
or U2540 (N_2540,N_2397,N_2174);
nand U2541 (N_2541,N_2068,N_2065);
nor U2542 (N_2542,N_2137,N_2035);
and U2543 (N_2543,N_2365,N_2111);
and U2544 (N_2544,N_2025,N_2221);
or U2545 (N_2545,N_2057,N_2259);
nor U2546 (N_2546,N_2170,N_2037);
nor U2547 (N_2547,N_2079,N_2107);
nor U2548 (N_2548,N_2420,N_2000);
or U2549 (N_2549,N_2007,N_2231);
nor U2550 (N_2550,N_2419,N_2261);
and U2551 (N_2551,N_2119,N_2468);
nor U2552 (N_2552,N_2086,N_2105);
nor U2553 (N_2553,N_2038,N_2471);
and U2554 (N_2554,N_2123,N_2288);
and U2555 (N_2555,N_2329,N_2267);
nand U2556 (N_2556,N_2251,N_2432);
nand U2557 (N_2557,N_2467,N_2186);
nor U2558 (N_2558,N_2456,N_2014);
and U2559 (N_2559,N_2010,N_2465);
nor U2560 (N_2560,N_2043,N_2378);
nand U2561 (N_2561,N_2127,N_2314);
and U2562 (N_2562,N_2498,N_2444);
and U2563 (N_2563,N_2292,N_2320);
or U2564 (N_2564,N_2045,N_2156);
nand U2565 (N_2565,N_2099,N_2149);
nand U2566 (N_2566,N_2110,N_2178);
or U2567 (N_2567,N_2476,N_2411);
and U2568 (N_2568,N_2446,N_2250);
or U2569 (N_2569,N_2439,N_2067);
nor U2570 (N_2570,N_2484,N_2206);
nand U2571 (N_2571,N_2096,N_2005);
nand U2572 (N_2572,N_2453,N_2140);
and U2573 (N_2573,N_2181,N_2021);
nand U2574 (N_2574,N_2071,N_2047);
or U2575 (N_2575,N_2169,N_2374);
nor U2576 (N_2576,N_2253,N_2337);
or U2577 (N_2577,N_2227,N_2328);
or U2578 (N_2578,N_2196,N_2348);
nand U2579 (N_2579,N_2294,N_2167);
or U2580 (N_2580,N_2249,N_2212);
or U2581 (N_2581,N_2070,N_2274);
nor U2582 (N_2582,N_2308,N_2303);
and U2583 (N_2583,N_2076,N_2226);
nor U2584 (N_2584,N_2492,N_2472);
nand U2585 (N_2585,N_2210,N_2089);
nand U2586 (N_2586,N_2331,N_2017);
and U2587 (N_2587,N_2384,N_2192);
and U2588 (N_2588,N_2113,N_2350);
nor U2589 (N_2589,N_2461,N_2074);
or U2590 (N_2590,N_2151,N_2321);
and U2591 (N_2591,N_2393,N_2050);
nor U2592 (N_2592,N_2166,N_2114);
or U2593 (N_2593,N_2059,N_2031);
xnor U2594 (N_2594,N_2310,N_2408);
nor U2595 (N_2595,N_2495,N_2116);
nor U2596 (N_2596,N_2297,N_2488);
and U2597 (N_2597,N_2060,N_2399);
or U2598 (N_2598,N_2028,N_2268);
or U2599 (N_2599,N_2041,N_2285);
and U2600 (N_2600,N_2269,N_2034);
nor U2601 (N_2601,N_2327,N_2217);
and U2602 (N_2602,N_2190,N_2478);
nor U2603 (N_2603,N_2128,N_2332);
or U2604 (N_2604,N_2039,N_2161);
nand U2605 (N_2605,N_2090,N_2030);
and U2606 (N_2606,N_2207,N_2413);
or U2607 (N_2607,N_2475,N_2032);
nand U2608 (N_2608,N_2276,N_2145);
nor U2609 (N_2609,N_2202,N_2163);
or U2610 (N_2610,N_2295,N_2082);
nand U2611 (N_2611,N_2302,N_2106);
or U2612 (N_2612,N_2496,N_2424);
and U2613 (N_2613,N_2152,N_2219);
and U2614 (N_2614,N_2490,N_2241);
or U2615 (N_2615,N_2088,N_2386);
or U2616 (N_2616,N_2485,N_2254);
nor U2617 (N_2617,N_2098,N_2448);
nor U2618 (N_2618,N_2359,N_2233);
nand U2619 (N_2619,N_2442,N_2198);
or U2620 (N_2620,N_2040,N_2434);
nand U2621 (N_2621,N_2279,N_2204);
xnor U2622 (N_2622,N_2200,N_2366);
or U2623 (N_2623,N_2343,N_2335);
or U2624 (N_2624,N_2316,N_2154);
or U2625 (N_2625,N_2338,N_2290);
nor U2626 (N_2626,N_2429,N_2497);
nand U2627 (N_2627,N_2022,N_2201);
and U2628 (N_2628,N_2470,N_2360);
xor U2629 (N_2629,N_2373,N_2454);
and U2630 (N_2630,N_2375,N_2133);
nand U2631 (N_2631,N_2462,N_2401);
nand U2632 (N_2632,N_2077,N_2441);
or U2633 (N_2633,N_2347,N_2125);
xor U2634 (N_2634,N_2148,N_2230);
or U2635 (N_2635,N_2138,N_2376);
and U2636 (N_2636,N_2438,N_2277);
or U2637 (N_2637,N_2271,N_2199);
xnor U2638 (N_2638,N_2255,N_2313);
nor U2639 (N_2639,N_2016,N_2412);
nand U2640 (N_2640,N_2120,N_2353);
nand U2641 (N_2641,N_2346,N_2162);
and U2642 (N_2642,N_2341,N_2457);
and U2643 (N_2643,N_2012,N_2405);
nor U2644 (N_2644,N_2240,N_2487);
and U2645 (N_2645,N_2415,N_2104);
nor U2646 (N_2646,N_2085,N_2307);
or U2647 (N_2647,N_2131,N_2215);
or U2648 (N_2648,N_2262,N_2426);
nor U2649 (N_2649,N_2208,N_2499);
nand U2650 (N_2650,N_2054,N_2402);
or U2651 (N_2651,N_2403,N_2001);
nand U2652 (N_2652,N_2141,N_2286);
or U2653 (N_2653,N_2306,N_2112);
or U2654 (N_2654,N_2371,N_2118);
and U2655 (N_2655,N_2213,N_2425);
and U2656 (N_2656,N_2362,N_2390);
and U2657 (N_2657,N_2298,N_2052);
or U2658 (N_2658,N_2195,N_2319);
and U2659 (N_2659,N_2340,N_2211);
xor U2660 (N_2660,N_2361,N_2400);
nor U2661 (N_2661,N_2029,N_2091);
nor U2662 (N_2662,N_2246,N_2483);
nand U2663 (N_2663,N_2435,N_2182);
nand U2664 (N_2664,N_2289,N_2389);
or U2665 (N_2665,N_2130,N_2352);
nor U2666 (N_2666,N_2301,N_2069);
or U2667 (N_2667,N_2173,N_2278);
or U2668 (N_2668,N_2299,N_2330);
nand U2669 (N_2669,N_2191,N_2282);
and U2670 (N_2670,N_2334,N_2159);
nand U2671 (N_2671,N_2242,N_2160);
or U2672 (N_2672,N_2381,N_2339);
nand U2673 (N_2673,N_2322,N_2354);
nor U2674 (N_2674,N_2394,N_2257);
nor U2675 (N_2675,N_2270,N_2477);
or U2676 (N_2676,N_2153,N_2019);
or U2677 (N_2677,N_2406,N_2236);
or U2678 (N_2678,N_2124,N_2232);
and U2679 (N_2679,N_2046,N_2229);
and U2680 (N_2680,N_2117,N_2146);
nand U2681 (N_2681,N_2417,N_2342);
nor U2682 (N_2682,N_2398,N_2423);
and U2683 (N_2683,N_2024,N_2493);
nor U2684 (N_2684,N_2458,N_2225);
and U2685 (N_2685,N_2180,N_2430);
nor U2686 (N_2686,N_2383,N_2256);
nor U2687 (N_2687,N_2092,N_2428);
nand U2688 (N_2688,N_2237,N_2479);
nand U2689 (N_2689,N_2193,N_2252);
nor U2690 (N_2690,N_2380,N_2064);
and U2691 (N_2691,N_2317,N_2094);
and U2692 (N_2692,N_2291,N_2026);
nor U2693 (N_2693,N_2392,N_2450);
or U2694 (N_2694,N_2377,N_2436);
xnor U2695 (N_2695,N_2443,N_2395);
nand U2696 (N_2696,N_2020,N_2184);
nand U2697 (N_2697,N_2002,N_2033);
nor U2698 (N_2698,N_2214,N_2387);
and U2699 (N_2699,N_2061,N_2265);
or U2700 (N_2700,N_2177,N_2056);
nor U2701 (N_2701,N_2318,N_2388);
nor U2702 (N_2702,N_2351,N_2147);
and U2703 (N_2703,N_2349,N_2247);
nand U2704 (N_2704,N_2281,N_2220);
and U2705 (N_2705,N_2244,N_2011);
and U2706 (N_2706,N_2391,N_2304);
and U2707 (N_2707,N_2055,N_2473);
or U2708 (N_2708,N_2081,N_2409);
or U2709 (N_2709,N_2469,N_2382);
nor U2710 (N_2710,N_2172,N_2036);
and U2711 (N_2711,N_2013,N_2325);
nor U2712 (N_2712,N_2323,N_2168);
nand U2713 (N_2713,N_2356,N_2491);
xnor U2714 (N_2714,N_2203,N_2205);
nor U2715 (N_2715,N_2480,N_2287);
and U2716 (N_2716,N_2440,N_2143);
nand U2717 (N_2717,N_2078,N_2309);
and U2718 (N_2718,N_2368,N_2464);
and U2719 (N_2719,N_2379,N_2494);
nor U2720 (N_2720,N_2053,N_2486);
and U2721 (N_2721,N_2108,N_2238);
and U2722 (N_2722,N_2235,N_2004);
nand U2723 (N_2723,N_2044,N_2175);
nand U2724 (N_2724,N_2009,N_2157);
nor U2725 (N_2725,N_2459,N_2084);
nand U2726 (N_2726,N_2194,N_2407);
nor U2727 (N_2727,N_2103,N_2109);
nor U2728 (N_2728,N_2239,N_2455);
or U2729 (N_2729,N_2095,N_2197);
or U2730 (N_2730,N_2042,N_2129);
xor U2731 (N_2731,N_2051,N_2357);
nor U2732 (N_2732,N_2080,N_2209);
or U2733 (N_2733,N_2100,N_2142);
nand U2734 (N_2734,N_2481,N_2273);
nor U2735 (N_2735,N_2048,N_2218);
nor U2736 (N_2736,N_2058,N_2073);
and U2737 (N_2737,N_2102,N_2171);
nor U2738 (N_2738,N_2311,N_2228);
or U2739 (N_2739,N_2144,N_2263);
nor U2740 (N_2740,N_2296,N_2101);
and U2741 (N_2741,N_2449,N_2179);
or U2742 (N_2742,N_2165,N_2300);
nand U2743 (N_2743,N_2223,N_2164);
and U2744 (N_2744,N_2305,N_2234);
nand U2745 (N_2745,N_2447,N_2266);
and U2746 (N_2746,N_2075,N_2176);
and U2747 (N_2747,N_2006,N_2344);
and U2748 (N_2748,N_2451,N_2155);
and U2749 (N_2749,N_2280,N_2188);
and U2750 (N_2750,N_2244,N_2183);
and U2751 (N_2751,N_2307,N_2135);
and U2752 (N_2752,N_2051,N_2223);
nand U2753 (N_2753,N_2361,N_2037);
or U2754 (N_2754,N_2342,N_2378);
nand U2755 (N_2755,N_2145,N_2330);
and U2756 (N_2756,N_2486,N_2064);
nand U2757 (N_2757,N_2348,N_2177);
or U2758 (N_2758,N_2324,N_2178);
or U2759 (N_2759,N_2352,N_2062);
nand U2760 (N_2760,N_2177,N_2265);
or U2761 (N_2761,N_2355,N_2051);
nand U2762 (N_2762,N_2094,N_2289);
nor U2763 (N_2763,N_2418,N_2180);
nand U2764 (N_2764,N_2391,N_2127);
or U2765 (N_2765,N_2026,N_2125);
nand U2766 (N_2766,N_2185,N_2243);
and U2767 (N_2767,N_2474,N_2048);
and U2768 (N_2768,N_2413,N_2201);
and U2769 (N_2769,N_2155,N_2255);
nor U2770 (N_2770,N_2402,N_2094);
nand U2771 (N_2771,N_2300,N_2138);
and U2772 (N_2772,N_2175,N_2321);
nand U2773 (N_2773,N_2216,N_2249);
nand U2774 (N_2774,N_2204,N_2374);
and U2775 (N_2775,N_2129,N_2320);
or U2776 (N_2776,N_2328,N_2215);
or U2777 (N_2777,N_2277,N_2383);
and U2778 (N_2778,N_2391,N_2256);
or U2779 (N_2779,N_2230,N_2194);
nand U2780 (N_2780,N_2417,N_2495);
nand U2781 (N_2781,N_2465,N_2380);
and U2782 (N_2782,N_2114,N_2420);
nand U2783 (N_2783,N_2076,N_2384);
or U2784 (N_2784,N_2457,N_2090);
nand U2785 (N_2785,N_2001,N_2458);
or U2786 (N_2786,N_2079,N_2364);
nor U2787 (N_2787,N_2431,N_2242);
nand U2788 (N_2788,N_2211,N_2427);
nor U2789 (N_2789,N_2188,N_2479);
and U2790 (N_2790,N_2154,N_2215);
nor U2791 (N_2791,N_2186,N_2033);
and U2792 (N_2792,N_2170,N_2254);
nor U2793 (N_2793,N_2178,N_2315);
nor U2794 (N_2794,N_2336,N_2192);
nor U2795 (N_2795,N_2292,N_2305);
or U2796 (N_2796,N_2482,N_2309);
nand U2797 (N_2797,N_2438,N_2177);
nor U2798 (N_2798,N_2322,N_2274);
and U2799 (N_2799,N_2060,N_2180);
nand U2800 (N_2800,N_2329,N_2153);
or U2801 (N_2801,N_2445,N_2289);
nand U2802 (N_2802,N_2256,N_2087);
nand U2803 (N_2803,N_2106,N_2048);
nand U2804 (N_2804,N_2376,N_2487);
and U2805 (N_2805,N_2412,N_2486);
nand U2806 (N_2806,N_2114,N_2381);
nor U2807 (N_2807,N_2133,N_2360);
nand U2808 (N_2808,N_2071,N_2330);
and U2809 (N_2809,N_2047,N_2029);
nand U2810 (N_2810,N_2198,N_2111);
nand U2811 (N_2811,N_2405,N_2209);
or U2812 (N_2812,N_2119,N_2369);
and U2813 (N_2813,N_2464,N_2329);
and U2814 (N_2814,N_2032,N_2049);
nor U2815 (N_2815,N_2346,N_2484);
nor U2816 (N_2816,N_2327,N_2386);
nand U2817 (N_2817,N_2186,N_2115);
nand U2818 (N_2818,N_2343,N_2084);
nor U2819 (N_2819,N_2147,N_2499);
and U2820 (N_2820,N_2098,N_2425);
nand U2821 (N_2821,N_2486,N_2440);
nand U2822 (N_2822,N_2230,N_2155);
or U2823 (N_2823,N_2024,N_2049);
nand U2824 (N_2824,N_2030,N_2193);
nor U2825 (N_2825,N_2199,N_2053);
and U2826 (N_2826,N_2389,N_2048);
and U2827 (N_2827,N_2147,N_2328);
nor U2828 (N_2828,N_2030,N_2129);
or U2829 (N_2829,N_2273,N_2118);
or U2830 (N_2830,N_2036,N_2125);
or U2831 (N_2831,N_2390,N_2011);
or U2832 (N_2832,N_2185,N_2320);
or U2833 (N_2833,N_2005,N_2319);
nand U2834 (N_2834,N_2360,N_2108);
and U2835 (N_2835,N_2270,N_2326);
or U2836 (N_2836,N_2285,N_2373);
nand U2837 (N_2837,N_2131,N_2324);
or U2838 (N_2838,N_2247,N_2309);
or U2839 (N_2839,N_2221,N_2103);
and U2840 (N_2840,N_2328,N_2365);
or U2841 (N_2841,N_2186,N_2490);
nand U2842 (N_2842,N_2125,N_2309);
nand U2843 (N_2843,N_2328,N_2146);
nor U2844 (N_2844,N_2139,N_2218);
or U2845 (N_2845,N_2456,N_2190);
nor U2846 (N_2846,N_2078,N_2454);
nand U2847 (N_2847,N_2191,N_2048);
nand U2848 (N_2848,N_2309,N_2083);
nand U2849 (N_2849,N_2484,N_2360);
nor U2850 (N_2850,N_2288,N_2198);
nand U2851 (N_2851,N_2101,N_2490);
nor U2852 (N_2852,N_2173,N_2014);
nor U2853 (N_2853,N_2275,N_2038);
xnor U2854 (N_2854,N_2269,N_2261);
or U2855 (N_2855,N_2412,N_2420);
or U2856 (N_2856,N_2295,N_2065);
or U2857 (N_2857,N_2218,N_2150);
or U2858 (N_2858,N_2237,N_2264);
nand U2859 (N_2859,N_2016,N_2390);
nor U2860 (N_2860,N_2195,N_2018);
nor U2861 (N_2861,N_2297,N_2263);
and U2862 (N_2862,N_2104,N_2149);
nor U2863 (N_2863,N_2172,N_2032);
nand U2864 (N_2864,N_2000,N_2407);
and U2865 (N_2865,N_2052,N_2015);
and U2866 (N_2866,N_2015,N_2024);
and U2867 (N_2867,N_2399,N_2054);
and U2868 (N_2868,N_2082,N_2469);
and U2869 (N_2869,N_2437,N_2239);
and U2870 (N_2870,N_2378,N_2182);
nand U2871 (N_2871,N_2415,N_2099);
or U2872 (N_2872,N_2016,N_2398);
nor U2873 (N_2873,N_2419,N_2276);
or U2874 (N_2874,N_2259,N_2202);
nor U2875 (N_2875,N_2458,N_2286);
nand U2876 (N_2876,N_2028,N_2190);
and U2877 (N_2877,N_2214,N_2349);
nor U2878 (N_2878,N_2009,N_2199);
and U2879 (N_2879,N_2374,N_2030);
nor U2880 (N_2880,N_2137,N_2023);
nor U2881 (N_2881,N_2249,N_2423);
and U2882 (N_2882,N_2032,N_2298);
nand U2883 (N_2883,N_2272,N_2148);
and U2884 (N_2884,N_2026,N_2039);
and U2885 (N_2885,N_2043,N_2259);
and U2886 (N_2886,N_2479,N_2238);
xor U2887 (N_2887,N_2160,N_2496);
nand U2888 (N_2888,N_2060,N_2320);
nand U2889 (N_2889,N_2122,N_2175);
nor U2890 (N_2890,N_2310,N_2010);
and U2891 (N_2891,N_2177,N_2343);
or U2892 (N_2892,N_2172,N_2148);
nand U2893 (N_2893,N_2444,N_2084);
nand U2894 (N_2894,N_2428,N_2005);
nand U2895 (N_2895,N_2303,N_2003);
or U2896 (N_2896,N_2399,N_2468);
nor U2897 (N_2897,N_2166,N_2075);
and U2898 (N_2898,N_2270,N_2260);
nor U2899 (N_2899,N_2357,N_2287);
nor U2900 (N_2900,N_2397,N_2208);
or U2901 (N_2901,N_2345,N_2448);
and U2902 (N_2902,N_2086,N_2236);
nor U2903 (N_2903,N_2249,N_2450);
or U2904 (N_2904,N_2136,N_2296);
nand U2905 (N_2905,N_2197,N_2117);
and U2906 (N_2906,N_2294,N_2475);
and U2907 (N_2907,N_2335,N_2129);
or U2908 (N_2908,N_2095,N_2442);
nor U2909 (N_2909,N_2441,N_2057);
or U2910 (N_2910,N_2368,N_2292);
nand U2911 (N_2911,N_2081,N_2187);
or U2912 (N_2912,N_2230,N_2013);
nor U2913 (N_2913,N_2302,N_2184);
and U2914 (N_2914,N_2296,N_2026);
nor U2915 (N_2915,N_2196,N_2061);
nor U2916 (N_2916,N_2141,N_2183);
nor U2917 (N_2917,N_2284,N_2292);
nor U2918 (N_2918,N_2287,N_2446);
and U2919 (N_2919,N_2187,N_2458);
and U2920 (N_2920,N_2122,N_2266);
or U2921 (N_2921,N_2341,N_2047);
nor U2922 (N_2922,N_2108,N_2086);
and U2923 (N_2923,N_2030,N_2331);
nand U2924 (N_2924,N_2351,N_2274);
or U2925 (N_2925,N_2230,N_2358);
and U2926 (N_2926,N_2476,N_2395);
or U2927 (N_2927,N_2263,N_2137);
and U2928 (N_2928,N_2036,N_2051);
nand U2929 (N_2929,N_2031,N_2135);
nor U2930 (N_2930,N_2375,N_2274);
nor U2931 (N_2931,N_2296,N_2292);
nand U2932 (N_2932,N_2352,N_2080);
and U2933 (N_2933,N_2290,N_2170);
nand U2934 (N_2934,N_2216,N_2392);
nand U2935 (N_2935,N_2132,N_2307);
nand U2936 (N_2936,N_2188,N_2087);
nor U2937 (N_2937,N_2469,N_2296);
nand U2938 (N_2938,N_2331,N_2087);
nor U2939 (N_2939,N_2148,N_2017);
or U2940 (N_2940,N_2166,N_2359);
and U2941 (N_2941,N_2050,N_2145);
or U2942 (N_2942,N_2284,N_2013);
or U2943 (N_2943,N_2308,N_2340);
and U2944 (N_2944,N_2040,N_2469);
nor U2945 (N_2945,N_2310,N_2058);
nor U2946 (N_2946,N_2354,N_2129);
and U2947 (N_2947,N_2361,N_2105);
nor U2948 (N_2948,N_2131,N_2231);
or U2949 (N_2949,N_2114,N_2095);
and U2950 (N_2950,N_2215,N_2106);
and U2951 (N_2951,N_2122,N_2076);
and U2952 (N_2952,N_2062,N_2464);
nand U2953 (N_2953,N_2089,N_2100);
and U2954 (N_2954,N_2102,N_2390);
or U2955 (N_2955,N_2400,N_2273);
or U2956 (N_2956,N_2412,N_2177);
or U2957 (N_2957,N_2092,N_2041);
and U2958 (N_2958,N_2135,N_2256);
or U2959 (N_2959,N_2074,N_2218);
nand U2960 (N_2960,N_2258,N_2236);
nand U2961 (N_2961,N_2089,N_2326);
nand U2962 (N_2962,N_2047,N_2464);
nor U2963 (N_2963,N_2334,N_2109);
nand U2964 (N_2964,N_2135,N_2165);
and U2965 (N_2965,N_2081,N_2023);
nor U2966 (N_2966,N_2487,N_2095);
nor U2967 (N_2967,N_2224,N_2195);
and U2968 (N_2968,N_2078,N_2334);
and U2969 (N_2969,N_2403,N_2060);
and U2970 (N_2970,N_2434,N_2053);
and U2971 (N_2971,N_2280,N_2186);
nor U2972 (N_2972,N_2395,N_2328);
nor U2973 (N_2973,N_2192,N_2212);
and U2974 (N_2974,N_2157,N_2356);
or U2975 (N_2975,N_2344,N_2115);
and U2976 (N_2976,N_2217,N_2468);
nor U2977 (N_2977,N_2124,N_2343);
nor U2978 (N_2978,N_2467,N_2032);
nand U2979 (N_2979,N_2153,N_2468);
nand U2980 (N_2980,N_2014,N_2425);
nand U2981 (N_2981,N_2061,N_2286);
and U2982 (N_2982,N_2144,N_2185);
or U2983 (N_2983,N_2000,N_2333);
and U2984 (N_2984,N_2448,N_2033);
or U2985 (N_2985,N_2368,N_2080);
and U2986 (N_2986,N_2081,N_2059);
and U2987 (N_2987,N_2487,N_2293);
or U2988 (N_2988,N_2082,N_2481);
nand U2989 (N_2989,N_2262,N_2238);
nand U2990 (N_2990,N_2264,N_2434);
nor U2991 (N_2991,N_2282,N_2478);
or U2992 (N_2992,N_2036,N_2389);
or U2993 (N_2993,N_2362,N_2277);
or U2994 (N_2994,N_2196,N_2015);
nor U2995 (N_2995,N_2016,N_2174);
nor U2996 (N_2996,N_2161,N_2146);
nor U2997 (N_2997,N_2115,N_2415);
and U2998 (N_2998,N_2319,N_2382);
nor U2999 (N_2999,N_2031,N_2492);
and U3000 (N_3000,N_2639,N_2817);
nor U3001 (N_3001,N_2997,N_2716);
nor U3002 (N_3002,N_2891,N_2668);
or U3003 (N_3003,N_2543,N_2978);
or U3004 (N_3004,N_2772,N_2833);
nand U3005 (N_3005,N_2719,N_2987);
and U3006 (N_3006,N_2746,N_2641);
or U3007 (N_3007,N_2620,N_2724);
nand U3008 (N_3008,N_2600,N_2929);
nor U3009 (N_3009,N_2524,N_2819);
nand U3010 (N_3010,N_2725,N_2932);
or U3011 (N_3011,N_2921,N_2871);
or U3012 (N_3012,N_2553,N_2878);
and U3013 (N_3013,N_2736,N_2571);
nor U3014 (N_3014,N_2866,N_2988);
or U3015 (N_3015,N_2936,N_2615);
and U3016 (N_3016,N_2589,N_2516);
nand U3017 (N_3017,N_2959,N_2602);
or U3018 (N_3018,N_2836,N_2843);
nand U3019 (N_3019,N_2791,N_2768);
or U3020 (N_3020,N_2928,N_2701);
or U3021 (N_3021,N_2713,N_2554);
and U3022 (N_3022,N_2688,N_2609);
or U3023 (N_3023,N_2678,N_2755);
and U3024 (N_3024,N_2839,N_2662);
nor U3025 (N_3025,N_2650,N_2608);
or U3026 (N_3026,N_2606,N_2757);
nand U3027 (N_3027,N_2914,N_2631);
or U3028 (N_3028,N_2733,N_2872);
nor U3029 (N_3029,N_2756,N_2773);
and U3030 (N_3030,N_2656,N_2938);
or U3031 (N_3031,N_2953,N_2810);
and U3032 (N_3032,N_2663,N_2973);
or U3033 (N_3033,N_2889,N_2882);
and U3034 (N_3034,N_2677,N_2542);
nor U3035 (N_3035,N_2536,N_2984);
or U3036 (N_3036,N_2831,N_2949);
nand U3037 (N_3037,N_2751,N_2550);
or U3038 (N_3038,N_2657,N_2513);
and U3039 (N_3039,N_2961,N_2728);
nand U3040 (N_3040,N_2884,N_2937);
nand U3041 (N_3041,N_2560,N_2894);
nor U3042 (N_3042,N_2853,N_2703);
nor U3043 (N_3043,N_2888,N_2841);
and U3044 (N_3044,N_2775,N_2590);
nor U3045 (N_3045,N_2501,N_2748);
xor U3046 (N_3046,N_2999,N_2729);
nand U3047 (N_3047,N_2511,N_2507);
or U3048 (N_3048,N_2770,N_2634);
nand U3049 (N_3049,N_2582,N_2812);
nor U3050 (N_3050,N_2789,N_2707);
and U3051 (N_3051,N_2907,N_2750);
xnor U3052 (N_3052,N_2799,N_2925);
or U3053 (N_3053,N_2875,N_2869);
nor U3054 (N_3054,N_2783,N_2623);
and U3055 (N_3055,N_2911,N_2573);
nand U3056 (N_3056,N_2661,N_2964);
and U3057 (N_3057,N_2548,N_2752);
nor U3058 (N_3058,N_2519,N_2723);
and U3059 (N_3059,N_2722,N_2828);
or U3060 (N_3060,N_2718,N_2950);
and U3061 (N_3061,N_2682,N_2672);
nand U3062 (N_3062,N_2933,N_2976);
nand U3063 (N_3063,N_2568,N_2885);
nand U3064 (N_3064,N_2693,N_2525);
nand U3065 (N_3065,N_2850,N_2971);
or U3066 (N_3066,N_2919,N_2764);
or U3067 (N_3067,N_2655,N_2510);
nor U3068 (N_3068,N_2636,N_2537);
or U3069 (N_3069,N_2823,N_2689);
and U3070 (N_3070,N_2643,N_2813);
nor U3071 (N_3071,N_2526,N_2908);
nor U3072 (N_3072,N_2780,N_2967);
nand U3073 (N_3073,N_2998,N_2506);
nor U3074 (N_3074,N_2659,N_2956);
nand U3075 (N_3075,N_2981,N_2926);
nand U3076 (N_3076,N_2881,N_2801);
nor U3077 (N_3077,N_2691,N_2715);
or U3078 (N_3078,N_2972,N_2845);
or U3079 (N_3079,N_2766,N_2547);
or U3080 (N_3080,N_2979,N_2931);
and U3081 (N_3081,N_2962,N_2697);
and U3082 (N_3082,N_2555,N_2753);
nand U3083 (N_3083,N_2787,N_2735);
nand U3084 (N_3084,N_2565,N_2905);
and U3085 (N_3085,N_2534,N_2870);
nand U3086 (N_3086,N_2622,N_2581);
nand U3087 (N_3087,N_2915,N_2977);
or U3088 (N_3088,N_2821,N_2575);
nand U3089 (N_3089,N_2686,N_2637);
nor U3090 (N_3090,N_2818,N_2648);
nor U3091 (N_3091,N_2569,N_2879);
and U3092 (N_3092,N_2830,N_2610);
and U3093 (N_3093,N_2954,N_2876);
and U3094 (N_3094,N_2683,N_2788);
nand U3095 (N_3095,N_2579,N_2712);
and U3096 (N_3096,N_2690,N_2539);
or U3097 (N_3097,N_2795,N_2842);
and U3098 (N_3098,N_2939,N_2706);
and U3099 (N_3099,N_2771,N_2709);
nor U3100 (N_3100,N_2852,N_2518);
or U3101 (N_3101,N_2617,N_2708);
nand U3102 (N_3102,N_2647,N_2532);
or U3103 (N_3103,N_2503,N_2627);
or U3104 (N_3104,N_2613,N_2749);
nand U3105 (N_3105,N_2528,N_2629);
and U3106 (N_3106,N_2667,N_2523);
or U3107 (N_3107,N_2898,N_2996);
and U3108 (N_3108,N_2603,N_2796);
or U3109 (N_3109,N_2727,N_2500);
nor U3110 (N_3110,N_2734,N_2805);
and U3111 (N_3111,N_2957,N_2856);
nor U3112 (N_3112,N_2868,N_2761);
nand U3113 (N_3113,N_2598,N_2848);
and U3114 (N_3114,N_2562,N_2564);
nor U3115 (N_3115,N_2803,N_2990);
and U3116 (N_3116,N_2893,N_2759);
nand U3117 (N_3117,N_2694,N_2587);
nand U3118 (N_3118,N_2685,N_2807);
or U3119 (N_3119,N_2741,N_2873);
and U3120 (N_3120,N_2742,N_2567);
or U3121 (N_3121,N_2994,N_2530);
nor U3122 (N_3122,N_2858,N_2955);
nand U3123 (N_3123,N_2597,N_2861);
nand U3124 (N_3124,N_2737,N_2681);
nor U3125 (N_3125,N_2857,N_2664);
and U3126 (N_3126,N_2592,N_2561);
and U3127 (N_3127,N_2824,N_2776);
nand U3128 (N_3128,N_2515,N_2778);
nand U3129 (N_3129,N_2612,N_2696);
and U3130 (N_3130,N_2811,N_2774);
or U3131 (N_3131,N_2963,N_2566);
or U3132 (N_3132,N_2533,N_2863);
and U3133 (N_3133,N_2540,N_2784);
nor U3134 (N_3134,N_2654,N_2745);
or U3135 (N_3135,N_2621,N_2522);
nand U3136 (N_3136,N_2844,N_2945);
or U3137 (N_3137,N_2680,N_2546);
or U3138 (N_3138,N_2563,N_2529);
or U3139 (N_3139,N_2601,N_2779);
or U3140 (N_3140,N_2556,N_2765);
or U3141 (N_3141,N_2910,N_2509);
nand U3142 (N_3142,N_2816,N_2985);
nor U3143 (N_3143,N_2942,N_2760);
nand U3144 (N_3144,N_2611,N_2698);
nor U3145 (N_3145,N_2903,N_2767);
nor U3146 (N_3146,N_2923,N_2785);
nor U3147 (N_3147,N_2798,N_2895);
nand U3148 (N_3148,N_2640,N_2982);
nand U3149 (N_3149,N_2541,N_2671);
and U3150 (N_3150,N_2628,N_2531);
nand U3151 (N_3151,N_2820,N_2646);
nor U3152 (N_3152,N_2652,N_2580);
or U3153 (N_3153,N_2520,N_2952);
nor U3154 (N_3154,N_2808,N_2595);
or U3155 (N_3155,N_2782,N_2934);
and U3156 (N_3156,N_2904,N_2695);
nand U3157 (N_3157,N_2538,N_2585);
and U3158 (N_3158,N_2747,N_2890);
or U3159 (N_3159,N_2527,N_2702);
and U3160 (N_3160,N_2838,N_2653);
nand U3161 (N_3161,N_2545,N_2673);
or U3162 (N_3162,N_2699,N_2679);
and U3163 (N_3163,N_2966,N_2892);
and U3164 (N_3164,N_2607,N_2754);
nand U3165 (N_3165,N_2544,N_2577);
and U3166 (N_3166,N_2593,N_2710);
or U3167 (N_3167,N_2864,N_2815);
nand U3168 (N_3168,N_2944,N_2992);
and U3169 (N_3169,N_2576,N_2599);
or U3170 (N_3170,N_2794,N_2840);
or U3171 (N_3171,N_2744,N_2951);
nand U3172 (N_3172,N_2762,N_2887);
nand U3173 (N_3173,N_2670,N_2574);
or U3174 (N_3174,N_2551,N_2809);
or U3175 (N_3175,N_2993,N_2605);
and U3176 (N_3176,N_2584,N_2859);
and U3177 (N_3177,N_2714,N_2632);
and U3178 (N_3178,N_2941,N_2860);
nor U3179 (N_3179,N_2705,N_2827);
nor U3180 (N_3180,N_2717,N_2591);
and U3181 (N_3181,N_2829,N_2552);
nand U3182 (N_3182,N_2927,N_2974);
nor U3183 (N_3183,N_2880,N_2867);
or U3184 (N_3184,N_2658,N_2517);
or U3185 (N_3185,N_2638,N_2721);
nand U3186 (N_3186,N_2943,N_2665);
nor U3187 (N_3187,N_2630,N_2583);
or U3188 (N_3188,N_2797,N_2535);
nor U3189 (N_3189,N_2633,N_2916);
and U3190 (N_3190,N_2930,N_2660);
or U3191 (N_3191,N_2777,N_2902);
and U3192 (N_3192,N_2918,N_2559);
or U3193 (N_3193,N_2730,N_2849);
nor U3194 (N_3194,N_2970,N_2588);
and U3195 (N_3195,N_2624,N_2769);
nand U3196 (N_3196,N_2505,N_2825);
nor U3197 (N_3197,N_2557,N_2642);
or U3198 (N_3198,N_2897,N_2837);
nor U3199 (N_3199,N_2687,N_2983);
xnor U3200 (N_3200,N_2651,N_2674);
nor U3201 (N_3201,N_2645,N_2619);
or U3202 (N_3202,N_2899,N_2802);
and U3203 (N_3203,N_2558,N_2739);
or U3204 (N_3204,N_2800,N_2935);
and U3205 (N_3205,N_2684,N_2814);
or U3206 (N_3206,N_2675,N_2855);
nand U3207 (N_3207,N_2570,N_2906);
nand U3208 (N_3208,N_2521,N_2793);
nand U3209 (N_3209,N_2790,N_2854);
nor U3210 (N_3210,N_2991,N_2851);
nand U3211 (N_3211,N_2804,N_2958);
nor U3212 (N_3212,N_2711,N_2549);
and U3213 (N_3213,N_2865,N_2822);
nand U3214 (N_3214,N_2832,N_2578);
and U3215 (N_3215,N_2900,N_2572);
nand U3216 (N_3216,N_2912,N_2743);
or U3217 (N_3217,N_2763,N_2965);
nand U3218 (N_3218,N_2980,N_2704);
nand U3219 (N_3219,N_2738,N_2504);
and U3220 (N_3220,N_2896,N_2960);
or U3221 (N_3221,N_2986,N_2806);
nor U3222 (N_3222,N_2614,N_2995);
nand U3223 (N_3223,N_2975,N_2514);
nor U3224 (N_3224,N_2826,N_2901);
nor U3225 (N_3225,N_2834,N_2924);
nand U3226 (N_3226,N_2700,N_2626);
or U3227 (N_3227,N_2781,N_2669);
nor U3228 (N_3228,N_2594,N_2913);
nor U3229 (N_3229,N_2922,N_2874);
nor U3230 (N_3230,N_2940,N_2847);
xor U3231 (N_3231,N_2969,N_2596);
or U3232 (N_3232,N_2625,N_2846);
nor U3233 (N_3233,N_2635,N_2909);
nor U3234 (N_3234,N_2618,N_2726);
and U3235 (N_3235,N_2758,N_2644);
nor U3236 (N_3236,N_2968,N_2886);
nor U3237 (N_3237,N_2948,N_2731);
nand U3238 (N_3238,N_2989,N_2917);
or U3239 (N_3239,N_2740,N_2862);
nand U3240 (N_3240,N_2512,N_2502);
nand U3241 (N_3241,N_2586,N_2692);
and U3242 (N_3242,N_2649,N_2508);
nand U3243 (N_3243,N_2720,N_2616);
and U3244 (N_3244,N_2877,N_2883);
and U3245 (N_3245,N_2666,N_2946);
or U3246 (N_3246,N_2786,N_2835);
and U3247 (N_3247,N_2792,N_2676);
or U3248 (N_3248,N_2947,N_2604);
nor U3249 (N_3249,N_2920,N_2732);
or U3250 (N_3250,N_2570,N_2871);
and U3251 (N_3251,N_2706,N_2536);
or U3252 (N_3252,N_2588,N_2884);
and U3253 (N_3253,N_2674,N_2834);
nor U3254 (N_3254,N_2534,N_2940);
nor U3255 (N_3255,N_2556,N_2858);
nor U3256 (N_3256,N_2662,N_2960);
xnor U3257 (N_3257,N_2616,N_2588);
and U3258 (N_3258,N_2974,N_2538);
nor U3259 (N_3259,N_2745,N_2706);
and U3260 (N_3260,N_2716,N_2695);
nor U3261 (N_3261,N_2517,N_2803);
nor U3262 (N_3262,N_2522,N_2878);
and U3263 (N_3263,N_2708,N_2738);
and U3264 (N_3264,N_2962,N_2797);
or U3265 (N_3265,N_2701,N_2834);
nand U3266 (N_3266,N_2519,N_2967);
nor U3267 (N_3267,N_2900,N_2637);
nand U3268 (N_3268,N_2682,N_2633);
nand U3269 (N_3269,N_2720,N_2679);
nor U3270 (N_3270,N_2847,N_2529);
and U3271 (N_3271,N_2694,N_2571);
nor U3272 (N_3272,N_2551,N_2885);
nand U3273 (N_3273,N_2561,N_2890);
and U3274 (N_3274,N_2785,N_2961);
or U3275 (N_3275,N_2979,N_2625);
nor U3276 (N_3276,N_2723,N_2871);
nand U3277 (N_3277,N_2672,N_2614);
or U3278 (N_3278,N_2578,N_2623);
nand U3279 (N_3279,N_2881,N_2665);
nor U3280 (N_3280,N_2838,N_2948);
nand U3281 (N_3281,N_2585,N_2909);
and U3282 (N_3282,N_2772,N_2826);
nor U3283 (N_3283,N_2814,N_2782);
nor U3284 (N_3284,N_2883,N_2857);
nand U3285 (N_3285,N_2648,N_2578);
nor U3286 (N_3286,N_2717,N_2734);
or U3287 (N_3287,N_2921,N_2522);
or U3288 (N_3288,N_2894,N_2812);
nor U3289 (N_3289,N_2578,N_2973);
and U3290 (N_3290,N_2646,N_2549);
and U3291 (N_3291,N_2879,N_2761);
or U3292 (N_3292,N_2541,N_2902);
and U3293 (N_3293,N_2777,N_2515);
or U3294 (N_3294,N_2736,N_2868);
nor U3295 (N_3295,N_2529,N_2796);
nand U3296 (N_3296,N_2903,N_2847);
and U3297 (N_3297,N_2680,N_2792);
or U3298 (N_3298,N_2713,N_2660);
and U3299 (N_3299,N_2890,N_2793);
or U3300 (N_3300,N_2545,N_2904);
and U3301 (N_3301,N_2667,N_2735);
nand U3302 (N_3302,N_2977,N_2935);
or U3303 (N_3303,N_2509,N_2507);
and U3304 (N_3304,N_2830,N_2888);
or U3305 (N_3305,N_2985,N_2869);
or U3306 (N_3306,N_2842,N_2646);
and U3307 (N_3307,N_2505,N_2644);
xnor U3308 (N_3308,N_2637,N_2847);
or U3309 (N_3309,N_2739,N_2926);
and U3310 (N_3310,N_2731,N_2799);
or U3311 (N_3311,N_2519,N_2671);
or U3312 (N_3312,N_2772,N_2783);
nand U3313 (N_3313,N_2663,N_2771);
nor U3314 (N_3314,N_2934,N_2579);
and U3315 (N_3315,N_2731,N_2890);
nand U3316 (N_3316,N_2619,N_2904);
or U3317 (N_3317,N_2974,N_2946);
nand U3318 (N_3318,N_2658,N_2948);
nor U3319 (N_3319,N_2583,N_2795);
or U3320 (N_3320,N_2701,N_2707);
and U3321 (N_3321,N_2710,N_2723);
nand U3322 (N_3322,N_2506,N_2873);
nand U3323 (N_3323,N_2749,N_2828);
nand U3324 (N_3324,N_2664,N_2598);
or U3325 (N_3325,N_2933,N_2514);
nand U3326 (N_3326,N_2586,N_2905);
nand U3327 (N_3327,N_2922,N_2524);
nor U3328 (N_3328,N_2969,N_2526);
and U3329 (N_3329,N_2552,N_2518);
and U3330 (N_3330,N_2835,N_2526);
nand U3331 (N_3331,N_2529,N_2969);
or U3332 (N_3332,N_2756,N_2791);
or U3333 (N_3333,N_2662,N_2894);
xnor U3334 (N_3334,N_2738,N_2941);
and U3335 (N_3335,N_2965,N_2543);
or U3336 (N_3336,N_2894,N_2605);
and U3337 (N_3337,N_2502,N_2989);
or U3338 (N_3338,N_2519,N_2645);
nor U3339 (N_3339,N_2716,N_2995);
nor U3340 (N_3340,N_2606,N_2820);
or U3341 (N_3341,N_2699,N_2680);
nand U3342 (N_3342,N_2769,N_2963);
nor U3343 (N_3343,N_2615,N_2852);
or U3344 (N_3344,N_2835,N_2851);
and U3345 (N_3345,N_2592,N_2860);
nand U3346 (N_3346,N_2963,N_2616);
nor U3347 (N_3347,N_2861,N_2911);
or U3348 (N_3348,N_2996,N_2890);
and U3349 (N_3349,N_2708,N_2699);
or U3350 (N_3350,N_2573,N_2638);
and U3351 (N_3351,N_2797,N_2642);
nor U3352 (N_3352,N_2509,N_2788);
nand U3353 (N_3353,N_2650,N_2567);
and U3354 (N_3354,N_2780,N_2922);
and U3355 (N_3355,N_2683,N_2934);
nor U3356 (N_3356,N_2755,N_2577);
nand U3357 (N_3357,N_2658,N_2983);
and U3358 (N_3358,N_2965,N_2675);
nand U3359 (N_3359,N_2560,N_2803);
and U3360 (N_3360,N_2658,N_2684);
nand U3361 (N_3361,N_2849,N_2882);
or U3362 (N_3362,N_2735,N_2943);
nand U3363 (N_3363,N_2731,N_2875);
or U3364 (N_3364,N_2786,N_2944);
nand U3365 (N_3365,N_2611,N_2817);
nor U3366 (N_3366,N_2836,N_2501);
and U3367 (N_3367,N_2887,N_2812);
or U3368 (N_3368,N_2661,N_2738);
nor U3369 (N_3369,N_2600,N_2703);
nand U3370 (N_3370,N_2920,N_2947);
nand U3371 (N_3371,N_2727,N_2647);
nor U3372 (N_3372,N_2550,N_2655);
or U3373 (N_3373,N_2574,N_2709);
nor U3374 (N_3374,N_2642,N_2727);
and U3375 (N_3375,N_2966,N_2721);
or U3376 (N_3376,N_2738,N_2530);
nor U3377 (N_3377,N_2592,N_2687);
and U3378 (N_3378,N_2622,N_2981);
nor U3379 (N_3379,N_2778,N_2524);
nand U3380 (N_3380,N_2622,N_2972);
and U3381 (N_3381,N_2693,N_2698);
nand U3382 (N_3382,N_2627,N_2764);
nand U3383 (N_3383,N_2779,N_2886);
or U3384 (N_3384,N_2981,N_2939);
or U3385 (N_3385,N_2659,N_2992);
nand U3386 (N_3386,N_2710,N_2715);
nand U3387 (N_3387,N_2812,N_2668);
and U3388 (N_3388,N_2695,N_2881);
or U3389 (N_3389,N_2616,N_2847);
or U3390 (N_3390,N_2681,N_2695);
and U3391 (N_3391,N_2557,N_2684);
nand U3392 (N_3392,N_2723,N_2686);
and U3393 (N_3393,N_2830,N_2710);
and U3394 (N_3394,N_2807,N_2834);
or U3395 (N_3395,N_2857,N_2768);
and U3396 (N_3396,N_2936,N_2837);
or U3397 (N_3397,N_2551,N_2805);
nor U3398 (N_3398,N_2682,N_2898);
or U3399 (N_3399,N_2521,N_2518);
nor U3400 (N_3400,N_2781,N_2909);
nor U3401 (N_3401,N_2645,N_2962);
or U3402 (N_3402,N_2740,N_2994);
nand U3403 (N_3403,N_2522,N_2590);
and U3404 (N_3404,N_2576,N_2613);
and U3405 (N_3405,N_2645,N_2701);
nor U3406 (N_3406,N_2844,N_2993);
and U3407 (N_3407,N_2564,N_2653);
nor U3408 (N_3408,N_2934,N_2843);
and U3409 (N_3409,N_2501,N_2945);
and U3410 (N_3410,N_2846,N_2723);
nand U3411 (N_3411,N_2609,N_2647);
xnor U3412 (N_3412,N_2690,N_2927);
nand U3413 (N_3413,N_2635,N_2691);
and U3414 (N_3414,N_2500,N_2876);
nor U3415 (N_3415,N_2880,N_2970);
and U3416 (N_3416,N_2806,N_2620);
and U3417 (N_3417,N_2728,N_2595);
nor U3418 (N_3418,N_2662,N_2872);
or U3419 (N_3419,N_2820,N_2711);
nand U3420 (N_3420,N_2699,N_2855);
nand U3421 (N_3421,N_2872,N_2782);
nor U3422 (N_3422,N_2651,N_2535);
or U3423 (N_3423,N_2779,N_2966);
nor U3424 (N_3424,N_2815,N_2930);
or U3425 (N_3425,N_2604,N_2957);
and U3426 (N_3426,N_2756,N_2872);
nor U3427 (N_3427,N_2791,N_2950);
nor U3428 (N_3428,N_2806,N_2892);
and U3429 (N_3429,N_2629,N_2896);
nor U3430 (N_3430,N_2768,N_2514);
nand U3431 (N_3431,N_2927,N_2761);
nand U3432 (N_3432,N_2978,N_2531);
or U3433 (N_3433,N_2744,N_2743);
and U3434 (N_3434,N_2577,N_2771);
or U3435 (N_3435,N_2521,N_2933);
and U3436 (N_3436,N_2591,N_2975);
or U3437 (N_3437,N_2525,N_2999);
nor U3438 (N_3438,N_2941,N_2798);
or U3439 (N_3439,N_2793,N_2638);
nor U3440 (N_3440,N_2686,N_2818);
nor U3441 (N_3441,N_2621,N_2857);
and U3442 (N_3442,N_2881,N_2994);
nor U3443 (N_3443,N_2906,N_2868);
nand U3444 (N_3444,N_2839,N_2667);
or U3445 (N_3445,N_2977,N_2714);
nand U3446 (N_3446,N_2860,N_2970);
nor U3447 (N_3447,N_2800,N_2687);
or U3448 (N_3448,N_2509,N_2783);
or U3449 (N_3449,N_2877,N_2680);
or U3450 (N_3450,N_2991,N_2816);
and U3451 (N_3451,N_2533,N_2858);
and U3452 (N_3452,N_2960,N_2992);
and U3453 (N_3453,N_2580,N_2867);
or U3454 (N_3454,N_2858,N_2875);
nand U3455 (N_3455,N_2601,N_2995);
or U3456 (N_3456,N_2751,N_2634);
or U3457 (N_3457,N_2696,N_2516);
nor U3458 (N_3458,N_2569,N_2637);
nand U3459 (N_3459,N_2988,N_2819);
nor U3460 (N_3460,N_2741,N_2847);
nor U3461 (N_3461,N_2983,N_2672);
or U3462 (N_3462,N_2640,N_2653);
or U3463 (N_3463,N_2774,N_2602);
or U3464 (N_3464,N_2708,N_2894);
and U3465 (N_3465,N_2522,N_2708);
or U3466 (N_3466,N_2677,N_2971);
nor U3467 (N_3467,N_2519,N_2730);
or U3468 (N_3468,N_2639,N_2500);
nand U3469 (N_3469,N_2851,N_2795);
nor U3470 (N_3470,N_2968,N_2841);
nand U3471 (N_3471,N_2935,N_2691);
or U3472 (N_3472,N_2555,N_2897);
nor U3473 (N_3473,N_2944,N_2611);
nand U3474 (N_3474,N_2979,N_2900);
nand U3475 (N_3475,N_2672,N_2824);
and U3476 (N_3476,N_2703,N_2683);
nand U3477 (N_3477,N_2730,N_2549);
and U3478 (N_3478,N_2515,N_2637);
nand U3479 (N_3479,N_2912,N_2966);
and U3480 (N_3480,N_2686,N_2890);
nand U3481 (N_3481,N_2656,N_2939);
nor U3482 (N_3482,N_2687,N_2554);
nand U3483 (N_3483,N_2990,N_2909);
nor U3484 (N_3484,N_2831,N_2802);
nor U3485 (N_3485,N_2709,N_2633);
nand U3486 (N_3486,N_2667,N_2795);
or U3487 (N_3487,N_2609,N_2680);
nor U3488 (N_3488,N_2989,N_2756);
nor U3489 (N_3489,N_2604,N_2838);
or U3490 (N_3490,N_2546,N_2620);
nor U3491 (N_3491,N_2507,N_2708);
nor U3492 (N_3492,N_2637,N_2589);
nand U3493 (N_3493,N_2749,N_2839);
nor U3494 (N_3494,N_2815,N_2833);
or U3495 (N_3495,N_2546,N_2713);
and U3496 (N_3496,N_2597,N_2656);
and U3497 (N_3497,N_2654,N_2753);
nor U3498 (N_3498,N_2694,N_2976);
or U3499 (N_3499,N_2644,N_2804);
nand U3500 (N_3500,N_3111,N_3080);
nand U3501 (N_3501,N_3057,N_3029);
nand U3502 (N_3502,N_3369,N_3065);
nand U3503 (N_3503,N_3190,N_3481);
and U3504 (N_3504,N_3416,N_3015);
nor U3505 (N_3505,N_3364,N_3415);
or U3506 (N_3506,N_3084,N_3116);
nand U3507 (N_3507,N_3449,N_3236);
nor U3508 (N_3508,N_3157,N_3192);
and U3509 (N_3509,N_3058,N_3028);
nand U3510 (N_3510,N_3455,N_3120);
nor U3511 (N_3511,N_3314,N_3278);
and U3512 (N_3512,N_3424,N_3471);
or U3513 (N_3513,N_3330,N_3174);
nor U3514 (N_3514,N_3326,N_3468);
and U3515 (N_3515,N_3127,N_3460);
nor U3516 (N_3516,N_3377,N_3279);
nand U3517 (N_3517,N_3323,N_3012);
and U3518 (N_3518,N_3207,N_3059);
and U3519 (N_3519,N_3394,N_3165);
or U3520 (N_3520,N_3143,N_3177);
and U3521 (N_3521,N_3422,N_3311);
nand U3522 (N_3522,N_3421,N_3123);
nor U3523 (N_3523,N_3488,N_3469);
and U3524 (N_3524,N_3193,N_3348);
nand U3525 (N_3525,N_3290,N_3434);
and U3526 (N_3526,N_3341,N_3401);
nand U3527 (N_3527,N_3266,N_3342);
and U3528 (N_3528,N_3117,N_3408);
or U3529 (N_3529,N_3362,N_3244);
nand U3530 (N_3530,N_3461,N_3350);
or U3531 (N_3531,N_3257,N_3289);
nor U3532 (N_3532,N_3126,N_3475);
or U3533 (N_3533,N_3349,N_3403);
nand U3534 (N_3534,N_3105,N_3071);
or U3535 (N_3535,N_3281,N_3067);
nor U3536 (N_3536,N_3285,N_3052);
and U3537 (N_3537,N_3405,N_3465);
nand U3538 (N_3538,N_3466,N_3173);
nor U3539 (N_3539,N_3114,N_3131);
and U3540 (N_3540,N_3083,N_3115);
or U3541 (N_3541,N_3081,N_3498);
or U3542 (N_3542,N_3370,N_3474);
nor U3543 (N_3543,N_3159,N_3354);
xor U3544 (N_3544,N_3176,N_3452);
nor U3545 (N_3545,N_3258,N_3448);
nor U3546 (N_3546,N_3163,N_3287);
nand U3547 (N_3547,N_3494,N_3194);
and U3548 (N_3548,N_3160,N_3245);
and U3549 (N_3549,N_3361,N_3156);
nand U3550 (N_3550,N_3056,N_3274);
and U3551 (N_3551,N_3484,N_3388);
nand U3552 (N_3552,N_3148,N_3486);
nor U3553 (N_3553,N_3049,N_3025);
or U3554 (N_3554,N_3164,N_3172);
or U3555 (N_3555,N_3208,N_3203);
nand U3556 (N_3556,N_3016,N_3187);
nor U3557 (N_3557,N_3396,N_3064);
or U3558 (N_3558,N_3136,N_3209);
and U3559 (N_3559,N_3368,N_3243);
and U3560 (N_3560,N_3231,N_3457);
and U3561 (N_3561,N_3138,N_3464);
nor U3562 (N_3562,N_3296,N_3150);
and U3563 (N_3563,N_3395,N_3476);
nor U3564 (N_3564,N_3041,N_3202);
or U3565 (N_3565,N_3134,N_3376);
or U3566 (N_3566,N_3053,N_3493);
or U3567 (N_3567,N_3227,N_3409);
and U3568 (N_3568,N_3072,N_3298);
and U3569 (N_3569,N_3068,N_3217);
and U3570 (N_3570,N_3318,N_3410);
and U3571 (N_3571,N_3079,N_3024);
xnor U3572 (N_3572,N_3035,N_3199);
and U3573 (N_3573,N_3276,N_3107);
nor U3574 (N_3574,N_3213,N_3099);
nor U3575 (N_3575,N_3215,N_3070);
nor U3576 (N_3576,N_3175,N_3479);
or U3577 (N_3577,N_3280,N_3344);
nor U3578 (N_3578,N_3122,N_3091);
or U3579 (N_3579,N_3275,N_3201);
nor U3580 (N_3580,N_3265,N_3003);
and U3581 (N_3581,N_3008,N_3291);
or U3582 (N_3582,N_3188,N_3295);
or U3583 (N_3583,N_3251,N_3022);
nor U3584 (N_3584,N_3441,N_3262);
nor U3585 (N_3585,N_3020,N_3145);
and U3586 (N_3586,N_3205,N_3332);
or U3587 (N_3587,N_3086,N_3229);
nor U3588 (N_3588,N_3212,N_3018);
nand U3589 (N_3589,N_3151,N_3168);
and U3590 (N_3590,N_3397,N_3007);
or U3591 (N_3591,N_3263,N_3011);
or U3592 (N_3592,N_3261,N_3382);
or U3593 (N_3593,N_3200,N_3306);
xor U3594 (N_3594,N_3030,N_3129);
nor U3595 (N_3595,N_3256,N_3470);
nor U3596 (N_3596,N_3100,N_3288);
nand U3597 (N_3597,N_3338,N_3305);
nor U3598 (N_3598,N_3125,N_3186);
and U3599 (N_3599,N_3496,N_3324);
nor U3600 (N_3600,N_3197,N_3169);
nor U3601 (N_3601,N_3109,N_3429);
or U3602 (N_3602,N_3363,N_3392);
or U3603 (N_3603,N_3247,N_3443);
nor U3604 (N_3604,N_3389,N_3155);
and U3605 (N_3605,N_3228,N_3238);
or U3606 (N_3606,N_3264,N_3218);
nor U3607 (N_3607,N_3268,N_3180);
nor U3608 (N_3608,N_3359,N_3412);
and U3609 (N_3609,N_3055,N_3034);
nor U3610 (N_3610,N_3343,N_3005);
nand U3611 (N_3611,N_3373,N_3427);
xnor U3612 (N_3612,N_3358,N_3004);
nor U3613 (N_3613,N_3050,N_3355);
nor U3614 (N_3614,N_3299,N_3185);
nand U3615 (N_3615,N_3000,N_3402);
or U3616 (N_3616,N_3346,N_3487);
nand U3617 (N_3617,N_3170,N_3032);
or U3618 (N_3618,N_3076,N_3152);
and U3619 (N_3619,N_3226,N_3327);
or U3620 (N_3620,N_3241,N_3432);
nor U3621 (N_3621,N_3304,N_3319);
or U3622 (N_3622,N_3260,N_3027);
nand U3623 (N_3623,N_3183,N_3356);
or U3624 (N_3624,N_3308,N_3423);
xor U3625 (N_3625,N_3378,N_3092);
and U3626 (N_3626,N_3144,N_3098);
and U3627 (N_3627,N_3237,N_3184);
nand U3628 (N_3628,N_3130,N_3335);
nor U3629 (N_3629,N_3339,N_3234);
and U3630 (N_3630,N_3090,N_3069);
or U3631 (N_3631,N_3482,N_3088);
nor U3632 (N_3632,N_3379,N_3300);
and U3633 (N_3633,N_3104,N_3273);
nand U3634 (N_3634,N_3492,N_3073);
nand U3635 (N_3635,N_3235,N_3031);
or U3636 (N_3636,N_3087,N_3446);
nor U3637 (N_3637,N_3042,N_3490);
nor U3638 (N_3638,N_3082,N_3267);
nand U3639 (N_3639,N_3210,N_3095);
or U3640 (N_3640,N_3062,N_3230);
and U3641 (N_3641,N_3096,N_3121);
or U3642 (N_3642,N_3413,N_3106);
nand U3643 (N_3643,N_3347,N_3407);
or U3644 (N_3644,N_3246,N_3371);
nand U3645 (N_3645,N_3112,N_3418);
or U3646 (N_3646,N_3473,N_3282);
and U3647 (N_3647,N_3398,N_3269);
or U3648 (N_3648,N_3045,N_3320);
and U3649 (N_3649,N_3309,N_3271);
and U3650 (N_3650,N_3206,N_3497);
and U3651 (N_3651,N_3181,N_3019);
and U3652 (N_3652,N_3297,N_3154);
nor U3653 (N_3653,N_3047,N_3224);
nand U3654 (N_3654,N_3002,N_3385);
nand U3655 (N_3655,N_3480,N_3312);
or U3656 (N_3656,N_3102,N_3146);
nor U3657 (N_3657,N_3171,N_3060);
or U3658 (N_3658,N_3317,N_3133);
nor U3659 (N_3659,N_3255,N_3303);
nand U3660 (N_3660,N_3435,N_3337);
nand U3661 (N_3661,N_3431,N_3137);
nand U3662 (N_3662,N_3259,N_3331);
or U3663 (N_3663,N_3037,N_3038);
or U3664 (N_3664,N_3239,N_3232);
nand U3665 (N_3665,N_3233,N_3414);
or U3666 (N_3666,N_3372,N_3094);
nor U3667 (N_3667,N_3310,N_3375);
nand U3668 (N_3668,N_3139,N_3078);
nand U3669 (N_3669,N_3046,N_3380);
or U3670 (N_3670,N_3179,N_3292);
nor U3671 (N_3671,N_3214,N_3485);
nor U3672 (N_3672,N_3043,N_3216);
nand U3673 (N_3673,N_3039,N_3110);
and U3674 (N_3674,N_3436,N_3017);
nand U3675 (N_3675,N_3438,N_3454);
or U3676 (N_3676,N_3428,N_3089);
or U3677 (N_3677,N_3253,N_3333);
nand U3678 (N_3678,N_3437,N_3430);
nand U3679 (N_3679,N_3499,N_3467);
and U3680 (N_3680,N_3103,N_3366);
or U3681 (N_3681,N_3097,N_3010);
nor U3682 (N_3682,N_3400,N_3383);
or U3683 (N_3683,N_3447,N_3124);
nor U3684 (N_3684,N_3294,N_3336);
or U3685 (N_3685,N_3367,N_3054);
or U3686 (N_3686,N_3381,N_3153);
or U3687 (N_3687,N_3451,N_3277);
nand U3688 (N_3688,N_3178,N_3093);
nand U3689 (N_3689,N_3036,N_3426);
or U3690 (N_3690,N_3272,N_3472);
and U3691 (N_3691,N_3167,N_3390);
and U3692 (N_3692,N_3462,N_3211);
or U3693 (N_3693,N_3147,N_3014);
nand U3694 (N_3694,N_3351,N_3450);
nor U3695 (N_3695,N_3302,N_3440);
nor U3696 (N_3696,N_3048,N_3458);
nor U3697 (N_3697,N_3417,N_3419);
nand U3698 (N_3698,N_3021,N_3051);
or U3699 (N_3699,N_3463,N_3254);
nand U3700 (N_3700,N_3196,N_3374);
or U3701 (N_3701,N_3353,N_3182);
or U3702 (N_3702,N_3453,N_3240);
and U3703 (N_3703,N_3286,N_3220);
nor U3704 (N_3704,N_3132,N_3495);
or U3705 (N_3705,N_3313,N_3033);
or U3706 (N_3706,N_3135,N_3283);
nand U3707 (N_3707,N_3101,N_3478);
nand U3708 (N_3708,N_3252,N_3433);
nor U3709 (N_3709,N_3158,N_3219);
and U3710 (N_3710,N_3321,N_3322);
nor U3711 (N_3711,N_3006,N_3248);
and U3712 (N_3712,N_3357,N_3442);
nor U3713 (N_3713,N_3189,N_3119);
or U3714 (N_3714,N_3340,N_3483);
or U3715 (N_3715,N_3113,N_3085);
nor U3716 (N_3716,N_3191,N_3140);
nor U3717 (N_3717,N_3001,N_3066);
and U3718 (N_3718,N_3459,N_3149);
nand U3719 (N_3719,N_3365,N_3387);
or U3720 (N_3720,N_3108,N_3393);
nor U3721 (N_3721,N_3128,N_3040);
or U3722 (N_3722,N_3166,N_3360);
and U3723 (N_3723,N_3444,N_3023);
nand U3724 (N_3724,N_3325,N_3063);
and U3725 (N_3725,N_3420,N_3077);
or U3726 (N_3726,N_3439,N_3315);
nor U3727 (N_3727,N_3061,N_3118);
and U3728 (N_3728,N_3026,N_3445);
or U3729 (N_3729,N_3074,N_3477);
or U3730 (N_3730,N_3386,N_3161);
and U3731 (N_3731,N_3307,N_3225);
and U3732 (N_3732,N_3270,N_3142);
nand U3733 (N_3733,N_3250,N_3204);
or U3734 (N_3734,N_3075,N_3328);
or U3735 (N_3735,N_3489,N_3222);
nor U3736 (N_3736,N_3491,N_3221);
and U3737 (N_3737,N_3223,N_3352);
or U3738 (N_3738,N_3198,N_3456);
or U3739 (N_3739,N_3404,N_3391);
nand U3740 (N_3740,N_3425,N_3009);
nand U3741 (N_3741,N_3162,N_3249);
nor U3742 (N_3742,N_3044,N_3345);
nor U3743 (N_3743,N_3399,N_3406);
or U3744 (N_3744,N_3293,N_3334);
and U3745 (N_3745,N_3013,N_3316);
or U3746 (N_3746,N_3384,N_3411);
nor U3747 (N_3747,N_3284,N_3242);
or U3748 (N_3748,N_3329,N_3195);
nand U3749 (N_3749,N_3141,N_3301);
and U3750 (N_3750,N_3217,N_3481);
and U3751 (N_3751,N_3322,N_3017);
or U3752 (N_3752,N_3478,N_3151);
or U3753 (N_3753,N_3056,N_3487);
or U3754 (N_3754,N_3213,N_3474);
and U3755 (N_3755,N_3499,N_3341);
or U3756 (N_3756,N_3448,N_3023);
nand U3757 (N_3757,N_3458,N_3239);
nor U3758 (N_3758,N_3324,N_3455);
and U3759 (N_3759,N_3071,N_3000);
nand U3760 (N_3760,N_3215,N_3306);
and U3761 (N_3761,N_3385,N_3393);
and U3762 (N_3762,N_3341,N_3105);
nor U3763 (N_3763,N_3113,N_3499);
or U3764 (N_3764,N_3497,N_3267);
nor U3765 (N_3765,N_3099,N_3351);
and U3766 (N_3766,N_3081,N_3453);
nor U3767 (N_3767,N_3101,N_3166);
and U3768 (N_3768,N_3109,N_3250);
nor U3769 (N_3769,N_3445,N_3152);
nor U3770 (N_3770,N_3157,N_3373);
or U3771 (N_3771,N_3345,N_3443);
or U3772 (N_3772,N_3106,N_3019);
or U3773 (N_3773,N_3306,N_3153);
or U3774 (N_3774,N_3386,N_3048);
and U3775 (N_3775,N_3368,N_3343);
or U3776 (N_3776,N_3463,N_3321);
and U3777 (N_3777,N_3385,N_3145);
and U3778 (N_3778,N_3443,N_3303);
or U3779 (N_3779,N_3036,N_3444);
and U3780 (N_3780,N_3156,N_3127);
and U3781 (N_3781,N_3067,N_3192);
nand U3782 (N_3782,N_3132,N_3112);
nor U3783 (N_3783,N_3284,N_3250);
and U3784 (N_3784,N_3397,N_3015);
nor U3785 (N_3785,N_3247,N_3495);
nor U3786 (N_3786,N_3310,N_3381);
and U3787 (N_3787,N_3429,N_3203);
and U3788 (N_3788,N_3383,N_3069);
or U3789 (N_3789,N_3088,N_3458);
nor U3790 (N_3790,N_3170,N_3118);
nor U3791 (N_3791,N_3103,N_3063);
or U3792 (N_3792,N_3402,N_3018);
xor U3793 (N_3793,N_3008,N_3051);
or U3794 (N_3794,N_3220,N_3420);
or U3795 (N_3795,N_3460,N_3067);
nand U3796 (N_3796,N_3393,N_3362);
nand U3797 (N_3797,N_3113,N_3453);
and U3798 (N_3798,N_3445,N_3178);
nor U3799 (N_3799,N_3017,N_3359);
nand U3800 (N_3800,N_3111,N_3200);
nand U3801 (N_3801,N_3008,N_3305);
or U3802 (N_3802,N_3151,N_3112);
xor U3803 (N_3803,N_3330,N_3054);
nor U3804 (N_3804,N_3180,N_3326);
nor U3805 (N_3805,N_3214,N_3061);
nor U3806 (N_3806,N_3191,N_3010);
nor U3807 (N_3807,N_3196,N_3234);
and U3808 (N_3808,N_3204,N_3234);
and U3809 (N_3809,N_3225,N_3311);
and U3810 (N_3810,N_3492,N_3312);
or U3811 (N_3811,N_3101,N_3366);
nor U3812 (N_3812,N_3316,N_3279);
nor U3813 (N_3813,N_3194,N_3310);
nor U3814 (N_3814,N_3429,N_3011);
nand U3815 (N_3815,N_3009,N_3290);
nor U3816 (N_3816,N_3109,N_3235);
and U3817 (N_3817,N_3249,N_3126);
nand U3818 (N_3818,N_3464,N_3081);
nor U3819 (N_3819,N_3011,N_3498);
nand U3820 (N_3820,N_3477,N_3288);
or U3821 (N_3821,N_3135,N_3091);
nor U3822 (N_3822,N_3195,N_3386);
or U3823 (N_3823,N_3402,N_3099);
and U3824 (N_3824,N_3219,N_3279);
nor U3825 (N_3825,N_3257,N_3171);
nand U3826 (N_3826,N_3178,N_3077);
or U3827 (N_3827,N_3040,N_3265);
or U3828 (N_3828,N_3214,N_3258);
nand U3829 (N_3829,N_3301,N_3200);
nand U3830 (N_3830,N_3217,N_3456);
nand U3831 (N_3831,N_3179,N_3194);
and U3832 (N_3832,N_3410,N_3038);
or U3833 (N_3833,N_3003,N_3282);
nand U3834 (N_3834,N_3236,N_3022);
nand U3835 (N_3835,N_3246,N_3011);
and U3836 (N_3836,N_3180,N_3014);
or U3837 (N_3837,N_3250,N_3254);
nor U3838 (N_3838,N_3242,N_3286);
nand U3839 (N_3839,N_3129,N_3170);
nand U3840 (N_3840,N_3252,N_3337);
nor U3841 (N_3841,N_3243,N_3164);
or U3842 (N_3842,N_3268,N_3207);
nand U3843 (N_3843,N_3369,N_3296);
or U3844 (N_3844,N_3215,N_3390);
and U3845 (N_3845,N_3235,N_3190);
and U3846 (N_3846,N_3040,N_3042);
or U3847 (N_3847,N_3033,N_3126);
and U3848 (N_3848,N_3270,N_3269);
or U3849 (N_3849,N_3485,N_3445);
nand U3850 (N_3850,N_3423,N_3461);
nor U3851 (N_3851,N_3377,N_3206);
or U3852 (N_3852,N_3083,N_3205);
and U3853 (N_3853,N_3436,N_3380);
nor U3854 (N_3854,N_3387,N_3442);
nor U3855 (N_3855,N_3249,N_3003);
or U3856 (N_3856,N_3367,N_3183);
nand U3857 (N_3857,N_3173,N_3487);
or U3858 (N_3858,N_3107,N_3009);
nand U3859 (N_3859,N_3312,N_3416);
nor U3860 (N_3860,N_3236,N_3475);
and U3861 (N_3861,N_3073,N_3470);
nand U3862 (N_3862,N_3074,N_3392);
and U3863 (N_3863,N_3203,N_3294);
nand U3864 (N_3864,N_3153,N_3207);
nand U3865 (N_3865,N_3045,N_3046);
or U3866 (N_3866,N_3107,N_3486);
nor U3867 (N_3867,N_3371,N_3125);
or U3868 (N_3868,N_3091,N_3333);
or U3869 (N_3869,N_3236,N_3294);
nand U3870 (N_3870,N_3392,N_3367);
and U3871 (N_3871,N_3046,N_3094);
and U3872 (N_3872,N_3251,N_3156);
nand U3873 (N_3873,N_3032,N_3105);
nand U3874 (N_3874,N_3236,N_3014);
nand U3875 (N_3875,N_3414,N_3237);
nor U3876 (N_3876,N_3198,N_3024);
or U3877 (N_3877,N_3486,N_3137);
and U3878 (N_3878,N_3170,N_3214);
or U3879 (N_3879,N_3234,N_3143);
or U3880 (N_3880,N_3281,N_3241);
nand U3881 (N_3881,N_3385,N_3232);
or U3882 (N_3882,N_3153,N_3295);
or U3883 (N_3883,N_3140,N_3097);
and U3884 (N_3884,N_3336,N_3328);
or U3885 (N_3885,N_3283,N_3413);
or U3886 (N_3886,N_3269,N_3276);
nor U3887 (N_3887,N_3137,N_3222);
and U3888 (N_3888,N_3168,N_3323);
or U3889 (N_3889,N_3245,N_3439);
nand U3890 (N_3890,N_3466,N_3487);
nand U3891 (N_3891,N_3221,N_3464);
and U3892 (N_3892,N_3085,N_3351);
nand U3893 (N_3893,N_3249,N_3380);
and U3894 (N_3894,N_3385,N_3024);
and U3895 (N_3895,N_3219,N_3074);
nor U3896 (N_3896,N_3459,N_3223);
nor U3897 (N_3897,N_3298,N_3095);
nand U3898 (N_3898,N_3460,N_3375);
nor U3899 (N_3899,N_3136,N_3248);
and U3900 (N_3900,N_3120,N_3458);
nor U3901 (N_3901,N_3010,N_3157);
nor U3902 (N_3902,N_3456,N_3073);
nor U3903 (N_3903,N_3159,N_3328);
nand U3904 (N_3904,N_3467,N_3478);
and U3905 (N_3905,N_3113,N_3025);
and U3906 (N_3906,N_3093,N_3079);
nor U3907 (N_3907,N_3320,N_3165);
nand U3908 (N_3908,N_3364,N_3222);
xnor U3909 (N_3909,N_3192,N_3439);
and U3910 (N_3910,N_3163,N_3464);
nand U3911 (N_3911,N_3042,N_3465);
nand U3912 (N_3912,N_3118,N_3146);
nand U3913 (N_3913,N_3069,N_3118);
nand U3914 (N_3914,N_3313,N_3449);
nand U3915 (N_3915,N_3243,N_3250);
nand U3916 (N_3916,N_3459,N_3047);
nand U3917 (N_3917,N_3384,N_3324);
and U3918 (N_3918,N_3085,N_3384);
nand U3919 (N_3919,N_3010,N_3456);
and U3920 (N_3920,N_3291,N_3419);
or U3921 (N_3921,N_3164,N_3137);
and U3922 (N_3922,N_3282,N_3213);
nand U3923 (N_3923,N_3444,N_3239);
nand U3924 (N_3924,N_3423,N_3220);
and U3925 (N_3925,N_3231,N_3019);
and U3926 (N_3926,N_3151,N_3079);
nand U3927 (N_3927,N_3201,N_3121);
and U3928 (N_3928,N_3225,N_3468);
nand U3929 (N_3929,N_3339,N_3423);
nor U3930 (N_3930,N_3487,N_3428);
or U3931 (N_3931,N_3247,N_3483);
nor U3932 (N_3932,N_3311,N_3392);
nor U3933 (N_3933,N_3222,N_3023);
nor U3934 (N_3934,N_3321,N_3013);
nand U3935 (N_3935,N_3164,N_3279);
nor U3936 (N_3936,N_3204,N_3458);
or U3937 (N_3937,N_3135,N_3294);
and U3938 (N_3938,N_3217,N_3214);
or U3939 (N_3939,N_3492,N_3448);
or U3940 (N_3940,N_3024,N_3210);
or U3941 (N_3941,N_3050,N_3322);
nand U3942 (N_3942,N_3398,N_3473);
nor U3943 (N_3943,N_3258,N_3185);
nor U3944 (N_3944,N_3058,N_3439);
or U3945 (N_3945,N_3284,N_3177);
nor U3946 (N_3946,N_3094,N_3104);
nor U3947 (N_3947,N_3364,N_3113);
or U3948 (N_3948,N_3105,N_3251);
nand U3949 (N_3949,N_3030,N_3252);
nor U3950 (N_3950,N_3416,N_3474);
nand U3951 (N_3951,N_3042,N_3289);
nor U3952 (N_3952,N_3457,N_3293);
nand U3953 (N_3953,N_3119,N_3372);
nor U3954 (N_3954,N_3089,N_3185);
nand U3955 (N_3955,N_3470,N_3255);
nor U3956 (N_3956,N_3362,N_3256);
and U3957 (N_3957,N_3454,N_3183);
nor U3958 (N_3958,N_3103,N_3420);
and U3959 (N_3959,N_3294,N_3470);
or U3960 (N_3960,N_3333,N_3464);
nand U3961 (N_3961,N_3466,N_3442);
nor U3962 (N_3962,N_3288,N_3291);
nor U3963 (N_3963,N_3145,N_3168);
nand U3964 (N_3964,N_3351,N_3280);
nor U3965 (N_3965,N_3105,N_3131);
nor U3966 (N_3966,N_3135,N_3498);
or U3967 (N_3967,N_3336,N_3400);
nand U3968 (N_3968,N_3252,N_3056);
or U3969 (N_3969,N_3214,N_3213);
nor U3970 (N_3970,N_3372,N_3425);
and U3971 (N_3971,N_3041,N_3367);
nand U3972 (N_3972,N_3340,N_3141);
nor U3973 (N_3973,N_3215,N_3327);
and U3974 (N_3974,N_3397,N_3443);
nand U3975 (N_3975,N_3358,N_3072);
or U3976 (N_3976,N_3242,N_3237);
nor U3977 (N_3977,N_3187,N_3485);
nor U3978 (N_3978,N_3150,N_3037);
nand U3979 (N_3979,N_3144,N_3091);
nand U3980 (N_3980,N_3433,N_3253);
or U3981 (N_3981,N_3170,N_3388);
or U3982 (N_3982,N_3048,N_3407);
nor U3983 (N_3983,N_3142,N_3283);
xnor U3984 (N_3984,N_3150,N_3062);
and U3985 (N_3985,N_3204,N_3185);
nor U3986 (N_3986,N_3373,N_3481);
nor U3987 (N_3987,N_3185,N_3202);
nor U3988 (N_3988,N_3429,N_3295);
nand U3989 (N_3989,N_3049,N_3390);
or U3990 (N_3990,N_3365,N_3146);
and U3991 (N_3991,N_3172,N_3471);
and U3992 (N_3992,N_3253,N_3398);
or U3993 (N_3993,N_3131,N_3319);
or U3994 (N_3994,N_3233,N_3325);
and U3995 (N_3995,N_3472,N_3378);
nor U3996 (N_3996,N_3322,N_3438);
and U3997 (N_3997,N_3480,N_3064);
or U3998 (N_3998,N_3230,N_3412);
nand U3999 (N_3999,N_3322,N_3152);
nand U4000 (N_4000,N_3651,N_3596);
or U4001 (N_4001,N_3695,N_3703);
nor U4002 (N_4002,N_3717,N_3776);
nand U4003 (N_4003,N_3927,N_3733);
or U4004 (N_4004,N_3983,N_3999);
and U4005 (N_4005,N_3917,N_3716);
or U4006 (N_4006,N_3548,N_3872);
or U4007 (N_4007,N_3754,N_3971);
or U4008 (N_4008,N_3541,N_3636);
and U4009 (N_4009,N_3663,N_3792);
and U4010 (N_4010,N_3712,N_3959);
or U4011 (N_4011,N_3827,N_3830);
and U4012 (N_4012,N_3678,N_3730);
nor U4013 (N_4013,N_3839,N_3883);
nor U4014 (N_4014,N_3648,N_3696);
or U4015 (N_4015,N_3553,N_3610);
or U4016 (N_4016,N_3879,N_3860);
and U4017 (N_4017,N_3990,N_3563);
nand U4018 (N_4018,N_3653,N_3924);
nand U4019 (N_4019,N_3940,N_3794);
and U4020 (N_4020,N_3930,N_3787);
or U4021 (N_4021,N_3685,N_3580);
nand U4022 (N_4022,N_3968,N_3600);
and U4023 (N_4023,N_3539,N_3744);
and U4024 (N_4024,N_3858,N_3944);
nand U4025 (N_4025,N_3649,N_3767);
nor U4026 (N_4026,N_3699,N_3774);
nand U4027 (N_4027,N_3997,N_3892);
nand U4028 (N_4028,N_3618,N_3813);
nand U4029 (N_4029,N_3627,N_3739);
and U4030 (N_4030,N_3764,N_3902);
nand U4031 (N_4031,N_3661,N_3547);
or U4032 (N_4032,N_3701,N_3668);
or U4033 (N_4033,N_3903,N_3840);
nor U4034 (N_4034,N_3756,N_3738);
or U4035 (N_4035,N_3743,N_3537);
or U4036 (N_4036,N_3808,N_3722);
nand U4037 (N_4037,N_3884,N_3876);
nor U4038 (N_4038,N_3597,N_3629);
or U4039 (N_4039,N_3612,N_3848);
nand U4040 (N_4040,N_3786,N_3688);
and U4041 (N_4041,N_3846,N_3804);
nand U4042 (N_4042,N_3535,N_3590);
nor U4043 (N_4043,N_3602,N_3953);
nor U4044 (N_4044,N_3992,N_3849);
nor U4045 (N_4045,N_3569,N_3766);
or U4046 (N_4046,N_3855,N_3615);
nand U4047 (N_4047,N_3975,N_3518);
or U4048 (N_4048,N_3877,N_3562);
and U4049 (N_4049,N_3785,N_3505);
nor U4050 (N_4050,N_3740,N_3735);
nor U4051 (N_4051,N_3891,N_3994);
or U4052 (N_4052,N_3727,N_3991);
nor U4053 (N_4053,N_3543,N_3556);
and U4054 (N_4054,N_3585,N_3622);
and U4055 (N_4055,N_3878,N_3851);
nor U4056 (N_4056,N_3502,N_3910);
xnor U4057 (N_4057,N_3709,N_3942);
nor U4058 (N_4058,N_3519,N_3885);
nor U4059 (N_4059,N_3868,N_3698);
nor U4060 (N_4060,N_3731,N_3573);
or U4061 (N_4061,N_3993,N_3824);
nand U4062 (N_4062,N_3647,N_3711);
nor U4063 (N_4063,N_3886,N_3669);
or U4064 (N_4064,N_3601,N_3915);
or U4065 (N_4065,N_3842,N_3591);
nor U4066 (N_4066,N_3859,N_3675);
nor U4067 (N_4067,N_3838,N_3864);
nand U4068 (N_4068,N_3586,N_3869);
xnor U4069 (N_4069,N_3987,N_3758);
nor U4070 (N_4070,N_3530,N_3689);
or U4071 (N_4071,N_3576,N_3962);
nand U4072 (N_4072,N_3707,N_3955);
nand U4073 (N_4073,N_3723,N_3963);
or U4074 (N_4074,N_3683,N_3835);
nand U4075 (N_4075,N_3866,N_3826);
nand U4076 (N_4076,N_3624,N_3800);
nand U4077 (N_4077,N_3687,N_3515);
or U4078 (N_4078,N_3524,N_3783);
nand U4079 (N_4079,N_3697,N_3901);
or U4080 (N_4080,N_3575,N_3939);
or U4081 (N_4081,N_3947,N_3603);
and U4082 (N_4082,N_3666,N_3873);
nor U4083 (N_4083,N_3728,N_3906);
and U4084 (N_4084,N_3510,N_3814);
nor U4085 (N_4085,N_3920,N_3880);
nor U4086 (N_4086,N_3751,N_3631);
or U4087 (N_4087,N_3934,N_3657);
and U4088 (N_4088,N_3941,N_3501);
and U4089 (N_4089,N_3907,N_3960);
nand U4090 (N_4090,N_3887,N_3888);
nor U4091 (N_4091,N_3644,N_3823);
nand U4092 (N_4092,N_3998,N_3718);
nand U4093 (N_4093,N_3755,N_3599);
or U4094 (N_4094,N_3558,N_3912);
and U4095 (N_4095,N_3807,N_3988);
nand U4096 (N_4096,N_3506,N_3784);
and U4097 (N_4097,N_3995,N_3904);
or U4098 (N_4098,N_3528,N_3554);
or U4099 (N_4099,N_3650,N_3522);
and U4100 (N_4100,N_3828,N_3978);
or U4101 (N_4101,N_3677,N_3704);
and U4102 (N_4102,N_3874,N_3825);
nor U4103 (N_4103,N_3625,N_3605);
nor U4104 (N_4104,N_3802,N_3936);
nor U4105 (N_4105,N_3692,N_3925);
nor U4106 (N_4106,N_3616,N_3761);
nand U4107 (N_4107,N_3911,N_3578);
and U4108 (N_4108,N_3882,N_3565);
nor U4109 (N_4109,N_3725,N_3742);
nor U4110 (N_4110,N_3979,N_3621);
or U4111 (N_4111,N_3900,N_3918);
nand U4112 (N_4112,N_3806,N_3822);
nand U4113 (N_4113,N_3641,N_3973);
nand U4114 (N_4114,N_3574,N_3513);
nand U4115 (N_4115,N_3659,N_3750);
nor U4116 (N_4116,N_3948,N_3760);
nand U4117 (N_4117,N_3665,N_3732);
nand U4118 (N_4118,N_3549,N_3771);
and U4119 (N_4119,N_3536,N_3977);
and U4120 (N_4120,N_3950,N_3749);
nor U4121 (N_4121,N_3844,N_3604);
and U4122 (N_4122,N_3980,N_3729);
and U4123 (N_4123,N_3817,N_3845);
and U4124 (N_4124,N_3655,N_3798);
nor U4125 (N_4125,N_3726,N_3639);
or U4126 (N_4126,N_3710,N_3832);
and U4127 (N_4127,N_3521,N_3926);
nor U4128 (N_4128,N_3966,N_3595);
or U4129 (N_4129,N_3670,N_3778);
or U4130 (N_4130,N_3759,N_3769);
or U4131 (N_4131,N_3818,N_3929);
and U4132 (N_4132,N_3662,N_3782);
nor U4133 (N_4133,N_3747,N_3945);
or U4134 (N_4134,N_3763,N_3633);
and U4135 (N_4135,N_3577,N_3555);
nor U4136 (N_4136,N_3635,N_3815);
nand U4137 (N_4137,N_3589,N_3789);
or U4138 (N_4138,N_3608,N_3854);
and U4139 (N_4139,N_3870,N_3606);
nor U4140 (N_4140,N_3875,N_3700);
nand U4141 (N_4141,N_3949,N_3871);
nor U4142 (N_4142,N_3748,N_3682);
nand U4143 (N_4143,N_3752,N_3588);
or U4144 (N_4144,N_3504,N_3834);
or U4145 (N_4145,N_3568,N_3544);
nor U4146 (N_4146,N_3542,N_3526);
and U4147 (N_4147,N_3922,N_3500);
nand U4148 (N_4148,N_3642,N_3693);
nand U4149 (N_4149,N_3974,N_3809);
nor U4150 (N_4150,N_3933,N_3520);
nand U4151 (N_4151,N_3793,N_3724);
and U4152 (N_4152,N_3637,N_3981);
nand U4153 (N_4153,N_3609,N_3923);
and U4154 (N_4154,N_3853,N_3741);
nor U4155 (N_4155,N_3705,N_3713);
nor U4156 (N_4156,N_3671,N_3570);
and U4157 (N_4157,N_3796,N_3531);
nand U4158 (N_4158,N_3736,N_3961);
and U4159 (N_4159,N_3567,N_3914);
nor U4160 (N_4160,N_3937,N_3928);
or U4161 (N_4161,N_3956,N_3538);
and U4162 (N_4162,N_3607,N_3852);
and U4163 (N_4163,N_3836,N_3989);
and U4164 (N_4164,N_3765,N_3921);
and U4165 (N_4165,N_3679,N_3564);
and U4166 (N_4166,N_3831,N_3856);
and U4167 (N_4167,N_3821,N_3656);
nor U4168 (N_4168,N_3511,N_3951);
and U4169 (N_4169,N_3617,N_3909);
and U4170 (N_4170,N_3811,N_3803);
nand U4171 (N_4171,N_3660,N_3819);
and U4172 (N_4172,N_3857,N_3720);
or U4173 (N_4173,N_3533,N_3954);
nor U4174 (N_4174,N_3626,N_3691);
nand U4175 (N_4175,N_3850,N_3516);
nand U4176 (N_4176,N_3634,N_3593);
nand U4177 (N_4177,N_3652,N_3583);
or U4178 (N_4178,N_3581,N_3630);
and U4179 (N_4179,N_3780,N_3805);
nand U4180 (N_4180,N_3781,N_3690);
nand U4181 (N_4181,N_3619,N_3594);
and U4182 (N_4182,N_3721,N_3841);
nor U4183 (N_4183,N_3847,N_3829);
and U4184 (N_4184,N_3791,N_3540);
nor U4185 (N_4185,N_3645,N_3664);
or U4186 (N_4186,N_3584,N_3579);
and U4187 (N_4187,N_3512,N_3938);
nand U4188 (N_4188,N_3587,N_3613);
nand U4189 (N_4189,N_3965,N_3790);
or U4190 (N_4190,N_3810,N_3517);
and U4191 (N_4191,N_3894,N_3714);
and U4192 (N_4192,N_3889,N_3514);
nand U4193 (N_4193,N_3946,N_3816);
nor U4194 (N_4194,N_3734,N_3757);
nor U4195 (N_4195,N_3620,N_3772);
and U4196 (N_4196,N_3932,N_3976);
and U4197 (N_4197,N_3908,N_3837);
or U4198 (N_4198,N_3913,N_3545);
nand U4199 (N_4199,N_3632,N_3865);
nor U4200 (N_4200,N_3561,N_3982);
nand U4201 (N_4201,N_3559,N_3638);
nor U4202 (N_4202,N_3905,N_3779);
nand U4203 (N_4203,N_3560,N_3935);
nor U4204 (N_4204,N_3996,N_3753);
nor U4205 (N_4205,N_3667,N_3985);
nor U4206 (N_4206,N_3557,N_3571);
xor U4207 (N_4207,N_3676,N_3551);
nor U4208 (N_4208,N_3762,N_3795);
nor U4209 (N_4209,N_3534,N_3529);
and U4210 (N_4210,N_3532,N_3943);
and U4211 (N_4211,N_3646,N_3843);
nor U4212 (N_4212,N_3694,N_3546);
nor U4213 (N_4213,N_3788,N_3552);
nand U4214 (N_4214,N_3673,N_3967);
nor U4215 (N_4215,N_3768,N_3820);
nor U4216 (N_4216,N_3986,N_3969);
nor U4217 (N_4217,N_3952,N_3895);
nand U4218 (N_4218,N_3863,N_3715);
and U4219 (N_4219,N_3702,N_3890);
nor U4220 (N_4220,N_3643,N_3706);
and U4221 (N_4221,N_3861,N_3623);
nor U4222 (N_4222,N_3686,N_3507);
or U4223 (N_4223,N_3777,N_3746);
nand U4224 (N_4224,N_3773,N_3674);
nor U4225 (N_4225,N_3899,N_3957);
nor U4226 (N_4226,N_3916,N_3897);
or U4227 (N_4227,N_3509,N_3801);
or U4228 (N_4228,N_3582,N_3898);
nand U4229 (N_4229,N_3508,N_3958);
or U4230 (N_4230,N_3684,N_3611);
nor U4231 (N_4231,N_3592,N_3681);
and U4232 (N_4232,N_3770,N_3598);
and U4233 (N_4233,N_3640,N_3614);
nand U4234 (N_4234,N_3672,N_3919);
nor U4235 (N_4235,N_3775,N_3984);
nand U4236 (N_4236,N_3867,N_3896);
or U4237 (N_4237,N_3572,N_3931);
nand U4238 (N_4238,N_3833,N_3881);
nand U4239 (N_4239,N_3550,N_3719);
or U4240 (N_4240,N_3523,N_3797);
or U4241 (N_4241,N_3525,N_3658);
nor U4242 (N_4242,N_3812,N_3964);
nor U4243 (N_4243,N_3799,N_3566);
nand U4244 (N_4244,N_3972,N_3737);
and U4245 (N_4245,N_3893,N_3708);
nand U4246 (N_4246,N_3503,N_3970);
or U4247 (N_4247,N_3628,N_3745);
nor U4248 (N_4248,N_3654,N_3527);
nor U4249 (N_4249,N_3862,N_3680);
nand U4250 (N_4250,N_3805,N_3510);
or U4251 (N_4251,N_3695,N_3594);
or U4252 (N_4252,N_3971,N_3915);
and U4253 (N_4253,N_3879,N_3842);
nand U4254 (N_4254,N_3690,N_3772);
nor U4255 (N_4255,N_3764,N_3981);
nand U4256 (N_4256,N_3909,N_3889);
or U4257 (N_4257,N_3809,N_3959);
nand U4258 (N_4258,N_3978,N_3994);
nand U4259 (N_4259,N_3962,N_3504);
nand U4260 (N_4260,N_3730,N_3934);
nand U4261 (N_4261,N_3978,N_3912);
and U4262 (N_4262,N_3735,N_3506);
and U4263 (N_4263,N_3792,N_3769);
and U4264 (N_4264,N_3617,N_3580);
nand U4265 (N_4265,N_3545,N_3638);
nand U4266 (N_4266,N_3910,N_3634);
nand U4267 (N_4267,N_3897,N_3689);
nand U4268 (N_4268,N_3849,N_3772);
nor U4269 (N_4269,N_3604,N_3652);
and U4270 (N_4270,N_3628,N_3772);
nand U4271 (N_4271,N_3756,N_3840);
and U4272 (N_4272,N_3774,N_3687);
or U4273 (N_4273,N_3967,N_3629);
nand U4274 (N_4274,N_3742,N_3933);
or U4275 (N_4275,N_3806,N_3504);
nand U4276 (N_4276,N_3526,N_3517);
or U4277 (N_4277,N_3927,N_3794);
and U4278 (N_4278,N_3605,N_3951);
and U4279 (N_4279,N_3692,N_3869);
and U4280 (N_4280,N_3735,N_3983);
or U4281 (N_4281,N_3951,N_3829);
nor U4282 (N_4282,N_3517,N_3757);
nor U4283 (N_4283,N_3805,N_3788);
or U4284 (N_4284,N_3862,N_3584);
nor U4285 (N_4285,N_3947,N_3572);
nand U4286 (N_4286,N_3977,N_3773);
or U4287 (N_4287,N_3560,N_3724);
nand U4288 (N_4288,N_3725,N_3762);
nand U4289 (N_4289,N_3696,N_3559);
or U4290 (N_4290,N_3875,N_3708);
nor U4291 (N_4291,N_3623,N_3848);
nand U4292 (N_4292,N_3748,N_3963);
nor U4293 (N_4293,N_3607,N_3610);
nor U4294 (N_4294,N_3751,N_3808);
nand U4295 (N_4295,N_3589,N_3882);
and U4296 (N_4296,N_3914,N_3555);
nor U4297 (N_4297,N_3576,N_3656);
or U4298 (N_4298,N_3659,N_3896);
nor U4299 (N_4299,N_3851,N_3778);
or U4300 (N_4300,N_3819,N_3992);
and U4301 (N_4301,N_3807,N_3775);
nor U4302 (N_4302,N_3879,N_3599);
and U4303 (N_4303,N_3640,N_3980);
nand U4304 (N_4304,N_3888,N_3738);
nand U4305 (N_4305,N_3604,N_3684);
nor U4306 (N_4306,N_3743,N_3721);
and U4307 (N_4307,N_3574,N_3807);
or U4308 (N_4308,N_3763,N_3765);
nor U4309 (N_4309,N_3582,N_3800);
nand U4310 (N_4310,N_3821,N_3950);
and U4311 (N_4311,N_3825,N_3847);
nor U4312 (N_4312,N_3783,N_3688);
and U4313 (N_4313,N_3711,N_3736);
nand U4314 (N_4314,N_3720,N_3787);
nor U4315 (N_4315,N_3814,N_3516);
nand U4316 (N_4316,N_3662,N_3988);
and U4317 (N_4317,N_3664,N_3831);
nor U4318 (N_4318,N_3635,N_3518);
or U4319 (N_4319,N_3835,N_3765);
and U4320 (N_4320,N_3525,N_3596);
and U4321 (N_4321,N_3830,N_3626);
nand U4322 (N_4322,N_3620,N_3740);
nand U4323 (N_4323,N_3693,N_3627);
and U4324 (N_4324,N_3908,N_3633);
nand U4325 (N_4325,N_3756,N_3533);
nand U4326 (N_4326,N_3803,N_3540);
nor U4327 (N_4327,N_3541,N_3832);
nand U4328 (N_4328,N_3551,N_3882);
or U4329 (N_4329,N_3997,N_3625);
nor U4330 (N_4330,N_3776,N_3794);
and U4331 (N_4331,N_3598,N_3654);
or U4332 (N_4332,N_3803,N_3737);
nand U4333 (N_4333,N_3977,N_3645);
nand U4334 (N_4334,N_3805,N_3856);
or U4335 (N_4335,N_3511,N_3885);
and U4336 (N_4336,N_3881,N_3974);
or U4337 (N_4337,N_3997,N_3999);
or U4338 (N_4338,N_3703,N_3737);
nor U4339 (N_4339,N_3794,N_3813);
and U4340 (N_4340,N_3566,N_3990);
nor U4341 (N_4341,N_3583,N_3642);
nor U4342 (N_4342,N_3771,N_3583);
and U4343 (N_4343,N_3596,N_3605);
and U4344 (N_4344,N_3554,N_3985);
or U4345 (N_4345,N_3785,N_3938);
nor U4346 (N_4346,N_3864,N_3593);
nand U4347 (N_4347,N_3673,N_3944);
nand U4348 (N_4348,N_3837,N_3819);
and U4349 (N_4349,N_3518,N_3621);
or U4350 (N_4350,N_3996,N_3677);
nor U4351 (N_4351,N_3633,N_3693);
nor U4352 (N_4352,N_3587,N_3692);
nor U4353 (N_4353,N_3769,N_3849);
nand U4354 (N_4354,N_3872,N_3883);
and U4355 (N_4355,N_3990,N_3623);
and U4356 (N_4356,N_3954,N_3627);
or U4357 (N_4357,N_3532,N_3593);
or U4358 (N_4358,N_3756,N_3927);
and U4359 (N_4359,N_3629,N_3722);
nand U4360 (N_4360,N_3831,N_3628);
nor U4361 (N_4361,N_3746,N_3838);
and U4362 (N_4362,N_3909,N_3706);
and U4363 (N_4363,N_3992,N_3954);
nand U4364 (N_4364,N_3933,N_3582);
nor U4365 (N_4365,N_3961,N_3698);
or U4366 (N_4366,N_3782,N_3958);
nand U4367 (N_4367,N_3879,N_3563);
and U4368 (N_4368,N_3558,N_3569);
nor U4369 (N_4369,N_3783,N_3634);
or U4370 (N_4370,N_3914,N_3505);
nand U4371 (N_4371,N_3664,N_3810);
and U4372 (N_4372,N_3673,N_3603);
nor U4373 (N_4373,N_3851,N_3576);
or U4374 (N_4374,N_3901,N_3748);
and U4375 (N_4375,N_3764,N_3821);
nand U4376 (N_4376,N_3525,N_3960);
nand U4377 (N_4377,N_3829,N_3810);
and U4378 (N_4378,N_3998,N_3852);
nand U4379 (N_4379,N_3635,N_3654);
nand U4380 (N_4380,N_3523,N_3942);
nor U4381 (N_4381,N_3648,N_3525);
and U4382 (N_4382,N_3597,N_3895);
nor U4383 (N_4383,N_3859,N_3866);
or U4384 (N_4384,N_3867,N_3750);
nor U4385 (N_4385,N_3904,N_3600);
or U4386 (N_4386,N_3667,N_3781);
or U4387 (N_4387,N_3872,N_3964);
nor U4388 (N_4388,N_3598,N_3720);
xnor U4389 (N_4389,N_3634,N_3960);
and U4390 (N_4390,N_3730,N_3875);
or U4391 (N_4391,N_3715,N_3922);
nand U4392 (N_4392,N_3987,N_3845);
and U4393 (N_4393,N_3680,N_3779);
nor U4394 (N_4394,N_3851,N_3560);
nor U4395 (N_4395,N_3870,N_3635);
and U4396 (N_4396,N_3764,N_3693);
nor U4397 (N_4397,N_3856,N_3578);
or U4398 (N_4398,N_3504,N_3707);
or U4399 (N_4399,N_3953,N_3710);
nor U4400 (N_4400,N_3598,N_3914);
and U4401 (N_4401,N_3886,N_3790);
nand U4402 (N_4402,N_3837,N_3682);
or U4403 (N_4403,N_3551,N_3973);
and U4404 (N_4404,N_3962,N_3877);
nor U4405 (N_4405,N_3986,N_3599);
nand U4406 (N_4406,N_3709,N_3784);
nand U4407 (N_4407,N_3611,N_3504);
and U4408 (N_4408,N_3912,N_3819);
and U4409 (N_4409,N_3636,N_3709);
or U4410 (N_4410,N_3500,N_3635);
nand U4411 (N_4411,N_3696,N_3524);
nor U4412 (N_4412,N_3580,N_3790);
nor U4413 (N_4413,N_3537,N_3950);
nor U4414 (N_4414,N_3820,N_3992);
or U4415 (N_4415,N_3579,N_3993);
or U4416 (N_4416,N_3504,N_3719);
nand U4417 (N_4417,N_3893,N_3770);
nand U4418 (N_4418,N_3549,N_3982);
nand U4419 (N_4419,N_3947,N_3783);
nand U4420 (N_4420,N_3614,N_3922);
nor U4421 (N_4421,N_3902,N_3826);
nand U4422 (N_4422,N_3864,N_3780);
nand U4423 (N_4423,N_3805,N_3588);
or U4424 (N_4424,N_3929,N_3988);
nor U4425 (N_4425,N_3737,N_3528);
or U4426 (N_4426,N_3514,N_3914);
nor U4427 (N_4427,N_3861,N_3945);
and U4428 (N_4428,N_3842,N_3969);
and U4429 (N_4429,N_3635,N_3910);
nor U4430 (N_4430,N_3762,N_3842);
nand U4431 (N_4431,N_3949,N_3940);
or U4432 (N_4432,N_3870,N_3977);
nand U4433 (N_4433,N_3822,N_3533);
or U4434 (N_4434,N_3587,N_3677);
and U4435 (N_4435,N_3962,N_3974);
nand U4436 (N_4436,N_3765,N_3750);
or U4437 (N_4437,N_3501,N_3971);
nand U4438 (N_4438,N_3949,N_3648);
xnor U4439 (N_4439,N_3517,N_3814);
or U4440 (N_4440,N_3538,N_3781);
and U4441 (N_4441,N_3828,N_3935);
and U4442 (N_4442,N_3559,N_3839);
or U4443 (N_4443,N_3840,N_3989);
or U4444 (N_4444,N_3532,N_3622);
nand U4445 (N_4445,N_3719,N_3913);
nand U4446 (N_4446,N_3818,N_3625);
nor U4447 (N_4447,N_3789,N_3577);
and U4448 (N_4448,N_3983,N_3678);
nor U4449 (N_4449,N_3507,N_3529);
and U4450 (N_4450,N_3804,N_3653);
or U4451 (N_4451,N_3844,N_3912);
and U4452 (N_4452,N_3922,N_3501);
nor U4453 (N_4453,N_3991,N_3916);
nor U4454 (N_4454,N_3546,N_3586);
and U4455 (N_4455,N_3839,N_3825);
nor U4456 (N_4456,N_3870,N_3550);
nor U4457 (N_4457,N_3593,N_3765);
nand U4458 (N_4458,N_3696,N_3542);
nand U4459 (N_4459,N_3749,N_3595);
nand U4460 (N_4460,N_3718,N_3999);
and U4461 (N_4461,N_3867,N_3928);
nand U4462 (N_4462,N_3844,N_3704);
nor U4463 (N_4463,N_3757,N_3893);
nor U4464 (N_4464,N_3557,N_3993);
nor U4465 (N_4465,N_3679,N_3620);
and U4466 (N_4466,N_3884,N_3571);
nor U4467 (N_4467,N_3891,N_3787);
and U4468 (N_4468,N_3780,N_3527);
nand U4469 (N_4469,N_3722,N_3533);
nand U4470 (N_4470,N_3863,N_3664);
nor U4471 (N_4471,N_3821,N_3943);
or U4472 (N_4472,N_3894,N_3872);
nand U4473 (N_4473,N_3965,N_3578);
nor U4474 (N_4474,N_3816,N_3705);
nand U4475 (N_4475,N_3554,N_3679);
nand U4476 (N_4476,N_3752,N_3811);
nor U4477 (N_4477,N_3514,N_3749);
nor U4478 (N_4478,N_3538,N_3606);
or U4479 (N_4479,N_3679,N_3640);
and U4480 (N_4480,N_3516,N_3717);
or U4481 (N_4481,N_3866,N_3621);
and U4482 (N_4482,N_3579,N_3879);
and U4483 (N_4483,N_3661,N_3767);
or U4484 (N_4484,N_3573,N_3806);
nand U4485 (N_4485,N_3983,N_3884);
nor U4486 (N_4486,N_3795,N_3965);
and U4487 (N_4487,N_3909,N_3581);
nand U4488 (N_4488,N_3695,N_3673);
and U4489 (N_4489,N_3775,N_3824);
and U4490 (N_4490,N_3738,N_3658);
nor U4491 (N_4491,N_3632,N_3695);
nand U4492 (N_4492,N_3701,N_3878);
nor U4493 (N_4493,N_3815,N_3887);
nand U4494 (N_4494,N_3575,N_3891);
nand U4495 (N_4495,N_3945,N_3614);
or U4496 (N_4496,N_3537,N_3750);
nand U4497 (N_4497,N_3512,N_3951);
nor U4498 (N_4498,N_3504,N_3624);
xor U4499 (N_4499,N_3666,N_3733);
xnor U4500 (N_4500,N_4016,N_4482);
and U4501 (N_4501,N_4076,N_4278);
nor U4502 (N_4502,N_4126,N_4494);
nand U4503 (N_4503,N_4224,N_4092);
nor U4504 (N_4504,N_4053,N_4008);
or U4505 (N_4505,N_4246,N_4364);
nand U4506 (N_4506,N_4153,N_4163);
or U4507 (N_4507,N_4478,N_4433);
nand U4508 (N_4508,N_4182,N_4345);
nand U4509 (N_4509,N_4237,N_4460);
and U4510 (N_4510,N_4006,N_4422);
nor U4511 (N_4511,N_4041,N_4238);
and U4512 (N_4512,N_4037,N_4347);
nor U4513 (N_4513,N_4324,N_4388);
nor U4514 (N_4514,N_4413,N_4356);
or U4515 (N_4515,N_4243,N_4461);
and U4516 (N_4516,N_4469,N_4265);
nand U4517 (N_4517,N_4430,N_4212);
and U4518 (N_4518,N_4112,N_4214);
nand U4519 (N_4519,N_4473,N_4048);
nand U4520 (N_4520,N_4401,N_4419);
xor U4521 (N_4521,N_4305,N_4299);
or U4522 (N_4522,N_4239,N_4011);
nand U4523 (N_4523,N_4458,N_4467);
or U4524 (N_4524,N_4102,N_4157);
or U4525 (N_4525,N_4408,N_4040);
nor U4526 (N_4526,N_4149,N_4176);
or U4527 (N_4527,N_4217,N_4403);
and U4528 (N_4528,N_4242,N_4317);
nor U4529 (N_4529,N_4141,N_4368);
or U4530 (N_4530,N_4121,N_4023);
nor U4531 (N_4531,N_4335,N_4385);
and U4532 (N_4532,N_4247,N_4327);
or U4533 (N_4533,N_4480,N_4470);
nor U4534 (N_4534,N_4028,N_4400);
and U4535 (N_4535,N_4117,N_4152);
nor U4536 (N_4536,N_4415,N_4491);
nand U4537 (N_4537,N_4154,N_4412);
nor U4538 (N_4538,N_4380,N_4236);
or U4539 (N_4539,N_4026,N_4424);
or U4540 (N_4540,N_4125,N_4098);
or U4541 (N_4541,N_4488,N_4373);
nor U4542 (N_4542,N_4358,N_4104);
nor U4543 (N_4543,N_4180,N_4199);
nor U4544 (N_4544,N_4302,N_4455);
nand U4545 (N_4545,N_4352,N_4484);
and U4546 (N_4546,N_4392,N_4096);
or U4547 (N_4547,N_4007,N_4267);
nor U4548 (N_4548,N_4277,N_4232);
and U4549 (N_4549,N_4304,N_4283);
or U4550 (N_4550,N_4273,N_4312);
nor U4551 (N_4551,N_4429,N_4326);
or U4552 (N_4552,N_4481,N_4492);
nor U4553 (N_4553,N_4393,N_4362);
and U4554 (N_4554,N_4116,N_4463);
or U4555 (N_4555,N_4086,N_4464);
nand U4556 (N_4556,N_4162,N_4418);
and U4557 (N_4557,N_4130,N_4017);
nand U4558 (N_4558,N_4213,N_4244);
or U4559 (N_4559,N_4235,N_4209);
or U4560 (N_4560,N_4161,N_4106);
nor U4561 (N_4561,N_4047,N_4128);
or U4562 (N_4562,N_4474,N_4348);
and U4563 (N_4563,N_4100,N_4428);
and U4564 (N_4564,N_4319,N_4334);
and U4565 (N_4565,N_4377,N_4120);
nand U4566 (N_4566,N_4268,N_4240);
or U4567 (N_4567,N_4483,N_4271);
or U4568 (N_4568,N_4002,N_4056);
nand U4569 (N_4569,N_4186,N_4067);
or U4570 (N_4570,N_4274,N_4350);
nand U4571 (N_4571,N_4349,N_4090);
nand U4572 (N_4572,N_4476,N_4499);
nor U4573 (N_4573,N_4179,N_4151);
and U4574 (N_4574,N_4168,N_4332);
nor U4575 (N_4575,N_4003,N_4000);
or U4576 (N_4576,N_4234,N_4328);
nor U4577 (N_4577,N_4147,N_4225);
nor U4578 (N_4578,N_4195,N_4343);
nand U4579 (N_4579,N_4105,N_4331);
and U4580 (N_4580,N_4009,N_4131);
and U4581 (N_4581,N_4389,N_4001);
nor U4582 (N_4582,N_4446,N_4457);
nand U4583 (N_4583,N_4160,N_4059);
or U4584 (N_4584,N_4063,N_4311);
nor U4585 (N_4585,N_4387,N_4034);
and U4586 (N_4586,N_4437,N_4293);
nand U4587 (N_4587,N_4218,N_4462);
nor U4588 (N_4588,N_4351,N_4353);
nor U4589 (N_4589,N_4253,N_4370);
nand U4590 (N_4590,N_4187,N_4044);
nor U4591 (N_4591,N_4431,N_4145);
nand U4592 (N_4592,N_4135,N_4230);
nor U4593 (N_4593,N_4489,N_4083);
nor U4594 (N_4594,N_4496,N_4261);
nand U4595 (N_4595,N_4307,N_4391);
or U4596 (N_4596,N_4136,N_4118);
nor U4597 (N_4597,N_4254,N_4490);
and U4598 (N_4598,N_4108,N_4078);
nor U4599 (N_4599,N_4405,N_4072);
nand U4600 (N_4600,N_4396,N_4306);
or U4601 (N_4601,N_4073,N_4318);
nor U4602 (N_4602,N_4325,N_4156);
nor U4603 (N_4603,N_4382,N_4027);
and U4604 (N_4604,N_4250,N_4185);
and U4605 (N_4605,N_4258,N_4101);
nor U4606 (N_4606,N_4447,N_4223);
nand U4607 (N_4607,N_4436,N_4084);
nor U4608 (N_4608,N_4216,N_4342);
or U4609 (N_4609,N_4226,N_4122);
or U4610 (N_4610,N_4004,N_4444);
and U4611 (N_4611,N_4115,N_4440);
and U4612 (N_4612,N_4365,N_4159);
and U4613 (N_4613,N_4256,N_4190);
or U4614 (N_4614,N_4414,N_4144);
nand U4615 (N_4615,N_4094,N_4251);
nor U4616 (N_4616,N_4089,N_4035);
or U4617 (N_4617,N_4219,N_4255);
or U4618 (N_4618,N_4322,N_4018);
xor U4619 (N_4619,N_4320,N_4200);
nand U4620 (N_4620,N_4171,N_4421);
nor U4621 (N_4621,N_4012,N_4184);
nand U4622 (N_4622,N_4498,N_4025);
nand U4623 (N_4623,N_4233,N_4289);
and U4624 (N_4624,N_4191,N_4398);
or U4625 (N_4625,N_4275,N_4280);
nand U4626 (N_4626,N_4207,N_4303);
and U4627 (N_4627,N_4381,N_4043);
nand U4628 (N_4628,N_4448,N_4409);
or U4629 (N_4629,N_4085,N_4222);
nor U4630 (N_4630,N_4060,N_4198);
nor U4631 (N_4631,N_4257,N_4142);
or U4632 (N_4632,N_4410,N_4245);
nor U4633 (N_4633,N_4315,N_4316);
nand U4634 (N_4634,N_4020,N_4417);
nand U4635 (N_4635,N_4344,N_4049);
nor U4636 (N_4636,N_4181,N_4390);
and U4637 (N_4637,N_4329,N_4087);
nor U4638 (N_4638,N_4402,N_4369);
and U4639 (N_4639,N_4459,N_4174);
nor U4640 (N_4640,N_4110,N_4450);
nor U4641 (N_4641,N_4140,N_4286);
nand U4642 (N_4642,N_4363,N_4252);
or U4643 (N_4643,N_4103,N_4074);
or U4644 (N_4644,N_4341,N_4263);
nor U4645 (N_4645,N_4384,N_4291);
nor U4646 (N_4646,N_4339,N_4124);
nor U4647 (N_4647,N_4472,N_4175);
and U4648 (N_4648,N_4134,N_4229);
and U4649 (N_4649,N_4138,N_4228);
nand U4650 (N_4650,N_4170,N_4301);
nor U4651 (N_4651,N_4071,N_4281);
nor U4652 (N_4652,N_4361,N_4081);
or U4653 (N_4653,N_4069,N_4150);
and U4654 (N_4654,N_4227,N_4355);
nor U4655 (N_4655,N_4133,N_4276);
or U4656 (N_4656,N_4132,N_4497);
and U4657 (N_4657,N_4285,N_4054);
and U4658 (N_4658,N_4337,N_4164);
or U4659 (N_4659,N_4336,N_4183);
or U4660 (N_4660,N_4068,N_4477);
or U4661 (N_4661,N_4443,N_4091);
and U4662 (N_4662,N_4050,N_4206);
or U4663 (N_4663,N_4367,N_4211);
and U4664 (N_4664,N_4374,N_4269);
nor U4665 (N_4665,N_4031,N_4434);
and U4666 (N_4666,N_4445,N_4158);
and U4667 (N_4667,N_4005,N_4204);
and U4668 (N_4668,N_4451,N_4137);
and U4669 (N_4669,N_4468,N_4340);
and U4670 (N_4670,N_4495,N_4479);
or U4671 (N_4671,N_4077,N_4260);
nor U4672 (N_4672,N_4061,N_4298);
and U4673 (N_4673,N_4177,N_4082);
nor U4674 (N_4674,N_4454,N_4172);
nand U4675 (N_4675,N_4292,N_4294);
nand U4676 (N_4676,N_4290,N_4399);
and U4677 (N_4677,N_4075,N_4475);
and U4678 (N_4678,N_4231,N_4192);
nand U4679 (N_4679,N_4221,N_4248);
nand U4680 (N_4680,N_4052,N_4129);
nor U4681 (N_4681,N_4169,N_4215);
nor U4682 (N_4682,N_4038,N_4021);
and U4683 (N_4683,N_4264,N_4178);
or U4684 (N_4684,N_4013,N_4423);
nor U4685 (N_4685,N_4194,N_4453);
nor U4686 (N_4686,N_4404,N_4146);
or U4687 (N_4687,N_4166,N_4383);
and U4688 (N_4688,N_4397,N_4282);
and U4689 (N_4689,N_4284,N_4080);
or U4690 (N_4690,N_4155,N_4189);
nand U4691 (N_4691,N_4360,N_4139);
or U4692 (N_4692,N_4024,N_4148);
nor U4693 (N_4693,N_4338,N_4471);
or U4694 (N_4694,N_4300,N_4193);
nor U4695 (N_4695,N_4107,N_4095);
and U4696 (N_4696,N_4039,N_4014);
or U4697 (N_4697,N_4220,N_4143);
nand U4698 (N_4698,N_4486,N_4079);
nor U4699 (N_4699,N_4466,N_4379);
or U4700 (N_4700,N_4313,N_4346);
or U4701 (N_4701,N_4119,N_4113);
and U4702 (N_4702,N_4066,N_4030);
or U4703 (N_4703,N_4287,N_4032);
or U4704 (N_4704,N_4057,N_4407);
and U4705 (N_4705,N_4452,N_4376);
and U4706 (N_4706,N_4241,N_4321);
nand U4707 (N_4707,N_4070,N_4062);
and U4708 (N_4708,N_4395,N_4330);
nor U4709 (N_4709,N_4297,N_4295);
or U4710 (N_4710,N_4259,N_4449);
nand U4711 (N_4711,N_4109,N_4357);
nor U4712 (N_4712,N_4371,N_4465);
and U4713 (N_4713,N_4173,N_4266);
or U4714 (N_4714,N_4308,N_4441);
or U4715 (N_4715,N_4099,N_4296);
nand U4716 (N_4716,N_4055,N_4411);
or U4717 (N_4717,N_4359,N_4188);
xnor U4718 (N_4718,N_4442,N_4427);
nand U4719 (N_4719,N_4019,N_4088);
and U4720 (N_4720,N_4438,N_4114);
and U4721 (N_4721,N_4420,N_4354);
or U4722 (N_4722,N_4485,N_4288);
or U4723 (N_4723,N_4065,N_4205);
or U4724 (N_4724,N_4033,N_4272);
nand U4725 (N_4725,N_4406,N_4097);
or U4726 (N_4726,N_4249,N_4456);
and U4727 (N_4727,N_4310,N_4203);
and U4728 (N_4728,N_4015,N_4036);
nor U4729 (N_4729,N_4093,N_4045);
and U4730 (N_4730,N_4314,N_4270);
nand U4731 (N_4731,N_4196,N_4058);
xnor U4732 (N_4732,N_4165,N_4323);
nand U4733 (N_4733,N_4366,N_4197);
or U4734 (N_4734,N_4435,N_4127);
or U4735 (N_4735,N_4432,N_4493);
nor U4736 (N_4736,N_4042,N_4394);
nor U4737 (N_4737,N_4123,N_4309);
nor U4738 (N_4738,N_4378,N_4201);
or U4739 (N_4739,N_4425,N_4029);
nand U4740 (N_4740,N_4426,N_4208);
nor U4741 (N_4741,N_4372,N_4167);
nand U4742 (N_4742,N_4051,N_4375);
and U4743 (N_4743,N_4064,N_4386);
or U4744 (N_4744,N_4333,N_4439);
nand U4745 (N_4745,N_4210,N_4416);
nor U4746 (N_4746,N_4010,N_4262);
and U4747 (N_4747,N_4046,N_4022);
nand U4748 (N_4748,N_4279,N_4111);
nor U4749 (N_4749,N_4202,N_4487);
nand U4750 (N_4750,N_4105,N_4086);
nand U4751 (N_4751,N_4113,N_4153);
nand U4752 (N_4752,N_4032,N_4427);
nand U4753 (N_4753,N_4254,N_4402);
and U4754 (N_4754,N_4475,N_4287);
xnor U4755 (N_4755,N_4343,N_4364);
nor U4756 (N_4756,N_4209,N_4325);
nand U4757 (N_4757,N_4114,N_4155);
and U4758 (N_4758,N_4064,N_4447);
nor U4759 (N_4759,N_4240,N_4134);
or U4760 (N_4760,N_4246,N_4224);
nand U4761 (N_4761,N_4234,N_4331);
nand U4762 (N_4762,N_4145,N_4243);
nor U4763 (N_4763,N_4384,N_4043);
nor U4764 (N_4764,N_4185,N_4360);
nor U4765 (N_4765,N_4169,N_4364);
and U4766 (N_4766,N_4243,N_4121);
nor U4767 (N_4767,N_4379,N_4343);
nand U4768 (N_4768,N_4402,N_4171);
and U4769 (N_4769,N_4380,N_4289);
or U4770 (N_4770,N_4055,N_4112);
nor U4771 (N_4771,N_4326,N_4136);
or U4772 (N_4772,N_4405,N_4079);
nor U4773 (N_4773,N_4390,N_4266);
nand U4774 (N_4774,N_4003,N_4251);
and U4775 (N_4775,N_4144,N_4107);
or U4776 (N_4776,N_4250,N_4311);
and U4777 (N_4777,N_4097,N_4373);
nor U4778 (N_4778,N_4059,N_4283);
nand U4779 (N_4779,N_4488,N_4154);
or U4780 (N_4780,N_4237,N_4016);
nor U4781 (N_4781,N_4177,N_4362);
nand U4782 (N_4782,N_4031,N_4448);
nand U4783 (N_4783,N_4319,N_4409);
or U4784 (N_4784,N_4411,N_4499);
and U4785 (N_4785,N_4496,N_4013);
nor U4786 (N_4786,N_4464,N_4100);
nor U4787 (N_4787,N_4097,N_4158);
and U4788 (N_4788,N_4443,N_4322);
nor U4789 (N_4789,N_4277,N_4457);
nand U4790 (N_4790,N_4358,N_4195);
nor U4791 (N_4791,N_4456,N_4430);
or U4792 (N_4792,N_4321,N_4397);
nor U4793 (N_4793,N_4116,N_4008);
or U4794 (N_4794,N_4208,N_4195);
nor U4795 (N_4795,N_4306,N_4403);
nor U4796 (N_4796,N_4388,N_4153);
nor U4797 (N_4797,N_4363,N_4045);
nand U4798 (N_4798,N_4351,N_4478);
and U4799 (N_4799,N_4110,N_4391);
nand U4800 (N_4800,N_4255,N_4438);
or U4801 (N_4801,N_4473,N_4399);
or U4802 (N_4802,N_4108,N_4048);
nand U4803 (N_4803,N_4208,N_4140);
nor U4804 (N_4804,N_4474,N_4035);
and U4805 (N_4805,N_4041,N_4259);
or U4806 (N_4806,N_4311,N_4233);
nor U4807 (N_4807,N_4138,N_4434);
nand U4808 (N_4808,N_4225,N_4122);
nor U4809 (N_4809,N_4131,N_4214);
or U4810 (N_4810,N_4002,N_4155);
nor U4811 (N_4811,N_4487,N_4306);
nor U4812 (N_4812,N_4226,N_4377);
or U4813 (N_4813,N_4005,N_4199);
nor U4814 (N_4814,N_4189,N_4456);
nand U4815 (N_4815,N_4097,N_4137);
or U4816 (N_4816,N_4425,N_4377);
nor U4817 (N_4817,N_4335,N_4374);
or U4818 (N_4818,N_4232,N_4107);
nor U4819 (N_4819,N_4023,N_4278);
and U4820 (N_4820,N_4114,N_4242);
and U4821 (N_4821,N_4469,N_4126);
nand U4822 (N_4822,N_4033,N_4248);
nand U4823 (N_4823,N_4255,N_4459);
or U4824 (N_4824,N_4208,N_4087);
nor U4825 (N_4825,N_4056,N_4174);
nor U4826 (N_4826,N_4051,N_4324);
and U4827 (N_4827,N_4336,N_4151);
nand U4828 (N_4828,N_4132,N_4125);
nor U4829 (N_4829,N_4413,N_4251);
nand U4830 (N_4830,N_4247,N_4101);
or U4831 (N_4831,N_4048,N_4277);
and U4832 (N_4832,N_4173,N_4058);
or U4833 (N_4833,N_4411,N_4131);
nor U4834 (N_4834,N_4358,N_4043);
and U4835 (N_4835,N_4325,N_4467);
or U4836 (N_4836,N_4006,N_4404);
and U4837 (N_4837,N_4174,N_4119);
nor U4838 (N_4838,N_4393,N_4311);
nor U4839 (N_4839,N_4400,N_4355);
nor U4840 (N_4840,N_4304,N_4263);
nand U4841 (N_4841,N_4255,N_4046);
nand U4842 (N_4842,N_4093,N_4161);
and U4843 (N_4843,N_4240,N_4499);
or U4844 (N_4844,N_4375,N_4104);
or U4845 (N_4845,N_4388,N_4056);
nand U4846 (N_4846,N_4147,N_4358);
nor U4847 (N_4847,N_4248,N_4352);
and U4848 (N_4848,N_4350,N_4308);
nor U4849 (N_4849,N_4369,N_4317);
or U4850 (N_4850,N_4353,N_4062);
nor U4851 (N_4851,N_4190,N_4084);
or U4852 (N_4852,N_4150,N_4051);
nand U4853 (N_4853,N_4426,N_4179);
or U4854 (N_4854,N_4403,N_4140);
and U4855 (N_4855,N_4011,N_4133);
and U4856 (N_4856,N_4333,N_4487);
and U4857 (N_4857,N_4085,N_4499);
nor U4858 (N_4858,N_4399,N_4169);
or U4859 (N_4859,N_4360,N_4143);
nand U4860 (N_4860,N_4010,N_4431);
nand U4861 (N_4861,N_4147,N_4406);
or U4862 (N_4862,N_4278,N_4292);
nor U4863 (N_4863,N_4413,N_4215);
nand U4864 (N_4864,N_4279,N_4213);
nor U4865 (N_4865,N_4144,N_4058);
nor U4866 (N_4866,N_4486,N_4270);
and U4867 (N_4867,N_4478,N_4467);
or U4868 (N_4868,N_4255,N_4258);
nor U4869 (N_4869,N_4141,N_4223);
or U4870 (N_4870,N_4427,N_4181);
or U4871 (N_4871,N_4225,N_4452);
nand U4872 (N_4872,N_4070,N_4114);
nor U4873 (N_4873,N_4181,N_4260);
nor U4874 (N_4874,N_4072,N_4451);
xor U4875 (N_4875,N_4074,N_4213);
and U4876 (N_4876,N_4275,N_4382);
xnor U4877 (N_4877,N_4462,N_4094);
nor U4878 (N_4878,N_4072,N_4454);
and U4879 (N_4879,N_4154,N_4492);
and U4880 (N_4880,N_4139,N_4197);
nor U4881 (N_4881,N_4203,N_4190);
and U4882 (N_4882,N_4322,N_4247);
or U4883 (N_4883,N_4114,N_4131);
nor U4884 (N_4884,N_4078,N_4427);
and U4885 (N_4885,N_4011,N_4096);
or U4886 (N_4886,N_4111,N_4293);
nand U4887 (N_4887,N_4131,N_4478);
and U4888 (N_4888,N_4007,N_4281);
or U4889 (N_4889,N_4366,N_4249);
or U4890 (N_4890,N_4354,N_4201);
nand U4891 (N_4891,N_4350,N_4278);
nand U4892 (N_4892,N_4034,N_4215);
nand U4893 (N_4893,N_4009,N_4362);
and U4894 (N_4894,N_4491,N_4262);
and U4895 (N_4895,N_4410,N_4430);
nand U4896 (N_4896,N_4011,N_4369);
nor U4897 (N_4897,N_4356,N_4287);
or U4898 (N_4898,N_4072,N_4426);
or U4899 (N_4899,N_4008,N_4487);
and U4900 (N_4900,N_4454,N_4135);
and U4901 (N_4901,N_4499,N_4482);
xor U4902 (N_4902,N_4359,N_4439);
nor U4903 (N_4903,N_4393,N_4253);
nand U4904 (N_4904,N_4423,N_4271);
or U4905 (N_4905,N_4445,N_4287);
or U4906 (N_4906,N_4115,N_4435);
and U4907 (N_4907,N_4078,N_4383);
nor U4908 (N_4908,N_4056,N_4284);
nor U4909 (N_4909,N_4345,N_4018);
or U4910 (N_4910,N_4425,N_4128);
nor U4911 (N_4911,N_4293,N_4292);
nor U4912 (N_4912,N_4448,N_4066);
or U4913 (N_4913,N_4006,N_4182);
or U4914 (N_4914,N_4153,N_4105);
nand U4915 (N_4915,N_4491,N_4413);
nor U4916 (N_4916,N_4405,N_4131);
nor U4917 (N_4917,N_4193,N_4191);
nand U4918 (N_4918,N_4317,N_4281);
or U4919 (N_4919,N_4134,N_4293);
and U4920 (N_4920,N_4054,N_4287);
and U4921 (N_4921,N_4055,N_4008);
nand U4922 (N_4922,N_4041,N_4258);
and U4923 (N_4923,N_4235,N_4244);
or U4924 (N_4924,N_4360,N_4365);
nand U4925 (N_4925,N_4367,N_4240);
nor U4926 (N_4926,N_4059,N_4415);
and U4927 (N_4927,N_4189,N_4111);
and U4928 (N_4928,N_4181,N_4001);
and U4929 (N_4929,N_4137,N_4337);
and U4930 (N_4930,N_4239,N_4172);
nor U4931 (N_4931,N_4195,N_4025);
nand U4932 (N_4932,N_4031,N_4215);
nand U4933 (N_4933,N_4004,N_4040);
nand U4934 (N_4934,N_4145,N_4116);
or U4935 (N_4935,N_4178,N_4346);
nor U4936 (N_4936,N_4104,N_4143);
or U4937 (N_4937,N_4261,N_4184);
and U4938 (N_4938,N_4133,N_4436);
nor U4939 (N_4939,N_4055,N_4278);
and U4940 (N_4940,N_4448,N_4256);
or U4941 (N_4941,N_4413,N_4446);
or U4942 (N_4942,N_4384,N_4018);
and U4943 (N_4943,N_4055,N_4477);
nand U4944 (N_4944,N_4056,N_4096);
or U4945 (N_4945,N_4029,N_4115);
and U4946 (N_4946,N_4134,N_4464);
nor U4947 (N_4947,N_4363,N_4240);
and U4948 (N_4948,N_4454,N_4079);
and U4949 (N_4949,N_4058,N_4250);
nand U4950 (N_4950,N_4462,N_4448);
nor U4951 (N_4951,N_4077,N_4370);
and U4952 (N_4952,N_4362,N_4308);
or U4953 (N_4953,N_4384,N_4235);
and U4954 (N_4954,N_4421,N_4032);
or U4955 (N_4955,N_4154,N_4106);
nand U4956 (N_4956,N_4343,N_4446);
nand U4957 (N_4957,N_4100,N_4354);
nor U4958 (N_4958,N_4285,N_4290);
nor U4959 (N_4959,N_4322,N_4049);
nor U4960 (N_4960,N_4248,N_4373);
nand U4961 (N_4961,N_4052,N_4440);
and U4962 (N_4962,N_4046,N_4035);
and U4963 (N_4963,N_4470,N_4370);
or U4964 (N_4964,N_4104,N_4141);
nand U4965 (N_4965,N_4004,N_4121);
nand U4966 (N_4966,N_4463,N_4045);
and U4967 (N_4967,N_4428,N_4364);
or U4968 (N_4968,N_4008,N_4171);
or U4969 (N_4969,N_4189,N_4186);
nor U4970 (N_4970,N_4182,N_4120);
or U4971 (N_4971,N_4234,N_4064);
and U4972 (N_4972,N_4341,N_4251);
nor U4973 (N_4973,N_4298,N_4324);
nor U4974 (N_4974,N_4000,N_4437);
nand U4975 (N_4975,N_4419,N_4333);
nor U4976 (N_4976,N_4315,N_4469);
nand U4977 (N_4977,N_4203,N_4292);
or U4978 (N_4978,N_4408,N_4225);
and U4979 (N_4979,N_4167,N_4102);
nand U4980 (N_4980,N_4433,N_4377);
nand U4981 (N_4981,N_4292,N_4326);
nand U4982 (N_4982,N_4299,N_4241);
nor U4983 (N_4983,N_4034,N_4419);
nand U4984 (N_4984,N_4246,N_4035);
or U4985 (N_4985,N_4254,N_4271);
or U4986 (N_4986,N_4307,N_4016);
or U4987 (N_4987,N_4180,N_4459);
and U4988 (N_4988,N_4411,N_4092);
nand U4989 (N_4989,N_4266,N_4322);
nor U4990 (N_4990,N_4198,N_4444);
or U4991 (N_4991,N_4001,N_4465);
and U4992 (N_4992,N_4382,N_4235);
and U4993 (N_4993,N_4223,N_4450);
nand U4994 (N_4994,N_4052,N_4090);
and U4995 (N_4995,N_4417,N_4013);
nor U4996 (N_4996,N_4224,N_4417);
nor U4997 (N_4997,N_4092,N_4392);
and U4998 (N_4998,N_4060,N_4337);
and U4999 (N_4999,N_4415,N_4085);
nor UO_0 (O_0,N_4996,N_4588);
or UO_1 (O_1,N_4838,N_4575);
nand UO_2 (O_2,N_4849,N_4783);
nor UO_3 (O_3,N_4720,N_4995);
or UO_4 (O_4,N_4816,N_4916);
nor UO_5 (O_5,N_4609,N_4704);
nand UO_6 (O_6,N_4794,N_4504);
nand UO_7 (O_7,N_4961,N_4812);
or UO_8 (O_8,N_4876,N_4625);
and UO_9 (O_9,N_4556,N_4841);
or UO_10 (O_10,N_4760,N_4569);
or UO_11 (O_11,N_4617,N_4712);
or UO_12 (O_12,N_4831,N_4796);
nand UO_13 (O_13,N_4857,N_4553);
and UO_14 (O_14,N_4748,N_4790);
nor UO_15 (O_15,N_4566,N_4829);
nand UO_16 (O_16,N_4886,N_4533);
nand UO_17 (O_17,N_4848,N_4826);
nor UO_18 (O_18,N_4589,N_4837);
nand UO_19 (O_19,N_4864,N_4576);
or UO_20 (O_20,N_4906,N_4510);
nand UO_21 (O_21,N_4847,N_4820);
nand UO_22 (O_22,N_4986,N_4762);
nand UO_23 (O_23,N_4622,N_4516);
or UO_24 (O_24,N_4726,N_4536);
nand UO_25 (O_25,N_4804,N_4844);
nand UO_26 (O_26,N_4861,N_4677);
nor UO_27 (O_27,N_4535,N_4978);
or UO_28 (O_28,N_4866,N_4949);
nand UO_29 (O_29,N_4803,N_4500);
or UO_30 (O_30,N_4945,N_4613);
nor UO_31 (O_31,N_4813,N_4534);
nor UO_32 (O_32,N_4667,N_4738);
or UO_33 (O_33,N_4618,N_4614);
nor UO_34 (O_34,N_4686,N_4843);
nand UO_35 (O_35,N_4963,N_4714);
nor UO_36 (O_36,N_4842,N_4532);
or UO_37 (O_37,N_4921,N_4811);
or UO_38 (O_38,N_4942,N_4970);
nor UO_39 (O_39,N_4935,N_4962);
nand UO_40 (O_40,N_4641,N_4693);
nand UO_41 (O_41,N_4854,N_4604);
or UO_42 (O_42,N_4889,N_4513);
nor UO_43 (O_43,N_4845,N_4885);
nand UO_44 (O_44,N_4694,N_4756);
nor UO_45 (O_45,N_4526,N_4665);
nand UO_46 (O_46,N_4926,N_4587);
nand UO_47 (O_47,N_4934,N_4666);
or UO_48 (O_48,N_4980,N_4967);
nor UO_49 (O_49,N_4636,N_4508);
and UO_50 (O_50,N_4697,N_4674);
nor UO_51 (O_51,N_4759,N_4994);
or UO_52 (O_52,N_4596,N_4805);
nand UO_53 (O_53,N_4913,N_4543);
nand UO_54 (O_54,N_4769,N_4912);
nor UO_55 (O_55,N_4895,N_4542);
nor UO_56 (O_56,N_4800,N_4633);
and UO_57 (O_57,N_4672,N_4715);
and UO_58 (O_58,N_4593,N_4778);
nor UO_59 (O_59,N_4993,N_4809);
and UO_60 (O_60,N_4668,N_4767);
nand UO_61 (O_61,N_4839,N_4872);
and UO_62 (O_62,N_4541,N_4675);
nand UO_63 (O_63,N_4632,N_4966);
and UO_64 (O_64,N_4975,N_4595);
nor UO_65 (O_65,N_4867,N_4890);
or UO_66 (O_66,N_4821,N_4643);
or UO_67 (O_67,N_4834,N_4631);
nor UO_68 (O_68,N_4528,N_4621);
or UO_69 (O_69,N_4554,N_4741);
nand UO_70 (O_70,N_4620,N_4571);
and UO_71 (O_71,N_4691,N_4507);
or UO_72 (O_72,N_4955,N_4865);
nor UO_73 (O_73,N_4608,N_4771);
nor UO_74 (O_74,N_4538,N_4754);
nor UO_75 (O_75,N_4773,N_4888);
and UO_76 (O_76,N_4789,N_4819);
nand UO_77 (O_77,N_4957,N_4860);
or UO_78 (O_78,N_4870,N_4544);
or UO_79 (O_79,N_4574,N_4882);
and UO_80 (O_80,N_4898,N_4551);
nand UO_81 (O_81,N_4965,N_4736);
nor UO_82 (O_82,N_4925,N_4808);
and UO_83 (O_83,N_4582,N_4594);
and UO_84 (O_84,N_4573,N_4937);
and UO_85 (O_85,N_4652,N_4610);
and UO_86 (O_86,N_4717,N_4518);
nand UO_87 (O_87,N_4522,N_4501);
nand UO_88 (O_88,N_4519,N_4629);
and UO_89 (O_89,N_4581,N_4933);
or UO_90 (O_90,N_4563,N_4817);
or UO_91 (O_91,N_4973,N_4892);
or UO_92 (O_92,N_4655,N_4863);
nor UO_93 (O_93,N_4572,N_4810);
nor UO_94 (O_94,N_4883,N_4584);
nor UO_95 (O_95,N_4787,N_4752);
and UO_96 (O_96,N_4798,N_4700);
or UO_97 (O_97,N_4701,N_4706);
or UO_98 (O_98,N_4710,N_4703);
and UO_99 (O_99,N_4974,N_4689);
or UO_100 (O_100,N_4678,N_4559);
nand UO_101 (O_101,N_4776,N_4683);
nor UO_102 (O_102,N_4830,N_4537);
nand UO_103 (O_103,N_4705,N_4669);
and UO_104 (O_104,N_4590,N_4658);
nand UO_105 (O_105,N_4661,N_4530);
nor UO_106 (O_106,N_4681,N_4733);
nand UO_107 (O_107,N_4753,N_4750);
nand UO_108 (O_108,N_4976,N_4585);
or UO_109 (O_109,N_4684,N_4793);
nor UO_110 (O_110,N_4646,N_4903);
nor UO_111 (O_111,N_4568,N_4662);
and UO_112 (O_112,N_4887,N_4984);
or UO_113 (O_113,N_4971,N_4982);
or UO_114 (O_114,N_4799,N_4567);
and UO_115 (O_115,N_4727,N_4987);
nor UO_116 (O_116,N_4941,N_4648);
nand UO_117 (O_117,N_4840,N_4988);
nor UO_118 (O_118,N_4827,N_4531);
nor UO_119 (O_119,N_4555,N_4517);
or UO_120 (O_120,N_4539,N_4868);
and UO_121 (O_121,N_4599,N_4774);
nand UO_122 (O_122,N_4605,N_4619);
or UO_123 (O_123,N_4832,N_4807);
nor UO_124 (O_124,N_4852,N_4899);
and UO_125 (O_125,N_4524,N_4664);
nor UO_126 (O_126,N_4547,N_4877);
or UO_127 (O_127,N_4953,N_4671);
nand UO_128 (O_128,N_4992,N_4644);
or UO_129 (O_129,N_4924,N_4855);
and UO_130 (O_130,N_4846,N_4959);
nor UO_131 (O_131,N_4969,N_4749);
and UO_132 (O_132,N_4611,N_4818);
nor UO_133 (O_133,N_4936,N_4999);
nand UO_134 (O_134,N_4977,N_4801);
nor UO_135 (O_135,N_4914,N_4891);
nor UO_136 (O_136,N_4732,N_4972);
and UO_137 (O_137,N_4859,N_4873);
and UO_138 (O_138,N_4502,N_4651);
or UO_139 (O_139,N_4964,N_4910);
and UO_140 (O_140,N_4660,N_4509);
nor UO_141 (O_141,N_4875,N_4853);
or UO_142 (O_142,N_4637,N_4731);
nor UO_143 (O_143,N_4772,N_4932);
nand UO_144 (O_144,N_4591,N_4670);
nor UO_145 (O_145,N_4792,N_4673);
nor UO_146 (O_146,N_4952,N_4983);
nand UO_147 (O_147,N_4645,N_4728);
or UO_148 (O_148,N_4784,N_4918);
nor UO_149 (O_149,N_4757,N_4630);
or UO_150 (O_150,N_4869,N_4920);
nor UO_151 (O_151,N_4968,N_4521);
nand UO_152 (O_152,N_4552,N_4751);
nor UO_153 (O_153,N_4602,N_4721);
nand UO_154 (O_154,N_4549,N_4739);
and UO_155 (O_155,N_4985,N_4525);
and UO_156 (O_156,N_4682,N_4833);
or UO_157 (O_157,N_4598,N_4881);
and UO_158 (O_158,N_4862,N_4814);
or UO_159 (O_159,N_4612,N_4785);
or UO_160 (O_160,N_4586,N_4725);
nor UO_161 (O_161,N_4825,N_4911);
or UO_162 (O_162,N_4561,N_4676);
nor UO_163 (O_163,N_4765,N_4615);
and UO_164 (O_164,N_4835,N_4577);
or UO_165 (O_165,N_4640,N_4506);
nor UO_166 (O_166,N_4989,N_4687);
nor UO_167 (O_167,N_4879,N_4742);
or UO_168 (O_168,N_4780,N_4740);
nor UO_169 (O_169,N_4558,N_4940);
or UO_170 (O_170,N_4616,N_4824);
nor UO_171 (O_171,N_4763,N_4806);
nor UO_172 (O_172,N_4919,N_4624);
or UO_173 (O_173,N_4929,N_4943);
or UO_174 (O_174,N_4514,N_4680);
or UO_175 (O_175,N_4570,N_4529);
nand UO_176 (O_176,N_4896,N_4729);
nor UO_177 (O_177,N_4579,N_4696);
nor UO_178 (O_178,N_4761,N_4902);
nand UO_179 (O_179,N_4850,N_4690);
and UO_180 (O_180,N_4894,N_4909);
and UO_181 (O_181,N_4540,N_4991);
nand UO_182 (O_182,N_4557,N_4716);
or UO_183 (O_183,N_4901,N_4564);
nor UO_184 (O_184,N_4947,N_4546);
or UO_185 (O_185,N_4997,N_4626);
nand UO_186 (O_186,N_4822,N_4642);
nand UO_187 (O_187,N_4634,N_4795);
nor UO_188 (O_188,N_4638,N_4927);
nand UO_189 (O_189,N_4764,N_4639);
nand UO_190 (O_190,N_4702,N_4583);
nand UO_191 (O_191,N_4663,N_4659);
nand UO_192 (O_192,N_4950,N_4592);
nor UO_193 (O_193,N_4915,N_4709);
or UO_194 (O_194,N_4656,N_4874);
or UO_195 (O_195,N_4730,N_4708);
and UO_196 (O_196,N_4743,N_4951);
or UO_197 (O_197,N_4930,N_4944);
nand UO_198 (O_198,N_4900,N_4755);
or UO_199 (O_199,N_4922,N_4550);
or UO_200 (O_200,N_4711,N_4685);
and UO_201 (O_201,N_4600,N_4503);
or UO_202 (O_202,N_4719,N_4956);
nand UO_203 (O_203,N_4722,N_4979);
nand UO_204 (O_204,N_4657,N_4623);
nor UO_205 (O_205,N_4923,N_4758);
and UO_206 (O_206,N_4523,N_4565);
nand UO_207 (O_207,N_4578,N_4905);
nor UO_208 (O_208,N_4828,N_4907);
and UO_209 (O_209,N_4635,N_4699);
or UO_210 (O_210,N_4836,N_4695);
nand UO_211 (O_211,N_4858,N_4948);
nand UO_212 (O_212,N_4724,N_4946);
and UO_213 (O_213,N_4908,N_4737);
or UO_214 (O_214,N_4960,N_4654);
nor UO_215 (O_215,N_4647,N_4745);
nor UO_216 (O_216,N_4515,N_4545);
or UO_217 (O_217,N_4904,N_4791);
nor UO_218 (O_218,N_4893,N_4768);
and UO_219 (O_219,N_4628,N_4878);
and UO_220 (O_220,N_4823,N_4580);
nand UO_221 (O_221,N_4746,N_4786);
nand UO_222 (O_222,N_4815,N_4802);
nor UO_223 (O_223,N_4884,N_4562);
and UO_224 (O_224,N_4601,N_4770);
nor UO_225 (O_225,N_4527,N_4981);
nand UO_226 (O_226,N_4505,N_4998);
and UO_227 (O_227,N_4931,N_4851);
or UO_228 (O_228,N_4679,N_4653);
or UO_229 (O_229,N_4781,N_4775);
nand UO_230 (O_230,N_4698,N_4744);
and UO_231 (O_231,N_4954,N_4707);
or UO_232 (O_232,N_4928,N_4606);
nand UO_233 (O_233,N_4782,N_4990);
nand UO_234 (O_234,N_4650,N_4603);
or UO_235 (O_235,N_4871,N_4788);
nand UO_236 (O_236,N_4779,N_4692);
or UO_237 (O_237,N_4880,N_4511);
nor UO_238 (O_238,N_4856,N_4607);
or UO_239 (O_239,N_4797,N_4777);
nand UO_240 (O_240,N_4718,N_4723);
or UO_241 (O_241,N_4649,N_4939);
or UO_242 (O_242,N_4627,N_4713);
nand UO_243 (O_243,N_4917,N_4735);
nor UO_244 (O_244,N_4512,N_4958);
nand UO_245 (O_245,N_4747,N_4597);
nor UO_246 (O_246,N_4897,N_4734);
nand UO_247 (O_247,N_4520,N_4560);
nand UO_248 (O_248,N_4766,N_4688);
or UO_249 (O_249,N_4938,N_4548);
nand UO_250 (O_250,N_4734,N_4887);
nor UO_251 (O_251,N_4996,N_4562);
nand UO_252 (O_252,N_4814,N_4799);
nand UO_253 (O_253,N_4517,N_4756);
or UO_254 (O_254,N_4574,N_4808);
or UO_255 (O_255,N_4686,N_4617);
and UO_256 (O_256,N_4680,N_4890);
nand UO_257 (O_257,N_4668,N_4954);
nor UO_258 (O_258,N_4911,N_4945);
nand UO_259 (O_259,N_4659,N_4777);
nand UO_260 (O_260,N_4534,N_4892);
nor UO_261 (O_261,N_4730,N_4740);
nor UO_262 (O_262,N_4978,N_4675);
or UO_263 (O_263,N_4581,N_4785);
nor UO_264 (O_264,N_4666,N_4769);
nand UO_265 (O_265,N_4707,N_4722);
nand UO_266 (O_266,N_4856,N_4546);
nand UO_267 (O_267,N_4612,N_4956);
and UO_268 (O_268,N_4571,N_4894);
and UO_269 (O_269,N_4982,N_4521);
nand UO_270 (O_270,N_4647,N_4754);
nand UO_271 (O_271,N_4549,N_4900);
nor UO_272 (O_272,N_4637,N_4833);
xnor UO_273 (O_273,N_4953,N_4702);
or UO_274 (O_274,N_4504,N_4981);
nor UO_275 (O_275,N_4852,N_4990);
nor UO_276 (O_276,N_4626,N_4958);
nor UO_277 (O_277,N_4684,N_4619);
or UO_278 (O_278,N_4756,N_4862);
or UO_279 (O_279,N_4530,N_4565);
nor UO_280 (O_280,N_4804,N_4889);
nor UO_281 (O_281,N_4683,N_4741);
nand UO_282 (O_282,N_4767,N_4777);
and UO_283 (O_283,N_4870,N_4984);
or UO_284 (O_284,N_4899,N_4559);
nor UO_285 (O_285,N_4769,N_4602);
nor UO_286 (O_286,N_4976,N_4878);
nor UO_287 (O_287,N_4902,N_4766);
or UO_288 (O_288,N_4526,N_4907);
nor UO_289 (O_289,N_4799,N_4852);
or UO_290 (O_290,N_4670,N_4736);
and UO_291 (O_291,N_4976,N_4782);
nor UO_292 (O_292,N_4954,N_4745);
nor UO_293 (O_293,N_4604,N_4739);
or UO_294 (O_294,N_4548,N_4558);
or UO_295 (O_295,N_4790,N_4925);
and UO_296 (O_296,N_4590,N_4589);
and UO_297 (O_297,N_4594,N_4621);
nor UO_298 (O_298,N_4559,N_4773);
nor UO_299 (O_299,N_4736,N_4946);
or UO_300 (O_300,N_4515,N_4693);
nor UO_301 (O_301,N_4655,N_4667);
and UO_302 (O_302,N_4870,N_4985);
nor UO_303 (O_303,N_4993,N_4611);
nand UO_304 (O_304,N_4892,N_4894);
xnor UO_305 (O_305,N_4625,N_4720);
or UO_306 (O_306,N_4956,N_4708);
or UO_307 (O_307,N_4549,N_4539);
and UO_308 (O_308,N_4504,N_4696);
nor UO_309 (O_309,N_4705,N_4948);
nand UO_310 (O_310,N_4958,N_4815);
and UO_311 (O_311,N_4886,N_4707);
nand UO_312 (O_312,N_4847,N_4973);
nor UO_313 (O_313,N_4887,N_4544);
nor UO_314 (O_314,N_4796,N_4931);
and UO_315 (O_315,N_4573,N_4975);
and UO_316 (O_316,N_4508,N_4564);
nor UO_317 (O_317,N_4638,N_4990);
or UO_318 (O_318,N_4749,N_4755);
or UO_319 (O_319,N_4866,N_4535);
nor UO_320 (O_320,N_4545,N_4743);
nand UO_321 (O_321,N_4833,N_4790);
and UO_322 (O_322,N_4559,N_4934);
nand UO_323 (O_323,N_4505,N_4865);
and UO_324 (O_324,N_4550,N_4619);
and UO_325 (O_325,N_4580,N_4703);
nand UO_326 (O_326,N_4569,N_4716);
or UO_327 (O_327,N_4865,N_4533);
and UO_328 (O_328,N_4759,N_4621);
or UO_329 (O_329,N_4884,N_4556);
and UO_330 (O_330,N_4887,N_4633);
or UO_331 (O_331,N_4979,N_4706);
and UO_332 (O_332,N_4689,N_4630);
nor UO_333 (O_333,N_4915,N_4632);
xor UO_334 (O_334,N_4697,N_4845);
or UO_335 (O_335,N_4654,N_4539);
nand UO_336 (O_336,N_4648,N_4751);
nor UO_337 (O_337,N_4929,N_4785);
nor UO_338 (O_338,N_4992,N_4813);
nand UO_339 (O_339,N_4660,N_4978);
nand UO_340 (O_340,N_4641,N_4569);
nor UO_341 (O_341,N_4767,N_4577);
nor UO_342 (O_342,N_4647,N_4588);
nand UO_343 (O_343,N_4953,N_4536);
and UO_344 (O_344,N_4810,N_4809);
nand UO_345 (O_345,N_4562,N_4812);
and UO_346 (O_346,N_4689,N_4943);
or UO_347 (O_347,N_4562,N_4988);
nand UO_348 (O_348,N_4879,N_4933);
nor UO_349 (O_349,N_4612,N_4709);
and UO_350 (O_350,N_4887,N_4691);
and UO_351 (O_351,N_4827,N_4936);
and UO_352 (O_352,N_4746,N_4600);
or UO_353 (O_353,N_4812,N_4501);
nor UO_354 (O_354,N_4859,N_4929);
nor UO_355 (O_355,N_4686,N_4952);
and UO_356 (O_356,N_4563,N_4694);
nor UO_357 (O_357,N_4542,N_4861);
nor UO_358 (O_358,N_4501,N_4641);
or UO_359 (O_359,N_4576,N_4775);
nand UO_360 (O_360,N_4563,N_4849);
or UO_361 (O_361,N_4900,N_4972);
and UO_362 (O_362,N_4783,N_4969);
nor UO_363 (O_363,N_4906,N_4758);
nand UO_364 (O_364,N_4936,N_4987);
and UO_365 (O_365,N_4708,N_4842);
nor UO_366 (O_366,N_4967,N_4547);
nand UO_367 (O_367,N_4627,N_4606);
and UO_368 (O_368,N_4821,N_4861);
nand UO_369 (O_369,N_4732,N_4996);
or UO_370 (O_370,N_4622,N_4796);
or UO_371 (O_371,N_4983,N_4680);
nand UO_372 (O_372,N_4543,N_4962);
nand UO_373 (O_373,N_4869,N_4616);
nand UO_374 (O_374,N_4520,N_4716);
or UO_375 (O_375,N_4558,N_4505);
or UO_376 (O_376,N_4651,N_4966);
nor UO_377 (O_377,N_4763,N_4621);
and UO_378 (O_378,N_4574,N_4857);
or UO_379 (O_379,N_4870,N_4913);
nor UO_380 (O_380,N_4576,N_4959);
or UO_381 (O_381,N_4952,N_4707);
nand UO_382 (O_382,N_4568,N_4554);
and UO_383 (O_383,N_4947,N_4936);
and UO_384 (O_384,N_4554,N_4939);
or UO_385 (O_385,N_4812,N_4942);
or UO_386 (O_386,N_4998,N_4784);
or UO_387 (O_387,N_4626,N_4562);
nand UO_388 (O_388,N_4869,N_4716);
or UO_389 (O_389,N_4807,N_4835);
and UO_390 (O_390,N_4544,N_4667);
and UO_391 (O_391,N_4938,N_4853);
or UO_392 (O_392,N_4616,N_4527);
and UO_393 (O_393,N_4524,N_4742);
and UO_394 (O_394,N_4565,N_4927);
or UO_395 (O_395,N_4888,N_4902);
nand UO_396 (O_396,N_4790,N_4671);
and UO_397 (O_397,N_4522,N_4559);
or UO_398 (O_398,N_4627,N_4933);
and UO_399 (O_399,N_4805,N_4673);
nor UO_400 (O_400,N_4553,N_4962);
nand UO_401 (O_401,N_4943,N_4819);
nand UO_402 (O_402,N_4544,N_4532);
nand UO_403 (O_403,N_4563,N_4940);
or UO_404 (O_404,N_4650,N_4555);
or UO_405 (O_405,N_4512,N_4751);
nor UO_406 (O_406,N_4508,N_4524);
nor UO_407 (O_407,N_4998,N_4604);
and UO_408 (O_408,N_4780,N_4564);
or UO_409 (O_409,N_4556,N_4614);
nor UO_410 (O_410,N_4593,N_4979);
nand UO_411 (O_411,N_4929,N_4654);
and UO_412 (O_412,N_4546,N_4982);
or UO_413 (O_413,N_4539,N_4930);
or UO_414 (O_414,N_4610,N_4560);
or UO_415 (O_415,N_4715,N_4905);
or UO_416 (O_416,N_4556,N_4792);
or UO_417 (O_417,N_4856,N_4522);
and UO_418 (O_418,N_4840,N_4814);
nand UO_419 (O_419,N_4574,N_4519);
or UO_420 (O_420,N_4924,N_4678);
and UO_421 (O_421,N_4504,N_4922);
and UO_422 (O_422,N_4817,N_4626);
nor UO_423 (O_423,N_4987,N_4734);
nand UO_424 (O_424,N_4606,N_4833);
and UO_425 (O_425,N_4562,N_4719);
and UO_426 (O_426,N_4795,N_4511);
nor UO_427 (O_427,N_4695,N_4519);
nand UO_428 (O_428,N_4986,N_4673);
or UO_429 (O_429,N_4727,N_4805);
nand UO_430 (O_430,N_4665,N_4595);
and UO_431 (O_431,N_4711,N_4814);
nand UO_432 (O_432,N_4950,N_4727);
or UO_433 (O_433,N_4976,N_4542);
and UO_434 (O_434,N_4917,N_4526);
or UO_435 (O_435,N_4680,N_4899);
or UO_436 (O_436,N_4979,N_4832);
and UO_437 (O_437,N_4915,N_4698);
or UO_438 (O_438,N_4722,N_4688);
or UO_439 (O_439,N_4819,N_4907);
and UO_440 (O_440,N_4584,N_4861);
and UO_441 (O_441,N_4548,N_4557);
nand UO_442 (O_442,N_4851,N_4776);
and UO_443 (O_443,N_4774,N_4653);
or UO_444 (O_444,N_4985,N_4883);
or UO_445 (O_445,N_4838,N_4601);
and UO_446 (O_446,N_4519,N_4674);
nand UO_447 (O_447,N_4911,N_4709);
nand UO_448 (O_448,N_4909,N_4945);
nand UO_449 (O_449,N_4744,N_4980);
nand UO_450 (O_450,N_4836,N_4667);
or UO_451 (O_451,N_4790,N_4586);
nor UO_452 (O_452,N_4952,N_4818);
or UO_453 (O_453,N_4657,N_4778);
and UO_454 (O_454,N_4597,N_4862);
and UO_455 (O_455,N_4713,N_4790);
nand UO_456 (O_456,N_4516,N_4856);
and UO_457 (O_457,N_4740,N_4647);
or UO_458 (O_458,N_4558,N_4514);
nor UO_459 (O_459,N_4505,N_4832);
nand UO_460 (O_460,N_4547,N_4697);
nand UO_461 (O_461,N_4788,N_4706);
and UO_462 (O_462,N_4953,N_4873);
or UO_463 (O_463,N_4503,N_4735);
nor UO_464 (O_464,N_4756,N_4829);
nand UO_465 (O_465,N_4727,N_4707);
or UO_466 (O_466,N_4773,N_4686);
nor UO_467 (O_467,N_4776,N_4917);
nand UO_468 (O_468,N_4801,N_4558);
nor UO_469 (O_469,N_4816,N_4809);
xor UO_470 (O_470,N_4987,N_4510);
and UO_471 (O_471,N_4507,N_4712);
nand UO_472 (O_472,N_4646,N_4628);
nor UO_473 (O_473,N_4956,N_4793);
and UO_474 (O_474,N_4505,N_4671);
nor UO_475 (O_475,N_4941,N_4814);
and UO_476 (O_476,N_4588,N_4767);
or UO_477 (O_477,N_4668,N_4919);
or UO_478 (O_478,N_4705,N_4895);
nand UO_479 (O_479,N_4520,N_4576);
or UO_480 (O_480,N_4908,N_4646);
or UO_481 (O_481,N_4735,N_4859);
or UO_482 (O_482,N_4855,N_4986);
or UO_483 (O_483,N_4768,N_4816);
nand UO_484 (O_484,N_4868,N_4765);
or UO_485 (O_485,N_4688,N_4691);
or UO_486 (O_486,N_4835,N_4624);
or UO_487 (O_487,N_4542,N_4652);
nor UO_488 (O_488,N_4932,N_4974);
and UO_489 (O_489,N_4547,N_4828);
nand UO_490 (O_490,N_4992,N_4987);
nand UO_491 (O_491,N_4569,N_4791);
and UO_492 (O_492,N_4772,N_4601);
nand UO_493 (O_493,N_4788,N_4694);
nand UO_494 (O_494,N_4840,N_4655);
xnor UO_495 (O_495,N_4554,N_4629);
nor UO_496 (O_496,N_4724,N_4701);
nand UO_497 (O_497,N_4821,N_4765);
nand UO_498 (O_498,N_4907,N_4543);
and UO_499 (O_499,N_4804,N_4903);
nor UO_500 (O_500,N_4914,N_4643);
nand UO_501 (O_501,N_4511,N_4755);
and UO_502 (O_502,N_4511,N_4750);
or UO_503 (O_503,N_4513,N_4699);
or UO_504 (O_504,N_4763,N_4980);
nor UO_505 (O_505,N_4784,N_4647);
or UO_506 (O_506,N_4543,N_4855);
and UO_507 (O_507,N_4847,N_4611);
nor UO_508 (O_508,N_4534,N_4552);
and UO_509 (O_509,N_4998,N_4698);
and UO_510 (O_510,N_4538,N_4671);
or UO_511 (O_511,N_4954,N_4525);
nor UO_512 (O_512,N_4630,N_4753);
and UO_513 (O_513,N_4779,N_4763);
nor UO_514 (O_514,N_4726,N_4753);
nor UO_515 (O_515,N_4669,N_4952);
nor UO_516 (O_516,N_4937,N_4835);
and UO_517 (O_517,N_4738,N_4505);
xor UO_518 (O_518,N_4760,N_4696);
nor UO_519 (O_519,N_4707,N_4758);
nor UO_520 (O_520,N_4579,N_4539);
or UO_521 (O_521,N_4802,N_4850);
nand UO_522 (O_522,N_4926,N_4969);
or UO_523 (O_523,N_4921,N_4807);
or UO_524 (O_524,N_4700,N_4994);
nor UO_525 (O_525,N_4860,N_4991);
and UO_526 (O_526,N_4649,N_4821);
nor UO_527 (O_527,N_4697,N_4665);
nand UO_528 (O_528,N_4611,N_4516);
nand UO_529 (O_529,N_4710,N_4702);
nor UO_530 (O_530,N_4849,N_4888);
and UO_531 (O_531,N_4729,N_4998);
nor UO_532 (O_532,N_4597,N_4724);
nor UO_533 (O_533,N_4781,N_4922);
nor UO_534 (O_534,N_4527,N_4999);
and UO_535 (O_535,N_4642,N_4510);
xor UO_536 (O_536,N_4568,N_4680);
and UO_537 (O_537,N_4729,N_4823);
and UO_538 (O_538,N_4884,N_4606);
nor UO_539 (O_539,N_4618,N_4916);
or UO_540 (O_540,N_4873,N_4708);
and UO_541 (O_541,N_4879,N_4540);
nand UO_542 (O_542,N_4901,N_4726);
nand UO_543 (O_543,N_4790,N_4928);
nand UO_544 (O_544,N_4539,N_4517);
and UO_545 (O_545,N_4984,N_4843);
and UO_546 (O_546,N_4969,N_4875);
and UO_547 (O_547,N_4758,N_4774);
or UO_548 (O_548,N_4758,N_4649);
nor UO_549 (O_549,N_4974,N_4534);
or UO_550 (O_550,N_4938,N_4937);
nand UO_551 (O_551,N_4918,N_4657);
nand UO_552 (O_552,N_4631,N_4950);
and UO_553 (O_553,N_4720,N_4763);
nand UO_554 (O_554,N_4885,N_4956);
nor UO_555 (O_555,N_4662,N_4823);
xor UO_556 (O_556,N_4977,N_4917);
nor UO_557 (O_557,N_4636,N_4836);
and UO_558 (O_558,N_4923,N_4944);
or UO_559 (O_559,N_4544,N_4791);
nand UO_560 (O_560,N_4543,N_4674);
nor UO_561 (O_561,N_4578,N_4739);
and UO_562 (O_562,N_4832,N_4882);
nand UO_563 (O_563,N_4746,N_4867);
nand UO_564 (O_564,N_4589,N_4743);
nor UO_565 (O_565,N_4773,N_4849);
or UO_566 (O_566,N_4911,N_4792);
nor UO_567 (O_567,N_4714,N_4517);
nor UO_568 (O_568,N_4883,N_4563);
nand UO_569 (O_569,N_4992,N_4751);
and UO_570 (O_570,N_4561,N_4990);
or UO_571 (O_571,N_4706,N_4696);
and UO_572 (O_572,N_4803,N_4591);
nor UO_573 (O_573,N_4903,N_4515);
and UO_574 (O_574,N_4763,N_4885);
and UO_575 (O_575,N_4902,N_4986);
nor UO_576 (O_576,N_4920,N_4816);
or UO_577 (O_577,N_4858,N_4795);
and UO_578 (O_578,N_4650,N_4926);
nand UO_579 (O_579,N_4812,N_4838);
or UO_580 (O_580,N_4628,N_4741);
and UO_581 (O_581,N_4555,N_4942);
nor UO_582 (O_582,N_4664,N_4657);
and UO_583 (O_583,N_4797,N_4827);
or UO_584 (O_584,N_4872,N_4922);
nor UO_585 (O_585,N_4817,N_4590);
nor UO_586 (O_586,N_4840,N_4608);
or UO_587 (O_587,N_4637,N_4820);
nor UO_588 (O_588,N_4776,N_4548);
nor UO_589 (O_589,N_4927,N_4523);
nor UO_590 (O_590,N_4752,N_4600);
nor UO_591 (O_591,N_4968,N_4929);
nand UO_592 (O_592,N_4928,N_4806);
or UO_593 (O_593,N_4881,N_4909);
nor UO_594 (O_594,N_4738,N_4590);
nor UO_595 (O_595,N_4943,N_4663);
or UO_596 (O_596,N_4517,N_4755);
nand UO_597 (O_597,N_4877,N_4989);
nand UO_598 (O_598,N_4911,N_4658);
nor UO_599 (O_599,N_4851,N_4615);
nor UO_600 (O_600,N_4555,N_4948);
nand UO_601 (O_601,N_4874,N_4663);
nor UO_602 (O_602,N_4694,N_4973);
and UO_603 (O_603,N_4652,N_4612);
or UO_604 (O_604,N_4689,N_4939);
nand UO_605 (O_605,N_4738,N_4809);
nand UO_606 (O_606,N_4813,N_4891);
nor UO_607 (O_607,N_4727,N_4965);
nand UO_608 (O_608,N_4925,N_4906);
or UO_609 (O_609,N_4676,N_4982);
or UO_610 (O_610,N_4878,N_4905);
or UO_611 (O_611,N_4987,N_4914);
or UO_612 (O_612,N_4889,N_4751);
xor UO_613 (O_613,N_4875,N_4530);
and UO_614 (O_614,N_4671,N_4808);
nor UO_615 (O_615,N_4797,N_4724);
nand UO_616 (O_616,N_4992,N_4684);
nor UO_617 (O_617,N_4705,N_4529);
and UO_618 (O_618,N_4563,N_4585);
nand UO_619 (O_619,N_4769,N_4606);
or UO_620 (O_620,N_4763,N_4892);
and UO_621 (O_621,N_4527,N_4861);
or UO_622 (O_622,N_4551,N_4573);
nor UO_623 (O_623,N_4653,N_4834);
nor UO_624 (O_624,N_4984,N_4747);
and UO_625 (O_625,N_4788,N_4828);
or UO_626 (O_626,N_4984,N_4911);
or UO_627 (O_627,N_4578,N_4520);
nand UO_628 (O_628,N_4697,N_4814);
nand UO_629 (O_629,N_4599,N_4896);
nand UO_630 (O_630,N_4985,N_4614);
or UO_631 (O_631,N_4726,N_4792);
nand UO_632 (O_632,N_4864,N_4697);
nand UO_633 (O_633,N_4686,N_4664);
nand UO_634 (O_634,N_4679,N_4665);
and UO_635 (O_635,N_4696,N_4521);
nand UO_636 (O_636,N_4965,N_4742);
or UO_637 (O_637,N_4880,N_4529);
and UO_638 (O_638,N_4891,N_4543);
nand UO_639 (O_639,N_4502,N_4744);
and UO_640 (O_640,N_4677,N_4693);
nand UO_641 (O_641,N_4914,N_4851);
or UO_642 (O_642,N_4549,N_4813);
or UO_643 (O_643,N_4861,N_4628);
and UO_644 (O_644,N_4757,N_4530);
or UO_645 (O_645,N_4931,N_4930);
nand UO_646 (O_646,N_4715,N_4674);
or UO_647 (O_647,N_4506,N_4863);
nor UO_648 (O_648,N_4774,N_4832);
or UO_649 (O_649,N_4749,N_4604);
nand UO_650 (O_650,N_4779,N_4785);
nand UO_651 (O_651,N_4591,N_4967);
and UO_652 (O_652,N_4748,N_4841);
nor UO_653 (O_653,N_4652,N_4706);
nor UO_654 (O_654,N_4768,N_4720);
and UO_655 (O_655,N_4949,N_4555);
nor UO_656 (O_656,N_4566,N_4964);
nand UO_657 (O_657,N_4509,N_4538);
nand UO_658 (O_658,N_4767,N_4776);
and UO_659 (O_659,N_4984,N_4695);
nand UO_660 (O_660,N_4688,N_4655);
or UO_661 (O_661,N_4860,N_4543);
nand UO_662 (O_662,N_4773,N_4926);
or UO_663 (O_663,N_4787,N_4542);
nor UO_664 (O_664,N_4833,N_4653);
nand UO_665 (O_665,N_4797,N_4955);
and UO_666 (O_666,N_4585,N_4912);
or UO_667 (O_667,N_4765,N_4694);
and UO_668 (O_668,N_4655,N_4943);
nor UO_669 (O_669,N_4644,N_4796);
nand UO_670 (O_670,N_4765,N_4565);
and UO_671 (O_671,N_4768,N_4642);
nor UO_672 (O_672,N_4837,N_4743);
and UO_673 (O_673,N_4767,N_4660);
nor UO_674 (O_674,N_4718,N_4526);
nand UO_675 (O_675,N_4746,N_4775);
and UO_676 (O_676,N_4676,N_4755);
and UO_677 (O_677,N_4786,N_4679);
nor UO_678 (O_678,N_4945,N_4688);
nor UO_679 (O_679,N_4990,N_4819);
nand UO_680 (O_680,N_4844,N_4546);
nor UO_681 (O_681,N_4660,N_4512);
or UO_682 (O_682,N_4705,N_4593);
and UO_683 (O_683,N_4536,N_4635);
nor UO_684 (O_684,N_4513,N_4598);
or UO_685 (O_685,N_4905,N_4800);
nor UO_686 (O_686,N_4826,N_4925);
and UO_687 (O_687,N_4598,N_4734);
and UO_688 (O_688,N_4788,N_4984);
nand UO_689 (O_689,N_4688,N_4868);
nand UO_690 (O_690,N_4823,N_4608);
or UO_691 (O_691,N_4880,N_4808);
nand UO_692 (O_692,N_4813,N_4973);
nor UO_693 (O_693,N_4543,N_4799);
or UO_694 (O_694,N_4802,N_4981);
or UO_695 (O_695,N_4849,N_4774);
and UO_696 (O_696,N_4976,N_4599);
and UO_697 (O_697,N_4737,N_4885);
nor UO_698 (O_698,N_4543,N_4512);
or UO_699 (O_699,N_4513,N_4962);
nor UO_700 (O_700,N_4879,N_4965);
or UO_701 (O_701,N_4756,N_4692);
and UO_702 (O_702,N_4837,N_4741);
nand UO_703 (O_703,N_4982,N_4603);
nand UO_704 (O_704,N_4651,N_4733);
nor UO_705 (O_705,N_4592,N_4737);
nor UO_706 (O_706,N_4726,N_4741);
nor UO_707 (O_707,N_4992,N_4613);
nand UO_708 (O_708,N_4755,N_4741);
or UO_709 (O_709,N_4835,N_4656);
nor UO_710 (O_710,N_4730,N_4615);
nor UO_711 (O_711,N_4921,N_4557);
nor UO_712 (O_712,N_4829,N_4892);
and UO_713 (O_713,N_4682,N_4673);
nand UO_714 (O_714,N_4749,N_4719);
and UO_715 (O_715,N_4878,N_4924);
or UO_716 (O_716,N_4802,N_4846);
and UO_717 (O_717,N_4550,N_4908);
nand UO_718 (O_718,N_4912,N_4689);
or UO_719 (O_719,N_4831,N_4746);
nand UO_720 (O_720,N_4875,N_4536);
nor UO_721 (O_721,N_4662,N_4778);
and UO_722 (O_722,N_4751,N_4919);
nor UO_723 (O_723,N_4880,N_4619);
nor UO_724 (O_724,N_4611,N_4937);
or UO_725 (O_725,N_4604,N_4926);
and UO_726 (O_726,N_4908,N_4911);
nand UO_727 (O_727,N_4962,N_4653);
nand UO_728 (O_728,N_4822,N_4935);
nand UO_729 (O_729,N_4840,N_4642);
or UO_730 (O_730,N_4983,N_4726);
nor UO_731 (O_731,N_4982,N_4720);
nand UO_732 (O_732,N_4944,N_4513);
and UO_733 (O_733,N_4739,N_4500);
nor UO_734 (O_734,N_4938,N_4890);
nor UO_735 (O_735,N_4904,N_4897);
nor UO_736 (O_736,N_4626,N_4973);
nand UO_737 (O_737,N_4920,N_4866);
and UO_738 (O_738,N_4645,N_4972);
or UO_739 (O_739,N_4522,N_4738);
nand UO_740 (O_740,N_4688,N_4550);
or UO_741 (O_741,N_4604,N_4876);
nor UO_742 (O_742,N_4695,N_4838);
or UO_743 (O_743,N_4858,N_4981);
and UO_744 (O_744,N_4592,N_4962);
or UO_745 (O_745,N_4916,N_4673);
nor UO_746 (O_746,N_4686,N_4527);
nor UO_747 (O_747,N_4863,N_4792);
or UO_748 (O_748,N_4518,N_4617);
nor UO_749 (O_749,N_4555,N_4652);
or UO_750 (O_750,N_4891,N_4907);
or UO_751 (O_751,N_4710,N_4787);
nor UO_752 (O_752,N_4912,N_4891);
or UO_753 (O_753,N_4776,N_4787);
or UO_754 (O_754,N_4553,N_4744);
nor UO_755 (O_755,N_4982,N_4558);
nand UO_756 (O_756,N_4908,N_4983);
and UO_757 (O_757,N_4576,N_4584);
nor UO_758 (O_758,N_4514,N_4828);
nand UO_759 (O_759,N_4574,N_4514);
xor UO_760 (O_760,N_4642,N_4913);
nor UO_761 (O_761,N_4509,N_4665);
and UO_762 (O_762,N_4548,N_4705);
or UO_763 (O_763,N_4654,N_4787);
or UO_764 (O_764,N_4893,N_4735);
and UO_765 (O_765,N_4889,N_4912);
and UO_766 (O_766,N_4655,N_4506);
xnor UO_767 (O_767,N_4922,N_4790);
or UO_768 (O_768,N_4711,N_4631);
nand UO_769 (O_769,N_4854,N_4742);
nor UO_770 (O_770,N_4915,N_4726);
and UO_771 (O_771,N_4597,N_4638);
nor UO_772 (O_772,N_4559,N_4688);
nor UO_773 (O_773,N_4912,N_4666);
and UO_774 (O_774,N_4511,N_4834);
nand UO_775 (O_775,N_4505,N_4601);
nand UO_776 (O_776,N_4568,N_4828);
nand UO_777 (O_777,N_4793,N_4516);
nand UO_778 (O_778,N_4607,N_4506);
nand UO_779 (O_779,N_4922,N_4857);
nand UO_780 (O_780,N_4631,N_4754);
and UO_781 (O_781,N_4784,N_4873);
nor UO_782 (O_782,N_4529,N_4890);
nor UO_783 (O_783,N_4526,N_4602);
or UO_784 (O_784,N_4730,N_4678);
and UO_785 (O_785,N_4883,N_4671);
nand UO_786 (O_786,N_4515,N_4675);
or UO_787 (O_787,N_4731,N_4693);
and UO_788 (O_788,N_4882,N_4522);
nor UO_789 (O_789,N_4512,N_4559);
and UO_790 (O_790,N_4871,N_4798);
nand UO_791 (O_791,N_4674,N_4852);
or UO_792 (O_792,N_4661,N_4694);
nand UO_793 (O_793,N_4995,N_4738);
nor UO_794 (O_794,N_4806,N_4809);
and UO_795 (O_795,N_4703,N_4756);
and UO_796 (O_796,N_4584,N_4980);
nor UO_797 (O_797,N_4931,N_4747);
and UO_798 (O_798,N_4597,N_4536);
nor UO_799 (O_799,N_4723,N_4951);
nor UO_800 (O_800,N_4784,N_4505);
or UO_801 (O_801,N_4788,N_4550);
or UO_802 (O_802,N_4531,N_4928);
nand UO_803 (O_803,N_4708,N_4530);
and UO_804 (O_804,N_4549,N_4828);
and UO_805 (O_805,N_4590,N_4673);
or UO_806 (O_806,N_4542,N_4987);
nand UO_807 (O_807,N_4748,N_4551);
and UO_808 (O_808,N_4689,N_4514);
or UO_809 (O_809,N_4790,N_4656);
or UO_810 (O_810,N_4604,N_4727);
and UO_811 (O_811,N_4996,N_4688);
nor UO_812 (O_812,N_4515,N_4970);
and UO_813 (O_813,N_4543,N_4568);
nor UO_814 (O_814,N_4659,N_4821);
nor UO_815 (O_815,N_4808,N_4613);
nor UO_816 (O_816,N_4954,N_4502);
nand UO_817 (O_817,N_4805,N_4680);
and UO_818 (O_818,N_4509,N_4980);
or UO_819 (O_819,N_4841,N_4807);
nand UO_820 (O_820,N_4562,N_4769);
and UO_821 (O_821,N_4752,N_4754);
and UO_822 (O_822,N_4670,N_4554);
nand UO_823 (O_823,N_4671,N_4675);
xnor UO_824 (O_824,N_4901,N_4769);
and UO_825 (O_825,N_4735,N_4943);
and UO_826 (O_826,N_4903,N_4913);
nor UO_827 (O_827,N_4733,N_4950);
and UO_828 (O_828,N_4876,N_4829);
nor UO_829 (O_829,N_4915,N_4680);
nand UO_830 (O_830,N_4748,N_4727);
nor UO_831 (O_831,N_4650,N_4818);
nand UO_832 (O_832,N_4801,N_4968);
and UO_833 (O_833,N_4514,N_4751);
or UO_834 (O_834,N_4934,N_4638);
and UO_835 (O_835,N_4641,N_4571);
or UO_836 (O_836,N_4702,N_4982);
nor UO_837 (O_837,N_4598,N_4500);
and UO_838 (O_838,N_4973,N_4866);
and UO_839 (O_839,N_4503,N_4846);
or UO_840 (O_840,N_4825,N_4656);
or UO_841 (O_841,N_4509,N_4882);
and UO_842 (O_842,N_4902,N_4545);
nor UO_843 (O_843,N_4830,N_4809);
and UO_844 (O_844,N_4966,N_4616);
nand UO_845 (O_845,N_4855,N_4812);
or UO_846 (O_846,N_4786,N_4732);
and UO_847 (O_847,N_4792,N_4980);
and UO_848 (O_848,N_4579,N_4784);
or UO_849 (O_849,N_4507,N_4573);
nor UO_850 (O_850,N_4645,N_4600);
nand UO_851 (O_851,N_4612,N_4679);
or UO_852 (O_852,N_4819,N_4739);
and UO_853 (O_853,N_4734,N_4888);
nand UO_854 (O_854,N_4645,N_4815);
nand UO_855 (O_855,N_4979,N_4957);
nor UO_856 (O_856,N_4551,N_4806);
nor UO_857 (O_857,N_4648,N_4777);
xor UO_858 (O_858,N_4639,N_4611);
or UO_859 (O_859,N_4722,N_4945);
or UO_860 (O_860,N_4971,N_4944);
nor UO_861 (O_861,N_4811,N_4705);
or UO_862 (O_862,N_4626,N_4628);
or UO_863 (O_863,N_4710,N_4514);
nor UO_864 (O_864,N_4707,N_4653);
and UO_865 (O_865,N_4914,N_4828);
nor UO_866 (O_866,N_4895,N_4767);
nor UO_867 (O_867,N_4790,N_4530);
and UO_868 (O_868,N_4864,N_4853);
nor UO_869 (O_869,N_4768,N_4740);
and UO_870 (O_870,N_4693,N_4884);
and UO_871 (O_871,N_4871,N_4520);
and UO_872 (O_872,N_4561,N_4846);
nor UO_873 (O_873,N_4699,N_4747);
or UO_874 (O_874,N_4988,N_4699);
nor UO_875 (O_875,N_4608,N_4999);
or UO_876 (O_876,N_4853,N_4508);
and UO_877 (O_877,N_4567,N_4960);
nor UO_878 (O_878,N_4889,N_4739);
and UO_879 (O_879,N_4518,N_4686);
or UO_880 (O_880,N_4757,N_4918);
and UO_881 (O_881,N_4763,N_4773);
nor UO_882 (O_882,N_4959,N_4789);
nor UO_883 (O_883,N_4815,N_4589);
nand UO_884 (O_884,N_4795,N_4514);
and UO_885 (O_885,N_4977,N_4939);
and UO_886 (O_886,N_4860,N_4514);
nand UO_887 (O_887,N_4802,N_4852);
and UO_888 (O_888,N_4636,N_4974);
nor UO_889 (O_889,N_4902,N_4885);
nand UO_890 (O_890,N_4508,N_4655);
nand UO_891 (O_891,N_4979,N_4881);
and UO_892 (O_892,N_4717,N_4583);
nor UO_893 (O_893,N_4721,N_4622);
or UO_894 (O_894,N_4758,N_4950);
or UO_895 (O_895,N_4935,N_4869);
or UO_896 (O_896,N_4598,N_4871);
and UO_897 (O_897,N_4954,N_4619);
or UO_898 (O_898,N_4989,N_4796);
xor UO_899 (O_899,N_4558,N_4715);
xor UO_900 (O_900,N_4944,N_4809);
or UO_901 (O_901,N_4749,N_4503);
nor UO_902 (O_902,N_4945,N_4860);
and UO_903 (O_903,N_4927,N_4640);
and UO_904 (O_904,N_4637,N_4938);
nand UO_905 (O_905,N_4594,N_4743);
nor UO_906 (O_906,N_4528,N_4505);
nor UO_907 (O_907,N_4804,N_4814);
or UO_908 (O_908,N_4843,N_4827);
nand UO_909 (O_909,N_4904,N_4801);
and UO_910 (O_910,N_4744,N_4936);
and UO_911 (O_911,N_4603,N_4610);
nor UO_912 (O_912,N_4691,N_4630);
nand UO_913 (O_913,N_4974,N_4632);
and UO_914 (O_914,N_4511,N_4914);
nor UO_915 (O_915,N_4523,N_4969);
nand UO_916 (O_916,N_4612,N_4799);
and UO_917 (O_917,N_4869,N_4504);
nor UO_918 (O_918,N_4653,N_4571);
nand UO_919 (O_919,N_4857,N_4984);
nor UO_920 (O_920,N_4976,N_4834);
and UO_921 (O_921,N_4804,N_4629);
and UO_922 (O_922,N_4554,N_4781);
nand UO_923 (O_923,N_4691,N_4827);
nor UO_924 (O_924,N_4730,N_4719);
or UO_925 (O_925,N_4721,N_4755);
or UO_926 (O_926,N_4507,N_4971);
nor UO_927 (O_927,N_4539,N_4561);
nor UO_928 (O_928,N_4926,N_4627);
or UO_929 (O_929,N_4685,N_4706);
and UO_930 (O_930,N_4555,N_4616);
nand UO_931 (O_931,N_4814,N_4956);
and UO_932 (O_932,N_4662,N_4668);
and UO_933 (O_933,N_4598,N_4603);
nand UO_934 (O_934,N_4789,N_4765);
and UO_935 (O_935,N_4936,N_4933);
nand UO_936 (O_936,N_4793,N_4765);
or UO_937 (O_937,N_4663,N_4842);
nor UO_938 (O_938,N_4975,N_4530);
nor UO_939 (O_939,N_4756,N_4852);
nand UO_940 (O_940,N_4689,N_4524);
nand UO_941 (O_941,N_4583,N_4600);
nor UO_942 (O_942,N_4665,N_4610);
nand UO_943 (O_943,N_4892,N_4601);
or UO_944 (O_944,N_4527,N_4747);
or UO_945 (O_945,N_4537,N_4887);
nand UO_946 (O_946,N_4556,N_4984);
and UO_947 (O_947,N_4515,N_4740);
nand UO_948 (O_948,N_4639,N_4641);
nand UO_949 (O_949,N_4761,N_4813);
and UO_950 (O_950,N_4669,N_4517);
and UO_951 (O_951,N_4656,N_4784);
and UO_952 (O_952,N_4954,N_4596);
or UO_953 (O_953,N_4802,N_4864);
nor UO_954 (O_954,N_4862,N_4885);
or UO_955 (O_955,N_4898,N_4778);
or UO_956 (O_956,N_4535,N_4664);
nor UO_957 (O_957,N_4553,N_4943);
xnor UO_958 (O_958,N_4789,N_4929);
nand UO_959 (O_959,N_4884,N_4921);
or UO_960 (O_960,N_4948,N_4799);
nor UO_961 (O_961,N_4776,N_4556);
or UO_962 (O_962,N_4538,N_4921);
or UO_963 (O_963,N_4517,N_4522);
and UO_964 (O_964,N_4545,N_4892);
nand UO_965 (O_965,N_4962,N_4600);
nor UO_966 (O_966,N_4656,N_4876);
or UO_967 (O_967,N_4673,N_4589);
and UO_968 (O_968,N_4680,N_4827);
and UO_969 (O_969,N_4748,N_4760);
nand UO_970 (O_970,N_4546,N_4594);
and UO_971 (O_971,N_4538,N_4791);
or UO_972 (O_972,N_4910,N_4574);
nor UO_973 (O_973,N_4706,N_4883);
nor UO_974 (O_974,N_4789,N_4643);
and UO_975 (O_975,N_4593,N_4867);
nand UO_976 (O_976,N_4782,N_4755);
and UO_977 (O_977,N_4620,N_4729);
nand UO_978 (O_978,N_4847,N_4607);
nand UO_979 (O_979,N_4971,N_4822);
nand UO_980 (O_980,N_4917,N_4763);
and UO_981 (O_981,N_4728,N_4588);
or UO_982 (O_982,N_4994,N_4907);
nor UO_983 (O_983,N_4738,N_4895);
nand UO_984 (O_984,N_4951,N_4977);
nor UO_985 (O_985,N_4538,N_4910);
nand UO_986 (O_986,N_4704,N_4524);
nor UO_987 (O_987,N_4631,N_4816);
nand UO_988 (O_988,N_4734,N_4576);
or UO_989 (O_989,N_4944,N_4759);
nor UO_990 (O_990,N_4813,N_4871);
nor UO_991 (O_991,N_4703,N_4953);
nor UO_992 (O_992,N_4693,N_4676);
nand UO_993 (O_993,N_4535,N_4549);
nand UO_994 (O_994,N_4972,N_4702);
and UO_995 (O_995,N_4915,N_4778);
nand UO_996 (O_996,N_4637,N_4539);
and UO_997 (O_997,N_4990,N_4737);
nor UO_998 (O_998,N_4832,N_4810);
nor UO_999 (O_999,N_4845,N_4711);
endmodule