module basic_1000_10000_1500_10_levels_1xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_18,In_750);
nor U1 (N_1,In_344,In_17);
and U2 (N_2,In_842,In_172);
nor U3 (N_3,In_761,In_918);
and U4 (N_4,In_351,In_223);
and U5 (N_5,In_101,In_495);
xor U6 (N_6,In_999,In_267);
nor U7 (N_7,In_785,In_292);
nand U8 (N_8,In_332,In_925);
nand U9 (N_9,In_961,In_437);
nand U10 (N_10,In_713,In_441);
or U11 (N_11,In_134,In_257);
or U12 (N_12,In_906,In_315);
and U13 (N_13,In_430,In_295);
or U14 (N_14,In_218,In_237);
nor U15 (N_15,In_775,In_791);
nand U16 (N_16,In_391,In_123);
nand U17 (N_17,In_362,In_623);
nor U18 (N_18,In_555,In_122);
nand U19 (N_19,In_929,In_600);
and U20 (N_20,In_135,In_656);
nor U21 (N_21,In_338,In_855);
and U22 (N_22,In_293,In_738);
nand U23 (N_23,In_119,In_660);
and U24 (N_24,In_987,In_685);
nand U25 (N_25,In_936,In_524);
and U26 (N_26,In_118,In_766);
or U27 (N_27,In_553,In_132);
or U28 (N_28,In_965,In_297);
nand U29 (N_29,In_424,In_498);
nand U30 (N_30,In_211,In_209);
and U31 (N_31,In_841,In_375);
nand U32 (N_32,In_889,In_802);
and U33 (N_33,In_635,In_300);
nor U34 (N_34,In_62,In_915);
or U35 (N_35,In_712,In_881);
and U36 (N_36,In_303,In_834);
nand U37 (N_37,In_336,In_125);
nand U38 (N_38,In_16,In_266);
or U39 (N_39,In_268,In_137);
and U40 (N_40,In_271,In_837);
and U41 (N_41,In_216,In_763);
and U42 (N_42,In_932,In_745);
nand U43 (N_43,In_171,In_217);
or U44 (N_44,In_556,In_769);
and U45 (N_45,In_507,In_420);
nand U46 (N_46,In_195,In_203);
nor U47 (N_47,In_423,In_730);
nand U48 (N_48,In_99,In_27);
nand U49 (N_49,In_24,In_898);
nor U50 (N_50,In_419,In_893);
nor U51 (N_51,In_408,In_457);
nor U52 (N_52,In_701,In_805);
nor U53 (N_53,In_497,In_835);
and U54 (N_54,In_803,In_819);
and U55 (N_55,In_201,In_272);
nand U56 (N_56,In_462,In_393);
nand U57 (N_57,In_684,In_341);
or U58 (N_58,In_175,In_156);
or U59 (N_59,In_288,In_523);
or U60 (N_60,In_709,In_824);
nand U61 (N_61,In_191,In_382);
or U62 (N_62,In_385,In_759);
nor U63 (N_63,In_215,In_251);
nor U64 (N_64,In_452,In_279);
and U65 (N_65,In_310,In_247);
and U66 (N_66,In_625,In_263);
nor U67 (N_67,In_659,In_696);
or U68 (N_68,In_586,In_964);
nand U69 (N_69,In_731,In_145);
and U70 (N_70,In_751,In_433);
or U71 (N_71,In_680,In_294);
nand U72 (N_72,In_595,In_96);
and U73 (N_73,In_417,In_314);
or U74 (N_74,In_230,In_867);
or U75 (N_75,In_374,In_945);
and U76 (N_76,In_29,In_492);
nor U77 (N_77,In_939,In_200);
and U78 (N_78,In_367,In_749);
nor U79 (N_79,In_951,In_818);
nor U80 (N_80,In_477,In_328);
or U81 (N_81,In_571,In_852);
and U82 (N_82,In_722,In_851);
nor U83 (N_83,In_346,In_493);
nor U84 (N_84,In_886,In_671);
nand U85 (N_85,In_853,In_827);
or U86 (N_86,In_113,In_318);
and U87 (N_87,In_102,In_645);
or U88 (N_88,In_980,In_776);
nand U89 (N_89,In_919,In_111);
nand U90 (N_90,In_883,In_800);
and U91 (N_91,In_690,In_655);
and U92 (N_92,In_90,In_952);
or U93 (N_93,In_468,In_427);
nand U94 (N_94,In_868,In_930);
nand U95 (N_95,In_583,In_161);
and U96 (N_96,In_325,In_164);
or U97 (N_97,In_447,In_782);
nor U98 (N_98,In_760,In_666);
or U99 (N_99,In_641,In_518);
or U100 (N_100,In_636,In_347);
or U101 (N_101,In_353,In_566);
nand U102 (N_102,In_202,In_993);
nor U103 (N_103,In_599,In_65);
xnor U104 (N_104,In_989,In_941);
or U105 (N_105,In_473,In_130);
or U106 (N_106,In_563,In_70);
or U107 (N_107,In_30,In_854);
nand U108 (N_108,In_753,In_21);
nand U109 (N_109,In_436,In_754);
and U110 (N_110,In_141,In_183);
and U111 (N_111,In_825,In_609);
nand U112 (N_112,In_770,In_466);
and U113 (N_113,In_320,In_312);
nor U114 (N_114,In_840,In_967);
nand U115 (N_115,In_923,In_801);
or U116 (N_116,In_98,In_364);
nand U117 (N_117,In_464,In_721);
nor U118 (N_118,In_662,In_545);
nor U119 (N_119,In_179,In_321);
nor U120 (N_120,In_559,In_110);
nand U121 (N_121,In_579,In_943);
and U122 (N_122,In_909,In_650);
nor U123 (N_123,In_587,In_574);
nor U124 (N_124,In_983,In_34);
or U125 (N_125,In_714,In_185);
nor U126 (N_126,In_259,In_632);
and U127 (N_127,In_284,In_529);
and U128 (N_128,In_527,In_736);
and U129 (N_129,In_658,In_42);
nand U130 (N_130,In_93,In_780);
and U131 (N_131,In_474,In_472);
or U132 (N_132,In_443,In_253);
or U133 (N_133,In_550,In_168);
and U134 (N_134,In_421,In_541);
nand U135 (N_135,In_705,In_2);
nand U136 (N_136,In_619,In_426);
nand U137 (N_137,In_544,In_789);
or U138 (N_138,In_585,In_904);
nor U139 (N_139,In_81,In_365);
nand U140 (N_140,In_675,In_928);
and U141 (N_141,In_549,In_764);
nor U142 (N_142,In_673,In_533);
nor U143 (N_143,In_304,In_148);
or U144 (N_144,In_407,In_72);
nor U145 (N_145,In_82,In_938);
or U146 (N_146,In_790,In_813);
or U147 (N_147,In_870,In_865);
nand U148 (N_148,In_615,In_740);
and U149 (N_149,In_604,In_12);
and U150 (N_150,In_395,In_914);
or U151 (N_151,In_167,In_565);
or U152 (N_152,In_719,In_717);
nor U153 (N_153,In_264,In_622);
or U154 (N_154,In_866,In_862);
nand U155 (N_155,In_494,In_843);
nor U156 (N_156,In_820,In_913);
and U157 (N_157,In_787,In_891);
or U158 (N_158,In_916,In_601);
and U159 (N_159,In_630,In_305);
and U160 (N_160,In_277,In_163);
nand U161 (N_161,In_100,In_535);
or U162 (N_162,In_948,In_301);
nand U163 (N_163,In_877,In_822);
nor U164 (N_164,In_439,In_143);
or U165 (N_165,In_706,In_910);
nor U166 (N_166,In_681,In_616);
and U167 (N_167,In_38,In_389);
nand U168 (N_168,In_536,In_84);
nand U169 (N_169,In_614,In_589);
and U170 (N_170,In_260,In_592);
or U171 (N_171,In_581,In_626);
nand U172 (N_172,In_124,In_155);
or U173 (N_173,In_323,In_922);
nor U174 (N_174,In_360,In_23);
nand U175 (N_175,In_463,In_235);
nand U176 (N_176,In_702,In_390);
and U177 (N_177,In_56,In_245);
or U178 (N_178,In_53,In_46);
and U179 (N_179,In_610,In_617);
and U180 (N_180,In_106,In_319);
nand U181 (N_181,In_104,In_977);
nand U182 (N_182,In_249,In_878);
nor U183 (N_183,In_514,In_548);
nor U184 (N_184,In_32,In_1);
nand U185 (N_185,In_368,In_376);
and U186 (N_186,In_401,In_349);
and U187 (N_187,In_434,In_611);
or U188 (N_188,In_151,In_220);
or U189 (N_189,In_520,In_783);
nand U190 (N_190,In_326,In_413);
and U191 (N_191,In_108,In_786);
or U192 (N_192,In_784,In_799);
and U193 (N_193,In_458,In_329);
nor U194 (N_194,In_665,In_949);
nand U195 (N_195,In_308,In_208);
and U196 (N_196,In_41,In_686);
and U197 (N_197,In_953,In_628);
nand U198 (N_198,In_265,In_63);
nor U199 (N_199,In_547,In_451);
nor U200 (N_200,In_757,In_744);
nor U201 (N_201,In_105,In_465);
and U202 (N_202,In_491,In_80);
and U203 (N_203,In_991,In_990);
nor U204 (N_204,In_89,In_154);
nor U205 (N_205,In_149,In_496);
nand U206 (N_206,In_821,In_222);
or U207 (N_207,In_695,In_501);
nand U208 (N_208,In_348,In_578);
or U209 (N_209,In_781,In_114);
nand U210 (N_210,In_572,In_661);
or U211 (N_211,In_152,In_399);
and U212 (N_212,In_109,In_689);
nand U213 (N_213,In_355,In_133);
nand U214 (N_214,In_598,In_704);
and U215 (N_215,In_359,In_159);
and U216 (N_216,In_697,In_902);
and U217 (N_217,In_988,In_729);
nor U218 (N_218,In_844,In_664);
and U219 (N_219,In_543,In_221);
nand U220 (N_220,In_997,In_752);
nand U221 (N_221,In_91,In_487);
or U222 (N_222,In_115,In_327);
and U223 (N_223,In_140,In_768);
or U224 (N_224,In_44,In_396);
and U225 (N_225,In_405,In_823);
nor U226 (N_226,In_937,In_334);
nand U227 (N_227,In_126,In_28);
or U228 (N_228,In_755,In_40);
nand U229 (N_229,In_299,In_252);
nor U230 (N_230,In_173,In_170);
nand U231 (N_231,In_933,In_994);
or U232 (N_232,In_682,In_181);
nor U233 (N_233,In_117,In_333);
nor U234 (N_234,In_817,In_54);
or U235 (N_235,In_828,In_788);
xor U236 (N_236,In_480,In_160);
or U237 (N_237,In_613,In_885);
nor U238 (N_238,In_189,In_76);
nand U239 (N_239,In_558,In_575);
or U240 (N_240,In_429,In_127);
or U241 (N_241,In_631,In_386);
nand U242 (N_242,In_475,In_739);
nand U243 (N_243,In_537,In_735);
nand U244 (N_244,In_43,In_370);
and U245 (N_245,In_187,In_435);
nand U246 (N_246,In_920,In_629);
and U247 (N_247,In_489,In_290);
and U248 (N_248,In_403,In_289);
or U249 (N_249,In_833,In_580);
nor U250 (N_250,In_459,In_311);
nor U251 (N_251,In_343,In_639);
or U252 (N_252,In_476,In_986);
nor U253 (N_253,In_49,In_234);
nor U254 (N_254,In_880,In_995);
and U255 (N_255,In_678,In_246);
nor U256 (N_256,In_551,In_792);
nor U257 (N_257,In_795,In_955);
nor U258 (N_258,In_888,In_37);
nor U259 (N_259,In_446,In_193);
nand U260 (N_260,In_363,In_88);
or U261 (N_261,In_177,In_643);
nand U262 (N_262,In_479,In_450);
or U263 (N_263,In_538,In_286);
and U264 (N_264,In_398,In_756);
nand U265 (N_265,In_486,In_471);
nor U266 (N_266,In_231,In_281);
and U267 (N_267,In_86,In_3);
or U268 (N_268,In_153,In_371);
nor U269 (N_269,In_369,In_55);
or U270 (N_270,In_388,In_207);
and U271 (N_271,In_248,In_174);
nor U272 (N_272,In_728,In_92);
or U273 (N_273,In_812,In_445);
and U274 (N_274,In_378,In_411);
or U275 (N_275,In_672,In_612);
nand U276 (N_276,In_488,In_469);
xor U277 (N_277,In_431,In_73);
or U278 (N_278,In_61,In_921);
nand U279 (N_279,In_269,In_940);
or U280 (N_280,In_568,In_860);
nand U281 (N_281,In_972,In_74);
nand U282 (N_282,In_50,In_150);
or U283 (N_283,In_966,In_772);
nand U284 (N_284,In_649,In_652);
nand U285 (N_285,In_718,In_564);
and U286 (N_286,In_380,In_857);
or U287 (N_287,In_942,In_723);
and U288 (N_288,In_47,In_849);
or U289 (N_289,In_693,In_642);
and U290 (N_290,In_506,In_283);
nor U291 (N_291,In_654,In_509);
nor U292 (N_292,In_897,In_255);
nand U293 (N_293,In_992,In_774);
nand U294 (N_294,In_815,In_384);
nor U295 (N_295,In_444,In_190);
or U296 (N_296,In_540,In_732);
or U297 (N_297,In_87,In_35);
nand U298 (N_298,In_20,In_241);
or U299 (N_299,In_663,In_900);
or U300 (N_300,In_95,In_121);
nor U301 (N_301,In_863,In_144);
nor U302 (N_302,In_316,In_956);
nand U303 (N_303,In_233,In_982);
nor U304 (N_304,In_120,In_317);
nand U305 (N_305,In_350,In_490);
nand U306 (N_306,In_958,In_287);
nor U307 (N_307,In_859,In_926);
nand U308 (N_308,In_924,In_58);
or U309 (N_309,In_845,In_19);
nand U310 (N_310,In_596,In_767);
or U311 (N_311,In_798,In_324);
and U312 (N_312,In_4,In_357);
and U313 (N_313,In_531,In_796);
nand U314 (N_314,In_48,In_8);
or U315 (N_315,In_85,In_861);
nand U316 (N_316,In_36,In_302);
or U317 (N_317,In_69,In_808);
nand U318 (N_318,In_892,In_169);
and U319 (N_319,In_165,In_778);
nand U320 (N_320,In_361,In_228);
nor U321 (N_321,In_392,In_605);
nor U322 (N_322,In_963,In_414);
nand U323 (N_323,In_146,In_77);
or U324 (N_324,In_358,In_669);
and U325 (N_325,In_64,In_748);
or U326 (N_326,In_703,In_521);
nor U327 (N_327,In_402,In_129);
and U328 (N_328,In_711,In_633);
nor U329 (N_329,In_515,In_794);
and U330 (N_330,In_428,In_773);
nor U331 (N_331,In_166,In_809);
and U332 (N_332,In_638,In_339);
and U333 (N_333,In_973,In_45);
and U334 (N_334,In_192,In_562);
nand U335 (N_335,In_131,In_214);
xnor U336 (N_336,In_875,In_905);
nor U337 (N_337,In_510,In_232);
or U338 (N_338,In_331,In_31);
and U339 (N_339,In_567,In_698);
nand U340 (N_340,In_969,In_0);
nand U341 (N_341,In_184,In_412);
nor U342 (N_342,In_404,In_683);
and U343 (N_343,In_270,In_449);
nor U344 (N_344,In_9,In_950);
nor U345 (N_345,In_528,In_432);
or U346 (N_346,In_513,In_627);
and U347 (N_347,In_552,In_882);
nand U348 (N_348,In_500,In_15);
and U349 (N_349,In_262,In_725);
nor U350 (N_350,In_624,In_743);
nand U351 (N_351,In_142,In_313);
and U352 (N_352,In_178,In_291);
or U353 (N_353,In_602,In_804);
xor U354 (N_354,In_67,In_887);
nand U355 (N_355,In_198,In_720);
or U356 (N_356,In_440,In_377);
or U357 (N_357,In_588,In_667);
nor U358 (N_358,In_206,In_668);
nand U359 (N_359,In_186,In_97);
nor U360 (N_360,In_453,In_10);
nor U361 (N_361,In_345,In_976);
or U362 (N_362,In_366,In_597);
and U363 (N_363,In_727,In_688);
nor U364 (N_364,In_250,In_651);
and U365 (N_365,In_864,In_275);
nand U366 (N_366,In_205,In_832);
or U367 (N_367,In_103,In_517);
nor U368 (N_368,In_383,In_470);
nand U369 (N_369,In_807,In_931);
or U370 (N_370,In_280,In_467);
or U371 (N_371,In_425,In_481);
or U372 (N_372,In_620,In_716);
nor U373 (N_373,In_679,In_944);
nand U374 (N_374,In_894,In_307);
nand U375 (N_375,In_158,In_525);
nor U376 (N_376,In_872,In_869);
nand U377 (N_377,In_814,In_646);
and U378 (N_378,In_779,In_691);
nor U379 (N_379,In_337,In_607);
nor U380 (N_380,In_59,In_442);
and U381 (N_381,In_79,In_653);
and U382 (N_382,In_850,In_901);
nand U383 (N_383,In_590,In_674);
and U384 (N_384,In_534,In_387);
nand U385 (N_385,In_846,In_136);
xnor U386 (N_386,In_197,In_907);
or U387 (N_387,In_677,In_454);
nand U388 (N_388,In_699,In_603);
xor U389 (N_389,In_726,In_415);
nand U390 (N_390,In_985,In_309);
xor U391 (N_391,In_116,In_692);
nor U392 (N_392,In_416,In_708);
and U393 (N_393,In_128,In_593);
and U394 (N_394,In_418,In_873);
nand U395 (N_395,In_811,In_746);
or U396 (N_396,In_569,In_946);
nand U397 (N_397,In_959,In_484);
nand U398 (N_398,In_68,In_608);
nand U399 (N_399,In_342,In_724);
nand U400 (N_400,In_372,In_188);
or U401 (N_401,In_573,In_647);
and U402 (N_402,In_83,In_51);
and U403 (N_403,In_644,In_478);
and U404 (N_404,In_25,In_874);
nand U405 (N_405,In_975,In_461);
xnor U406 (N_406,In_670,In_276);
and U407 (N_407,In_715,In_899);
nor U408 (N_408,In_895,In_199);
nand U409 (N_409,In_618,In_542);
nor U410 (N_410,In_60,In_577);
nor U411 (N_411,In_561,In_7);
or U412 (N_412,In_298,In_676);
and U413 (N_413,In_78,In_742);
and U414 (N_414,In_606,In_954);
or U415 (N_415,In_57,In_657);
nor U416 (N_416,In_225,In_499);
nor U417 (N_417,In_557,In_296);
nand U418 (N_418,In_22,In_455);
and U419 (N_419,In_210,In_871);
nand U420 (N_420,In_322,In_962);
nand U421 (N_421,In_243,In_274);
or U422 (N_422,In_511,In_957);
or U423 (N_423,In_409,In_830);
nand U424 (N_424,In_194,In_876);
and U425 (N_425,In_584,In_406);
or U426 (N_426,In_758,In_998);
and U427 (N_427,In_648,In_213);
and U428 (N_428,In_13,In_694);
and U429 (N_429,In_848,In_826);
nor U430 (N_430,In_974,In_816);
nand U431 (N_431,In_278,In_637);
and U432 (N_432,In_112,In_512);
or U433 (N_433,In_14,In_762);
and U434 (N_434,In_227,In_710);
and U435 (N_435,In_379,In_908);
and U436 (N_436,In_707,In_139);
and U437 (N_437,In_258,In_978);
nor U438 (N_438,In_554,In_797);
nand U439 (N_439,In_162,In_482);
and U440 (N_440,In_968,In_335);
nand U441 (N_441,In_504,In_11);
or U442 (N_442,In_381,In_546);
nand U443 (N_443,In_75,In_505);
or U444 (N_444,In_147,In_741);
and U445 (N_445,In_456,In_984);
nand U446 (N_446,In_960,In_747);
nand U447 (N_447,In_52,In_570);
nor U448 (N_448,In_981,In_594);
nor U449 (N_449,In_204,In_522);
or U450 (N_450,In_239,In_793);
nand U451 (N_451,In_530,In_733);
or U452 (N_452,In_306,In_971);
and U453 (N_453,In_502,In_884);
nand U454 (N_454,In_839,In_256);
and U455 (N_455,In_394,In_934);
and U456 (N_456,In_180,In_508);
and U457 (N_457,In_224,In_6);
and U458 (N_458,In_196,In_460);
nand U459 (N_459,In_879,In_373);
nand U460 (N_460,In_771,In_911);
nand U461 (N_461,In_282,In_532);
and U462 (N_462,In_254,In_896);
and U463 (N_463,In_634,In_912);
or U464 (N_464,In_397,In_244);
or U465 (N_465,In_526,In_970);
or U466 (N_466,In_238,In_66);
and U467 (N_467,In_700,In_400);
and U468 (N_468,In_591,In_438);
nor U469 (N_469,In_273,In_236);
nor U470 (N_470,In_71,In_519);
nor U471 (N_471,In_212,In_734);
or U472 (N_472,In_890,In_979);
nor U473 (N_473,In_806,In_777);
or U474 (N_474,In_903,In_621);
nor U475 (N_475,In_157,In_947);
nor U476 (N_476,In_765,In_640);
and U477 (N_477,In_352,In_836);
or U478 (N_478,In_829,In_94);
or U479 (N_479,In_485,In_582);
nand U480 (N_480,In_176,In_26);
and U481 (N_481,In_219,In_107);
and U482 (N_482,In_576,In_503);
nand U483 (N_483,In_847,In_448);
or U484 (N_484,In_5,In_340);
and U485 (N_485,In_261,In_285);
nor U486 (N_486,In_182,In_422);
nand U487 (N_487,In_917,In_935);
nand U488 (N_488,In_356,In_410);
nor U489 (N_489,In_831,In_560);
or U490 (N_490,In_539,In_242);
nand U491 (N_491,In_354,In_33);
nor U492 (N_492,In_483,In_856);
and U493 (N_493,In_240,In_858);
xnor U494 (N_494,In_229,In_138);
nor U495 (N_495,In_737,In_838);
and U496 (N_496,In_687,In_330);
or U497 (N_497,In_810,In_927);
and U498 (N_498,In_39,In_996);
and U499 (N_499,In_226,In_516);
nand U500 (N_500,In_670,In_502);
or U501 (N_501,In_244,In_68);
nor U502 (N_502,In_403,In_123);
or U503 (N_503,In_208,In_834);
nor U504 (N_504,In_951,In_266);
nor U505 (N_505,In_385,In_366);
or U506 (N_506,In_560,In_475);
and U507 (N_507,In_710,In_900);
or U508 (N_508,In_878,In_171);
or U509 (N_509,In_327,In_219);
and U510 (N_510,In_721,In_129);
nor U511 (N_511,In_269,In_185);
nor U512 (N_512,In_208,In_459);
nand U513 (N_513,In_999,In_344);
and U514 (N_514,In_489,In_507);
or U515 (N_515,In_497,In_904);
nand U516 (N_516,In_396,In_398);
and U517 (N_517,In_483,In_958);
nor U518 (N_518,In_494,In_388);
nor U519 (N_519,In_317,In_558);
nor U520 (N_520,In_338,In_869);
or U521 (N_521,In_532,In_496);
and U522 (N_522,In_413,In_668);
and U523 (N_523,In_767,In_406);
and U524 (N_524,In_102,In_721);
nor U525 (N_525,In_51,In_21);
nand U526 (N_526,In_874,In_414);
and U527 (N_527,In_529,In_224);
nand U528 (N_528,In_138,In_924);
and U529 (N_529,In_547,In_442);
or U530 (N_530,In_8,In_71);
and U531 (N_531,In_73,In_417);
nand U532 (N_532,In_213,In_895);
nor U533 (N_533,In_822,In_399);
nand U534 (N_534,In_58,In_391);
nor U535 (N_535,In_797,In_285);
or U536 (N_536,In_628,In_255);
nor U537 (N_537,In_483,In_357);
or U538 (N_538,In_822,In_373);
and U539 (N_539,In_224,In_760);
nand U540 (N_540,In_241,In_770);
or U541 (N_541,In_916,In_110);
nor U542 (N_542,In_969,In_892);
or U543 (N_543,In_915,In_811);
nand U544 (N_544,In_953,In_963);
and U545 (N_545,In_687,In_406);
or U546 (N_546,In_579,In_216);
nand U547 (N_547,In_21,In_826);
or U548 (N_548,In_481,In_655);
nor U549 (N_549,In_566,In_942);
nor U550 (N_550,In_217,In_399);
or U551 (N_551,In_564,In_957);
nand U552 (N_552,In_725,In_745);
nand U553 (N_553,In_214,In_104);
or U554 (N_554,In_107,In_9);
or U555 (N_555,In_113,In_692);
nand U556 (N_556,In_672,In_159);
and U557 (N_557,In_553,In_10);
nand U558 (N_558,In_950,In_236);
nor U559 (N_559,In_600,In_290);
nand U560 (N_560,In_925,In_111);
nand U561 (N_561,In_945,In_340);
nor U562 (N_562,In_615,In_763);
nor U563 (N_563,In_220,In_828);
nand U564 (N_564,In_640,In_528);
or U565 (N_565,In_857,In_580);
nor U566 (N_566,In_450,In_236);
or U567 (N_567,In_872,In_733);
or U568 (N_568,In_394,In_676);
and U569 (N_569,In_473,In_401);
nor U570 (N_570,In_576,In_871);
nand U571 (N_571,In_819,In_677);
xnor U572 (N_572,In_476,In_193);
or U573 (N_573,In_322,In_628);
or U574 (N_574,In_15,In_120);
and U575 (N_575,In_636,In_92);
nor U576 (N_576,In_725,In_879);
nand U577 (N_577,In_926,In_898);
nor U578 (N_578,In_279,In_187);
nand U579 (N_579,In_582,In_334);
and U580 (N_580,In_988,In_663);
and U581 (N_581,In_372,In_925);
nand U582 (N_582,In_689,In_994);
and U583 (N_583,In_159,In_164);
or U584 (N_584,In_722,In_428);
nor U585 (N_585,In_120,In_955);
nand U586 (N_586,In_911,In_132);
nand U587 (N_587,In_524,In_184);
nor U588 (N_588,In_494,In_171);
nor U589 (N_589,In_900,In_359);
nor U590 (N_590,In_325,In_947);
or U591 (N_591,In_564,In_589);
or U592 (N_592,In_707,In_122);
or U593 (N_593,In_891,In_740);
nand U594 (N_594,In_716,In_893);
nor U595 (N_595,In_594,In_221);
nand U596 (N_596,In_506,In_415);
or U597 (N_597,In_105,In_566);
or U598 (N_598,In_96,In_328);
and U599 (N_599,In_257,In_501);
and U600 (N_600,In_729,In_833);
nand U601 (N_601,In_623,In_214);
or U602 (N_602,In_583,In_598);
nand U603 (N_603,In_80,In_327);
or U604 (N_604,In_551,In_644);
and U605 (N_605,In_842,In_692);
or U606 (N_606,In_689,In_737);
nand U607 (N_607,In_308,In_202);
and U608 (N_608,In_752,In_168);
nor U609 (N_609,In_238,In_826);
nor U610 (N_610,In_292,In_26);
or U611 (N_611,In_528,In_975);
nor U612 (N_612,In_159,In_982);
nor U613 (N_613,In_456,In_741);
nand U614 (N_614,In_312,In_786);
nand U615 (N_615,In_19,In_942);
nor U616 (N_616,In_376,In_78);
or U617 (N_617,In_851,In_489);
and U618 (N_618,In_431,In_679);
and U619 (N_619,In_371,In_825);
and U620 (N_620,In_189,In_521);
or U621 (N_621,In_191,In_855);
nand U622 (N_622,In_947,In_40);
or U623 (N_623,In_339,In_995);
or U624 (N_624,In_633,In_606);
and U625 (N_625,In_348,In_181);
nor U626 (N_626,In_30,In_703);
or U627 (N_627,In_498,In_210);
or U628 (N_628,In_823,In_953);
nor U629 (N_629,In_909,In_418);
and U630 (N_630,In_222,In_623);
or U631 (N_631,In_381,In_708);
or U632 (N_632,In_516,In_916);
or U633 (N_633,In_865,In_81);
or U634 (N_634,In_680,In_309);
and U635 (N_635,In_10,In_196);
nor U636 (N_636,In_230,In_316);
or U637 (N_637,In_601,In_680);
nor U638 (N_638,In_685,In_814);
and U639 (N_639,In_634,In_930);
nand U640 (N_640,In_698,In_160);
nor U641 (N_641,In_987,In_959);
or U642 (N_642,In_148,In_997);
nor U643 (N_643,In_270,In_65);
and U644 (N_644,In_799,In_718);
nor U645 (N_645,In_451,In_4);
or U646 (N_646,In_703,In_710);
nor U647 (N_647,In_938,In_986);
nand U648 (N_648,In_98,In_424);
and U649 (N_649,In_708,In_604);
and U650 (N_650,In_108,In_410);
nand U651 (N_651,In_409,In_908);
and U652 (N_652,In_313,In_564);
or U653 (N_653,In_809,In_126);
nor U654 (N_654,In_602,In_416);
or U655 (N_655,In_481,In_55);
or U656 (N_656,In_202,In_773);
nand U657 (N_657,In_103,In_293);
nand U658 (N_658,In_261,In_872);
or U659 (N_659,In_825,In_51);
nand U660 (N_660,In_418,In_637);
nor U661 (N_661,In_269,In_470);
nand U662 (N_662,In_942,In_658);
nor U663 (N_663,In_957,In_909);
nor U664 (N_664,In_559,In_218);
nor U665 (N_665,In_310,In_432);
or U666 (N_666,In_974,In_680);
and U667 (N_667,In_580,In_431);
nand U668 (N_668,In_745,In_21);
nand U669 (N_669,In_52,In_635);
and U670 (N_670,In_626,In_973);
nor U671 (N_671,In_67,In_525);
or U672 (N_672,In_433,In_274);
nand U673 (N_673,In_791,In_135);
or U674 (N_674,In_339,In_821);
nand U675 (N_675,In_110,In_307);
nor U676 (N_676,In_848,In_786);
nor U677 (N_677,In_439,In_380);
or U678 (N_678,In_461,In_608);
nor U679 (N_679,In_271,In_494);
nor U680 (N_680,In_768,In_627);
nor U681 (N_681,In_546,In_226);
or U682 (N_682,In_892,In_5);
nand U683 (N_683,In_435,In_811);
and U684 (N_684,In_444,In_710);
or U685 (N_685,In_159,In_724);
or U686 (N_686,In_23,In_325);
nor U687 (N_687,In_143,In_467);
or U688 (N_688,In_97,In_714);
or U689 (N_689,In_12,In_843);
nand U690 (N_690,In_821,In_959);
and U691 (N_691,In_40,In_761);
nor U692 (N_692,In_746,In_926);
or U693 (N_693,In_987,In_634);
or U694 (N_694,In_457,In_33);
nor U695 (N_695,In_590,In_884);
or U696 (N_696,In_90,In_467);
and U697 (N_697,In_863,In_62);
and U698 (N_698,In_881,In_487);
nor U699 (N_699,In_25,In_42);
nor U700 (N_700,In_842,In_220);
nor U701 (N_701,In_462,In_110);
nor U702 (N_702,In_494,In_789);
nor U703 (N_703,In_961,In_312);
or U704 (N_704,In_58,In_200);
xnor U705 (N_705,In_74,In_775);
or U706 (N_706,In_36,In_574);
nor U707 (N_707,In_156,In_194);
nor U708 (N_708,In_956,In_988);
and U709 (N_709,In_558,In_771);
or U710 (N_710,In_263,In_871);
nand U711 (N_711,In_826,In_637);
or U712 (N_712,In_154,In_60);
nand U713 (N_713,In_925,In_583);
and U714 (N_714,In_83,In_973);
and U715 (N_715,In_394,In_833);
nor U716 (N_716,In_261,In_298);
nor U717 (N_717,In_577,In_324);
and U718 (N_718,In_339,In_136);
or U719 (N_719,In_330,In_778);
or U720 (N_720,In_676,In_744);
nor U721 (N_721,In_991,In_246);
and U722 (N_722,In_320,In_266);
or U723 (N_723,In_56,In_857);
nand U724 (N_724,In_609,In_764);
or U725 (N_725,In_608,In_2);
nand U726 (N_726,In_338,In_694);
xnor U727 (N_727,In_797,In_224);
nor U728 (N_728,In_488,In_484);
or U729 (N_729,In_923,In_427);
nand U730 (N_730,In_293,In_332);
and U731 (N_731,In_152,In_552);
and U732 (N_732,In_415,In_959);
and U733 (N_733,In_58,In_220);
and U734 (N_734,In_701,In_715);
nor U735 (N_735,In_214,In_536);
nand U736 (N_736,In_153,In_893);
and U737 (N_737,In_265,In_76);
nand U738 (N_738,In_733,In_834);
nand U739 (N_739,In_641,In_815);
and U740 (N_740,In_550,In_595);
or U741 (N_741,In_729,In_199);
or U742 (N_742,In_893,In_391);
and U743 (N_743,In_522,In_534);
or U744 (N_744,In_283,In_431);
nand U745 (N_745,In_825,In_647);
nor U746 (N_746,In_680,In_193);
and U747 (N_747,In_705,In_906);
nand U748 (N_748,In_562,In_141);
and U749 (N_749,In_248,In_467);
or U750 (N_750,In_477,In_834);
or U751 (N_751,In_421,In_150);
nand U752 (N_752,In_241,In_308);
nor U753 (N_753,In_843,In_777);
and U754 (N_754,In_611,In_661);
or U755 (N_755,In_62,In_374);
nor U756 (N_756,In_85,In_661);
and U757 (N_757,In_806,In_427);
nor U758 (N_758,In_583,In_445);
and U759 (N_759,In_30,In_635);
and U760 (N_760,In_666,In_253);
nor U761 (N_761,In_656,In_645);
or U762 (N_762,In_430,In_869);
nand U763 (N_763,In_36,In_237);
nor U764 (N_764,In_980,In_523);
nand U765 (N_765,In_990,In_422);
nor U766 (N_766,In_820,In_238);
nor U767 (N_767,In_129,In_764);
nand U768 (N_768,In_364,In_60);
or U769 (N_769,In_680,In_649);
nor U770 (N_770,In_5,In_918);
and U771 (N_771,In_733,In_764);
and U772 (N_772,In_232,In_756);
and U773 (N_773,In_622,In_117);
and U774 (N_774,In_442,In_937);
or U775 (N_775,In_721,In_585);
nor U776 (N_776,In_933,In_992);
and U777 (N_777,In_936,In_967);
nand U778 (N_778,In_630,In_327);
or U779 (N_779,In_843,In_191);
nand U780 (N_780,In_392,In_116);
nand U781 (N_781,In_789,In_894);
nor U782 (N_782,In_727,In_210);
nor U783 (N_783,In_703,In_965);
and U784 (N_784,In_931,In_216);
nand U785 (N_785,In_837,In_880);
or U786 (N_786,In_845,In_761);
nand U787 (N_787,In_171,In_142);
nor U788 (N_788,In_157,In_156);
nand U789 (N_789,In_471,In_122);
or U790 (N_790,In_701,In_126);
nand U791 (N_791,In_494,In_397);
nand U792 (N_792,In_964,In_571);
and U793 (N_793,In_787,In_421);
nor U794 (N_794,In_67,In_680);
or U795 (N_795,In_868,In_28);
and U796 (N_796,In_406,In_139);
or U797 (N_797,In_45,In_106);
nand U798 (N_798,In_26,In_42);
nand U799 (N_799,In_916,In_173);
and U800 (N_800,In_516,In_790);
nand U801 (N_801,In_772,In_879);
nor U802 (N_802,In_616,In_300);
and U803 (N_803,In_147,In_318);
or U804 (N_804,In_87,In_606);
nand U805 (N_805,In_409,In_250);
nand U806 (N_806,In_619,In_694);
nand U807 (N_807,In_564,In_39);
nand U808 (N_808,In_798,In_682);
nor U809 (N_809,In_666,In_65);
xnor U810 (N_810,In_838,In_973);
nor U811 (N_811,In_498,In_9);
nor U812 (N_812,In_60,In_885);
nor U813 (N_813,In_117,In_391);
or U814 (N_814,In_296,In_759);
and U815 (N_815,In_998,In_136);
or U816 (N_816,In_499,In_653);
nand U817 (N_817,In_904,In_343);
nand U818 (N_818,In_483,In_561);
nor U819 (N_819,In_80,In_370);
and U820 (N_820,In_849,In_921);
and U821 (N_821,In_711,In_147);
nor U822 (N_822,In_976,In_968);
nand U823 (N_823,In_309,In_923);
nand U824 (N_824,In_8,In_807);
and U825 (N_825,In_771,In_136);
or U826 (N_826,In_437,In_490);
nor U827 (N_827,In_153,In_171);
nor U828 (N_828,In_878,In_91);
nor U829 (N_829,In_669,In_546);
nand U830 (N_830,In_641,In_809);
nand U831 (N_831,In_944,In_510);
and U832 (N_832,In_670,In_821);
nand U833 (N_833,In_247,In_627);
or U834 (N_834,In_266,In_326);
and U835 (N_835,In_905,In_933);
or U836 (N_836,In_904,In_934);
nand U837 (N_837,In_98,In_367);
and U838 (N_838,In_753,In_235);
and U839 (N_839,In_603,In_34);
or U840 (N_840,In_732,In_299);
nor U841 (N_841,In_79,In_654);
nand U842 (N_842,In_610,In_114);
nor U843 (N_843,In_103,In_350);
nand U844 (N_844,In_220,In_320);
or U845 (N_845,In_282,In_219);
and U846 (N_846,In_363,In_507);
nor U847 (N_847,In_400,In_714);
or U848 (N_848,In_499,In_861);
nand U849 (N_849,In_849,In_375);
nand U850 (N_850,In_200,In_873);
and U851 (N_851,In_81,In_940);
nor U852 (N_852,In_616,In_150);
nand U853 (N_853,In_352,In_229);
nor U854 (N_854,In_903,In_866);
and U855 (N_855,In_264,In_41);
or U856 (N_856,In_54,In_798);
and U857 (N_857,In_952,In_532);
or U858 (N_858,In_23,In_549);
nor U859 (N_859,In_311,In_690);
and U860 (N_860,In_243,In_603);
nand U861 (N_861,In_217,In_64);
or U862 (N_862,In_948,In_505);
or U863 (N_863,In_860,In_170);
nand U864 (N_864,In_165,In_87);
or U865 (N_865,In_171,In_824);
nor U866 (N_866,In_298,In_690);
nor U867 (N_867,In_599,In_182);
and U868 (N_868,In_221,In_518);
or U869 (N_869,In_649,In_895);
nor U870 (N_870,In_190,In_180);
nor U871 (N_871,In_477,In_398);
and U872 (N_872,In_354,In_206);
nor U873 (N_873,In_520,In_810);
nor U874 (N_874,In_309,In_115);
and U875 (N_875,In_892,In_848);
nand U876 (N_876,In_110,In_285);
nand U877 (N_877,In_710,In_685);
nand U878 (N_878,In_670,In_736);
or U879 (N_879,In_182,In_637);
or U880 (N_880,In_998,In_243);
or U881 (N_881,In_558,In_719);
or U882 (N_882,In_851,In_880);
nor U883 (N_883,In_693,In_198);
nand U884 (N_884,In_891,In_874);
nand U885 (N_885,In_766,In_27);
and U886 (N_886,In_584,In_385);
or U887 (N_887,In_340,In_866);
or U888 (N_888,In_484,In_512);
nor U889 (N_889,In_821,In_526);
or U890 (N_890,In_961,In_813);
or U891 (N_891,In_451,In_455);
nand U892 (N_892,In_174,In_964);
or U893 (N_893,In_3,In_635);
and U894 (N_894,In_981,In_722);
nand U895 (N_895,In_993,In_146);
nand U896 (N_896,In_61,In_67);
or U897 (N_897,In_501,In_707);
nor U898 (N_898,In_855,In_23);
or U899 (N_899,In_216,In_31);
nand U900 (N_900,In_376,In_288);
nand U901 (N_901,In_41,In_437);
or U902 (N_902,In_940,In_846);
nand U903 (N_903,In_758,In_92);
nor U904 (N_904,In_266,In_374);
or U905 (N_905,In_695,In_24);
nor U906 (N_906,In_567,In_697);
nor U907 (N_907,In_538,In_274);
nor U908 (N_908,In_273,In_842);
nand U909 (N_909,In_943,In_702);
and U910 (N_910,In_377,In_412);
and U911 (N_911,In_30,In_36);
or U912 (N_912,In_217,In_491);
or U913 (N_913,In_29,In_624);
nor U914 (N_914,In_599,In_427);
and U915 (N_915,In_186,In_318);
nand U916 (N_916,In_995,In_394);
or U917 (N_917,In_654,In_534);
nor U918 (N_918,In_993,In_337);
nand U919 (N_919,In_354,In_707);
and U920 (N_920,In_805,In_676);
nor U921 (N_921,In_675,In_264);
and U922 (N_922,In_226,In_688);
xor U923 (N_923,In_985,In_841);
and U924 (N_924,In_831,In_471);
and U925 (N_925,In_271,In_937);
nor U926 (N_926,In_249,In_87);
and U927 (N_927,In_914,In_343);
nor U928 (N_928,In_98,In_296);
nand U929 (N_929,In_491,In_400);
nor U930 (N_930,In_338,In_268);
and U931 (N_931,In_236,In_366);
nand U932 (N_932,In_183,In_370);
nand U933 (N_933,In_335,In_956);
or U934 (N_934,In_755,In_816);
nor U935 (N_935,In_359,In_982);
and U936 (N_936,In_91,In_595);
nand U937 (N_937,In_709,In_462);
and U938 (N_938,In_653,In_732);
nand U939 (N_939,In_969,In_404);
nor U940 (N_940,In_21,In_308);
and U941 (N_941,In_251,In_437);
or U942 (N_942,In_683,In_887);
or U943 (N_943,In_225,In_907);
and U944 (N_944,In_182,In_866);
nand U945 (N_945,In_622,In_16);
or U946 (N_946,In_648,In_938);
nor U947 (N_947,In_751,In_937);
nor U948 (N_948,In_923,In_24);
nor U949 (N_949,In_281,In_807);
nand U950 (N_950,In_783,In_661);
nor U951 (N_951,In_219,In_916);
nand U952 (N_952,In_773,In_811);
or U953 (N_953,In_239,In_576);
or U954 (N_954,In_74,In_210);
nor U955 (N_955,In_32,In_734);
or U956 (N_956,In_183,In_450);
nor U957 (N_957,In_512,In_872);
nor U958 (N_958,In_239,In_837);
and U959 (N_959,In_493,In_655);
or U960 (N_960,In_429,In_401);
nor U961 (N_961,In_445,In_494);
or U962 (N_962,In_529,In_527);
nor U963 (N_963,In_530,In_930);
or U964 (N_964,In_711,In_921);
and U965 (N_965,In_816,In_642);
or U966 (N_966,In_661,In_259);
nand U967 (N_967,In_151,In_581);
or U968 (N_968,In_69,In_903);
nor U969 (N_969,In_795,In_94);
or U970 (N_970,In_141,In_916);
and U971 (N_971,In_28,In_917);
or U972 (N_972,In_619,In_686);
nand U973 (N_973,In_131,In_836);
nand U974 (N_974,In_26,In_108);
nor U975 (N_975,In_376,In_351);
nand U976 (N_976,In_873,In_474);
and U977 (N_977,In_199,In_644);
nand U978 (N_978,In_11,In_2);
nand U979 (N_979,In_333,In_491);
nand U980 (N_980,In_352,In_76);
nand U981 (N_981,In_781,In_78);
or U982 (N_982,In_861,In_551);
xor U983 (N_983,In_829,In_568);
or U984 (N_984,In_54,In_958);
nand U985 (N_985,In_207,In_211);
and U986 (N_986,In_645,In_267);
nand U987 (N_987,In_858,In_539);
or U988 (N_988,In_959,In_619);
nand U989 (N_989,In_517,In_160);
nor U990 (N_990,In_991,In_338);
nor U991 (N_991,In_27,In_228);
nand U992 (N_992,In_775,In_234);
or U993 (N_993,In_526,In_185);
and U994 (N_994,In_316,In_857);
and U995 (N_995,In_546,In_362);
or U996 (N_996,In_115,In_999);
or U997 (N_997,In_351,In_81);
nor U998 (N_998,In_788,In_661);
nand U999 (N_999,In_331,In_380);
and U1000 (N_1000,N_0,N_565);
nand U1001 (N_1001,N_814,N_224);
nor U1002 (N_1002,N_414,N_885);
and U1003 (N_1003,N_989,N_664);
or U1004 (N_1004,N_98,N_43);
nor U1005 (N_1005,N_539,N_941);
or U1006 (N_1006,N_732,N_415);
or U1007 (N_1007,N_643,N_581);
or U1008 (N_1008,N_940,N_293);
or U1009 (N_1009,N_708,N_49);
or U1010 (N_1010,N_891,N_689);
or U1011 (N_1011,N_783,N_321);
or U1012 (N_1012,N_560,N_629);
nor U1013 (N_1013,N_217,N_747);
and U1014 (N_1014,N_406,N_786);
nor U1015 (N_1015,N_3,N_880);
and U1016 (N_1016,N_151,N_713);
nor U1017 (N_1017,N_192,N_384);
nor U1018 (N_1018,N_930,N_805);
and U1019 (N_1019,N_846,N_834);
or U1020 (N_1020,N_503,N_420);
and U1021 (N_1021,N_286,N_662);
or U1022 (N_1022,N_199,N_407);
nand U1023 (N_1023,N_934,N_781);
nor U1024 (N_1024,N_787,N_370);
nand U1025 (N_1025,N_889,N_301);
nor U1026 (N_1026,N_433,N_493);
and U1027 (N_1027,N_990,N_150);
and U1028 (N_1028,N_167,N_588);
nor U1029 (N_1029,N_669,N_660);
nor U1030 (N_1030,N_602,N_774);
or U1031 (N_1031,N_211,N_35);
nand U1032 (N_1032,N_633,N_559);
nand U1033 (N_1033,N_145,N_120);
or U1034 (N_1034,N_634,N_296);
nand U1035 (N_1035,N_163,N_1);
nor U1036 (N_1036,N_209,N_147);
and U1037 (N_1037,N_811,N_182);
or U1038 (N_1038,N_975,N_96);
nor U1039 (N_1039,N_677,N_297);
or U1040 (N_1040,N_339,N_412);
or U1041 (N_1041,N_850,N_491);
nor U1042 (N_1042,N_733,N_349);
nand U1043 (N_1043,N_695,N_482);
and U1044 (N_1044,N_920,N_128);
nand U1045 (N_1045,N_443,N_70);
and U1046 (N_1046,N_603,N_121);
and U1047 (N_1047,N_290,N_952);
nor U1048 (N_1048,N_912,N_427);
or U1049 (N_1049,N_612,N_607);
or U1050 (N_1050,N_939,N_99);
nand U1051 (N_1051,N_827,N_76);
nor U1052 (N_1052,N_968,N_678);
and U1053 (N_1053,N_337,N_379);
nand U1054 (N_1054,N_874,N_501);
xor U1055 (N_1055,N_248,N_39);
nor U1056 (N_1056,N_102,N_777);
or U1057 (N_1057,N_294,N_212);
nor U1058 (N_1058,N_135,N_426);
and U1059 (N_1059,N_674,N_470);
nor U1060 (N_1060,N_778,N_116);
nor U1061 (N_1061,N_508,N_382);
nand U1062 (N_1062,N_769,N_84);
and U1063 (N_1063,N_467,N_568);
nand U1064 (N_1064,N_574,N_410);
nand U1065 (N_1065,N_276,N_46);
and U1066 (N_1066,N_620,N_567);
and U1067 (N_1067,N_916,N_861);
and U1068 (N_1068,N_396,N_269);
or U1069 (N_1069,N_868,N_10);
nor U1070 (N_1070,N_762,N_447);
nor U1071 (N_1071,N_322,N_621);
nand U1072 (N_1072,N_108,N_802);
nor U1073 (N_1073,N_551,N_970);
xnor U1074 (N_1074,N_562,N_441);
nor U1075 (N_1075,N_373,N_71);
nand U1076 (N_1076,N_820,N_275);
or U1077 (N_1077,N_371,N_899);
nor U1078 (N_1078,N_41,N_942);
nor U1079 (N_1079,N_174,N_351);
and U1080 (N_1080,N_37,N_927);
nand U1081 (N_1081,N_91,N_268);
nand U1082 (N_1082,N_526,N_854);
and U1083 (N_1083,N_530,N_318);
xnor U1084 (N_1084,N_255,N_724);
and U1085 (N_1085,N_515,N_595);
nor U1086 (N_1086,N_364,N_188);
nand U1087 (N_1087,N_655,N_399);
or U1088 (N_1088,N_862,N_273);
nor U1089 (N_1089,N_401,N_578);
and U1090 (N_1090,N_898,N_830);
or U1091 (N_1091,N_59,N_334);
or U1092 (N_1092,N_89,N_50);
and U1093 (N_1093,N_693,N_254);
nor U1094 (N_1094,N_859,N_863);
nand U1095 (N_1095,N_365,N_32);
nor U1096 (N_1096,N_881,N_274);
nand U1097 (N_1097,N_137,N_969);
nand U1098 (N_1098,N_743,N_536);
nand U1099 (N_1099,N_234,N_68);
or U1100 (N_1100,N_505,N_516);
nand U1101 (N_1101,N_718,N_625);
nor U1102 (N_1102,N_421,N_358);
nor U1103 (N_1103,N_598,N_40);
and U1104 (N_1104,N_913,N_646);
or U1105 (N_1105,N_701,N_134);
and U1106 (N_1106,N_237,N_519);
nor U1107 (N_1107,N_973,N_395);
nand U1108 (N_1108,N_178,N_631);
and U1109 (N_1109,N_492,N_672);
and U1110 (N_1110,N_146,N_24);
nand U1111 (N_1111,N_23,N_205);
nand U1112 (N_1112,N_459,N_264);
nor U1113 (N_1113,N_311,N_465);
or U1114 (N_1114,N_618,N_887);
and U1115 (N_1115,N_753,N_51);
nand U1116 (N_1116,N_538,N_330);
and U1117 (N_1117,N_183,N_152);
nand U1118 (N_1118,N_79,N_947);
nand U1119 (N_1119,N_717,N_902);
and U1120 (N_1120,N_408,N_511);
nand U1121 (N_1121,N_184,N_550);
nor U1122 (N_1122,N_36,N_833);
and U1123 (N_1123,N_794,N_908);
and U1124 (N_1124,N_796,N_791);
or U1125 (N_1125,N_488,N_865);
nand U1126 (N_1126,N_935,N_844);
or U1127 (N_1127,N_422,N_556);
and U1128 (N_1128,N_552,N_261);
nor U1129 (N_1129,N_176,N_142);
and U1130 (N_1130,N_469,N_139);
nand U1131 (N_1131,N_162,N_265);
nand U1132 (N_1132,N_309,N_510);
or U1133 (N_1133,N_165,N_333);
and U1134 (N_1134,N_876,N_586);
nand U1135 (N_1135,N_615,N_476);
nand U1136 (N_1136,N_57,N_825);
and U1137 (N_1137,N_428,N_460);
or U1138 (N_1138,N_292,N_55);
nor U1139 (N_1139,N_374,N_991);
nor U1140 (N_1140,N_231,N_228);
nor U1141 (N_1141,N_676,N_792);
nand U1142 (N_1142,N_785,N_189);
nor U1143 (N_1143,N_534,N_543);
and U1144 (N_1144,N_700,N_303);
nand U1145 (N_1145,N_155,N_573);
or U1146 (N_1146,N_438,N_62);
and U1147 (N_1147,N_285,N_434);
nand U1148 (N_1148,N_808,N_979);
nor U1149 (N_1149,N_557,N_996);
and U1150 (N_1150,N_517,N_824);
nor U1151 (N_1151,N_725,N_613);
nor U1152 (N_1152,N_685,N_879);
nor U1153 (N_1153,N_886,N_64);
or U1154 (N_1154,N_338,N_627);
and U1155 (N_1155,N_432,N_749);
and U1156 (N_1156,N_957,N_981);
nor U1157 (N_1157,N_316,N_815);
or U1158 (N_1158,N_765,N_113);
or U1159 (N_1159,N_649,N_226);
or U1160 (N_1160,N_962,N_897);
and U1161 (N_1161,N_352,N_362);
nor U1162 (N_1162,N_400,N_439);
nand U1163 (N_1163,N_263,N_727);
nor U1164 (N_1164,N_809,N_758);
or U1165 (N_1165,N_473,N_754);
nor U1166 (N_1166,N_33,N_463);
nor U1167 (N_1167,N_249,N_936);
nand U1168 (N_1168,N_85,N_350);
nor U1169 (N_1169,N_2,N_435);
nand U1170 (N_1170,N_838,N_326);
and U1171 (N_1171,N_30,N_673);
nor U1172 (N_1172,N_101,N_699);
nor U1173 (N_1173,N_983,N_992);
and U1174 (N_1174,N_911,N_54);
or U1175 (N_1175,N_641,N_768);
nor U1176 (N_1176,N_284,N_583);
nor U1177 (N_1177,N_784,N_654);
nand U1178 (N_1178,N_525,N_741);
nand U1179 (N_1179,N_289,N_164);
or U1180 (N_1180,N_506,N_766);
and U1181 (N_1181,N_393,N_715);
or U1182 (N_1182,N_481,N_88);
and U1183 (N_1183,N_616,N_884);
or U1184 (N_1184,N_215,N_335);
nand U1185 (N_1185,N_256,N_949);
nand U1186 (N_1186,N_353,N_458);
or U1187 (N_1187,N_582,N_974);
nand U1188 (N_1188,N_26,N_245);
nand U1189 (N_1189,N_545,N_580);
nand U1190 (N_1190,N_278,N_214);
and U1191 (N_1191,N_186,N_541);
nand U1192 (N_1192,N_168,N_999);
and U1193 (N_1193,N_806,N_247);
nand U1194 (N_1194,N_721,N_319);
or U1195 (N_1195,N_728,N_735);
nand U1196 (N_1196,N_376,N_527);
and U1197 (N_1197,N_836,N_789);
and U1198 (N_1198,N_489,N_356);
nand U1199 (N_1199,N_775,N_687);
nand U1200 (N_1200,N_124,N_663);
nand U1201 (N_1201,N_544,N_67);
or U1202 (N_1202,N_554,N_93);
or U1203 (N_1203,N_956,N_344);
nand U1204 (N_1204,N_771,N_388);
and U1205 (N_1205,N_698,N_7);
nand U1206 (N_1206,N_72,N_853);
nor U1207 (N_1207,N_558,N_471);
and U1208 (N_1208,N_608,N_829);
nand U1209 (N_1209,N_227,N_922);
nand U1210 (N_1210,N_115,N_590);
or U1211 (N_1211,N_16,N_12);
nand U1212 (N_1212,N_528,N_266);
and U1213 (N_1213,N_710,N_524);
nand U1214 (N_1214,N_206,N_372);
or U1215 (N_1215,N_359,N_252);
and U1216 (N_1216,N_900,N_295);
or U1217 (N_1217,N_203,N_790);
or U1218 (N_1218,N_591,N_976);
nand U1219 (N_1219,N_5,N_832);
or U1220 (N_1220,N_800,N_716);
nor U1221 (N_1221,N_213,N_682);
or U1222 (N_1222,N_100,N_823);
nor U1223 (N_1223,N_965,N_614);
or U1224 (N_1224,N_60,N_759);
and U1225 (N_1225,N_204,N_866);
and U1226 (N_1226,N_229,N_915);
nor U1227 (N_1227,N_392,N_628);
nand U1228 (N_1228,N_430,N_657);
nand U1229 (N_1229,N_703,N_816);
nor U1230 (N_1230,N_720,N_149);
and U1231 (N_1231,N_380,N_65);
or U1232 (N_1232,N_734,N_253);
nand U1233 (N_1233,N_890,N_925);
nor U1234 (N_1234,N_684,N_175);
and U1235 (N_1235,N_485,N_757);
nor U1236 (N_1236,N_619,N_332);
and U1237 (N_1237,N_413,N_737);
and U1238 (N_1238,N_875,N_112);
and U1239 (N_1239,N_325,N_110);
nor U1240 (N_1240,N_719,N_455);
and U1241 (N_1241,N_445,N_444);
nand U1242 (N_1242,N_161,N_118);
and U1243 (N_1243,N_86,N_540);
nand U1244 (N_1244,N_196,N_869);
nand U1245 (N_1245,N_394,N_532);
nor U1246 (N_1246,N_202,N_688);
nand U1247 (N_1247,N_431,N_232);
or U1248 (N_1248,N_772,N_369);
nand U1249 (N_1249,N_377,N_883);
nand U1250 (N_1250,N_592,N_826);
and U1251 (N_1251,N_529,N_730);
and U1252 (N_1252,N_222,N_236);
nor U1253 (N_1253,N_642,N_726);
or U1254 (N_1254,N_328,N_281);
and U1255 (N_1255,N_129,N_917);
and U1256 (N_1256,N_773,N_748);
nand U1257 (N_1257,N_675,N_450);
nor U1258 (N_1258,N_92,N_429);
or U1259 (N_1259,N_804,N_670);
nand U1260 (N_1260,N_363,N_442);
or U1261 (N_1261,N_610,N_200);
or U1262 (N_1262,N_244,N_323);
nor U1263 (N_1263,N_819,N_304);
and U1264 (N_1264,N_90,N_307);
nand U1265 (N_1265,N_645,N_170);
or U1266 (N_1266,N_453,N_52);
and U1267 (N_1267,N_402,N_136);
xor U1268 (N_1268,N_15,N_343);
nor U1269 (N_1269,N_653,N_896);
nor U1270 (N_1270,N_324,N_951);
or U1271 (N_1271,N_13,N_190);
and U1272 (N_1272,N_533,N_801);
or U1273 (N_1273,N_490,N_246);
nand U1274 (N_1274,N_572,N_746);
and U1275 (N_1275,N_667,N_597);
or U1276 (N_1276,N_843,N_822);
nand U1277 (N_1277,N_988,N_767);
or U1278 (N_1278,N_74,N_243);
nor U1279 (N_1279,N_187,N_53);
or U1280 (N_1280,N_484,N_561);
nand U1281 (N_1281,N_357,N_694);
nor U1282 (N_1282,N_740,N_346);
nand U1283 (N_1283,N_872,N_260);
xor U1284 (N_1284,N_919,N_122);
nand U1285 (N_1285,N_873,N_456);
and U1286 (N_1286,N_61,N_201);
or U1287 (N_1287,N_622,N_867);
and U1288 (N_1288,N_738,N_918);
nor U1289 (N_1289,N_223,N_666);
nand U1290 (N_1290,N_739,N_812);
nor U1291 (N_1291,N_953,N_821);
or U1292 (N_1292,N_605,N_640);
nand U1293 (N_1293,N_810,N_665);
or U1294 (N_1294,N_994,N_302);
xnor U1295 (N_1295,N_141,N_436);
nand U1296 (N_1296,N_828,N_195);
or U1297 (N_1297,N_119,N_692);
nand U1298 (N_1298,N_144,N_966);
nand U1299 (N_1299,N_18,N_87);
nand U1300 (N_1300,N_709,N_271);
nand U1301 (N_1301,N_950,N_892);
nand U1302 (N_1302,N_690,N_258);
and U1303 (N_1303,N_702,N_305);
and U1304 (N_1304,N_239,N_138);
nand U1305 (N_1305,N_932,N_73);
or U1306 (N_1306,N_272,N_417);
nor U1307 (N_1307,N_345,N_914);
nor U1308 (N_1308,N_893,N_924);
xnor U1309 (N_1309,N_910,N_472);
nand U1310 (N_1310,N_44,N_241);
and U1311 (N_1311,N_423,N_986);
nor U1312 (N_1312,N_398,N_107);
and U1313 (N_1313,N_210,N_750);
and U1314 (N_1314,N_331,N_977);
and U1315 (N_1315,N_300,N_287);
or U1316 (N_1316,N_596,N_20);
or U1317 (N_1317,N_267,N_982);
nor U1318 (N_1318,N_587,N_440);
and U1319 (N_1319,N_779,N_995);
nand U1320 (N_1320,N_475,N_114);
nor U1321 (N_1321,N_944,N_926);
nor U1322 (N_1322,N_327,N_83);
and U1323 (N_1323,N_509,N_943);
or U1324 (N_1324,N_133,N_230);
nand U1325 (N_1325,N_28,N_360);
nand U1326 (N_1326,N_166,N_208);
and U1327 (N_1327,N_148,N_523);
and U1328 (N_1328,N_960,N_419);
nor U1329 (N_1329,N_9,N_75);
and U1330 (N_1330,N_466,N_817);
and U1331 (N_1331,N_803,N_894);
nand U1332 (N_1332,N_385,N_126);
or U1333 (N_1333,N_909,N_576);
nor U1334 (N_1334,N_548,N_831);
nand U1335 (N_1335,N_348,N_946);
or U1336 (N_1336,N_668,N_797);
and U1337 (N_1337,N_594,N_159);
nand U1338 (N_1338,N_366,N_888);
and U1339 (N_1339,N_948,N_630);
and U1340 (N_1340,N_347,N_11);
and U1341 (N_1341,N_298,N_744);
nand U1342 (N_1342,N_937,N_585);
or U1343 (N_1343,N_848,N_375);
nor U1344 (N_1344,N_78,N_27);
or U1345 (N_1345,N_604,N_745);
xor U1346 (N_1346,N_468,N_870);
nor U1347 (N_1347,N_81,N_570);
and U1348 (N_1348,N_218,N_635);
and U1349 (N_1349,N_923,N_354);
xnor U1350 (N_1350,N_25,N_457);
nor U1351 (N_1351,N_17,N_381);
or U1352 (N_1352,N_140,N_707);
nand U1353 (N_1353,N_462,N_221);
nor U1354 (N_1354,N_499,N_632);
or U1355 (N_1355,N_411,N_279);
and U1356 (N_1356,N_104,N_63);
or U1357 (N_1357,N_21,N_479);
nand U1358 (N_1358,N_569,N_575);
nand U1359 (N_1359,N_967,N_593);
nand U1360 (N_1360,N_626,N_555);
and U1361 (N_1361,N_907,N_714);
or U1362 (N_1362,N_959,N_842);
and U1363 (N_1363,N_242,N_259);
and U1364 (N_1364,N_696,N_277);
or U1365 (N_1365,N_518,N_66);
or U1366 (N_1366,N_520,N_882);
and U1367 (N_1367,N_6,N_452);
nand U1368 (N_1368,N_798,N_644);
nor U1369 (N_1369,N_931,N_955);
or U1370 (N_1370,N_405,N_314);
or U1371 (N_1371,N_845,N_310);
or U1372 (N_1372,N_34,N_95);
and U1373 (N_1373,N_609,N_171);
or U1374 (N_1374,N_425,N_424);
nand U1375 (N_1375,N_513,N_340);
or U1376 (N_1376,N_185,N_22);
nor U1377 (N_1377,N_160,N_451);
or U1378 (N_1378,N_97,N_507);
and U1379 (N_1379,N_980,N_599);
and U1380 (N_1380,N_722,N_963);
and U1381 (N_1381,N_542,N_378);
and U1382 (N_1382,N_742,N_764);
and U1383 (N_1383,N_45,N_387);
nor U1384 (N_1384,N_198,N_193);
or U1385 (N_1385,N_220,N_82);
nor U1386 (N_1386,N_125,N_928);
nor U1387 (N_1387,N_601,N_958);
and U1388 (N_1388,N_47,N_656);
nand U1389 (N_1389,N_961,N_156);
nand U1390 (N_1390,N_905,N_240);
nand U1391 (N_1391,N_502,N_871);
nor U1392 (N_1392,N_409,N_933);
nor U1393 (N_1393,N_282,N_29);
or U1394 (N_1394,N_477,N_807);
or U1395 (N_1395,N_130,N_997);
and U1396 (N_1396,N_712,N_761);
nor U1397 (N_1397,N_404,N_449);
nand U1398 (N_1398,N_31,N_855);
or U1399 (N_1399,N_751,N_480);
and U1400 (N_1400,N_317,N_571);
nor U1401 (N_1401,N_782,N_257);
or U1402 (N_1402,N_547,N_857);
nand U1403 (N_1403,N_535,N_877);
nor U1404 (N_1404,N_904,N_341);
nand U1405 (N_1405,N_799,N_180);
or U1406 (N_1406,N_978,N_238);
nor U1407 (N_1407,N_624,N_964);
nand U1408 (N_1408,N_756,N_839);
nor U1409 (N_1409,N_531,N_658);
nor U1410 (N_1410,N_549,N_383);
and U1411 (N_1411,N_397,N_197);
or U1412 (N_1412,N_522,N_512);
or U1413 (N_1413,N_921,N_671);
and U1414 (N_1414,N_878,N_906);
and U1415 (N_1415,N_111,N_474);
and U1416 (N_1416,N_4,N_19);
nor U1417 (N_1417,N_320,N_945);
and U1418 (N_1418,N_683,N_313);
nand U1419 (N_1419,N_901,N_563);
or U1420 (N_1420,N_851,N_355);
or U1421 (N_1421,N_250,N_342);
nor U1422 (N_1422,N_752,N_483);
nor U1423 (N_1423,N_858,N_418);
nand U1424 (N_1424,N_566,N_390);
nor U1425 (N_1425,N_659,N_391);
or U1426 (N_1426,N_611,N_938);
nor U1427 (N_1427,N_650,N_280);
or U1428 (N_1428,N_486,N_731);
and U1429 (N_1429,N_661,N_299);
or U1430 (N_1430,N_971,N_852);
nor U1431 (N_1431,N_686,N_308);
nor U1432 (N_1432,N_216,N_14);
or U1433 (N_1433,N_361,N_153);
or U1434 (N_1434,N_389,N_172);
nor U1435 (N_1435,N_315,N_648);
nor U1436 (N_1436,N_521,N_584);
or U1437 (N_1437,N_312,N_984);
nand U1438 (N_1438,N_169,N_793);
and U1439 (N_1439,N_94,N_579);
nand U1440 (N_1440,N_847,N_157);
or U1441 (N_1441,N_127,N_8);
nor U1442 (N_1442,N_763,N_514);
nand U1443 (N_1443,N_58,N_494);
and U1444 (N_1444,N_132,N_623);
or U1445 (N_1445,N_207,N_697);
and U1446 (N_1446,N_705,N_651);
or U1447 (N_1447,N_291,N_813);
and U1448 (N_1448,N_564,N_849);
and U1449 (N_1449,N_818,N_235);
nor U1450 (N_1450,N_448,N_639);
nor U1451 (N_1451,N_856,N_446);
or U1452 (N_1452,N_788,N_283);
and U1453 (N_1453,N_498,N_553);
nor U1454 (N_1454,N_77,N_454);
nor U1455 (N_1455,N_841,N_497);
and U1456 (N_1456,N_589,N_181);
and U1457 (N_1457,N_679,N_681);
nand U1458 (N_1458,N_600,N_367);
and U1459 (N_1459,N_478,N_251);
nand U1460 (N_1460,N_680,N_106);
or U1461 (N_1461,N_306,N_770);
and U1462 (N_1462,N_537,N_80);
and U1463 (N_1463,N_416,N_606);
nand U1464 (N_1464,N_336,N_48);
nor U1465 (N_1465,N_500,N_903);
nor U1466 (N_1466,N_496,N_56);
nand U1467 (N_1467,N_495,N_103);
nor U1468 (N_1468,N_636,N_191);
and U1469 (N_1469,N_895,N_225);
and U1470 (N_1470,N_131,N_42);
nor U1471 (N_1471,N_487,N_329);
nor U1472 (N_1472,N_617,N_109);
nand U1473 (N_1473,N_638,N_706);
nand U1474 (N_1474,N_736,N_577);
or U1475 (N_1475,N_158,N_647);
nand U1476 (N_1476,N_173,N_38);
and U1477 (N_1477,N_755,N_864);
nand U1478 (N_1478,N_546,N_840);
and U1479 (N_1479,N_760,N_117);
or U1480 (N_1480,N_723,N_177);
nor U1481 (N_1481,N_504,N_929);
nand U1482 (N_1482,N_652,N_437);
or U1483 (N_1483,N_233,N_219);
or U1484 (N_1484,N_860,N_123);
or U1485 (N_1485,N_998,N_837);
or U1486 (N_1486,N_795,N_711);
nand U1487 (N_1487,N_69,N_262);
or U1488 (N_1488,N_461,N_403);
and U1489 (N_1489,N_985,N_704);
xor U1490 (N_1490,N_835,N_776);
or U1491 (N_1491,N_691,N_464);
or U1492 (N_1492,N_987,N_105);
and U1493 (N_1493,N_729,N_993);
nand U1494 (N_1494,N_780,N_386);
or U1495 (N_1495,N_368,N_954);
nor U1496 (N_1496,N_288,N_972);
and U1497 (N_1497,N_194,N_637);
or U1498 (N_1498,N_154,N_179);
nor U1499 (N_1499,N_270,N_143);
nand U1500 (N_1500,N_273,N_40);
or U1501 (N_1501,N_228,N_944);
nand U1502 (N_1502,N_9,N_893);
or U1503 (N_1503,N_20,N_984);
nand U1504 (N_1504,N_288,N_311);
or U1505 (N_1505,N_590,N_421);
nand U1506 (N_1506,N_658,N_67);
or U1507 (N_1507,N_566,N_335);
and U1508 (N_1508,N_722,N_426);
and U1509 (N_1509,N_821,N_962);
or U1510 (N_1510,N_522,N_786);
nand U1511 (N_1511,N_571,N_161);
and U1512 (N_1512,N_258,N_614);
and U1513 (N_1513,N_269,N_577);
nand U1514 (N_1514,N_588,N_345);
nor U1515 (N_1515,N_335,N_332);
nand U1516 (N_1516,N_102,N_793);
nor U1517 (N_1517,N_655,N_788);
nand U1518 (N_1518,N_900,N_140);
nor U1519 (N_1519,N_597,N_567);
or U1520 (N_1520,N_777,N_56);
or U1521 (N_1521,N_210,N_973);
nand U1522 (N_1522,N_829,N_447);
nand U1523 (N_1523,N_131,N_1);
or U1524 (N_1524,N_261,N_417);
nor U1525 (N_1525,N_598,N_462);
or U1526 (N_1526,N_474,N_193);
nand U1527 (N_1527,N_161,N_675);
nand U1528 (N_1528,N_900,N_808);
nor U1529 (N_1529,N_507,N_531);
and U1530 (N_1530,N_685,N_940);
nand U1531 (N_1531,N_686,N_761);
or U1532 (N_1532,N_50,N_533);
nand U1533 (N_1533,N_285,N_158);
or U1534 (N_1534,N_966,N_741);
and U1535 (N_1535,N_934,N_968);
and U1536 (N_1536,N_649,N_272);
nor U1537 (N_1537,N_507,N_557);
nand U1538 (N_1538,N_697,N_982);
nor U1539 (N_1539,N_274,N_632);
or U1540 (N_1540,N_322,N_688);
nand U1541 (N_1541,N_930,N_744);
nor U1542 (N_1542,N_587,N_74);
and U1543 (N_1543,N_538,N_760);
nor U1544 (N_1544,N_700,N_106);
and U1545 (N_1545,N_155,N_893);
nor U1546 (N_1546,N_639,N_462);
nand U1547 (N_1547,N_450,N_366);
or U1548 (N_1548,N_63,N_146);
or U1549 (N_1549,N_208,N_28);
nor U1550 (N_1550,N_434,N_589);
and U1551 (N_1551,N_263,N_52);
or U1552 (N_1552,N_220,N_150);
or U1553 (N_1553,N_104,N_448);
nand U1554 (N_1554,N_872,N_574);
nand U1555 (N_1555,N_998,N_318);
nand U1556 (N_1556,N_119,N_461);
or U1557 (N_1557,N_552,N_731);
and U1558 (N_1558,N_429,N_484);
nor U1559 (N_1559,N_216,N_722);
nand U1560 (N_1560,N_682,N_970);
and U1561 (N_1561,N_328,N_434);
nand U1562 (N_1562,N_316,N_211);
or U1563 (N_1563,N_169,N_796);
or U1564 (N_1564,N_610,N_456);
nor U1565 (N_1565,N_445,N_68);
or U1566 (N_1566,N_965,N_278);
and U1567 (N_1567,N_586,N_3);
nand U1568 (N_1568,N_968,N_460);
nand U1569 (N_1569,N_353,N_952);
nor U1570 (N_1570,N_790,N_74);
or U1571 (N_1571,N_824,N_437);
or U1572 (N_1572,N_473,N_512);
nor U1573 (N_1573,N_707,N_646);
nand U1574 (N_1574,N_409,N_263);
and U1575 (N_1575,N_771,N_835);
and U1576 (N_1576,N_800,N_702);
nand U1577 (N_1577,N_592,N_737);
and U1578 (N_1578,N_747,N_934);
or U1579 (N_1579,N_474,N_509);
nand U1580 (N_1580,N_460,N_149);
or U1581 (N_1581,N_105,N_244);
nor U1582 (N_1582,N_4,N_769);
nand U1583 (N_1583,N_546,N_96);
nor U1584 (N_1584,N_883,N_100);
nand U1585 (N_1585,N_338,N_602);
or U1586 (N_1586,N_713,N_818);
and U1587 (N_1587,N_732,N_461);
or U1588 (N_1588,N_82,N_128);
nor U1589 (N_1589,N_241,N_29);
nor U1590 (N_1590,N_426,N_860);
or U1591 (N_1591,N_743,N_497);
nand U1592 (N_1592,N_333,N_190);
xor U1593 (N_1593,N_103,N_272);
nand U1594 (N_1594,N_246,N_621);
nor U1595 (N_1595,N_986,N_925);
and U1596 (N_1596,N_353,N_551);
and U1597 (N_1597,N_483,N_477);
or U1598 (N_1598,N_977,N_248);
nand U1599 (N_1599,N_719,N_638);
nor U1600 (N_1600,N_837,N_213);
and U1601 (N_1601,N_109,N_117);
nand U1602 (N_1602,N_464,N_356);
or U1603 (N_1603,N_720,N_196);
and U1604 (N_1604,N_452,N_116);
or U1605 (N_1605,N_83,N_224);
or U1606 (N_1606,N_261,N_920);
or U1607 (N_1607,N_89,N_101);
nor U1608 (N_1608,N_517,N_582);
nand U1609 (N_1609,N_676,N_398);
or U1610 (N_1610,N_163,N_455);
nor U1611 (N_1611,N_522,N_13);
nor U1612 (N_1612,N_128,N_579);
or U1613 (N_1613,N_360,N_447);
nor U1614 (N_1614,N_772,N_267);
nor U1615 (N_1615,N_919,N_846);
or U1616 (N_1616,N_858,N_254);
nor U1617 (N_1617,N_970,N_353);
or U1618 (N_1618,N_896,N_642);
nand U1619 (N_1619,N_696,N_881);
and U1620 (N_1620,N_311,N_287);
nand U1621 (N_1621,N_414,N_619);
nand U1622 (N_1622,N_799,N_157);
nor U1623 (N_1623,N_306,N_319);
nand U1624 (N_1624,N_42,N_776);
or U1625 (N_1625,N_363,N_786);
and U1626 (N_1626,N_833,N_404);
and U1627 (N_1627,N_609,N_197);
nor U1628 (N_1628,N_300,N_625);
nand U1629 (N_1629,N_585,N_204);
or U1630 (N_1630,N_184,N_545);
or U1631 (N_1631,N_88,N_924);
or U1632 (N_1632,N_112,N_449);
and U1633 (N_1633,N_901,N_536);
nand U1634 (N_1634,N_439,N_542);
nand U1635 (N_1635,N_346,N_230);
or U1636 (N_1636,N_371,N_659);
or U1637 (N_1637,N_799,N_176);
and U1638 (N_1638,N_6,N_222);
or U1639 (N_1639,N_719,N_854);
or U1640 (N_1640,N_781,N_566);
nand U1641 (N_1641,N_910,N_119);
nor U1642 (N_1642,N_356,N_326);
nand U1643 (N_1643,N_908,N_879);
or U1644 (N_1644,N_472,N_538);
or U1645 (N_1645,N_831,N_431);
nor U1646 (N_1646,N_908,N_102);
nor U1647 (N_1647,N_190,N_587);
nand U1648 (N_1648,N_641,N_149);
and U1649 (N_1649,N_709,N_377);
or U1650 (N_1650,N_845,N_727);
and U1651 (N_1651,N_761,N_950);
or U1652 (N_1652,N_847,N_652);
nand U1653 (N_1653,N_165,N_20);
nor U1654 (N_1654,N_789,N_32);
nor U1655 (N_1655,N_125,N_586);
nand U1656 (N_1656,N_840,N_206);
and U1657 (N_1657,N_250,N_913);
nand U1658 (N_1658,N_919,N_414);
nand U1659 (N_1659,N_849,N_26);
nor U1660 (N_1660,N_606,N_404);
nand U1661 (N_1661,N_924,N_16);
nand U1662 (N_1662,N_715,N_385);
nor U1663 (N_1663,N_867,N_138);
or U1664 (N_1664,N_159,N_873);
nor U1665 (N_1665,N_891,N_360);
nor U1666 (N_1666,N_450,N_432);
nor U1667 (N_1667,N_883,N_862);
or U1668 (N_1668,N_926,N_287);
nand U1669 (N_1669,N_180,N_424);
nor U1670 (N_1670,N_835,N_589);
nand U1671 (N_1671,N_879,N_11);
or U1672 (N_1672,N_856,N_908);
nand U1673 (N_1673,N_120,N_89);
and U1674 (N_1674,N_853,N_94);
or U1675 (N_1675,N_437,N_889);
nand U1676 (N_1676,N_471,N_146);
or U1677 (N_1677,N_515,N_772);
nor U1678 (N_1678,N_993,N_298);
nand U1679 (N_1679,N_439,N_571);
and U1680 (N_1680,N_558,N_403);
and U1681 (N_1681,N_16,N_485);
and U1682 (N_1682,N_685,N_537);
and U1683 (N_1683,N_984,N_772);
nand U1684 (N_1684,N_288,N_109);
nor U1685 (N_1685,N_261,N_403);
nor U1686 (N_1686,N_544,N_165);
nor U1687 (N_1687,N_886,N_355);
nor U1688 (N_1688,N_845,N_463);
or U1689 (N_1689,N_963,N_753);
nand U1690 (N_1690,N_285,N_520);
nor U1691 (N_1691,N_128,N_130);
or U1692 (N_1692,N_392,N_104);
and U1693 (N_1693,N_498,N_399);
nor U1694 (N_1694,N_183,N_512);
or U1695 (N_1695,N_512,N_90);
and U1696 (N_1696,N_850,N_539);
and U1697 (N_1697,N_172,N_548);
nor U1698 (N_1698,N_917,N_187);
nand U1699 (N_1699,N_990,N_180);
or U1700 (N_1700,N_557,N_603);
nor U1701 (N_1701,N_605,N_994);
or U1702 (N_1702,N_129,N_11);
nand U1703 (N_1703,N_371,N_310);
nand U1704 (N_1704,N_404,N_895);
and U1705 (N_1705,N_328,N_805);
or U1706 (N_1706,N_262,N_823);
or U1707 (N_1707,N_11,N_367);
and U1708 (N_1708,N_106,N_661);
and U1709 (N_1709,N_446,N_251);
and U1710 (N_1710,N_159,N_526);
nor U1711 (N_1711,N_200,N_478);
nand U1712 (N_1712,N_177,N_142);
or U1713 (N_1713,N_180,N_547);
nor U1714 (N_1714,N_37,N_996);
nor U1715 (N_1715,N_801,N_452);
nand U1716 (N_1716,N_158,N_244);
and U1717 (N_1717,N_128,N_379);
nor U1718 (N_1718,N_987,N_154);
or U1719 (N_1719,N_110,N_382);
nand U1720 (N_1720,N_360,N_789);
xor U1721 (N_1721,N_674,N_176);
and U1722 (N_1722,N_306,N_713);
or U1723 (N_1723,N_956,N_968);
xnor U1724 (N_1724,N_914,N_830);
nand U1725 (N_1725,N_615,N_784);
nor U1726 (N_1726,N_310,N_793);
nor U1727 (N_1727,N_851,N_134);
and U1728 (N_1728,N_244,N_875);
and U1729 (N_1729,N_556,N_733);
nor U1730 (N_1730,N_164,N_19);
or U1731 (N_1731,N_905,N_351);
and U1732 (N_1732,N_187,N_843);
or U1733 (N_1733,N_412,N_193);
nand U1734 (N_1734,N_781,N_565);
nand U1735 (N_1735,N_307,N_453);
and U1736 (N_1736,N_363,N_388);
nand U1737 (N_1737,N_705,N_46);
or U1738 (N_1738,N_65,N_615);
nand U1739 (N_1739,N_958,N_814);
or U1740 (N_1740,N_320,N_253);
or U1741 (N_1741,N_278,N_393);
and U1742 (N_1742,N_436,N_546);
or U1743 (N_1743,N_379,N_734);
nand U1744 (N_1744,N_270,N_958);
nor U1745 (N_1745,N_392,N_658);
nor U1746 (N_1746,N_744,N_898);
nor U1747 (N_1747,N_79,N_466);
and U1748 (N_1748,N_510,N_790);
and U1749 (N_1749,N_673,N_312);
or U1750 (N_1750,N_604,N_597);
nor U1751 (N_1751,N_55,N_455);
nand U1752 (N_1752,N_569,N_810);
nand U1753 (N_1753,N_170,N_15);
nor U1754 (N_1754,N_58,N_747);
nor U1755 (N_1755,N_75,N_818);
nor U1756 (N_1756,N_960,N_938);
or U1757 (N_1757,N_935,N_103);
nand U1758 (N_1758,N_877,N_966);
and U1759 (N_1759,N_662,N_756);
and U1760 (N_1760,N_921,N_950);
or U1761 (N_1761,N_240,N_960);
and U1762 (N_1762,N_275,N_649);
or U1763 (N_1763,N_596,N_121);
and U1764 (N_1764,N_846,N_787);
and U1765 (N_1765,N_934,N_412);
and U1766 (N_1766,N_691,N_26);
nor U1767 (N_1767,N_698,N_353);
nand U1768 (N_1768,N_102,N_547);
or U1769 (N_1769,N_869,N_527);
and U1770 (N_1770,N_959,N_660);
nand U1771 (N_1771,N_345,N_651);
nand U1772 (N_1772,N_891,N_662);
nand U1773 (N_1773,N_710,N_930);
nor U1774 (N_1774,N_6,N_388);
nor U1775 (N_1775,N_815,N_855);
nor U1776 (N_1776,N_796,N_983);
nand U1777 (N_1777,N_235,N_376);
or U1778 (N_1778,N_27,N_3);
and U1779 (N_1779,N_34,N_77);
and U1780 (N_1780,N_661,N_153);
or U1781 (N_1781,N_46,N_774);
nor U1782 (N_1782,N_988,N_661);
or U1783 (N_1783,N_661,N_248);
nor U1784 (N_1784,N_980,N_90);
and U1785 (N_1785,N_805,N_258);
and U1786 (N_1786,N_64,N_457);
nor U1787 (N_1787,N_680,N_757);
nor U1788 (N_1788,N_182,N_102);
or U1789 (N_1789,N_36,N_783);
nor U1790 (N_1790,N_742,N_29);
or U1791 (N_1791,N_684,N_731);
or U1792 (N_1792,N_866,N_309);
and U1793 (N_1793,N_172,N_663);
and U1794 (N_1794,N_797,N_984);
or U1795 (N_1795,N_679,N_804);
and U1796 (N_1796,N_626,N_221);
nor U1797 (N_1797,N_769,N_737);
nor U1798 (N_1798,N_171,N_778);
and U1799 (N_1799,N_5,N_976);
or U1800 (N_1800,N_156,N_976);
nand U1801 (N_1801,N_839,N_382);
nor U1802 (N_1802,N_671,N_88);
and U1803 (N_1803,N_131,N_184);
nor U1804 (N_1804,N_189,N_27);
xnor U1805 (N_1805,N_197,N_946);
and U1806 (N_1806,N_979,N_422);
nand U1807 (N_1807,N_370,N_287);
and U1808 (N_1808,N_977,N_395);
nor U1809 (N_1809,N_989,N_864);
and U1810 (N_1810,N_172,N_753);
nor U1811 (N_1811,N_65,N_857);
nor U1812 (N_1812,N_580,N_57);
nand U1813 (N_1813,N_945,N_433);
nor U1814 (N_1814,N_760,N_714);
and U1815 (N_1815,N_628,N_812);
nand U1816 (N_1816,N_583,N_971);
and U1817 (N_1817,N_848,N_95);
nand U1818 (N_1818,N_103,N_915);
nand U1819 (N_1819,N_890,N_910);
nand U1820 (N_1820,N_396,N_57);
nand U1821 (N_1821,N_166,N_855);
or U1822 (N_1822,N_23,N_333);
nand U1823 (N_1823,N_236,N_55);
and U1824 (N_1824,N_166,N_844);
nand U1825 (N_1825,N_30,N_299);
nor U1826 (N_1826,N_722,N_362);
nand U1827 (N_1827,N_642,N_505);
and U1828 (N_1828,N_79,N_342);
or U1829 (N_1829,N_378,N_663);
and U1830 (N_1830,N_837,N_452);
or U1831 (N_1831,N_3,N_927);
or U1832 (N_1832,N_311,N_158);
or U1833 (N_1833,N_951,N_799);
nand U1834 (N_1834,N_318,N_964);
nand U1835 (N_1835,N_28,N_385);
nor U1836 (N_1836,N_41,N_317);
and U1837 (N_1837,N_364,N_756);
nor U1838 (N_1838,N_460,N_385);
nor U1839 (N_1839,N_990,N_582);
nand U1840 (N_1840,N_917,N_509);
and U1841 (N_1841,N_361,N_137);
nand U1842 (N_1842,N_456,N_921);
or U1843 (N_1843,N_949,N_774);
nor U1844 (N_1844,N_14,N_904);
nor U1845 (N_1845,N_690,N_881);
or U1846 (N_1846,N_328,N_643);
or U1847 (N_1847,N_29,N_421);
nand U1848 (N_1848,N_808,N_248);
or U1849 (N_1849,N_208,N_506);
and U1850 (N_1850,N_543,N_734);
and U1851 (N_1851,N_455,N_798);
and U1852 (N_1852,N_934,N_645);
and U1853 (N_1853,N_124,N_301);
and U1854 (N_1854,N_888,N_587);
and U1855 (N_1855,N_375,N_508);
and U1856 (N_1856,N_227,N_41);
nand U1857 (N_1857,N_720,N_542);
nand U1858 (N_1858,N_589,N_676);
nand U1859 (N_1859,N_466,N_605);
nor U1860 (N_1860,N_350,N_674);
nand U1861 (N_1861,N_709,N_80);
and U1862 (N_1862,N_138,N_845);
or U1863 (N_1863,N_59,N_854);
and U1864 (N_1864,N_931,N_366);
or U1865 (N_1865,N_836,N_657);
nor U1866 (N_1866,N_341,N_425);
or U1867 (N_1867,N_441,N_37);
and U1868 (N_1868,N_368,N_141);
nand U1869 (N_1869,N_935,N_392);
nor U1870 (N_1870,N_926,N_644);
or U1871 (N_1871,N_817,N_478);
and U1872 (N_1872,N_936,N_631);
xnor U1873 (N_1873,N_882,N_816);
nand U1874 (N_1874,N_299,N_892);
nand U1875 (N_1875,N_304,N_649);
or U1876 (N_1876,N_704,N_593);
and U1877 (N_1877,N_909,N_666);
or U1878 (N_1878,N_928,N_769);
nor U1879 (N_1879,N_109,N_227);
or U1880 (N_1880,N_421,N_53);
nor U1881 (N_1881,N_327,N_330);
and U1882 (N_1882,N_15,N_434);
or U1883 (N_1883,N_407,N_34);
and U1884 (N_1884,N_405,N_62);
nor U1885 (N_1885,N_579,N_73);
nand U1886 (N_1886,N_167,N_846);
and U1887 (N_1887,N_0,N_781);
and U1888 (N_1888,N_322,N_532);
and U1889 (N_1889,N_546,N_867);
or U1890 (N_1890,N_450,N_989);
and U1891 (N_1891,N_470,N_955);
or U1892 (N_1892,N_351,N_811);
nand U1893 (N_1893,N_598,N_300);
and U1894 (N_1894,N_591,N_116);
or U1895 (N_1895,N_415,N_514);
nand U1896 (N_1896,N_190,N_411);
nor U1897 (N_1897,N_776,N_26);
or U1898 (N_1898,N_475,N_30);
or U1899 (N_1899,N_513,N_791);
or U1900 (N_1900,N_168,N_995);
or U1901 (N_1901,N_478,N_110);
and U1902 (N_1902,N_292,N_403);
nand U1903 (N_1903,N_58,N_191);
nor U1904 (N_1904,N_964,N_570);
nor U1905 (N_1905,N_18,N_864);
and U1906 (N_1906,N_275,N_53);
nand U1907 (N_1907,N_366,N_709);
nand U1908 (N_1908,N_788,N_193);
nor U1909 (N_1909,N_612,N_399);
and U1910 (N_1910,N_678,N_474);
or U1911 (N_1911,N_128,N_195);
and U1912 (N_1912,N_266,N_639);
nand U1913 (N_1913,N_810,N_417);
nor U1914 (N_1914,N_650,N_866);
and U1915 (N_1915,N_979,N_373);
and U1916 (N_1916,N_358,N_413);
or U1917 (N_1917,N_246,N_659);
or U1918 (N_1918,N_571,N_978);
and U1919 (N_1919,N_138,N_730);
nor U1920 (N_1920,N_593,N_33);
nor U1921 (N_1921,N_285,N_670);
and U1922 (N_1922,N_139,N_59);
nand U1923 (N_1923,N_405,N_517);
and U1924 (N_1924,N_272,N_89);
nor U1925 (N_1925,N_75,N_921);
and U1926 (N_1926,N_451,N_482);
or U1927 (N_1927,N_867,N_896);
or U1928 (N_1928,N_317,N_16);
or U1929 (N_1929,N_966,N_621);
nor U1930 (N_1930,N_523,N_662);
nand U1931 (N_1931,N_259,N_916);
or U1932 (N_1932,N_330,N_186);
nand U1933 (N_1933,N_182,N_933);
nand U1934 (N_1934,N_758,N_690);
nor U1935 (N_1935,N_377,N_505);
nand U1936 (N_1936,N_302,N_23);
or U1937 (N_1937,N_325,N_902);
nand U1938 (N_1938,N_526,N_942);
or U1939 (N_1939,N_513,N_658);
and U1940 (N_1940,N_122,N_959);
nand U1941 (N_1941,N_974,N_726);
nand U1942 (N_1942,N_848,N_176);
and U1943 (N_1943,N_182,N_573);
or U1944 (N_1944,N_48,N_561);
and U1945 (N_1945,N_908,N_661);
nand U1946 (N_1946,N_901,N_877);
nand U1947 (N_1947,N_160,N_490);
nor U1948 (N_1948,N_866,N_233);
nand U1949 (N_1949,N_651,N_448);
nand U1950 (N_1950,N_901,N_807);
nand U1951 (N_1951,N_748,N_572);
or U1952 (N_1952,N_141,N_21);
nand U1953 (N_1953,N_203,N_128);
or U1954 (N_1954,N_333,N_945);
and U1955 (N_1955,N_671,N_514);
or U1956 (N_1956,N_882,N_86);
nand U1957 (N_1957,N_771,N_909);
or U1958 (N_1958,N_588,N_507);
nand U1959 (N_1959,N_488,N_379);
nor U1960 (N_1960,N_850,N_684);
nand U1961 (N_1961,N_373,N_133);
nand U1962 (N_1962,N_909,N_983);
or U1963 (N_1963,N_223,N_104);
nor U1964 (N_1964,N_204,N_375);
nor U1965 (N_1965,N_808,N_547);
and U1966 (N_1966,N_814,N_708);
or U1967 (N_1967,N_684,N_688);
or U1968 (N_1968,N_105,N_368);
or U1969 (N_1969,N_500,N_35);
nor U1970 (N_1970,N_520,N_971);
nand U1971 (N_1971,N_63,N_319);
and U1972 (N_1972,N_660,N_911);
or U1973 (N_1973,N_259,N_604);
and U1974 (N_1974,N_20,N_461);
nor U1975 (N_1975,N_996,N_691);
or U1976 (N_1976,N_575,N_789);
or U1977 (N_1977,N_106,N_361);
and U1978 (N_1978,N_208,N_765);
nand U1979 (N_1979,N_673,N_37);
and U1980 (N_1980,N_613,N_676);
and U1981 (N_1981,N_18,N_9);
or U1982 (N_1982,N_196,N_622);
and U1983 (N_1983,N_608,N_456);
or U1984 (N_1984,N_414,N_786);
or U1985 (N_1985,N_607,N_62);
and U1986 (N_1986,N_981,N_304);
or U1987 (N_1987,N_555,N_773);
nor U1988 (N_1988,N_754,N_701);
and U1989 (N_1989,N_242,N_266);
nor U1990 (N_1990,N_925,N_48);
or U1991 (N_1991,N_232,N_571);
or U1992 (N_1992,N_442,N_71);
and U1993 (N_1993,N_405,N_33);
or U1994 (N_1994,N_378,N_576);
nor U1995 (N_1995,N_772,N_860);
nor U1996 (N_1996,N_51,N_586);
nor U1997 (N_1997,N_389,N_749);
nor U1998 (N_1998,N_501,N_754);
nor U1999 (N_1999,N_774,N_47);
or U2000 (N_2000,N_1306,N_1452);
nand U2001 (N_2001,N_1982,N_1495);
nand U2002 (N_2002,N_1110,N_1261);
or U2003 (N_2003,N_1672,N_1044);
nor U2004 (N_2004,N_1830,N_1393);
nor U2005 (N_2005,N_1757,N_1781);
or U2006 (N_2006,N_1161,N_1555);
nor U2007 (N_2007,N_1285,N_1947);
nand U2008 (N_2008,N_1405,N_1398);
nand U2009 (N_2009,N_1800,N_1963);
nor U2010 (N_2010,N_1547,N_1014);
nand U2011 (N_2011,N_1116,N_1584);
nor U2012 (N_2012,N_1346,N_1128);
nand U2013 (N_2013,N_1862,N_1323);
and U2014 (N_2014,N_1365,N_1904);
and U2015 (N_2015,N_1391,N_1666);
nor U2016 (N_2016,N_1430,N_1386);
nor U2017 (N_2017,N_1630,N_1651);
or U2018 (N_2018,N_1887,N_1321);
nor U2019 (N_2019,N_1929,N_1154);
nor U2020 (N_2020,N_1156,N_1092);
and U2021 (N_2021,N_1545,N_1582);
and U2022 (N_2022,N_1200,N_1373);
nand U2023 (N_2023,N_1871,N_1911);
nor U2024 (N_2024,N_1277,N_1780);
nor U2025 (N_2025,N_1629,N_1111);
and U2026 (N_2026,N_1708,N_1475);
xor U2027 (N_2027,N_1662,N_1791);
nor U2028 (N_2028,N_1675,N_1444);
and U2029 (N_2029,N_1951,N_1600);
nor U2030 (N_2030,N_1889,N_1726);
or U2031 (N_2031,N_1442,N_1840);
nand U2032 (N_2032,N_1440,N_1741);
nand U2033 (N_2033,N_1981,N_1308);
or U2034 (N_2034,N_1097,N_1687);
nand U2035 (N_2035,N_1934,N_1139);
nand U2036 (N_2036,N_1160,N_1715);
and U2037 (N_2037,N_1855,N_1586);
or U2038 (N_2038,N_1606,N_1641);
and U2039 (N_2039,N_1618,N_1478);
or U2040 (N_2040,N_1621,N_1607);
nor U2041 (N_2041,N_1048,N_1267);
nor U2042 (N_2042,N_1260,N_1471);
nor U2043 (N_2043,N_1583,N_1140);
or U2044 (N_2044,N_1221,N_1297);
and U2045 (N_2045,N_1252,N_1512);
nor U2046 (N_2046,N_1249,N_1222);
and U2047 (N_2047,N_1322,N_1098);
and U2048 (N_2048,N_1157,N_1822);
nor U2049 (N_2049,N_1169,N_1223);
nand U2050 (N_2050,N_1113,N_1719);
nor U2051 (N_2051,N_1553,N_1100);
nand U2052 (N_2052,N_1036,N_1681);
nand U2053 (N_2053,N_1387,N_1885);
and U2054 (N_2054,N_1886,N_1109);
and U2055 (N_2055,N_1955,N_1538);
or U2056 (N_2056,N_1534,N_1419);
nor U2057 (N_2057,N_1435,N_1890);
nand U2058 (N_2058,N_1552,N_1505);
nor U2059 (N_2059,N_1711,N_1759);
and U2060 (N_2060,N_1670,N_1774);
or U2061 (N_2061,N_1500,N_1604);
and U2062 (N_2062,N_1399,N_1043);
and U2063 (N_2063,N_1273,N_1596);
or U2064 (N_2064,N_1357,N_1038);
nand U2065 (N_2065,N_1228,N_1377);
or U2066 (N_2066,N_1164,N_1404);
nand U2067 (N_2067,N_1674,N_1354);
and U2068 (N_2068,N_1022,N_1465);
or U2069 (N_2069,N_1577,N_1546);
or U2070 (N_2070,N_1779,N_1931);
nor U2071 (N_2071,N_1028,N_1507);
nand U2072 (N_2072,N_1216,N_1806);
and U2073 (N_2073,N_1016,N_1150);
nand U2074 (N_2074,N_1688,N_1698);
nand U2075 (N_2075,N_1166,N_1334);
nand U2076 (N_2076,N_1634,N_1343);
or U2077 (N_2077,N_1530,N_1006);
nor U2078 (N_2078,N_1335,N_1163);
or U2079 (N_2079,N_1747,N_1299);
nand U2080 (N_2080,N_1699,N_1665);
nand U2081 (N_2081,N_1753,N_1650);
or U2082 (N_2082,N_1589,N_1197);
or U2083 (N_2083,N_1230,N_1782);
or U2084 (N_2084,N_1259,N_1085);
or U2085 (N_2085,N_1420,N_1272);
nor U2086 (N_2086,N_1498,N_1455);
and U2087 (N_2087,N_1513,N_1107);
and U2088 (N_2088,N_1412,N_1418);
nand U2089 (N_2089,N_1917,N_1953);
and U2090 (N_2090,N_1176,N_1434);
and U2091 (N_2091,N_1787,N_1338);
or U2092 (N_2092,N_1183,N_1985);
or U2093 (N_2093,N_1049,N_1879);
nor U2094 (N_2094,N_1668,N_1397);
or U2095 (N_2095,N_1853,N_1810);
xnor U2096 (N_2096,N_1793,N_1180);
nand U2097 (N_2097,N_1777,N_1842);
nand U2098 (N_2098,N_1439,N_1579);
nand U2099 (N_2099,N_1511,N_1250);
nor U2100 (N_2100,N_1986,N_1202);
or U2101 (N_2101,N_1739,N_1123);
and U2102 (N_2102,N_1358,N_1380);
and U2103 (N_2103,N_1214,N_1704);
nand U2104 (N_2104,N_1271,N_1570);
or U2105 (N_2105,N_1317,N_1523);
nand U2106 (N_2106,N_1926,N_1432);
nand U2107 (N_2107,N_1789,N_1104);
nor U2108 (N_2108,N_1746,N_1030);
nand U2109 (N_2109,N_1479,N_1900);
and U2110 (N_2110,N_1848,N_1903);
nand U2111 (N_2111,N_1188,N_1775);
or U2112 (N_2112,N_1408,N_1256);
or U2113 (N_2113,N_1120,N_1590);
nand U2114 (N_2114,N_1952,N_1496);
nand U2115 (N_2115,N_1155,N_1783);
nand U2116 (N_2116,N_1730,N_1227);
or U2117 (N_2117,N_1005,N_1413);
and U2118 (N_2118,N_1248,N_1244);
xnor U2119 (N_2119,N_1426,N_1633);
nor U2120 (N_2120,N_1979,N_1300);
or U2121 (N_2121,N_1385,N_1959);
nor U2122 (N_2122,N_1018,N_1205);
or U2123 (N_2123,N_1563,N_1126);
and U2124 (N_2124,N_1697,N_1204);
and U2125 (N_2125,N_1501,N_1178);
nand U2126 (N_2126,N_1960,N_1499);
nor U2127 (N_2127,N_1165,N_1694);
nor U2128 (N_2128,N_1593,N_1443);
nand U2129 (N_2129,N_1752,N_1020);
nor U2130 (N_2130,N_1910,N_1191);
xor U2131 (N_2131,N_1012,N_1770);
nand U2132 (N_2132,N_1280,N_1972);
nor U2133 (N_2133,N_1026,N_1517);
nor U2134 (N_2134,N_1591,N_1146);
and U2135 (N_2135,N_1624,N_1870);
or U2136 (N_2136,N_1655,N_1893);
or U2137 (N_2137,N_1002,N_1211);
or U2138 (N_2138,N_1461,N_1967);
nor U2139 (N_2139,N_1134,N_1502);
nor U2140 (N_2140,N_1874,N_1971);
nand U2141 (N_2141,N_1376,N_1785);
or U2142 (N_2142,N_1429,N_1945);
nand U2143 (N_2143,N_1623,N_1878);
and U2144 (N_2144,N_1587,N_1859);
nor U2145 (N_2145,N_1406,N_1756);
nand U2146 (N_2146,N_1595,N_1922);
nand U2147 (N_2147,N_1218,N_1663);
xnor U2148 (N_2148,N_1340,N_1573);
nand U2149 (N_2149,N_1283,N_1556);
nand U2150 (N_2150,N_1061,N_1436);
nand U2151 (N_2151,N_1091,N_1686);
nand U2152 (N_2152,N_1700,N_1896);
or U2153 (N_2153,N_1867,N_1152);
and U2154 (N_2154,N_1836,N_1074);
and U2155 (N_2155,N_1433,N_1720);
and U2156 (N_2156,N_1743,N_1640);
or U2157 (N_2157,N_1309,N_1009);
or U2158 (N_2158,N_1243,N_1918);
or U2159 (N_2159,N_1549,N_1866);
nand U2160 (N_2160,N_1923,N_1013);
or U2161 (N_2161,N_1410,N_1987);
nand U2162 (N_2162,N_1384,N_1213);
and U2163 (N_2163,N_1275,N_1325);
nand U2164 (N_2164,N_1937,N_1816);
nand U2165 (N_2165,N_1734,N_1835);
and U2166 (N_2166,N_1186,N_1291);
nor U2167 (N_2167,N_1751,N_1264);
or U2168 (N_2168,N_1510,N_1516);
nor U2169 (N_2169,N_1033,N_1854);
nand U2170 (N_2170,N_1492,N_1310);
or U2171 (N_2171,N_1246,N_1737);
or U2172 (N_2172,N_1560,N_1333);
nand U2173 (N_2173,N_1316,N_1899);
nand U2174 (N_2174,N_1869,N_1023);
or U2175 (N_2175,N_1490,N_1010);
nor U2176 (N_2176,N_1326,N_1695);
and U2177 (N_2177,N_1997,N_1425);
nand U2178 (N_2178,N_1802,N_1941);
and U2179 (N_2179,N_1056,N_1193);
nand U2180 (N_2180,N_1265,N_1276);
and U2181 (N_2181,N_1301,N_1628);
nor U2182 (N_2182,N_1144,N_1701);
nand U2183 (N_2183,N_1850,N_1807);
or U2184 (N_2184,N_1046,N_1201);
nand U2185 (N_2185,N_1281,N_1849);
or U2186 (N_2186,N_1231,N_1619);
or U2187 (N_2187,N_1474,N_1122);
nor U2188 (N_2188,N_1920,N_1151);
nor U2189 (N_2189,N_1808,N_1684);
nand U2190 (N_2190,N_1347,N_1915);
and U2191 (N_2191,N_1395,N_1718);
or U2192 (N_2192,N_1551,N_1564);
or U2193 (N_2193,N_1838,N_1084);
nand U2194 (N_2194,N_1532,N_1247);
or U2195 (N_2195,N_1565,N_1124);
nor U2196 (N_2196,N_1571,N_1764);
nand U2197 (N_2197,N_1368,N_1677);
and U2198 (N_2198,N_1060,N_1153);
nand U2199 (N_2199,N_1379,N_1921);
or U2200 (N_2200,N_1554,N_1860);
or U2201 (N_2201,N_1678,N_1314);
nand U2202 (N_2202,N_1821,N_1237);
or U2203 (N_2203,N_1488,N_1792);
nor U2204 (N_2204,N_1531,N_1270);
and U2205 (N_2205,N_1927,N_1045);
and U2206 (N_2206,N_1833,N_1302);
nand U2207 (N_2207,N_1936,N_1646);
and U2208 (N_2208,N_1143,N_1788);
or U2209 (N_2209,N_1503,N_1361);
nor U2210 (N_2210,N_1664,N_1882);
or U2211 (N_2211,N_1401,N_1293);
and U2212 (N_2212,N_1990,N_1796);
or U2213 (N_2213,N_1631,N_1818);
or U2214 (N_2214,N_1279,N_1642);
nand U2215 (N_2215,N_1212,N_1598);
nand U2216 (N_2216,N_1238,N_1491);
or U2217 (N_2217,N_1957,N_1173);
and U2218 (N_2218,N_1978,N_1636);
nor U2219 (N_2219,N_1182,N_1776);
nor U2220 (N_2220,N_1627,N_1327);
nor U2221 (N_2221,N_1892,N_1797);
nand U2222 (N_2222,N_1011,N_1041);
nor U2223 (N_2223,N_1313,N_1129);
nand U2224 (N_2224,N_1992,N_1864);
nor U2225 (N_2225,N_1245,N_1812);
and U2226 (N_2226,N_1181,N_1605);
and U2227 (N_2227,N_1127,N_1360);
nor U2228 (N_2228,N_1572,N_1263);
nor U2229 (N_2229,N_1266,N_1177);
and U2230 (N_2230,N_1476,N_1149);
nor U2231 (N_2231,N_1965,N_1856);
nand U2232 (N_2232,N_1255,N_1328);
xor U2233 (N_2233,N_1620,N_1034);
or U2234 (N_2234,N_1844,N_1529);
and U2235 (N_2235,N_1518,N_1112);
nor U2236 (N_2236,N_1374,N_1485);
nand U2237 (N_2237,N_1196,N_1162);
and U2238 (N_2238,N_1147,N_1449);
or U2239 (N_2239,N_1611,N_1094);
nand U2240 (N_2240,N_1875,N_1993);
and U2241 (N_2241,N_1745,N_1135);
nand U2242 (N_2242,N_1712,N_1241);
or U2243 (N_2243,N_1451,N_1072);
nor U2244 (N_2244,N_1407,N_1829);
nand U2245 (N_2245,N_1103,N_1969);
and U2246 (N_2246,N_1114,N_1190);
and U2247 (N_2247,N_1909,N_1690);
or U2248 (N_2248,N_1613,N_1561);
or U2249 (N_2249,N_1716,N_1970);
or U2250 (N_2250,N_1071,N_1661);
or U2251 (N_2251,N_1880,N_1159);
and U2252 (N_2252,N_1839,N_1567);
nor U2253 (N_2253,N_1576,N_1585);
and U2254 (N_2254,N_1400,N_1390);
or U2255 (N_2255,N_1544,N_1671);
nor U2256 (N_2256,N_1363,N_1075);
or U2257 (N_2257,N_1095,N_1076);
and U2258 (N_2258,N_1602,N_1610);
nand U2259 (N_2259,N_1954,N_1765);
nor U2260 (N_2260,N_1804,N_1138);
or U2261 (N_2261,N_1943,N_1846);
nand U2262 (N_2262,N_1388,N_1722);
and U2263 (N_2263,N_1481,N_1203);
and U2264 (N_2264,N_1657,N_1115);
nor U2265 (N_2265,N_1320,N_1515);
or U2266 (N_2266,N_1438,N_1251);
nor U2267 (N_2267,N_1268,N_1240);
nand U2268 (N_2268,N_1070,N_1446);
and U2269 (N_2269,N_1437,N_1784);
nor U2270 (N_2270,N_1614,N_1187);
nor U2271 (N_2271,N_1557,N_1232);
nor U2272 (N_2272,N_1928,N_1145);
and U2273 (N_2273,N_1578,N_1933);
or U2274 (N_2274,N_1815,N_1996);
and U2275 (N_2275,N_1524,N_1742);
nor U2276 (N_2276,N_1318,N_1845);
or U2277 (N_2277,N_1458,N_1089);
nand U2278 (N_2278,N_1102,N_1950);
nand U2279 (N_2279,N_1622,N_1643);
and U2280 (N_2280,N_1736,N_1814);
nor U2281 (N_2281,N_1226,N_1142);
nor U2282 (N_2282,N_1654,N_1351);
or U2283 (N_2283,N_1210,N_1052);
nor U2284 (N_2284,N_1339,N_1031);
nand U2285 (N_2285,N_1108,N_1858);
and U2286 (N_2286,N_1863,N_1888);
or U2287 (N_2287,N_1079,N_1966);
xnor U2288 (N_2288,N_1964,N_1637);
and U2289 (N_2289,N_1184,N_1274);
nand U2290 (N_2290,N_1758,N_1315);
or U2291 (N_2291,N_1375,N_1771);
nor U2292 (N_2292,N_1396,N_1409);
nand U2293 (N_2293,N_1527,N_1378);
nor U2294 (N_2294,N_1902,N_1287);
or U2295 (N_2295,N_1065,N_1001);
nand U2296 (N_2296,N_1514,N_1239);
nand U2297 (N_2297,N_1486,N_1944);
or U2298 (N_2298,N_1068,N_1424);
nor U2299 (N_2299,N_1235,N_1463);
nand U2300 (N_2300,N_1289,N_1801);
nor U2301 (N_2301,N_1344,N_1137);
and U2302 (N_2302,N_1055,N_1760);
nand U2303 (N_2303,N_1508,N_1447);
and U2304 (N_2304,N_1148,N_1336);
or U2305 (N_2305,N_1961,N_1962);
nor U2306 (N_2306,N_1819,N_1541);
and U2307 (N_2307,N_1766,N_1868);
or U2308 (N_2308,N_1087,N_1362);
or U2309 (N_2309,N_1861,N_1989);
nor U2310 (N_2310,N_1581,N_1949);
and U2311 (N_2311,N_1660,N_1367);
nor U2312 (N_2312,N_1653,N_1894);
or U2313 (N_2313,N_1004,N_1473);
nand U2314 (N_2314,N_1025,N_1521);
nand U2315 (N_2315,N_1170,N_1345);
and U2316 (N_2316,N_1422,N_1062);
and U2317 (N_2317,N_1017,N_1286);
or U2318 (N_2318,N_1769,N_1296);
and U2319 (N_2319,N_1003,N_1415);
or U2320 (N_2320,N_1035,N_1257);
or U2321 (N_2321,N_1575,N_1450);
nand U2322 (N_2322,N_1469,N_1905);
nand U2323 (N_2323,N_1939,N_1298);
and U2324 (N_2324,N_1872,N_1324);
nor U2325 (N_2325,N_1847,N_1828);
or U2326 (N_2326,N_1794,N_1913);
or U2327 (N_2327,N_1428,N_1168);
nand U2328 (N_2328,N_1976,N_1656);
and U2329 (N_2329,N_1948,N_1768);
and U2330 (N_2330,N_1738,N_1487);
nor U2331 (N_2331,N_1883,N_1403);
or U2332 (N_2332,N_1703,N_1394);
xor U2333 (N_2333,N_1938,N_1562);
nand U2334 (N_2334,N_1483,N_1494);
and U2335 (N_2335,N_1907,N_1891);
and U2336 (N_2336,N_1550,N_1799);
or U2337 (N_2337,N_1983,N_1192);
nand U2338 (N_2338,N_1064,N_1369);
and U2339 (N_2339,N_1647,N_1175);
and U2340 (N_2340,N_1691,N_1710);
nor U2341 (N_2341,N_1057,N_1229);
nand U2342 (N_2342,N_1749,N_1356);
nor U2343 (N_2343,N_1713,N_1884);
nor U2344 (N_2344,N_1083,N_1852);
nor U2345 (N_2345,N_1919,N_1912);
or U2346 (N_2346,N_1209,N_1171);
and U2347 (N_2347,N_1615,N_1994);
nand U2348 (N_2348,N_1592,N_1402);
nor U2349 (N_2349,N_1727,N_1658);
or U2350 (N_2350,N_1980,N_1027);
and U2351 (N_2351,N_1762,N_1597);
nor U2352 (N_2352,N_1709,N_1382);
and U2353 (N_2353,N_1877,N_1609);
nand U2354 (N_2354,N_1925,N_1522);
nand U2355 (N_2355,N_1294,N_1811);
or U2356 (N_2356,N_1370,N_1714);
nor U2357 (N_2357,N_1608,N_1189);
nor U2358 (N_2358,N_1895,N_1568);
or U2359 (N_2359,N_1693,N_1696);
or U2360 (N_2360,N_1303,N_1705);
nor U2361 (N_2361,N_1548,N_1208);
nor U2362 (N_2362,N_1755,N_1132);
nand U2363 (N_2363,N_1644,N_1988);
nor U2364 (N_2364,N_1763,N_1706);
and U2365 (N_2365,N_1118,N_1652);
and U2366 (N_2366,N_1873,N_1566);
or U2367 (N_2367,N_1106,N_1051);
or U2368 (N_2368,N_1638,N_1411);
nand U2369 (N_2369,N_1054,N_1509);
nor U2370 (N_2370,N_1778,N_1185);
and U2371 (N_2371,N_1635,N_1625);
and U2372 (N_2372,N_1050,N_1198);
nand U2373 (N_2373,N_1464,N_1117);
nor U2374 (N_2374,N_1359,N_1790);
or U2375 (N_2375,N_1282,N_1832);
nor U2376 (N_2376,N_1342,N_1195);
nand U2377 (N_2377,N_1825,N_1649);
and U2378 (N_2378,N_1729,N_1467);
nand U2379 (N_2379,N_1682,N_1685);
or U2380 (N_2380,N_1307,N_1817);
nor U2381 (N_2381,N_1723,N_1372);
or U2382 (N_2382,N_1717,N_1105);
or U2383 (N_2383,N_1133,N_1416);
nand U2384 (N_2384,N_1823,N_1857);
nor U2385 (N_2385,N_1136,N_1220);
and U2386 (N_2386,N_1067,N_1000);
nand U2387 (N_2387,N_1468,N_1813);
and U2388 (N_2388,N_1242,N_1805);
and U2389 (N_2389,N_1998,N_1352);
nand U2390 (N_2390,N_1506,N_1841);
or U2391 (N_2391,N_1466,N_1667);
or U2392 (N_2392,N_1225,N_1482);
and U2393 (N_2393,N_1066,N_1459);
and U2394 (N_2394,N_1594,N_1906);
or U2395 (N_2395,N_1088,N_1311);
and U2396 (N_2396,N_1974,N_1269);
nor U2397 (N_2397,N_1292,N_1968);
and U2398 (N_2398,N_1381,N_1441);
nand U2399 (N_2399,N_1304,N_1528);
nand U2400 (N_2400,N_1984,N_1047);
or U2401 (N_2401,N_1707,N_1588);
and U2402 (N_2402,N_1574,N_1824);
nand U2403 (N_2403,N_1331,N_1253);
and U2404 (N_2404,N_1167,N_1460);
and U2405 (N_2405,N_1119,N_1341);
nand U2406 (N_2406,N_1725,N_1721);
or U2407 (N_2407,N_1999,N_1207);
or U2408 (N_2408,N_1470,N_1520);
nand U2409 (N_2409,N_1078,N_1535);
or U2410 (N_2410,N_1007,N_1234);
or U2411 (N_2411,N_1093,N_1932);
and U2412 (N_2412,N_1366,N_1090);
nand U2413 (N_2413,N_1786,N_1820);
or U2414 (N_2414,N_1924,N_1462);
and U2415 (N_2415,N_1617,N_1616);
and U2416 (N_2416,N_1015,N_1099);
nor U2417 (N_2417,N_1851,N_1612);
nand U2418 (N_2418,N_1121,N_1991);
and U2419 (N_2419,N_1073,N_1526);
nor U2420 (N_2420,N_1632,N_1233);
nand U2421 (N_2421,N_1539,N_1329);
nand U2422 (N_2422,N_1278,N_1946);
nor U2423 (N_2423,N_1645,N_1683);
or U2424 (N_2424,N_1081,N_1053);
nor U2425 (N_2425,N_1740,N_1457);
and U2426 (N_2426,N_1733,N_1542);
or U2427 (N_2427,N_1454,N_1383);
xnor U2428 (N_2428,N_1477,N_1558);
or U2429 (N_2429,N_1559,N_1897);
nor U2430 (N_2430,N_1731,N_1975);
and U2431 (N_2431,N_1021,N_1037);
and U2432 (N_2432,N_1956,N_1773);
or U2433 (N_2433,N_1199,N_1421);
nand U2434 (N_2434,N_1332,N_1069);
nor U2435 (N_2435,N_1826,N_1364);
nand U2436 (N_2436,N_1427,N_1930);
nand U2437 (N_2437,N_1809,N_1024);
nand U2438 (N_2438,N_1803,N_1330);
nor U2439 (N_2439,N_1569,N_1973);
nand U2440 (N_2440,N_1679,N_1543);
nor U2441 (N_2441,N_1288,N_1217);
nand U2442 (N_2442,N_1445,N_1580);
and U2443 (N_2443,N_1676,N_1353);
and U2444 (N_2444,N_1337,N_1995);
nand U2445 (N_2445,N_1032,N_1754);
nand U2446 (N_2446,N_1172,N_1837);
or U2447 (N_2447,N_1101,N_1914);
or U2448 (N_2448,N_1086,N_1659);
and U2449 (N_2449,N_1448,N_1371);
nand U2450 (N_2450,N_1493,N_1236);
nand U2451 (N_2451,N_1349,N_1131);
xnor U2452 (N_2452,N_1312,N_1348);
nor U2453 (N_2453,N_1431,N_1540);
or U2454 (N_2454,N_1603,N_1601);
nand U2455 (N_2455,N_1673,N_1519);
nor U2456 (N_2456,N_1876,N_1077);
or U2457 (N_2457,N_1772,N_1831);
or U2458 (N_2458,N_1898,N_1039);
nand U2459 (N_2459,N_1798,N_1881);
nor U2460 (N_2460,N_1305,N_1724);
and U2461 (N_2461,N_1525,N_1497);
nand U2462 (N_2462,N_1748,N_1319);
and U2463 (N_2463,N_1744,N_1179);
and U2464 (N_2464,N_1626,N_1082);
and U2465 (N_2465,N_1295,N_1504);
nor U2466 (N_2466,N_1489,N_1008);
nor U2467 (N_2467,N_1834,N_1692);
nor U2468 (N_2468,N_1843,N_1141);
nand U2469 (N_2469,N_1019,N_1029);
nor U2470 (N_2470,N_1480,N_1537);
nor U2471 (N_2471,N_1689,N_1865);
nor U2472 (N_2472,N_1827,N_1219);
or U2473 (N_2473,N_1669,N_1215);
nor U2474 (N_2474,N_1206,N_1290);
or U2475 (N_2475,N_1639,N_1767);
and U2476 (N_2476,N_1958,N_1472);
nand U2477 (N_2477,N_1063,N_1908);
or U2478 (N_2478,N_1735,N_1350);
nor U2479 (N_2479,N_1262,N_1456);
nand U2480 (N_2480,N_1599,N_1058);
nor U2481 (N_2481,N_1977,N_1059);
or U2482 (N_2482,N_1392,N_1750);
nand U2483 (N_2483,N_1680,N_1732);
nand U2484 (N_2484,N_1158,N_1258);
or U2485 (N_2485,N_1942,N_1423);
and U2486 (N_2486,N_1355,N_1130);
or U2487 (N_2487,N_1453,N_1096);
or U2488 (N_2488,N_1901,N_1080);
and U2489 (N_2489,N_1040,N_1935);
nor U2490 (N_2490,N_1042,N_1414);
nand U2491 (N_2491,N_1174,N_1417);
nand U2492 (N_2492,N_1916,N_1940);
or U2493 (N_2493,N_1533,N_1389);
or U2494 (N_2494,N_1702,N_1284);
nand U2495 (N_2495,N_1194,N_1648);
or U2496 (N_2496,N_1795,N_1254);
or U2497 (N_2497,N_1761,N_1728);
nor U2498 (N_2498,N_1224,N_1125);
and U2499 (N_2499,N_1536,N_1484);
or U2500 (N_2500,N_1434,N_1386);
nand U2501 (N_2501,N_1276,N_1322);
or U2502 (N_2502,N_1390,N_1075);
and U2503 (N_2503,N_1221,N_1742);
and U2504 (N_2504,N_1230,N_1086);
nand U2505 (N_2505,N_1873,N_1206);
and U2506 (N_2506,N_1397,N_1252);
or U2507 (N_2507,N_1758,N_1483);
nor U2508 (N_2508,N_1401,N_1124);
nand U2509 (N_2509,N_1118,N_1847);
nor U2510 (N_2510,N_1608,N_1656);
nor U2511 (N_2511,N_1814,N_1073);
nor U2512 (N_2512,N_1495,N_1171);
nor U2513 (N_2513,N_1391,N_1406);
or U2514 (N_2514,N_1241,N_1706);
nand U2515 (N_2515,N_1980,N_1438);
nor U2516 (N_2516,N_1051,N_1668);
nor U2517 (N_2517,N_1798,N_1841);
or U2518 (N_2518,N_1411,N_1539);
or U2519 (N_2519,N_1267,N_1960);
or U2520 (N_2520,N_1911,N_1245);
nor U2521 (N_2521,N_1471,N_1520);
nor U2522 (N_2522,N_1339,N_1534);
nand U2523 (N_2523,N_1565,N_1748);
nor U2524 (N_2524,N_1979,N_1146);
or U2525 (N_2525,N_1884,N_1936);
and U2526 (N_2526,N_1151,N_1528);
or U2527 (N_2527,N_1299,N_1520);
nor U2528 (N_2528,N_1026,N_1915);
or U2529 (N_2529,N_1074,N_1843);
or U2530 (N_2530,N_1223,N_1378);
nor U2531 (N_2531,N_1207,N_1901);
nand U2532 (N_2532,N_1279,N_1245);
or U2533 (N_2533,N_1538,N_1843);
nor U2534 (N_2534,N_1044,N_1564);
and U2535 (N_2535,N_1868,N_1395);
and U2536 (N_2536,N_1284,N_1184);
and U2537 (N_2537,N_1384,N_1625);
or U2538 (N_2538,N_1719,N_1967);
or U2539 (N_2539,N_1354,N_1849);
nand U2540 (N_2540,N_1836,N_1585);
or U2541 (N_2541,N_1081,N_1918);
nor U2542 (N_2542,N_1465,N_1090);
xnor U2543 (N_2543,N_1197,N_1894);
nor U2544 (N_2544,N_1713,N_1559);
nor U2545 (N_2545,N_1399,N_1967);
or U2546 (N_2546,N_1019,N_1796);
nand U2547 (N_2547,N_1915,N_1961);
nor U2548 (N_2548,N_1505,N_1363);
or U2549 (N_2549,N_1524,N_1068);
nand U2550 (N_2550,N_1595,N_1477);
nor U2551 (N_2551,N_1315,N_1734);
or U2552 (N_2552,N_1583,N_1997);
or U2553 (N_2553,N_1759,N_1785);
nand U2554 (N_2554,N_1256,N_1123);
xor U2555 (N_2555,N_1239,N_1578);
or U2556 (N_2556,N_1637,N_1402);
nand U2557 (N_2557,N_1530,N_1117);
nand U2558 (N_2558,N_1530,N_1064);
or U2559 (N_2559,N_1692,N_1803);
or U2560 (N_2560,N_1511,N_1185);
and U2561 (N_2561,N_1917,N_1786);
or U2562 (N_2562,N_1197,N_1988);
and U2563 (N_2563,N_1569,N_1915);
or U2564 (N_2564,N_1176,N_1209);
or U2565 (N_2565,N_1211,N_1942);
nand U2566 (N_2566,N_1875,N_1330);
or U2567 (N_2567,N_1517,N_1502);
and U2568 (N_2568,N_1111,N_1779);
or U2569 (N_2569,N_1848,N_1429);
or U2570 (N_2570,N_1292,N_1537);
nand U2571 (N_2571,N_1334,N_1839);
xnor U2572 (N_2572,N_1069,N_1317);
and U2573 (N_2573,N_1311,N_1922);
and U2574 (N_2574,N_1742,N_1469);
nand U2575 (N_2575,N_1830,N_1662);
nor U2576 (N_2576,N_1128,N_1876);
and U2577 (N_2577,N_1918,N_1049);
or U2578 (N_2578,N_1764,N_1407);
nand U2579 (N_2579,N_1667,N_1774);
nor U2580 (N_2580,N_1937,N_1013);
nand U2581 (N_2581,N_1421,N_1157);
xor U2582 (N_2582,N_1778,N_1766);
or U2583 (N_2583,N_1275,N_1345);
and U2584 (N_2584,N_1250,N_1974);
nand U2585 (N_2585,N_1584,N_1981);
nor U2586 (N_2586,N_1773,N_1242);
nor U2587 (N_2587,N_1720,N_1296);
nor U2588 (N_2588,N_1887,N_1230);
nor U2589 (N_2589,N_1283,N_1597);
and U2590 (N_2590,N_1413,N_1482);
nor U2591 (N_2591,N_1035,N_1828);
nand U2592 (N_2592,N_1255,N_1350);
nand U2593 (N_2593,N_1964,N_1628);
and U2594 (N_2594,N_1080,N_1287);
and U2595 (N_2595,N_1682,N_1120);
and U2596 (N_2596,N_1164,N_1544);
and U2597 (N_2597,N_1424,N_1183);
and U2598 (N_2598,N_1143,N_1174);
nor U2599 (N_2599,N_1909,N_1910);
nor U2600 (N_2600,N_1588,N_1368);
nand U2601 (N_2601,N_1289,N_1057);
and U2602 (N_2602,N_1676,N_1877);
or U2603 (N_2603,N_1223,N_1876);
and U2604 (N_2604,N_1975,N_1212);
or U2605 (N_2605,N_1041,N_1028);
nor U2606 (N_2606,N_1385,N_1463);
nor U2607 (N_2607,N_1473,N_1858);
and U2608 (N_2608,N_1236,N_1203);
and U2609 (N_2609,N_1854,N_1242);
and U2610 (N_2610,N_1638,N_1503);
nand U2611 (N_2611,N_1756,N_1305);
and U2612 (N_2612,N_1601,N_1688);
and U2613 (N_2613,N_1584,N_1277);
nor U2614 (N_2614,N_1326,N_1787);
and U2615 (N_2615,N_1582,N_1360);
or U2616 (N_2616,N_1715,N_1719);
or U2617 (N_2617,N_1289,N_1314);
or U2618 (N_2618,N_1898,N_1020);
or U2619 (N_2619,N_1424,N_1152);
nor U2620 (N_2620,N_1173,N_1767);
or U2621 (N_2621,N_1966,N_1166);
or U2622 (N_2622,N_1804,N_1890);
nor U2623 (N_2623,N_1023,N_1322);
or U2624 (N_2624,N_1223,N_1986);
or U2625 (N_2625,N_1605,N_1680);
and U2626 (N_2626,N_1220,N_1439);
nor U2627 (N_2627,N_1430,N_1266);
nor U2628 (N_2628,N_1634,N_1834);
nand U2629 (N_2629,N_1583,N_1883);
nor U2630 (N_2630,N_1953,N_1204);
and U2631 (N_2631,N_1727,N_1845);
or U2632 (N_2632,N_1187,N_1389);
and U2633 (N_2633,N_1599,N_1109);
nand U2634 (N_2634,N_1933,N_1052);
or U2635 (N_2635,N_1449,N_1222);
and U2636 (N_2636,N_1467,N_1004);
xor U2637 (N_2637,N_1497,N_1635);
xnor U2638 (N_2638,N_1463,N_1340);
nor U2639 (N_2639,N_1655,N_1585);
or U2640 (N_2640,N_1544,N_1652);
or U2641 (N_2641,N_1374,N_1084);
or U2642 (N_2642,N_1314,N_1850);
or U2643 (N_2643,N_1966,N_1906);
xnor U2644 (N_2644,N_1850,N_1510);
and U2645 (N_2645,N_1665,N_1847);
nand U2646 (N_2646,N_1511,N_1997);
nor U2647 (N_2647,N_1391,N_1676);
and U2648 (N_2648,N_1112,N_1918);
or U2649 (N_2649,N_1144,N_1649);
xor U2650 (N_2650,N_1044,N_1390);
and U2651 (N_2651,N_1605,N_1611);
nor U2652 (N_2652,N_1471,N_1459);
and U2653 (N_2653,N_1048,N_1207);
or U2654 (N_2654,N_1349,N_1161);
nor U2655 (N_2655,N_1012,N_1388);
nand U2656 (N_2656,N_1744,N_1406);
and U2657 (N_2657,N_1722,N_1930);
nor U2658 (N_2658,N_1680,N_1644);
nor U2659 (N_2659,N_1121,N_1408);
or U2660 (N_2660,N_1503,N_1084);
nand U2661 (N_2661,N_1687,N_1340);
and U2662 (N_2662,N_1589,N_1411);
or U2663 (N_2663,N_1191,N_1577);
nor U2664 (N_2664,N_1521,N_1588);
or U2665 (N_2665,N_1753,N_1985);
and U2666 (N_2666,N_1770,N_1114);
nor U2667 (N_2667,N_1730,N_1711);
and U2668 (N_2668,N_1067,N_1040);
nand U2669 (N_2669,N_1000,N_1963);
or U2670 (N_2670,N_1536,N_1637);
nand U2671 (N_2671,N_1176,N_1495);
nor U2672 (N_2672,N_1376,N_1869);
and U2673 (N_2673,N_1418,N_1396);
nor U2674 (N_2674,N_1585,N_1929);
and U2675 (N_2675,N_1394,N_1010);
and U2676 (N_2676,N_1035,N_1491);
nand U2677 (N_2677,N_1099,N_1550);
or U2678 (N_2678,N_1550,N_1247);
nand U2679 (N_2679,N_1084,N_1383);
or U2680 (N_2680,N_1112,N_1389);
nand U2681 (N_2681,N_1976,N_1054);
and U2682 (N_2682,N_1520,N_1973);
and U2683 (N_2683,N_1782,N_1746);
or U2684 (N_2684,N_1855,N_1237);
or U2685 (N_2685,N_1443,N_1487);
or U2686 (N_2686,N_1614,N_1247);
and U2687 (N_2687,N_1079,N_1651);
and U2688 (N_2688,N_1453,N_1589);
and U2689 (N_2689,N_1646,N_1653);
nor U2690 (N_2690,N_1736,N_1007);
nor U2691 (N_2691,N_1643,N_1771);
nor U2692 (N_2692,N_1218,N_1828);
nand U2693 (N_2693,N_1799,N_1671);
nor U2694 (N_2694,N_1534,N_1539);
and U2695 (N_2695,N_1223,N_1885);
nor U2696 (N_2696,N_1390,N_1624);
or U2697 (N_2697,N_1323,N_1530);
nand U2698 (N_2698,N_1206,N_1040);
nand U2699 (N_2699,N_1652,N_1022);
nor U2700 (N_2700,N_1914,N_1591);
or U2701 (N_2701,N_1884,N_1584);
nand U2702 (N_2702,N_1658,N_1299);
or U2703 (N_2703,N_1809,N_1918);
or U2704 (N_2704,N_1243,N_1896);
and U2705 (N_2705,N_1696,N_1897);
or U2706 (N_2706,N_1916,N_1611);
nor U2707 (N_2707,N_1856,N_1968);
nor U2708 (N_2708,N_1462,N_1914);
or U2709 (N_2709,N_1342,N_1201);
nand U2710 (N_2710,N_1127,N_1916);
nor U2711 (N_2711,N_1628,N_1811);
nor U2712 (N_2712,N_1915,N_1618);
nand U2713 (N_2713,N_1881,N_1247);
or U2714 (N_2714,N_1836,N_1851);
nand U2715 (N_2715,N_1302,N_1646);
or U2716 (N_2716,N_1550,N_1782);
and U2717 (N_2717,N_1101,N_1955);
and U2718 (N_2718,N_1913,N_1646);
or U2719 (N_2719,N_1688,N_1322);
or U2720 (N_2720,N_1025,N_1687);
nor U2721 (N_2721,N_1463,N_1171);
nor U2722 (N_2722,N_1440,N_1154);
nand U2723 (N_2723,N_1311,N_1751);
nand U2724 (N_2724,N_1412,N_1949);
or U2725 (N_2725,N_1793,N_1629);
and U2726 (N_2726,N_1739,N_1337);
nor U2727 (N_2727,N_1781,N_1386);
nand U2728 (N_2728,N_1436,N_1113);
nor U2729 (N_2729,N_1692,N_1075);
nand U2730 (N_2730,N_1252,N_1811);
xor U2731 (N_2731,N_1875,N_1654);
xor U2732 (N_2732,N_1535,N_1900);
and U2733 (N_2733,N_1380,N_1807);
nand U2734 (N_2734,N_1028,N_1951);
or U2735 (N_2735,N_1585,N_1531);
or U2736 (N_2736,N_1008,N_1232);
or U2737 (N_2737,N_1804,N_1448);
or U2738 (N_2738,N_1374,N_1972);
or U2739 (N_2739,N_1038,N_1686);
nor U2740 (N_2740,N_1785,N_1453);
and U2741 (N_2741,N_1495,N_1508);
nor U2742 (N_2742,N_1006,N_1201);
and U2743 (N_2743,N_1208,N_1583);
nand U2744 (N_2744,N_1976,N_1989);
or U2745 (N_2745,N_1276,N_1820);
nand U2746 (N_2746,N_1809,N_1322);
nor U2747 (N_2747,N_1195,N_1553);
or U2748 (N_2748,N_1932,N_1601);
or U2749 (N_2749,N_1527,N_1580);
and U2750 (N_2750,N_1281,N_1609);
nor U2751 (N_2751,N_1379,N_1387);
nand U2752 (N_2752,N_1401,N_1109);
or U2753 (N_2753,N_1915,N_1062);
or U2754 (N_2754,N_1199,N_1410);
nand U2755 (N_2755,N_1753,N_1666);
nor U2756 (N_2756,N_1493,N_1034);
nand U2757 (N_2757,N_1211,N_1519);
nor U2758 (N_2758,N_1070,N_1985);
or U2759 (N_2759,N_1251,N_1003);
or U2760 (N_2760,N_1930,N_1591);
and U2761 (N_2761,N_1762,N_1934);
nor U2762 (N_2762,N_1980,N_1219);
nand U2763 (N_2763,N_1582,N_1892);
or U2764 (N_2764,N_1484,N_1167);
nand U2765 (N_2765,N_1966,N_1320);
nand U2766 (N_2766,N_1663,N_1999);
and U2767 (N_2767,N_1682,N_1095);
and U2768 (N_2768,N_1167,N_1354);
nor U2769 (N_2769,N_1273,N_1256);
or U2770 (N_2770,N_1187,N_1684);
nand U2771 (N_2771,N_1779,N_1479);
or U2772 (N_2772,N_1049,N_1724);
or U2773 (N_2773,N_1127,N_1620);
nor U2774 (N_2774,N_1704,N_1755);
nand U2775 (N_2775,N_1287,N_1347);
nand U2776 (N_2776,N_1183,N_1404);
nor U2777 (N_2777,N_1068,N_1602);
and U2778 (N_2778,N_1159,N_1480);
nand U2779 (N_2779,N_1250,N_1696);
nor U2780 (N_2780,N_1554,N_1962);
or U2781 (N_2781,N_1688,N_1016);
or U2782 (N_2782,N_1274,N_1828);
and U2783 (N_2783,N_1024,N_1039);
and U2784 (N_2784,N_1142,N_1277);
or U2785 (N_2785,N_1107,N_1962);
nand U2786 (N_2786,N_1085,N_1796);
nand U2787 (N_2787,N_1011,N_1542);
nor U2788 (N_2788,N_1323,N_1803);
nand U2789 (N_2789,N_1436,N_1159);
or U2790 (N_2790,N_1732,N_1070);
nand U2791 (N_2791,N_1321,N_1263);
nand U2792 (N_2792,N_1393,N_1389);
and U2793 (N_2793,N_1602,N_1420);
xnor U2794 (N_2794,N_1262,N_1395);
nand U2795 (N_2795,N_1750,N_1959);
and U2796 (N_2796,N_1404,N_1807);
nand U2797 (N_2797,N_1905,N_1872);
nand U2798 (N_2798,N_1429,N_1797);
nand U2799 (N_2799,N_1235,N_1992);
nor U2800 (N_2800,N_1065,N_1327);
or U2801 (N_2801,N_1406,N_1583);
nand U2802 (N_2802,N_1859,N_1437);
or U2803 (N_2803,N_1474,N_1116);
and U2804 (N_2804,N_1472,N_1145);
and U2805 (N_2805,N_1393,N_1519);
nor U2806 (N_2806,N_1692,N_1299);
nand U2807 (N_2807,N_1941,N_1465);
nor U2808 (N_2808,N_1576,N_1524);
nand U2809 (N_2809,N_1493,N_1847);
nand U2810 (N_2810,N_1214,N_1719);
nand U2811 (N_2811,N_1346,N_1381);
nand U2812 (N_2812,N_1622,N_1421);
nor U2813 (N_2813,N_1584,N_1132);
nand U2814 (N_2814,N_1605,N_1962);
or U2815 (N_2815,N_1204,N_1336);
and U2816 (N_2816,N_1064,N_1400);
xnor U2817 (N_2817,N_1488,N_1985);
xnor U2818 (N_2818,N_1759,N_1645);
and U2819 (N_2819,N_1730,N_1362);
and U2820 (N_2820,N_1007,N_1952);
nor U2821 (N_2821,N_1092,N_1095);
nand U2822 (N_2822,N_1185,N_1247);
nor U2823 (N_2823,N_1335,N_1112);
or U2824 (N_2824,N_1252,N_1549);
and U2825 (N_2825,N_1396,N_1044);
nor U2826 (N_2826,N_1776,N_1716);
or U2827 (N_2827,N_1027,N_1284);
nor U2828 (N_2828,N_1661,N_1185);
nand U2829 (N_2829,N_1057,N_1156);
or U2830 (N_2830,N_1009,N_1459);
or U2831 (N_2831,N_1343,N_1237);
and U2832 (N_2832,N_1395,N_1054);
and U2833 (N_2833,N_1734,N_1947);
nand U2834 (N_2834,N_1549,N_1461);
nor U2835 (N_2835,N_1770,N_1614);
or U2836 (N_2836,N_1128,N_1903);
or U2837 (N_2837,N_1046,N_1371);
or U2838 (N_2838,N_1439,N_1938);
and U2839 (N_2839,N_1317,N_1444);
or U2840 (N_2840,N_1230,N_1934);
or U2841 (N_2841,N_1636,N_1369);
nand U2842 (N_2842,N_1307,N_1531);
or U2843 (N_2843,N_1800,N_1904);
and U2844 (N_2844,N_1304,N_1578);
and U2845 (N_2845,N_1805,N_1846);
nand U2846 (N_2846,N_1939,N_1373);
nor U2847 (N_2847,N_1497,N_1102);
or U2848 (N_2848,N_1260,N_1985);
nand U2849 (N_2849,N_1822,N_1858);
nand U2850 (N_2850,N_1325,N_1439);
and U2851 (N_2851,N_1281,N_1485);
and U2852 (N_2852,N_1472,N_1636);
nand U2853 (N_2853,N_1544,N_1781);
nor U2854 (N_2854,N_1529,N_1038);
nor U2855 (N_2855,N_1232,N_1601);
or U2856 (N_2856,N_1434,N_1254);
and U2857 (N_2857,N_1702,N_1812);
nand U2858 (N_2858,N_1883,N_1071);
and U2859 (N_2859,N_1700,N_1070);
and U2860 (N_2860,N_1012,N_1279);
and U2861 (N_2861,N_1642,N_1426);
nor U2862 (N_2862,N_1264,N_1467);
and U2863 (N_2863,N_1385,N_1472);
nand U2864 (N_2864,N_1245,N_1012);
or U2865 (N_2865,N_1623,N_1764);
and U2866 (N_2866,N_1986,N_1836);
or U2867 (N_2867,N_1317,N_1356);
or U2868 (N_2868,N_1455,N_1927);
nand U2869 (N_2869,N_1054,N_1542);
or U2870 (N_2870,N_1338,N_1723);
or U2871 (N_2871,N_1848,N_1166);
nand U2872 (N_2872,N_1163,N_1906);
or U2873 (N_2873,N_1473,N_1202);
nand U2874 (N_2874,N_1815,N_1806);
nand U2875 (N_2875,N_1120,N_1351);
and U2876 (N_2876,N_1627,N_1229);
nand U2877 (N_2877,N_1045,N_1235);
and U2878 (N_2878,N_1201,N_1832);
and U2879 (N_2879,N_1361,N_1759);
or U2880 (N_2880,N_1899,N_1828);
or U2881 (N_2881,N_1704,N_1379);
and U2882 (N_2882,N_1352,N_1809);
nor U2883 (N_2883,N_1455,N_1537);
or U2884 (N_2884,N_1262,N_1612);
nand U2885 (N_2885,N_1314,N_1237);
or U2886 (N_2886,N_1851,N_1349);
or U2887 (N_2887,N_1574,N_1266);
nor U2888 (N_2888,N_1499,N_1514);
nand U2889 (N_2889,N_1355,N_1031);
nor U2890 (N_2890,N_1426,N_1479);
nand U2891 (N_2891,N_1894,N_1245);
or U2892 (N_2892,N_1562,N_1201);
and U2893 (N_2893,N_1514,N_1047);
and U2894 (N_2894,N_1033,N_1696);
nand U2895 (N_2895,N_1544,N_1329);
nor U2896 (N_2896,N_1845,N_1494);
nand U2897 (N_2897,N_1845,N_1704);
and U2898 (N_2898,N_1327,N_1111);
and U2899 (N_2899,N_1438,N_1619);
or U2900 (N_2900,N_1660,N_1979);
nand U2901 (N_2901,N_1503,N_1032);
nand U2902 (N_2902,N_1745,N_1449);
or U2903 (N_2903,N_1066,N_1982);
and U2904 (N_2904,N_1203,N_1660);
or U2905 (N_2905,N_1970,N_1973);
xor U2906 (N_2906,N_1551,N_1436);
and U2907 (N_2907,N_1954,N_1304);
nor U2908 (N_2908,N_1972,N_1393);
nand U2909 (N_2909,N_1917,N_1686);
nor U2910 (N_2910,N_1844,N_1679);
or U2911 (N_2911,N_1982,N_1963);
nor U2912 (N_2912,N_1285,N_1720);
nand U2913 (N_2913,N_1453,N_1701);
or U2914 (N_2914,N_1943,N_1930);
and U2915 (N_2915,N_1374,N_1057);
nor U2916 (N_2916,N_1684,N_1691);
nor U2917 (N_2917,N_1010,N_1798);
or U2918 (N_2918,N_1996,N_1149);
nor U2919 (N_2919,N_1432,N_1935);
nand U2920 (N_2920,N_1930,N_1386);
nand U2921 (N_2921,N_1209,N_1249);
nor U2922 (N_2922,N_1334,N_1226);
or U2923 (N_2923,N_1707,N_1191);
or U2924 (N_2924,N_1443,N_1779);
and U2925 (N_2925,N_1685,N_1894);
nor U2926 (N_2926,N_1546,N_1310);
nand U2927 (N_2927,N_1459,N_1938);
and U2928 (N_2928,N_1178,N_1193);
nor U2929 (N_2929,N_1145,N_1390);
nor U2930 (N_2930,N_1542,N_1752);
and U2931 (N_2931,N_1637,N_1748);
nand U2932 (N_2932,N_1746,N_1124);
and U2933 (N_2933,N_1279,N_1281);
and U2934 (N_2934,N_1397,N_1597);
nor U2935 (N_2935,N_1132,N_1744);
or U2936 (N_2936,N_1277,N_1589);
and U2937 (N_2937,N_1880,N_1530);
nand U2938 (N_2938,N_1403,N_1776);
or U2939 (N_2939,N_1710,N_1095);
xor U2940 (N_2940,N_1850,N_1908);
and U2941 (N_2941,N_1364,N_1956);
or U2942 (N_2942,N_1831,N_1049);
and U2943 (N_2943,N_1890,N_1860);
or U2944 (N_2944,N_1307,N_1656);
and U2945 (N_2945,N_1728,N_1733);
or U2946 (N_2946,N_1892,N_1949);
and U2947 (N_2947,N_1950,N_1523);
and U2948 (N_2948,N_1678,N_1318);
nand U2949 (N_2949,N_1123,N_1729);
nand U2950 (N_2950,N_1423,N_1398);
nor U2951 (N_2951,N_1189,N_1013);
and U2952 (N_2952,N_1303,N_1634);
nor U2953 (N_2953,N_1987,N_1198);
nor U2954 (N_2954,N_1203,N_1259);
nand U2955 (N_2955,N_1794,N_1648);
nor U2956 (N_2956,N_1255,N_1045);
or U2957 (N_2957,N_1840,N_1744);
nor U2958 (N_2958,N_1901,N_1692);
nand U2959 (N_2959,N_1315,N_1296);
nor U2960 (N_2960,N_1351,N_1843);
and U2961 (N_2961,N_1767,N_1037);
and U2962 (N_2962,N_1392,N_1919);
nor U2963 (N_2963,N_1943,N_1280);
nand U2964 (N_2964,N_1718,N_1669);
nand U2965 (N_2965,N_1717,N_1741);
nand U2966 (N_2966,N_1484,N_1579);
or U2967 (N_2967,N_1887,N_1161);
and U2968 (N_2968,N_1119,N_1219);
nor U2969 (N_2969,N_1336,N_1859);
and U2970 (N_2970,N_1629,N_1734);
xnor U2971 (N_2971,N_1269,N_1309);
nand U2972 (N_2972,N_1576,N_1787);
nand U2973 (N_2973,N_1691,N_1846);
or U2974 (N_2974,N_1371,N_1885);
and U2975 (N_2975,N_1415,N_1285);
or U2976 (N_2976,N_1581,N_1537);
nand U2977 (N_2977,N_1421,N_1707);
and U2978 (N_2978,N_1474,N_1753);
and U2979 (N_2979,N_1606,N_1438);
and U2980 (N_2980,N_1107,N_1088);
nor U2981 (N_2981,N_1237,N_1378);
and U2982 (N_2982,N_1641,N_1364);
and U2983 (N_2983,N_1114,N_1787);
and U2984 (N_2984,N_1779,N_1398);
nand U2985 (N_2985,N_1068,N_1572);
or U2986 (N_2986,N_1892,N_1921);
nor U2987 (N_2987,N_1294,N_1100);
and U2988 (N_2988,N_1882,N_1517);
or U2989 (N_2989,N_1583,N_1005);
nand U2990 (N_2990,N_1769,N_1130);
nor U2991 (N_2991,N_1280,N_1552);
nor U2992 (N_2992,N_1502,N_1143);
nand U2993 (N_2993,N_1846,N_1879);
and U2994 (N_2994,N_1169,N_1618);
and U2995 (N_2995,N_1478,N_1677);
nor U2996 (N_2996,N_1836,N_1355);
and U2997 (N_2997,N_1485,N_1830);
or U2998 (N_2998,N_1254,N_1369);
nand U2999 (N_2999,N_1208,N_1260);
and U3000 (N_3000,N_2319,N_2943);
and U3001 (N_3001,N_2232,N_2992);
nand U3002 (N_3002,N_2686,N_2807);
nor U3003 (N_3003,N_2736,N_2853);
and U3004 (N_3004,N_2627,N_2732);
nand U3005 (N_3005,N_2510,N_2682);
or U3006 (N_3006,N_2747,N_2188);
and U3007 (N_3007,N_2879,N_2673);
or U3008 (N_3008,N_2438,N_2269);
or U3009 (N_3009,N_2267,N_2551);
nor U3010 (N_3010,N_2579,N_2541);
nor U3011 (N_3011,N_2256,N_2959);
nor U3012 (N_3012,N_2053,N_2578);
and U3013 (N_3013,N_2058,N_2638);
nor U3014 (N_3014,N_2937,N_2076);
or U3015 (N_3015,N_2544,N_2954);
or U3016 (N_3016,N_2873,N_2713);
or U3017 (N_3017,N_2146,N_2972);
nand U3018 (N_3018,N_2710,N_2831);
and U3019 (N_3019,N_2082,N_2254);
and U3020 (N_3020,N_2022,N_2392);
nor U3021 (N_3021,N_2208,N_2095);
and U3022 (N_3022,N_2289,N_2786);
nor U3023 (N_3023,N_2584,N_2397);
nor U3024 (N_3024,N_2801,N_2123);
or U3025 (N_3025,N_2539,N_2855);
or U3026 (N_3026,N_2883,N_2446);
nor U3027 (N_3027,N_2947,N_2344);
nand U3028 (N_3028,N_2362,N_2419);
and U3029 (N_3029,N_2019,N_2488);
nor U3030 (N_3030,N_2923,N_2555);
and U3031 (N_3031,N_2635,N_2859);
or U3032 (N_3032,N_2622,N_2485);
nand U3033 (N_3033,N_2039,N_2444);
and U3034 (N_3034,N_2910,N_2078);
nand U3035 (N_3035,N_2998,N_2926);
and U3036 (N_3036,N_2052,N_2315);
nand U3037 (N_3037,N_2200,N_2387);
nor U3038 (N_3038,N_2401,N_2154);
nand U3039 (N_3039,N_2901,N_2467);
nand U3040 (N_3040,N_2535,N_2817);
nor U3041 (N_3041,N_2089,N_2004);
and U3042 (N_3042,N_2288,N_2935);
or U3043 (N_3043,N_2865,N_2716);
nand U3044 (N_3044,N_2517,N_2083);
nand U3045 (N_3045,N_2618,N_2588);
nand U3046 (N_3046,N_2008,N_2814);
nand U3047 (N_3047,N_2258,N_2586);
nand U3048 (N_3048,N_2536,N_2382);
nand U3049 (N_3049,N_2385,N_2688);
nor U3050 (N_3050,N_2163,N_2305);
and U3051 (N_3051,N_2820,N_2689);
nand U3052 (N_3052,N_2354,N_2006);
nand U3053 (N_3053,N_2509,N_2270);
nor U3054 (N_3054,N_2511,N_2044);
or U3055 (N_3055,N_2648,N_2455);
or U3056 (N_3056,N_2667,N_2702);
nand U3057 (N_3057,N_2989,N_2028);
and U3058 (N_3058,N_2300,N_2913);
nand U3059 (N_3059,N_2169,N_2180);
nand U3060 (N_3060,N_2133,N_2693);
and U3061 (N_3061,N_2715,N_2091);
and U3062 (N_3062,N_2612,N_2582);
nor U3063 (N_3063,N_2669,N_2925);
and U3064 (N_3064,N_2152,N_2764);
nor U3065 (N_3065,N_2869,N_2224);
nand U3066 (N_3066,N_2007,N_2216);
nor U3067 (N_3067,N_2888,N_2748);
nand U3068 (N_3068,N_2366,N_2808);
or U3069 (N_3069,N_2338,N_2896);
and U3070 (N_3070,N_2283,N_2616);
nor U3071 (N_3071,N_2178,N_2632);
or U3072 (N_3072,N_2112,N_2376);
and U3073 (N_3073,N_2050,N_2184);
nand U3074 (N_3074,N_2166,N_2677);
and U3075 (N_3075,N_2065,N_2601);
nor U3076 (N_3076,N_2605,N_2294);
nor U3077 (N_3077,N_2404,N_2225);
nand U3078 (N_3078,N_2727,N_2221);
nor U3079 (N_3079,N_2029,N_2835);
nor U3080 (N_3080,N_2255,N_2212);
or U3081 (N_3081,N_2962,N_2381);
nor U3082 (N_3082,N_2378,N_2528);
and U3083 (N_3083,N_2406,N_2930);
nand U3084 (N_3084,N_2391,N_2646);
nand U3085 (N_3085,N_2505,N_2002);
nand U3086 (N_3086,N_2785,N_2529);
and U3087 (N_3087,N_2690,N_2563);
nand U3088 (N_3088,N_2661,N_2885);
nand U3089 (N_3089,N_2265,N_2778);
and U3090 (N_3090,N_2623,N_2779);
nor U3091 (N_3091,N_2754,N_2096);
or U3092 (N_3092,N_2183,N_2851);
and U3093 (N_3093,N_2304,N_2591);
nand U3094 (N_3094,N_2985,N_2033);
or U3095 (N_3095,N_2607,N_2284);
or U3096 (N_3096,N_2102,N_2629);
and U3097 (N_3097,N_2384,N_2461);
nor U3098 (N_3098,N_2922,N_2124);
and U3099 (N_3099,N_2068,N_2470);
nand U3100 (N_3100,N_2685,N_2651);
nand U3101 (N_3101,N_2633,N_2776);
and U3102 (N_3102,N_2904,N_2264);
xnor U3103 (N_3103,N_2171,N_2696);
nand U3104 (N_3104,N_2659,N_2099);
nor U3105 (N_3105,N_2457,N_2059);
nor U3106 (N_3106,N_2834,N_2558);
or U3107 (N_3107,N_2531,N_2781);
nand U3108 (N_3108,N_2513,N_2072);
or U3109 (N_3109,N_2608,N_2238);
nor U3110 (N_3110,N_2223,N_2365);
and U3111 (N_3111,N_2583,N_2156);
and U3112 (N_3112,N_2328,N_2905);
nor U3113 (N_3113,N_2186,N_2369);
nand U3114 (N_3114,N_2324,N_2699);
and U3115 (N_3115,N_2720,N_2092);
nor U3116 (N_3116,N_2427,N_2860);
or U3117 (N_3117,N_2540,N_2203);
or U3118 (N_3118,N_2011,N_2977);
nor U3119 (N_3119,N_2233,N_2897);
xor U3120 (N_3120,N_2405,N_2833);
nor U3121 (N_3121,N_2310,N_2014);
and U3122 (N_3122,N_2542,N_2527);
and U3123 (N_3123,N_2750,N_2486);
or U3124 (N_3124,N_2519,N_2088);
or U3125 (N_3125,N_2936,N_2818);
nand U3126 (N_3126,N_2295,N_2120);
nand U3127 (N_3127,N_2143,N_2230);
or U3128 (N_3128,N_2861,N_2347);
nand U3129 (N_3129,N_2386,N_2243);
nand U3130 (N_3130,N_2292,N_2744);
and U3131 (N_3131,N_2504,N_2458);
nand U3132 (N_3132,N_2423,N_2409);
nand U3133 (N_3133,N_2280,N_2440);
or U3134 (N_3134,N_2759,N_2692);
nor U3135 (N_3135,N_2062,N_2581);
and U3136 (N_3136,N_2085,N_2153);
nor U3137 (N_3137,N_2740,N_2484);
nor U3138 (N_3138,N_2907,N_2864);
or U3139 (N_3139,N_2260,N_2771);
or U3140 (N_3140,N_2017,N_2676);
and U3141 (N_3141,N_2164,N_2978);
nor U3142 (N_3142,N_2031,N_2312);
nor U3143 (N_3143,N_2891,N_2021);
and U3144 (N_3144,N_2982,N_2886);
nand U3145 (N_3145,N_2707,N_2594);
and U3146 (N_3146,N_2435,N_2613);
and U3147 (N_3147,N_2367,N_2137);
nor U3148 (N_3148,N_2887,N_2942);
nand U3149 (N_3149,N_2032,N_2195);
and U3150 (N_3150,N_2734,N_2698);
and U3151 (N_3151,N_2970,N_2924);
nor U3152 (N_3152,N_2953,N_2566);
and U3153 (N_3153,N_2552,N_2619);
and U3154 (N_3154,N_2567,N_2572);
nor U3155 (N_3155,N_2706,N_2986);
or U3156 (N_3156,N_2691,N_2657);
or U3157 (N_3157,N_2190,N_2168);
xnor U3158 (N_3158,N_2758,N_2139);
or U3159 (N_3159,N_2144,N_2912);
or U3160 (N_3160,N_2063,N_2589);
nor U3161 (N_3161,N_2900,N_2674);
nor U3162 (N_3162,N_2079,N_2823);
nor U3163 (N_3163,N_2104,N_2979);
or U3164 (N_3164,N_2080,N_2398);
nand U3165 (N_3165,N_2148,N_2729);
nand U3166 (N_3166,N_2162,N_2849);
and U3167 (N_3167,N_2497,N_2760);
nand U3168 (N_3168,N_2523,N_2441);
nand U3169 (N_3169,N_2334,N_2739);
nor U3170 (N_3170,N_2991,N_2422);
and U3171 (N_3171,N_2201,N_2797);
or U3172 (N_3172,N_2332,N_2279);
nand U3173 (N_3173,N_2695,N_2330);
nand U3174 (N_3174,N_2066,N_2590);
nor U3175 (N_3175,N_2150,N_2556);
nand U3176 (N_3176,N_2013,N_2945);
nand U3177 (N_3177,N_2671,N_2030);
nand U3178 (N_3178,N_2631,N_2389);
and U3179 (N_3179,N_2246,N_2737);
or U3180 (N_3180,N_2287,N_2165);
or U3181 (N_3181,N_2210,N_2755);
nor U3182 (N_3182,N_2857,N_2122);
nand U3183 (N_3183,N_2048,N_2890);
nand U3184 (N_3184,N_2973,N_2198);
or U3185 (N_3185,N_2323,N_2463);
or U3186 (N_3186,N_2027,N_2805);
nand U3187 (N_3187,N_2316,N_2878);
nor U3188 (N_3188,N_2342,N_2204);
nand U3189 (N_3189,N_2763,N_2575);
and U3190 (N_3190,N_2432,N_2561);
or U3191 (N_3191,N_2838,N_2103);
or U3192 (N_3192,N_2158,N_2037);
nor U3193 (N_3193,N_2918,N_2061);
nor U3194 (N_3194,N_2051,N_2533);
nor U3195 (N_3195,N_2009,N_2309);
and U3196 (N_3196,N_2241,N_2626);
nand U3197 (N_3197,N_2955,N_2217);
nand U3198 (N_3198,N_2351,N_2850);
and U3199 (N_3199,N_2129,N_2275);
nand U3200 (N_3200,N_2360,N_2532);
nor U3201 (N_3201,N_2705,N_2147);
nor U3202 (N_3202,N_2487,N_2653);
nor U3203 (N_3203,N_2452,N_2361);
and U3204 (N_3204,N_2866,N_2100);
and U3205 (N_3205,N_2215,N_2917);
or U3206 (N_3206,N_2055,N_2483);
or U3207 (N_3207,N_2664,N_2403);
nor U3208 (N_3208,N_2408,N_2311);
nor U3209 (N_3209,N_2704,N_2421);
nor U3210 (N_3210,N_2862,N_2291);
or U3211 (N_3211,N_2209,N_2473);
nand U3212 (N_3212,N_2848,N_2666);
nor U3213 (N_3213,N_2253,N_2709);
and U3214 (N_3214,N_2116,N_2562);
or U3215 (N_3215,N_2714,N_2783);
nor U3216 (N_3216,N_2380,N_2250);
and U3217 (N_3217,N_2757,N_2546);
nor U3218 (N_3218,N_2000,N_2717);
or U3219 (N_3219,N_2073,N_2557);
and U3220 (N_3220,N_2293,N_2167);
or U3221 (N_3221,N_2114,N_2239);
and U3222 (N_3222,N_2041,N_2161);
and U3223 (N_3223,N_2784,N_2802);
or U3224 (N_3224,N_2313,N_2719);
nand U3225 (N_3225,N_2822,N_2951);
nor U3226 (N_3226,N_2881,N_2018);
nor U3227 (N_3227,N_2762,N_2151);
nor U3228 (N_3228,N_2663,N_2595);
or U3229 (N_3229,N_2346,N_2222);
or U3230 (N_3230,N_2624,N_2498);
nand U3231 (N_3231,N_2654,N_2773);
and U3232 (N_3232,N_2414,N_2573);
nor U3233 (N_3233,N_2500,N_2554);
nand U3234 (N_3234,N_2495,N_2597);
and U3235 (N_3235,N_2046,N_2026);
and U3236 (N_3236,N_2374,N_2956);
xor U3237 (N_3237,N_2938,N_2769);
and U3238 (N_3238,N_2454,N_2852);
and U3239 (N_3239,N_2520,N_2155);
or U3240 (N_3240,N_2585,N_2894);
and U3241 (N_3241,N_2273,N_2966);
nand U3242 (N_3242,N_2816,N_2827);
or U3243 (N_3243,N_2606,N_2325);
nand U3244 (N_3244,N_2110,N_2772);
nor U3245 (N_3245,N_2811,N_2206);
or U3246 (N_3246,N_2761,N_2242);
nor U3247 (N_3247,N_2262,N_2348);
and U3248 (N_3248,N_2842,N_2994);
and U3249 (N_3249,N_2940,N_2550);
or U3250 (N_3250,N_2929,N_2074);
nand U3251 (N_3251,N_2796,N_2396);
and U3252 (N_3252,N_2649,N_2756);
or U3253 (N_3253,N_2824,N_2069);
or U3254 (N_3254,N_2399,N_2415);
nand U3255 (N_3255,N_2482,N_2577);
nand U3256 (N_3256,N_2742,N_2798);
and U3257 (N_3257,N_2679,N_2218);
and U3258 (N_3258,N_2263,N_2126);
or U3259 (N_3259,N_2314,N_2571);
and U3260 (N_3260,N_2479,N_2106);
nor U3261 (N_3261,N_2899,N_2636);
nand U3262 (N_3262,N_2508,N_2064);
and U3263 (N_3263,N_2569,N_2281);
or U3264 (N_3264,N_2298,N_2060);
or U3265 (N_3265,N_2620,N_2322);
nor U3266 (N_3266,N_2057,N_2416);
and U3267 (N_3267,N_2788,N_2113);
and U3268 (N_3268,N_2919,N_2521);
and U3269 (N_3269,N_2799,N_2548);
xnor U3270 (N_3270,N_2199,N_2368);
nor U3271 (N_3271,N_2803,N_2678);
and U3272 (N_3272,N_2191,N_2854);
or U3273 (N_3273,N_2261,N_2042);
nand U3274 (N_3274,N_2024,N_2352);
or U3275 (N_3275,N_2410,N_2196);
or U3276 (N_3276,N_2081,N_2559);
or U3277 (N_3277,N_2173,N_2700);
or U3278 (N_3278,N_2634,N_2214);
nand U3279 (N_3279,N_2839,N_2600);
and U3280 (N_3280,N_2302,N_2856);
nand U3281 (N_3281,N_2812,N_2274);
nand U3282 (N_3282,N_2920,N_2400);
or U3283 (N_3283,N_2506,N_2468);
nor U3284 (N_3284,N_2456,N_2297);
nand U3285 (N_3285,N_2449,N_2832);
and U3286 (N_3286,N_2429,N_2968);
and U3287 (N_3287,N_2170,N_2117);
or U3288 (N_3288,N_2433,N_2372);
or U3289 (N_3289,N_2160,N_2645);
nand U3290 (N_3290,N_2639,N_2522);
or U3291 (N_3291,N_2375,N_2040);
and U3292 (N_3292,N_2988,N_2118);
or U3293 (N_3293,N_2765,N_2127);
nor U3294 (N_3294,N_2743,N_2967);
and U3295 (N_3295,N_2753,N_2580);
and U3296 (N_3296,N_2981,N_2576);
nor U3297 (N_3297,N_2921,N_2047);
nand U3298 (N_3298,N_2472,N_2202);
and U3299 (N_3299,N_2038,N_2290);
and U3300 (N_3300,N_2628,N_2383);
nor U3301 (N_3301,N_2830,N_2359);
nor U3302 (N_3302,N_2308,N_2697);
and U3303 (N_3303,N_2229,N_2983);
or U3304 (N_3304,N_2643,N_2708);
nand U3305 (N_3305,N_2355,N_2098);
nor U3306 (N_3306,N_2418,N_2430);
nand U3307 (N_3307,N_2931,N_2526);
or U3308 (N_3308,N_2231,N_2189);
and U3309 (N_3309,N_2932,N_2684);
and U3310 (N_3310,N_2553,N_2777);
nand U3311 (N_3311,N_2880,N_2428);
nor U3312 (N_3312,N_2592,N_2448);
nand U3313 (N_3313,N_2725,N_2244);
nand U3314 (N_3314,N_2530,N_2094);
nor U3315 (N_3315,N_2658,N_2278);
nor U3316 (N_3316,N_2889,N_2240);
nand U3317 (N_3317,N_2565,N_2105);
or U3318 (N_3318,N_2035,N_2775);
or U3319 (N_3319,N_2711,N_2303);
and U3320 (N_3320,N_2791,N_2211);
nor U3321 (N_3321,N_2701,N_2436);
nand U3322 (N_3322,N_2902,N_2642);
nor U3323 (N_3323,N_2426,N_2996);
nand U3324 (N_3324,N_2752,N_2395);
or U3325 (N_3325,N_2847,N_2949);
nand U3326 (N_3326,N_2491,N_2075);
nor U3327 (N_3327,N_2015,N_2373);
nand U3328 (N_3328,N_2538,N_2413);
nor U3329 (N_3329,N_2599,N_2837);
or U3330 (N_3330,N_2474,N_2445);
and U3331 (N_3331,N_2045,N_2939);
nand U3332 (N_3332,N_2895,N_2809);
and U3333 (N_3333,N_2172,N_2875);
or U3334 (N_3334,N_2543,N_2974);
and U3335 (N_3335,N_2990,N_2829);
nand U3336 (N_3336,N_2906,N_2515);
nor U3337 (N_3337,N_2142,N_2192);
or U3338 (N_3338,N_2615,N_2141);
or U3339 (N_3339,N_2025,N_2272);
or U3340 (N_3340,N_2794,N_2140);
nand U3341 (N_3341,N_2345,N_2101);
and U3342 (N_3342,N_2412,N_2249);
nor U3343 (N_3343,N_2054,N_2234);
nor U3344 (N_3344,N_2093,N_2841);
or U3345 (N_3345,N_2999,N_2207);
or U3346 (N_3346,N_2872,N_2726);
nand U3347 (N_3347,N_2687,N_2969);
and U3348 (N_3348,N_2478,N_2915);
or U3349 (N_3349,N_2020,N_2010);
nor U3350 (N_3350,N_2388,N_2537);
or U3351 (N_3351,N_2349,N_2787);
nor U3352 (N_3352,N_2251,N_2276);
nand U3353 (N_3353,N_2898,N_2795);
and U3354 (N_3354,N_2975,N_2723);
or U3355 (N_3355,N_2681,N_2683);
and U3356 (N_3356,N_2928,N_2724);
or U3357 (N_3357,N_2247,N_2703);
or U3358 (N_3358,N_2145,N_2296);
and U3359 (N_3359,N_2644,N_2656);
nor U3360 (N_3360,N_2460,N_2194);
or U3361 (N_3361,N_2877,N_2135);
nor U3362 (N_3362,N_2547,N_2489);
and U3363 (N_3363,N_2317,N_2252);
or U3364 (N_3364,N_2916,N_2950);
nor U3365 (N_3365,N_2205,N_2131);
or U3366 (N_3366,N_2181,N_2863);
nand U3367 (N_3367,N_2514,N_2005);
nand U3368 (N_3368,N_2179,N_2662);
nand U3369 (N_3369,N_2774,N_2259);
and U3370 (N_3370,N_2793,N_2884);
or U3371 (N_3371,N_2003,N_2086);
and U3372 (N_3372,N_2425,N_2944);
nand U3373 (N_3373,N_2672,N_2503);
or U3374 (N_3374,N_2333,N_2335);
or U3375 (N_3375,N_2282,N_2927);
nor U3376 (N_3376,N_2957,N_2023);
and U3377 (N_3377,N_2876,N_2496);
nor U3378 (N_3378,N_2868,N_2545);
xnor U3379 (N_3379,N_2892,N_2176);
and U3380 (N_3380,N_2908,N_2652);
or U3381 (N_3381,N_2665,N_2320);
nor U3382 (N_3382,N_2668,N_2364);
nand U3383 (N_3383,N_2193,N_2903);
nand U3384 (N_3384,N_2993,N_2056);
nor U3385 (N_3385,N_2825,N_2718);
nor U3386 (N_3386,N_2987,N_2749);
nor U3387 (N_3387,N_2434,N_2268);
or U3388 (N_3388,N_2329,N_2712);
nand U3389 (N_3389,N_2109,N_2012);
nand U3390 (N_3390,N_2507,N_2437);
nand U3391 (N_3391,N_2358,N_2431);
or U3392 (N_3392,N_2828,N_2286);
or U3393 (N_3393,N_2941,N_2331);
and U3394 (N_3394,N_2464,N_2130);
and U3395 (N_3395,N_2735,N_2070);
xnor U3396 (N_3396,N_2134,N_2840);
or U3397 (N_3397,N_2976,N_2768);
nand U3398 (N_3398,N_2893,N_2603);
nand U3399 (N_3399,N_2958,N_2997);
or U3400 (N_3400,N_2961,N_2914);
nor U3401 (N_3401,N_2227,N_2071);
and U3402 (N_3402,N_2640,N_2933);
nor U3403 (N_3403,N_2442,N_2236);
nor U3404 (N_3404,N_2821,N_2655);
nor U3405 (N_3405,N_2318,N_2459);
and U3406 (N_3406,N_2471,N_2266);
nand U3407 (N_3407,N_2336,N_2450);
and U3408 (N_3408,N_2248,N_2469);
and U3409 (N_3409,N_2534,N_2560);
nand U3410 (N_3410,N_2647,N_2353);
nand U3411 (N_3411,N_2271,N_2043);
nor U3412 (N_3412,N_2843,N_2077);
or U3413 (N_3413,N_2306,N_2477);
nor U3414 (N_3414,N_2237,N_2327);
or U3415 (N_3415,N_2049,N_2371);
or U3416 (N_3416,N_2357,N_2466);
and U3417 (N_3417,N_2277,N_2845);
or U3418 (N_3418,N_2617,N_2034);
or U3419 (N_3419,N_2858,N_2731);
nor U3420 (N_3420,N_2402,N_2965);
nand U3421 (N_3421,N_2637,N_2157);
nand U3422 (N_3422,N_2213,N_2159);
and U3423 (N_3423,N_2670,N_2728);
nor U3424 (N_3424,N_2393,N_2465);
or U3425 (N_3425,N_2394,N_2524);
or U3426 (N_3426,N_2340,N_2995);
or U3427 (N_3427,N_2946,N_2766);
nand U3428 (N_3428,N_2611,N_2767);
nand U3429 (N_3429,N_2115,N_2525);
and U3430 (N_3430,N_2596,N_2789);
or U3431 (N_3431,N_2307,N_2090);
nand U3432 (N_3432,N_2480,N_2462);
or U3433 (N_3433,N_2326,N_2136);
and U3434 (N_3434,N_2343,N_2447);
and U3435 (N_3435,N_2614,N_2417);
nor U3436 (N_3436,N_2602,N_2097);
nor U3437 (N_3437,N_2219,N_2518);
and U3438 (N_3438,N_2481,N_2245);
nor U3439 (N_3439,N_2337,N_2871);
and U3440 (N_3440,N_2493,N_2197);
and U3441 (N_3441,N_2502,N_2494);
and U3442 (N_3442,N_2813,N_2257);
nor U3443 (N_3443,N_2439,N_2108);
nand U3444 (N_3444,N_2490,N_2948);
nand U3445 (N_3445,N_2621,N_2138);
and U3446 (N_3446,N_2630,N_2492);
nor U3447 (N_3447,N_2604,N_2870);
or U3448 (N_3448,N_2960,N_2370);
nor U3449 (N_3449,N_2844,N_2733);
or U3450 (N_3450,N_2356,N_2836);
nor U3451 (N_3451,N_2815,N_2660);
and U3452 (N_3452,N_2751,N_2549);
or U3453 (N_3453,N_2730,N_2377);
nor U3454 (N_3454,N_2084,N_2512);
nand U3455 (N_3455,N_2182,N_2390);
nand U3456 (N_3456,N_2220,N_2187);
nand U3457 (N_3457,N_2177,N_2909);
or U3458 (N_3458,N_2800,N_2453);
xor U3459 (N_3459,N_2721,N_2185);
xnor U3460 (N_3460,N_2285,N_2121);
and U3461 (N_3461,N_2228,N_2610);
nor U3462 (N_3462,N_2411,N_2443);
and U3463 (N_3463,N_2971,N_2598);
nor U3464 (N_3464,N_2980,N_2379);
nor U3465 (N_3465,N_2174,N_2867);
and U3466 (N_3466,N_2516,N_2424);
or U3467 (N_3467,N_2568,N_2593);
nor U3468 (N_3468,N_2363,N_2746);
nor U3469 (N_3469,N_2119,N_2321);
nand U3470 (N_3470,N_2339,N_2111);
nand U3471 (N_3471,N_2036,N_2650);
nor U3472 (N_3472,N_2128,N_2846);
nand U3473 (N_3473,N_2934,N_2738);
nor U3474 (N_3474,N_2806,N_2819);
or U3475 (N_3475,N_2826,N_2570);
nor U3476 (N_3476,N_2722,N_2574);
or U3477 (N_3477,N_2780,N_2782);
nor U3478 (N_3478,N_2609,N_2226);
nand U3479 (N_3479,N_2882,N_2420);
and U3480 (N_3480,N_2790,N_2125);
and U3481 (N_3481,N_2984,N_2963);
and U3482 (N_3482,N_2175,N_2132);
nand U3483 (N_3483,N_2675,N_2235);
or U3484 (N_3484,N_2625,N_2067);
or U3485 (N_3485,N_2001,N_2804);
nand U3486 (N_3486,N_2476,N_2407);
nand U3487 (N_3487,N_2770,N_2501);
nor U3488 (N_3488,N_2301,N_2745);
or U3489 (N_3489,N_2564,N_2499);
nor U3490 (N_3490,N_2587,N_2741);
nor U3491 (N_3491,N_2451,N_2964);
nand U3492 (N_3492,N_2680,N_2087);
nor U3493 (N_3493,N_2016,N_2475);
nor U3494 (N_3494,N_2149,N_2874);
nor U3495 (N_3495,N_2107,N_2641);
nor U3496 (N_3496,N_2341,N_2299);
nand U3497 (N_3497,N_2694,N_2952);
nand U3498 (N_3498,N_2350,N_2792);
nor U3499 (N_3499,N_2911,N_2810);
nor U3500 (N_3500,N_2365,N_2524);
nand U3501 (N_3501,N_2387,N_2244);
or U3502 (N_3502,N_2383,N_2635);
and U3503 (N_3503,N_2554,N_2529);
or U3504 (N_3504,N_2948,N_2130);
nand U3505 (N_3505,N_2134,N_2884);
nor U3506 (N_3506,N_2956,N_2295);
nor U3507 (N_3507,N_2077,N_2729);
nand U3508 (N_3508,N_2115,N_2349);
nand U3509 (N_3509,N_2978,N_2324);
nand U3510 (N_3510,N_2360,N_2902);
and U3511 (N_3511,N_2055,N_2713);
nand U3512 (N_3512,N_2450,N_2178);
or U3513 (N_3513,N_2153,N_2702);
nor U3514 (N_3514,N_2889,N_2879);
and U3515 (N_3515,N_2980,N_2381);
and U3516 (N_3516,N_2045,N_2234);
and U3517 (N_3517,N_2714,N_2025);
nand U3518 (N_3518,N_2419,N_2611);
nand U3519 (N_3519,N_2543,N_2089);
and U3520 (N_3520,N_2052,N_2001);
nand U3521 (N_3521,N_2861,N_2671);
or U3522 (N_3522,N_2586,N_2291);
nand U3523 (N_3523,N_2646,N_2506);
and U3524 (N_3524,N_2274,N_2705);
and U3525 (N_3525,N_2692,N_2549);
nor U3526 (N_3526,N_2632,N_2541);
or U3527 (N_3527,N_2392,N_2806);
nor U3528 (N_3528,N_2204,N_2453);
nand U3529 (N_3529,N_2671,N_2290);
and U3530 (N_3530,N_2941,N_2921);
nand U3531 (N_3531,N_2687,N_2281);
and U3532 (N_3532,N_2444,N_2079);
xnor U3533 (N_3533,N_2653,N_2817);
and U3534 (N_3534,N_2440,N_2099);
and U3535 (N_3535,N_2276,N_2911);
or U3536 (N_3536,N_2012,N_2978);
nor U3537 (N_3537,N_2043,N_2553);
nand U3538 (N_3538,N_2586,N_2714);
and U3539 (N_3539,N_2335,N_2589);
or U3540 (N_3540,N_2590,N_2811);
and U3541 (N_3541,N_2480,N_2278);
nand U3542 (N_3542,N_2236,N_2853);
or U3543 (N_3543,N_2792,N_2396);
nor U3544 (N_3544,N_2074,N_2938);
and U3545 (N_3545,N_2883,N_2280);
nand U3546 (N_3546,N_2585,N_2445);
or U3547 (N_3547,N_2692,N_2161);
nand U3548 (N_3548,N_2489,N_2130);
or U3549 (N_3549,N_2538,N_2025);
nand U3550 (N_3550,N_2511,N_2777);
and U3551 (N_3551,N_2659,N_2365);
nand U3552 (N_3552,N_2397,N_2038);
or U3553 (N_3553,N_2857,N_2396);
or U3554 (N_3554,N_2859,N_2196);
or U3555 (N_3555,N_2089,N_2802);
nand U3556 (N_3556,N_2367,N_2920);
nor U3557 (N_3557,N_2213,N_2714);
nor U3558 (N_3558,N_2298,N_2938);
and U3559 (N_3559,N_2587,N_2366);
and U3560 (N_3560,N_2543,N_2232);
nand U3561 (N_3561,N_2182,N_2302);
and U3562 (N_3562,N_2417,N_2787);
and U3563 (N_3563,N_2438,N_2332);
and U3564 (N_3564,N_2481,N_2701);
nor U3565 (N_3565,N_2503,N_2554);
nand U3566 (N_3566,N_2659,N_2548);
nand U3567 (N_3567,N_2836,N_2735);
or U3568 (N_3568,N_2662,N_2571);
nor U3569 (N_3569,N_2892,N_2254);
nand U3570 (N_3570,N_2876,N_2762);
or U3571 (N_3571,N_2111,N_2127);
nor U3572 (N_3572,N_2275,N_2689);
and U3573 (N_3573,N_2660,N_2857);
and U3574 (N_3574,N_2434,N_2798);
nand U3575 (N_3575,N_2978,N_2489);
nor U3576 (N_3576,N_2596,N_2221);
or U3577 (N_3577,N_2519,N_2958);
or U3578 (N_3578,N_2648,N_2953);
or U3579 (N_3579,N_2446,N_2210);
nor U3580 (N_3580,N_2432,N_2241);
nor U3581 (N_3581,N_2156,N_2269);
nor U3582 (N_3582,N_2904,N_2258);
and U3583 (N_3583,N_2320,N_2618);
nor U3584 (N_3584,N_2364,N_2571);
nand U3585 (N_3585,N_2745,N_2807);
or U3586 (N_3586,N_2002,N_2831);
and U3587 (N_3587,N_2864,N_2837);
nand U3588 (N_3588,N_2463,N_2065);
and U3589 (N_3589,N_2444,N_2552);
nand U3590 (N_3590,N_2327,N_2330);
or U3591 (N_3591,N_2597,N_2569);
nand U3592 (N_3592,N_2973,N_2627);
and U3593 (N_3593,N_2971,N_2390);
nor U3594 (N_3594,N_2138,N_2285);
nand U3595 (N_3595,N_2221,N_2203);
nor U3596 (N_3596,N_2121,N_2719);
nand U3597 (N_3597,N_2648,N_2620);
and U3598 (N_3598,N_2487,N_2660);
or U3599 (N_3599,N_2314,N_2507);
and U3600 (N_3600,N_2336,N_2485);
and U3601 (N_3601,N_2239,N_2667);
nand U3602 (N_3602,N_2134,N_2203);
or U3603 (N_3603,N_2629,N_2671);
nand U3604 (N_3604,N_2166,N_2038);
and U3605 (N_3605,N_2750,N_2169);
nand U3606 (N_3606,N_2008,N_2758);
nor U3607 (N_3607,N_2796,N_2835);
or U3608 (N_3608,N_2603,N_2930);
nand U3609 (N_3609,N_2557,N_2445);
nand U3610 (N_3610,N_2102,N_2754);
and U3611 (N_3611,N_2557,N_2426);
or U3612 (N_3612,N_2082,N_2374);
and U3613 (N_3613,N_2514,N_2211);
nor U3614 (N_3614,N_2718,N_2589);
or U3615 (N_3615,N_2551,N_2914);
nand U3616 (N_3616,N_2406,N_2110);
nor U3617 (N_3617,N_2953,N_2620);
nand U3618 (N_3618,N_2067,N_2062);
and U3619 (N_3619,N_2960,N_2308);
xor U3620 (N_3620,N_2576,N_2684);
nand U3621 (N_3621,N_2699,N_2344);
nor U3622 (N_3622,N_2652,N_2722);
nor U3623 (N_3623,N_2299,N_2020);
or U3624 (N_3624,N_2167,N_2335);
nand U3625 (N_3625,N_2403,N_2381);
nor U3626 (N_3626,N_2013,N_2745);
nand U3627 (N_3627,N_2255,N_2215);
nor U3628 (N_3628,N_2877,N_2111);
or U3629 (N_3629,N_2084,N_2044);
xor U3630 (N_3630,N_2833,N_2286);
or U3631 (N_3631,N_2820,N_2279);
nor U3632 (N_3632,N_2225,N_2789);
nor U3633 (N_3633,N_2738,N_2474);
nor U3634 (N_3634,N_2235,N_2290);
nor U3635 (N_3635,N_2920,N_2102);
and U3636 (N_3636,N_2516,N_2269);
nand U3637 (N_3637,N_2549,N_2530);
and U3638 (N_3638,N_2852,N_2751);
or U3639 (N_3639,N_2183,N_2519);
and U3640 (N_3640,N_2384,N_2068);
nor U3641 (N_3641,N_2764,N_2274);
or U3642 (N_3642,N_2347,N_2428);
nand U3643 (N_3643,N_2696,N_2044);
nor U3644 (N_3644,N_2560,N_2993);
or U3645 (N_3645,N_2469,N_2581);
nand U3646 (N_3646,N_2965,N_2231);
or U3647 (N_3647,N_2590,N_2067);
and U3648 (N_3648,N_2728,N_2227);
and U3649 (N_3649,N_2892,N_2516);
nand U3650 (N_3650,N_2103,N_2098);
or U3651 (N_3651,N_2450,N_2151);
nand U3652 (N_3652,N_2605,N_2582);
nor U3653 (N_3653,N_2193,N_2857);
or U3654 (N_3654,N_2989,N_2526);
and U3655 (N_3655,N_2191,N_2150);
nor U3656 (N_3656,N_2530,N_2680);
nand U3657 (N_3657,N_2714,N_2330);
nor U3658 (N_3658,N_2844,N_2944);
or U3659 (N_3659,N_2084,N_2829);
or U3660 (N_3660,N_2721,N_2331);
nand U3661 (N_3661,N_2049,N_2546);
nand U3662 (N_3662,N_2337,N_2469);
and U3663 (N_3663,N_2064,N_2373);
nand U3664 (N_3664,N_2339,N_2005);
or U3665 (N_3665,N_2731,N_2610);
and U3666 (N_3666,N_2746,N_2092);
nand U3667 (N_3667,N_2062,N_2909);
and U3668 (N_3668,N_2958,N_2292);
and U3669 (N_3669,N_2377,N_2432);
nor U3670 (N_3670,N_2652,N_2599);
and U3671 (N_3671,N_2596,N_2516);
nand U3672 (N_3672,N_2277,N_2521);
xor U3673 (N_3673,N_2437,N_2815);
nor U3674 (N_3674,N_2441,N_2258);
nand U3675 (N_3675,N_2583,N_2798);
nand U3676 (N_3676,N_2405,N_2968);
or U3677 (N_3677,N_2807,N_2176);
or U3678 (N_3678,N_2497,N_2394);
nand U3679 (N_3679,N_2567,N_2557);
nor U3680 (N_3680,N_2596,N_2528);
or U3681 (N_3681,N_2493,N_2929);
or U3682 (N_3682,N_2863,N_2770);
and U3683 (N_3683,N_2357,N_2652);
or U3684 (N_3684,N_2335,N_2405);
nor U3685 (N_3685,N_2715,N_2101);
nor U3686 (N_3686,N_2260,N_2472);
or U3687 (N_3687,N_2905,N_2742);
and U3688 (N_3688,N_2219,N_2930);
or U3689 (N_3689,N_2706,N_2697);
and U3690 (N_3690,N_2723,N_2317);
or U3691 (N_3691,N_2355,N_2321);
nor U3692 (N_3692,N_2557,N_2275);
nand U3693 (N_3693,N_2704,N_2739);
and U3694 (N_3694,N_2953,N_2741);
and U3695 (N_3695,N_2066,N_2008);
nor U3696 (N_3696,N_2677,N_2216);
xnor U3697 (N_3697,N_2863,N_2197);
nor U3698 (N_3698,N_2924,N_2171);
or U3699 (N_3699,N_2228,N_2144);
nor U3700 (N_3700,N_2781,N_2208);
and U3701 (N_3701,N_2718,N_2673);
nand U3702 (N_3702,N_2647,N_2100);
or U3703 (N_3703,N_2640,N_2178);
nor U3704 (N_3704,N_2765,N_2891);
or U3705 (N_3705,N_2731,N_2762);
nor U3706 (N_3706,N_2237,N_2267);
and U3707 (N_3707,N_2204,N_2045);
nor U3708 (N_3708,N_2700,N_2758);
nor U3709 (N_3709,N_2380,N_2088);
or U3710 (N_3710,N_2218,N_2399);
nand U3711 (N_3711,N_2744,N_2440);
or U3712 (N_3712,N_2987,N_2183);
or U3713 (N_3713,N_2147,N_2175);
nor U3714 (N_3714,N_2452,N_2583);
nand U3715 (N_3715,N_2754,N_2911);
and U3716 (N_3716,N_2587,N_2030);
nor U3717 (N_3717,N_2754,N_2779);
nand U3718 (N_3718,N_2798,N_2106);
nor U3719 (N_3719,N_2827,N_2252);
or U3720 (N_3720,N_2784,N_2685);
or U3721 (N_3721,N_2092,N_2065);
and U3722 (N_3722,N_2095,N_2266);
and U3723 (N_3723,N_2591,N_2693);
or U3724 (N_3724,N_2476,N_2612);
or U3725 (N_3725,N_2368,N_2273);
and U3726 (N_3726,N_2093,N_2625);
and U3727 (N_3727,N_2815,N_2553);
nand U3728 (N_3728,N_2711,N_2341);
nand U3729 (N_3729,N_2044,N_2863);
nor U3730 (N_3730,N_2290,N_2199);
nand U3731 (N_3731,N_2004,N_2748);
and U3732 (N_3732,N_2510,N_2176);
and U3733 (N_3733,N_2357,N_2446);
or U3734 (N_3734,N_2343,N_2463);
nand U3735 (N_3735,N_2667,N_2949);
and U3736 (N_3736,N_2445,N_2672);
and U3737 (N_3737,N_2973,N_2298);
or U3738 (N_3738,N_2289,N_2932);
and U3739 (N_3739,N_2109,N_2903);
nand U3740 (N_3740,N_2636,N_2793);
nor U3741 (N_3741,N_2106,N_2084);
nand U3742 (N_3742,N_2329,N_2616);
or U3743 (N_3743,N_2044,N_2700);
and U3744 (N_3744,N_2720,N_2691);
and U3745 (N_3745,N_2612,N_2565);
or U3746 (N_3746,N_2516,N_2146);
and U3747 (N_3747,N_2483,N_2560);
and U3748 (N_3748,N_2584,N_2323);
and U3749 (N_3749,N_2202,N_2504);
and U3750 (N_3750,N_2876,N_2589);
or U3751 (N_3751,N_2691,N_2765);
nand U3752 (N_3752,N_2534,N_2918);
or U3753 (N_3753,N_2149,N_2496);
and U3754 (N_3754,N_2334,N_2809);
nor U3755 (N_3755,N_2909,N_2984);
nor U3756 (N_3756,N_2215,N_2330);
nor U3757 (N_3757,N_2521,N_2730);
nor U3758 (N_3758,N_2470,N_2772);
nand U3759 (N_3759,N_2043,N_2344);
nand U3760 (N_3760,N_2377,N_2436);
nand U3761 (N_3761,N_2326,N_2420);
nand U3762 (N_3762,N_2360,N_2517);
nand U3763 (N_3763,N_2249,N_2923);
nand U3764 (N_3764,N_2387,N_2743);
nor U3765 (N_3765,N_2960,N_2886);
and U3766 (N_3766,N_2370,N_2550);
nand U3767 (N_3767,N_2721,N_2461);
and U3768 (N_3768,N_2168,N_2704);
and U3769 (N_3769,N_2671,N_2267);
nor U3770 (N_3770,N_2695,N_2352);
or U3771 (N_3771,N_2923,N_2732);
and U3772 (N_3772,N_2477,N_2114);
or U3773 (N_3773,N_2749,N_2585);
nand U3774 (N_3774,N_2620,N_2595);
nor U3775 (N_3775,N_2285,N_2930);
nand U3776 (N_3776,N_2045,N_2924);
or U3777 (N_3777,N_2667,N_2752);
and U3778 (N_3778,N_2001,N_2800);
and U3779 (N_3779,N_2712,N_2910);
and U3780 (N_3780,N_2662,N_2080);
nand U3781 (N_3781,N_2291,N_2899);
nor U3782 (N_3782,N_2128,N_2979);
nor U3783 (N_3783,N_2592,N_2566);
nor U3784 (N_3784,N_2950,N_2840);
or U3785 (N_3785,N_2336,N_2048);
nand U3786 (N_3786,N_2722,N_2767);
or U3787 (N_3787,N_2283,N_2044);
nand U3788 (N_3788,N_2856,N_2396);
nor U3789 (N_3789,N_2952,N_2234);
nor U3790 (N_3790,N_2327,N_2829);
nor U3791 (N_3791,N_2632,N_2117);
nor U3792 (N_3792,N_2395,N_2788);
xor U3793 (N_3793,N_2327,N_2949);
nand U3794 (N_3794,N_2988,N_2858);
and U3795 (N_3795,N_2383,N_2981);
and U3796 (N_3796,N_2978,N_2517);
nand U3797 (N_3797,N_2774,N_2566);
xnor U3798 (N_3798,N_2196,N_2707);
or U3799 (N_3799,N_2129,N_2355);
and U3800 (N_3800,N_2639,N_2902);
nor U3801 (N_3801,N_2246,N_2007);
and U3802 (N_3802,N_2245,N_2609);
or U3803 (N_3803,N_2181,N_2784);
and U3804 (N_3804,N_2773,N_2930);
or U3805 (N_3805,N_2634,N_2636);
and U3806 (N_3806,N_2879,N_2622);
and U3807 (N_3807,N_2367,N_2753);
nor U3808 (N_3808,N_2186,N_2052);
and U3809 (N_3809,N_2280,N_2057);
nand U3810 (N_3810,N_2001,N_2610);
and U3811 (N_3811,N_2136,N_2437);
nand U3812 (N_3812,N_2159,N_2112);
xor U3813 (N_3813,N_2310,N_2946);
nor U3814 (N_3814,N_2495,N_2376);
nor U3815 (N_3815,N_2870,N_2980);
or U3816 (N_3816,N_2223,N_2059);
and U3817 (N_3817,N_2298,N_2422);
nand U3818 (N_3818,N_2596,N_2843);
or U3819 (N_3819,N_2237,N_2913);
and U3820 (N_3820,N_2703,N_2893);
nor U3821 (N_3821,N_2932,N_2518);
nor U3822 (N_3822,N_2287,N_2077);
or U3823 (N_3823,N_2963,N_2300);
nand U3824 (N_3824,N_2522,N_2274);
nor U3825 (N_3825,N_2248,N_2343);
nor U3826 (N_3826,N_2196,N_2948);
nand U3827 (N_3827,N_2609,N_2726);
or U3828 (N_3828,N_2387,N_2258);
and U3829 (N_3829,N_2452,N_2789);
nand U3830 (N_3830,N_2389,N_2473);
nor U3831 (N_3831,N_2725,N_2682);
nor U3832 (N_3832,N_2014,N_2805);
and U3833 (N_3833,N_2926,N_2695);
or U3834 (N_3834,N_2754,N_2893);
or U3835 (N_3835,N_2333,N_2139);
and U3836 (N_3836,N_2504,N_2780);
or U3837 (N_3837,N_2059,N_2747);
and U3838 (N_3838,N_2790,N_2681);
nand U3839 (N_3839,N_2005,N_2610);
nand U3840 (N_3840,N_2156,N_2263);
and U3841 (N_3841,N_2609,N_2699);
nor U3842 (N_3842,N_2785,N_2665);
or U3843 (N_3843,N_2023,N_2650);
nand U3844 (N_3844,N_2315,N_2398);
nand U3845 (N_3845,N_2608,N_2911);
and U3846 (N_3846,N_2620,N_2208);
or U3847 (N_3847,N_2772,N_2553);
nand U3848 (N_3848,N_2746,N_2374);
or U3849 (N_3849,N_2818,N_2364);
nand U3850 (N_3850,N_2296,N_2648);
or U3851 (N_3851,N_2630,N_2005);
nor U3852 (N_3852,N_2144,N_2950);
nor U3853 (N_3853,N_2210,N_2926);
xnor U3854 (N_3854,N_2223,N_2857);
nor U3855 (N_3855,N_2421,N_2353);
or U3856 (N_3856,N_2942,N_2324);
nand U3857 (N_3857,N_2773,N_2329);
or U3858 (N_3858,N_2028,N_2539);
and U3859 (N_3859,N_2585,N_2293);
or U3860 (N_3860,N_2429,N_2320);
nand U3861 (N_3861,N_2594,N_2979);
nand U3862 (N_3862,N_2063,N_2339);
nand U3863 (N_3863,N_2154,N_2736);
nand U3864 (N_3864,N_2755,N_2658);
xnor U3865 (N_3865,N_2113,N_2312);
and U3866 (N_3866,N_2882,N_2922);
nand U3867 (N_3867,N_2072,N_2694);
nor U3868 (N_3868,N_2181,N_2244);
nand U3869 (N_3869,N_2462,N_2548);
or U3870 (N_3870,N_2072,N_2691);
and U3871 (N_3871,N_2697,N_2289);
nor U3872 (N_3872,N_2546,N_2923);
nor U3873 (N_3873,N_2525,N_2228);
nor U3874 (N_3874,N_2906,N_2265);
and U3875 (N_3875,N_2205,N_2328);
nand U3876 (N_3876,N_2002,N_2984);
and U3877 (N_3877,N_2939,N_2062);
nor U3878 (N_3878,N_2951,N_2519);
nand U3879 (N_3879,N_2582,N_2551);
or U3880 (N_3880,N_2296,N_2533);
and U3881 (N_3881,N_2068,N_2841);
or U3882 (N_3882,N_2044,N_2795);
or U3883 (N_3883,N_2477,N_2482);
nand U3884 (N_3884,N_2659,N_2066);
or U3885 (N_3885,N_2710,N_2418);
or U3886 (N_3886,N_2172,N_2171);
or U3887 (N_3887,N_2308,N_2718);
nand U3888 (N_3888,N_2081,N_2457);
or U3889 (N_3889,N_2238,N_2092);
and U3890 (N_3890,N_2374,N_2414);
or U3891 (N_3891,N_2749,N_2232);
or U3892 (N_3892,N_2223,N_2475);
nand U3893 (N_3893,N_2425,N_2301);
or U3894 (N_3894,N_2308,N_2629);
and U3895 (N_3895,N_2816,N_2535);
or U3896 (N_3896,N_2267,N_2207);
nand U3897 (N_3897,N_2161,N_2693);
or U3898 (N_3898,N_2346,N_2934);
and U3899 (N_3899,N_2114,N_2552);
or U3900 (N_3900,N_2650,N_2511);
or U3901 (N_3901,N_2211,N_2367);
or U3902 (N_3902,N_2225,N_2155);
and U3903 (N_3903,N_2886,N_2674);
nor U3904 (N_3904,N_2988,N_2854);
or U3905 (N_3905,N_2230,N_2360);
nand U3906 (N_3906,N_2362,N_2428);
and U3907 (N_3907,N_2255,N_2544);
nor U3908 (N_3908,N_2113,N_2956);
and U3909 (N_3909,N_2265,N_2336);
and U3910 (N_3910,N_2875,N_2084);
nand U3911 (N_3911,N_2318,N_2744);
and U3912 (N_3912,N_2403,N_2186);
or U3913 (N_3913,N_2469,N_2448);
or U3914 (N_3914,N_2580,N_2050);
and U3915 (N_3915,N_2736,N_2203);
nor U3916 (N_3916,N_2795,N_2146);
nand U3917 (N_3917,N_2693,N_2477);
and U3918 (N_3918,N_2276,N_2758);
nand U3919 (N_3919,N_2116,N_2919);
nand U3920 (N_3920,N_2488,N_2801);
and U3921 (N_3921,N_2238,N_2843);
nand U3922 (N_3922,N_2665,N_2469);
or U3923 (N_3923,N_2905,N_2679);
and U3924 (N_3924,N_2847,N_2765);
nor U3925 (N_3925,N_2883,N_2500);
nor U3926 (N_3926,N_2325,N_2090);
xor U3927 (N_3927,N_2298,N_2231);
or U3928 (N_3928,N_2362,N_2408);
and U3929 (N_3929,N_2453,N_2095);
nand U3930 (N_3930,N_2772,N_2457);
nand U3931 (N_3931,N_2118,N_2699);
nor U3932 (N_3932,N_2672,N_2083);
or U3933 (N_3933,N_2694,N_2965);
or U3934 (N_3934,N_2207,N_2670);
or U3935 (N_3935,N_2858,N_2458);
or U3936 (N_3936,N_2955,N_2482);
nand U3937 (N_3937,N_2551,N_2600);
or U3938 (N_3938,N_2386,N_2196);
or U3939 (N_3939,N_2481,N_2430);
nand U3940 (N_3940,N_2503,N_2727);
or U3941 (N_3941,N_2900,N_2168);
or U3942 (N_3942,N_2498,N_2268);
nor U3943 (N_3943,N_2854,N_2514);
and U3944 (N_3944,N_2027,N_2804);
xor U3945 (N_3945,N_2759,N_2527);
nand U3946 (N_3946,N_2971,N_2002);
nand U3947 (N_3947,N_2571,N_2060);
or U3948 (N_3948,N_2183,N_2245);
nor U3949 (N_3949,N_2248,N_2267);
nor U3950 (N_3950,N_2385,N_2338);
or U3951 (N_3951,N_2934,N_2910);
nand U3952 (N_3952,N_2074,N_2675);
nor U3953 (N_3953,N_2237,N_2955);
xnor U3954 (N_3954,N_2266,N_2244);
nand U3955 (N_3955,N_2852,N_2890);
or U3956 (N_3956,N_2311,N_2960);
nor U3957 (N_3957,N_2787,N_2891);
nand U3958 (N_3958,N_2899,N_2534);
and U3959 (N_3959,N_2365,N_2610);
and U3960 (N_3960,N_2626,N_2905);
or U3961 (N_3961,N_2652,N_2626);
and U3962 (N_3962,N_2779,N_2659);
or U3963 (N_3963,N_2746,N_2489);
and U3964 (N_3964,N_2224,N_2008);
or U3965 (N_3965,N_2371,N_2034);
nor U3966 (N_3966,N_2121,N_2886);
or U3967 (N_3967,N_2740,N_2958);
and U3968 (N_3968,N_2766,N_2417);
and U3969 (N_3969,N_2909,N_2143);
and U3970 (N_3970,N_2648,N_2412);
nor U3971 (N_3971,N_2627,N_2751);
nor U3972 (N_3972,N_2991,N_2130);
nor U3973 (N_3973,N_2634,N_2357);
nor U3974 (N_3974,N_2226,N_2858);
and U3975 (N_3975,N_2157,N_2876);
or U3976 (N_3976,N_2528,N_2250);
and U3977 (N_3977,N_2976,N_2786);
nand U3978 (N_3978,N_2726,N_2472);
nand U3979 (N_3979,N_2079,N_2882);
or U3980 (N_3980,N_2543,N_2113);
or U3981 (N_3981,N_2313,N_2754);
or U3982 (N_3982,N_2083,N_2222);
nand U3983 (N_3983,N_2666,N_2854);
nor U3984 (N_3984,N_2482,N_2369);
nor U3985 (N_3985,N_2432,N_2755);
nand U3986 (N_3986,N_2395,N_2986);
nor U3987 (N_3987,N_2599,N_2454);
nand U3988 (N_3988,N_2972,N_2545);
nor U3989 (N_3989,N_2060,N_2736);
and U3990 (N_3990,N_2152,N_2849);
and U3991 (N_3991,N_2479,N_2532);
and U3992 (N_3992,N_2858,N_2335);
or U3993 (N_3993,N_2729,N_2343);
or U3994 (N_3994,N_2013,N_2074);
and U3995 (N_3995,N_2386,N_2268);
and U3996 (N_3996,N_2005,N_2374);
or U3997 (N_3997,N_2663,N_2237);
and U3998 (N_3998,N_2170,N_2385);
and U3999 (N_3999,N_2350,N_2763);
or U4000 (N_4000,N_3823,N_3301);
and U4001 (N_4001,N_3002,N_3524);
nor U4002 (N_4002,N_3529,N_3239);
xnor U4003 (N_4003,N_3272,N_3518);
or U4004 (N_4004,N_3581,N_3038);
and U4005 (N_4005,N_3563,N_3662);
nand U4006 (N_4006,N_3300,N_3615);
and U4007 (N_4007,N_3220,N_3631);
nand U4008 (N_4008,N_3539,N_3015);
nor U4009 (N_4009,N_3785,N_3051);
and U4010 (N_4010,N_3171,N_3116);
nor U4011 (N_4011,N_3462,N_3277);
nand U4012 (N_4012,N_3311,N_3659);
nor U4013 (N_4013,N_3123,N_3621);
nand U4014 (N_4014,N_3401,N_3134);
nand U4015 (N_4015,N_3212,N_3299);
or U4016 (N_4016,N_3445,N_3256);
and U4017 (N_4017,N_3879,N_3587);
nand U4018 (N_4018,N_3538,N_3297);
and U4019 (N_4019,N_3818,N_3592);
and U4020 (N_4020,N_3309,N_3020);
nor U4021 (N_4021,N_3618,N_3996);
nor U4022 (N_4022,N_3578,N_3450);
nor U4023 (N_4023,N_3656,N_3866);
nor U4024 (N_4024,N_3897,N_3365);
nor U4025 (N_4025,N_3672,N_3479);
or U4026 (N_4026,N_3726,N_3834);
and U4027 (N_4027,N_3429,N_3630);
and U4028 (N_4028,N_3333,N_3037);
nor U4029 (N_4029,N_3155,N_3279);
nor U4030 (N_4030,N_3318,N_3503);
nand U4031 (N_4031,N_3419,N_3749);
nand U4032 (N_4032,N_3736,N_3213);
nand U4033 (N_4033,N_3515,N_3453);
nand U4034 (N_4034,N_3531,N_3676);
or U4035 (N_4035,N_3810,N_3308);
and U4036 (N_4036,N_3557,N_3101);
nand U4037 (N_4037,N_3642,N_3109);
or U4038 (N_4038,N_3759,N_3667);
nor U4039 (N_4039,N_3612,N_3701);
and U4040 (N_4040,N_3022,N_3035);
and U4041 (N_4041,N_3168,N_3635);
and U4042 (N_4042,N_3252,N_3902);
or U4043 (N_4043,N_3291,N_3968);
nand U4044 (N_4044,N_3704,N_3822);
and U4045 (N_4045,N_3454,N_3679);
nor U4046 (N_4046,N_3686,N_3156);
and U4047 (N_4047,N_3438,N_3657);
nor U4048 (N_4048,N_3043,N_3476);
nand U4049 (N_4049,N_3120,N_3164);
nand U4050 (N_4050,N_3236,N_3577);
or U4051 (N_4051,N_3629,N_3098);
nor U4052 (N_4052,N_3328,N_3077);
or U4053 (N_4053,N_3225,N_3148);
nor U4054 (N_4054,N_3521,N_3214);
nor U4055 (N_4055,N_3179,N_3888);
xor U4056 (N_4056,N_3568,N_3203);
or U4057 (N_4057,N_3858,N_3100);
or U4058 (N_4058,N_3268,N_3224);
nor U4059 (N_4059,N_3725,N_3458);
and U4060 (N_4060,N_3139,N_3674);
nor U4061 (N_4061,N_3535,N_3122);
or U4062 (N_4062,N_3233,N_3170);
nand U4063 (N_4063,N_3791,N_3840);
nor U4064 (N_4064,N_3547,N_3954);
or U4065 (N_4065,N_3856,N_3124);
or U4066 (N_4066,N_3378,N_3843);
nor U4067 (N_4067,N_3989,N_3663);
and U4068 (N_4068,N_3567,N_3293);
and U4069 (N_4069,N_3430,N_3505);
and U4070 (N_4070,N_3444,N_3697);
nand U4071 (N_4071,N_3979,N_3755);
nor U4072 (N_4072,N_3319,N_3865);
and U4073 (N_4073,N_3157,N_3808);
nor U4074 (N_4074,N_3330,N_3492);
nand U4075 (N_4075,N_3924,N_3584);
nand U4076 (N_4076,N_3934,N_3661);
nor U4077 (N_4077,N_3602,N_3741);
and U4078 (N_4078,N_3210,N_3732);
or U4079 (N_4079,N_3779,N_3972);
and U4080 (N_4080,N_3811,N_3498);
or U4081 (N_4081,N_3861,N_3588);
or U4082 (N_4082,N_3836,N_3243);
nor U4083 (N_4083,N_3008,N_3707);
xnor U4084 (N_4084,N_3281,N_3730);
and U4085 (N_4085,N_3130,N_3698);
nand U4086 (N_4086,N_3922,N_3951);
and U4087 (N_4087,N_3219,N_3542);
and U4088 (N_4088,N_3350,N_3081);
nand U4089 (N_4089,N_3396,N_3145);
and U4090 (N_4090,N_3315,N_3228);
and U4091 (N_4091,N_3017,N_3864);
and U4092 (N_4092,N_3942,N_3187);
nand U4093 (N_4093,N_3324,N_3893);
or U4094 (N_4094,N_3691,N_3906);
and U4095 (N_4095,N_3411,N_3862);
and U4096 (N_4096,N_3694,N_3606);
or U4097 (N_4097,N_3738,N_3706);
or U4098 (N_4098,N_3807,N_3937);
nand U4099 (N_4099,N_3267,N_3534);
nand U4100 (N_4100,N_3891,N_3094);
and U4101 (N_4101,N_3264,N_3889);
nand U4102 (N_4102,N_3414,N_3231);
nand U4103 (N_4103,N_3824,N_3447);
nand U4104 (N_4104,N_3000,N_3728);
nand U4105 (N_4105,N_3408,N_3747);
and U4106 (N_4106,N_3034,N_3623);
nor U4107 (N_4107,N_3446,N_3898);
and U4108 (N_4108,N_3377,N_3056);
nor U4109 (N_4109,N_3079,N_3522);
and U4110 (N_4110,N_3543,N_3734);
nand U4111 (N_4111,N_3669,N_3347);
or U4112 (N_4112,N_3312,N_3780);
nor U4113 (N_4113,N_3537,N_3711);
nor U4114 (N_4114,N_3456,N_3533);
nand U4115 (N_4115,N_3792,N_3467);
and U4116 (N_4116,N_3513,N_3677);
nand U4117 (N_4117,N_3371,N_3911);
nand U4118 (N_4118,N_3416,N_3607);
or U4119 (N_4119,N_3226,N_3923);
nand U4120 (N_4120,N_3245,N_3201);
or U4121 (N_4121,N_3649,N_3549);
or U4122 (N_4122,N_3742,N_3799);
nor U4123 (N_4123,N_3682,N_3582);
or U4124 (N_4124,N_3280,N_3192);
nor U4125 (N_4125,N_3143,N_3142);
nor U4126 (N_4126,N_3947,N_3975);
nor U4127 (N_4127,N_3658,N_3695);
nand U4128 (N_4128,N_3827,N_3980);
nor U4129 (N_4129,N_3527,N_3275);
nor U4130 (N_4130,N_3845,N_3604);
or U4131 (N_4131,N_3573,N_3571);
nor U4132 (N_4132,N_3422,N_3285);
nand U4133 (N_4133,N_3455,N_3193);
nand U4134 (N_4134,N_3135,N_3227);
and U4135 (N_4135,N_3765,N_3205);
nor U4136 (N_4136,N_3044,N_3617);
or U4137 (N_4137,N_3717,N_3407);
nor U4138 (N_4138,N_3758,N_3718);
and U4139 (N_4139,N_3525,N_3483);
nand U4140 (N_4140,N_3383,N_3241);
nor U4141 (N_4141,N_3781,N_3619);
and U4142 (N_4142,N_3198,N_3580);
and U4143 (N_4143,N_3036,N_3796);
nand U4144 (N_4144,N_3006,N_3919);
nor U4145 (N_4145,N_3912,N_3260);
nand U4146 (N_4146,N_3772,N_3217);
nand U4147 (N_4147,N_3232,N_3833);
or U4148 (N_4148,N_3962,N_3255);
and U4149 (N_4149,N_3990,N_3388);
nand U4150 (N_4150,N_3102,N_3119);
or U4151 (N_4151,N_3723,N_3992);
nand U4152 (N_4152,N_3999,N_3069);
or U4153 (N_4153,N_3355,N_3194);
and U4154 (N_4154,N_3128,N_3605);
nand U4155 (N_4155,N_3851,N_3775);
nor U4156 (N_4156,N_3838,N_3459);
nand U4157 (N_4157,N_3434,N_3640);
and U4158 (N_4158,N_3341,N_3366);
and U4159 (N_4159,N_3913,N_3372);
and U4160 (N_4160,N_3023,N_3868);
nor U4161 (N_4161,N_3511,N_3909);
nand U4162 (N_4162,N_3501,N_3976);
nand U4163 (N_4163,N_3819,N_3175);
nor U4164 (N_4164,N_3085,N_3837);
nand U4165 (N_4165,N_3042,N_3786);
or U4166 (N_4166,N_3121,N_3965);
and U4167 (N_4167,N_3141,N_3108);
or U4168 (N_4168,N_3565,N_3393);
or U4169 (N_4169,N_3334,N_3905);
or U4170 (N_4170,N_3439,N_3614);
nor U4171 (N_4171,N_3594,N_3502);
nor U4172 (N_4172,N_3849,N_3821);
nand U4173 (N_4173,N_3546,N_3544);
and U4174 (N_4174,N_3551,N_3065);
and U4175 (N_4175,N_3561,N_3952);
nor U4176 (N_4176,N_3288,N_3960);
nand U4177 (N_4177,N_3714,N_3787);
nor U4178 (N_4178,N_3722,N_3668);
nand U4179 (N_4179,N_3223,N_3579);
nor U4180 (N_4180,N_3877,N_3353);
and U4181 (N_4181,N_3673,N_3296);
and U4182 (N_4182,N_3744,N_3655);
or U4183 (N_4183,N_3111,N_3971);
or U4184 (N_4184,N_3391,N_3757);
or U4185 (N_4185,N_3364,N_3943);
and U4186 (N_4186,N_3046,N_3559);
and U4187 (N_4187,N_3977,N_3519);
and U4188 (N_4188,N_3251,N_3025);
and U4189 (N_4189,N_3392,N_3415);
nor U4190 (N_4190,N_3825,N_3835);
or U4191 (N_4191,N_3753,N_3746);
or U4192 (N_4192,N_3080,N_3215);
nand U4193 (N_4193,N_3553,N_3152);
nand U4194 (N_4194,N_3872,N_3941);
or U4195 (N_4195,N_3813,N_3165);
or U4196 (N_4196,N_3191,N_3751);
nand U4197 (N_4197,N_3093,N_3469);
nand U4198 (N_4198,N_3494,N_3465);
and U4199 (N_4199,N_3748,N_3622);
nor U4200 (N_4200,N_3370,N_3988);
nor U4201 (N_4201,N_3389,N_3316);
or U4202 (N_4202,N_3853,N_3591);
nor U4203 (N_4203,N_3063,N_3995);
or U4204 (N_4204,N_3910,N_3367);
or U4205 (N_4205,N_3981,N_3666);
and U4206 (N_4206,N_3530,N_3678);
and U4207 (N_4207,N_3814,N_3495);
or U4208 (N_4208,N_3671,N_3998);
nand U4209 (N_4209,N_3441,N_3274);
or U4210 (N_4210,N_3878,N_3869);
and U4211 (N_4211,N_3359,N_3013);
nand U4212 (N_4212,N_3600,N_3883);
and U4213 (N_4213,N_3499,N_3306);
and U4214 (N_4214,N_3335,N_3448);
nand U4215 (N_4215,N_3112,N_3766);
nor U4216 (N_4216,N_3871,N_3208);
and U4217 (N_4217,N_3735,N_3406);
and U4218 (N_4218,N_3461,N_3342);
nor U4219 (N_4219,N_3729,N_3027);
or U4220 (N_4220,N_3940,N_3860);
and U4221 (N_4221,N_3532,N_3183);
or U4222 (N_4222,N_3460,N_3481);
nand U4223 (N_4223,N_3442,N_3249);
and U4224 (N_4224,N_3696,N_3485);
nand U4225 (N_4225,N_3985,N_3918);
and U4226 (N_4226,N_3639,N_3830);
nand U4227 (N_4227,N_3806,N_3409);
or U4228 (N_4228,N_3030,N_3273);
nand U4229 (N_4229,N_3506,N_3204);
nor U4230 (N_4230,N_3693,N_3105);
and U4231 (N_4231,N_3449,N_3715);
and U4232 (N_4232,N_3049,N_3368);
or U4233 (N_4233,N_3826,N_3180);
and U4234 (N_4234,N_3059,N_3638);
and U4235 (N_4235,N_3993,N_3731);
and U4236 (N_4236,N_3084,N_3259);
nand U4237 (N_4237,N_3452,N_3764);
nand U4238 (N_4238,N_3554,N_3437);
and U4239 (N_4239,N_3457,N_3144);
and U4240 (N_4240,N_3727,N_3938);
nand U4241 (N_4241,N_3805,N_3174);
or U4242 (N_4242,N_3650,N_3558);
nand U4243 (N_4243,N_3054,N_3875);
or U4244 (N_4244,N_3946,N_3574);
nor U4245 (N_4245,N_3555,N_3903);
nand U4246 (N_4246,N_3881,N_3195);
or U4247 (N_4247,N_3379,N_3660);
or U4248 (N_4248,N_3514,N_3939);
and U4249 (N_4249,N_3894,N_3159);
or U4250 (N_4250,N_3705,N_3583);
nand U4251 (N_4251,N_3848,N_3490);
nor U4252 (N_4252,N_3762,N_3949);
nand U4253 (N_4253,N_3855,N_3859);
nand U4254 (N_4254,N_3138,N_3097);
or U4255 (N_4255,N_3890,N_3708);
nor U4256 (N_4256,N_3598,N_3047);
nand U4257 (N_4257,N_3320,N_3520);
nor U4258 (N_4258,N_3257,N_3340);
nand U4259 (N_4259,N_3776,N_3209);
nand U4260 (N_4260,N_3794,N_3003);
nor U4261 (N_4261,N_3254,N_3405);
or U4262 (N_4262,N_3160,N_3589);
and U4263 (N_4263,N_3244,N_3162);
nand U4264 (N_4264,N_3289,N_3750);
nand U4265 (N_4265,N_3634,N_3436);
or U4266 (N_4266,N_3899,N_3154);
nor U4267 (N_4267,N_3493,N_3637);
and U4268 (N_4268,N_3303,N_3424);
nor U4269 (N_4269,N_3181,N_3647);
nor U4270 (N_4270,N_3173,N_3106);
or U4271 (N_4271,N_3646,N_3062);
nor U4272 (N_4272,N_3354,N_3804);
nand U4273 (N_4273,N_3153,N_3018);
nor U4274 (N_4274,N_3852,N_3050);
nand U4275 (N_4275,N_3468,N_3048);
nand U4276 (N_4276,N_3474,N_3218);
nor U4277 (N_4277,N_3509,N_3246);
nand U4278 (N_4278,N_3473,N_3107);
or U4279 (N_4279,N_3278,N_3394);
nand U4280 (N_4280,N_3376,N_3817);
nand U4281 (N_4281,N_3126,N_3029);
xnor U4282 (N_4282,N_3351,N_3361);
or U4283 (N_4283,N_3550,N_3014);
nand U4284 (N_4284,N_3739,N_3031);
and U4285 (N_4285,N_3305,N_3828);
nand U4286 (N_4286,N_3375,N_3374);
nand U4287 (N_4287,N_3795,N_3643);
and U4288 (N_4288,N_3016,N_3681);
or U4289 (N_4289,N_3147,N_3433);
or U4290 (N_4290,N_3329,N_3876);
nand U4291 (N_4291,N_3240,N_3925);
nand U4292 (N_4292,N_3276,N_3435);
nor U4293 (N_4293,N_3071,N_3616);
or U4294 (N_4294,N_3541,N_3692);
nor U4295 (N_4295,N_3927,N_3752);
nand U4296 (N_4296,N_3398,N_3055);
or U4297 (N_4297,N_3724,N_3185);
nor U4298 (N_4298,N_3386,N_3075);
nor U4299 (N_4299,N_3060,N_3700);
nor U4300 (N_4300,N_3863,N_3778);
and U4301 (N_4301,N_3440,N_3095);
nand U4302 (N_4302,N_3788,N_3963);
or U4303 (N_4303,N_3358,N_3099);
and U4304 (N_4304,N_3137,N_3295);
and U4305 (N_4305,N_3713,N_3688);
nand U4306 (N_4306,N_3325,N_3200);
and U4307 (N_4307,N_3644,N_3294);
nor U4308 (N_4308,N_3104,N_3745);
and U4309 (N_4309,N_3763,N_3242);
or U4310 (N_4310,N_3585,N_3431);
nand U4311 (N_4311,N_3664,N_3167);
nor U4312 (N_4312,N_3207,N_3983);
nor U4313 (N_4313,N_3322,N_3345);
nand U4314 (N_4314,N_3427,N_3028);
and U4315 (N_4315,N_3633,N_3432);
or U4316 (N_4316,N_3874,N_3508);
or U4317 (N_4317,N_3338,N_3399);
nor U4318 (N_4318,N_3117,N_3512);
nand U4319 (N_4319,N_3072,N_3948);
and U4320 (N_4320,N_3332,N_3400);
nand U4321 (N_4321,N_3323,N_3994);
and U4322 (N_4322,N_3841,N_3052);
nor U4323 (N_4323,N_3058,N_3488);
nor U4324 (N_4324,N_3327,N_3884);
nand U4325 (N_4325,N_3412,N_3624);
nand U4326 (N_4326,N_3425,N_3395);
and U4327 (N_4327,N_3382,N_3870);
nand U4328 (N_4328,N_3045,N_3222);
nor U4329 (N_4329,N_3186,N_3074);
and U4330 (N_4330,N_3286,N_3188);
and U4331 (N_4331,N_3176,N_3712);
nor U4332 (N_4332,N_3090,N_3892);
nand U4333 (N_4333,N_3402,N_3966);
nand U4334 (N_4334,N_3978,N_3850);
or U4335 (N_4335,N_3463,N_3916);
nor U4336 (N_4336,N_3073,N_3645);
nor U4337 (N_4337,N_3936,N_3771);
nand U4338 (N_4338,N_3475,N_3944);
nor U4339 (N_4339,N_3783,N_3997);
nor U4340 (N_4340,N_3178,N_3011);
or U4341 (N_4341,N_3782,N_3613);
and U4342 (N_4342,N_3846,N_3304);
and U4343 (N_4343,N_3932,N_3070);
or U4344 (N_4344,N_3907,N_3928);
or U4345 (N_4345,N_3007,N_3648);
or U4346 (N_4346,N_3920,N_3313);
nand U4347 (N_4347,N_3504,N_3789);
or U4348 (N_4348,N_3917,N_3675);
and U4349 (N_4349,N_3896,N_3238);
and U4350 (N_4350,N_3873,N_3854);
and U4351 (N_4351,N_3428,N_3287);
and U4352 (N_4352,N_3829,N_3466);
and U4353 (N_4353,N_3720,N_3777);
and U4354 (N_4354,N_3410,N_3019);
or U4355 (N_4355,N_3163,N_3510);
nor U4356 (N_4356,N_3970,N_3536);
nand U4357 (N_4357,N_3348,N_3576);
or U4358 (N_4358,N_3302,N_3754);
nor U4359 (N_4359,N_3221,N_3211);
and U4360 (N_4360,N_3685,N_3767);
or U4361 (N_4361,N_3958,N_3092);
and U4362 (N_4362,N_3061,N_3959);
and U4363 (N_4363,N_3146,N_3344);
nand U4364 (N_4364,N_3710,N_3608);
nor U4365 (N_4365,N_3336,N_3247);
nor U4366 (N_4366,N_3339,N_3670);
and U4367 (N_4367,N_3477,N_3556);
or U4368 (N_4368,N_3169,N_3343);
or U4369 (N_4369,N_3307,N_3721);
nor U4370 (N_4370,N_3283,N_3769);
xnor U4371 (N_4371,N_3001,N_3689);
nor U4372 (N_4372,N_3262,N_3831);
or U4373 (N_4373,N_3683,N_3471);
and U4374 (N_4374,N_3387,N_3282);
or U4375 (N_4375,N_3687,N_3352);
or U4376 (N_4376,N_3626,N_3507);
nand U4377 (N_4377,N_3381,N_3196);
nor U4378 (N_4378,N_3362,N_3740);
nor U4379 (N_4379,N_3956,N_3690);
or U4380 (N_4380,N_3129,N_3802);
and U4381 (N_4381,N_3500,N_3258);
nand U4382 (N_4382,N_3253,N_3575);
xnor U4383 (N_4383,N_3610,N_3470);
nor U4384 (N_4384,N_3935,N_3041);
or U4385 (N_4385,N_3632,N_3699);
nor U4386 (N_4386,N_3839,N_3032);
nor U4387 (N_4387,N_3150,N_3967);
or U4388 (N_4388,N_3189,N_3206);
nor U4389 (N_4389,N_3057,N_3974);
and U4390 (N_4390,N_3653,N_3820);
nand U4391 (N_4391,N_3263,N_3651);
or U4392 (N_4392,N_3844,N_3380);
or U4393 (N_4393,N_3284,N_3184);
and U4394 (N_4394,N_3451,N_3867);
or U4395 (N_4395,N_3773,N_3526);
and U4396 (N_4396,N_3076,N_3161);
nand U4397 (N_4397,N_3847,N_3040);
nand U4398 (N_4398,N_3926,N_3012);
or U4399 (N_4399,N_3933,N_3832);
nand U4400 (N_4400,N_3140,N_3654);
nand U4401 (N_4401,N_3760,N_3815);
nand U4402 (N_4402,N_3373,N_3480);
nor U4403 (N_4403,N_3487,N_3929);
nand U4404 (N_4404,N_3290,N_3572);
nand U4405 (N_4405,N_3420,N_3314);
nor U4406 (N_4406,N_3709,N_3039);
or U4407 (N_4407,N_3784,N_3586);
nor U4408 (N_4408,N_3774,N_3986);
nand U4409 (N_4409,N_3271,N_3010);
nand U4410 (N_4410,N_3229,N_3596);
or U4411 (N_4411,N_3172,N_3953);
nand U4412 (N_4412,N_3908,N_3931);
nor U4413 (N_4413,N_3703,N_3113);
nor U4414 (N_4414,N_3895,N_3005);
nor U4415 (N_4415,N_3761,N_3096);
or U4416 (N_4416,N_3882,N_3816);
and U4417 (N_4417,N_3593,N_3114);
or U4418 (N_4418,N_3151,N_3930);
or U4419 (N_4419,N_3945,N_3321);
nand U4420 (N_4420,N_3298,N_3087);
nand U4421 (N_4421,N_3800,N_3793);
nand U4422 (N_4422,N_3955,N_3548);
or U4423 (N_4423,N_3957,N_3482);
or U4424 (N_4424,N_3756,N_3914);
nor U4425 (N_4425,N_3067,N_3516);
nor U4426 (N_4426,N_3472,N_3770);
and U4427 (N_4427,N_3950,N_3857);
and U4428 (N_4428,N_3250,N_3915);
and U4429 (N_4429,N_3982,N_3064);
and U4430 (N_4430,N_3118,N_3921);
nor U4431 (N_4431,N_3356,N_3234);
nor U4432 (N_4432,N_3743,N_3545);
and U4433 (N_4433,N_3641,N_3216);
or U4434 (N_4434,N_3880,N_3798);
nand U4435 (N_4435,N_3292,N_3357);
nor U4436 (N_4436,N_3131,N_3797);
nand U4437 (N_4437,N_3790,N_3603);
nand U4438 (N_4438,N_3363,N_3904);
nor U4439 (N_4439,N_3900,N_3125);
or U4440 (N_4440,N_3418,N_3021);
nor U4441 (N_4441,N_3423,N_3984);
or U4442 (N_4442,N_3346,N_3842);
nand U4443 (N_4443,N_3369,N_3136);
nor U4444 (N_4444,N_3540,N_3166);
and U4445 (N_4445,N_3803,N_3266);
nand U4446 (N_4446,N_3609,N_3569);
nand U4447 (N_4447,N_3235,N_3384);
nor U4448 (N_4448,N_3089,N_3496);
nor U4449 (N_4449,N_3489,N_3197);
and U4450 (N_4450,N_3360,N_3110);
and U4451 (N_4451,N_3620,N_3665);
nor U4452 (N_4452,N_3809,N_3611);
nand U4453 (N_4453,N_3237,N_3053);
nand U4454 (N_4454,N_3088,N_3182);
or U4455 (N_4455,N_3326,N_3397);
nand U4456 (N_4456,N_3404,N_3413);
nor U4457 (N_4457,N_3991,N_3570);
nand U4458 (N_4458,N_3443,N_3417);
or U4459 (N_4459,N_3627,N_3068);
nor U4460 (N_4460,N_3269,N_3270);
and U4461 (N_4461,N_3680,N_3497);
or U4462 (N_4462,N_3964,N_3684);
and U4463 (N_4463,N_3310,N_3024);
nand U4464 (N_4464,N_3331,N_3261);
or U4465 (N_4465,N_3158,N_3317);
or U4466 (N_4466,N_3082,N_3566);
or U4467 (N_4467,N_3523,N_3552);
nand U4468 (N_4468,N_3737,N_3628);
nand U4469 (N_4469,N_3083,N_3528);
and U4470 (N_4470,N_3337,N_3801);
and U4471 (N_4471,N_3478,N_3177);
or U4472 (N_4472,N_3265,N_3597);
nor U4473 (N_4473,N_3733,N_3517);
or U4474 (N_4474,N_3403,N_3103);
or U4475 (N_4475,N_3564,N_3887);
nand U4476 (N_4476,N_3560,N_3230);
nand U4477 (N_4477,N_3426,N_3149);
or U4478 (N_4478,N_3961,N_3486);
and U4479 (N_4479,N_3590,N_3595);
and U4480 (N_4480,N_3248,N_3464);
and U4481 (N_4481,N_3091,N_3385);
or U4482 (N_4482,N_3702,N_3115);
nor U4483 (N_4483,N_3199,N_3078);
nand U4484 (N_4484,N_3625,N_3886);
nand U4485 (N_4485,N_3421,N_3009);
or U4486 (N_4486,N_3026,N_3349);
nand U4487 (N_4487,N_3190,N_3599);
nand U4488 (N_4488,N_3987,N_3033);
nand U4489 (N_4489,N_3004,N_3901);
nand U4490 (N_4490,N_3133,N_3127);
and U4491 (N_4491,N_3973,N_3086);
nand U4492 (N_4492,N_3491,N_3484);
and U4493 (N_4493,N_3716,N_3768);
nand U4494 (N_4494,N_3719,N_3601);
or U4495 (N_4495,N_3132,N_3562);
or U4496 (N_4496,N_3636,N_3885);
and U4497 (N_4497,N_3969,N_3652);
or U4498 (N_4498,N_3390,N_3202);
and U4499 (N_4499,N_3812,N_3066);
or U4500 (N_4500,N_3440,N_3625);
nor U4501 (N_4501,N_3551,N_3971);
nand U4502 (N_4502,N_3636,N_3841);
nor U4503 (N_4503,N_3265,N_3802);
or U4504 (N_4504,N_3490,N_3276);
and U4505 (N_4505,N_3157,N_3103);
and U4506 (N_4506,N_3244,N_3576);
nor U4507 (N_4507,N_3170,N_3357);
or U4508 (N_4508,N_3398,N_3006);
and U4509 (N_4509,N_3655,N_3969);
or U4510 (N_4510,N_3381,N_3870);
nand U4511 (N_4511,N_3802,N_3768);
nand U4512 (N_4512,N_3356,N_3273);
or U4513 (N_4513,N_3785,N_3329);
nor U4514 (N_4514,N_3208,N_3715);
or U4515 (N_4515,N_3197,N_3823);
nand U4516 (N_4516,N_3400,N_3545);
or U4517 (N_4517,N_3040,N_3318);
nand U4518 (N_4518,N_3459,N_3468);
nor U4519 (N_4519,N_3917,N_3461);
or U4520 (N_4520,N_3482,N_3008);
nor U4521 (N_4521,N_3678,N_3195);
and U4522 (N_4522,N_3662,N_3554);
nor U4523 (N_4523,N_3485,N_3611);
nand U4524 (N_4524,N_3470,N_3710);
or U4525 (N_4525,N_3053,N_3115);
nand U4526 (N_4526,N_3288,N_3069);
nor U4527 (N_4527,N_3390,N_3550);
nor U4528 (N_4528,N_3371,N_3142);
and U4529 (N_4529,N_3372,N_3048);
nor U4530 (N_4530,N_3458,N_3290);
nor U4531 (N_4531,N_3621,N_3523);
or U4532 (N_4532,N_3109,N_3778);
or U4533 (N_4533,N_3379,N_3410);
or U4534 (N_4534,N_3028,N_3688);
or U4535 (N_4535,N_3309,N_3120);
nor U4536 (N_4536,N_3201,N_3060);
and U4537 (N_4537,N_3306,N_3132);
xnor U4538 (N_4538,N_3715,N_3550);
and U4539 (N_4539,N_3522,N_3344);
and U4540 (N_4540,N_3014,N_3063);
nor U4541 (N_4541,N_3879,N_3372);
nand U4542 (N_4542,N_3354,N_3395);
and U4543 (N_4543,N_3802,N_3395);
nand U4544 (N_4544,N_3536,N_3130);
and U4545 (N_4545,N_3288,N_3670);
and U4546 (N_4546,N_3579,N_3658);
nor U4547 (N_4547,N_3591,N_3888);
nand U4548 (N_4548,N_3648,N_3359);
or U4549 (N_4549,N_3768,N_3249);
or U4550 (N_4550,N_3780,N_3575);
nand U4551 (N_4551,N_3924,N_3533);
nand U4552 (N_4552,N_3815,N_3442);
nand U4553 (N_4553,N_3701,N_3424);
nor U4554 (N_4554,N_3678,N_3320);
or U4555 (N_4555,N_3420,N_3783);
or U4556 (N_4556,N_3130,N_3606);
nor U4557 (N_4557,N_3452,N_3409);
nand U4558 (N_4558,N_3521,N_3028);
nor U4559 (N_4559,N_3914,N_3462);
and U4560 (N_4560,N_3087,N_3019);
and U4561 (N_4561,N_3590,N_3136);
and U4562 (N_4562,N_3169,N_3386);
nand U4563 (N_4563,N_3028,N_3391);
nor U4564 (N_4564,N_3825,N_3967);
or U4565 (N_4565,N_3166,N_3759);
nor U4566 (N_4566,N_3848,N_3574);
nand U4567 (N_4567,N_3743,N_3849);
nor U4568 (N_4568,N_3925,N_3443);
or U4569 (N_4569,N_3779,N_3689);
nand U4570 (N_4570,N_3965,N_3280);
and U4571 (N_4571,N_3321,N_3487);
or U4572 (N_4572,N_3366,N_3595);
nor U4573 (N_4573,N_3761,N_3775);
or U4574 (N_4574,N_3948,N_3188);
nor U4575 (N_4575,N_3206,N_3018);
or U4576 (N_4576,N_3338,N_3953);
or U4577 (N_4577,N_3333,N_3737);
or U4578 (N_4578,N_3772,N_3961);
nor U4579 (N_4579,N_3064,N_3866);
or U4580 (N_4580,N_3766,N_3107);
nor U4581 (N_4581,N_3315,N_3747);
nor U4582 (N_4582,N_3425,N_3327);
or U4583 (N_4583,N_3745,N_3008);
nor U4584 (N_4584,N_3290,N_3563);
or U4585 (N_4585,N_3382,N_3841);
and U4586 (N_4586,N_3984,N_3743);
or U4587 (N_4587,N_3928,N_3433);
nor U4588 (N_4588,N_3212,N_3468);
or U4589 (N_4589,N_3087,N_3495);
and U4590 (N_4590,N_3707,N_3617);
and U4591 (N_4591,N_3316,N_3234);
and U4592 (N_4592,N_3805,N_3838);
nor U4593 (N_4593,N_3029,N_3243);
and U4594 (N_4594,N_3121,N_3263);
or U4595 (N_4595,N_3397,N_3855);
and U4596 (N_4596,N_3433,N_3593);
and U4597 (N_4597,N_3096,N_3991);
nand U4598 (N_4598,N_3764,N_3638);
and U4599 (N_4599,N_3050,N_3392);
nor U4600 (N_4600,N_3313,N_3527);
nor U4601 (N_4601,N_3886,N_3355);
and U4602 (N_4602,N_3226,N_3939);
or U4603 (N_4603,N_3717,N_3307);
nand U4604 (N_4604,N_3489,N_3640);
and U4605 (N_4605,N_3303,N_3053);
or U4606 (N_4606,N_3888,N_3013);
or U4607 (N_4607,N_3635,N_3905);
or U4608 (N_4608,N_3861,N_3524);
nor U4609 (N_4609,N_3582,N_3584);
or U4610 (N_4610,N_3310,N_3941);
nor U4611 (N_4611,N_3833,N_3948);
or U4612 (N_4612,N_3362,N_3584);
and U4613 (N_4613,N_3442,N_3643);
and U4614 (N_4614,N_3120,N_3755);
and U4615 (N_4615,N_3246,N_3698);
and U4616 (N_4616,N_3108,N_3560);
xor U4617 (N_4617,N_3419,N_3726);
and U4618 (N_4618,N_3693,N_3034);
or U4619 (N_4619,N_3173,N_3139);
and U4620 (N_4620,N_3783,N_3948);
and U4621 (N_4621,N_3710,N_3366);
nand U4622 (N_4622,N_3504,N_3423);
nand U4623 (N_4623,N_3184,N_3725);
nand U4624 (N_4624,N_3310,N_3960);
nor U4625 (N_4625,N_3386,N_3764);
and U4626 (N_4626,N_3528,N_3478);
nor U4627 (N_4627,N_3977,N_3995);
and U4628 (N_4628,N_3588,N_3520);
or U4629 (N_4629,N_3894,N_3697);
nand U4630 (N_4630,N_3607,N_3132);
nand U4631 (N_4631,N_3310,N_3813);
and U4632 (N_4632,N_3270,N_3858);
and U4633 (N_4633,N_3754,N_3602);
or U4634 (N_4634,N_3409,N_3799);
nor U4635 (N_4635,N_3715,N_3810);
nor U4636 (N_4636,N_3083,N_3520);
nor U4637 (N_4637,N_3575,N_3976);
and U4638 (N_4638,N_3479,N_3779);
and U4639 (N_4639,N_3427,N_3847);
nand U4640 (N_4640,N_3163,N_3872);
and U4641 (N_4641,N_3476,N_3180);
nand U4642 (N_4642,N_3474,N_3781);
or U4643 (N_4643,N_3120,N_3965);
and U4644 (N_4644,N_3703,N_3199);
and U4645 (N_4645,N_3654,N_3925);
or U4646 (N_4646,N_3624,N_3012);
and U4647 (N_4647,N_3235,N_3331);
nand U4648 (N_4648,N_3154,N_3730);
nand U4649 (N_4649,N_3014,N_3468);
nand U4650 (N_4650,N_3201,N_3383);
nand U4651 (N_4651,N_3248,N_3550);
and U4652 (N_4652,N_3419,N_3082);
nor U4653 (N_4653,N_3779,N_3907);
and U4654 (N_4654,N_3450,N_3645);
nor U4655 (N_4655,N_3350,N_3761);
or U4656 (N_4656,N_3392,N_3116);
nand U4657 (N_4657,N_3759,N_3124);
or U4658 (N_4658,N_3096,N_3653);
nand U4659 (N_4659,N_3527,N_3440);
or U4660 (N_4660,N_3862,N_3152);
nand U4661 (N_4661,N_3839,N_3221);
or U4662 (N_4662,N_3305,N_3928);
and U4663 (N_4663,N_3145,N_3587);
xor U4664 (N_4664,N_3527,N_3836);
and U4665 (N_4665,N_3954,N_3603);
or U4666 (N_4666,N_3820,N_3605);
or U4667 (N_4667,N_3597,N_3666);
nor U4668 (N_4668,N_3354,N_3198);
or U4669 (N_4669,N_3283,N_3418);
nor U4670 (N_4670,N_3028,N_3669);
nand U4671 (N_4671,N_3623,N_3544);
nand U4672 (N_4672,N_3240,N_3409);
or U4673 (N_4673,N_3725,N_3748);
nor U4674 (N_4674,N_3255,N_3788);
or U4675 (N_4675,N_3135,N_3106);
or U4676 (N_4676,N_3639,N_3233);
and U4677 (N_4677,N_3102,N_3358);
nor U4678 (N_4678,N_3687,N_3761);
and U4679 (N_4679,N_3168,N_3421);
or U4680 (N_4680,N_3079,N_3626);
nor U4681 (N_4681,N_3074,N_3734);
xor U4682 (N_4682,N_3181,N_3004);
nor U4683 (N_4683,N_3697,N_3762);
nor U4684 (N_4684,N_3289,N_3245);
and U4685 (N_4685,N_3063,N_3307);
and U4686 (N_4686,N_3133,N_3711);
or U4687 (N_4687,N_3621,N_3358);
and U4688 (N_4688,N_3737,N_3890);
nand U4689 (N_4689,N_3049,N_3228);
nand U4690 (N_4690,N_3501,N_3992);
nand U4691 (N_4691,N_3328,N_3342);
or U4692 (N_4692,N_3659,N_3507);
nand U4693 (N_4693,N_3505,N_3018);
nor U4694 (N_4694,N_3095,N_3478);
or U4695 (N_4695,N_3461,N_3089);
nor U4696 (N_4696,N_3972,N_3956);
nand U4697 (N_4697,N_3272,N_3088);
nor U4698 (N_4698,N_3216,N_3123);
and U4699 (N_4699,N_3245,N_3980);
or U4700 (N_4700,N_3316,N_3180);
or U4701 (N_4701,N_3736,N_3802);
nand U4702 (N_4702,N_3089,N_3382);
or U4703 (N_4703,N_3820,N_3872);
nor U4704 (N_4704,N_3706,N_3855);
or U4705 (N_4705,N_3140,N_3960);
and U4706 (N_4706,N_3233,N_3007);
nand U4707 (N_4707,N_3961,N_3549);
or U4708 (N_4708,N_3506,N_3915);
nand U4709 (N_4709,N_3683,N_3551);
nand U4710 (N_4710,N_3895,N_3885);
nor U4711 (N_4711,N_3187,N_3964);
or U4712 (N_4712,N_3931,N_3688);
and U4713 (N_4713,N_3802,N_3138);
nand U4714 (N_4714,N_3393,N_3269);
nor U4715 (N_4715,N_3185,N_3999);
and U4716 (N_4716,N_3871,N_3120);
and U4717 (N_4717,N_3920,N_3188);
or U4718 (N_4718,N_3358,N_3791);
and U4719 (N_4719,N_3642,N_3334);
and U4720 (N_4720,N_3986,N_3015);
or U4721 (N_4721,N_3299,N_3600);
and U4722 (N_4722,N_3706,N_3539);
nor U4723 (N_4723,N_3884,N_3248);
and U4724 (N_4724,N_3015,N_3699);
nand U4725 (N_4725,N_3703,N_3812);
and U4726 (N_4726,N_3417,N_3779);
nor U4727 (N_4727,N_3479,N_3163);
nand U4728 (N_4728,N_3577,N_3670);
or U4729 (N_4729,N_3965,N_3790);
nand U4730 (N_4730,N_3117,N_3058);
and U4731 (N_4731,N_3788,N_3195);
or U4732 (N_4732,N_3878,N_3936);
nand U4733 (N_4733,N_3588,N_3353);
and U4734 (N_4734,N_3673,N_3206);
and U4735 (N_4735,N_3600,N_3015);
nor U4736 (N_4736,N_3678,N_3256);
nor U4737 (N_4737,N_3303,N_3994);
or U4738 (N_4738,N_3018,N_3052);
nor U4739 (N_4739,N_3276,N_3614);
and U4740 (N_4740,N_3816,N_3119);
nor U4741 (N_4741,N_3139,N_3755);
nand U4742 (N_4742,N_3526,N_3385);
or U4743 (N_4743,N_3342,N_3322);
or U4744 (N_4744,N_3322,N_3275);
nor U4745 (N_4745,N_3725,N_3714);
nand U4746 (N_4746,N_3352,N_3481);
or U4747 (N_4747,N_3369,N_3821);
nor U4748 (N_4748,N_3844,N_3602);
or U4749 (N_4749,N_3940,N_3639);
nor U4750 (N_4750,N_3198,N_3055);
nand U4751 (N_4751,N_3025,N_3013);
and U4752 (N_4752,N_3821,N_3860);
and U4753 (N_4753,N_3866,N_3407);
nor U4754 (N_4754,N_3381,N_3854);
and U4755 (N_4755,N_3975,N_3049);
nor U4756 (N_4756,N_3346,N_3376);
and U4757 (N_4757,N_3302,N_3429);
nand U4758 (N_4758,N_3549,N_3916);
or U4759 (N_4759,N_3908,N_3284);
nand U4760 (N_4760,N_3069,N_3303);
nor U4761 (N_4761,N_3066,N_3598);
nor U4762 (N_4762,N_3881,N_3274);
nand U4763 (N_4763,N_3857,N_3995);
nand U4764 (N_4764,N_3299,N_3423);
nor U4765 (N_4765,N_3034,N_3615);
nor U4766 (N_4766,N_3702,N_3916);
nor U4767 (N_4767,N_3637,N_3051);
and U4768 (N_4768,N_3820,N_3336);
and U4769 (N_4769,N_3829,N_3249);
and U4770 (N_4770,N_3954,N_3388);
nor U4771 (N_4771,N_3977,N_3141);
and U4772 (N_4772,N_3101,N_3769);
or U4773 (N_4773,N_3200,N_3539);
nand U4774 (N_4774,N_3852,N_3178);
nor U4775 (N_4775,N_3702,N_3140);
and U4776 (N_4776,N_3017,N_3105);
nor U4777 (N_4777,N_3367,N_3071);
nand U4778 (N_4778,N_3923,N_3974);
and U4779 (N_4779,N_3547,N_3001);
and U4780 (N_4780,N_3245,N_3953);
nor U4781 (N_4781,N_3597,N_3798);
and U4782 (N_4782,N_3812,N_3852);
nand U4783 (N_4783,N_3334,N_3606);
and U4784 (N_4784,N_3001,N_3817);
nor U4785 (N_4785,N_3831,N_3842);
and U4786 (N_4786,N_3941,N_3890);
or U4787 (N_4787,N_3486,N_3353);
nor U4788 (N_4788,N_3069,N_3188);
nor U4789 (N_4789,N_3536,N_3941);
and U4790 (N_4790,N_3154,N_3560);
or U4791 (N_4791,N_3104,N_3144);
and U4792 (N_4792,N_3312,N_3441);
nor U4793 (N_4793,N_3314,N_3610);
nor U4794 (N_4794,N_3482,N_3724);
nand U4795 (N_4795,N_3165,N_3982);
and U4796 (N_4796,N_3114,N_3926);
nor U4797 (N_4797,N_3831,N_3754);
nor U4798 (N_4798,N_3985,N_3665);
and U4799 (N_4799,N_3727,N_3017);
nand U4800 (N_4800,N_3706,N_3258);
or U4801 (N_4801,N_3359,N_3857);
nand U4802 (N_4802,N_3402,N_3756);
nand U4803 (N_4803,N_3185,N_3731);
nand U4804 (N_4804,N_3710,N_3032);
nor U4805 (N_4805,N_3016,N_3035);
nand U4806 (N_4806,N_3194,N_3625);
or U4807 (N_4807,N_3806,N_3822);
and U4808 (N_4808,N_3127,N_3608);
and U4809 (N_4809,N_3223,N_3700);
nor U4810 (N_4810,N_3013,N_3206);
and U4811 (N_4811,N_3614,N_3726);
nor U4812 (N_4812,N_3028,N_3858);
nor U4813 (N_4813,N_3284,N_3925);
nor U4814 (N_4814,N_3301,N_3240);
or U4815 (N_4815,N_3348,N_3643);
nor U4816 (N_4816,N_3133,N_3519);
or U4817 (N_4817,N_3325,N_3674);
nor U4818 (N_4818,N_3563,N_3078);
nor U4819 (N_4819,N_3727,N_3928);
nand U4820 (N_4820,N_3339,N_3023);
nor U4821 (N_4821,N_3594,N_3604);
or U4822 (N_4822,N_3775,N_3355);
or U4823 (N_4823,N_3088,N_3633);
or U4824 (N_4824,N_3114,N_3517);
nor U4825 (N_4825,N_3873,N_3584);
nand U4826 (N_4826,N_3940,N_3652);
nand U4827 (N_4827,N_3688,N_3001);
nand U4828 (N_4828,N_3518,N_3174);
nand U4829 (N_4829,N_3182,N_3512);
nand U4830 (N_4830,N_3999,N_3722);
or U4831 (N_4831,N_3407,N_3028);
nor U4832 (N_4832,N_3394,N_3479);
and U4833 (N_4833,N_3041,N_3648);
and U4834 (N_4834,N_3852,N_3937);
and U4835 (N_4835,N_3068,N_3926);
nor U4836 (N_4836,N_3380,N_3245);
and U4837 (N_4837,N_3950,N_3366);
nand U4838 (N_4838,N_3758,N_3954);
nand U4839 (N_4839,N_3853,N_3894);
nor U4840 (N_4840,N_3906,N_3524);
nor U4841 (N_4841,N_3091,N_3194);
nor U4842 (N_4842,N_3571,N_3279);
or U4843 (N_4843,N_3145,N_3139);
nand U4844 (N_4844,N_3978,N_3470);
or U4845 (N_4845,N_3221,N_3298);
or U4846 (N_4846,N_3159,N_3631);
nand U4847 (N_4847,N_3190,N_3843);
and U4848 (N_4848,N_3258,N_3959);
and U4849 (N_4849,N_3144,N_3609);
nor U4850 (N_4850,N_3183,N_3250);
or U4851 (N_4851,N_3016,N_3761);
nor U4852 (N_4852,N_3194,N_3305);
or U4853 (N_4853,N_3002,N_3393);
or U4854 (N_4854,N_3754,N_3541);
xor U4855 (N_4855,N_3429,N_3537);
or U4856 (N_4856,N_3682,N_3586);
xnor U4857 (N_4857,N_3102,N_3213);
or U4858 (N_4858,N_3328,N_3899);
and U4859 (N_4859,N_3464,N_3565);
and U4860 (N_4860,N_3389,N_3961);
and U4861 (N_4861,N_3671,N_3262);
nand U4862 (N_4862,N_3017,N_3070);
and U4863 (N_4863,N_3383,N_3633);
nand U4864 (N_4864,N_3049,N_3825);
nand U4865 (N_4865,N_3302,N_3769);
and U4866 (N_4866,N_3971,N_3464);
nor U4867 (N_4867,N_3593,N_3315);
nor U4868 (N_4868,N_3071,N_3276);
and U4869 (N_4869,N_3449,N_3481);
and U4870 (N_4870,N_3061,N_3281);
and U4871 (N_4871,N_3670,N_3277);
nor U4872 (N_4872,N_3594,N_3613);
nor U4873 (N_4873,N_3460,N_3855);
or U4874 (N_4874,N_3095,N_3125);
and U4875 (N_4875,N_3165,N_3297);
and U4876 (N_4876,N_3317,N_3732);
nand U4877 (N_4877,N_3736,N_3896);
or U4878 (N_4878,N_3164,N_3540);
nor U4879 (N_4879,N_3954,N_3236);
or U4880 (N_4880,N_3137,N_3884);
nand U4881 (N_4881,N_3391,N_3661);
and U4882 (N_4882,N_3629,N_3537);
and U4883 (N_4883,N_3012,N_3260);
nor U4884 (N_4884,N_3175,N_3570);
nand U4885 (N_4885,N_3504,N_3225);
and U4886 (N_4886,N_3890,N_3414);
nand U4887 (N_4887,N_3488,N_3512);
and U4888 (N_4888,N_3495,N_3134);
nand U4889 (N_4889,N_3114,N_3135);
or U4890 (N_4890,N_3780,N_3564);
or U4891 (N_4891,N_3074,N_3536);
and U4892 (N_4892,N_3214,N_3263);
and U4893 (N_4893,N_3738,N_3260);
and U4894 (N_4894,N_3428,N_3304);
and U4895 (N_4895,N_3909,N_3795);
or U4896 (N_4896,N_3809,N_3137);
or U4897 (N_4897,N_3633,N_3082);
and U4898 (N_4898,N_3407,N_3812);
and U4899 (N_4899,N_3502,N_3985);
and U4900 (N_4900,N_3110,N_3888);
and U4901 (N_4901,N_3632,N_3692);
nand U4902 (N_4902,N_3369,N_3712);
or U4903 (N_4903,N_3652,N_3977);
and U4904 (N_4904,N_3736,N_3834);
nor U4905 (N_4905,N_3616,N_3756);
and U4906 (N_4906,N_3647,N_3223);
nand U4907 (N_4907,N_3303,N_3392);
or U4908 (N_4908,N_3771,N_3844);
nor U4909 (N_4909,N_3951,N_3127);
nor U4910 (N_4910,N_3458,N_3631);
nand U4911 (N_4911,N_3371,N_3506);
and U4912 (N_4912,N_3294,N_3062);
or U4913 (N_4913,N_3578,N_3660);
nor U4914 (N_4914,N_3290,N_3466);
and U4915 (N_4915,N_3157,N_3257);
and U4916 (N_4916,N_3491,N_3513);
nor U4917 (N_4917,N_3859,N_3434);
nor U4918 (N_4918,N_3134,N_3910);
or U4919 (N_4919,N_3063,N_3144);
and U4920 (N_4920,N_3609,N_3532);
nor U4921 (N_4921,N_3751,N_3695);
and U4922 (N_4922,N_3333,N_3163);
nor U4923 (N_4923,N_3075,N_3359);
and U4924 (N_4924,N_3381,N_3729);
nand U4925 (N_4925,N_3681,N_3205);
nor U4926 (N_4926,N_3857,N_3698);
nand U4927 (N_4927,N_3732,N_3918);
or U4928 (N_4928,N_3500,N_3973);
or U4929 (N_4929,N_3409,N_3576);
nor U4930 (N_4930,N_3003,N_3076);
nand U4931 (N_4931,N_3070,N_3446);
nor U4932 (N_4932,N_3420,N_3836);
and U4933 (N_4933,N_3226,N_3541);
or U4934 (N_4934,N_3740,N_3316);
nand U4935 (N_4935,N_3181,N_3135);
nand U4936 (N_4936,N_3675,N_3364);
nor U4937 (N_4937,N_3752,N_3132);
and U4938 (N_4938,N_3553,N_3982);
nand U4939 (N_4939,N_3833,N_3974);
nor U4940 (N_4940,N_3996,N_3691);
nand U4941 (N_4941,N_3932,N_3713);
nand U4942 (N_4942,N_3784,N_3043);
and U4943 (N_4943,N_3622,N_3356);
and U4944 (N_4944,N_3978,N_3488);
and U4945 (N_4945,N_3151,N_3374);
and U4946 (N_4946,N_3440,N_3283);
nand U4947 (N_4947,N_3570,N_3015);
or U4948 (N_4948,N_3119,N_3642);
and U4949 (N_4949,N_3249,N_3678);
nand U4950 (N_4950,N_3318,N_3521);
or U4951 (N_4951,N_3840,N_3562);
nand U4952 (N_4952,N_3497,N_3185);
and U4953 (N_4953,N_3934,N_3853);
and U4954 (N_4954,N_3851,N_3240);
and U4955 (N_4955,N_3384,N_3654);
nor U4956 (N_4956,N_3273,N_3262);
nand U4957 (N_4957,N_3639,N_3746);
or U4958 (N_4958,N_3046,N_3617);
nand U4959 (N_4959,N_3555,N_3901);
nor U4960 (N_4960,N_3823,N_3968);
nor U4961 (N_4961,N_3935,N_3759);
nand U4962 (N_4962,N_3041,N_3541);
nor U4963 (N_4963,N_3695,N_3409);
and U4964 (N_4964,N_3823,N_3564);
and U4965 (N_4965,N_3716,N_3101);
or U4966 (N_4966,N_3837,N_3507);
nor U4967 (N_4967,N_3349,N_3070);
or U4968 (N_4968,N_3050,N_3497);
nor U4969 (N_4969,N_3757,N_3169);
nand U4970 (N_4970,N_3752,N_3773);
xor U4971 (N_4971,N_3035,N_3689);
nand U4972 (N_4972,N_3110,N_3818);
or U4973 (N_4973,N_3740,N_3727);
and U4974 (N_4974,N_3953,N_3223);
and U4975 (N_4975,N_3771,N_3031);
nand U4976 (N_4976,N_3501,N_3194);
or U4977 (N_4977,N_3544,N_3001);
nand U4978 (N_4978,N_3013,N_3442);
or U4979 (N_4979,N_3489,N_3462);
and U4980 (N_4980,N_3773,N_3389);
nor U4981 (N_4981,N_3689,N_3658);
nand U4982 (N_4982,N_3456,N_3238);
and U4983 (N_4983,N_3983,N_3233);
nor U4984 (N_4984,N_3632,N_3826);
nor U4985 (N_4985,N_3955,N_3463);
nor U4986 (N_4986,N_3799,N_3641);
or U4987 (N_4987,N_3679,N_3570);
or U4988 (N_4988,N_3436,N_3464);
and U4989 (N_4989,N_3134,N_3547);
nand U4990 (N_4990,N_3010,N_3458);
nand U4991 (N_4991,N_3234,N_3461);
and U4992 (N_4992,N_3331,N_3362);
or U4993 (N_4993,N_3300,N_3485);
nand U4994 (N_4994,N_3143,N_3077);
nand U4995 (N_4995,N_3925,N_3100);
or U4996 (N_4996,N_3305,N_3786);
and U4997 (N_4997,N_3902,N_3510);
nand U4998 (N_4998,N_3626,N_3167);
and U4999 (N_4999,N_3987,N_3246);
and U5000 (N_5000,N_4788,N_4182);
nor U5001 (N_5001,N_4479,N_4366);
and U5002 (N_5002,N_4031,N_4512);
or U5003 (N_5003,N_4938,N_4945);
or U5004 (N_5004,N_4698,N_4865);
nor U5005 (N_5005,N_4626,N_4534);
nand U5006 (N_5006,N_4995,N_4800);
and U5007 (N_5007,N_4671,N_4746);
and U5008 (N_5008,N_4187,N_4809);
or U5009 (N_5009,N_4734,N_4267);
or U5010 (N_5010,N_4271,N_4404);
or U5011 (N_5011,N_4414,N_4230);
nand U5012 (N_5012,N_4381,N_4364);
and U5013 (N_5013,N_4039,N_4694);
nor U5014 (N_5014,N_4955,N_4577);
nand U5015 (N_5015,N_4637,N_4470);
and U5016 (N_5016,N_4873,N_4243);
and U5017 (N_5017,N_4360,N_4554);
nand U5018 (N_5018,N_4193,N_4987);
nor U5019 (N_5019,N_4067,N_4572);
and U5020 (N_5020,N_4318,N_4767);
nor U5021 (N_5021,N_4736,N_4260);
and U5022 (N_5022,N_4084,N_4921);
and U5023 (N_5023,N_4881,N_4427);
or U5024 (N_5024,N_4225,N_4612);
and U5025 (N_5025,N_4455,N_4622);
nor U5026 (N_5026,N_4802,N_4602);
or U5027 (N_5027,N_4019,N_4023);
nor U5028 (N_5028,N_4239,N_4748);
or U5029 (N_5029,N_4306,N_4310);
nor U5030 (N_5030,N_4365,N_4505);
and U5031 (N_5031,N_4652,N_4482);
and U5032 (N_5032,N_4200,N_4466);
nor U5033 (N_5033,N_4308,N_4847);
nor U5034 (N_5034,N_4695,N_4386);
nor U5035 (N_5035,N_4901,N_4538);
nor U5036 (N_5036,N_4887,N_4475);
nand U5037 (N_5037,N_4008,N_4131);
or U5038 (N_5038,N_4598,N_4165);
nand U5039 (N_5039,N_4400,N_4620);
and U5040 (N_5040,N_4049,N_4823);
or U5041 (N_5041,N_4026,N_4891);
nand U5042 (N_5042,N_4486,N_4269);
nor U5043 (N_5043,N_4774,N_4914);
or U5044 (N_5044,N_4937,N_4493);
xnor U5045 (N_5045,N_4720,N_4523);
and U5046 (N_5046,N_4359,N_4483);
nor U5047 (N_5047,N_4043,N_4457);
nand U5048 (N_5048,N_4605,N_4883);
and U5049 (N_5049,N_4643,N_4540);
nand U5050 (N_5050,N_4147,N_4932);
nor U5051 (N_5051,N_4928,N_4152);
or U5052 (N_5052,N_4875,N_4755);
nand U5053 (N_5053,N_4003,N_4964);
or U5054 (N_5054,N_4940,N_4839);
nand U5055 (N_5055,N_4357,N_4993);
or U5056 (N_5056,N_4218,N_4996);
and U5057 (N_5057,N_4775,N_4321);
nand U5058 (N_5058,N_4122,N_4034);
nand U5059 (N_5059,N_4056,N_4051);
or U5060 (N_5060,N_4744,N_4275);
nor U5061 (N_5061,N_4676,N_4781);
or U5062 (N_5062,N_4974,N_4918);
nand U5063 (N_5063,N_4545,N_4630);
or U5064 (N_5064,N_4579,N_4764);
nand U5065 (N_5065,N_4521,N_4172);
nor U5066 (N_5066,N_4002,N_4737);
or U5067 (N_5067,N_4681,N_4378);
and U5068 (N_5068,N_4356,N_4487);
and U5069 (N_5069,N_4819,N_4053);
nor U5070 (N_5070,N_4732,N_4441);
nor U5071 (N_5071,N_4343,N_4220);
or U5072 (N_5072,N_4494,N_4578);
nand U5073 (N_5073,N_4477,N_4634);
nand U5074 (N_5074,N_4687,N_4525);
nor U5075 (N_5075,N_4666,N_4708);
and U5076 (N_5076,N_4556,N_4596);
or U5077 (N_5077,N_4902,N_4586);
nand U5078 (N_5078,N_4134,N_4362);
nand U5079 (N_5079,N_4613,N_4735);
or U5080 (N_5080,N_4130,N_4768);
and U5081 (N_5081,N_4702,N_4078);
nand U5082 (N_5082,N_4190,N_4992);
and U5083 (N_5083,N_4428,N_4785);
and U5084 (N_5084,N_4725,N_4238);
and U5085 (N_5085,N_4363,N_4824);
and U5086 (N_5086,N_4433,N_4536);
and U5087 (N_5087,N_4226,N_4247);
and U5088 (N_5088,N_4944,N_4813);
nand U5089 (N_5089,N_4971,N_4291);
and U5090 (N_5090,N_4970,N_4168);
nand U5091 (N_5091,N_4422,N_4097);
nand U5092 (N_5092,N_4154,N_4565);
or U5093 (N_5093,N_4690,N_4266);
and U5094 (N_5094,N_4217,N_4001);
nor U5095 (N_5095,N_4094,N_4942);
and U5096 (N_5096,N_4765,N_4038);
or U5097 (N_5097,N_4953,N_4617);
or U5098 (N_5098,N_4115,N_4329);
or U5099 (N_5099,N_4183,N_4423);
and U5100 (N_5100,N_4608,N_4710);
and U5101 (N_5101,N_4432,N_4091);
and U5102 (N_5102,N_4777,N_4361);
nand U5103 (N_5103,N_4621,N_4389);
nor U5104 (N_5104,N_4370,N_4095);
and U5105 (N_5105,N_4917,N_4403);
nand U5106 (N_5106,N_4314,N_4185);
and U5107 (N_5107,N_4391,N_4281);
xnor U5108 (N_5108,N_4629,N_4495);
nor U5109 (N_5109,N_4843,N_4059);
nand U5110 (N_5110,N_4135,N_4196);
and U5111 (N_5111,N_4397,N_4782);
nor U5112 (N_5112,N_4575,N_4593);
nor U5113 (N_5113,N_4803,N_4826);
and U5114 (N_5114,N_4439,N_4346);
or U5115 (N_5115,N_4189,N_4128);
or U5116 (N_5116,N_4814,N_4611);
nor U5117 (N_5117,N_4715,N_4840);
or U5118 (N_5118,N_4029,N_4162);
or U5119 (N_5119,N_4300,N_4478);
or U5120 (N_5120,N_4568,N_4212);
nor U5121 (N_5121,N_4195,N_4730);
nor U5122 (N_5122,N_4589,N_4142);
and U5123 (N_5123,N_4639,N_4529);
nand U5124 (N_5124,N_4573,N_4551);
nand U5125 (N_5125,N_4713,N_4327);
and U5126 (N_5126,N_4526,N_4533);
nor U5127 (N_5127,N_4820,N_4237);
nor U5128 (N_5128,N_4390,N_4811);
nand U5129 (N_5129,N_4858,N_4743);
or U5130 (N_5130,N_4015,N_4245);
nor U5131 (N_5131,N_4885,N_4770);
or U5132 (N_5132,N_4828,N_4436);
or U5133 (N_5133,N_4170,N_4975);
or U5134 (N_5134,N_4194,N_4595);
and U5135 (N_5135,N_4492,N_4264);
or U5136 (N_5136,N_4157,N_4372);
nor U5137 (N_5137,N_4119,N_4060);
nor U5138 (N_5138,N_4377,N_4419);
nor U5139 (N_5139,N_4398,N_4462);
nand U5140 (N_5140,N_4209,N_4718);
or U5141 (N_5141,N_4345,N_4133);
nand U5142 (N_5142,N_4151,N_4651);
and U5143 (N_5143,N_4919,N_4005);
nand U5144 (N_5144,N_4440,N_4334);
nand U5145 (N_5145,N_4807,N_4654);
or U5146 (N_5146,N_4679,N_4600);
nand U5147 (N_5147,N_4552,N_4032);
or U5148 (N_5148,N_4369,N_4333);
nand U5149 (N_5149,N_4303,N_4009);
and U5150 (N_5150,N_4298,N_4956);
or U5151 (N_5151,N_4878,N_4197);
nor U5152 (N_5152,N_4606,N_4675);
nand U5153 (N_5153,N_4778,N_4065);
nand U5154 (N_5154,N_4438,N_4465);
or U5155 (N_5155,N_4740,N_4776);
nand U5156 (N_5156,N_4714,N_4160);
or U5157 (N_5157,N_4962,N_4640);
nand U5158 (N_5158,N_4831,N_4180);
nor U5159 (N_5159,N_4272,N_4036);
or U5160 (N_5160,N_4913,N_4434);
and U5161 (N_5161,N_4907,N_4751);
nand U5162 (N_5162,N_4549,N_4186);
and U5163 (N_5163,N_4110,N_4888);
nand U5164 (N_5164,N_4066,N_4326);
nor U5165 (N_5165,N_4752,N_4876);
and U5166 (N_5166,N_4924,N_4042);
or U5167 (N_5167,N_4931,N_4520);
and U5168 (N_5168,N_4382,N_4544);
nand U5169 (N_5169,N_4724,N_4559);
and U5170 (N_5170,N_4402,N_4144);
and U5171 (N_5171,N_4192,N_4830);
nor U5172 (N_5172,N_4783,N_4635);
nand U5173 (N_5173,N_4044,N_4516);
and U5174 (N_5174,N_4331,N_4158);
nand U5175 (N_5175,N_4836,N_4355);
and U5176 (N_5176,N_4421,N_4517);
nor U5177 (N_5177,N_4779,N_4650);
or U5178 (N_5178,N_4176,N_4668);
and U5179 (N_5179,N_4799,N_4786);
nand U5180 (N_5180,N_4846,N_4412);
nor U5181 (N_5181,N_4191,N_4408);
nand U5182 (N_5182,N_4978,N_4040);
nor U5183 (N_5183,N_4085,N_4252);
and U5184 (N_5184,N_4396,N_4712);
nor U5185 (N_5185,N_4242,N_4075);
nor U5186 (N_5186,N_4844,N_4817);
nand U5187 (N_5187,N_4892,N_4063);
nor U5188 (N_5188,N_4503,N_4105);
and U5189 (N_5189,N_4214,N_4205);
and U5190 (N_5190,N_4150,N_4050);
nor U5191 (N_5191,N_4371,N_4295);
and U5192 (N_5192,N_4805,N_4124);
or U5193 (N_5193,N_4335,N_4979);
nand U5194 (N_5194,N_4889,N_4092);
or U5195 (N_5195,N_4825,N_4862);
or U5196 (N_5196,N_4213,N_4215);
and U5197 (N_5197,N_4988,N_4121);
nor U5198 (N_5198,N_4757,N_4149);
nor U5199 (N_5199,N_4472,N_4219);
nand U5200 (N_5200,N_4723,N_4090);
nand U5201 (N_5201,N_4851,N_4570);
nor U5202 (N_5202,N_4244,N_4787);
nor U5203 (N_5203,N_4903,N_4283);
or U5204 (N_5204,N_4703,N_4977);
or U5205 (N_5205,N_4541,N_4104);
nand U5206 (N_5206,N_4895,N_4447);
nor U5207 (N_5207,N_4489,N_4347);
or U5208 (N_5208,N_4114,N_4101);
nand U5209 (N_5209,N_4341,N_4546);
or U5210 (N_5210,N_4967,N_4206);
nor U5211 (N_5211,N_4968,N_4502);
nor U5212 (N_5212,N_4431,N_4017);
nand U5213 (N_5213,N_4961,N_4481);
nand U5214 (N_5214,N_4474,N_4416);
nand U5215 (N_5215,N_4393,N_4437);
and U5216 (N_5216,N_4927,N_4276);
or U5217 (N_5217,N_4616,N_4256);
nor U5218 (N_5218,N_4262,N_4615);
nor U5219 (N_5219,N_4574,N_4729);
or U5220 (N_5220,N_4072,N_4286);
or U5221 (N_5221,N_4672,N_4376);
or U5222 (N_5222,N_4665,N_4870);
and U5223 (N_5223,N_4125,N_4709);
nand U5224 (N_5224,N_4818,N_4012);
nand U5225 (N_5225,N_4986,N_4407);
or U5226 (N_5226,N_4273,N_4509);
nor U5227 (N_5227,N_4395,N_4759);
nor U5228 (N_5228,N_4936,N_4352);
and U5229 (N_5229,N_4628,N_4951);
or U5230 (N_5230,N_4827,N_4897);
nand U5231 (N_5231,N_4083,N_4728);
and U5232 (N_5232,N_4353,N_4394);
nor U5233 (N_5233,N_4859,N_4120);
nor U5234 (N_5234,N_4553,N_4904);
and U5235 (N_5235,N_4425,N_4860);
or U5236 (N_5236,N_4284,N_4719);
or U5237 (N_5237,N_4342,N_4171);
nand U5238 (N_5238,N_4057,N_4688);
nor U5239 (N_5239,N_4358,N_4905);
and U5240 (N_5240,N_4076,N_4941);
nor U5241 (N_5241,N_4006,N_4086);
nor U5242 (N_5242,N_4202,N_4417);
and U5243 (N_5243,N_4296,N_4093);
or U5244 (N_5244,N_4207,N_4791);
nor U5245 (N_5245,N_4164,N_4580);
or U5246 (N_5246,N_4835,N_4780);
or U5247 (N_5247,N_4255,N_4476);
nor U5248 (N_5248,N_4893,N_4801);
and U5249 (N_5249,N_4584,N_4669);
nor U5250 (N_5250,N_4204,N_4991);
and U5251 (N_5251,N_4340,N_4277);
nor U5252 (N_5252,N_4241,N_4211);
nor U5253 (N_5253,N_4738,N_4312);
or U5254 (N_5254,N_4771,N_4024);
or U5255 (N_5255,N_4623,N_4375);
nand U5256 (N_5256,N_4102,N_4344);
nand U5257 (N_5257,N_4409,N_4045);
nand U5258 (N_5258,N_4106,N_4011);
or U5259 (N_5259,N_4911,N_4963);
nor U5260 (N_5260,N_4337,N_4025);
and U5261 (N_5261,N_4463,N_4514);
or U5262 (N_5262,N_4235,N_4137);
or U5263 (N_5263,N_4199,N_4070);
and U5264 (N_5264,N_4330,N_4789);
nand U5265 (N_5265,N_4446,N_4451);
nor U5266 (N_5266,N_4401,N_4188);
nand U5267 (N_5267,N_4886,N_4146);
or U5268 (N_5268,N_4233,N_4251);
or U5269 (N_5269,N_4754,N_4089);
or U5270 (N_5270,N_4037,N_4319);
nor U5271 (N_5271,N_4107,N_4999);
or U5272 (N_5272,N_4804,N_4542);
nand U5273 (N_5273,N_4792,N_4567);
and U5274 (N_5274,N_4550,N_4614);
nand U5275 (N_5275,N_4726,N_4126);
and U5276 (N_5276,N_4856,N_4322);
or U5277 (N_5277,N_4965,N_4721);
nand U5278 (N_5278,N_4959,N_4822);
nand U5279 (N_5279,N_4228,N_4073);
and U5280 (N_5280,N_4046,N_4597);
and U5281 (N_5281,N_4208,N_4430);
nor U5282 (N_5282,N_4501,N_4848);
or U5283 (N_5283,N_4184,N_4625);
and U5284 (N_5284,N_4320,N_4981);
nor U5285 (N_5285,N_4943,N_4773);
nor U5286 (N_5286,N_4677,N_4530);
nor U5287 (N_5287,N_4784,N_4884);
nor U5288 (N_5288,N_4522,N_4282);
or U5289 (N_5289,N_4223,N_4960);
and U5290 (N_5290,N_4841,N_4473);
nor U5291 (N_5291,N_4795,N_4849);
and U5292 (N_5292,N_4156,N_4560);
and U5293 (N_5293,N_4488,N_4561);
and U5294 (N_5294,N_4763,N_4969);
nand U5295 (N_5295,N_4872,N_4415);
nor U5296 (N_5296,N_4898,N_4018);
nand U5297 (N_5297,N_4108,N_4599);
or U5298 (N_5298,N_4354,N_4497);
and U5299 (N_5299,N_4535,N_4000);
or U5300 (N_5300,N_4490,N_4254);
or U5301 (N_5301,N_4632,N_4664);
nand U5302 (N_5302,N_4449,N_4109);
nor U5303 (N_5303,N_4812,N_4739);
nand U5304 (N_5304,N_4984,N_4198);
and U5305 (N_5305,N_4062,N_4683);
or U5306 (N_5306,N_4815,N_4864);
or U5307 (N_5307,N_4504,N_4506);
nor U5308 (N_5308,N_4435,N_4659);
and U5309 (N_5309,N_4954,N_4351);
nand U5310 (N_5310,N_4633,N_4169);
or U5311 (N_5311,N_4603,N_4112);
nor U5312 (N_5312,N_4555,N_4248);
or U5313 (N_5313,N_4673,N_4148);
nand U5314 (N_5314,N_4588,N_4653);
and U5315 (N_5315,N_4950,N_4949);
nand U5316 (N_5316,N_4068,N_4467);
nor U5317 (N_5317,N_4014,N_4790);
nor U5318 (N_5318,N_4590,N_4947);
nor U5319 (N_5319,N_4661,N_4080);
and U5320 (N_5320,N_4464,N_4882);
nor U5321 (N_5321,N_4145,N_4307);
nor U5322 (N_5322,N_4532,N_4539);
nor U5323 (N_5323,N_4564,N_4380);
or U5324 (N_5324,N_4258,N_4636);
nor U5325 (N_5325,N_4508,N_4136);
nand U5326 (N_5326,N_4177,N_4527);
nor U5327 (N_5327,N_4662,N_4684);
nand U5328 (N_5328,N_4758,N_4772);
and U5329 (N_5329,N_4899,N_4499);
and U5330 (N_5330,N_4460,N_4129);
nor U5331 (N_5331,N_4021,N_4385);
or U5332 (N_5332,N_4418,N_4100);
or U5333 (N_5333,N_4459,N_4696);
nand U5334 (N_5334,N_4317,N_4649);
and U5335 (N_5335,N_4656,N_4693);
or U5336 (N_5336,N_4166,N_4915);
or U5337 (N_5337,N_4691,N_4304);
nand U5338 (N_5338,N_4022,N_4268);
or U5339 (N_5339,N_4760,N_4173);
nor U5340 (N_5340,N_4845,N_4581);
nor U5341 (N_5341,N_4231,N_4982);
nor U5342 (N_5342,N_4916,N_4935);
nor U5343 (N_5343,N_4201,N_4077);
or U5344 (N_5344,N_4657,N_4762);
or U5345 (N_5345,N_4627,N_4966);
and U5346 (N_5346,N_4302,N_4667);
or U5347 (N_5347,N_4280,N_4221);
nor U5348 (N_5348,N_4444,N_4387);
and U5349 (N_5349,N_4980,N_4644);
or U5350 (N_5350,N_4141,N_4468);
or U5351 (N_5351,N_4793,N_4880);
or U5352 (N_5352,N_4569,N_4159);
nand U5353 (N_5353,N_4537,N_4861);
and U5354 (N_5354,N_4013,N_4692);
xnor U5355 (N_5355,N_4655,N_4699);
or U5356 (N_5356,N_4576,N_4663);
nand U5357 (N_5357,N_4181,N_4745);
nand U5358 (N_5358,N_4140,N_4480);
nor U5359 (N_5359,N_4706,N_4583);
and U5360 (N_5360,N_4934,N_4816);
and U5361 (N_5361,N_4610,N_4139);
nand U5362 (N_5362,N_4458,N_4117);
nor U5363 (N_5363,N_4113,N_4456);
and U5364 (N_5364,N_4641,N_4328);
nand U5365 (N_5365,N_4349,N_4624);
nor U5366 (N_5366,N_4642,N_4498);
nand U5367 (N_5367,N_4519,N_4410);
nand U5368 (N_5368,N_4682,N_4047);
nand U5369 (N_5369,N_4413,N_4222);
nor U5370 (N_5370,N_4007,N_4405);
or U5371 (N_5371,N_4957,N_4646);
nor U5372 (N_5372,N_4925,N_4513);
nand U5373 (N_5373,N_4680,N_4855);
nor U5374 (N_5374,N_4920,N_4563);
nand U5375 (N_5375,N_4253,N_4618);
nor U5376 (N_5376,N_4087,N_4896);
nor U5377 (N_5377,N_4316,N_4647);
nor U5378 (N_5378,N_4350,N_4524);
or U5379 (N_5379,N_4035,N_4016);
nand U5380 (N_5380,N_4557,N_4518);
nor U5381 (N_5381,N_4592,N_4420);
nand U5382 (N_5382,N_4741,N_4178);
or U5383 (N_5383,N_4454,N_4339);
or U5384 (N_5384,N_4797,N_4929);
or U5385 (N_5385,N_4030,N_4543);
nor U5386 (N_5386,N_4411,N_4041);
nor U5387 (N_5387,N_4081,N_4167);
and U5388 (N_5388,N_4069,N_4323);
or U5389 (N_5389,N_4704,N_4685);
and U5390 (N_5390,N_4842,N_4877);
nand U5391 (N_5391,N_4453,N_4443);
or U5392 (N_5392,N_4426,N_4794);
and U5393 (N_5393,N_4336,N_4548);
or U5394 (N_5394,N_4367,N_4368);
nand U5395 (N_5395,N_4123,N_4939);
or U5396 (N_5396,N_4491,N_4591);
or U5397 (N_5397,N_4722,N_4232);
and U5398 (N_5398,N_4571,N_4868);
nand U5399 (N_5399,N_4798,N_4392);
nand U5400 (N_5400,N_4088,N_4853);
nor U5401 (N_5401,N_4265,N_4250);
and U5402 (N_5402,N_4054,N_4325);
nor U5403 (N_5403,N_4871,N_4863);
nor U5404 (N_5404,N_4289,N_4852);
nor U5405 (N_5405,N_4894,N_4619);
or U5406 (N_5406,N_4292,N_4711);
and U5407 (N_5407,N_4594,N_4496);
nand U5408 (N_5408,N_4033,N_4607);
and U5409 (N_5409,N_4731,N_4933);
nor U5410 (N_5410,N_4952,N_4922);
nand U5411 (N_5411,N_4111,N_4910);
and U5412 (N_5412,N_4750,N_4203);
or U5413 (N_5413,N_4155,N_4082);
or U5414 (N_5414,N_4028,N_4461);
nand U5415 (N_5415,N_4379,N_4263);
nor U5416 (N_5416,N_4810,N_4926);
and U5417 (N_5417,N_4210,N_4293);
or U5418 (N_5418,N_4829,N_4373);
or U5419 (N_5419,N_4658,N_4890);
and U5420 (N_5420,N_4585,N_4099);
nor U5421 (N_5421,N_4116,N_4727);
and U5422 (N_5422,N_4912,N_4384);
or U5423 (N_5423,N_4442,N_4869);
nor U5424 (N_5424,N_4879,N_4867);
and U5425 (N_5425,N_4471,N_4285);
nand U5426 (N_5426,N_4717,N_4224);
or U5427 (N_5427,N_4374,N_4528);
nor U5428 (N_5428,N_4098,N_4808);
nand U5429 (N_5429,N_4689,N_4832);
nor U5430 (N_5430,N_4609,N_4648);
nor U5431 (N_5431,N_4270,N_4052);
or U5432 (N_5432,N_4701,N_4216);
and U5433 (N_5433,N_4531,N_4994);
and U5434 (N_5434,N_4246,N_4445);
or U5435 (N_5435,N_4866,N_4055);
or U5436 (N_5436,N_4096,N_4686);
nor U5437 (N_5437,N_4976,N_4716);
and U5438 (N_5438,N_4906,N_4697);
nand U5439 (N_5439,N_4469,N_4500);
nand U5440 (N_5440,N_4153,N_4753);
and U5441 (N_5441,N_4313,N_4678);
nand U5442 (N_5442,N_4821,N_4796);
nand U5443 (N_5443,N_4288,N_4174);
or U5444 (N_5444,N_4733,N_4229);
nor U5445 (N_5445,N_4587,N_4670);
and U5446 (N_5446,N_4118,N_4834);
nor U5447 (N_5447,N_4278,N_4429);
or U5448 (N_5448,N_4604,N_4132);
or U5449 (N_5449,N_4010,N_4985);
nand U5450 (N_5450,N_4074,N_4249);
and U5451 (N_5451,N_4756,N_4287);
and U5452 (N_5452,N_4761,N_4507);
nor U5453 (N_5453,N_4299,N_4027);
nand U5454 (N_5454,N_4020,N_4274);
and U5455 (N_5455,N_4908,N_4511);
and U5456 (N_5456,N_4997,N_4742);
nor U5457 (N_5457,N_4259,N_4297);
nor U5458 (N_5458,N_4127,N_4837);
or U5459 (N_5459,N_4631,N_4900);
nor U5460 (N_5460,N_4058,N_4958);
and U5461 (N_5461,N_4874,N_4562);
nand U5462 (N_5462,N_4388,N_4103);
and U5463 (N_5463,N_4946,N_4290);
nor U5464 (N_5464,N_4452,N_4769);
and U5465 (N_5465,N_4332,N_4948);
nand U5466 (N_5466,N_4833,N_4558);
or U5467 (N_5467,N_4989,N_4311);
and U5468 (N_5468,N_4240,N_4707);
or U5469 (N_5469,N_4705,N_4079);
and U5470 (N_5470,N_4582,N_4972);
nor U5471 (N_5471,N_4257,N_4261);
nor U5472 (N_5472,N_4766,N_4749);
nor U5473 (N_5473,N_4838,N_4179);
or U5474 (N_5474,N_4163,N_4806);
and U5475 (N_5475,N_4485,N_4484);
nand U5476 (N_5476,N_4143,N_4424);
xor U5477 (N_5477,N_4674,N_4175);
nor U5478 (N_5478,N_4161,N_4909);
or U5479 (N_5479,N_4515,N_4406);
nor U5480 (N_5480,N_4510,N_4227);
nor U5481 (N_5481,N_4309,N_4305);
nand U5482 (N_5482,N_4601,N_4645);
and U5483 (N_5483,N_4700,N_4338);
nor U5484 (N_5484,N_4236,N_4324);
or U5485 (N_5485,N_4294,N_4061);
xor U5486 (N_5486,N_4383,N_4854);
nand U5487 (N_5487,N_4071,N_4315);
nor U5488 (N_5488,N_4857,N_4004);
nor U5489 (N_5489,N_4930,N_4064);
nor U5490 (N_5490,N_4450,N_4983);
nor U5491 (N_5491,N_4138,N_4973);
nor U5492 (N_5492,N_4301,N_4348);
or U5493 (N_5493,N_4566,N_4048);
or U5494 (N_5494,N_4279,N_4448);
or U5495 (N_5495,N_4990,N_4547);
nor U5496 (N_5496,N_4638,N_4660);
nor U5497 (N_5497,N_4923,N_4850);
nand U5498 (N_5498,N_4747,N_4234);
or U5499 (N_5499,N_4998,N_4399);
nand U5500 (N_5500,N_4889,N_4546);
and U5501 (N_5501,N_4657,N_4274);
and U5502 (N_5502,N_4779,N_4253);
nand U5503 (N_5503,N_4220,N_4887);
nand U5504 (N_5504,N_4811,N_4951);
nand U5505 (N_5505,N_4090,N_4270);
and U5506 (N_5506,N_4600,N_4418);
or U5507 (N_5507,N_4284,N_4006);
or U5508 (N_5508,N_4261,N_4847);
or U5509 (N_5509,N_4126,N_4353);
and U5510 (N_5510,N_4653,N_4039);
nor U5511 (N_5511,N_4981,N_4907);
and U5512 (N_5512,N_4622,N_4860);
and U5513 (N_5513,N_4346,N_4119);
nand U5514 (N_5514,N_4006,N_4178);
nand U5515 (N_5515,N_4238,N_4088);
nand U5516 (N_5516,N_4423,N_4119);
and U5517 (N_5517,N_4112,N_4937);
xnor U5518 (N_5518,N_4932,N_4580);
nand U5519 (N_5519,N_4702,N_4434);
nor U5520 (N_5520,N_4042,N_4234);
nand U5521 (N_5521,N_4555,N_4272);
nand U5522 (N_5522,N_4309,N_4264);
or U5523 (N_5523,N_4004,N_4834);
or U5524 (N_5524,N_4951,N_4831);
nand U5525 (N_5525,N_4306,N_4280);
and U5526 (N_5526,N_4231,N_4647);
and U5527 (N_5527,N_4067,N_4081);
or U5528 (N_5528,N_4922,N_4948);
or U5529 (N_5529,N_4180,N_4538);
and U5530 (N_5530,N_4240,N_4185);
and U5531 (N_5531,N_4519,N_4266);
or U5532 (N_5532,N_4561,N_4816);
nand U5533 (N_5533,N_4167,N_4511);
or U5534 (N_5534,N_4068,N_4103);
or U5535 (N_5535,N_4243,N_4542);
nor U5536 (N_5536,N_4344,N_4307);
or U5537 (N_5537,N_4855,N_4757);
nor U5538 (N_5538,N_4536,N_4493);
nor U5539 (N_5539,N_4585,N_4321);
or U5540 (N_5540,N_4447,N_4855);
or U5541 (N_5541,N_4034,N_4086);
and U5542 (N_5542,N_4349,N_4718);
or U5543 (N_5543,N_4720,N_4490);
nand U5544 (N_5544,N_4725,N_4123);
and U5545 (N_5545,N_4482,N_4306);
nor U5546 (N_5546,N_4311,N_4399);
nand U5547 (N_5547,N_4068,N_4966);
or U5548 (N_5548,N_4290,N_4574);
or U5549 (N_5549,N_4590,N_4219);
nor U5550 (N_5550,N_4146,N_4506);
nand U5551 (N_5551,N_4539,N_4552);
nand U5552 (N_5552,N_4402,N_4572);
and U5553 (N_5553,N_4473,N_4485);
nand U5554 (N_5554,N_4903,N_4737);
or U5555 (N_5555,N_4508,N_4882);
and U5556 (N_5556,N_4938,N_4507);
nor U5557 (N_5557,N_4467,N_4458);
or U5558 (N_5558,N_4428,N_4192);
or U5559 (N_5559,N_4042,N_4754);
nand U5560 (N_5560,N_4042,N_4701);
and U5561 (N_5561,N_4517,N_4904);
or U5562 (N_5562,N_4933,N_4376);
nand U5563 (N_5563,N_4771,N_4682);
nand U5564 (N_5564,N_4058,N_4395);
nor U5565 (N_5565,N_4568,N_4131);
nor U5566 (N_5566,N_4669,N_4883);
nand U5567 (N_5567,N_4017,N_4631);
and U5568 (N_5568,N_4171,N_4497);
and U5569 (N_5569,N_4866,N_4944);
nand U5570 (N_5570,N_4498,N_4062);
nand U5571 (N_5571,N_4865,N_4536);
and U5572 (N_5572,N_4336,N_4489);
or U5573 (N_5573,N_4708,N_4025);
nor U5574 (N_5574,N_4328,N_4512);
and U5575 (N_5575,N_4949,N_4657);
and U5576 (N_5576,N_4735,N_4201);
or U5577 (N_5577,N_4598,N_4224);
or U5578 (N_5578,N_4856,N_4066);
nor U5579 (N_5579,N_4969,N_4849);
nand U5580 (N_5580,N_4907,N_4234);
nand U5581 (N_5581,N_4501,N_4671);
nand U5582 (N_5582,N_4213,N_4274);
nor U5583 (N_5583,N_4956,N_4649);
or U5584 (N_5584,N_4143,N_4726);
nand U5585 (N_5585,N_4085,N_4552);
and U5586 (N_5586,N_4711,N_4004);
nand U5587 (N_5587,N_4253,N_4888);
and U5588 (N_5588,N_4958,N_4354);
nor U5589 (N_5589,N_4550,N_4069);
or U5590 (N_5590,N_4807,N_4594);
nand U5591 (N_5591,N_4083,N_4876);
and U5592 (N_5592,N_4555,N_4635);
nor U5593 (N_5593,N_4285,N_4668);
nor U5594 (N_5594,N_4583,N_4017);
and U5595 (N_5595,N_4157,N_4409);
and U5596 (N_5596,N_4524,N_4829);
and U5597 (N_5597,N_4004,N_4096);
nand U5598 (N_5598,N_4796,N_4512);
nor U5599 (N_5599,N_4325,N_4340);
or U5600 (N_5600,N_4510,N_4859);
nor U5601 (N_5601,N_4050,N_4589);
nor U5602 (N_5602,N_4429,N_4234);
or U5603 (N_5603,N_4502,N_4710);
nand U5604 (N_5604,N_4029,N_4220);
and U5605 (N_5605,N_4274,N_4288);
or U5606 (N_5606,N_4865,N_4672);
nor U5607 (N_5607,N_4979,N_4741);
or U5608 (N_5608,N_4110,N_4660);
and U5609 (N_5609,N_4354,N_4846);
and U5610 (N_5610,N_4931,N_4570);
or U5611 (N_5611,N_4965,N_4282);
or U5612 (N_5612,N_4745,N_4283);
or U5613 (N_5613,N_4401,N_4474);
nor U5614 (N_5614,N_4048,N_4267);
nand U5615 (N_5615,N_4424,N_4638);
or U5616 (N_5616,N_4149,N_4511);
nor U5617 (N_5617,N_4672,N_4120);
and U5618 (N_5618,N_4022,N_4590);
or U5619 (N_5619,N_4179,N_4334);
and U5620 (N_5620,N_4454,N_4315);
nand U5621 (N_5621,N_4047,N_4991);
or U5622 (N_5622,N_4325,N_4622);
nand U5623 (N_5623,N_4002,N_4439);
nand U5624 (N_5624,N_4249,N_4586);
and U5625 (N_5625,N_4391,N_4280);
nand U5626 (N_5626,N_4338,N_4850);
or U5627 (N_5627,N_4309,N_4318);
or U5628 (N_5628,N_4655,N_4914);
or U5629 (N_5629,N_4448,N_4410);
and U5630 (N_5630,N_4408,N_4510);
nor U5631 (N_5631,N_4334,N_4581);
and U5632 (N_5632,N_4284,N_4286);
or U5633 (N_5633,N_4945,N_4876);
nand U5634 (N_5634,N_4396,N_4657);
nand U5635 (N_5635,N_4137,N_4860);
and U5636 (N_5636,N_4424,N_4006);
nor U5637 (N_5637,N_4415,N_4884);
and U5638 (N_5638,N_4860,N_4187);
or U5639 (N_5639,N_4742,N_4241);
nor U5640 (N_5640,N_4924,N_4701);
nor U5641 (N_5641,N_4792,N_4183);
nand U5642 (N_5642,N_4040,N_4191);
or U5643 (N_5643,N_4559,N_4910);
nand U5644 (N_5644,N_4025,N_4925);
nor U5645 (N_5645,N_4286,N_4821);
and U5646 (N_5646,N_4282,N_4502);
nor U5647 (N_5647,N_4311,N_4832);
and U5648 (N_5648,N_4062,N_4272);
and U5649 (N_5649,N_4118,N_4435);
or U5650 (N_5650,N_4378,N_4391);
and U5651 (N_5651,N_4708,N_4050);
nand U5652 (N_5652,N_4425,N_4268);
nor U5653 (N_5653,N_4044,N_4683);
nor U5654 (N_5654,N_4358,N_4420);
nor U5655 (N_5655,N_4655,N_4648);
and U5656 (N_5656,N_4674,N_4828);
and U5657 (N_5657,N_4393,N_4182);
nand U5658 (N_5658,N_4600,N_4569);
or U5659 (N_5659,N_4153,N_4017);
nor U5660 (N_5660,N_4409,N_4896);
and U5661 (N_5661,N_4289,N_4128);
or U5662 (N_5662,N_4894,N_4309);
nand U5663 (N_5663,N_4362,N_4402);
or U5664 (N_5664,N_4305,N_4713);
and U5665 (N_5665,N_4048,N_4798);
nand U5666 (N_5666,N_4562,N_4618);
nor U5667 (N_5667,N_4581,N_4157);
or U5668 (N_5668,N_4540,N_4756);
nand U5669 (N_5669,N_4288,N_4381);
nand U5670 (N_5670,N_4804,N_4311);
nand U5671 (N_5671,N_4769,N_4365);
nand U5672 (N_5672,N_4964,N_4747);
nor U5673 (N_5673,N_4210,N_4515);
nor U5674 (N_5674,N_4401,N_4594);
nor U5675 (N_5675,N_4430,N_4570);
or U5676 (N_5676,N_4416,N_4595);
and U5677 (N_5677,N_4438,N_4885);
nand U5678 (N_5678,N_4418,N_4559);
and U5679 (N_5679,N_4797,N_4050);
or U5680 (N_5680,N_4430,N_4193);
nor U5681 (N_5681,N_4080,N_4405);
or U5682 (N_5682,N_4906,N_4246);
or U5683 (N_5683,N_4481,N_4411);
or U5684 (N_5684,N_4420,N_4253);
nor U5685 (N_5685,N_4252,N_4881);
nor U5686 (N_5686,N_4863,N_4392);
and U5687 (N_5687,N_4978,N_4964);
nor U5688 (N_5688,N_4473,N_4402);
nand U5689 (N_5689,N_4648,N_4704);
nor U5690 (N_5690,N_4068,N_4939);
or U5691 (N_5691,N_4986,N_4391);
nor U5692 (N_5692,N_4556,N_4570);
and U5693 (N_5693,N_4286,N_4084);
nand U5694 (N_5694,N_4791,N_4924);
xor U5695 (N_5695,N_4330,N_4900);
nor U5696 (N_5696,N_4446,N_4233);
nand U5697 (N_5697,N_4399,N_4855);
nand U5698 (N_5698,N_4804,N_4223);
nor U5699 (N_5699,N_4214,N_4380);
and U5700 (N_5700,N_4272,N_4013);
nand U5701 (N_5701,N_4984,N_4586);
nor U5702 (N_5702,N_4430,N_4079);
xnor U5703 (N_5703,N_4542,N_4580);
or U5704 (N_5704,N_4418,N_4952);
and U5705 (N_5705,N_4151,N_4267);
or U5706 (N_5706,N_4288,N_4850);
nor U5707 (N_5707,N_4580,N_4983);
and U5708 (N_5708,N_4729,N_4464);
nand U5709 (N_5709,N_4165,N_4661);
nor U5710 (N_5710,N_4817,N_4128);
nor U5711 (N_5711,N_4977,N_4007);
nand U5712 (N_5712,N_4228,N_4859);
nand U5713 (N_5713,N_4205,N_4318);
or U5714 (N_5714,N_4959,N_4125);
xor U5715 (N_5715,N_4054,N_4087);
and U5716 (N_5716,N_4327,N_4663);
nand U5717 (N_5717,N_4358,N_4768);
and U5718 (N_5718,N_4772,N_4675);
nor U5719 (N_5719,N_4071,N_4004);
nor U5720 (N_5720,N_4415,N_4977);
nor U5721 (N_5721,N_4200,N_4448);
or U5722 (N_5722,N_4133,N_4138);
nand U5723 (N_5723,N_4727,N_4003);
or U5724 (N_5724,N_4853,N_4830);
nand U5725 (N_5725,N_4038,N_4395);
nand U5726 (N_5726,N_4427,N_4344);
and U5727 (N_5727,N_4611,N_4980);
and U5728 (N_5728,N_4698,N_4158);
or U5729 (N_5729,N_4240,N_4719);
nand U5730 (N_5730,N_4698,N_4080);
nand U5731 (N_5731,N_4480,N_4394);
and U5732 (N_5732,N_4341,N_4701);
nand U5733 (N_5733,N_4004,N_4900);
and U5734 (N_5734,N_4271,N_4273);
nand U5735 (N_5735,N_4408,N_4037);
or U5736 (N_5736,N_4934,N_4144);
or U5737 (N_5737,N_4825,N_4984);
nand U5738 (N_5738,N_4848,N_4951);
nor U5739 (N_5739,N_4644,N_4511);
and U5740 (N_5740,N_4145,N_4366);
or U5741 (N_5741,N_4619,N_4782);
or U5742 (N_5742,N_4988,N_4966);
xor U5743 (N_5743,N_4710,N_4904);
and U5744 (N_5744,N_4572,N_4521);
or U5745 (N_5745,N_4413,N_4977);
and U5746 (N_5746,N_4856,N_4284);
nand U5747 (N_5747,N_4108,N_4489);
and U5748 (N_5748,N_4447,N_4790);
nand U5749 (N_5749,N_4314,N_4654);
and U5750 (N_5750,N_4730,N_4592);
nor U5751 (N_5751,N_4785,N_4067);
or U5752 (N_5752,N_4799,N_4150);
or U5753 (N_5753,N_4969,N_4158);
and U5754 (N_5754,N_4328,N_4546);
and U5755 (N_5755,N_4264,N_4733);
and U5756 (N_5756,N_4458,N_4680);
or U5757 (N_5757,N_4908,N_4859);
nand U5758 (N_5758,N_4858,N_4401);
and U5759 (N_5759,N_4309,N_4281);
and U5760 (N_5760,N_4171,N_4466);
nand U5761 (N_5761,N_4020,N_4252);
nand U5762 (N_5762,N_4464,N_4246);
nand U5763 (N_5763,N_4455,N_4338);
and U5764 (N_5764,N_4902,N_4133);
or U5765 (N_5765,N_4553,N_4689);
and U5766 (N_5766,N_4082,N_4068);
and U5767 (N_5767,N_4466,N_4307);
or U5768 (N_5768,N_4728,N_4508);
xnor U5769 (N_5769,N_4074,N_4552);
or U5770 (N_5770,N_4376,N_4956);
nor U5771 (N_5771,N_4648,N_4723);
nand U5772 (N_5772,N_4493,N_4449);
nor U5773 (N_5773,N_4804,N_4153);
nand U5774 (N_5774,N_4698,N_4094);
or U5775 (N_5775,N_4056,N_4680);
or U5776 (N_5776,N_4049,N_4087);
and U5777 (N_5777,N_4094,N_4245);
nor U5778 (N_5778,N_4720,N_4172);
and U5779 (N_5779,N_4230,N_4254);
and U5780 (N_5780,N_4042,N_4751);
or U5781 (N_5781,N_4539,N_4689);
xnor U5782 (N_5782,N_4871,N_4417);
and U5783 (N_5783,N_4442,N_4861);
or U5784 (N_5784,N_4986,N_4303);
or U5785 (N_5785,N_4030,N_4459);
nand U5786 (N_5786,N_4691,N_4273);
nor U5787 (N_5787,N_4770,N_4177);
nand U5788 (N_5788,N_4540,N_4957);
or U5789 (N_5789,N_4052,N_4426);
and U5790 (N_5790,N_4426,N_4352);
nor U5791 (N_5791,N_4452,N_4522);
nor U5792 (N_5792,N_4255,N_4021);
nand U5793 (N_5793,N_4245,N_4731);
or U5794 (N_5794,N_4654,N_4391);
and U5795 (N_5795,N_4399,N_4194);
or U5796 (N_5796,N_4997,N_4105);
nor U5797 (N_5797,N_4002,N_4082);
nor U5798 (N_5798,N_4693,N_4415);
nor U5799 (N_5799,N_4616,N_4315);
nor U5800 (N_5800,N_4770,N_4304);
nand U5801 (N_5801,N_4755,N_4664);
or U5802 (N_5802,N_4798,N_4351);
or U5803 (N_5803,N_4771,N_4930);
nor U5804 (N_5804,N_4645,N_4405);
nand U5805 (N_5805,N_4378,N_4633);
and U5806 (N_5806,N_4592,N_4311);
nand U5807 (N_5807,N_4491,N_4668);
or U5808 (N_5808,N_4498,N_4708);
or U5809 (N_5809,N_4316,N_4630);
nand U5810 (N_5810,N_4550,N_4133);
or U5811 (N_5811,N_4291,N_4639);
or U5812 (N_5812,N_4892,N_4987);
and U5813 (N_5813,N_4302,N_4602);
nor U5814 (N_5814,N_4176,N_4156);
and U5815 (N_5815,N_4093,N_4096);
and U5816 (N_5816,N_4194,N_4754);
nand U5817 (N_5817,N_4323,N_4423);
or U5818 (N_5818,N_4566,N_4162);
or U5819 (N_5819,N_4042,N_4848);
or U5820 (N_5820,N_4361,N_4002);
and U5821 (N_5821,N_4110,N_4191);
nand U5822 (N_5822,N_4051,N_4712);
nand U5823 (N_5823,N_4407,N_4060);
and U5824 (N_5824,N_4764,N_4425);
nor U5825 (N_5825,N_4209,N_4445);
nand U5826 (N_5826,N_4003,N_4426);
or U5827 (N_5827,N_4877,N_4264);
nor U5828 (N_5828,N_4089,N_4519);
nand U5829 (N_5829,N_4754,N_4793);
and U5830 (N_5830,N_4215,N_4863);
or U5831 (N_5831,N_4974,N_4984);
nand U5832 (N_5832,N_4415,N_4074);
nand U5833 (N_5833,N_4627,N_4022);
or U5834 (N_5834,N_4716,N_4540);
nor U5835 (N_5835,N_4196,N_4722);
nand U5836 (N_5836,N_4438,N_4894);
xnor U5837 (N_5837,N_4302,N_4099);
nor U5838 (N_5838,N_4242,N_4851);
or U5839 (N_5839,N_4887,N_4363);
and U5840 (N_5840,N_4634,N_4543);
nand U5841 (N_5841,N_4105,N_4296);
nor U5842 (N_5842,N_4554,N_4210);
and U5843 (N_5843,N_4480,N_4567);
and U5844 (N_5844,N_4275,N_4080);
and U5845 (N_5845,N_4199,N_4469);
or U5846 (N_5846,N_4176,N_4917);
nand U5847 (N_5847,N_4881,N_4985);
and U5848 (N_5848,N_4152,N_4757);
nor U5849 (N_5849,N_4308,N_4747);
and U5850 (N_5850,N_4808,N_4390);
or U5851 (N_5851,N_4743,N_4071);
nor U5852 (N_5852,N_4877,N_4365);
or U5853 (N_5853,N_4123,N_4921);
nor U5854 (N_5854,N_4716,N_4312);
nand U5855 (N_5855,N_4126,N_4404);
or U5856 (N_5856,N_4650,N_4461);
nand U5857 (N_5857,N_4857,N_4652);
or U5858 (N_5858,N_4472,N_4579);
or U5859 (N_5859,N_4816,N_4785);
and U5860 (N_5860,N_4460,N_4682);
or U5861 (N_5861,N_4929,N_4107);
and U5862 (N_5862,N_4844,N_4486);
or U5863 (N_5863,N_4840,N_4654);
or U5864 (N_5864,N_4074,N_4584);
nand U5865 (N_5865,N_4916,N_4992);
and U5866 (N_5866,N_4254,N_4828);
and U5867 (N_5867,N_4991,N_4373);
xnor U5868 (N_5868,N_4187,N_4364);
or U5869 (N_5869,N_4953,N_4799);
or U5870 (N_5870,N_4194,N_4154);
and U5871 (N_5871,N_4454,N_4228);
or U5872 (N_5872,N_4396,N_4551);
nor U5873 (N_5873,N_4289,N_4317);
or U5874 (N_5874,N_4728,N_4258);
or U5875 (N_5875,N_4513,N_4579);
or U5876 (N_5876,N_4661,N_4602);
or U5877 (N_5877,N_4812,N_4636);
or U5878 (N_5878,N_4351,N_4484);
nor U5879 (N_5879,N_4423,N_4640);
and U5880 (N_5880,N_4598,N_4483);
nand U5881 (N_5881,N_4708,N_4026);
nor U5882 (N_5882,N_4848,N_4745);
nor U5883 (N_5883,N_4994,N_4445);
nor U5884 (N_5884,N_4050,N_4087);
nor U5885 (N_5885,N_4522,N_4478);
xnor U5886 (N_5886,N_4747,N_4190);
nor U5887 (N_5887,N_4936,N_4455);
and U5888 (N_5888,N_4010,N_4827);
nor U5889 (N_5889,N_4562,N_4892);
nor U5890 (N_5890,N_4254,N_4518);
nor U5891 (N_5891,N_4877,N_4816);
or U5892 (N_5892,N_4884,N_4331);
nand U5893 (N_5893,N_4712,N_4638);
and U5894 (N_5894,N_4163,N_4598);
nor U5895 (N_5895,N_4586,N_4373);
nand U5896 (N_5896,N_4481,N_4818);
nor U5897 (N_5897,N_4990,N_4257);
or U5898 (N_5898,N_4338,N_4725);
and U5899 (N_5899,N_4562,N_4175);
or U5900 (N_5900,N_4698,N_4131);
and U5901 (N_5901,N_4341,N_4030);
or U5902 (N_5902,N_4164,N_4423);
nor U5903 (N_5903,N_4185,N_4514);
or U5904 (N_5904,N_4059,N_4863);
nor U5905 (N_5905,N_4114,N_4615);
or U5906 (N_5906,N_4284,N_4457);
nor U5907 (N_5907,N_4425,N_4343);
nand U5908 (N_5908,N_4878,N_4746);
and U5909 (N_5909,N_4499,N_4738);
nand U5910 (N_5910,N_4071,N_4543);
or U5911 (N_5911,N_4226,N_4986);
xnor U5912 (N_5912,N_4904,N_4618);
nand U5913 (N_5913,N_4114,N_4042);
and U5914 (N_5914,N_4569,N_4191);
or U5915 (N_5915,N_4280,N_4785);
xnor U5916 (N_5916,N_4480,N_4065);
or U5917 (N_5917,N_4450,N_4058);
or U5918 (N_5918,N_4908,N_4403);
nand U5919 (N_5919,N_4921,N_4170);
nand U5920 (N_5920,N_4747,N_4755);
or U5921 (N_5921,N_4818,N_4200);
nand U5922 (N_5922,N_4369,N_4617);
nor U5923 (N_5923,N_4660,N_4422);
nand U5924 (N_5924,N_4129,N_4337);
or U5925 (N_5925,N_4185,N_4847);
and U5926 (N_5926,N_4232,N_4889);
nand U5927 (N_5927,N_4987,N_4513);
nor U5928 (N_5928,N_4768,N_4996);
and U5929 (N_5929,N_4706,N_4816);
and U5930 (N_5930,N_4649,N_4630);
or U5931 (N_5931,N_4867,N_4988);
or U5932 (N_5932,N_4186,N_4229);
nand U5933 (N_5933,N_4482,N_4558);
nor U5934 (N_5934,N_4987,N_4238);
and U5935 (N_5935,N_4150,N_4189);
nor U5936 (N_5936,N_4942,N_4020);
nand U5937 (N_5937,N_4163,N_4560);
or U5938 (N_5938,N_4882,N_4967);
or U5939 (N_5939,N_4566,N_4977);
nor U5940 (N_5940,N_4610,N_4625);
nor U5941 (N_5941,N_4723,N_4852);
nand U5942 (N_5942,N_4655,N_4576);
nor U5943 (N_5943,N_4870,N_4649);
nor U5944 (N_5944,N_4363,N_4407);
nor U5945 (N_5945,N_4662,N_4100);
or U5946 (N_5946,N_4987,N_4350);
or U5947 (N_5947,N_4051,N_4984);
nor U5948 (N_5948,N_4324,N_4440);
and U5949 (N_5949,N_4633,N_4542);
and U5950 (N_5950,N_4990,N_4596);
nor U5951 (N_5951,N_4344,N_4998);
nand U5952 (N_5952,N_4106,N_4267);
nand U5953 (N_5953,N_4789,N_4384);
or U5954 (N_5954,N_4838,N_4665);
xnor U5955 (N_5955,N_4414,N_4333);
or U5956 (N_5956,N_4736,N_4688);
nor U5957 (N_5957,N_4556,N_4438);
and U5958 (N_5958,N_4543,N_4546);
nor U5959 (N_5959,N_4770,N_4466);
nand U5960 (N_5960,N_4578,N_4168);
or U5961 (N_5961,N_4192,N_4510);
nand U5962 (N_5962,N_4163,N_4158);
and U5963 (N_5963,N_4263,N_4683);
nor U5964 (N_5964,N_4517,N_4611);
nand U5965 (N_5965,N_4222,N_4000);
or U5966 (N_5966,N_4918,N_4045);
nand U5967 (N_5967,N_4081,N_4688);
nor U5968 (N_5968,N_4940,N_4442);
nand U5969 (N_5969,N_4510,N_4677);
nor U5970 (N_5970,N_4970,N_4155);
or U5971 (N_5971,N_4234,N_4667);
and U5972 (N_5972,N_4124,N_4310);
and U5973 (N_5973,N_4224,N_4462);
and U5974 (N_5974,N_4686,N_4076);
nor U5975 (N_5975,N_4509,N_4974);
nor U5976 (N_5976,N_4435,N_4859);
nand U5977 (N_5977,N_4491,N_4998);
or U5978 (N_5978,N_4014,N_4874);
nor U5979 (N_5979,N_4249,N_4722);
nor U5980 (N_5980,N_4751,N_4919);
nor U5981 (N_5981,N_4244,N_4443);
nand U5982 (N_5982,N_4886,N_4881);
nor U5983 (N_5983,N_4136,N_4148);
or U5984 (N_5984,N_4411,N_4955);
and U5985 (N_5985,N_4854,N_4639);
nor U5986 (N_5986,N_4598,N_4050);
nor U5987 (N_5987,N_4124,N_4905);
nand U5988 (N_5988,N_4604,N_4844);
nand U5989 (N_5989,N_4538,N_4331);
nor U5990 (N_5990,N_4032,N_4927);
or U5991 (N_5991,N_4153,N_4539);
and U5992 (N_5992,N_4548,N_4354);
and U5993 (N_5993,N_4128,N_4978);
nor U5994 (N_5994,N_4001,N_4535);
nor U5995 (N_5995,N_4468,N_4640);
xnor U5996 (N_5996,N_4372,N_4111);
nor U5997 (N_5997,N_4207,N_4923);
or U5998 (N_5998,N_4103,N_4545);
and U5999 (N_5999,N_4984,N_4890);
nand U6000 (N_6000,N_5297,N_5880);
nor U6001 (N_6001,N_5876,N_5820);
nand U6002 (N_6002,N_5281,N_5072);
nand U6003 (N_6003,N_5196,N_5200);
or U6004 (N_6004,N_5346,N_5197);
nand U6005 (N_6005,N_5728,N_5009);
nand U6006 (N_6006,N_5415,N_5039);
and U6007 (N_6007,N_5082,N_5012);
nand U6008 (N_6008,N_5267,N_5307);
nand U6009 (N_6009,N_5336,N_5738);
or U6010 (N_6010,N_5438,N_5428);
or U6011 (N_6011,N_5611,N_5688);
nor U6012 (N_6012,N_5277,N_5757);
and U6013 (N_6013,N_5450,N_5592);
nand U6014 (N_6014,N_5842,N_5984);
nor U6015 (N_6015,N_5961,N_5531);
nand U6016 (N_6016,N_5858,N_5520);
and U6017 (N_6017,N_5526,N_5478);
nor U6018 (N_6018,N_5373,N_5529);
or U6019 (N_6019,N_5476,N_5750);
or U6020 (N_6020,N_5989,N_5488);
and U6021 (N_6021,N_5691,N_5530);
and U6022 (N_6022,N_5953,N_5483);
and U6023 (N_6023,N_5209,N_5495);
or U6024 (N_6024,N_5033,N_5058);
nand U6025 (N_6025,N_5812,N_5958);
or U6026 (N_6026,N_5096,N_5440);
or U6027 (N_6027,N_5845,N_5223);
or U6028 (N_6028,N_5290,N_5952);
nand U6029 (N_6029,N_5780,N_5610);
or U6030 (N_6030,N_5258,N_5299);
or U6031 (N_6031,N_5005,N_5312);
and U6032 (N_6032,N_5800,N_5318);
nor U6033 (N_6033,N_5413,N_5316);
or U6034 (N_6034,N_5805,N_5322);
and U6035 (N_6035,N_5003,N_5525);
nand U6036 (N_6036,N_5455,N_5268);
nor U6037 (N_6037,N_5499,N_5252);
and U6038 (N_6038,N_5016,N_5519);
or U6039 (N_6039,N_5636,N_5090);
nand U6040 (N_6040,N_5212,N_5062);
and U6041 (N_6041,N_5954,N_5042);
or U6042 (N_6042,N_5945,N_5759);
nand U6043 (N_6043,N_5790,N_5020);
nor U6044 (N_6044,N_5872,N_5470);
nand U6045 (N_6045,N_5425,N_5421);
nand U6046 (N_6046,N_5128,N_5703);
nand U6047 (N_6047,N_5347,N_5816);
xnor U6048 (N_6048,N_5539,N_5881);
nor U6049 (N_6049,N_5768,N_5049);
nor U6050 (N_6050,N_5018,N_5202);
or U6051 (N_6051,N_5949,N_5515);
nand U6052 (N_6052,N_5206,N_5720);
nand U6053 (N_6053,N_5771,N_5753);
nor U6054 (N_6054,N_5030,N_5095);
nand U6055 (N_6055,N_5484,N_5325);
and U6056 (N_6056,N_5973,N_5433);
nor U6057 (N_6057,N_5372,N_5752);
and U6058 (N_6058,N_5356,N_5349);
and U6059 (N_6059,N_5376,N_5054);
and U6060 (N_6060,N_5809,N_5405);
nand U6061 (N_6061,N_5069,N_5060);
nor U6062 (N_6062,N_5195,N_5735);
nand U6063 (N_6063,N_5510,N_5137);
and U6064 (N_6064,N_5287,N_5660);
and U6065 (N_6065,N_5627,N_5622);
nand U6066 (N_6066,N_5852,N_5010);
or U6067 (N_6067,N_5679,N_5940);
nand U6068 (N_6068,N_5232,N_5092);
nor U6069 (N_6069,N_5417,N_5785);
nor U6070 (N_6070,N_5295,N_5004);
and U6071 (N_6071,N_5250,N_5723);
and U6072 (N_6072,N_5279,N_5310);
and U6073 (N_6073,N_5485,N_5221);
or U6074 (N_6074,N_5533,N_5065);
and U6075 (N_6075,N_5167,N_5762);
or U6076 (N_6076,N_5333,N_5112);
nand U6077 (N_6077,N_5794,N_5390);
and U6078 (N_6078,N_5630,N_5557);
or U6079 (N_6079,N_5225,N_5035);
or U6080 (N_6080,N_5199,N_5142);
or U6081 (N_6081,N_5150,N_5629);
and U6082 (N_6082,N_5183,N_5867);
nor U6083 (N_6083,N_5781,N_5001);
and U6084 (N_6084,N_5758,N_5754);
nor U6085 (N_6085,N_5644,N_5079);
nand U6086 (N_6086,N_5456,N_5542);
nor U6087 (N_6087,N_5791,N_5903);
or U6088 (N_6088,N_5409,N_5576);
nand U6089 (N_6089,N_5936,N_5987);
and U6090 (N_6090,N_5840,N_5761);
or U6091 (N_6091,N_5574,N_5094);
nor U6092 (N_6092,N_5102,N_5658);
nand U6093 (N_6093,N_5496,N_5220);
and U6094 (N_6094,N_5793,N_5523);
and U6095 (N_6095,N_5260,N_5229);
nor U6096 (N_6096,N_5383,N_5243);
nand U6097 (N_6097,N_5308,N_5700);
nor U6098 (N_6098,N_5399,N_5395);
nor U6099 (N_6099,N_5412,N_5912);
nor U6100 (N_6100,N_5806,N_5571);
nor U6101 (N_6101,N_5344,N_5974);
xor U6102 (N_6102,N_5481,N_5546);
nor U6103 (N_6103,N_5575,N_5222);
nor U6104 (N_6104,N_5437,N_5050);
and U6105 (N_6105,N_5655,N_5146);
nor U6106 (N_6106,N_5198,N_5391);
nor U6107 (N_6107,N_5013,N_5505);
and U6108 (N_6108,N_5898,N_5014);
nand U6109 (N_6109,N_5783,N_5901);
or U6110 (N_6110,N_5883,N_5751);
and U6111 (N_6111,N_5767,N_5219);
nor U6112 (N_6112,N_5578,N_5775);
nand U6113 (N_6113,N_5788,N_5797);
nand U6114 (N_6114,N_5602,N_5827);
and U6115 (N_6115,N_5733,N_5570);
or U6116 (N_6116,N_5321,N_5429);
and U6117 (N_6117,N_5593,N_5491);
or U6118 (N_6118,N_5676,N_5831);
nand U6119 (N_6119,N_5408,N_5273);
nor U6120 (N_6120,N_5911,N_5846);
and U6121 (N_6121,N_5628,N_5100);
nand U6122 (N_6122,N_5416,N_5897);
nor U6123 (N_6123,N_5895,N_5176);
and U6124 (N_6124,N_5148,N_5819);
nor U6125 (N_6125,N_5443,N_5763);
and U6126 (N_6126,N_5381,N_5214);
nand U6127 (N_6127,N_5853,N_5374);
or U6128 (N_6128,N_5259,N_5037);
nand U6129 (N_6129,N_5254,N_5657);
and U6130 (N_6130,N_5311,N_5185);
and U6131 (N_6131,N_5105,N_5215);
or U6132 (N_6132,N_5547,N_5830);
and U6133 (N_6133,N_5745,N_5847);
nand U6134 (N_6134,N_5778,N_5432);
nor U6135 (N_6135,N_5889,N_5015);
nand U6136 (N_6136,N_5908,N_5920);
nor U6137 (N_6137,N_5131,N_5040);
nor U6138 (N_6138,N_5303,N_5717);
or U6139 (N_6139,N_5048,N_5869);
or U6140 (N_6140,N_5704,N_5149);
or U6141 (N_6141,N_5471,N_5111);
nand U6142 (N_6142,N_5494,N_5969);
nor U6143 (N_6143,N_5888,N_5851);
and U6144 (N_6144,N_5482,N_5514);
or U6145 (N_6145,N_5130,N_5765);
and U6146 (N_6146,N_5850,N_5359);
xnor U6147 (N_6147,N_5586,N_5088);
nand U6148 (N_6148,N_5475,N_5139);
and U6149 (N_6149,N_5075,N_5388);
and U6150 (N_6150,N_5501,N_5103);
and U6151 (N_6151,N_5264,N_5216);
and U6152 (N_6152,N_5875,N_5906);
and U6153 (N_6153,N_5302,N_5330);
nor U6154 (N_6154,N_5580,N_5230);
nor U6155 (N_6155,N_5518,N_5122);
or U6156 (N_6156,N_5694,N_5191);
and U6157 (N_6157,N_5179,N_5726);
and U6158 (N_6158,N_5055,N_5357);
nand U6159 (N_6159,N_5787,N_5174);
or U6160 (N_6160,N_5600,N_5561);
and U6161 (N_6161,N_5737,N_5568);
and U6162 (N_6162,N_5887,N_5159);
nand U6163 (N_6163,N_5210,N_5451);
and U6164 (N_6164,N_5274,N_5948);
nand U6165 (N_6165,N_5564,N_5589);
and U6166 (N_6166,N_5832,N_5411);
and U6167 (N_6167,N_5234,N_5617);
nand U6168 (N_6168,N_5366,N_5782);
and U6169 (N_6169,N_5923,N_5052);
and U6170 (N_6170,N_5152,N_5272);
and U6171 (N_6171,N_5369,N_5528);
or U6172 (N_6172,N_5414,N_5459);
nor U6173 (N_6173,N_5296,N_5071);
and U6174 (N_6174,N_5991,N_5305);
nand U6175 (N_6175,N_5671,N_5235);
nor U6176 (N_6176,N_5022,N_5899);
nand U6177 (N_6177,N_5567,N_5021);
and U6178 (N_6178,N_5169,N_5692);
or U6179 (N_6179,N_5682,N_5626);
and U6180 (N_6180,N_5885,N_5687);
and U6181 (N_6181,N_5817,N_5674);
or U6182 (N_6182,N_5544,N_5201);
or U6183 (N_6183,N_5334,N_5160);
or U6184 (N_6184,N_5132,N_5172);
nand U6185 (N_6185,N_5400,N_5848);
and U6186 (N_6186,N_5749,N_5263);
and U6187 (N_6187,N_5224,N_5086);
nor U6188 (N_6188,N_5266,N_5620);
and U6189 (N_6189,N_5747,N_5449);
nor U6190 (N_6190,N_5981,N_5980);
nand U6191 (N_6191,N_5970,N_5882);
nor U6192 (N_6192,N_5862,N_5653);
or U6193 (N_6193,N_5615,N_5804);
and U6194 (N_6194,N_5545,N_5667);
nand U6195 (N_6195,N_5777,N_5217);
and U6196 (N_6196,N_5493,N_5916);
or U6197 (N_6197,N_5304,N_5032);
and U6198 (N_6198,N_5073,N_5659);
and U6199 (N_6199,N_5551,N_5354);
or U6200 (N_6200,N_5151,N_5382);
nor U6201 (N_6201,N_5384,N_5447);
and U6202 (N_6202,N_5902,N_5540);
nand U6203 (N_6203,N_5844,N_5686);
nor U6204 (N_6204,N_5672,N_5572);
nand U6205 (N_6205,N_5326,N_5007);
and U6206 (N_6206,N_5900,N_5314);
nand U6207 (N_6207,N_5826,N_5743);
nor U6208 (N_6208,N_5256,N_5070);
nor U6209 (N_6209,N_5925,N_5651);
or U6210 (N_6210,N_5943,N_5635);
and U6211 (N_6211,N_5158,N_5950);
nor U6212 (N_6212,N_5472,N_5722);
or U6213 (N_6213,N_5594,N_5975);
nor U6214 (N_6214,N_5255,N_5652);
nor U6215 (N_6215,N_5996,N_5716);
or U6216 (N_6216,N_5746,N_5978);
and U6217 (N_6217,N_5638,N_5238);
xor U6218 (N_6218,N_5410,N_5621);
nand U6219 (N_6219,N_5666,N_5824);
or U6220 (N_6220,N_5769,N_5664);
nor U6221 (N_6221,N_5119,N_5113);
or U6222 (N_6222,N_5959,N_5563);
or U6223 (N_6223,N_5890,N_5731);
and U6224 (N_6224,N_5623,N_5244);
or U6225 (N_6225,N_5080,N_5935);
nand U6226 (N_6226,N_5045,N_5527);
and U6227 (N_6227,N_5742,N_5632);
and U6228 (N_6228,N_5669,N_5982);
nand U6229 (N_6229,N_5927,N_5914);
nor U6230 (N_6230,N_5309,N_5907);
and U6231 (N_6231,N_5854,N_5964);
or U6232 (N_6232,N_5684,N_5998);
and U6233 (N_6233,N_5057,N_5891);
or U6234 (N_6234,N_5799,N_5327);
and U6235 (N_6235,N_5188,N_5587);
nand U6236 (N_6236,N_5841,N_5461);
or U6237 (N_6237,N_5596,N_5521);
and U6238 (N_6238,N_5207,N_5053);
and U6239 (N_6239,N_5170,N_5937);
and U6240 (N_6240,N_5083,N_5000);
nand U6241 (N_6241,N_5507,N_5795);
nand U6242 (N_6242,N_5813,N_5734);
or U6243 (N_6243,N_5145,N_5239);
or U6244 (N_6244,N_5324,N_5856);
nor U6245 (N_6245,N_5121,N_5690);
nor U6246 (N_6246,N_5041,N_5162);
nor U6247 (N_6247,N_5894,N_5051);
or U6248 (N_6248,N_5597,N_5941);
or U6249 (N_6249,N_5331,N_5656);
or U6250 (N_6250,N_5836,N_5504);
nor U6251 (N_6251,N_5956,N_5061);
and U6252 (N_6252,N_5386,N_5968);
nor U6253 (N_6253,N_5101,N_5559);
nor U6254 (N_6254,N_5426,N_5835);
or U6255 (N_6255,N_5802,N_5618);
nand U6256 (N_6256,N_5203,N_5161);
nor U6257 (N_6257,N_5689,N_5764);
nand U6258 (N_6258,N_5059,N_5960);
nor U6259 (N_6259,N_5859,N_5590);
xnor U6260 (N_6260,N_5965,N_5019);
and U6261 (N_6261,N_5915,N_5818);
nand U6262 (N_6262,N_5995,N_5718);
nand U6263 (N_6263,N_5419,N_5253);
or U6264 (N_6264,N_5976,N_5538);
and U6265 (N_6265,N_5967,N_5803);
and U6266 (N_6266,N_5601,N_5865);
or U6267 (N_6267,N_5343,N_5537);
nor U6268 (N_6268,N_5228,N_5227);
or U6269 (N_6269,N_5766,N_5192);
nand U6270 (N_6270,N_5573,N_5918);
or U6271 (N_6271,N_5289,N_5822);
and U6272 (N_6272,N_5427,N_5680);
nor U6273 (N_6273,N_5550,N_5994);
and U6274 (N_6274,N_5650,N_5190);
nor U6275 (N_6275,N_5106,N_5884);
nand U6276 (N_6276,N_5084,N_5946);
or U6277 (N_6277,N_5164,N_5140);
or U6278 (N_6278,N_5448,N_5467);
and U6279 (N_6279,N_5930,N_5077);
and U6280 (N_6280,N_5300,N_5839);
and U6281 (N_6281,N_5457,N_5099);
nor U6282 (N_6282,N_5487,N_5878);
nand U6283 (N_6283,N_5786,N_5023);
and U6284 (N_6284,N_5337,N_5270);
nand U6285 (N_6285,N_5284,N_5114);
nor U6286 (N_6286,N_5442,N_5934);
nor U6287 (N_6287,N_5760,N_5624);
nor U6288 (N_6288,N_5532,N_5193);
nor U6289 (N_6289,N_5631,N_5654);
or U6290 (N_6290,N_5008,N_5939);
or U6291 (N_6291,N_5246,N_5896);
or U6292 (N_6292,N_5002,N_5814);
nor U6293 (N_6293,N_5598,N_5988);
nand U6294 (N_6294,N_5834,N_5315);
nand U6295 (N_6295,N_5418,N_5251);
nand U6296 (N_6296,N_5933,N_5905);
nor U6297 (N_6297,N_5857,N_5707);
or U6298 (N_6298,N_5328,N_5047);
nand U6299 (N_6299,N_5497,N_5625);
and U6300 (N_6300,N_5719,N_5406);
nor U6301 (N_6301,N_5056,N_5770);
or U6302 (N_6302,N_5017,N_5157);
or U6303 (N_6303,N_5093,N_5541);
nor U6304 (N_6304,N_5715,N_5534);
nor U6305 (N_6305,N_5338,N_5074);
nor U6306 (N_6306,N_5298,N_5345);
nand U6307 (N_6307,N_5278,N_5599);
or U6308 (N_6308,N_5640,N_5508);
and U6309 (N_6309,N_5962,N_5569);
and U6310 (N_6310,N_5319,N_5189);
nor U6311 (N_6311,N_5466,N_5257);
or U6312 (N_6312,N_5031,N_5662);
nand U6313 (N_6313,N_5509,N_5892);
nand U6314 (N_6314,N_5683,N_5744);
or U6315 (N_6315,N_5917,N_5825);
or U6316 (N_6316,N_5739,N_5163);
nor U6317 (N_6317,N_5153,N_5725);
nor U6318 (N_6318,N_5705,N_5616);
nor U6319 (N_6319,N_5306,N_5365);
or U6320 (N_6320,N_5670,N_5932);
nand U6321 (N_6321,N_5585,N_5454);
nand U6322 (N_6322,N_5681,N_5706);
or U6323 (N_6323,N_5377,N_5389);
nor U6324 (N_6324,N_5614,N_5595);
nand U6325 (N_6325,N_5997,N_5696);
nand U6326 (N_6326,N_5125,N_5498);
nor U6327 (N_6327,N_5156,N_5554);
nor U6328 (N_6328,N_5489,N_5979);
and U6329 (N_6329,N_5942,N_5361);
nand U6330 (N_6330,N_5136,N_5972);
and U6331 (N_6331,N_5661,N_5133);
or U6332 (N_6332,N_5364,N_5603);
nor U6333 (N_6333,N_5643,N_5929);
nor U6334 (N_6334,N_5977,N_5067);
nand U6335 (N_6335,N_5261,N_5877);
nand U6336 (N_6336,N_5127,N_5604);
and U6337 (N_6337,N_5177,N_5313);
or U6338 (N_6338,N_5028,N_5126);
xor U6339 (N_6339,N_5473,N_5789);
and U6340 (N_6340,N_5773,N_5874);
nand U6341 (N_6341,N_5178,N_5713);
nor U6342 (N_6342,N_5807,N_5516);
nor U6343 (N_6343,N_5107,N_5011);
and U6344 (N_6344,N_5524,N_5194);
nor U6345 (N_6345,N_5171,N_5434);
nand U6346 (N_6346,N_5721,N_5556);
and U6347 (N_6347,N_5397,N_5135);
and U6348 (N_6348,N_5124,N_5063);
and U6349 (N_6349,N_5463,N_5709);
nor U6350 (N_6350,N_5317,N_5076);
and U6351 (N_6351,N_5291,N_5422);
nand U6352 (N_6352,N_5944,N_5245);
nor U6353 (N_6353,N_5549,N_5724);
and U6354 (N_6354,N_5535,N_5360);
or U6355 (N_6355,N_5605,N_5702);
nand U6356 (N_6356,N_5486,N_5469);
nor U6357 (N_6357,N_5120,N_5685);
and U6358 (N_6358,N_5971,N_5710);
and U6359 (N_6359,N_5218,N_5490);
or U6360 (N_6360,N_5606,N_5999);
nor U6361 (N_6361,N_5340,N_5144);
and U6362 (N_6362,N_5271,N_5168);
and U6363 (N_6363,N_5843,N_5465);
nand U6364 (N_6364,N_5211,N_5957);
and U6365 (N_6365,N_5341,N_5863);
nor U6366 (N_6366,N_5581,N_5714);
nand U6367 (N_6367,N_5026,N_5755);
nand U6368 (N_6368,N_5375,N_5134);
and U6369 (N_6369,N_5904,N_5861);
or U6370 (N_6370,N_5619,N_5184);
nor U6371 (N_6371,N_5784,N_5236);
and U6372 (N_6372,N_5029,N_5378);
nand U6373 (N_6373,N_5924,N_5821);
and U6374 (N_6374,N_5776,N_5612);
and U6375 (N_6375,N_5522,N_5849);
and U6376 (N_6376,N_5363,N_5503);
nand U6377 (N_6377,N_5548,N_5097);
nor U6378 (N_6378,N_5362,N_5729);
nor U6379 (N_6379,N_5241,N_5247);
nor U6380 (N_6380,N_5286,N_5452);
nor U6381 (N_6381,N_5024,N_5444);
or U6382 (N_6382,N_5992,N_5558);
or U6383 (N_6383,N_5801,N_5394);
and U6384 (N_6384,N_5909,N_5808);
nand U6385 (N_6385,N_5886,N_5129);
nand U6386 (N_6386,N_5913,N_5698);
or U6387 (N_6387,N_5637,N_5983);
nand U6388 (N_6388,N_5104,N_5648);
nor U6389 (N_6389,N_5693,N_5293);
and U6390 (N_6390,N_5108,N_5393);
nand U6391 (N_6391,N_5562,N_5633);
nor U6392 (N_6392,N_5921,N_5385);
or U6393 (N_6393,N_5458,N_5403);
nor U6394 (N_6394,N_5342,N_5282);
nand U6395 (N_6395,N_5085,N_5608);
nor U6396 (N_6396,N_5675,N_5828);
nand U6397 (N_6397,N_5237,N_5453);
nor U6398 (N_6398,N_5423,N_5701);
nand U6399 (N_6399,N_5955,N_5186);
nand U6400 (N_6400,N_5138,N_5928);
and U6401 (N_6401,N_5329,N_5552);
nor U6402 (N_6402,N_5323,N_5833);
nor U6403 (N_6403,N_5123,N_5985);
or U6404 (N_6404,N_5871,N_5175);
or U6405 (N_6405,N_5779,N_5371);
nor U6406 (N_6406,N_5205,N_5265);
and U6407 (N_6407,N_5634,N_5064);
and U6408 (N_6408,N_5430,N_5436);
nand U6409 (N_6409,N_5166,N_5280);
and U6410 (N_6410,N_5283,N_5294);
and U6411 (N_6411,N_5919,N_5368);
or U6412 (N_6412,N_5446,N_5736);
nor U6413 (N_6413,N_5512,N_5677);
nor U6414 (N_6414,N_5553,N_5838);
nor U6415 (N_6415,N_5240,N_5242);
or U6416 (N_6416,N_5091,N_5034);
and U6417 (N_6417,N_5098,N_5922);
nor U6418 (N_6418,N_5613,N_5046);
nand U6419 (N_6419,N_5798,N_5262);
or U6420 (N_6420,N_5639,N_5699);
or U6421 (N_6421,N_5609,N_5774);
or U6422 (N_6422,N_5380,N_5043);
or U6423 (N_6423,N_5500,N_5089);
nor U6424 (N_6424,N_5479,N_5647);
nor U6425 (N_6425,N_5320,N_5963);
nand U6426 (N_6426,N_5864,N_5301);
nand U6427 (N_6427,N_5868,N_5370);
nand U6428 (N_6428,N_5565,N_5511);
xor U6429 (N_6429,N_5431,N_5860);
nand U6430 (N_6430,N_5355,N_5815);
nand U6431 (N_6431,N_5645,N_5464);
nand U6432 (N_6432,N_5213,N_5543);
nand U6433 (N_6433,N_5811,N_5350);
nor U6434 (N_6434,N_5748,N_5044);
and U6435 (N_6435,N_5730,N_5352);
nand U6436 (N_6436,N_5335,N_5697);
nand U6437 (N_6437,N_5441,N_5555);
and U6438 (N_6438,N_5182,N_5025);
and U6439 (N_6439,N_5379,N_5292);
nand U6440 (N_6440,N_5741,N_5926);
or U6441 (N_6441,N_5480,N_5141);
nor U6442 (N_6442,N_5893,N_5087);
nor U6443 (N_6443,N_5460,N_5226);
nor U6444 (N_6444,N_5712,N_5560);
nand U6445 (N_6445,N_5285,N_5038);
nor U6446 (N_6446,N_5641,N_5339);
and U6447 (N_6447,N_5424,N_5866);
or U6448 (N_6448,N_5966,N_5387);
nand U6449 (N_6449,N_5154,N_5116);
and U6450 (N_6450,N_5506,N_5879);
or U6451 (N_6451,N_5036,N_5249);
nand U6452 (N_6452,N_5181,N_5649);
or U6453 (N_6453,N_5248,N_5204);
or U6454 (N_6454,N_5517,N_5792);
nor U6455 (N_6455,N_5358,N_5678);
nor U6456 (N_6456,N_5810,N_5947);
nor U6457 (N_6457,N_5269,N_5986);
nor U6458 (N_6458,N_5588,N_5439);
nor U6459 (N_6459,N_5231,N_5110);
nand U6460 (N_6460,N_5642,N_5027);
nand U6461 (N_6461,N_5993,N_5582);
nand U6462 (N_6462,N_5367,N_5165);
or U6463 (N_6463,N_5081,N_5756);
nand U6464 (N_6464,N_5829,N_5566);
nand U6465 (N_6465,N_5951,N_5663);
or U6466 (N_6466,N_5006,N_5396);
and U6467 (N_6467,N_5353,N_5492);
xnor U6468 (N_6468,N_5796,N_5173);
nor U6469 (N_6469,N_5646,N_5208);
or U6470 (N_6470,N_5584,N_5155);
nor U6471 (N_6471,N_5695,N_5477);
nand U6472 (N_6472,N_5579,N_5348);
nor U6473 (N_6473,N_5407,N_5583);
nor U6474 (N_6474,N_5740,N_5068);
and U6475 (N_6475,N_5332,N_5536);
and U6476 (N_6476,N_5435,N_5990);
and U6477 (N_6477,N_5727,N_5276);
and U6478 (N_6478,N_5931,N_5402);
nand U6479 (N_6479,N_5117,N_5474);
or U6480 (N_6480,N_5351,N_5577);
nor U6481 (N_6481,N_5115,N_5118);
and U6482 (N_6482,N_5938,N_5870);
or U6483 (N_6483,N_5502,N_5445);
nand U6484 (N_6484,N_5392,N_5665);
nor U6485 (N_6485,N_5513,N_5143);
and U6486 (N_6486,N_5147,N_5288);
and U6487 (N_6487,N_5708,N_5910);
or U6488 (N_6488,N_5420,N_5233);
nor U6489 (N_6489,N_5066,N_5673);
nor U6490 (N_6490,N_5668,N_5711);
or U6491 (N_6491,N_5823,N_5398);
or U6492 (N_6492,N_5187,N_5607);
and U6493 (N_6493,N_5732,N_5180);
or U6494 (N_6494,N_5468,N_5855);
or U6495 (N_6495,N_5837,N_5873);
and U6496 (N_6496,N_5772,N_5078);
nor U6497 (N_6497,N_5591,N_5462);
and U6498 (N_6498,N_5109,N_5275);
and U6499 (N_6499,N_5404,N_5401);
nand U6500 (N_6500,N_5036,N_5014);
or U6501 (N_6501,N_5680,N_5115);
or U6502 (N_6502,N_5952,N_5128);
and U6503 (N_6503,N_5223,N_5493);
nand U6504 (N_6504,N_5973,N_5580);
xnor U6505 (N_6505,N_5940,N_5413);
and U6506 (N_6506,N_5618,N_5799);
nor U6507 (N_6507,N_5487,N_5658);
nor U6508 (N_6508,N_5164,N_5980);
or U6509 (N_6509,N_5355,N_5105);
nand U6510 (N_6510,N_5099,N_5586);
and U6511 (N_6511,N_5584,N_5314);
and U6512 (N_6512,N_5621,N_5472);
nand U6513 (N_6513,N_5429,N_5648);
or U6514 (N_6514,N_5209,N_5867);
nor U6515 (N_6515,N_5509,N_5524);
or U6516 (N_6516,N_5976,N_5543);
nand U6517 (N_6517,N_5132,N_5966);
nor U6518 (N_6518,N_5607,N_5978);
or U6519 (N_6519,N_5068,N_5980);
or U6520 (N_6520,N_5128,N_5985);
nor U6521 (N_6521,N_5231,N_5162);
nor U6522 (N_6522,N_5768,N_5121);
nand U6523 (N_6523,N_5957,N_5365);
and U6524 (N_6524,N_5209,N_5611);
and U6525 (N_6525,N_5533,N_5951);
and U6526 (N_6526,N_5016,N_5940);
or U6527 (N_6527,N_5785,N_5013);
or U6528 (N_6528,N_5939,N_5035);
or U6529 (N_6529,N_5753,N_5406);
nand U6530 (N_6530,N_5163,N_5867);
nand U6531 (N_6531,N_5243,N_5011);
xnor U6532 (N_6532,N_5211,N_5852);
and U6533 (N_6533,N_5680,N_5446);
or U6534 (N_6534,N_5348,N_5210);
nand U6535 (N_6535,N_5681,N_5081);
nor U6536 (N_6536,N_5563,N_5195);
nand U6537 (N_6537,N_5175,N_5653);
or U6538 (N_6538,N_5151,N_5042);
or U6539 (N_6539,N_5817,N_5630);
and U6540 (N_6540,N_5776,N_5450);
nor U6541 (N_6541,N_5834,N_5002);
and U6542 (N_6542,N_5130,N_5243);
nand U6543 (N_6543,N_5933,N_5946);
nor U6544 (N_6544,N_5199,N_5748);
or U6545 (N_6545,N_5466,N_5744);
nor U6546 (N_6546,N_5629,N_5638);
nor U6547 (N_6547,N_5406,N_5122);
nand U6548 (N_6548,N_5522,N_5313);
nor U6549 (N_6549,N_5747,N_5654);
nor U6550 (N_6550,N_5699,N_5227);
or U6551 (N_6551,N_5271,N_5891);
and U6552 (N_6552,N_5156,N_5615);
nor U6553 (N_6553,N_5823,N_5577);
and U6554 (N_6554,N_5674,N_5851);
or U6555 (N_6555,N_5985,N_5589);
and U6556 (N_6556,N_5365,N_5908);
or U6557 (N_6557,N_5751,N_5720);
and U6558 (N_6558,N_5034,N_5060);
nor U6559 (N_6559,N_5840,N_5297);
nor U6560 (N_6560,N_5915,N_5254);
nor U6561 (N_6561,N_5856,N_5906);
or U6562 (N_6562,N_5502,N_5328);
nor U6563 (N_6563,N_5560,N_5136);
or U6564 (N_6564,N_5870,N_5813);
nand U6565 (N_6565,N_5811,N_5240);
nor U6566 (N_6566,N_5560,N_5228);
and U6567 (N_6567,N_5807,N_5728);
or U6568 (N_6568,N_5981,N_5145);
nor U6569 (N_6569,N_5124,N_5426);
nand U6570 (N_6570,N_5721,N_5195);
and U6571 (N_6571,N_5721,N_5468);
and U6572 (N_6572,N_5601,N_5838);
nor U6573 (N_6573,N_5787,N_5299);
nor U6574 (N_6574,N_5465,N_5341);
or U6575 (N_6575,N_5719,N_5085);
nand U6576 (N_6576,N_5434,N_5732);
nor U6577 (N_6577,N_5868,N_5200);
xor U6578 (N_6578,N_5121,N_5984);
or U6579 (N_6579,N_5737,N_5767);
and U6580 (N_6580,N_5595,N_5048);
and U6581 (N_6581,N_5051,N_5239);
nand U6582 (N_6582,N_5937,N_5563);
nor U6583 (N_6583,N_5273,N_5165);
and U6584 (N_6584,N_5452,N_5037);
nand U6585 (N_6585,N_5254,N_5504);
nor U6586 (N_6586,N_5889,N_5994);
nor U6587 (N_6587,N_5288,N_5314);
nor U6588 (N_6588,N_5826,N_5846);
nand U6589 (N_6589,N_5200,N_5703);
nor U6590 (N_6590,N_5015,N_5131);
and U6591 (N_6591,N_5456,N_5305);
or U6592 (N_6592,N_5357,N_5145);
nor U6593 (N_6593,N_5228,N_5145);
nand U6594 (N_6594,N_5003,N_5512);
and U6595 (N_6595,N_5058,N_5242);
nand U6596 (N_6596,N_5443,N_5788);
and U6597 (N_6597,N_5001,N_5239);
nor U6598 (N_6598,N_5984,N_5597);
nand U6599 (N_6599,N_5081,N_5354);
or U6600 (N_6600,N_5078,N_5038);
nor U6601 (N_6601,N_5846,N_5652);
nand U6602 (N_6602,N_5895,N_5172);
and U6603 (N_6603,N_5257,N_5637);
or U6604 (N_6604,N_5714,N_5861);
nor U6605 (N_6605,N_5129,N_5002);
nand U6606 (N_6606,N_5403,N_5333);
nand U6607 (N_6607,N_5380,N_5169);
nand U6608 (N_6608,N_5759,N_5768);
nor U6609 (N_6609,N_5418,N_5300);
nor U6610 (N_6610,N_5117,N_5297);
nand U6611 (N_6611,N_5644,N_5235);
nor U6612 (N_6612,N_5231,N_5234);
or U6613 (N_6613,N_5267,N_5334);
or U6614 (N_6614,N_5233,N_5134);
and U6615 (N_6615,N_5470,N_5572);
nor U6616 (N_6616,N_5487,N_5773);
and U6617 (N_6617,N_5652,N_5653);
or U6618 (N_6618,N_5775,N_5537);
and U6619 (N_6619,N_5988,N_5184);
and U6620 (N_6620,N_5213,N_5903);
or U6621 (N_6621,N_5520,N_5739);
and U6622 (N_6622,N_5512,N_5936);
and U6623 (N_6623,N_5123,N_5967);
or U6624 (N_6624,N_5725,N_5474);
nand U6625 (N_6625,N_5622,N_5361);
or U6626 (N_6626,N_5853,N_5456);
nor U6627 (N_6627,N_5005,N_5777);
nand U6628 (N_6628,N_5025,N_5518);
and U6629 (N_6629,N_5356,N_5404);
or U6630 (N_6630,N_5493,N_5529);
nand U6631 (N_6631,N_5206,N_5605);
nor U6632 (N_6632,N_5319,N_5256);
and U6633 (N_6633,N_5981,N_5550);
and U6634 (N_6634,N_5015,N_5314);
nand U6635 (N_6635,N_5192,N_5773);
or U6636 (N_6636,N_5422,N_5718);
or U6637 (N_6637,N_5819,N_5508);
and U6638 (N_6638,N_5230,N_5250);
nor U6639 (N_6639,N_5070,N_5112);
or U6640 (N_6640,N_5792,N_5646);
and U6641 (N_6641,N_5251,N_5211);
nand U6642 (N_6642,N_5685,N_5524);
nand U6643 (N_6643,N_5277,N_5006);
and U6644 (N_6644,N_5463,N_5689);
or U6645 (N_6645,N_5316,N_5341);
and U6646 (N_6646,N_5886,N_5045);
and U6647 (N_6647,N_5117,N_5615);
nand U6648 (N_6648,N_5332,N_5523);
nor U6649 (N_6649,N_5314,N_5388);
nor U6650 (N_6650,N_5427,N_5068);
and U6651 (N_6651,N_5190,N_5761);
nor U6652 (N_6652,N_5170,N_5925);
or U6653 (N_6653,N_5484,N_5800);
nor U6654 (N_6654,N_5737,N_5796);
and U6655 (N_6655,N_5093,N_5416);
nand U6656 (N_6656,N_5839,N_5560);
nand U6657 (N_6657,N_5482,N_5185);
and U6658 (N_6658,N_5349,N_5339);
and U6659 (N_6659,N_5623,N_5448);
nor U6660 (N_6660,N_5996,N_5102);
nor U6661 (N_6661,N_5669,N_5649);
nor U6662 (N_6662,N_5731,N_5203);
or U6663 (N_6663,N_5604,N_5042);
or U6664 (N_6664,N_5671,N_5930);
nor U6665 (N_6665,N_5283,N_5003);
nor U6666 (N_6666,N_5595,N_5906);
or U6667 (N_6667,N_5177,N_5655);
nor U6668 (N_6668,N_5906,N_5476);
nor U6669 (N_6669,N_5209,N_5001);
or U6670 (N_6670,N_5040,N_5654);
nor U6671 (N_6671,N_5193,N_5323);
or U6672 (N_6672,N_5531,N_5249);
and U6673 (N_6673,N_5943,N_5137);
nand U6674 (N_6674,N_5613,N_5509);
and U6675 (N_6675,N_5619,N_5618);
or U6676 (N_6676,N_5305,N_5500);
nand U6677 (N_6677,N_5625,N_5928);
and U6678 (N_6678,N_5888,N_5122);
nor U6679 (N_6679,N_5909,N_5757);
and U6680 (N_6680,N_5757,N_5730);
or U6681 (N_6681,N_5129,N_5902);
or U6682 (N_6682,N_5850,N_5342);
nor U6683 (N_6683,N_5987,N_5793);
nand U6684 (N_6684,N_5006,N_5665);
or U6685 (N_6685,N_5929,N_5863);
or U6686 (N_6686,N_5718,N_5450);
or U6687 (N_6687,N_5214,N_5997);
and U6688 (N_6688,N_5355,N_5714);
or U6689 (N_6689,N_5554,N_5214);
nand U6690 (N_6690,N_5231,N_5426);
nor U6691 (N_6691,N_5859,N_5094);
and U6692 (N_6692,N_5773,N_5296);
xor U6693 (N_6693,N_5672,N_5522);
nand U6694 (N_6694,N_5335,N_5497);
nand U6695 (N_6695,N_5924,N_5745);
and U6696 (N_6696,N_5813,N_5327);
and U6697 (N_6697,N_5480,N_5208);
and U6698 (N_6698,N_5567,N_5635);
or U6699 (N_6699,N_5434,N_5129);
nor U6700 (N_6700,N_5912,N_5471);
and U6701 (N_6701,N_5753,N_5437);
nand U6702 (N_6702,N_5533,N_5350);
nor U6703 (N_6703,N_5344,N_5075);
nor U6704 (N_6704,N_5892,N_5318);
nand U6705 (N_6705,N_5727,N_5161);
nor U6706 (N_6706,N_5418,N_5443);
nor U6707 (N_6707,N_5290,N_5769);
nor U6708 (N_6708,N_5910,N_5756);
nor U6709 (N_6709,N_5071,N_5264);
and U6710 (N_6710,N_5229,N_5569);
nand U6711 (N_6711,N_5048,N_5486);
and U6712 (N_6712,N_5486,N_5543);
or U6713 (N_6713,N_5169,N_5871);
or U6714 (N_6714,N_5369,N_5334);
xnor U6715 (N_6715,N_5202,N_5166);
nand U6716 (N_6716,N_5804,N_5063);
and U6717 (N_6717,N_5534,N_5012);
or U6718 (N_6718,N_5786,N_5765);
nand U6719 (N_6719,N_5383,N_5423);
nor U6720 (N_6720,N_5014,N_5369);
nand U6721 (N_6721,N_5598,N_5639);
nor U6722 (N_6722,N_5676,N_5320);
nor U6723 (N_6723,N_5622,N_5558);
nor U6724 (N_6724,N_5297,N_5250);
xor U6725 (N_6725,N_5229,N_5951);
or U6726 (N_6726,N_5447,N_5983);
and U6727 (N_6727,N_5909,N_5268);
nand U6728 (N_6728,N_5719,N_5853);
nand U6729 (N_6729,N_5758,N_5100);
nand U6730 (N_6730,N_5923,N_5738);
or U6731 (N_6731,N_5374,N_5573);
nor U6732 (N_6732,N_5992,N_5593);
nand U6733 (N_6733,N_5378,N_5967);
nor U6734 (N_6734,N_5323,N_5572);
or U6735 (N_6735,N_5528,N_5326);
nor U6736 (N_6736,N_5451,N_5787);
nor U6737 (N_6737,N_5865,N_5331);
and U6738 (N_6738,N_5980,N_5304);
nand U6739 (N_6739,N_5363,N_5483);
or U6740 (N_6740,N_5343,N_5236);
and U6741 (N_6741,N_5795,N_5423);
or U6742 (N_6742,N_5472,N_5228);
nor U6743 (N_6743,N_5215,N_5909);
and U6744 (N_6744,N_5064,N_5479);
nand U6745 (N_6745,N_5259,N_5322);
nand U6746 (N_6746,N_5069,N_5763);
nor U6747 (N_6747,N_5981,N_5506);
nor U6748 (N_6748,N_5165,N_5421);
or U6749 (N_6749,N_5860,N_5789);
and U6750 (N_6750,N_5259,N_5667);
nor U6751 (N_6751,N_5955,N_5290);
or U6752 (N_6752,N_5154,N_5684);
nand U6753 (N_6753,N_5647,N_5114);
nand U6754 (N_6754,N_5958,N_5622);
nor U6755 (N_6755,N_5323,N_5370);
nand U6756 (N_6756,N_5022,N_5645);
nor U6757 (N_6757,N_5787,N_5004);
or U6758 (N_6758,N_5479,N_5096);
and U6759 (N_6759,N_5999,N_5686);
nor U6760 (N_6760,N_5095,N_5017);
or U6761 (N_6761,N_5137,N_5863);
xor U6762 (N_6762,N_5057,N_5483);
nand U6763 (N_6763,N_5774,N_5302);
and U6764 (N_6764,N_5122,N_5157);
nand U6765 (N_6765,N_5049,N_5793);
nor U6766 (N_6766,N_5904,N_5795);
or U6767 (N_6767,N_5694,N_5276);
nand U6768 (N_6768,N_5798,N_5099);
and U6769 (N_6769,N_5510,N_5275);
and U6770 (N_6770,N_5819,N_5795);
and U6771 (N_6771,N_5121,N_5996);
nor U6772 (N_6772,N_5453,N_5424);
or U6773 (N_6773,N_5097,N_5796);
and U6774 (N_6774,N_5582,N_5173);
and U6775 (N_6775,N_5286,N_5134);
or U6776 (N_6776,N_5793,N_5383);
nor U6777 (N_6777,N_5985,N_5110);
or U6778 (N_6778,N_5233,N_5759);
nor U6779 (N_6779,N_5476,N_5046);
or U6780 (N_6780,N_5707,N_5053);
nand U6781 (N_6781,N_5246,N_5008);
nand U6782 (N_6782,N_5117,N_5505);
and U6783 (N_6783,N_5621,N_5875);
and U6784 (N_6784,N_5519,N_5073);
and U6785 (N_6785,N_5478,N_5981);
and U6786 (N_6786,N_5240,N_5267);
and U6787 (N_6787,N_5042,N_5959);
xor U6788 (N_6788,N_5984,N_5343);
nand U6789 (N_6789,N_5848,N_5807);
nand U6790 (N_6790,N_5913,N_5293);
nand U6791 (N_6791,N_5186,N_5254);
and U6792 (N_6792,N_5704,N_5844);
or U6793 (N_6793,N_5447,N_5696);
nand U6794 (N_6794,N_5302,N_5920);
nand U6795 (N_6795,N_5095,N_5180);
nor U6796 (N_6796,N_5769,N_5599);
and U6797 (N_6797,N_5226,N_5815);
and U6798 (N_6798,N_5358,N_5836);
xor U6799 (N_6799,N_5246,N_5743);
nand U6800 (N_6800,N_5981,N_5326);
nor U6801 (N_6801,N_5122,N_5042);
nand U6802 (N_6802,N_5289,N_5075);
nand U6803 (N_6803,N_5946,N_5768);
or U6804 (N_6804,N_5161,N_5584);
and U6805 (N_6805,N_5912,N_5800);
and U6806 (N_6806,N_5341,N_5682);
and U6807 (N_6807,N_5818,N_5094);
nor U6808 (N_6808,N_5296,N_5116);
or U6809 (N_6809,N_5640,N_5541);
and U6810 (N_6810,N_5420,N_5082);
nand U6811 (N_6811,N_5799,N_5796);
nor U6812 (N_6812,N_5372,N_5043);
and U6813 (N_6813,N_5497,N_5797);
and U6814 (N_6814,N_5128,N_5319);
or U6815 (N_6815,N_5504,N_5920);
nor U6816 (N_6816,N_5851,N_5787);
or U6817 (N_6817,N_5825,N_5489);
nor U6818 (N_6818,N_5173,N_5930);
nor U6819 (N_6819,N_5980,N_5348);
or U6820 (N_6820,N_5885,N_5033);
nor U6821 (N_6821,N_5559,N_5463);
nand U6822 (N_6822,N_5186,N_5474);
or U6823 (N_6823,N_5030,N_5992);
nand U6824 (N_6824,N_5577,N_5734);
nand U6825 (N_6825,N_5641,N_5945);
nand U6826 (N_6826,N_5501,N_5581);
and U6827 (N_6827,N_5615,N_5601);
nand U6828 (N_6828,N_5522,N_5512);
nor U6829 (N_6829,N_5421,N_5967);
or U6830 (N_6830,N_5929,N_5365);
nor U6831 (N_6831,N_5167,N_5115);
nand U6832 (N_6832,N_5018,N_5094);
nand U6833 (N_6833,N_5929,N_5734);
or U6834 (N_6834,N_5192,N_5065);
or U6835 (N_6835,N_5689,N_5220);
and U6836 (N_6836,N_5292,N_5397);
or U6837 (N_6837,N_5006,N_5744);
or U6838 (N_6838,N_5050,N_5208);
nor U6839 (N_6839,N_5844,N_5299);
nor U6840 (N_6840,N_5092,N_5853);
or U6841 (N_6841,N_5108,N_5436);
nand U6842 (N_6842,N_5481,N_5812);
nor U6843 (N_6843,N_5721,N_5129);
nor U6844 (N_6844,N_5705,N_5323);
nand U6845 (N_6845,N_5227,N_5889);
nand U6846 (N_6846,N_5277,N_5805);
or U6847 (N_6847,N_5947,N_5344);
nand U6848 (N_6848,N_5509,N_5904);
and U6849 (N_6849,N_5371,N_5519);
and U6850 (N_6850,N_5261,N_5595);
and U6851 (N_6851,N_5912,N_5049);
nand U6852 (N_6852,N_5186,N_5388);
nor U6853 (N_6853,N_5529,N_5149);
nor U6854 (N_6854,N_5420,N_5845);
or U6855 (N_6855,N_5734,N_5605);
nor U6856 (N_6856,N_5382,N_5239);
nand U6857 (N_6857,N_5577,N_5009);
and U6858 (N_6858,N_5566,N_5421);
nand U6859 (N_6859,N_5168,N_5282);
or U6860 (N_6860,N_5992,N_5741);
or U6861 (N_6861,N_5965,N_5297);
nor U6862 (N_6862,N_5914,N_5404);
or U6863 (N_6863,N_5942,N_5466);
or U6864 (N_6864,N_5783,N_5366);
nand U6865 (N_6865,N_5773,N_5815);
and U6866 (N_6866,N_5102,N_5423);
nor U6867 (N_6867,N_5317,N_5016);
nor U6868 (N_6868,N_5255,N_5490);
and U6869 (N_6869,N_5082,N_5971);
or U6870 (N_6870,N_5853,N_5592);
and U6871 (N_6871,N_5051,N_5013);
nand U6872 (N_6872,N_5675,N_5289);
nor U6873 (N_6873,N_5693,N_5561);
or U6874 (N_6874,N_5813,N_5857);
and U6875 (N_6875,N_5202,N_5448);
or U6876 (N_6876,N_5585,N_5738);
nand U6877 (N_6877,N_5313,N_5058);
or U6878 (N_6878,N_5196,N_5894);
or U6879 (N_6879,N_5020,N_5349);
nor U6880 (N_6880,N_5920,N_5747);
xnor U6881 (N_6881,N_5645,N_5015);
nor U6882 (N_6882,N_5308,N_5254);
or U6883 (N_6883,N_5154,N_5077);
and U6884 (N_6884,N_5630,N_5848);
or U6885 (N_6885,N_5853,N_5397);
nand U6886 (N_6886,N_5340,N_5567);
nor U6887 (N_6887,N_5219,N_5122);
nor U6888 (N_6888,N_5933,N_5476);
or U6889 (N_6889,N_5318,N_5424);
nand U6890 (N_6890,N_5354,N_5419);
nand U6891 (N_6891,N_5463,N_5208);
and U6892 (N_6892,N_5557,N_5442);
and U6893 (N_6893,N_5113,N_5681);
and U6894 (N_6894,N_5647,N_5966);
and U6895 (N_6895,N_5435,N_5170);
nand U6896 (N_6896,N_5207,N_5826);
or U6897 (N_6897,N_5592,N_5811);
or U6898 (N_6898,N_5308,N_5365);
and U6899 (N_6899,N_5893,N_5716);
nand U6900 (N_6900,N_5134,N_5094);
nor U6901 (N_6901,N_5995,N_5593);
and U6902 (N_6902,N_5748,N_5530);
or U6903 (N_6903,N_5090,N_5084);
and U6904 (N_6904,N_5393,N_5494);
nand U6905 (N_6905,N_5056,N_5174);
nand U6906 (N_6906,N_5682,N_5842);
nor U6907 (N_6907,N_5133,N_5595);
nor U6908 (N_6908,N_5721,N_5404);
or U6909 (N_6909,N_5217,N_5214);
or U6910 (N_6910,N_5975,N_5903);
or U6911 (N_6911,N_5928,N_5113);
nand U6912 (N_6912,N_5596,N_5019);
nor U6913 (N_6913,N_5161,N_5223);
nor U6914 (N_6914,N_5675,N_5357);
nand U6915 (N_6915,N_5301,N_5941);
and U6916 (N_6916,N_5527,N_5838);
and U6917 (N_6917,N_5250,N_5262);
nor U6918 (N_6918,N_5978,N_5693);
and U6919 (N_6919,N_5087,N_5697);
nor U6920 (N_6920,N_5242,N_5490);
nand U6921 (N_6921,N_5384,N_5317);
nand U6922 (N_6922,N_5425,N_5949);
or U6923 (N_6923,N_5617,N_5430);
and U6924 (N_6924,N_5238,N_5477);
or U6925 (N_6925,N_5231,N_5915);
nor U6926 (N_6926,N_5696,N_5518);
nand U6927 (N_6927,N_5793,N_5398);
nand U6928 (N_6928,N_5489,N_5329);
and U6929 (N_6929,N_5106,N_5771);
nor U6930 (N_6930,N_5578,N_5099);
or U6931 (N_6931,N_5233,N_5113);
and U6932 (N_6932,N_5947,N_5614);
and U6933 (N_6933,N_5097,N_5438);
and U6934 (N_6934,N_5166,N_5698);
nor U6935 (N_6935,N_5964,N_5322);
nand U6936 (N_6936,N_5898,N_5977);
nand U6937 (N_6937,N_5593,N_5085);
or U6938 (N_6938,N_5576,N_5249);
and U6939 (N_6939,N_5077,N_5003);
and U6940 (N_6940,N_5665,N_5149);
nor U6941 (N_6941,N_5516,N_5763);
nor U6942 (N_6942,N_5015,N_5564);
nor U6943 (N_6943,N_5616,N_5167);
nand U6944 (N_6944,N_5920,N_5977);
nor U6945 (N_6945,N_5915,N_5452);
and U6946 (N_6946,N_5646,N_5279);
nor U6947 (N_6947,N_5336,N_5050);
and U6948 (N_6948,N_5641,N_5469);
and U6949 (N_6949,N_5422,N_5387);
nor U6950 (N_6950,N_5043,N_5408);
nor U6951 (N_6951,N_5192,N_5224);
and U6952 (N_6952,N_5492,N_5796);
nand U6953 (N_6953,N_5609,N_5518);
nor U6954 (N_6954,N_5042,N_5486);
or U6955 (N_6955,N_5825,N_5480);
or U6956 (N_6956,N_5370,N_5993);
nor U6957 (N_6957,N_5345,N_5251);
and U6958 (N_6958,N_5514,N_5938);
and U6959 (N_6959,N_5022,N_5185);
or U6960 (N_6960,N_5707,N_5127);
nand U6961 (N_6961,N_5464,N_5587);
and U6962 (N_6962,N_5787,N_5809);
nor U6963 (N_6963,N_5101,N_5261);
nand U6964 (N_6964,N_5574,N_5478);
nor U6965 (N_6965,N_5749,N_5297);
or U6966 (N_6966,N_5205,N_5806);
and U6967 (N_6967,N_5965,N_5705);
nand U6968 (N_6968,N_5031,N_5524);
nor U6969 (N_6969,N_5812,N_5260);
nand U6970 (N_6970,N_5990,N_5253);
or U6971 (N_6971,N_5662,N_5075);
and U6972 (N_6972,N_5389,N_5807);
or U6973 (N_6973,N_5251,N_5124);
and U6974 (N_6974,N_5952,N_5108);
or U6975 (N_6975,N_5681,N_5958);
or U6976 (N_6976,N_5644,N_5770);
nor U6977 (N_6977,N_5024,N_5771);
and U6978 (N_6978,N_5582,N_5064);
nor U6979 (N_6979,N_5053,N_5035);
and U6980 (N_6980,N_5056,N_5452);
or U6981 (N_6981,N_5654,N_5585);
nor U6982 (N_6982,N_5397,N_5072);
nand U6983 (N_6983,N_5269,N_5215);
xor U6984 (N_6984,N_5748,N_5290);
nor U6985 (N_6985,N_5972,N_5452);
nor U6986 (N_6986,N_5696,N_5797);
nand U6987 (N_6987,N_5897,N_5901);
nand U6988 (N_6988,N_5346,N_5409);
nor U6989 (N_6989,N_5384,N_5950);
or U6990 (N_6990,N_5307,N_5592);
or U6991 (N_6991,N_5587,N_5760);
nand U6992 (N_6992,N_5311,N_5298);
nor U6993 (N_6993,N_5993,N_5715);
or U6994 (N_6994,N_5699,N_5724);
nand U6995 (N_6995,N_5904,N_5917);
xor U6996 (N_6996,N_5882,N_5967);
nor U6997 (N_6997,N_5507,N_5255);
nor U6998 (N_6998,N_5209,N_5712);
nor U6999 (N_6999,N_5085,N_5330);
nor U7000 (N_7000,N_6967,N_6758);
nand U7001 (N_7001,N_6998,N_6172);
nor U7002 (N_7002,N_6466,N_6954);
or U7003 (N_7003,N_6706,N_6960);
nand U7004 (N_7004,N_6043,N_6997);
nand U7005 (N_7005,N_6500,N_6638);
nand U7006 (N_7006,N_6124,N_6527);
or U7007 (N_7007,N_6881,N_6114);
and U7008 (N_7008,N_6193,N_6574);
or U7009 (N_7009,N_6417,N_6957);
and U7010 (N_7010,N_6811,N_6641);
nor U7011 (N_7011,N_6864,N_6838);
xnor U7012 (N_7012,N_6244,N_6129);
or U7013 (N_7013,N_6693,N_6478);
and U7014 (N_7014,N_6137,N_6982);
nor U7015 (N_7015,N_6068,N_6661);
and U7016 (N_7016,N_6804,N_6782);
nand U7017 (N_7017,N_6635,N_6825);
and U7018 (N_7018,N_6475,N_6840);
or U7019 (N_7019,N_6090,N_6945);
nand U7020 (N_7020,N_6057,N_6007);
xor U7021 (N_7021,N_6666,N_6927);
nand U7022 (N_7022,N_6257,N_6887);
nor U7023 (N_7023,N_6824,N_6353);
and U7024 (N_7024,N_6367,N_6792);
nor U7025 (N_7025,N_6710,N_6085);
or U7026 (N_7026,N_6951,N_6676);
and U7027 (N_7027,N_6533,N_6276);
nand U7028 (N_7028,N_6911,N_6769);
nand U7029 (N_7029,N_6664,N_6182);
nor U7030 (N_7030,N_6802,N_6272);
nor U7031 (N_7031,N_6070,N_6657);
and U7032 (N_7032,N_6966,N_6465);
nand U7033 (N_7033,N_6322,N_6499);
nand U7034 (N_7034,N_6262,N_6397);
nor U7035 (N_7035,N_6695,N_6235);
nand U7036 (N_7036,N_6368,N_6698);
or U7037 (N_7037,N_6819,N_6246);
nor U7038 (N_7038,N_6827,N_6469);
and U7039 (N_7039,N_6471,N_6513);
and U7040 (N_7040,N_6948,N_6569);
nor U7041 (N_7041,N_6504,N_6071);
nand U7042 (N_7042,N_6249,N_6134);
or U7043 (N_7043,N_6680,N_6509);
or U7044 (N_7044,N_6535,N_6364);
nand U7045 (N_7045,N_6391,N_6679);
and U7046 (N_7046,N_6521,N_6107);
and U7047 (N_7047,N_6485,N_6697);
and U7048 (N_7048,N_6362,N_6100);
and U7049 (N_7049,N_6320,N_6946);
nor U7050 (N_7050,N_6361,N_6280);
or U7051 (N_7051,N_6601,N_6645);
nand U7052 (N_7052,N_6221,N_6999);
and U7053 (N_7053,N_6739,N_6433);
or U7054 (N_7054,N_6561,N_6772);
and U7055 (N_7055,N_6563,N_6347);
or U7056 (N_7056,N_6776,N_6315);
nand U7057 (N_7057,N_6744,N_6801);
nor U7058 (N_7058,N_6095,N_6024);
or U7059 (N_7059,N_6806,N_6269);
or U7060 (N_7060,N_6783,N_6577);
nor U7061 (N_7061,N_6786,N_6628);
and U7062 (N_7062,N_6926,N_6143);
nand U7063 (N_7063,N_6828,N_6356);
and U7064 (N_7064,N_6295,N_6943);
or U7065 (N_7065,N_6876,N_6463);
and U7066 (N_7066,N_6459,N_6903);
nand U7067 (N_7067,N_6299,N_6472);
and U7068 (N_7068,N_6492,N_6524);
and U7069 (N_7069,N_6899,N_6120);
or U7070 (N_7070,N_6436,N_6343);
or U7071 (N_7071,N_6800,N_6649);
nor U7072 (N_7072,N_6117,N_6968);
nand U7073 (N_7073,N_6460,N_6684);
nor U7074 (N_7074,N_6534,N_6282);
or U7075 (N_7075,N_6423,N_6742);
and U7076 (N_7076,N_6201,N_6757);
and U7077 (N_7077,N_6467,N_6351);
nand U7078 (N_7078,N_6089,N_6302);
nand U7079 (N_7079,N_6750,N_6022);
nand U7080 (N_7080,N_6001,N_6528);
or U7081 (N_7081,N_6025,N_6133);
or U7082 (N_7082,N_6588,N_6452);
nand U7083 (N_7083,N_6583,N_6634);
nor U7084 (N_7084,N_6181,N_6456);
nand U7085 (N_7085,N_6484,N_6369);
nand U7086 (N_7086,N_6755,N_6650);
and U7087 (N_7087,N_6516,N_6377);
and U7088 (N_7088,N_6681,N_6329);
nand U7089 (N_7089,N_6690,N_6974);
nand U7090 (N_7090,N_6489,N_6217);
or U7091 (N_7091,N_6596,N_6342);
or U7092 (N_7092,N_6514,N_6384);
nor U7093 (N_7093,N_6863,N_6875);
or U7094 (N_7094,N_6425,N_6510);
and U7095 (N_7095,N_6430,N_6422);
nand U7096 (N_7096,N_6765,N_6242);
and U7097 (N_7097,N_6613,N_6185);
nand U7098 (N_7098,N_6200,N_6515);
and U7099 (N_7099,N_6046,N_6402);
and U7100 (N_7100,N_6556,N_6570);
or U7101 (N_7101,N_6206,N_6701);
and U7102 (N_7102,N_6223,N_6495);
and U7103 (N_7103,N_6247,N_6625);
nor U7104 (N_7104,N_6788,N_6157);
and U7105 (N_7105,N_6880,N_6713);
or U7106 (N_7106,N_6985,N_6851);
and U7107 (N_7107,N_6216,N_6891);
and U7108 (N_7108,N_6905,N_6831);
nor U7109 (N_7109,N_6944,N_6033);
or U7110 (N_7110,N_6300,N_6953);
nand U7111 (N_7111,N_6963,N_6077);
and U7112 (N_7112,N_6021,N_6624);
or U7113 (N_7113,N_6405,N_6284);
and U7114 (N_7114,N_6365,N_6759);
or U7115 (N_7115,N_6198,N_6842);
nand U7116 (N_7116,N_6580,N_6894);
nand U7117 (N_7117,N_6323,N_6623);
and U7118 (N_7118,N_6155,N_6050);
nor U7119 (N_7119,N_6862,N_6526);
and U7120 (N_7120,N_6752,N_6018);
and U7121 (N_7121,N_6297,N_6626);
nor U7122 (N_7122,N_6633,N_6308);
or U7123 (N_7123,N_6063,N_6052);
nand U7124 (N_7124,N_6565,N_6131);
nand U7125 (N_7125,N_6861,N_6464);
nand U7126 (N_7126,N_6969,N_6871);
nand U7127 (N_7127,N_6820,N_6303);
or U7128 (N_7128,N_6075,N_6823);
and U7129 (N_7129,N_6670,N_6034);
or U7130 (N_7130,N_6537,N_6003);
nand U7131 (N_7131,N_6784,N_6956);
or U7132 (N_7132,N_6686,N_6258);
and U7133 (N_7133,N_6164,N_6045);
xnor U7134 (N_7134,N_6689,N_6311);
nand U7135 (N_7135,N_6251,N_6011);
nor U7136 (N_7136,N_6376,N_6448);
and U7137 (N_7137,N_6403,N_6176);
or U7138 (N_7138,N_6371,N_6918);
or U7139 (N_7139,N_6180,N_6008);
nor U7140 (N_7140,N_6379,N_6844);
nor U7141 (N_7141,N_6572,N_6126);
nand U7142 (N_7142,N_6073,N_6672);
nor U7143 (N_7143,N_6506,N_6614);
nor U7144 (N_7144,N_6408,N_6768);
and U7145 (N_7145,N_6138,N_6644);
nand U7146 (N_7146,N_6910,N_6330);
nand U7147 (N_7147,N_6058,N_6546);
or U7148 (N_7148,N_6543,N_6812);
and U7149 (N_7149,N_6445,N_6805);
nor U7150 (N_7150,N_6976,N_6219);
or U7151 (N_7151,N_6971,N_6410);
nor U7152 (N_7152,N_6290,N_6890);
nor U7153 (N_7153,N_6798,N_6699);
nand U7154 (N_7154,N_6518,N_6162);
and U7155 (N_7155,N_6813,N_6988);
and U7156 (N_7156,N_6947,N_6069);
or U7157 (N_7157,N_6540,N_6105);
nand U7158 (N_7158,N_6908,N_6762);
nor U7159 (N_7159,N_6749,N_6333);
nand U7160 (N_7160,N_6076,N_6677);
nand U7161 (N_7161,N_6933,N_6035);
or U7162 (N_7162,N_6421,N_6026);
nand U7163 (N_7163,N_6177,N_6632);
and U7164 (N_7164,N_6121,N_6847);
or U7165 (N_7165,N_6643,N_6923);
nand U7166 (N_7166,N_6196,N_6738);
nor U7167 (N_7167,N_6959,N_6846);
nand U7168 (N_7168,N_6902,N_6617);
nand U7169 (N_7169,N_6538,N_6156);
and U7170 (N_7170,N_6934,N_6132);
or U7171 (N_7171,N_6080,N_6413);
nand U7172 (N_7172,N_6158,N_6883);
or U7173 (N_7173,N_6065,N_6525);
nor U7174 (N_7174,N_6064,N_6396);
nor U7175 (N_7175,N_6724,N_6150);
and U7176 (N_7176,N_6288,N_6836);
nand U7177 (N_7177,N_6858,N_6503);
and U7178 (N_7178,N_6594,N_6748);
and U7179 (N_7179,N_6019,N_6291);
nand U7180 (N_7180,N_6669,N_6931);
or U7181 (N_7181,N_6111,N_6253);
and U7182 (N_7182,N_6938,N_6327);
or U7183 (N_7183,N_6787,N_6639);
or U7184 (N_7184,N_6979,N_6778);
and U7185 (N_7185,N_6366,N_6834);
nor U7186 (N_7186,N_6455,N_6047);
nand U7187 (N_7187,N_6659,N_6312);
or U7188 (N_7188,N_6989,N_6213);
or U7189 (N_7189,N_6882,N_6897);
or U7190 (N_7190,N_6508,N_6383);
and U7191 (N_7191,N_6093,N_6994);
or U7192 (N_7192,N_6273,N_6208);
or U7193 (N_7193,N_6381,N_6568);
nand U7194 (N_7194,N_6239,N_6675);
and U7195 (N_7195,N_6919,N_6855);
nor U7196 (N_7196,N_6854,N_6474);
nor U7197 (N_7197,N_6061,N_6874);
and U7198 (N_7198,N_6852,N_6865);
and U7199 (N_7199,N_6160,N_6547);
nand U7200 (N_7200,N_6892,N_6306);
and U7201 (N_7201,N_6372,N_6562);
nor U7202 (N_7202,N_6000,N_6937);
and U7203 (N_7203,N_6993,N_6390);
nand U7204 (N_7204,N_6404,N_6502);
and U7205 (N_7205,N_6289,N_6990);
nand U7206 (N_7206,N_6554,N_6551);
or U7207 (N_7207,N_6142,N_6996);
nand U7208 (N_7208,N_6780,N_6431);
nand U7209 (N_7209,N_6231,N_6777);
nor U7210 (N_7210,N_6764,N_6074);
nor U7211 (N_7211,N_6557,N_6924);
or U7212 (N_7212,N_6833,N_6737);
nor U7213 (N_7213,N_6274,N_6298);
or U7214 (N_7214,N_6728,N_6210);
nor U7215 (N_7215,N_6346,N_6708);
or U7216 (N_7216,N_6277,N_6536);
nand U7217 (N_7217,N_6860,N_6037);
nor U7218 (N_7218,N_6191,N_6331);
nor U7219 (N_7219,N_6378,N_6393);
nor U7220 (N_7220,N_6420,N_6382);
nor U7221 (N_7221,N_6889,N_6949);
or U7222 (N_7222,N_6939,N_6775);
or U7223 (N_7223,N_6779,N_6730);
and U7224 (N_7224,N_6726,N_6721);
or U7225 (N_7225,N_6714,N_6961);
nand U7226 (N_7226,N_6548,N_6853);
nand U7227 (N_7227,N_6694,N_6211);
nor U7228 (N_7228,N_6468,N_6496);
or U7229 (N_7229,N_6224,N_6461);
and U7230 (N_7230,N_6770,N_6581);
and U7231 (N_7231,N_6116,N_6549);
or U7232 (N_7232,N_6349,N_6481);
or U7233 (N_7233,N_6148,N_6906);
or U7234 (N_7234,N_6789,N_6491);
nor U7235 (N_7235,N_6444,N_6088);
nor U7236 (N_7236,N_6795,N_6900);
and U7237 (N_7237,N_6578,N_6663);
nor U7238 (N_7238,N_6305,N_6531);
and U7239 (N_7239,N_6809,N_6530);
and U7240 (N_7240,N_6817,N_6703);
nand U7241 (N_7241,N_6187,N_6281);
or U7242 (N_7242,N_6980,N_6793);
nor U7243 (N_7243,N_6041,N_6119);
and U7244 (N_7244,N_6341,N_6539);
nand U7245 (N_7245,N_6363,N_6715);
and U7246 (N_7246,N_6983,N_6743);
and U7247 (N_7247,N_6579,N_6204);
and U7248 (N_7248,N_6110,N_6886);
and U7249 (N_7249,N_6673,N_6048);
nand U7250 (N_7250,N_6595,N_6559);
nand U7251 (N_7251,N_6720,N_6582);
or U7252 (N_7252,N_6409,N_6810);
nand U7253 (N_7253,N_6407,N_6821);
nand U7254 (N_7254,N_6773,N_6416);
and U7255 (N_7255,N_6942,N_6428);
nand U7256 (N_7256,N_6166,N_6760);
and U7257 (N_7257,N_6986,N_6727);
nand U7258 (N_7258,N_6197,N_6081);
nand U7259 (N_7259,N_6375,N_6108);
or U7260 (N_7260,N_6352,N_6978);
nor U7261 (N_7261,N_6292,N_6092);
nor U7262 (N_7262,N_6031,N_6012);
and U7263 (N_7263,N_6955,N_6103);
or U7264 (N_7264,N_6925,N_6631);
nor U7265 (N_7265,N_6051,N_6912);
or U7266 (N_7266,N_6140,N_6324);
and U7267 (N_7267,N_6036,N_6279);
nand U7268 (N_7268,N_6104,N_6896);
nand U7269 (N_7269,N_6808,N_6683);
nor U7270 (N_7270,N_6794,N_6545);
nand U7271 (N_7271,N_6866,N_6053);
or U7272 (N_7272,N_6096,N_6822);
xor U7273 (N_7273,N_6294,N_6437);
and U7274 (N_7274,N_6358,N_6552);
nand U7275 (N_7275,N_6700,N_6418);
or U7276 (N_7276,N_6640,N_6154);
or U7277 (N_7277,N_6236,N_6973);
nor U7278 (N_7278,N_6250,N_6040);
or U7279 (N_7279,N_6380,N_6885);
and U7280 (N_7280,N_6682,N_6932);
nor U7281 (N_7281,N_6179,N_6328);
nand U7282 (N_7282,N_6627,N_6020);
nand U7283 (N_7283,N_6992,N_6656);
or U7284 (N_7284,N_6774,N_6141);
nand U7285 (N_7285,N_6230,N_6411);
nor U7286 (N_7286,N_6754,N_6803);
and U7287 (N_7287,N_6270,N_6275);
nand U7288 (N_7288,N_6214,N_6790);
and U7289 (N_7289,N_6458,N_6203);
nand U7290 (N_7290,N_6360,N_6194);
and U7291 (N_7291,N_6149,N_6082);
or U7292 (N_7292,N_6002,N_6152);
or U7293 (N_7293,N_6245,N_6086);
xor U7294 (N_7294,N_6286,N_6135);
or U7295 (N_7295,N_6442,N_6326);
or U7296 (N_7296,N_6029,N_6667);
nand U7297 (N_7297,N_6869,N_6220);
nand U7298 (N_7298,N_6835,N_6977);
nand U7299 (N_7299,N_6332,N_6237);
or U7300 (N_7300,N_6147,N_6845);
nor U7301 (N_7301,N_6712,N_6486);
xor U7302 (N_7302,N_6373,N_6567);
nor U7303 (N_7303,N_6161,N_6056);
nand U7304 (N_7304,N_6856,N_6113);
nor U7305 (N_7305,N_6564,N_6006);
nand U7306 (N_7306,N_6928,N_6254);
nor U7307 (N_7307,N_6094,N_6427);
nand U7308 (N_7308,N_6734,N_6317);
nor U7309 (N_7309,N_6443,N_6573);
or U7310 (N_7310,N_6265,N_6125);
nor U7311 (N_7311,N_6914,N_6599);
or U7312 (N_7312,N_6898,N_6370);
and U7313 (N_7313,N_6604,N_6316);
nand U7314 (N_7314,N_6023,N_6941);
nor U7315 (N_7315,N_6243,N_6654);
and U7316 (N_7316,N_6587,N_6517);
nor U7317 (N_7317,N_6202,N_6646);
nand U7318 (N_7318,N_6450,N_6873);
nor U7319 (N_7319,N_6717,N_6584);
or U7320 (N_7320,N_6271,N_6153);
and U7321 (N_7321,N_6532,N_6877);
nand U7322 (N_7322,N_6745,N_6339);
nor U7323 (N_7323,N_6916,N_6529);
or U7324 (N_7324,N_6446,N_6816);
and U7325 (N_7325,N_6174,N_6477);
or U7326 (N_7326,N_6746,N_6060);
nand U7327 (N_7327,N_6505,N_6586);
and U7328 (N_7328,N_6122,N_6618);
or U7329 (N_7329,N_6837,N_6385);
or U7330 (N_7330,N_6732,N_6839);
or U7331 (N_7331,N_6829,N_6662);
nand U7332 (N_7332,N_6066,N_6207);
nor U7333 (N_7333,N_6340,N_6260);
or U7334 (N_7334,N_6415,N_6039);
and U7335 (N_7335,N_6814,N_6435);
and U7336 (N_7336,N_6167,N_6612);
nor U7337 (N_7337,N_6238,N_6815);
nand U7338 (N_7338,N_6336,N_6304);
or U7339 (N_7339,N_6542,N_6611);
or U7340 (N_7340,N_6042,N_6597);
and U7341 (N_7341,N_6929,N_6169);
nand U7342 (N_7342,N_6118,N_6849);
nor U7343 (N_7343,N_6962,N_6130);
or U7344 (N_7344,N_6589,N_6653);
and U7345 (N_7345,N_6479,N_6620);
and U7346 (N_7346,N_6429,N_6044);
nor U7347 (N_7347,N_6190,N_6619);
or U7348 (N_7348,N_6921,N_6936);
or U7349 (N_7349,N_6602,N_6259);
or U7350 (N_7350,N_6451,N_6175);
and U7351 (N_7351,N_6884,N_6241);
and U7352 (N_7352,N_6761,N_6622);
nor U7353 (N_7353,N_6796,N_6310);
nand U7354 (N_7354,N_6389,N_6665);
and U7355 (N_7355,N_6189,N_6541);
nor U7356 (N_7356,N_6763,N_6171);
and U7357 (N_7357,N_6867,N_6395);
nor U7358 (N_7358,N_6482,N_6859);
nand U7359 (N_7359,N_6248,N_6084);
nor U7360 (N_7360,N_6637,N_6857);
nand U7361 (N_7361,N_6733,N_6054);
nand U7362 (N_7362,N_6412,N_6909);
or U7363 (N_7363,N_6711,N_6462);
or U7364 (N_7364,N_6480,N_6032);
or U7365 (N_7365,N_6687,N_6826);
nor U7366 (N_7366,N_6401,N_6128);
nor U7367 (N_7367,N_6483,N_6605);
nand U7368 (N_7368,N_6392,N_6544);
nand U7369 (N_7369,N_6497,N_6359);
nor U7370 (N_7370,N_6498,N_6419);
nand U7371 (N_7371,N_6374,N_6205);
and U7372 (N_7372,N_6512,N_6165);
and U7373 (N_7373,N_6729,N_6751);
and U7374 (N_7374,N_6178,N_6671);
nand U7375 (N_7375,N_6691,N_6736);
nand U7376 (N_7376,N_6832,N_6170);
nand U7377 (N_7377,N_6807,N_6901);
nor U7378 (N_7378,N_6747,N_6293);
and U7379 (N_7379,N_6441,N_6072);
nand U7380 (N_7380,N_6922,N_6571);
and U7381 (N_7381,N_6964,N_6766);
nand U7382 (N_7382,N_6872,N_6685);
and U7383 (N_7383,N_6501,N_6227);
and U7384 (N_7384,N_6457,N_6144);
or U7385 (N_7385,N_6655,N_6426);
nand U7386 (N_7386,N_6799,N_6593);
nand U7387 (N_7387,N_6240,N_6895);
nor U7388 (N_7388,N_6127,N_6688);
nor U7389 (N_7389,N_6350,N_6476);
and U7390 (N_7390,N_6097,N_6266);
or U7391 (N_7391,N_6719,N_6355);
nor U7392 (N_7392,N_6432,N_6079);
nor U7393 (N_7393,N_6606,N_6030);
nand U7394 (N_7394,N_6309,N_6283);
or U7395 (N_7395,N_6600,N_6186);
nor U7396 (N_7396,N_6753,N_6307);
nand U7397 (N_7397,N_6091,N_6106);
nand U7398 (N_7398,N_6038,N_6668);
or U7399 (N_7399,N_6674,N_6731);
or U7400 (N_7400,N_6984,N_6652);
nand U7401 (N_7401,N_6893,N_6314);
nor U7402 (N_7402,N_6139,N_6215);
nor U7403 (N_7403,N_6005,N_6608);
and U7404 (N_7404,N_6232,N_6168);
nand U7405 (N_7405,N_6439,N_6335);
nor U7406 (N_7406,N_6488,N_6028);
or U7407 (N_7407,N_6915,N_6658);
nand U7408 (N_7408,N_6558,N_6692);
and U7409 (N_7409,N_6083,N_6490);
or U7410 (N_7410,N_6725,N_6609);
or U7411 (N_7411,N_6981,N_6566);
and U7412 (N_7412,N_6940,N_6229);
nand U7413 (N_7413,N_6263,N_6267);
nor U7414 (N_7414,N_6145,N_6015);
or U7415 (N_7415,N_6398,N_6354);
nor U7416 (N_7416,N_6621,N_6301);
nand U7417 (N_7417,N_6049,N_6319);
nand U7418 (N_7418,N_6440,N_6878);
nand U7419 (N_7419,N_6325,N_6192);
or U7420 (N_7420,N_6473,N_6337);
nand U7421 (N_7421,N_6630,N_6101);
or U7422 (N_7422,N_6348,N_6102);
xor U7423 (N_7423,N_6087,N_6519);
and U7424 (N_7424,N_6592,N_6183);
or U7425 (N_7425,N_6470,N_6453);
nor U7426 (N_7426,N_6287,N_6321);
and U7427 (N_7427,N_6560,N_6722);
nand U7428 (N_7428,N_6151,N_6424);
nor U7429 (N_7429,N_6590,N_6704);
nor U7430 (N_7430,N_6705,N_6907);
or U7431 (N_7431,N_6702,N_6678);
nor U7432 (N_7432,N_6013,N_6222);
and U7433 (N_7433,N_6136,N_6781);
nand U7434 (N_7434,N_6226,N_6062);
nand U7435 (N_7435,N_6059,N_6791);
nand U7436 (N_7436,N_6109,N_6709);
or U7437 (N_7437,N_6888,N_6576);
or U7438 (N_7438,N_6209,N_6555);
and U7439 (N_7439,N_6987,N_6507);
nand U7440 (N_7440,N_6598,N_6648);
nand U7441 (N_7441,N_6841,N_6920);
and U7442 (N_7442,N_6647,N_6264);
nand U7443 (N_7443,N_6636,N_6487);
or U7444 (N_7444,N_6017,N_6009);
nand U7445 (N_7445,N_6188,N_6660);
nor U7446 (N_7446,N_6146,N_6256);
nand U7447 (N_7447,N_6818,N_6112);
nand U7448 (N_7448,N_6318,N_6741);
nor U7449 (N_7449,N_6591,N_6848);
nand U7450 (N_7450,N_6184,N_6523);
nor U7451 (N_7451,N_6233,N_6494);
or U7452 (N_7452,N_6386,N_6735);
nand U7453 (N_7453,N_6952,N_6913);
and U7454 (N_7454,N_6707,N_6740);
and U7455 (N_7455,N_6607,N_6406);
nand U7456 (N_7456,N_6970,N_6930);
nand U7457 (N_7457,N_6313,N_6991);
nand U7458 (N_7458,N_6522,N_6278);
nand U7459 (N_7459,N_6629,N_6447);
and U7460 (N_7460,N_6357,N_6575);
or U7461 (N_7461,N_6255,N_6234);
nand U7462 (N_7462,N_6268,N_6716);
or U7463 (N_7463,N_6449,N_6718);
or U7464 (N_7464,N_6159,N_6218);
and U7465 (N_7465,N_6261,N_6553);
nor U7466 (N_7466,N_6195,N_6123);
nand U7467 (N_7467,N_6723,N_6163);
nor U7468 (N_7468,N_6603,N_6642);
nor U7469 (N_7469,N_6388,N_6399);
nand U7470 (N_7470,N_6225,N_6334);
nor U7471 (N_7471,N_6338,N_6756);
or U7472 (N_7472,N_6616,N_6414);
nand U7473 (N_7473,N_6965,N_6434);
or U7474 (N_7474,N_6585,N_6870);
and U7475 (N_7475,N_6078,N_6868);
nand U7476 (N_7476,N_6975,N_6055);
nand U7477 (N_7477,N_6493,N_6771);
nor U7478 (N_7478,N_6016,N_6879);
or U7479 (N_7479,N_6610,N_6830);
and U7480 (N_7480,N_6520,N_6252);
nor U7481 (N_7481,N_6935,N_6173);
nand U7482 (N_7482,N_6067,N_6696);
nand U7483 (N_7483,N_6285,N_6843);
nor U7484 (N_7484,N_6850,N_6651);
or U7485 (N_7485,N_6115,N_6972);
xor U7486 (N_7486,N_6615,N_6345);
and U7487 (N_7487,N_6904,N_6212);
and U7488 (N_7488,N_6785,N_6454);
and U7489 (N_7489,N_6098,N_6995);
nand U7490 (N_7490,N_6027,N_6767);
nor U7491 (N_7491,N_6004,N_6394);
and U7492 (N_7492,N_6387,N_6958);
and U7493 (N_7493,N_6550,N_6511);
nand U7494 (N_7494,N_6400,N_6296);
nor U7495 (N_7495,N_6797,N_6010);
nand U7496 (N_7496,N_6199,N_6917);
nor U7497 (N_7497,N_6099,N_6344);
nor U7498 (N_7498,N_6438,N_6228);
nor U7499 (N_7499,N_6950,N_6014);
and U7500 (N_7500,N_6149,N_6392);
and U7501 (N_7501,N_6809,N_6053);
nor U7502 (N_7502,N_6374,N_6572);
nand U7503 (N_7503,N_6870,N_6977);
nor U7504 (N_7504,N_6365,N_6465);
and U7505 (N_7505,N_6175,N_6683);
nor U7506 (N_7506,N_6196,N_6022);
nor U7507 (N_7507,N_6163,N_6012);
and U7508 (N_7508,N_6522,N_6832);
xor U7509 (N_7509,N_6523,N_6770);
or U7510 (N_7510,N_6291,N_6502);
and U7511 (N_7511,N_6226,N_6440);
or U7512 (N_7512,N_6827,N_6100);
and U7513 (N_7513,N_6383,N_6853);
nand U7514 (N_7514,N_6905,N_6620);
and U7515 (N_7515,N_6092,N_6858);
or U7516 (N_7516,N_6541,N_6958);
nand U7517 (N_7517,N_6086,N_6139);
or U7518 (N_7518,N_6769,N_6993);
nand U7519 (N_7519,N_6141,N_6910);
and U7520 (N_7520,N_6821,N_6957);
nor U7521 (N_7521,N_6345,N_6560);
nor U7522 (N_7522,N_6391,N_6746);
or U7523 (N_7523,N_6212,N_6548);
or U7524 (N_7524,N_6476,N_6470);
nand U7525 (N_7525,N_6328,N_6856);
nor U7526 (N_7526,N_6980,N_6403);
and U7527 (N_7527,N_6687,N_6625);
nand U7528 (N_7528,N_6927,N_6884);
nand U7529 (N_7529,N_6358,N_6454);
and U7530 (N_7530,N_6089,N_6441);
or U7531 (N_7531,N_6531,N_6052);
or U7532 (N_7532,N_6506,N_6053);
nor U7533 (N_7533,N_6094,N_6596);
nor U7534 (N_7534,N_6466,N_6566);
and U7535 (N_7535,N_6776,N_6597);
nor U7536 (N_7536,N_6203,N_6038);
nand U7537 (N_7537,N_6547,N_6694);
nand U7538 (N_7538,N_6739,N_6335);
or U7539 (N_7539,N_6808,N_6902);
or U7540 (N_7540,N_6524,N_6269);
and U7541 (N_7541,N_6466,N_6084);
nor U7542 (N_7542,N_6409,N_6930);
or U7543 (N_7543,N_6814,N_6051);
or U7544 (N_7544,N_6324,N_6015);
or U7545 (N_7545,N_6045,N_6563);
nand U7546 (N_7546,N_6939,N_6301);
or U7547 (N_7547,N_6626,N_6980);
nand U7548 (N_7548,N_6903,N_6210);
and U7549 (N_7549,N_6734,N_6464);
nand U7550 (N_7550,N_6358,N_6555);
and U7551 (N_7551,N_6922,N_6076);
nand U7552 (N_7552,N_6008,N_6287);
nand U7553 (N_7553,N_6653,N_6330);
and U7554 (N_7554,N_6754,N_6138);
nand U7555 (N_7555,N_6296,N_6602);
and U7556 (N_7556,N_6619,N_6472);
nor U7557 (N_7557,N_6739,N_6877);
and U7558 (N_7558,N_6789,N_6499);
nand U7559 (N_7559,N_6008,N_6423);
and U7560 (N_7560,N_6739,N_6595);
nor U7561 (N_7561,N_6914,N_6899);
and U7562 (N_7562,N_6256,N_6415);
and U7563 (N_7563,N_6906,N_6091);
nor U7564 (N_7564,N_6604,N_6236);
nand U7565 (N_7565,N_6580,N_6339);
nand U7566 (N_7566,N_6918,N_6735);
nor U7567 (N_7567,N_6158,N_6647);
or U7568 (N_7568,N_6907,N_6962);
and U7569 (N_7569,N_6297,N_6112);
nor U7570 (N_7570,N_6420,N_6286);
nand U7571 (N_7571,N_6333,N_6403);
nand U7572 (N_7572,N_6770,N_6678);
nand U7573 (N_7573,N_6772,N_6925);
or U7574 (N_7574,N_6143,N_6725);
and U7575 (N_7575,N_6053,N_6378);
and U7576 (N_7576,N_6380,N_6579);
or U7577 (N_7577,N_6043,N_6121);
or U7578 (N_7578,N_6441,N_6975);
or U7579 (N_7579,N_6350,N_6043);
and U7580 (N_7580,N_6939,N_6331);
nand U7581 (N_7581,N_6946,N_6297);
or U7582 (N_7582,N_6188,N_6303);
nand U7583 (N_7583,N_6789,N_6542);
nor U7584 (N_7584,N_6519,N_6572);
nor U7585 (N_7585,N_6053,N_6287);
or U7586 (N_7586,N_6445,N_6688);
nor U7587 (N_7587,N_6503,N_6752);
nand U7588 (N_7588,N_6817,N_6780);
or U7589 (N_7589,N_6467,N_6864);
nand U7590 (N_7590,N_6063,N_6973);
and U7591 (N_7591,N_6991,N_6920);
and U7592 (N_7592,N_6500,N_6072);
nor U7593 (N_7593,N_6738,N_6779);
and U7594 (N_7594,N_6575,N_6792);
or U7595 (N_7595,N_6740,N_6729);
nor U7596 (N_7596,N_6972,N_6561);
nand U7597 (N_7597,N_6525,N_6456);
and U7598 (N_7598,N_6751,N_6965);
or U7599 (N_7599,N_6586,N_6962);
or U7600 (N_7600,N_6714,N_6527);
nand U7601 (N_7601,N_6088,N_6251);
and U7602 (N_7602,N_6131,N_6720);
and U7603 (N_7603,N_6676,N_6202);
and U7604 (N_7604,N_6089,N_6407);
nor U7605 (N_7605,N_6490,N_6511);
nand U7606 (N_7606,N_6172,N_6911);
nor U7607 (N_7607,N_6257,N_6172);
and U7608 (N_7608,N_6307,N_6221);
and U7609 (N_7609,N_6934,N_6318);
and U7610 (N_7610,N_6721,N_6427);
nand U7611 (N_7611,N_6959,N_6102);
and U7612 (N_7612,N_6497,N_6979);
nor U7613 (N_7613,N_6959,N_6875);
nor U7614 (N_7614,N_6840,N_6878);
nand U7615 (N_7615,N_6323,N_6403);
nor U7616 (N_7616,N_6198,N_6982);
nand U7617 (N_7617,N_6947,N_6635);
nand U7618 (N_7618,N_6870,N_6016);
or U7619 (N_7619,N_6079,N_6628);
or U7620 (N_7620,N_6642,N_6097);
nand U7621 (N_7621,N_6869,N_6190);
or U7622 (N_7622,N_6098,N_6628);
or U7623 (N_7623,N_6159,N_6228);
and U7624 (N_7624,N_6803,N_6344);
nor U7625 (N_7625,N_6936,N_6916);
nor U7626 (N_7626,N_6751,N_6976);
or U7627 (N_7627,N_6399,N_6425);
nand U7628 (N_7628,N_6532,N_6748);
and U7629 (N_7629,N_6417,N_6808);
and U7630 (N_7630,N_6004,N_6863);
or U7631 (N_7631,N_6771,N_6462);
nor U7632 (N_7632,N_6411,N_6951);
nor U7633 (N_7633,N_6033,N_6009);
nor U7634 (N_7634,N_6413,N_6618);
nor U7635 (N_7635,N_6974,N_6307);
nor U7636 (N_7636,N_6237,N_6177);
nand U7637 (N_7637,N_6350,N_6659);
nor U7638 (N_7638,N_6401,N_6797);
or U7639 (N_7639,N_6393,N_6362);
nand U7640 (N_7640,N_6279,N_6079);
nand U7641 (N_7641,N_6513,N_6076);
and U7642 (N_7642,N_6463,N_6501);
or U7643 (N_7643,N_6593,N_6534);
nand U7644 (N_7644,N_6126,N_6767);
nand U7645 (N_7645,N_6166,N_6303);
and U7646 (N_7646,N_6900,N_6639);
nor U7647 (N_7647,N_6150,N_6823);
and U7648 (N_7648,N_6787,N_6159);
nand U7649 (N_7649,N_6849,N_6373);
nand U7650 (N_7650,N_6536,N_6182);
nor U7651 (N_7651,N_6103,N_6660);
or U7652 (N_7652,N_6657,N_6578);
and U7653 (N_7653,N_6189,N_6414);
nor U7654 (N_7654,N_6767,N_6013);
and U7655 (N_7655,N_6822,N_6731);
nor U7656 (N_7656,N_6790,N_6120);
or U7657 (N_7657,N_6921,N_6634);
or U7658 (N_7658,N_6836,N_6356);
or U7659 (N_7659,N_6862,N_6118);
or U7660 (N_7660,N_6195,N_6971);
nor U7661 (N_7661,N_6580,N_6351);
nand U7662 (N_7662,N_6925,N_6832);
or U7663 (N_7663,N_6135,N_6051);
and U7664 (N_7664,N_6554,N_6508);
nand U7665 (N_7665,N_6734,N_6967);
or U7666 (N_7666,N_6826,N_6469);
nand U7667 (N_7667,N_6576,N_6477);
or U7668 (N_7668,N_6594,N_6253);
and U7669 (N_7669,N_6703,N_6855);
nor U7670 (N_7670,N_6405,N_6793);
nand U7671 (N_7671,N_6142,N_6799);
or U7672 (N_7672,N_6030,N_6934);
xnor U7673 (N_7673,N_6332,N_6052);
or U7674 (N_7674,N_6179,N_6872);
nor U7675 (N_7675,N_6494,N_6336);
and U7676 (N_7676,N_6834,N_6943);
nand U7677 (N_7677,N_6968,N_6313);
nand U7678 (N_7678,N_6122,N_6025);
or U7679 (N_7679,N_6834,N_6913);
and U7680 (N_7680,N_6311,N_6209);
or U7681 (N_7681,N_6868,N_6370);
nor U7682 (N_7682,N_6611,N_6530);
nand U7683 (N_7683,N_6574,N_6275);
or U7684 (N_7684,N_6531,N_6775);
nor U7685 (N_7685,N_6223,N_6728);
nand U7686 (N_7686,N_6135,N_6072);
nand U7687 (N_7687,N_6059,N_6101);
xor U7688 (N_7688,N_6123,N_6472);
nor U7689 (N_7689,N_6807,N_6127);
nor U7690 (N_7690,N_6313,N_6076);
or U7691 (N_7691,N_6481,N_6986);
or U7692 (N_7692,N_6726,N_6658);
nor U7693 (N_7693,N_6167,N_6884);
nand U7694 (N_7694,N_6235,N_6142);
and U7695 (N_7695,N_6454,N_6501);
or U7696 (N_7696,N_6247,N_6567);
and U7697 (N_7697,N_6389,N_6021);
or U7698 (N_7698,N_6094,N_6116);
or U7699 (N_7699,N_6352,N_6747);
nor U7700 (N_7700,N_6047,N_6128);
nor U7701 (N_7701,N_6951,N_6597);
or U7702 (N_7702,N_6398,N_6646);
or U7703 (N_7703,N_6706,N_6363);
nand U7704 (N_7704,N_6595,N_6937);
nand U7705 (N_7705,N_6956,N_6366);
nand U7706 (N_7706,N_6141,N_6784);
or U7707 (N_7707,N_6582,N_6669);
xnor U7708 (N_7708,N_6905,N_6096);
xnor U7709 (N_7709,N_6247,N_6635);
nand U7710 (N_7710,N_6089,N_6644);
and U7711 (N_7711,N_6824,N_6603);
nand U7712 (N_7712,N_6959,N_6026);
nand U7713 (N_7713,N_6264,N_6367);
or U7714 (N_7714,N_6272,N_6504);
nand U7715 (N_7715,N_6725,N_6711);
or U7716 (N_7716,N_6075,N_6996);
or U7717 (N_7717,N_6546,N_6585);
nand U7718 (N_7718,N_6334,N_6589);
nand U7719 (N_7719,N_6097,N_6930);
or U7720 (N_7720,N_6049,N_6546);
and U7721 (N_7721,N_6289,N_6898);
nor U7722 (N_7722,N_6666,N_6250);
nand U7723 (N_7723,N_6235,N_6574);
or U7724 (N_7724,N_6313,N_6770);
nand U7725 (N_7725,N_6967,N_6837);
or U7726 (N_7726,N_6365,N_6356);
or U7727 (N_7727,N_6135,N_6832);
or U7728 (N_7728,N_6925,N_6971);
or U7729 (N_7729,N_6104,N_6361);
and U7730 (N_7730,N_6832,N_6151);
or U7731 (N_7731,N_6716,N_6120);
and U7732 (N_7732,N_6497,N_6863);
and U7733 (N_7733,N_6157,N_6853);
xnor U7734 (N_7734,N_6146,N_6941);
nor U7735 (N_7735,N_6175,N_6639);
xnor U7736 (N_7736,N_6475,N_6450);
nand U7737 (N_7737,N_6460,N_6809);
or U7738 (N_7738,N_6971,N_6969);
nand U7739 (N_7739,N_6219,N_6954);
nor U7740 (N_7740,N_6790,N_6568);
and U7741 (N_7741,N_6075,N_6793);
and U7742 (N_7742,N_6492,N_6244);
nor U7743 (N_7743,N_6865,N_6530);
and U7744 (N_7744,N_6375,N_6698);
or U7745 (N_7745,N_6188,N_6418);
or U7746 (N_7746,N_6137,N_6974);
nor U7747 (N_7747,N_6989,N_6493);
or U7748 (N_7748,N_6513,N_6162);
and U7749 (N_7749,N_6839,N_6691);
nor U7750 (N_7750,N_6379,N_6638);
nand U7751 (N_7751,N_6368,N_6023);
nand U7752 (N_7752,N_6140,N_6144);
nand U7753 (N_7753,N_6882,N_6801);
nor U7754 (N_7754,N_6417,N_6270);
and U7755 (N_7755,N_6978,N_6360);
or U7756 (N_7756,N_6737,N_6358);
or U7757 (N_7757,N_6041,N_6723);
nand U7758 (N_7758,N_6081,N_6484);
nand U7759 (N_7759,N_6836,N_6724);
nor U7760 (N_7760,N_6785,N_6589);
or U7761 (N_7761,N_6540,N_6506);
or U7762 (N_7762,N_6973,N_6253);
and U7763 (N_7763,N_6509,N_6867);
nand U7764 (N_7764,N_6408,N_6802);
and U7765 (N_7765,N_6763,N_6102);
and U7766 (N_7766,N_6308,N_6226);
nand U7767 (N_7767,N_6272,N_6614);
nand U7768 (N_7768,N_6432,N_6621);
or U7769 (N_7769,N_6371,N_6058);
nor U7770 (N_7770,N_6356,N_6735);
nand U7771 (N_7771,N_6379,N_6855);
or U7772 (N_7772,N_6604,N_6147);
nor U7773 (N_7773,N_6911,N_6746);
nand U7774 (N_7774,N_6434,N_6152);
nor U7775 (N_7775,N_6007,N_6583);
nor U7776 (N_7776,N_6198,N_6101);
or U7777 (N_7777,N_6369,N_6942);
and U7778 (N_7778,N_6350,N_6404);
nor U7779 (N_7779,N_6754,N_6904);
or U7780 (N_7780,N_6554,N_6887);
nand U7781 (N_7781,N_6161,N_6767);
or U7782 (N_7782,N_6693,N_6321);
or U7783 (N_7783,N_6181,N_6062);
and U7784 (N_7784,N_6485,N_6328);
or U7785 (N_7785,N_6785,N_6725);
and U7786 (N_7786,N_6623,N_6384);
or U7787 (N_7787,N_6537,N_6803);
nand U7788 (N_7788,N_6228,N_6333);
or U7789 (N_7789,N_6777,N_6814);
nand U7790 (N_7790,N_6374,N_6544);
nand U7791 (N_7791,N_6298,N_6782);
nand U7792 (N_7792,N_6448,N_6225);
nand U7793 (N_7793,N_6741,N_6626);
and U7794 (N_7794,N_6509,N_6620);
nand U7795 (N_7795,N_6195,N_6669);
nor U7796 (N_7796,N_6630,N_6794);
nand U7797 (N_7797,N_6737,N_6760);
nor U7798 (N_7798,N_6395,N_6928);
nand U7799 (N_7799,N_6580,N_6000);
and U7800 (N_7800,N_6316,N_6270);
xnor U7801 (N_7801,N_6636,N_6444);
or U7802 (N_7802,N_6704,N_6836);
nand U7803 (N_7803,N_6353,N_6098);
nor U7804 (N_7804,N_6273,N_6609);
or U7805 (N_7805,N_6744,N_6889);
and U7806 (N_7806,N_6925,N_6324);
or U7807 (N_7807,N_6189,N_6861);
and U7808 (N_7808,N_6208,N_6711);
nor U7809 (N_7809,N_6686,N_6317);
nor U7810 (N_7810,N_6568,N_6209);
or U7811 (N_7811,N_6671,N_6747);
nand U7812 (N_7812,N_6103,N_6091);
or U7813 (N_7813,N_6186,N_6220);
nand U7814 (N_7814,N_6107,N_6181);
nand U7815 (N_7815,N_6412,N_6191);
nor U7816 (N_7816,N_6075,N_6127);
nor U7817 (N_7817,N_6421,N_6907);
or U7818 (N_7818,N_6001,N_6617);
and U7819 (N_7819,N_6033,N_6896);
and U7820 (N_7820,N_6638,N_6630);
nand U7821 (N_7821,N_6472,N_6986);
nor U7822 (N_7822,N_6778,N_6310);
nor U7823 (N_7823,N_6620,N_6434);
nand U7824 (N_7824,N_6603,N_6716);
or U7825 (N_7825,N_6770,N_6355);
or U7826 (N_7826,N_6225,N_6219);
nor U7827 (N_7827,N_6396,N_6620);
or U7828 (N_7828,N_6105,N_6206);
and U7829 (N_7829,N_6500,N_6419);
nor U7830 (N_7830,N_6634,N_6557);
and U7831 (N_7831,N_6645,N_6745);
nand U7832 (N_7832,N_6110,N_6047);
nor U7833 (N_7833,N_6882,N_6311);
or U7834 (N_7834,N_6003,N_6412);
nor U7835 (N_7835,N_6548,N_6914);
nor U7836 (N_7836,N_6825,N_6406);
nor U7837 (N_7837,N_6269,N_6167);
nand U7838 (N_7838,N_6645,N_6820);
nor U7839 (N_7839,N_6573,N_6472);
or U7840 (N_7840,N_6582,N_6758);
nor U7841 (N_7841,N_6860,N_6736);
or U7842 (N_7842,N_6187,N_6779);
or U7843 (N_7843,N_6962,N_6822);
and U7844 (N_7844,N_6673,N_6205);
or U7845 (N_7845,N_6469,N_6391);
nor U7846 (N_7846,N_6221,N_6551);
nor U7847 (N_7847,N_6997,N_6413);
nor U7848 (N_7848,N_6630,N_6319);
nor U7849 (N_7849,N_6358,N_6022);
or U7850 (N_7850,N_6921,N_6737);
nor U7851 (N_7851,N_6059,N_6441);
nor U7852 (N_7852,N_6842,N_6518);
and U7853 (N_7853,N_6743,N_6434);
nand U7854 (N_7854,N_6548,N_6441);
nor U7855 (N_7855,N_6178,N_6190);
and U7856 (N_7856,N_6130,N_6162);
or U7857 (N_7857,N_6067,N_6154);
and U7858 (N_7858,N_6845,N_6935);
nor U7859 (N_7859,N_6344,N_6658);
and U7860 (N_7860,N_6845,N_6444);
nor U7861 (N_7861,N_6927,N_6782);
nor U7862 (N_7862,N_6600,N_6543);
xnor U7863 (N_7863,N_6705,N_6291);
nor U7864 (N_7864,N_6632,N_6127);
and U7865 (N_7865,N_6797,N_6596);
nor U7866 (N_7866,N_6167,N_6179);
or U7867 (N_7867,N_6978,N_6248);
xnor U7868 (N_7868,N_6427,N_6238);
or U7869 (N_7869,N_6877,N_6299);
nand U7870 (N_7870,N_6390,N_6825);
or U7871 (N_7871,N_6291,N_6161);
and U7872 (N_7872,N_6157,N_6355);
nand U7873 (N_7873,N_6664,N_6394);
or U7874 (N_7874,N_6896,N_6426);
and U7875 (N_7875,N_6284,N_6341);
and U7876 (N_7876,N_6055,N_6322);
and U7877 (N_7877,N_6707,N_6095);
nand U7878 (N_7878,N_6558,N_6787);
nor U7879 (N_7879,N_6700,N_6595);
nand U7880 (N_7880,N_6629,N_6376);
or U7881 (N_7881,N_6420,N_6049);
nor U7882 (N_7882,N_6998,N_6779);
nor U7883 (N_7883,N_6756,N_6238);
nor U7884 (N_7884,N_6056,N_6945);
nor U7885 (N_7885,N_6051,N_6441);
or U7886 (N_7886,N_6896,N_6936);
or U7887 (N_7887,N_6114,N_6244);
nand U7888 (N_7888,N_6694,N_6285);
nand U7889 (N_7889,N_6847,N_6687);
and U7890 (N_7890,N_6270,N_6047);
or U7891 (N_7891,N_6342,N_6540);
nor U7892 (N_7892,N_6068,N_6096);
or U7893 (N_7893,N_6841,N_6204);
nand U7894 (N_7894,N_6264,N_6120);
nand U7895 (N_7895,N_6176,N_6475);
and U7896 (N_7896,N_6664,N_6678);
nand U7897 (N_7897,N_6354,N_6439);
nor U7898 (N_7898,N_6121,N_6608);
or U7899 (N_7899,N_6849,N_6441);
or U7900 (N_7900,N_6105,N_6185);
or U7901 (N_7901,N_6078,N_6543);
nand U7902 (N_7902,N_6803,N_6452);
or U7903 (N_7903,N_6631,N_6135);
or U7904 (N_7904,N_6138,N_6867);
and U7905 (N_7905,N_6970,N_6546);
xor U7906 (N_7906,N_6182,N_6872);
nand U7907 (N_7907,N_6542,N_6537);
nor U7908 (N_7908,N_6824,N_6693);
nand U7909 (N_7909,N_6578,N_6805);
nand U7910 (N_7910,N_6690,N_6300);
nor U7911 (N_7911,N_6667,N_6241);
nor U7912 (N_7912,N_6062,N_6617);
and U7913 (N_7913,N_6659,N_6710);
nor U7914 (N_7914,N_6695,N_6957);
xnor U7915 (N_7915,N_6742,N_6504);
and U7916 (N_7916,N_6581,N_6785);
and U7917 (N_7917,N_6515,N_6630);
and U7918 (N_7918,N_6906,N_6314);
nand U7919 (N_7919,N_6816,N_6387);
or U7920 (N_7920,N_6402,N_6921);
and U7921 (N_7921,N_6720,N_6493);
and U7922 (N_7922,N_6414,N_6710);
or U7923 (N_7923,N_6536,N_6124);
or U7924 (N_7924,N_6382,N_6497);
and U7925 (N_7925,N_6668,N_6989);
or U7926 (N_7926,N_6087,N_6816);
or U7927 (N_7927,N_6229,N_6188);
nand U7928 (N_7928,N_6984,N_6294);
and U7929 (N_7929,N_6749,N_6790);
and U7930 (N_7930,N_6292,N_6832);
and U7931 (N_7931,N_6098,N_6026);
nor U7932 (N_7932,N_6313,N_6760);
and U7933 (N_7933,N_6506,N_6672);
nand U7934 (N_7934,N_6082,N_6879);
nand U7935 (N_7935,N_6481,N_6606);
nand U7936 (N_7936,N_6118,N_6718);
and U7937 (N_7937,N_6245,N_6366);
nor U7938 (N_7938,N_6638,N_6248);
and U7939 (N_7939,N_6699,N_6991);
xor U7940 (N_7940,N_6004,N_6677);
and U7941 (N_7941,N_6000,N_6617);
nand U7942 (N_7942,N_6450,N_6254);
nor U7943 (N_7943,N_6020,N_6262);
nand U7944 (N_7944,N_6175,N_6291);
and U7945 (N_7945,N_6944,N_6616);
and U7946 (N_7946,N_6074,N_6553);
nand U7947 (N_7947,N_6076,N_6060);
nand U7948 (N_7948,N_6873,N_6380);
or U7949 (N_7949,N_6108,N_6529);
nand U7950 (N_7950,N_6514,N_6954);
or U7951 (N_7951,N_6458,N_6248);
and U7952 (N_7952,N_6311,N_6875);
or U7953 (N_7953,N_6080,N_6791);
or U7954 (N_7954,N_6018,N_6672);
nand U7955 (N_7955,N_6565,N_6890);
nand U7956 (N_7956,N_6576,N_6611);
nand U7957 (N_7957,N_6165,N_6164);
and U7958 (N_7958,N_6595,N_6092);
nand U7959 (N_7959,N_6963,N_6759);
and U7960 (N_7960,N_6661,N_6966);
and U7961 (N_7961,N_6282,N_6263);
nand U7962 (N_7962,N_6720,N_6346);
nand U7963 (N_7963,N_6091,N_6357);
and U7964 (N_7964,N_6676,N_6332);
nand U7965 (N_7965,N_6158,N_6509);
or U7966 (N_7966,N_6091,N_6488);
and U7967 (N_7967,N_6569,N_6510);
and U7968 (N_7968,N_6412,N_6111);
nand U7969 (N_7969,N_6817,N_6853);
xor U7970 (N_7970,N_6584,N_6887);
and U7971 (N_7971,N_6496,N_6319);
and U7972 (N_7972,N_6598,N_6279);
nand U7973 (N_7973,N_6437,N_6564);
xor U7974 (N_7974,N_6157,N_6303);
nand U7975 (N_7975,N_6308,N_6504);
and U7976 (N_7976,N_6135,N_6673);
or U7977 (N_7977,N_6183,N_6950);
or U7978 (N_7978,N_6306,N_6290);
nor U7979 (N_7979,N_6067,N_6694);
or U7980 (N_7980,N_6108,N_6556);
nand U7981 (N_7981,N_6815,N_6099);
or U7982 (N_7982,N_6590,N_6231);
and U7983 (N_7983,N_6804,N_6581);
nor U7984 (N_7984,N_6925,N_6300);
nand U7985 (N_7985,N_6025,N_6399);
nand U7986 (N_7986,N_6636,N_6532);
or U7987 (N_7987,N_6537,N_6717);
or U7988 (N_7988,N_6306,N_6389);
nand U7989 (N_7989,N_6984,N_6334);
nand U7990 (N_7990,N_6613,N_6499);
or U7991 (N_7991,N_6685,N_6633);
nor U7992 (N_7992,N_6844,N_6346);
nand U7993 (N_7993,N_6099,N_6103);
and U7994 (N_7994,N_6615,N_6298);
and U7995 (N_7995,N_6469,N_6066);
or U7996 (N_7996,N_6359,N_6687);
nor U7997 (N_7997,N_6553,N_6126);
nand U7998 (N_7998,N_6206,N_6016);
nor U7999 (N_7999,N_6092,N_6766);
or U8000 (N_8000,N_7334,N_7019);
nor U8001 (N_8001,N_7615,N_7795);
or U8002 (N_8002,N_7843,N_7147);
or U8003 (N_8003,N_7776,N_7181);
nor U8004 (N_8004,N_7996,N_7386);
or U8005 (N_8005,N_7909,N_7339);
nor U8006 (N_8006,N_7313,N_7180);
nor U8007 (N_8007,N_7579,N_7040);
and U8008 (N_8008,N_7924,N_7985);
nand U8009 (N_8009,N_7130,N_7533);
nand U8010 (N_8010,N_7497,N_7511);
nand U8011 (N_8011,N_7954,N_7193);
nand U8012 (N_8012,N_7126,N_7506);
nor U8013 (N_8013,N_7343,N_7659);
nand U8014 (N_8014,N_7914,N_7588);
and U8015 (N_8015,N_7944,N_7308);
nor U8016 (N_8016,N_7173,N_7875);
or U8017 (N_8017,N_7791,N_7075);
or U8018 (N_8018,N_7369,N_7200);
nand U8019 (N_8019,N_7488,N_7738);
nand U8020 (N_8020,N_7543,N_7089);
nor U8021 (N_8021,N_7810,N_7933);
or U8022 (N_8022,N_7640,N_7046);
or U8023 (N_8023,N_7793,N_7146);
or U8024 (N_8024,N_7805,N_7893);
or U8025 (N_8025,N_7912,N_7621);
nor U8026 (N_8026,N_7743,N_7017);
nand U8027 (N_8027,N_7063,N_7184);
nor U8028 (N_8028,N_7225,N_7629);
and U8029 (N_8029,N_7548,N_7709);
nand U8030 (N_8030,N_7101,N_7554);
nand U8031 (N_8031,N_7323,N_7735);
or U8032 (N_8032,N_7142,N_7301);
nand U8033 (N_8033,N_7674,N_7680);
or U8034 (N_8034,N_7752,N_7387);
nand U8035 (N_8035,N_7410,N_7405);
and U8036 (N_8036,N_7941,N_7218);
nand U8037 (N_8037,N_7797,N_7982);
nor U8038 (N_8038,N_7698,N_7578);
and U8039 (N_8039,N_7054,N_7731);
nand U8040 (N_8040,N_7898,N_7445);
or U8041 (N_8041,N_7549,N_7043);
nor U8042 (N_8042,N_7788,N_7639);
and U8043 (N_8043,N_7446,N_7178);
nand U8044 (N_8044,N_7468,N_7160);
nand U8045 (N_8045,N_7902,N_7508);
nor U8046 (N_8046,N_7792,N_7449);
and U8047 (N_8047,N_7913,N_7097);
nand U8048 (N_8048,N_7668,N_7963);
nor U8049 (N_8049,N_7813,N_7612);
nand U8050 (N_8050,N_7604,N_7018);
and U8051 (N_8051,N_7310,N_7037);
nand U8052 (N_8052,N_7189,N_7027);
and U8053 (N_8053,N_7627,N_7357);
or U8054 (N_8054,N_7920,N_7164);
nor U8055 (N_8055,N_7161,N_7916);
nor U8056 (N_8056,N_7790,N_7266);
nor U8057 (N_8057,N_7513,N_7887);
nand U8058 (N_8058,N_7083,N_7910);
nand U8059 (N_8059,N_7885,N_7118);
or U8060 (N_8060,N_7960,N_7441);
nand U8061 (N_8061,N_7849,N_7727);
and U8062 (N_8062,N_7952,N_7165);
nand U8063 (N_8063,N_7501,N_7945);
and U8064 (N_8064,N_7248,N_7412);
nand U8065 (N_8065,N_7626,N_7447);
or U8066 (N_8066,N_7229,N_7451);
nand U8067 (N_8067,N_7450,N_7486);
nor U8068 (N_8068,N_7082,N_7419);
nor U8069 (N_8069,N_7479,N_7679);
nor U8070 (N_8070,N_7438,N_7264);
nand U8071 (N_8071,N_7532,N_7110);
or U8072 (N_8072,N_7072,N_7570);
nand U8073 (N_8073,N_7256,N_7871);
or U8074 (N_8074,N_7757,N_7827);
and U8075 (N_8075,N_7551,N_7705);
nor U8076 (N_8076,N_7775,N_7465);
nand U8077 (N_8077,N_7879,N_7759);
and U8078 (N_8078,N_7732,N_7074);
nor U8079 (N_8079,N_7806,N_7584);
nor U8080 (N_8080,N_7926,N_7762);
and U8081 (N_8081,N_7362,N_7836);
nor U8082 (N_8082,N_7948,N_7300);
nor U8083 (N_8083,N_7550,N_7587);
nand U8084 (N_8084,N_7758,N_7416);
nor U8085 (N_8085,N_7677,N_7864);
nand U8086 (N_8086,N_7581,N_7121);
nor U8087 (N_8087,N_7992,N_7107);
and U8088 (N_8088,N_7900,N_7411);
or U8089 (N_8089,N_7657,N_7056);
or U8090 (N_8090,N_7474,N_7574);
nand U8091 (N_8091,N_7383,N_7342);
or U8092 (N_8092,N_7254,N_7232);
or U8093 (N_8093,N_7038,N_7318);
or U8094 (N_8094,N_7528,N_7456);
or U8095 (N_8095,N_7865,N_7039);
or U8096 (N_8096,N_7919,N_7669);
nor U8097 (N_8097,N_7482,N_7653);
and U8098 (N_8098,N_7031,N_7713);
or U8099 (N_8099,N_7966,N_7319);
nor U8100 (N_8100,N_7157,N_7923);
nor U8101 (N_8101,N_7141,N_7003);
nand U8102 (N_8102,N_7702,N_7304);
nor U8103 (N_8103,N_7053,N_7891);
or U8104 (N_8104,N_7077,N_7377);
or U8105 (N_8105,N_7568,N_7324);
or U8106 (N_8106,N_7086,N_7594);
nor U8107 (N_8107,N_7841,N_7991);
nor U8108 (N_8108,N_7580,N_7403);
nor U8109 (N_8109,N_7703,N_7523);
nand U8110 (N_8110,N_7971,N_7290);
nor U8111 (N_8111,N_7974,N_7719);
or U8112 (N_8112,N_7191,N_7279);
xor U8113 (N_8113,N_7768,N_7375);
or U8114 (N_8114,N_7517,N_7443);
or U8115 (N_8115,N_7564,N_7278);
nand U8116 (N_8116,N_7648,N_7995);
nor U8117 (N_8117,N_7736,N_7502);
and U8118 (N_8118,N_7878,N_7823);
and U8119 (N_8119,N_7744,N_7483);
or U8120 (N_8120,N_7485,N_7880);
nor U8121 (N_8121,N_7590,N_7346);
or U8122 (N_8122,N_7395,N_7745);
and U8123 (N_8123,N_7062,N_7041);
xnor U8124 (N_8124,N_7964,N_7182);
nor U8125 (N_8125,N_7714,N_7239);
nand U8126 (N_8126,N_7658,N_7022);
or U8127 (N_8127,N_7382,N_7049);
nor U8128 (N_8128,N_7922,N_7609);
nor U8129 (N_8129,N_7496,N_7473);
or U8130 (N_8130,N_7662,N_7903);
nor U8131 (N_8131,N_7822,N_7350);
nand U8132 (N_8132,N_7614,N_7076);
nor U8133 (N_8133,N_7135,N_7915);
and U8134 (N_8134,N_7837,N_7093);
nand U8135 (N_8135,N_7381,N_7959);
or U8136 (N_8136,N_7807,N_7600);
or U8137 (N_8137,N_7844,N_7859);
or U8138 (N_8138,N_7299,N_7080);
and U8139 (N_8139,N_7556,N_7060);
and U8140 (N_8140,N_7721,N_7437);
nand U8141 (N_8141,N_7651,N_7355);
and U8142 (N_8142,N_7666,N_7454);
nor U8143 (N_8143,N_7618,N_7616);
nor U8144 (N_8144,N_7487,N_7812);
nand U8145 (N_8145,N_7457,N_7009);
nand U8146 (N_8146,N_7881,N_7630);
and U8147 (N_8147,N_7316,N_7407);
and U8148 (N_8148,N_7582,N_7071);
nand U8149 (N_8149,N_7785,N_7575);
or U8150 (N_8150,N_7185,N_7802);
and U8151 (N_8151,N_7004,N_7128);
or U8152 (N_8152,N_7633,N_7809);
and U8153 (N_8153,N_7529,N_7842);
nor U8154 (N_8154,N_7695,N_7675);
and U8155 (N_8155,N_7955,N_7979);
or U8156 (N_8156,N_7320,N_7632);
or U8157 (N_8157,N_7749,N_7149);
and U8158 (N_8158,N_7460,N_7665);
or U8159 (N_8159,N_7655,N_7469);
and U8160 (N_8160,N_7002,N_7845);
nor U8161 (N_8161,N_7722,N_7011);
and U8162 (N_8162,N_7379,N_7390);
nor U8163 (N_8163,N_7282,N_7710);
nor U8164 (N_8164,N_7862,N_7398);
or U8165 (N_8165,N_7918,N_7092);
nand U8166 (N_8166,N_7811,N_7650);
and U8167 (N_8167,N_7977,N_7030);
nand U8168 (N_8168,N_7817,N_7592);
nor U8169 (N_8169,N_7777,N_7925);
nor U8170 (N_8170,N_7249,N_7127);
nor U8171 (N_8171,N_7751,N_7409);
and U8172 (N_8172,N_7839,N_7471);
and U8173 (N_8173,N_7183,N_7882);
and U8174 (N_8174,N_7928,N_7832);
nand U8175 (N_8175,N_7322,N_7644);
and U8176 (N_8176,N_7593,N_7760);
nand U8177 (N_8177,N_7997,N_7470);
nand U8178 (N_8178,N_7641,N_7628);
or U8179 (N_8179,N_7771,N_7515);
nand U8180 (N_8180,N_7453,N_7289);
and U8181 (N_8181,N_7492,N_7159);
or U8182 (N_8182,N_7253,N_7888);
or U8183 (N_8183,N_7269,N_7190);
or U8184 (N_8184,N_7421,N_7246);
or U8185 (N_8185,N_7904,N_7341);
or U8186 (N_8186,N_7167,N_7534);
nor U8187 (N_8187,N_7032,N_7001);
and U8188 (N_8188,N_7286,N_7380);
nand U8189 (N_8189,N_7188,N_7602);
nand U8190 (N_8190,N_7868,N_7064);
nand U8191 (N_8191,N_7539,N_7569);
nand U8192 (N_8192,N_7678,N_7148);
and U8193 (N_8193,N_7957,N_7434);
nor U8194 (N_8194,N_7877,N_7026);
nand U8195 (N_8195,N_7786,N_7134);
or U8196 (N_8196,N_7230,N_7544);
nand U8197 (N_8197,N_7078,N_7417);
nor U8198 (N_8198,N_7363,N_7883);
and U8199 (N_8199,N_7047,N_7195);
xnor U8200 (N_8200,N_7537,N_7664);
nand U8201 (N_8201,N_7563,N_7023);
nand U8202 (N_8202,N_7660,N_7541);
nor U8203 (N_8203,N_7654,N_7228);
and U8204 (N_8204,N_7284,N_7696);
nand U8205 (N_8205,N_7969,N_7586);
nand U8206 (N_8206,N_7129,N_7965);
or U8207 (N_8207,N_7661,N_7467);
nand U8208 (N_8208,N_7427,N_7431);
and U8209 (N_8209,N_7998,N_7667);
nand U8210 (N_8210,N_7152,N_7156);
nand U8211 (N_8211,N_7572,N_7858);
nand U8212 (N_8212,N_7252,N_7692);
nand U8213 (N_8213,N_7436,N_7521);
nor U8214 (N_8214,N_7756,N_7087);
nand U8215 (N_8215,N_7336,N_7365);
and U8216 (N_8216,N_7361,N_7988);
and U8217 (N_8217,N_7444,N_7413);
nand U8218 (N_8218,N_7088,N_7294);
and U8219 (N_8219,N_7729,N_7934);
and U8220 (N_8220,N_7784,N_7459);
nor U8221 (N_8221,N_7136,N_7247);
or U8222 (N_8222,N_7504,N_7605);
and U8223 (N_8223,N_7192,N_7671);
nor U8224 (N_8224,N_7981,N_7226);
nor U8225 (N_8225,N_7065,N_7682);
and U8226 (N_8226,N_7275,N_7013);
nor U8227 (N_8227,N_7908,N_7234);
nand U8228 (N_8228,N_7936,N_7939);
or U8229 (N_8229,N_7950,N_7907);
or U8230 (N_8230,N_7404,N_7866);
or U8231 (N_8231,N_7006,N_7068);
nor U8232 (N_8232,N_7617,N_7516);
nor U8233 (N_8233,N_7553,N_7799);
or U8234 (N_8234,N_7422,N_7400);
or U8235 (N_8235,N_7546,N_7863);
or U8236 (N_8236,N_7987,N_7808);
and U8237 (N_8237,N_7712,N_7646);
and U8238 (N_8238,N_7297,N_7601);
or U8239 (N_8239,N_7138,N_7857);
and U8240 (N_8240,N_7057,N_7267);
nand U8241 (N_8241,N_7111,N_7619);
nor U8242 (N_8242,N_7287,N_7772);
nand U8243 (N_8243,N_7690,N_7733);
or U8244 (N_8244,N_7137,N_7163);
or U8245 (N_8245,N_7358,N_7099);
nor U8246 (N_8246,N_7623,N_7351);
nor U8247 (N_8247,N_7753,N_7697);
nand U8248 (N_8248,N_7498,N_7545);
xnor U8249 (N_8249,N_7789,N_7820);
and U8250 (N_8250,N_7035,N_7084);
nand U8251 (N_8251,N_7905,N_7458);
or U8252 (N_8252,N_7143,N_7746);
or U8253 (N_8253,N_7689,N_7391);
nand U8254 (N_8254,N_7921,N_7270);
or U8255 (N_8255,N_7566,N_7384);
or U8256 (N_8256,N_7894,N_7773);
and U8257 (N_8257,N_7231,N_7472);
nor U8258 (N_8258,N_7367,N_7684);
or U8259 (N_8259,N_7741,N_7114);
or U8260 (N_8260,N_7886,N_7154);
and U8261 (N_8261,N_7884,N_7973);
nor U8262 (N_8262,N_7061,N_7937);
nor U8263 (N_8263,N_7825,N_7115);
and U8264 (N_8264,N_7847,N_7368);
nand U8265 (N_8265,N_7800,N_7603);
and U8266 (N_8266,N_7798,N_7120);
and U8267 (N_8267,N_7376,N_7425);
and U8268 (N_8268,N_7538,N_7199);
xnor U8269 (N_8269,N_7024,N_7599);
or U8270 (N_8270,N_7364,N_7105);
xnor U8271 (N_8271,N_7207,N_7899);
nor U8272 (N_8272,N_7432,N_7175);
and U8273 (N_8273,N_7774,N_7214);
and U8274 (N_8274,N_7663,N_7734);
nand U8275 (N_8275,N_7510,N_7329);
or U8276 (N_8276,N_7356,N_7325);
or U8277 (N_8277,N_7874,N_7613);
nand U8278 (N_8278,N_7237,N_7834);
nor U8279 (N_8279,N_7274,N_7079);
and U8280 (N_8280,N_7423,N_7565);
nand U8281 (N_8281,N_7860,N_7327);
or U8282 (N_8282,N_7930,N_7853);
or U8283 (N_8283,N_7596,N_7206);
nor U8284 (N_8284,N_7686,N_7524);
or U8285 (N_8285,N_7642,N_7635);
xor U8286 (N_8286,N_7829,N_7321);
or U8287 (N_8287,N_7525,N_7067);
and U8288 (N_8288,N_7833,N_7691);
and U8289 (N_8289,N_7475,N_7428);
nor U8290 (N_8290,N_7058,N_7020);
and U8291 (N_8291,N_7708,N_7840);
or U8292 (N_8292,N_7025,N_7370);
and U8293 (N_8293,N_7507,N_7104);
nor U8294 (N_8294,N_7656,N_7761);
nand U8295 (N_8295,N_7172,N_7889);
nor U8296 (N_8296,N_7331,N_7268);
nand U8297 (N_8297,N_7312,N_7589);
nand U8298 (N_8298,N_7693,N_7448);
nand U8299 (N_8299,N_7787,N_7051);
nand U8300 (N_8300,N_7637,N_7177);
and U8301 (N_8301,N_7610,N_7867);
or U8302 (N_8302,N_7309,N_7452);
and U8303 (N_8303,N_7034,N_7306);
nor U8304 (N_8304,N_7917,N_7463);
or U8305 (N_8305,N_7091,N_7242);
or U8306 (N_8306,N_7131,N_7804);
and U8307 (N_8307,N_7766,N_7975);
xor U8308 (N_8308,N_7174,N_7781);
and U8309 (N_8309,N_7166,N_7958);
or U8310 (N_8310,N_7372,N_7393);
nand U8311 (N_8311,N_7014,N_7491);
nor U8312 (N_8312,N_7150,N_7527);
or U8313 (N_8313,N_7835,N_7298);
or U8314 (N_8314,N_7850,N_7724);
nand U8315 (N_8315,N_7241,N_7796);
nand U8316 (N_8316,N_7010,N_7169);
nand U8317 (N_8317,N_7503,N_7258);
or U8318 (N_8318,N_7830,N_7953);
nor U8319 (N_8319,N_7095,N_7332);
and U8320 (N_8320,N_7273,N_7782);
nor U8321 (N_8321,N_7935,N_7462);
or U8322 (N_8322,N_7480,N_7326);
nand U8323 (N_8323,N_7821,N_7558);
or U8324 (N_8324,N_7720,N_7081);
and U8325 (N_8325,N_7763,N_7622);
or U8326 (N_8326,N_7119,N_7162);
nand U8327 (N_8327,N_7755,N_7132);
and U8328 (N_8328,N_7967,N_7276);
or U8329 (N_8329,N_7385,N_7489);
nor U8330 (N_8330,N_7624,N_7052);
and U8331 (N_8331,N_7495,N_7576);
nand U8332 (N_8332,N_7221,N_7694);
and U8333 (N_8333,N_7345,N_7942);
nand U8334 (N_8334,N_7747,N_7122);
or U8335 (N_8335,N_7435,N_7901);
nor U8336 (N_8336,N_7337,N_7700);
or U8337 (N_8337,N_7238,N_7870);
nor U8338 (N_8338,N_7406,N_7028);
and U8339 (N_8339,N_7726,N_7250);
nand U8340 (N_8340,N_7036,N_7424);
nor U8341 (N_8341,N_7402,N_7033);
nor U8342 (N_8342,N_7993,N_7949);
nand U8343 (N_8343,N_7140,N_7396);
nand U8344 (N_8344,N_7378,N_7531);
and U8345 (N_8345,N_7359,N_7272);
nand U8346 (N_8346,N_7439,N_7490);
nor U8347 (N_8347,N_7389,N_7194);
or U8348 (N_8348,N_7509,N_7186);
nand U8349 (N_8349,N_7701,N_7911);
and U8350 (N_8350,N_7227,N_7305);
nand U8351 (N_8351,N_7968,N_7704);
or U8352 (N_8352,N_7293,N_7737);
or U8353 (N_8353,N_7461,N_7567);
and U8354 (N_8354,N_7429,N_7723);
nand U8355 (N_8355,N_7100,N_7366);
and U8356 (N_8356,N_7133,N_7518);
nand U8357 (N_8357,N_7643,N_7938);
and U8358 (N_8358,N_7240,N_7611);
nand U8359 (N_8359,N_7838,N_7536);
and U8360 (N_8360,N_7906,N_7478);
and U8361 (N_8361,N_7244,N_7989);
nor U8362 (N_8362,N_7262,N_7947);
or U8363 (N_8363,N_7303,N_7295);
nor U8364 (N_8364,N_7869,N_7314);
and U8365 (N_8365,N_7855,N_7263);
or U8366 (N_8366,N_7233,N_7285);
nand U8367 (N_8367,N_7846,N_7042);
and U8368 (N_8368,N_7715,N_7598);
or U8369 (N_8369,N_7373,N_7330);
or U8370 (N_8370,N_7251,N_7414);
or U8371 (N_8371,N_7291,N_7962);
and U8372 (N_8372,N_7591,N_7069);
and U8373 (N_8373,N_7255,N_7828);
and U8374 (N_8374,N_7890,N_7371);
nand U8375 (N_8375,N_7607,N_7055);
and U8376 (N_8376,N_7711,N_7770);
nand U8377 (N_8377,N_7571,N_7005);
and U8378 (N_8378,N_7197,N_7929);
nand U8379 (N_8379,N_7716,N_7505);
or U8380 (N_8380,N_7986,N_7983);
nand U8381 (N_8381,N_7895,N_7706);
nor U8382 (N_8382,N_7283,N_7990);
or U8383 (N_8383,N_7352,N_7271);
nand U8384 (N_8384,N_7399,N_7347);
and U8385 (N_8385,N_7205,N_7956);
nor U8386 (N_8386,N_7261,N_7212);
or U8387 (N_8387,N_7338,N_7420);
and U8388 (N_8388,N_7535,N_7464);
or U8389 (N_8389,N_7494,N_7519);
and U8390 (N_8390,N_7315,N_7943);
nor U8391 (N_8391,N_7260,N_7717);
and U8392 (N_8392,N_7748,N_7045);
nor U8393 (N_8393,N_7856,N_7547);
and U8394 (N_8394,N_7652,N_7335);
nand U8395 (N_8395,N_7151,N_7198);
nand U8396 (N_8396,N_7292,N_7070);
nand U8397 (N_8397,N_7526,N_7876);
xnor U8398 (N_8398,N_7211,N_7302);
and U8399 (N_8399,N_7585,N_7562);
nand U8400 (N_8400,N_7730,N_7976);
nor U8401 (N_8401,N_7265,N_7442);
or U8402 (N_8402,N_7728,N_7257);
and U8403 (N_8403,N_7408,N_7854);
and U8404 (N_8404,N_7780,N_7606);
or U8405 (N_8405,N_7560,N_7073);
nor U8406 (N_8406,N_7360,N_7213);
nor U8407 (N_8407,N_7094,N_7848);
and U8408 (N_8408,N_7951,N_7202);
nor U8409 (N_8409,N_7259,N_7209);
and U8410 (N_8410,N_7096,N_7109);
nand U8411 (N_8411,N_7561,N_7008);
or U8412 (N_8412,N_7573,N_7634);
nand U8413 (N_8413,N_7235,N_7946);
or U8414 (N_8414,N_7401,N_7219);
xnor U8415 (N_8415,N_7552,N_7455);
and U8416 (N_8416,N_7892,N_7649);
nand U8417 (N_8417,N_7852,N_7725);
or U8418 (N_8418,N_7978,N_7029);
and U8419 (N_8419,N_7631,N_7015);
or U8420 (N_8420,N_7897,N_7348);
nand U8421 (N_8421,N_7645,N_7392);
or U8422 (N_8422,N_7223,N_7217);
or U8423 (N_8423,N_7220,N_7718);
and U8424 (N_8424,N_7106,N_7831);
nand U8425 (N_8425,N_7769,N_7426);
nor U8426 (N_8426,N_7961,N_7873);
and U8427 (N_8427,N_7144,N_7123);
nand U8428 (N_8428,N_7636,N_7685);
nor U8429 (N_8429,N_7196,N_7044);
or U8430 (N_8430,N_7155,N_7583);
or U8431 (N_8431,N_7168,N_7801);
nand U8432 (N_8432,N_7994,N_7374);
nand U8433 (N_8433,N_7245,N_7940);
nand U8434 (N_8434,N_7103,N_7625);
nor U8435 (N_8435,N_7493,N_7676);
nor U8436 (N_8436,N_7179,N_7520);
and U8437 (N_8437,N_7638,N_7707);
nor U8438 (N_8438,N_7739,N_7125);
nand U8439 (N_8439,N_7433,N_7824);
nand U8440 (N_8440,N_7803,N_7595);
or U8441 (N_8441,N_7222,N_7117);
nor U8442 (N_8442,N_7980,N_7007);
nor U8443 (N_8443,N_7816,N_7466);
nor U8444 (N_8444,N_7764,N_7066);
and U8445 (N_8445,N_7216,N_7085);
and U8446 (N_8446,N_7016,N_7112);
and U8447 (N_8447,N_7397,N_7932);
nand U8448 (N_8448,N_7999,N_7972);
and U8449 (N_8449,N_7281,N_7688);
nand U8450 (N_8450,N_7514,N_7145);
nand U8451 (N_8451,N_7765,N_7328);
and U8452 (N_8452,N_7477,N_7687);
nor U8453 (N_8453,N_7208,N_7742);
and U8454 (N_8454,N_7484,N_7158);
or U8455 (N_8455,N_7333,N_7296);
and U8456 (N_8456,N_7388,N_7814);
or U8457 (N_8457,N_7555,N_7394);
and U8458 (N_8458,N_7740,N_7215);
nor U8459 (N_8459,N_7896,N_7344);
nand U8460 (N_8460,N_7108,N_7970);
nand U8461 (N_8461,N_7851,N_7277);
and U8462 (N_8462,N_7354,N_7418);
nand U8463 (N_8463,N_7012,N_7559);
and U8464 (N_8464,N_7340,N_7415);
nor U8465 (N_8465,N_7754,N_7476);
nor U8466 (N_8466,N_7349,N_7826);
or U8467 (N_8467,N_7750,N_7059);
nand U8468 (N_8468,N_7672,N_7577);
nor U8469 (N_8469,N_7819,N_7818);
and U8470 (N_8470,N_7307,N_7512);
xnor U8471 (N_8471,N_7203,N_7139);
nor U8472 (N_8472,N_7681,N_7440);
nand U8473 (N_8473,N_7499,N_7557);
or U8474 (N_8474,N_7620,N_7931);
nor U8475 (N_8475,N_7815,N_7187);
nand U8476 (N_8476,N_7224,N_7204);
nor U8477 (N_8477,N_7861,N_7236);
nand U8478 (N_8478,N_7597,N_7201);
nand U8479 (N_8479,N_7522,N_7021);
nor U8480 (N_8480,N_7243,N_7311);
nor U8481 (N_8481,N_7153,N_7090);
nor U8482 (N_8482,N_7670,N_7699);
or U8483 (N_8483,N_7116,N_7500);
nor U8484 (N_8484,N_7647,N_7000);
nand U8485 (N_8485,N_7530,N_7288);
or U8486 (N_8486,N_7779,N_7102);
nand U8487 (N_8487,N_7048,N_7481);
nor U8488 (N_8488,N_7683,N_7783);
nand U8489 (N_8489,N_7098,N_7872);
and U8490 (N_8490,N_7927,N_7608);
nor U8491 (N_8491,N_7794,N_7113);
and U8492 (N_8492,N_7210,N_7353);
nand U8493 (N_8493,N_7430,N_7984);
and U8494 (N_8494,N_7050,N_7767);
nor U8495 (N_8495,N_7317,N_7540);
nor U8496 (N_8496,N_7542,N_7170);
and U8497 (N_8497,N_7673,N_7280);
and U8498 (N_8498,N_7778,N_7124);
nand U8499 (N_8499,N_7176,N_7171);
or U8500 (N_8500,N_7644,N_7414);
and U8501 (N_8501,N_7393,N_7216);
and U8502 (N_8502,N_7914,N_7815);
or U8503 (N_8503,N_7970,N_7870);
nor U8504 (N_8504,N_7852,N_7538);
nand U8505 (N_8505,N_7161,N_7504);
or U8506 (N_8506,N_7243,N_7483);
nor U8507 (N_8507,N_7040,N_7392);
nand U8508 (N_8508,N_7621,N_7598);
nand U8509 (N_8509,N_7258,N_7027);
nor U8510 (N_8510,N_7735,N_7754);
or U8511 (N_8511,N_7742,N_7260);
and U8512 (N_8512,N_7140,N_7615);
nand U8513 (N_8513,N_7809,N_7674);
nand U8514 (N_8514,N_7141,N_7070);
or U8515 (N_8515,N_7153,N_7564);
nor U8516 (N_8516,N_7789,N_7388);
nor U8517 (N_8517,N_7425,N_7645);
nand U8518 (N_8518,N_7374,N_7658);
nor U8519 (N_8519,N_7074,N_7011);
or U8520 (N_8520,N_7238,N_7847);
nor U8521 (N_8521,N_7720,N_7310);
nor U8522 (N_8522,N_7432,N_7791);
and U8523 (N_8523,N_7975,N_7273);
nand U8524 (N_8524,N_7499,N_7119);
nor U8525 (N_8525,N_7203,N_7404);
nor U8526 (N_8526,N_7432,N_7792);
and U8527 (N_8527,N_7833,N_7396);
xnor U8528 (N_8528,N_7225,N_7160);
nand U8529 (N_8529,N_7243,N_7630);
and U8530 (N_8530,N_7166,N_7204);
and U8531 (N_8531,N_7340,N_7697);
or U8532 (N_8532,N_7265,N_7898);
and U8533 (N_8533,N_7417,N_7309);
or U8534 (N_8534,N_7159,N_7116);
or U8535 (N_8535,N_7370,N_7876);
nor U8536 (N_8536,N_7572,N_7640);
or U8537 (N_8537,N_7348,N_7264);
nand U8538 (N_8538,N_7448,N_7465);
nor U8539 (N_8539,N_7933,N_7541);
and U8540 (N_8540,N_7359,N_7369);
nor U8541 (N_8541,N_7979,N_7841);
and U8542 (N_8542,N_7415,N_7411);
nand U8543 (N_8543,N_7126,N_7899);
nor U8544 (N_8544,N_7167,N_7583);
and U8545 (N_8545,N_7526,N_7956);
or U8546 (N_8546,N_7742,N_7675);
nor U8547 (N_8547,N_7741,N_7229);
nand U8548 (N_8548,N_7447,N_7407);
nand U8549 (N_8549,N_7872,N_7893);
nand U8550 (N_8550,N_7357,N_7005);
and U8551 (N_8551,N_7675,N_7869);
xor U8552 (N_8552,N_7321,N_7276);
and U8553 (N_8553,N_7329,N_7309);
nand U8554 (N_8554,N_7725,N_7650);
nor U8555 (N_8555,N_7878,N_7730);
nor U8556 (N_8556,N_7295,N_7575);
nor U8557 (N_8557,N_7152,N_7385);
or U8558 (N_8558,N_7034,N_7516);
or U8559 (N_8559,N_7013,N_7404);
xor U8560 (N_8560,N_7326,N_7904);
nor U8561 (N_8561,N_7087,N_7800);
nand U8562 (N_8562,N_7119,N_7559);
or U8563 (N_8563,N_7261,N_7621);
nor U8564 (N_8564,N_7312,N_7388);
nand U8565 (N_8565,N_7617,N_7153);
and U8566 (N_8566,N_7037,N_7169);
nor U8567 (N_8567,N_7128,N_7620);
and U8568 (N_8568,N_7553,N_7824);
and U8569 (N_8569,N_7930,N_7160);
and U8570 (N_8570,N_7861,N_7867);
or U8571 (N_8571,N_7817,N_7595);
nor U8572 (N_8572,N_7238,N_7856);
and U8573 (N_8573,N_7240,N_7958);
and U8574 (N_8574,N_7618,N_7826);
and U8575 (N_8575,N_7162,N_7280);
or U8576 (N_8576,N_7007,N_7868);
or U8577 (N_8577,N_7668,N_7399);
nand U8578 (N_8578,N_7886,N_7142);
or U8579 (N_8579,N_7100,N_7532);
nand U8580 (N_8580,N_7829,N_7503);
nor U8581 (N_8581,N_7679,N_7585);
and U8582 (N_8582,N_7308,N_7715);
or U8583 (N_8583,N_7616,N_7902);
nor U8584 (N_8584,N_7349,N_7509);
nand U8585 (N_8585,N_7080,N_7319);
or U8586 (N_8586,N_7435,N_7053);
and U8587 (N_8587,N_7839,N_7348);
and U8588 (N_8588,N_7073,N_7027);
nor U8589 (N_8589,N_7645,N_7122);
and U8590 (N_8590,N_7696,N_7069);
or U8591 (N_8591,N_7606,N_7054);
or U8592 (N_8592,N_7743,N_7269);
or U8593 (N_8593,N_7444,N_7910);
and U8594 (N_8594,N_7584,N_7743);
nand U8595 (N_8595,N_7559,N_7138);
or U8596 (N_8596,N_7308,N_7411);
nor U8597 (N_8597,N_7554,N_7898);
and U8598 (N_8598,N_7955,N_7099);
nor U8599 (N_8599,N_7362,N_7578);
and U8600 (N_8600,N_7812,N_7216);
nand U8601 (N_8601,N_7281,N_7694);
nand U8602 (N_8602,N_7558,N_7979);
and U8603 (N_8603,N_7327,N_7435);
nand U8604 (N_8604,N_7402,N_7826);
nand U8605 (N_8605,N_7907,N_7099);
nand U8606 (N_8606,N_7666,N_7085);
nand U8607 (N_8607,N_7493,N_7266);
nand U8608 (N_8608,N_7532,N_7238);
and U8609 (N_8609,N_7920,N_7892);
or U8610 (N_8610,N_7572,N_7488);
or U8611 (N_8611,N_7073,N_7960);
nor U8612 (N_8612,N_7651,N_7185);
or U8613 (N_8613,N_7587,N_7446);
nand U8614 (N_8614,N_7027,N_7532);
or U8615 (N_8615,N_7397,N_7994);
or U8616 (N_8616,N_7336,N_7507);
and U8617 (N_8617,N_7556,N_7781);
nand U8618 (N_8618,N_7246,N_7334);
and U8619 (N_8619,N_7315,N_7961);
or U8620 (N_8620,N_7844,N_7693);
and U8621 (N_8621,N_7075,N_7062);
nand U8622 (N_8622,N_7071,N_7070);
or U8623 (N_8623,N_7233,N_7744);
and U8624 (N_8624,N_7539,N_7172);
nor U8625 (N_8625,N_7412,N_7000);
and U8626 (N_8626,N_7339,N_7470);
or U8627 (N_8627,N_7403,N_7098);
nand U8628 (N_8628,N_7304,N_7154);
nand U8629 (N_8629,N_7115,N_7850);
nor U8630 (N_8630,N_7992,N_7767);
nand U8631 (N_8631,N_7758,N_7263);
or U8632 (N_8632,N_7249,N_7084);
nor U8633 (N_8633,N_7948,N_7161);
or U8634 (N_8634,N_7417,N_7132);
or U8635 (N_8635,N_7023,N_7280);
nand U8636 (N_8636,N_7227,N_7169);
or U8637 (N_8637,N_7358,N_7243);
or U8638 (N_8638,N_7046,N_7821);
or U8639 (N_8639,N_7933,N_7555);
or U8640 (N_8640,N_7105,N_7104);
nor U8641 (N_8641,N_7090,N_7801);
nor U8642 (N_8642,N_7452,N_7326);
or U8643 (N_8643,N_7736,N_7304);
xnor U8644 (N_8644,N_7998,N_7940);
or U8645 (N_8645,N_7272,N_7457);
nand U8646 (N_8646,N_7569,N_7923);
or U8647 (N_8647,N_7086,N_7954);
nor U8648 (N_8648,N_7858,N_7451);
and U8649 (N_8649,N_7588,N_7947);
and U8650 (N_8650,N_7219,N_7654);
or U8651 (N_8651,N_7529,N_7403);
and U8652 (N_8652,N_7195,N_7163);
nor U8653 (N_8653,N_7002,N_7434);
nand U8654 (N_8654,N_7619,N_7135);
or U8655 (N_8655,N_7418,N_7470);
or U8656 (N_8656,N_7838,N_7682);
and U8657 (N_8657,N_7096,N_7361);
or U8658 (N_8658,N_7712,N_7323);
nor U8659 (N_8659,N_7404,N_7461);
nand U8660 (N_8660,N_7209,N_7034);
xor U8661 (N_8661,N_7306,N_7405);
and U8662 (N_8662,N_7833,N_7746);
and U8663 (N_8663,N_7631,N_7775);
or U8664 (N_8664,N_7961,N_7272);
and U8665 (N_8665,N_7745,N_7404);
nor U8666 (N_8666,N_7812,N_7360);
nor U8667 (N_8667,N_7300,N_7587);
nand U8668 (N_8668,N_7274,N_7638);
nor U8669 (N_8669,N_7617,N_7808);
or U8670 (N_8670,N_7152,N_7636);
nand U8671 (N_8671,N_7440,N_7576);
nor U8672 (N_8672,N_7762,N_7680);
and U8673 (N_8673,N_7264,N_7279);
nor U8674 (N_8674,N_7021,N_7763);
nand U8675 (N_8675,N_7138,N_7166);
nor U8676 (N_8676,N_7536,N_7829);
and U8677 (N_8677,N_7752,N_7211);
nand U8678 (N_8678,N_7127,N_7872);
nor U8679 (N_8679,N_7153,N_7242);
and U8680 (N_8680,N_7512,N_7864);
or U8681 (N_8681,N_7566,N_7530);
nor U8682 (N_8682,N_7190,N_7242);
nand U8683 (N_8683,N_7876,N_7102);
nand U8684 (N_8684,N_7358,N_7661);
nor U8685 (N_8685,N_7673,N_7544);
nor U8686 (N_8686,N_7878,N_7659);
nor U8687 (N_8687,N_7330,N_7807);
nor U8688 (N_8688,N_7819,N_7682);
nand U8689 (N_8689,N_7620,N_7380);
nor U8690 (N_8690,N_7306,N_7207);
nor U8691 (N_8691,N_7656,N_7900);
nor U8692 (N_8692,N_7126,N_7759);
nand U8693 (N_8693,N_7358,N_7522);
nand U8694 (N_8694,N_7336,N_7441);
nand U8695 (N_8695,N_7622,N_7785);
and U8696 (N_8696,N_7276,N_7329);
and U8697 (N_8697,N_7550,N_7911);
nor U8698 (N_8698,N_7469,N_7717);
or U8699 (N_8699,N_7889,N_7121);
or U8700 (N_8700,N_7852,N_7345);
and U8701 (N_8701,N_7903,N_7644);
nor U8702 (N_8702,N_7435,N_7179);
or U8703 (N_8703,N_7442,N_7659);
nor U8704 (N_8704,N_7194,N_7232);
or U8705 (N_8705,N_7700,N_7661);
nor U8706 (N_8706,N_7717,N_7521);
and U8707 (N_8707,N_7062,N_7808);
and U8708 (N_8708,N_7086,N_7552);
nand U8709 (N_8709,N_7824,N_7919);
nand U8710 (N_8710,N_7415,N_7690);
nor U8711 (N_8711,N_7574,N_7341);
xnor U8712 (N_8712,N_7301,N_7723);
and U8713 (N_8713,N_7088,N_7208);
and U8714 (N_8714,N_7095,N_7228);
or U8715 (N_8715,N_7558,N_7652);
or U8716 (N_8716,N_7220,N_7166);
nor U8717 (N_8717,N_7272,N_7291);
nand U8718 (N_8718,N_7706,N_7109);
and U8719 (N_8719,N_7127,N_7833);
nor U8720 (N_8720,N_7120,N_7053);
nand U8721 (N_8721,N_7894,N_7393);
nand U8722 (N_8722,N_7595,N_7409);
and U8723 (N_8723,N_7109,N_7225);
or U8724 (N_8724,N_7308,N_7733);
nor U8725 (N_8725,N_7654,N_7027);
and U8726 (N_8726,N_7692,N_7350);
nand U8727 (N_8727,N_7136,N_7278);
or U8728 (N_8728,N_7064,N_7558);
nor U8729 (N_8729,N_7105,N_7257);
nand U8730 (N_8730,N_7101,N_7054);
nor U8731 (N_8731,N_7713,N_7115);
nor U8732 (N_8732,N_7298,N_7305);
nor U8733 (N_8733,N_7321,N_7187);
and U8734 (N_8734,N_7595,N_7533);
and U8735 (N_8735,N_7607,N_7097);
nand U8736 (N_8736,N_7332,N_7200);
nand U8737 (N_8737,N_7797,N_7147);
nand U8738 (N_8738,N_7556,N_7526);
nand U8739 (N_8739,N_7497,N_7454);
nand U8740 (N_8740,N_7828,N_7822);
and U8741 (N_8741,N_7246,N_7526);
nor U8742 (N_8742,N_7746,N_7857);
or U8743 (N_8743,N_7554,N_7436);
and U8744 (N_8744,N_7813,N_7828);
nor U8745 (N_8745,N_7830,N_7726);
and U8746 (N_8746,N_7980,N_7559);
nand U8747 (N_8747,N_7873,N_7739);
and U8748 (N_8748,N_7479,N_7524);
and U8749 (N_8749,N_7493,N_7428);
nand U8750 (N_8750,N_7265,N_7803);
nand U8751 (N_8751,N_7675,N_7579);
nand U8752 (N_8752,N_7594,N_7868);
nor U8753 (N_8753,N_7068,N_7751);
nor U8754 (N_8754,N_7062,N_7339);
and U8755 (N_8755,N_7580,N_7968);
and U8756 (N_8756,N_7463,N_7683);
xnor U8757 (N_8757,N_7789,N_7946);
nor U8758 (N_8758,N_7636,N_7728);
or U8759 (N_8759,N_7402,N_7703);
nand U8760 (N_8760,N_7543,N_7523);
nor U8761 (N_8761,N_7451,N_7006);
or U8762 (N_8762,N_7889,N_7249);
and U8763 (N_8763,N_7660,N_7779);
nor U8764 (N_8764,N_7524,N_7332);
or U8765 (N_8765,N_7073,N_7958);
nor U8766 (N_8766,N_7646,N_7896);
nand U8767 (N_8767,N_7008,N_7529);
or U8768 (N_8768,N_7865,N_7394);
nand U8769 (N_8769,N_7364,N_7204);
nor U8770 (N_8770,N_7057,N_7909);
nand U8771 (N_8771,N_7996,N_7919);
or U8772 (N_8772,N_7432,N_7430);
nor U8773 (N_8773,N_7128,N_7493);
and U8774 (N_8774,N_7860,N_7322);
nand U8775 (N_8775,N_7235,N_7683);
and U8776 (N_8776,N_7056,N_7992);
nand U8777 (N_8777,N_7662,N_7158);
and U8778 (N_8778,N_7947,N_7887);
and U8779 (N_8779,N_7820,N_7857);
nor U8780 (N_8780,N_7839,N_7827);
and U8781 (N_8781,N_7020,N_7029);
and U8782 (N_8782,N_7292,N_7305);
nor U8783 (N_8783,N_7597,N_7438);
or U8784 (N_8784,N_7887,N_7721);
or U8785 (N_8785,N_7136,N_7200);
and U8786 (N_8786,N_7251,N_7449);
nand U8787 (N_8787,N_7978,N_7519);
nand U8788 (N_8788,N_7766,N_7805);
nor U8789 (N_8789,N_7990,N_7579);
nand U8790 (N_8790,N_7077,N_7902);
or U8791 (N_8791,N_7967,N_7971);
and U8792 (N_8792,N_7219,N_7299);
and U8793 (N_8793,N_7667,N_7672);
or U8794 (N_8794,N_7369,N_7544);
or U8795 (N_8795,N_7175,N_7717);
nand U8796 (N_8796,N_7668,N_7051);
or U8797 (N_8797,N_7754,N_7195);
and U8798 (N_8798,N_7058,N_7082);
nor U8799 (N_8799,N_7127,N_7147);
or U8800 (N_8800,N_7296,N_7620);
nor U8801 (N_8801,N_7317,N_7364);
or U8802 (N_8802,N_7965,N_7091);
and U8803 (N_8803,N_7621,N_7519);
and U8804 (N_8804,N_7215,N_7883);
and U8805 (N_8805,N_7924,N_7225);
or U8806 (N_8806,N_7745,N_7052);
and U8807 (N_8807,N_7895,N_7225);
and U8808 (N_8808,N_7881,N_7442);
nand U8809 (N_8809,N_7873,N_7372);
and U8810 (N_8810,N_7946,N_7625);
nand U8811 (N_8811,N_7609,N_7989);
nor U8812 (N_8812,N_7438,N_7742);
nand U8813 (N_8813,N_7869,N_7263);
nand U8814 (N_8814,N_7240,N_7831);
or U8815 (N_8815,N_7191,N_7880);
and U8816 (N_8816,N_7757,N_7452);
and U8817 (N_8817,N_7799,N_7129);
nand U8818 (N_8818,N_7201,N_7174);
nand U8819 (N_8819,N_7171,N_7774);
nand U8820 (N_8820,N_7217,N_7406);
or U8821 (N_8821,N_7079,N_7135);
nand U8822 (N_8822,N_7073,N_7112);
and U8823 (N_8823,N_7224,N_7678);
or U8824 (N_8824,N_7822,N_7596);
or U8825 (N_8825,N_7695,N_7704);
nor U8826 (N_8826,N_7247,N_7033);
nand U8827 (N_8827,N_7078,N_7161);
nor U8828 (N_8828,N_7510,N_7629);
and U8829 (N_8829,N_7252,N_7587);
nor U8830 (N_8830,N_7753,N_7271);
nor U8831 (N_8831,N_7586,N_7455);
nand U8832 (N_8832,N_7588,N_7022);
or U8833 (N_8833,N_7456,N_7504);
and U8834 (N_8834,N_7614,N_7354);
and U8835 (N_8835,N_7769,N_7531);
nand U8836 (N_8836,N_7152,N_7117);
nand U8837 (N_8837,N_7665,N_7515);
nor U8838 (N_8838,N_7339,N_7411);
and U8839 (N_8839,N_7982,N_7757);
and U8840 (N_8840,N_7800,N_7067);
or U8841 (N_8841,N_7407,N_7366);
nand U8842 (N_8842,N_7985,N_7792);
xnor U8843 (N_8843,N_7055,N_7967);
and U8844 (N_8844,N_7043,N_7390);
nand U8845 (N_8845,N_7764,N_7399);
nand U8846 (N_8846,N_7484,N_7894);
and U8847 (N_8847,N_7373,N_7157);
nand U8848 (N_8848,N_7480,N_7093);
nand U8849 (N_8849,N_7574,N_7330);
and U8850 (N_8850,N_7124,N_7927);
nand U8851 (N_8851,N_7476,N_7453);
nand U8852 (N_8852,N_7729,N_7073);
or U8853 (N_8853,N_7253,N_7430);
and U8854 (N_8854,N_7546,N_7311);
nand U8855 (N_8855,N_7356,N_7723);
nand U8856 (N_8856,N_7665,N_7613);
or U8857 (N_8857,N_7891,N_7103);
nor U8858 (N_8858,N_7308,N_7266);
and U8859 (N_8859,N_7841,N_7032);
or U8860 (N_8860,N_7384,N_7776);
and U8861 (N_8861,N_7252,N_7152);
or U8862 (N_8862,N_7882,N_7938);
nand U8863 (N_8863,N_7355,N_7011);
nor U8864 (N_8864,N_7656,N_7910);
nor U8865 (N_8865,N_7654,N_7071);
nand U8866 (N_8866,N_7903,N_7769);
and U8867 (N_8867,N_7307,N_7598);
and U8868 (N_8868,N_7675,N_7272);
nor U8869 (N_8869,N_7348,N_7838);
or U8870 (N_8870,N_7914,N_7929);
nor U8871 (N_8871,N_7729,N_7651);
nand U8872 (N_8872,N_7174,N_7909);
and U8873 (N_8873,N_7005,N_7580);
nor U8874 (N_8874,N_7931,N_7941);
nand U8875 (N_8875,N_7553,N_7060);
nor U8876 (N_8876,N_7786,N_7633);
nor U8877 (N_8877,N_7913,N_7657);
and U8878 (N_8878,N_7772,N_7537);
nand U8879 (N_8879,N_7743,N_7137);
and U8880 (N_8880,N_7766,N_7815);
or U8881 (N_8881,N_7326,N_7648);
nor U8882 (N_8882,N_7712,N_7051);
and U8883 (N_8883,N_7675,N_7746);
nand U8884 (N_8884,N_7268,N_7567);
nor U8885 (N_8885,N_7959,N_7990);
nand U8886 (N_8886,N_7176,N_7905);
or U8887 (N_8887,N_7147,N_7247);
or U8888 (N_8888,N_7195,N_7442);
nor U8889 (N_8889,N_7072,N_7488);
nor U8890 (N_8890,N_7816,N_7919);
nor U8891 (N_8891,N_7450,N_7769);
nand U8892 (N_8892,N_7821,N_7516);
or U8893 (N_8893,N_7496,N_7152);
and U8894 (N_8894,N_7950,N_7250);
and U8895 (N_8895,N_7639,N_7470);
xor U8896 (N_8896,N_7040,N_7987);
nand U8897 (N_8897,N_7838,N_7113);
nand U8898 (N_8898,N_7292,N_7128);
and U8899 (N_8899,N_7623,N_7881);
nor U8900 (N_8900,N_7759,N_7565);
nand U8901 (N_8901,N_7476,N_7100);
or U8902 (N_8902,N_7987,N_7016);
or U8903 (N_8903,N_7555,N_7870);
or U8904 (N_8904,N_7593,N_7135);
and U8905 (N_8905,N_7262,N_7665);
nand U8906 (N_8906,N_7032,N_7291);
or U8907 (N_8907,N_7069,N_7329);
nand U8908 (N_8908,N_7532,N_7800);
nor U8909 (N_8909,N_7549,N_7457);
nor U8910 (N_8910,N_7061,N_7132);
or U8911 (N_8911,N_7862,N_7570);
nand U8912 (N_8912,N_7619,N_7022);
nor U8913 (N_8913,N_7074,N_7878);
nand U8914 (N_8914,N_7672,N_7684);
and U8915 (N_8915,N_7729,N_7356);
and U8916 (N_8916,N_7776,N_7775);
nor U8917 (N_8917,N_7205,N_7258);
and U8918 (N_8918,N_7482,N_7441);
nand U8919 (N_8919,N_7146,N_7630);
and U8920 (N_8920,N_7147,N_7653);
and U8921 (N_8921,N_7615,N_7183);
nor U8922 (N_8922,N_7680,N_7811);
nor U8923 (N_8923,N_7464,N_7042);
nor U8924 (N_8924,N_7862,N_7972);
or U8925 (N_8925,N_7413,N_7038);
or U8926 (N_8926,N_7009,N_7786);
or U8927 (N_8927,N_7688,N_7273);
or U8928 (N_8928,N_7798,N_7291);
nand U8929 (N_8929,N_7822,N_7146);
or U8930 (N_8930,N_7377,N_7741);
and U8931 (N_8931,N_7717,N_7333);
nand U8932 (N_8932,N_7622,N_7255);
nand U8933 (N_8933,N_7520,N_7483);
or U8934 (N_8934,N_7708,N_7834);
nand U8935 (N_8935,N_7801,N_7176);
nor U8936 (N_8936,N_7357,N_7496);
and U8937 (N_8937,N_7094,N_7339);
and U8938 (N_8938,N_7995,N_7425);
or U8939 (N_8939,N_7300,N_7690);
nand U8940 (N_8940,N_7767,N_7732);
or U8941 (N_8941,N_7936,N_7010);
nand U8942 (N_8942,N_7935,N_7191);
nand U8943 (N_8943,N_7027,N_7414);
nand U8944 (N_8944,N_7575,N_7354);
nor U8945 (N_8945,N_7457,N_7748);
or U8946 (N_8946,N_7172,N_7086);
nand U8947 (N_8947,N_7690,N_7325);
and U8948 (N_8948,N_7082,N_7291);
or U8949 (N_8949,N_7360,N_7055);
nor U8950 (N_8950,N_7884,N_7918);
nand U8951 (N_8951,N_7261,N_7682);
nand U8952 (N_8952,N_7697,N_7198);
nand U8953 (N_8953,N_7562,N_7231);
or U8954 (N_8954,N_7613,N_7223);
and U8955 (N_8955,N_7942,N_7891);
nand U8956 (N_8956,N_7170,N_7093);
nand U8957 (N_8957,N_7688,N_7824);
and U8958 (N_8958,N_7729,N_7498);
or U8959 (N_8959,N_7574,N_7865);
nand U8960 (N_8960,N_7375,N_7945);
nor U8961 (N_8961,N_7612,N_7529);
or U8962 (N_8962,N_7661,N_7539);
and U8963 (N_8963,N_7932,N_7339);
and U8964 (N_8964,N_7910,N_7189);
and U8965 (N_8965,N_7751,N_7714);
and U8966 (N_8966,N_7535,N_7910);
nor U8967 (N_8967,N_7424,N_7613);
nor U8968 (N_8968,N_7991,N_7577);
and U8969 (N_8969,N_7404,N_7444);
nor U8970 (N_8970,N_7967,N_7102);
and U8971 (N_8971,N_7666,N_7491);
nand U8972 (N_8972,N_7133,N_7976);
or U8973 (N_8973,N_7320,N_7316);
nand U8974 (N_8974,N_7260,N_7647);
or U8975 (N_8975,N_7469,N_7666);
nor U8976 (N_8976,N_7547,N_7130);
or U8977 (N_8977,N_7258,N_7593);
and U8978 (N_8978,N_7540,N_7528);
or U8979 (N_8979,N_7146,N_7798);
and U8980 (N_8980,N_7605,N_7542);
nand U8981 (N_8981,N_7576,N_7256);
nor U8982 (N_8982,N_7673,N_7005);
or U8983 (N_8983,N_7680,N_7532);
nor U8984 (N_8984,N_7822,N_7259);
or U8985 (N_8985,N_7998,N_7897);
nand U8986 (N_8986,N_7086,N_7429);
nand U8987 (N_8987,N_7977,N_7972);
and U8988 (N_8988,N_7225,N_7745);
nor U8989 (N_8989,N_7776,N_7475);
and U8990 (N_8990,N_7813,N_7248);
and U8991 (N_8991,N_7916,N_7401);
nand U8992 (N_8992,N_7562,N_7275);
or U8993 (N_8993,N_7304,N_7068);
and U8994 (N_8994,N_7926,N_7788);
or U8995 (N_8995,N_7868,N_7923);
nand U8996 (N_8996,N_7779,N_7972);
nand U8997 (N_8997,N_7282,N_7247);
or U8998 (N_8998,N_7350,N_7768);
nor U8999 (N_8999,N_7375,N_7898);
nor U9000 (N_9000,N_8063,N_8720);
nor U9001 (N_9001,N_8170,N_8835);
and U9002 (N_9002,N_8397,N_8301);
nor U9003 (N_9003,N_8084,N_8514);
nor U9004 (N_9004,N_8161,N_8991);
nand U9005 (N_9005,N_8249,N_8127);
and U9006 (N_9006,N_8052,N_8317);
nand U9007 (N_9007,N_8351,N_8340);
or U9008 (N_9008,N_8878,N_8474);
nand U9009 (N_9009,N_8173,N_8768);
nor U9010 (N_9010,N_8691,N_8714);
nor U9011 (N_9011,N_8056,N_8080);
nor U9012 (N_9012,N_8907,N_8734);
nand U9013 (N_9013,N_8130,N_8954);
and U9014 (N_9014,N_8535,N_8430);
nor U9015 (N_9015,N_8947,N_8431);
and U9016 (N_9016,N_8944,N_8721);
and U9017 (N_9017,N_8157,N_8282);
and U9018 (N_9018,N_8796,N_8264);
nor U9019 (N_9019,N_8769,N_8632);
nor U9020 (N_9020,N_8412,N_8744);
or U9021 (N_9021,N_8837,N_8812);
nand U9022 (N_9022,N_8700,N_8171);
or U9023 (N_9023,N_8682,N_8808);
and U9024 (N_9024,N_8458,N_8990);
and U9025 (N_9025,N_8165,N_8386);
or U9026 (N_9026,N_8807,N_8135);
nand U9027 (N_9027,N_8472,N_8133);
and U9028 (N_9028,N_8091,N_8755);
nor U9029 (N_9029,N_8746,N_8414);
or U9030 (N_9030,N_8492,N_8302);
nand U9031 (N_9031,N_8176,N_8263);
nor U9032 (N_9032,N_8996,N_8434);
or U9033 (N_9033,N_8220,N_8110);
xor U9034 (N_9034,N_8087,N_8182);
or U9035 (N_9035,N_8693,N_8490);
nor U9036 (N_9036,N_8992,N_8318);
nor U9037 (N_9037,N_8899,N_8191);
and U9038 (N_9038,N_8373,N_8497);
nand U9039 (N_9039,N_8071,N_8113);
nor U9040 (N_9040,N_8505,N_8801);
xnor U9041 (N_9041,N_8209,N_8009);
and U9042 (N_9042,N_8297,N_8387);
and U9043 (N_9043,N_8903,N_8851);
or U9044 (N_9044,N_8201,N_8399);
or U9045 (N_9045,N_8262,N_8139);
nor U9046 (N_9046,N_8315,N_8172);
and U9047 (N_9047,N_8998,N_8369);
and U9048 (N_9048,N_8537,N_8293);
nand U9049 (N_9049,N_8076,N_8875);
and U9050 (N_9050,N_8763,N_8539);
and U9051 (N_9051,N_8961,N_8473);
nor U9052 (N_9052,N_8417,N_8493);
and U9053 (N_9053,N_8927,N_8384);
nor U9054 (N_9054,N_8544,N_8061);
nor U9055 (N_9055,N_8147,N_8745);
nand U9056 (N_9056,N_8733,N_8123);
nor U9057 (N_9057,N_8832,N_8489);
and U9058 (N_9058,N_8971,N_8348);
or U9059 (N_9059,N_8443,N_8802);
nor U9060 (N_9060,N_8070,N_8677);
nand U9061 (N_9061,N_8500,N_8739);
or U9062 (N_9062,N_8749,N_8271);
nand U9063 (N_9063,N_8603,N_8000);
nand U9064 (N_9064,N_8688,N_8482);
or U9065 (N_9065,N_8477,N_8900);
nand U9066 (N_9066,N_8987,N_8050);
and U9067 (N_9067,N_8868,N_8115);
or U9068 (N_9068,N_8082,N_8494);
nor U9069 (N_9069,N_8842,N_8227);
xnor U9070 (N_9070,N_8766,N_8783);
nor U9071 (N_9071,N_8021,N_8444);
nor U9072 (N_9072,N_8328,N_8457);
and U9073 (N_9073,N_8447,N_8413);
nor U9074 (N_9074,N_8977,N_8923);
and U9075 (N_9075,N_8156,N_8794);
nor U9076 (N_9076,N_8057,N_8967);
nand U9077 (N_9077,N_8086,N_8501);
or U9078 (N_9078,N_8138,N_8940);
or U9079 (N_9079,N_8966,N_8510);
or U9080 (N_9080,N_8356,N_8699);
nand U9081 (N_9081,N_8642,N_8306);
nand U9082 (N_9082,N_8719,N_8450);
nand U9083 (N_9083,N_8598,N_8174);
and U9084 (N_9084,N_8935,N_8828);
nand U9085 (N_9085,N_8914,N_8392);
nor U9086 (N_9086,N_8552,N_8952);
nand U9087 (N_9087,N_8010,N_8612);
or U9088 (N_9088,N_8031,N_8527);
nand U9089 (N_9089,N_8625,N_8664);
or U9090 (N_9090,N_8622,N_8407);
nor U9091 (N_9091,N_8058,N_8459);
nand U9092 (N_9092,N_8327,N_8155);
nand U9093 (N_9093,N_8452,N_8132);
or U9094 (N_9094,N_8377,N_8665);
nand U9095 (N_9095,N_8303,N_8819);
and U9096 (N_9096,N_8591,N_8706);
or U9097 (N_9097,N_8352,N_8040);
nand U9098 (N_9098,N_8777,N_8666);
nor U9099 (N_9099,N_8781,N_8461);
nand U9100 (N_9100,N_8462,N_8852);
nor U9101 (N_9101,N_8797,N_8566);
or U9102 (N_9102,N_8605,N_8752);
and U9103 (N_9103,N_8083,N_8879);
nand U9104 (N_9104,N_8571,N_8279);
nor U9105 (N_9105,N_8003,N_8519);
and U9106 (N_9106,N_8583,N_8806);
or U9107 (N_9107,N_8560,N_8169);
nor U9108 (N_9108,N_8901,N_8820);
and U9109 (N_9109,N_8761,N_8518);
and U9110 (N_9110,N_8988,N_8793);
or U9111 (N_9111,N_8895,N_8460);
nor U9112 (N_9112,N_8782,N_8513);
or U9113 (N_9113,N_8830,N_8385);
or U9114 (N_9114,N_8320,N_8499);
or U9115 (N_9115,N_8107,N_8886);
nand U9116 (N_9116,N_8144,N_8696);
or U9117 (N_9117,N_8008,N_8231);
or U9118 (N_9118,N_8390,N_8244);
nor U9119 (N_9119,N_8873,N_8818);
or U9120 (N_9120,N_8836,N_8710);
and U9121 (N_9121,N_8840,N_8643);
and U9122 (N_9122,N_8222,N_8241);
and U9123 (N_9123,N_8958,N_8649);
nor U9124 (N_9124,N_8627,N_8545);
nand U9125 (N_9125,N_8234,N_8281);
nor U9126 (N_9126,N_8375,N_8564);
nand U9127 (N_9127,N_8861,N_8338);
and U9128 (N_9128,N_8788,N_8592);
and U9129 (N_9129,N_8981,N_8711);
nand U9130 (N_9130,N_8307,N_8403);
nand U9131 (N_9131,N_8073,N_8296);
nand U9132 (N_9132,N_8379,N_8396);
nand U9133 (N_9133,N_8308,N_8738);
nor U9134 (N_9134,N_8680,N_8673);
or U9135 (N_9135,N_8476,N_8055);
and U9136 (N_9136,N_8286,N_8573);
nor U9137 (N_9137,N_8162,N_8043);
or U9138 (N_9138,N_8607,N_8599);
or U9139 (N_9139,N_8790,N_8218);
nor U9140 (N_9140,N_8148,N_8672);
or U9141 (N_9141,N_8874,N_8951);
nor U9142 (N_9142,N_8743,N_8233);
and U9143 (N_9143,N_8361,N_8863);
and U9144 (N_9144,N_8065,N_8116);
or U9145 (N_9145,N_8650,N_8969);
and U9146 (N_9146,N_8041,N_8324);
or U9147 (N_9147,N_8330,N_8270);
nor U9148 (N_9148,N_8433,N_8776);
nand U9149 (N_9149,N_8930,N_8919);
and U9150 (N_9150,N_8465,N_8645);
nor U9151 (N_9151,N_8154,N_8345);
and U9152 (N_9152,N_8454,N_8026);
and U9153 (N_9153,N_8124,N_8554);
nor U9154 (N_9154,N_8446,N_8813);
nor U9155 (N_9155,N_8674,N_8942);
and U9156 (N_9156,N_8758,N_8805);
nand U9157 (N_9157,N_8770,N_8986);
or U9158 (N_9158,N_8093,N_8617);
nand U9159 (N_9159,N_8678,N_8437);
or U9160 (N_9160,N_8533,N_8689);
and U9161 (N_9161,N_8335,N_8284);
and U9162 (N_9162,N_8005,N_8736);
or U9163 (N_9163,N_8588,N_8737);
and U9164 (N_9164,N_8079,N_8735);
nand U9165 (N_9165,N_8621,N_8099);
nor U9166 (N_9166,N_8648,N_8215);
nand U9167 (N_9167,N_8239,N_8810);
nor U9168 (N_9168,N_8311,N_8855);
nor U9169 (N_9169,N_8287,N_8230);
or U9170 (N_9170,N_8329,N_8159);
nor U9171 (N_9171,N_8053,N_8804);
and U9172 (N_9172,N_8251,N_8341);
or U9173 (N_9173,N_8644,N_8857);
or U9174 (N_9174,N_8530,N_8634);
and U9175 (N_9175,N_8695,N_8506);
nor U9176 (N_9176,N_8889,N_8631);
nor U9177 (N_9177,N_8498,N_8449);
and U9178 (N_9178,N_8725,N_8532);
nor U9179 (N_9179,N_8027,N_8484);
nand U9180 (N_9180,N_8751,N_8979);
or U9181 (N_9181,N_8398,N_8859);
or U9182 (N_9182,N_8421,N_8298);
nand U9183 (N_9183,N_8636,N_8193);
nor U9184 (N_9184,N_8798,N_8980);
nor U9185 (N_9185,N_8724,N_8686);
nand U9186 (N_9186,N_8829,N_8884);
and U9187 (N_9187,N_8168,N_8915);
nor U9188 (N_9188,N_8389,N_8997);
nand U9189 (N_9189,N_8321,N_8372);
and U9190 (N_9190,N_8119,N_8887);
or U9191 (N_9191,N_8512,N_8871);
nand U9192 (N_9192,N_8274,N_8205);
nor U9193 (N_9193,N_8833,N_8956);
nand U9194 (N_9194,N_8718,N_8618);
and U9195 (N_9195,N_8595,N_8750);
nand U9196 (N_9196,N_8206,N_8197);
and U9197 (N_9197,N_8475,N_8020);
nor U9198 (N_9198,N_8240,N_8424);
nor U9199 (N_9199,N_8198,N_8196);
and U9200 (N_9200,N_8838,N_8470);
and U9201 (N_9201,N_8312,N_8567);
and U9202 (N_9202,N_8265,N_8704);
nor U9203 (N_9203,N_8092,N_8368);
or U9204 (N_9204,N_8326,N_8960);
and U9205 (N_9205,N_8078,N_8019);
nand U9206 (N_9206,N_8393,N_8100);
nand U9207 (N_9207,N_8276,N_8141);
or U9208 (N_9208,N_8604,N_8917);
and U9209 (N_9209,N_8847,N_8468);
or U9210 (N_9210,N_8984,N_8902);
and U9211 (N_9211,N_8563,N_8867);
or U9212 (N_9212,N_8671,N_8232);
nor U9213 (N_9213,N_8024,N_8496);
nand U9214 (N_9214,N_8382,N_8486);
nor U9215 (N_9215,N_8294,N_8690);
nand U9216 (N_9216,N_8740,N_8022);
and U9217 (N_9217,N_8295,N_8408);
nand U9218 (N_9218,N_8623,N_8151);
or U9219 (N_9219,N_8072,N_8620);
or U9220 (N_9220,N_8955,N_8562);
or U9221 (N_9221,N_8485,N_8635);
nor U9222 (N_9222,N_8697,N_8035);
or U9223 (N_9223,N_8692,N_8362);
or U9224 (N_9224,N_8028,N_8225);
or U9225 (N_9225,N_8355,N_8597);
nor U9226 (N_9226,N_8004,N_8226);
or U9227 (N_9227,N_8601,N_8074);
nor U9228 (N_9228,N_8609,N_8953);
and U9229 (N_9229,N_8202,N_8681);
and U9230 (N_9230,N_8419,N_8784);
or U9231 (N_9231,N_8358,N_8380);
and U9232 (N_9232,N_8237,N_8432);
or U9233 (N_9233,N_8976,N_8557);
or U9234 (N_9234,N_8464,N_8153);
nor U9235 (N_9235,N_8025,N_8931);
and U9236 (N_9236,N_8655,N_8897);
nand U9237 (N_9237,N_8872,N_8219);
nor U9238 (N_9238,N_8325,N_8280);
and U9239 (N_9239,N_8939,N_8186);
nor U9240 (N_9240,N_8120,N_8047);
nor U9241 (N_9241,N_8723,N_8062);
nor U9242 (N_9242,N_8442,N_8579);
nor U9243 (N_9243,N_8933,N_8007);
nand U9244 (N_9244,N_8929,N_8762);
or U9245 (N_9245,N_8164,N_8023);
or U9246 (N_9246,N_8509,N_8626);
or U9247 (N_9247,N_8416,N_8791);
and U9248 (N_9248,N_8542,N_8189);
or U9249 (N_9249,N_8789,N_8012);
nor U9250 (N_9250,N_8337,N_8679);
nand U9251 (N_9251,N_8823,N_8516);
nand U9252 (N_9252,N_8570,N_8364);
or U9253 (N_9253,N_8016,N_8131);
nor U9254 (N_9254,N_8880,N_8126);
and U9255 (N_9255,N_8463,N_8925);
nor U9256 (N_9256,N_8252,N_8180);
or U9257 (N_9257,N_8551,N_8077);
and U9258 (N_9258,N_8466,N_8962);
and U9259 (N_9259,N_8524,N_8676);
nor U9260 (N_9260,N_8729,N_8223);
nand U9261 (N_9261,N_8435,N_8285);
nand U9262 (N_9262,N_8816,N_8118);
and U9263 (N_9263,N_8869,N_8068);
nor U9264 (N_9264,N_8970,N_8268);
and U9265 (N_9265,N_8896,N_8322);
nand U9266 (N_9266,N_8965,N_8034);
xnor U9267 (N_9267,N_8508,N_8378);
and U9268 (N_9268,N_8038,N_8985);
nor U9269 (N_9269,N_8406,N_8550);
nor U9270 (N_9270,N_8204,N_8728);
nand U9271 (N_9271,N_8095,N_8870);
or U9272 (N_9272,N_8576,N_8780);
and U9273 (N_9273,N_8032,N_8742);
nor U9274 (N_9274,N_8292,N_8716);
and U9275 (N_9275,N_8343,N_8973);
nand U9276 (N_9276,N_8060,N_8608);
or U9277 (N_9277,N_8891,N_8754);
nand U9278 (N_9278,N_8959,N_8339);
nor U9279 (N_9279,N_8548,N_8905);
or U9280 (N_9280,N_8975,N_8972);
nor U9281 (N_9281,N_8538,N_8654);
nand U9282 (N_9282,N_8584,N_8366);
nand U9283 (N_9283,N_8507,N_8085);
or U9284 (N_9284,N_8236,N_8075);
nor U9285 (N_9285,N_8616,N_8229);
nor U9286 (N_9286,N_8192,N_8090);
and U9287 (N_9287,N_8748,N_8316);
and U9288 (N_9288,N_8849,N_8698);
nand U9289 (N_9289,N_8715,N_8850);
and U9290 (N_9290,N_8300,N_8888);
and U9291 (N_9291,N_8323,N_8129);
or U9292 (N_9292,N_8224,N_8210);
or U9293 (N_9293,N_8349,N_8821);
nand U9294 (N_9294,N_8675,N_8668);
and U9295 (N_9295,N_8827,N_8898);
or U9296 (N_9296,N_8950,N_8883);
nor U9297 (N_9297,N_8949,N_8195);
nand U9298 (N_9298,N_8253,N_8633);
nand U9299 (N_9299,N_8394,N_8152);
and U9300 (N_9300,N_8054,N_8937);
and U9301 (N_9301,N_8614,N_8864);
and U9302 (N_9302,N_8289,N_8685);
nor U9303 (N_9303,N_8974,N_8255);
nand U9304 (N_9304,N_8381,N_8628);
or U9305 (N_9305,N_8438,N_8596);
or U9306 (N_9306,N_8150,N_8048);
or U9307 (N_9307,N_8190,N_8491);
nor U9308 (N_9308,N_8213,N_8314);
nand U9309 (N_9309,N_8122,N_8418);
or U9310 (N_9310,N_8453,N_8243);
or U9311 (N_9311,N_8051,N_8275);
nand U9312 (N_9312,N_8831,N_8278);
nor U9313 (N_9313,N_8824,N_8167);
and U9314 (N_9314,N_8117,N_8893);
and U9315 (N_9315,N_8656,N_8342);
or U9316 (N_9316,N_8904,N_8002);
and U9317 (N_9317,N_8703,N_8044);
xor U9318 (N_9318,N_8064,N_8257);
and U9319 (N_9319,N_8456,N_8921);
xnor U9320 (N_9320,N_8787,N_8701);
nor U9321 (N_9321,N_8683,N_8405);
nand U9322 (N_9322,N_8522,N_8978);
nand U9323 (N_9323,N_8918,N_8448);
and U9324 (N_9324,N_8606,N_8926);
and U9325 (N_9325,N_8684,N_8344);
nand U9326 (N_9326,N_8360,N_8694);
or U9327 (N_9327,N_8815,N_8753);
or U9328 (N_9328,N_8511,N_8067);
and U9329 (N_9329,N_8478,N_8574);
nand U9330 (N_9330,N_8160,N_8890);
nand U9331 (N_9331,N_8247,N_8238);
nand U9332 (N_9332,N_8333,N_8017);
and U9333 (N_9333,N_8964,N_8908);
nor U9334 (N_9334,N_8097,N_8401);
nand U9335 (N_9335,N_8799,N_8488);
nor U9336 (N_9336,N_8658,N_8221);
nand U9337 (N_9337,N_8938,N_8288);
or U9338 (N_9338,N_8702,N_8811);
and U9339 (N_9339,N_8246,N_8877);
nor U9340 (N_9340,N_8261,N_8647);
or U9341 (N_9341,N_8367,N_8540);
or U9342 (N_9342,N_8096,N_8841);
and U9343 (N_9343,N_8580,N_8146);
and U9344 (N_9344,N_8371,N_8036);
nor U9345 (N_9345,N_8088,N_8529);
and U9346 (N_9346,N_8309,N_8480);
nor U9347 (N_9347,N_8319,N_8305);
nor U9348 (N_9348,N_8304,N_8549);
nor U9349 (N_9349,N_8528,N_8659);
or U9350 (N_9350,N_8217,N_8332);
or U9351 (N_9351,N_8001,N_8862);
or U9352 (N_9352,N_8553,N_8011);
nor U9353 (N_9353,N_8374,N_8881);
nor U9354 (N_9354,N_8839,N_8657);
and U9355 (N_9355,N_8142,N_8114);
nand U9356 (N_9356,N_8611,N_8809);
nand U9357 (N_9357,N_8602,N_8313);
and U9358 (N_9358,N_8803,N_8451);
or U9359 (N_9359,N_8479,N_8646);
nand U9360 (N_9360,N_8272,N_8504);
nand U9361 (N_9361,N_8860,N_8726);
and U9362 (N_9362,N_8290,N_8854);
and U9363 (N_9363,N_8845,N_8081);
nor U9364 (N_9364,N_8029,N_8235);
and U9365 (N_9365,N_8610,N_8188);
nand U9366 (N_9366,N_8211,N_8593);
and U9367 (N_9367,N_8347,N_8187);
or U9368 (N_9368,N_8558,N_8517);
or U9369 (N_9369,N_8892,N_8128);
nand U9370 (N_9370,N_8922,N_8826);
nor U9371 (N_9371,N_8181,N_8334);
and U9372 (N_9372,N_8410,N_8045);
and U9373 (N_9373,N_8291,N_8640);
and U9374 (N_9374,N_8134,N_8543);
nand U9375 (N_9375,N_8911,N_8910);
nand U9376 (N_9376,N_8759,N_8876);
nand U9377 (N_9377,N_8411,N_8732);
nor U9378 (N_9378,N_8731,N_8523);
nand U9379 (N_9379,N_8525,N_8481);
or U9380 (N_9380,N_8121,N_8066);
or U9381 (N_9381,N_8982,N_8248);
and U9382 (N_9382,N_8559,N_8541);
or U9383 (N_9383,N_8767,N_8346);
nor U9384 (N_9384,N_8844,N_8989);
and U9385 (N_9385,N_8993,N_8531);
and U9386 (N_9386,N_8894,N_8561);
nor U9387 (N_9387,N_8906,N_8037);
or U9388 (N_9388,N_8515,N_8365);
or U9389 (N_9389,N_8353,N_8670);
or U9390 (N_9390,N_8865,N_8166);
nand U9391 (N_9391,N_8946,N_8590);
or U9392 (N_9392,N_8775,N_8555);
and U9393 (N_9393,N_8402,N_8577);
nand U9394 (N_9394,N_8713,N_8882);
or U9395 (N_9395,N_8089,N_8277);
or U9396 (N_9396,N_8429,N_8885);
xor U9397 (N_9397,N_8662,N_8928);
and U9398 (N_9398,N_8125,N_8568);
nand U9399 (N_9399,N_8030,N_8630);
nor U9400 (N_9400,N_8471,N_8199);
and U9401 (N_9401,N_8547,N_8983);
and U9402 (N_9402,N_8042,N_8059);
and U9403 (N_9403,N_8727,N_8163);
nor U9404 (N_9404,N_8254,N_8943);
nand U9405 (N_9405,N_8357,N_8354);
nor U9406 (N_9406,N_8145,N_8483);
and U9407 (N_9407,N_8469,N_8179);
nor U9408 (N_9408,N_8376,N_8383);
nand U9409 (N_9409,N_8999,N_8817);
nand U9410 (N_9410,N_8741,N_8203);
nor U9411 (N_9411,N_8069,N_8404);
and U9412 (N_9412,N_8814,N_8422);
nor U9413 (N_9413,N_8600,N_8932);
nand U9414 (N_9414,N_8687,N_8439);
nand U9415 (N_9415,N_8260,N_8638);
nand U9416 (N_9416,N_8242,N_8534);
nand U9417 (N_9417,N_8575,N_8585);
nand U9418 (N_9418,N_8536,N_8521);
and U9419 (N_9419,N_8409,N_8400);
nor U9420 (N_9420,N_8968,N_8094);
nor U9421 (N_9421,N_8267,N_8415);
nand U9422 (N_9422,N_8774,N_8015);
nor U9423 (N_9423,N_8395,N_8178);
or U9424 (N_9424,N_8660,N_8995);
and U9425 (N_9425,N_8228,N_8105);
nor U9426 (N_9426,N_8013,N_8800);
and U9427 (N_9427,N_8214,N_8503);
or U9428 (N_9428,N_8112,N_8578);
and U9429 (N_9429,N_8269,N_8661);
nor U9430 (N_9430,N_8273,N_8594);
or U9431 (N_9431,N_8912,N_8565);
nor U9432 (N_9432,N_8848,N_8846);
nand U9433 (N_9433,N_8445,N_8639);
and U9434 (N_9434,N_8336,N_8194);
and U9435 (N_9435,N_8143,N_8109);
or U9436 (N_9436,N_8772,N_8712);
nand U9437 (N_9437,N_8667,N_8359);
nand U9438 (N_9438,N_8948,N_8208);
nand U9439 (N_9439,N_8370,N_8207);
nor U9440 (N_9440,N_8924,N_8520);
and U9441 (N_9441,N_8200,N_8866);
or U9442 (N_9442,N_8708,N_8916);
or U9443 (N_9443,N_8185,N_8764);
nor U9444 (N_9444,N_8299,N_8103);
nor U9445 (N_9445,N_8572,N_8569);
or U9446 (N_9446,N_8216,N_8834);
or U9447 (N_9447,N_8391,N_8589);
or U9448 (N_9448,N_8653,N_8792);
and U9449 (N_9449,N_8106,N_8049);
and U9450 (N_9450,N_8425,N_8420);
nand U9451 (N_9451,N_8822,N_8747);
and U9452 (N_9452,N_8556,N_8388);
nor U9453 (N_9453,N_8363,N_8245);
or U9454 (N_9454,N_8177,N_8184);
nor U9455 (N_9455,N_8046,N_8250);
nor U9456 (N_9456,N_8587,N_8957);
nand U9457 (N_9457,N_8705,N_8014);
nor U9458 (N_9458,N_8104,N_8526);
nor U9459 (N_9459,N_8140,N_8310);
nand U9460 (N_9460,N_8111,N_8175);
and U9461 (N_9461,N_8033,N_8795);
nor U9462 (N_9462,N_8652,N_8613);
or U9463 (N_9463,N_8615,N_8582);
nor U9464 (N_9464,N_8136,N_8913);
or U9465 (N_9465,N_8006,N_8331);
or U9466 (N_9466,N_8546,N_8266);
nand U9467 (N_9467,N_8756,N_8259);
nand U9468 (N_9468,N_8467,N_8936);
nand U9469 (N_9469,N_8669,N_8858);
nand U9470 (N_9470,N_8428,N_8765);
and U9471 (N_9471,N_8350,N_8137);
and U9472 (N_9472,N_8786,N_8709);
nor U9473 (N_9473,N_8934,N_8771);
nand U9474 (N_9474,N_8427,N_8778);
and U9475 (N_9475,N_8212,N_8637);
nand U9476 (N_9476,N_8619,N_8651);
nand U9477 (N_9477,N_8757,N_8825);
nor U9478 (N_9478,N_8856,N_8108);
nand U9479 (N_9479,N_8101,N_8436);
and U9480 (N_9480,N_8994,N_8487);
and U9481 (N_9481,N_8760,N_8586);
nor U9482 (N_9482,N_8941,N_8730);
and U9483 (N_9483,N_8707,N_8853);
nor U9484 (N_9484,N_8256,N_8455);
and U9485 (N_9485,N_8773,N_8843);
or U9486 (N_9486,N_8039,N_8779);
or U9487 (N_9487,N_8785,N_8098);
nor U9488 (N_9488,N_8629,N_8502);
and U9489 (N_9489,N_8722,N_8440);
and U9490 (N_9490,N_8641,N_8258);
nand U9491 (N_9491,N_8495,N_8158);
nand U9492 (N_9492,N_8426,N_8920);
or U9493 (N_9493,N_8581,N_8283);
and U9494 (N_9494,N_8963,N_8423);
or U9495 (N_9495,N_8663,N_8018);
and U9496 (N_9496,N_8945,N_8183);
or U9497 (N_9497,N_8717,N_8441);
nand U9498 (N_9498,N_8102,N_8909);
and U9499 (N_9499,N_8624,N_8149);
and U9500 (N_9500,N_8290,N_8995);
or U9501 (N_9501,N_8562,N_8338);
and U9502 (N_9502,N_8086,N_8967);
nor U9503 (N_9503,N_8814,N_8817);
or U9504 (N_9504,N_8369,N_8964);
nor U9505 (N_9505,N_8828,N_8659);
and U9506 (N_9506,N_8559,N_8098);
nor U9507 (N_9507,N_8561,N_8139);
nor U9508 (N_9508,N_8215,N_8758);
or U9509 (N_9509,N_8844,N_8087);
nor U9510 (N_9510,N_8836,N_8504);
nand U9511 (N_9511,N_8356,N_8919);
nor U9512 (N_9512,N_8097,N_8719);
nor U9513 (N_9513,N_8892,N_8921);
and U9514 (N_9514,N_8197,N_8275);
nand U9515 (N_9515,N_8817,N_8813);
nand U9516 (N_9516,N_8558,N_8552);
or U9517 (N_9517,N_8405,N_8432);
nor U9518 (N_9518,N_8485,N_8331);
and U9519 (N_9519,N_8432,N_8353);
nor U9520 (N_9520,N_8628,N_8920);
nor U9521 (N_9521,N_8996,N_8090);
nand U9522 (N_9522,N_8044,N_8181);
or U9523 (N_9523,N_8797,N_8497);
and U9524 (N_9524,N_8629,N_8171);
and U9525 (N_9525,N_8416,N_8947);
nand U9526 (N_9526,N_8325,N_8095);
and U9527 (N_9527,N_8276,N_8202);
and U9528 (N_9528,N_8193,N_8603);
nor U9529 (N_9529,N_8446,N_8820);
or U9530 (N_9530,N_8865,N_8016);
nor U9531 (N_9531,N_8609,N_8826);
nor U9532 (N_9532,N_8302,N_8855);
nand U9533 (N_9533,N_8491,N_8184);
nand U9534 (N_9534,N_8154,N_8954);
nand U9535 (N_9535,N_8640,N_8431);
or U9536 (N_9536,N_8638,N_8603);
and U9537 (N_9537,N_8914,N_8089);
or U9538 (N_9538,N_8188,N_8220);
and U9539 (N_9539,N_8075,N_8004);
nand U9540 (N_9540,N_8730,N_8686);
nor U9541 (N_9541,N_8633,N_8115);
and U9542 (N_9542,N_8409,N_8307);
or U9543 (N_9543,N_8062,N_8661);
and U9544 (N_9544,N_8909,N_8008);
nand U9545 (N_9545,N_8456,N_8592);
and U9546 (N_9546,N_8113,N_8745);
nor U9547 (N_9547,N_8344,N_8752);
xnor U9548 (N_9548,N_8365,N_8632);
nor U9549 (N_9549,N_8045,N_8480);
nand U9550 (N_9550,N_8690,N_8092);
nand U9551 (N_9551,N_8342,N_8685);
nor U9552 (N_9552,N_8832,N_8889);
nor U9553 (N_9553,N_8388,N_8238);
nor U9554 (N_9554,N_8958,N_8708);
nand U9555 (N_9555,N_8557,N_8660);
or U9556 (N_9556,N_8143,N_8423);
nor U9557 (N_9557,N_8334,N_8792);
nor U9558 (N_9558,N_8580,N_8093);
nor U9559 (N_9559,N_8221,N_8829);
nor U9560 (N_9560,N_8321,N_8145);
nand U9561 (N_9561,N_8712,N_8100);
and U9562 (N_9562,N_8362,N_8858);
or U9563 (N_9563,N_8617,N_8745);
and U9564 (N_9564,N_8326,N_8468);
nand U9565 (N_9565,N_8927,N_8359);
and U9566 (N_9566,N_8727,N_8473);
or U9567 (N_9567,N_8845,N_8669);
and U9568 (N_9568,N_8405,N_8610);
or U9569 (N_9569,N_8721,N_8134);
nor U9570 (N_9570,N_8366,N_8447);
and U9571 (N_9571,N_8107,N_8606);
or U9572 (N_9572,N_8731,N_8741);
and U9573 (N_9573,N_8119,N_8923);
or U9574 (N_9574,N_8269,N_8237);
and U9575 (N_9575,N_8748,N_8524);
nand U9576 (N_9576,N_8507,N_8637);
and U9577 (N_9577,N_8907,N_8716);
nand U9578 (N_9578,N_8931,N_8108);
nand U9579 (N_9579,N_8418,N_8669);
nand U9580 (N_9580,N_8791,N_8458);
nand U9581 (N_9581,N_8988,N_8975);
or U9582 (N_9582,N_8199,N_8281);
and U9583 (N_9583,N_8698,N_8267);
nand U9584 (N_9584,N_8793,N_8476);
nor U9585 (N_9585,N_8094,N_8340);
or U9586 (N_9586,N_8974,N_8790);
nor U9587 (N_9587,N_8178,N_8762);
or U9588 (N_9588,N_8709,N_8862);
or U9589 (N_9589,N_8683,N_8973);
and U9590 (N_9590,N_8889,N_8732);
or U9591 (N_9591,N_8061,N_8955);
and U9592 (N_9592,N_8854,N_8230);
nand U9593 (N_9593,N_8161,N_8047);
or U9594 (N_9594,N_8082,N_8191);
or U9595 (N_9595,N_8612,N_8086);
and U9596 (N_9596,N_8435,N_8524);
nand U9597 (N_9597,N_8669,N_8833);
or U9598 (N_9598,N_8441,N_8785);
nor U9599 (N_9599,N_8101,N_8633);
nand U9600 (N_9600,N_8441,N_8430);
nand U9601 (N_9601,N_8904,N_8814);
nor U9602 (N_9602,N_8782,N_8043);
or U9603 (N_9603,N_8944,N_8662);
nand U9604 (N_9604,N_8327,N_8676);
nor U9605 (N_9605,N_8249,N_8168);
and U9606 (N_9606,N_8586,N_8968);
nand U9607 (N_9607,N_8055,N_8266);
or U9608 (N_9608,N_8667,N_8961);
nor U9609 (N_9609,N_8221,N_8990);
nand U9610 (N_9610,N_8295,N_8587);
or U9611 (N_9611,N_8962,N_8793);
nand U9612 (N_9612,N_8873,N_8524);
nand U9613 (N_9613,N_8671,N_8884);
or U9614 (N_9614,N_8711,N_8156);
or U9615 (N_9615,N_8512,N_8698);
and U9616 (N_9616,N_8848,N_8724);
nor U9617 (N_9617,N_8187,N_8998);
nand U9618 (N_9618,N_8220,N_8793);
nand U9619 (N_9619,N_8173,N_8097);
and U9620 (N_9620,N_8908,N_8578);
or U9621 (N_9621,N_8299,N_8423);
nand U9622 (N_9622,N_8884,N_8454);
and U9623 (N_9623,N_8829,N_8704);
and U9624 (N_9624,N_8105,N_8143);
and U9625 (N_9625,N_8731,N_8961);
or U9626 (N_9626,N_8849,N_8859);
nand U9627 (N_9627,N_8533,N_8628);
or U9628 (N_9628,N_8749,N_8991);
nand U9629 (N_9629,N_8531,N_8486);
nor U9630 (N_9630,N_8443,N_8311);
or U9631 (N_9631,N_8504,N_8298);
or U9632 (N_9632,N_8982,N_8349);
or U9633 (N_9633,N_8163,N_8667);
nand U9634 (N_9634,N_8662,N_8645);
nand U9635 (N_9635,N_8390,N_8906);
and U9636 (N_9636,N_8543,N_8923);
nand U9637 (N_9637,N_8423,N_8111);
nor U9638 (N_9638,N_8077,N_8457);
or U9639 (N_9639,N_8923,N_8597);
or U9640 (N_9640,N_8669,N_8873);
or U9641 (N_9641,N_8338,N_8748);
or U9642 (N_9642,N_8805,N_8423);
nor U9643 (N_9643,N_8591,N_8577);
nand U9644 (N_9644,N_8745,N_8069);
nand U9645 (N_9645,N_8454,N_8070);
or U9646 (N_9646,N_8499,N_8483);
nand U9647 (N_9647,N_8119,N_8500);
nor U9648 (N_9648,N_8267,N_8451);
nand U9649 (N_9649,N_8910,N_8333);
and U9650 (N_9650,N_8485,N_8708);
nand U9651 (N_9651,N_8374,N_8148);
and U9652 (N_9652,N_8669,N_8583);
nor U9653 (N_9653,N_8921,N_8631);
and U9654 (N_9654,N_8336,N_8214);
and U9655 (N_9655,N_8694,N_8171);
and U9656 (N_9656,N_8923,N_8208);
nand U9657 (N_9657,N_8125,N_8165);
nor U9658 (N_9658,N_8439,N_8609);
nor U9659 (N_9659,N_8268,N_8776);
or U9660 (N_9660,N_8759,N_8160);
xor U9661 (N_9661,N_8060,N_8188);
and U9662 (N_9662,N_8412,N_8551);
nand U9663 (N_9663,N_8451,N_8566);
nand U9664 (N_9664,N_8274,N_8529);
nor U9665 (N_9665,N_8872,N_8724);
or U9666 (N_9666,N_8395,N_8127);
nand U9667 (N_9667,N_8994,N_8222);
xnor U9668 (N_9668,N_8205,N_8947);
nor U9669 (N_9669,N_8367,N_8014);
and U9670 (N_9670,N_8478,N_8460);
nor U9671 (N_9671,N_8492,N_8247);
or U9672 (N_9672,N_8251,N_8410);
and U9673 (N_9673,N_8856,N_8004);
and U9674 (N_9674,N_8047,N_8637);
nand U9675 (N_9675,N_8282,N_8380);
nor U9676 (N_9676,N_8673,N_8487);
nand U9677 (N_9677,N_8505,N_8976);
or U9678 (N_9678,N_8081,N_8272);
nand U9679 (N_9679,N_8845,N_8192);
or U9680 (N_9680,N_8900,N_8971);
nor U9681 (N_9681,N_8763,N_8266);
and U9682 (N_9682,N_8082,N_8305);
or U9683 (N_9683,N_8157,N_8839);
xor U9684 (N_9684,N_8362,N_8720);
nand U9685 (N_9685,N_8404,N_8682);
nor U9686 (N_9686,N_8581,N_8437);
or U9687 (N_9687,N_8165,N_8049);
nand U9688 (N_9688,N_8786,N_8672);
and U9689 (N_9689,N_8307,N_8434);
nor U9690 (N_9690,N_8600,N_8755);
nand U9691 (N_9691,N_8794,N_8624);
and U9692 (N_9692,N_8079,N_8747);
nand U9693 (N_9693,N_8225,N_8953);
or U9694 (N_9694,N_8064,N_8946);
nand U9695 (N_9695,N_8295,N_8238);
nand U9696 (N_9696,N_8550,N_8427);
nand U9697 (N_9697,N_8358,N_8142);
xor U9698 (N_9698,N_8527,N_8999);
nor U9699 (N_9699,N_8501,N_8238);
and U9700 (N_9700,N_8963,N_8607);
or U9701 (N_9701,N_8121,N_8297);
or U9702 (N_9702,N_8855,N_8870);
nor U9703 (N_9703,N_8724,N_8679);
nand U9704 (N_9704,N_8034,N_8394);
nor U9705 (N_9705,N_8532,N_8673);
nor U9706 (N_9706,N_8021,N_8160);
nor U9707 (N_9707,N_8818,N_8216);
or U9708 (N_9708,N_8298,N_8803);
or U9709 (N_9709,N_8936,N_8901);
nand U9710 (N_9710,N_8339,N_8948);
or U9711 (N_9711,N_8701,N_8470);
nand U9712 (N_9712,N_8471,N_8711);
nor U9713 (N_9713,N_8533,N_8252);
and U9714 (N_9714,N_8476,N_8024);
nor U9715 (N_9715,N_8803,N_8820);
nor U9716 (N_9716,N_8838,N_8462);
nor U9717 (N_9717,N_8134,N_8749);
nand U9718 (N_9718,N_8786,N_8386);
and U9719 (N_9719,N_8729,N_8644);
and U9720 (N_9720,N_8268,N_8162);
and U9721 (N_9721,N_8991,N_8814);
nand U9722 (N_9722,N_8225,N_8809);
and U9723 (N_9723,N_8478,N_8971);
or U9724 (N_9724,N_8926,N_8528);
and U9725 (N_9725,N_8809,N_8776);
or U9726 (N_9726,N_8647,N_8070);
or U9727 (N_9727,N_8226,N_8076);
or U9728 (N_9728,N_8681,N_8256);
nand U9729 (N_9729,N_8481,N_8516);
nand U9730 (N_9730,N_8218,N_8722);
or U9731 (N_9731,N_8550,N_8057);
nor U9732 (N_9732,N_8029,N_8023);
nand U9733 (N_9733,N_8331,N_8885);
and U9734 (N_9734,N_8252,N_8525);
nor U9735 (N_9735,N_8787,N_8501);
and U9736 (N_9736,N_8491,N_8256);
and U9737 (N_9737,N_8371,N_8855);
nand U9738 (N_9738,N_8369,N_8703);
or U9739 (N_9739,N_8974,N_8085);
nor U9740 (N_9740,N_8494,N_8385);
and U9741 (N_9741,N_8888,N_8242);
or U9742 (N_9742,N_8233,N_8103);
nand U9743 (N_9743,N_8573,N_8311);
nand U9744 (N_9744,N_8425,N_8823);
nor U9745 (N_9745,N_8799,N_8393);
or U9746 (N_9746,N_8473,N_8795);
xor U9747 (N_9747,N_8426,N_8374);
or U9748 (N_9748,N_8110,N_8378);
and U9749 (N_9749,N_8797,N_8295);
nand U9750 (N_9750,N_8352,N_8444);
nand U9751 (N_9751,N_8296,N_8329);
nand U9752 (N_9752,N_8007,N_8564);
nor U9753 (N_9753,N_8645,N_8583);
and U9754 (N_9754,N_8911,N_8462);
and U9755 (N_9755,N_8444,N_8285);
and U9756 (N_9756,N_8686,N_8803);
and U9757 (N_9757,N_8140,N_8808);
or U9758 (N_9758,N_8697,N_8088);
nor U9759 (N_9759,N_8332,N_8696);
and U9760 (N_9760,N_8760,N_8585);
or U9761 (N_9761,N_8296,N_8224);
nand U9762 (N_9762,N_8907,N_8831);
and U9763 (N_9763,N_8009,N_8122);
or U9764 (N_9764,N_8771,N_8871);
and U9765 (N_9765,N_8622,N_8351);
nor U9766 (N_9766,N_8710,N_8419);
nand U9767 (N_9767,N_8757,N_8597);
and U9768 (N_9768,N_8078,N_8882);
nor U9769 (N_9769,N_8970,N_8537);
and U9770 (N_9770,N_8110,N_8099);
nand U9771 (N_9771,N_8198,N_8611);
and U9772 (N_9772,N_8987,N_8713);
or U9773 (N_9773,N_8070,N_8538);
nor U9774 (N_9774,N_8212,N_8449);
and U9775 (N_9775,N_8313,N_8607);
nand U9776 (N_9776,N_8629,N_8995);
nor U9777 (N_9777,N_8617,N_8180);
or U9778 (N_9778,N_8575,N_8406);
and U9779 (N_9779,N_8323,N_8506);
nor U9780 (N_9780,N_8610,N_8581);
nor U9781 (N_9781,N_8729,N_8929);
nand U9782 (N_9782,N_8096,N_8784);
nor U9783 (N_9783,N_8571,N_8604);
nand U9784 (N_9784,N_8969,N_8987);
nor U9785 (N_9785,N_8937,N_8501);
or U9786 (N_9786,N_8608,N_8936);
nand U9787 (N_9787,N_8164,N_8842);
and U9788 (N_9788,N_8508,N_8245);
or U9789 (N_9789,N_8372,N_8490);
nor U9790 (N_9790,N_8797,N_8342);
nand U9791 (N_9791,N_8868,N_8820);
or U9792 (N_9792,N_8715,N_8377);
nand U9793 (N_9793,N_8274,N_8136);
nor U9794 (N_9794,N_8313,N_8915);
and U9795 (N_9795,N_8033,N_8045);
nor U9796 (N_9796,N_8862,N_8386);
nand U9797 (N_9797,N_8133,N_8132);
nor U9798 (N_9798,N_8566,N_8243);
nand U9799 (N_9799,N_8671,N_8339);
and U9800 (N_9800,N_8775,N_8433);
nand U9801 (N_9801,N_8394,N_8554);
nor U9802 (N_9802,N_8115,N_8825);
nand U9803 (N_9803,N_8345,N_8421);
or U9804 (N_9804,N_8969,N_8826);
or U9805 (N_9805,N_8059,N_8965);
and U9806 (N_9806,N_8664,N_8018);
or U9807 (N_9807,N_8899,N_8879);
and U9808 (N_9808,N_8117,N_8871);
xnor U9809 (N_9809,N_8853,N_8290);
nor U9810 (N_9810,N_8090,N_8557);
or U9811 (N_9811,N_8278,N_8238);
and U9812 (N_9812,N_8199,N_8062);
or U9813 (N_9813,N_8625,N_8528);
nor U9814 (N_9814,N_8172,N_8505);
nand U9815 (N_9815,N_8614,N_8549);
and U9816 (N_9816,N_8248,N_8214);
and U9817 (N_9817,N_8550,N_8875);
or U9818 (N_9818,N_8659,N_8955);
nand U9819 (N_9819,N_8326,N_8373);
nor U9820 (N_9820,N_8696,N_8663);
nor U9821 (N_9821,N_8291,N_8148);
nand U9822 (N_9822,N_8019,N_8750);
and U9823 (N_9823,N_8720,N_8887);
nand U9824 (N_9824,N_8687,N_8749);
and U9825 (N_9825,N_8616,N_8907);
nor U9826 (N_9826,N_8646,N_8186);
or U9827 (N_9827,N_8244,N_8647);
nand U9828 (N_9828,N_8056,N_8104);
nand U9829 (N_9829,N_8559,N_8637);
nand U9830 (N_9830,N_8145,N_8669);
or U9831 (N_9831,N_8554,N_8884);
or U9832 (N_9832,N_8629,N_8873);
nand U9833 (N_9833,N_8236,N_8826);
nand U9834 (N_9834,N_8200,N_8075);
nand U9835 (N_9835,N_8941,N_8575);
nor U9836 (N_9836,N_8412,N_8260);
or U9837 (N_9837,N_8962,N_8436);
xor U9838 (N_9838,N_8387,N_8318);
nor U9839 (N_9839,N_8096,N_8974);
nand U9840 (N_9840,N_8621,N_8797);
or U9841 (N_9841,N_8823,N_8561);
and U9842 (N_9842,N_8518,N_8082);
xor U9843 (N_9843,N_8040,N_8174);
nor U9844 (N_9844,N_8259,N_8895);
and U9845 (N_9845,N_8571,N_8302);
and U9846 (N_9846,N_8170,N_8893);
nand U9847 (N_9847,N_8209,N_8395);
or U9848 (N_9848,N_8311,N_8738);
nand U9849 (N_9849,N_8524,N_8358);
and U9850 (N_9850,N_8881,N_8449);
or U9851 (N_9851,N_8731,N_8449);
and U9852 (N_9852,N_8539,N_8853);
nand U9853 (N_9853,N_8013,N_8600);
and U9854 (N_9854,N_8642,N_8919);
nand U9855 (N_9855,N_8847,N_8360);
nand U9856 (N_9856,N_8349,N_8233);
nand U9857 (N_9857,N_8581,N_8062);
or U9858 (N_9858,N_8991,N_8336);
and U9859 (N_9859,N_8597,N_8271);
nor U9860 (N_9860,N_8250,N_8001);
nand U9861 (N_9861,N_8916,N_8904);
and U9862 (N_9862,N_8737,N_8326);
nand U9863 (N_9863,N_8949,N_8703);
nor U9864 (N_9864,N_8392,N_8590);
nor U9865 (N_9865,N_8433,N_8254);
and U9866 (N_9866,N_8407,N_8073);
and U9867 (N_9867,N_8056,N_8619);
xor U9868 (N_9868,N_8753,N_8076);
and U9869 (N_9869,N_8476,N_8267);
or U9870 (N_9870,N_8335,N_8844);
and U9871 (N_9871,N_8799,N_8245);
or U9872 (N_9872,N_8173,N_8787);
nand U9873 (N_9873,N_8568,N_8522);
nor U9874 (N_9874,N_8739,N_8808);
nor U9875 (N_9875,N_8572,N_8481);
nor U9876 (N_9876,N_8339,N_8131);
nand U9877 (N_9877,N_8727,N_8064);
or U9878 (N_9878,N_8630,N_8206);
or U9879 (N_9879,N_8725,N_8250);
nor U9880 (N_9880,N_8807,N_8463);
nand U9881 (N_9881,N_8861,N_8692);
and U9882 (N_9882,N_8681,N_8741);
and U9883 (N_9883,N_8985,N_8722);
nor U9884 (N_9884,N_8358,N_8162);
or U9885 (N_9885,N_8683,N_8636);
or U9886 (N_9886,N_8166,N_8750);
or U9887 (N_9887,N_8848,N_8931);
nand U9888 (N_9888,N_8832,N_8497);
nand U9889 (N_9889,N_8200,N_8049);
nand U9890 (N_9890,N_8763,N_8481);
and U9891 (N_9891,N_8123,N_8048);
xnor U9892 (N_9892,N_8339,N_8082);
nor U9893 (N_9893,N_8325,N_8509);
nand U9894 (N_9894,N_8160,N_8361);
nor U9895 (N_9895,N_8561,N_8328);
or U9896 (N_9896,N_8466,N_8061);
nor U9897 (N_9897,N_8308,N_8486);
and U9898 (N_9898,N_8174,N_8747);
nand U9899 (N_9899,N_8319,N_8311);
nand U9900 (N_9900,N_8161,N_8810);
nand U9901 (N_9901,N_8424,N_8680);
and U9902 (N_9902,N_8608,N_8755);
nor U9903 (N_9903,N_8328,N_8450);
nand U9904 (N_9904,N_8223,N_8140);
and U9905 (N_9905,N_8660,N_8750);
nand U9906 (N_9906,N_8358,N_8237);
and U9907 (N_9907,N_8536,N_8177);
and U9908 (N_9908,N_8744,N_8486);
nor U9909 (N_9909,N_8490,N_8472);
nor U9910 (N_9910,N_8130,N_8528);
nor U9911 (N_9911,N_8604,N_8568);
nor U9912 (N_9912,N_8655,N_8612);
or U9913 (N_9913,N_8903,N_8852);
nor U9914 (N_9914,N_8114,N_8056);
nand U9915 (N_9915,N_8899,N_8873);
and U9916 (N_9916,N_8722,N_8652);
nand U9917 (N_9917,N_8556,N_8628);
nor U9918 (N_9918,N_8528,N_8459);
nor U9919 (N_9919,N_8613,N_8448);
nand U9920 (N_9920,N_8109,N_8314);
or U9921 (N_9921,N_8259,N_8253);
or U9922 (N_9922,N_8841,N_8362);
or U9923 (N_9923,N_8432,N_8265);
or U9924 (N_9924,N_8826,N_8258);
nor U9925 (N_9925,N_8176,N_8068);
or U9926 (N_9926,N_8931,N_8409);
or U9927 (N_9927,N_8327,N_8040);
and U9928 (N_9928,N_8730,N_8540);
or U9929 (N_9929,N_8188,N_8812);
and U9930 (N_9930,N_8053,N_8746);
or U9931 (N_9931,N_8296,N_8897);
nor U9932 (N_9932,N_8367,N_8672);
or U9933 (N_9933,N_8111,N_8967);
or U9934 (N_9934,N_8956,N_8973);
nand U9935 (N_9935,N_8662,N_8816);
or U9936 (N_9936,N_8794,N_8887);
nor U9937 (N_9937,N_8402,N_8868);
and U9938 (N_9938,N_8507,N_8021);
nand U9939 (N_9939,N_8808,N_8942);
or U9940 (N_9940,N_8384,N_8146);
nor U9941 (N_9941,N_8751,N_8184);
or U9942 (N_9942,N_8908,N_8936);
and U9943 (N_9943,N_8816,N_8639);
and U9944 (N_9944,N_8493,N_8598);
or U9945 (N_9945,N_8604,N_8539);
and U9946 (N_9946,N_8176,N_8241);
or U9947 (N_9947,N_8654,N_8501);
nand U9948 (N_9948,N_8905,N_8629);
or U9949 (N_9949,N_8408,N_8308);
nand U9950 (N_9950,N_8666,N_8210);
and U9951 (N_9951,N_8619,N_8266);
nor U9952 (N_9952,N_8767,N_8568);
or U9953 (N_9953,N_8036,N_8021);
nor U9954 (N_9954,N_8350,N_8607);
nand U9955 (N_9955,N_8374,N_8380);
and U9956 (N_9956,N_8036,N_8899);
and U9957 (N_9957,N_8367,N_8310);
nor U9958 (N_9958,N_8172,N_8953);
or U9959 (N_9959,N_8156,N_8365);
nor U9960 (N_9960,N_8382,N_8194);
or U9961 (N_9961,N_8457,N_8334);
nand U9962 (N_9962,N_8963,N_8013);
and U9963 (N_9963,N_8551,N_8358);
and U9964 (N_9964,N_8966,N_8315);
nor U9965 (N_9965,N_8781,N_8675);
nand U9966 (N_9966,N_8498,N_8679);
and U9967 (N_9967,N_8631,N_8164);
or U9968 (N_9968,N_8117,N_8341);
and U9969 (N_9969,N_8656,N_8496);
and U9970 (N_9970,N_8018,N_8084);
nand U9971 (N_9971,N_8141,N_8353);
nand U9972 (N_9972,N_8578,N_8789);
and U9973 (N_9973,N_8690,N_8696);
or U9974 (N_9974,N_8317,N_8414);
or U9975 (N_9975,N_8497,N_8900);
nor U9976 (N_9976,N_8801,N_8392);
nor U9977 (N_9977,N_8676,N_8857);
nand U9978 (N_9978,N_8252,N_8333);
nor U9979 (N_9979,N_8823,N_8782);
nor U9980 (N_9980,N_8616,N_8496);
nand U9981 (N_9981,N_8338,N_8093);
and U9982 (N_9982,N_8676,N_8691);
nor U9983 (N_9983,N_8722,N_8713);
or U9984 (N_9984,N_8602,N_8287);
and U9985 (N_9985,N_8064,N_8618);
or U9986 (N_9986,N_8867,N_8171);
nor U9987 (N_9987,N_8938,N_8210);
and U9988 (N_9988,N_8474,N_8804);
nand U9989 (N_9989,N_8818,N_8032);
and U9990 (N_9990,N_8955,N_8942);
nor U9991 (N_9991,N_8985,N_8524);
nor U9992 (N_9992,N_8016,N_8909);
and U9993 (N_9993,N_8734,N_8283);
and U9994 (N_9994,N_8261,N_8351);
or U9995 (N_9995,N_8991,N_8562);
and U9996 (N_9996,N_8193,N_8352);
nand U9997 (N_9997,N_8519,N_8110);
or U9998 (N_9998,N_8163,N_8881);
nand U9999 (N_9999,N_8621,N_8832);
or UO_0 (O_0,N_9538,N_9999);
or UO_1 (O_1,N_9054,N_9730);
nor UO_2 (O_2,N_9523,N_9807);
nor UO_3 (O_3,N_9699,N_9343);
or UO_4 (O_4,N_9536,N_9843);
and UO_5 (O_5,N_9308,N_9004);
and UO_6 (O_6,N_9342,N_9927);
nor UO_7 (O_7,N_9787,N_9026);
or UO_8 (O_8,N_9240,N_9478);
nor UO_9 (O_9,N_9090,N_9713);
nor UO_10 (O_10,N_9182,N_9610);
or UO_11 (O_11,N_9663,N_9047);
nand UO_12 (O_12,N_9042,N_9269);
and UO_13 (O_13,N_9388,N_9371);
or UO_14 (O_14,N_9684,N_9448);
nand UO_15 (O_15,N_9035,N_9970);
or UO_16 (O_16,N_9349,N_9802);
or UO_17 (O_17,N_9016,N_9548);
nand UO_18 (O_18,N_9301,N_9134);
nor UO_19 (O_19,N_9854,N_9592);
or UO_20 (O_20,N_9074,N_9630);
nor UO_21 (O_21,N_9245,N_9409);
or UO_22 (O_22,N_9763,N_9627);
or UO_23 (O_23,N_9121,N_9726);
nor UO_24 (O_24,N_9049,N_9119);
or UO_25 (O_25,N_9877,N_9836);
nand UO_26 (O_26,N_9268,N_9833);
and UO_27 (O_27,N_9552,N_9487);
and UO_28 (O_28,N_9594,N_9465);
nor UO_29 (O_29,N_9283,N_9602);
and UO_30 (O_30,N_9991,N_9468);
and UO_31 (O_31,N_9702,N_9230);
and UO_32 (O_32,N_9775,N_9011);
or UO_33 (O_33,N_9814,N_9431);
nand UO_34 (O_34,N_9876,N_9104);
nand UO_35 (O_35,N_9467,N_9980);
and UO_36 (O_36,N_9369,N_9483);
nor UO_37 (O_37,N_9660,N_9391);
and UO_38 (O_38,N_9373,N_9540);
nand UO_39 (O_39,N_9088,N_9709);
or UO_40 (O_40,N_9399,N_9239);
xor UO_41 (O_41,N_9312,N_9828);
nand UO_42 (O_42,N_9274,N_9733);
nor UO_43 (O_43,N_9822,N_9915);
or UO_44 (O_44,N_9194,N_9103);
and UO_45 (O_45,N_9385,N_9958);
or UO_46 (O_46,N_9493,N_9394);
and UO_47 (O_47,N_9585,N_9278);
or UO_48 (O_48,N_9938,N_9347);
and UO_49 (O_49,N_9811,N_9213);
and UO_50 (O_50,N_9866,N_9637);
or UO_51 (O_51,N_9514,N_9438);
or UO_52 (O_52,N_9595,N_9755);
nand UO_53 (O_53,N_9537,N_9508);
nor UO_54 (O_54,N_9719,N_9325);
and UO_55 (O_55,N_9341,N_9275);
and UO_56 (O_56,N_9251,N_9056);
or UO_57 (O_57,N_9234,N_9737);
nand UO_58 (O_58,N_9912,N_9148);
nand UO_59 (O_59,N_9307,N_9521);
nor UO_60 (O_60,N_9524,N_9174);
or UO_61 (O_61,N_9113,N_9625);
nand UO_62 (O_62,N_9293,N_9815);
or UO_63 (O_63,N_9977,N_9222);
and UO_64 (O_64,N_9582,N_9471);
nor UO_65 (O_65,N_9550,N_9058);
or UO_66 (O_66,N_9850,N_9348);
and UO_67 (O_67,N_9507,N_9855);
nand UO_68 (O_68,N_9377,N_9392);
nor UO_69 (O_69,N_9135,N_9241);
nand UO_70 (O_70,N_9800,N_9764);
or UO_71 (O_71,N_9416,N_9674);
or UO_72 (O_72,N_9365,N_9698);
and UO_73 (O_73,N_9987,N_9107);
or UO_74 (O_74,N_9920,N_9151);
and UO_75 (O_75,N_9414,N_9351);
nand UO_76 (O_76,N_9769,N_9979);
and UO_77 (O_77,N_9258,N_9028);
or UO_78 (O_78,N_9354,N_9573);
or UO_79 (O_79,N_9204,N_9082);
nand UO_80 (O_80,N_9045,N_9212);
and UO_81 (O_81,N_9893,N_9873);
and UO_82 (O_82,N_9050,N_9848);
nor UO_83 (O_83,N_9662,N_9505);
xnor UO_84 (O_84,N_9243,N_9973);
and UO_85 (O_85,N_9306,N_9694);
nor UO_86 (O_86,N_9302,N_9951);
or UO_87 (O_87,N_9485,N_9128);
nand UO_88 (O_88,N_9650,N_9863);
nand UO_89 (O_89,N_9060,N_9799);
and UO_90 (O_90,N_9604,N_9007);
or UO_91 (O_91,N_9109,N_9491);
nor UO_92 (O_92,N_9422,N_9984);
nand UO_93 (O_93,N_9321,N_9398);
and UO_94 (O_94,N_9535,N_9430);
and UO_95 (O_95,N_9449,N_9681);
or UO_96 (O_96,N_9942,N_9612);
nand UO_97 (O_97,N_9638,N_9395);
nor UO_98 (O_98,N_9770,N_9350);
or UO_99 (O_99,N_9804,N_9580);
or UO_100 (O_100,N_9296,N_9932);
or UO_101 (O_101,N_9840,N_9677);
nand UO_102 (O_102,N_9631,N_9288);
nand UO_103 (O_103,N_9735,N_9139);
or UO_104 (O_104,N_9919,N_9598);
and UO_105 (O_105,N_9327,N_9117);
and UO_106 (O_106,N_9599,N_9534);
or UO_107 (O_107,N_9158,N_9618);
or UO_108 (O_108,N_9994,N_9516);
nor UO_109 (O_109,N_9683,N_9330);
or UO_110 (O_110,N_9853,N_9995);
and UO_111 (O_111,N_9290,N_9701);
and UO_112 (O_112,N_9098,N_9295);
nand UO_113 (O_113,N_9503,N_9929);
and UO_114 (O_114,N_9765,N_9486);
nand UO_115 (O_115,N_9820,N_9639);
or UO_116 (O_116,N_9412,N_9874);
nor UO_117 (O_117,N_9197,N_9383);
nand UO_118 (O_118,N_9586,N_9621);
nor UO_119 (O_119,N_9137,N_9242);
nor UO_120 (O_120,N_9732,N_9703);
nand UO_121 (O_121,N_9632,N_9808);
nor UO_122 (O_122,N_9962,N_9813);
and UO_123 (O_123,N_9156,N_9459);
or UO_124 (O_124,N_9436,N_9164);
nand UO_125 (O_125,N_9555,N_9905);
nand UO_126 (O_126,N_9896,N_9511);
nand UO_127 (O_127,N_9577,N_9972);
nand UO_128 (O_128,N_9944,N_9669);
and UO_129 (O_129,N_9433,N_9917);
or UO_130 (O_130,N_9767,N_9457);
and UO_131 (O_131,N_9057,N_9869);
nand UO_132 (O_132,N_9364,N_9363);
nand UO_133 (O_133,N_9300,N_9731);
or UO_134 (O_134,N_9943,N_9214);
nand UO_135 (O_135,N_9806,N_9444);
nor UO_136 (O_136,N_9185,N_9931);
nor UO_137 (O_137,N_9901,N_9076);
or UO_138 (O_138,N_9891,N_9055);
or UO_139 (O_139,N_9191,N_9077);
nand UO_140 (O_140,N_9221,N_9928);
nand UO_141 (O_141,N_9607,N_9324);
or UO_142 (O_142,N_9183,N_9884);
or UO_143 (O_143,N_9784,N_9169);
nor UO_144 (O_144,N_9829,N_9781);
and UO_145 (O_145,N_9032,N_9635);
and UO_146 (O_146,N_9291,N_9360);
nand UO_147 (O_147,N_9458,N_9689);
and UO_148 (O_148,N_9738,N_9380);
and UO_149 (O_149,N_9340,N_9100);
or UO_150 (O_150,N_9666,N_9426);
or UO_151 (O_151,N_9883,N_9177);
and UO_152 (O_152,N_9790,N_9149);
nor UO_153 (O_153,N_9742,N_9101);
nand UO_154 (O_154,N_9624,N_9320);
nand UO_155 (O_155,N_9129,N_9574);
and UO_156 (O_156,N_9659,N_9219);
and UO_157 (O_157,N_9532,N_9333);
and UO_158 (O_158,N_9309,N_9376);
nor UO_159 (O_159,N_9093,N_9447);
or UO_160 (O_160,N_9115,N_9679);
or UO_161 (O_161,N_9130,N_9334);
nand UO_162 (O_162,N_9081,N_9879);
and UO_163 (O_163,N_9329,N_9397);
and UO_164 (O_164,N_9506,N_9331);
or UO_165 (O_165,N_9998,N_9424);
and UO_166 (O_166,N_9480,N_9993);
nor UO_167 (O_167,N_9696,N_9492);
xor UO_168 (O_168,N_9670,N_9909);
nor UO_169 (O_169,N_9600,N_9318);
and UO_170 (O_170,N_9978,N_9299);
nand UO_171 (O_171,N_9345,N_9125);
or UO_172 (O_172,N_9882,N_9895);
nor UO_173 (O_173,N_9440,N_9661);
nand UO_174 (O_174,N_9207,N_9849);
nor UO_175 (O_175,N_9649,N_9556);
nor UO_176 (O_176,N_9885,N_9721);
and UO_177 (O_177,N_9722,N_9856);
and UO_178 (O_178,N_9952,N_9445);
nor UO_179 (O_179,N_9179,N_9289);
and UO_180 (O_180,N_9469,N_9746);
or UO_181 (O_181,N_9563,N_9704);
nor UO_182 (O_182,N_9015,N_9509);
or UO_183 (O_183,N_9561,N_9851);
or UO_184 (O_184,N_9261,N_9569);
or UO_185 (O_185,N_9688,N_9611);
nand UO_186 (O_186,N_9894,N_9078);
nor UO_187 (O_187,N_9565,N_9572);
nor UO_188 (O_188,N_9140,N_9954);
or UO_189 (O_189,N_9379,N_9489);
and UO_190 (O_190,N_9052,N_9323);
nor UO_191 (O_191,N_9691,N_9934);
and UO_192 (O_192,N_9678,N_9797);
and UO_193 (O_193,N_9857,N_9039);
nor UO_194 (O_194,N_9542,N_9044);
nand UO_195 (O_195,N_9462,N_9898);
and UO_196 (O_196,N_9157,N_9190);
or UO_197 (O_197,N_9622,N_9969);
or UO_198 (O_198,N_9839,N_9001);
and UO_199 (O_199,N_9974,N_9652);
nor UO_200 (O_200,N_9539,N_9727);
or UO_201 (O_201,N_9803,N_9165);
and UO_202 (O_202,N_9723,N_9097);
nand UO_203 (O_203,N_9362,N_9712);
nand UO_204 (O_204,N_9921,N_9798);
nand UO_205 (O_205,N_9564,N_9428);
nor UO_206 (O_206,N_9531,N_9358);
nor UO_207 (O_207,N_9313,N_9933);
nor UO_208 (O_208,N_9361,N_9690);
nand UO_209 (O_209,N_9260,N_9027);
nand UO_210 (O_210,N_9619,N_9826);
and UO_211 (O_211,N_9461,N_9188);
or UO_212 (O_212,N_9238,N_9454);
nand UO_213 (O_213,N_9583,N_9037);
xor UO_214 (O_214,N_9346,N_9941);
nor UO_215 (O_215,N_9758,N_9903);
nand UO_216 (O_216,N_9982,N_9263);
and UO_217 (O_217,N_9114,N_9147);
and UO_218 (O_218,N_9824,N_9533);
or UO_219 (O_219,N_9996,N_9225);
nand UO_220 (O_220,N_9617,N_9588);
nand UO_221 (O_221,N_9025,N_9910);
or UO_222 (O_222,N_9945,N_9435);
and UO_223 (O_223,N_9581,N_9500);
nor UO_224 (O_224,N_9918,N_9199);
nand UO_225 (O_225,N_9629,N_9888);
and UO_226 (O_226,N_9418,N_9372);
nand UO_227 (O_227,N_9378,N_9682);
and UO_228 (O_228,N_9859,N_9757);
nand UO_229 (O_229,N_9860,N_9284);
nand UO_230 (O_230,N_9153,N_9837);
or UO_231 (O_231,N_9132,N_9481);
and UO_232 (O_232,N_9750,N_9591);
nor UO_233 (O_233,N_9626,N_9845);
nor UO_234 (O_234,N_9370,N_9867);
nand UO_235 (O_235,N_9788,N_9844);
nor UO_236 (O_236,N_9601,N_9069);
nor UO_237 (O_237,N_9695,N_9823);
nand UO_238 (O_238,N_9606,N_9587);
nor UO_239 (O_239,N_9776,N_9064);
nand UO_240 (O_240,N_9181,N_9720);
or UO_241 (O_241,N_9072,N_9106);
nor UO_242 (O_242,N_9687,N_9184);
or UO_243 (O_243,N_9452,N_9916);
or UO_244 (O_244,N_9785,N_9675);
nand UO_245 (O_245,N_9402,N_9075);
nor UO_246 (O_246,N_9053,N_9473);
nand UO_247 (O_247,N_9739,N_9759);
or UO_248 (O_248,N_9279,N_9123);
and UO_249 (O_249,N_9761,N_9748);
and UO_250 (O_250,N_9249,N_9861);
xor UO_251 (O_251,N_9091,N_9220);
nand UO_252 (O_252,N_9217,N_9355);
nand UO_253 (O_253,N_9644,N_9983);
nand UO_254 (O_254,N_9266,N_9831);
nand UO_255 (O_255,N_9322,N_9417);
or UO_256 (O_256,N_9603,N_9198);
and UO_257 (O_257,N_9878,N_9762);
nor UO_258 (O_258,N_9172,N_9832);
nand UO_259 (O_259,N_9178,N_9252);
and UO_260 (O_260,N_9167,N_9658);
nor UO_261 (O_261,N_9825,N_9120);
nor UO_262 (O_262,N_9124,N_9450);
or UO_263 (O_263,N_9768,N_9236);
nand UO_264 (O_264,N_9724,N_9809);
or UO_265 (O_265,N_9110,N_9443);
nand UO_266 (O_266,N_9253,N_9558);
or UO_267 (O_267,N_9566,N_9868);
nor UO_268 (O_268,N_9717,N_9287);
nor UO_269 (O_269,N_9453,N_9940);
or UO_270 (O_270,N_9890,N_9567);
nor UO_271 (O_271,N_9686,N_9640);
and UO_272 (O_272,N_9281,N_9881);
and UO_273 (O_273,N_9314,N_9294);
or UO_274 (O_274,N_9170,N_9557);
nor UO_275 (O_275,N_9773,N_9374);
or UO_276 (O_276,N_9636,N_9946);
nor UO_277 (O_277,N_9841,N_9957);
and UO_278 (O_278,N_9728,N_9387);
or UO_279 (O_279,N_9046,N_9019);
nor UO_280 (O_280,N_9925,N_9842);
and UO_281 (O_281,N_9189,N_9643);
nor UO_282 (O_282,N_9623,N_9482);
nand UO_283 (O_283,N_9159,N_9216);
nor UO_284 (O_284,N_9280,N_9111);
nor UO_285 (O_285,N_9700,N_9051);
nand UO_286 (O_286,N_9745,N_9858);
nand UO_287 (O_287,N_9013,N_9096);
or UO_288 (O_288,N_9549,N_9965);
and UO_289 (O_289,N_9789,N_9835);
nand UO_290 (O_290,N_9609,N_9171);
nor UO_291 (O_291,N_9203,N_9112);
nor UO_292 (O_292,N_9810,N_9515);
or UO_293 (O_293,N_9255,N_9571);
or UO_294 (O_294,N_9907,N_9226);
or UO_295 (O_295,N_9161,N_9655);
and UO_296 (O_296,N_9136,N_9922);
nand UO_297 (O_297,N_9176,N_9512);
nand UO_298 (O_298,N_9146,N_9305);
nor UO_299 (O_299,N_9259,N_9367);
nor UO_300 (O_300,N_9529,N_9070);
and UO_301 (O_301,N_9162,N_9419);
nor UO_302 (O_302,N_9795,N_9315);
nor UO_303 (O_303,N_9145,N_9272);
nand UO_304 (O_304,N_9396,N_9956);
nand UO_305 (O_305,N_9389,N_9546);
nand UO_306 (O_306,N_9743,N_9964);
nand UO_307 (O_307,N_9211,N_9740);
nor UO_308 (O_308,N_9817,N_9427);
nor UO_309 (O_309,N_9749,N_9285);
and UO_310 (O_310,N_9479,N_9021);
or UO_311 (O_311,N_9009,N_9911);
nor UO_312 (O_312,N_9180,N_9410);
or UO_313 (O_313,N_9846,N_9005);
nand UO_314 (O_314,N_9408,N_9900);
nand UO_315 (O_315,N_9886,N_9924);
nand UO_316 (O_316,N_9834,N_9411);
nor UO_317 (O_317,N_9282,N_9304);
or UO_318 (O_318,N_9935,N_9705);
and UO_319 (O_319,N_9576,N_9384);
nand UO_320 (O_320,N_9233,N_9830);
and UO_321 (O_321,N_9708,N_9783);
nor UO_322 (O_322,N_9989,N_9852);
and UO_323 (O_323,N_9332,N_9277);
and UO_324 (O_324,N_9499,N_9464);
or UO_325 (O_325,N_9008,N_9560);
nor UO_326 (O_326,N_9036,N_9000);
nand UO_327 (O_327,N_9201,N_9244);
nand UO_328 (O_328,N_9229,N_9421);
nand UO_329 (O_329,N_9760,N_9033);
or UO_330 (O_330,N_9526,N_9166);
nor UO_331 (O_331,N_9676,N_9337);
nor UO_332 (O_332,N_9404,N_9892);
xnor UO_333 (O_333,N_9297,N_9522);
and UO_334 (O_334,N_9257,N_9771);
nor UO_335 (O_335,N_9975,N_9985);
or UO_336 (O_336,N_9904,N_9960);
or UO_337 (O_337,N_9642,N_9476);
or UO_338 (O_338,N_9870,N_9210);
nor UO_339 (O_339,N_9756,N_9022);
nand UO_340 (O_340,N_9215,N_9990);
and UO_341 (O_341,N_9142,N_9310);
xnor UO_342 (O_342,N_9752,N_9232);
and UO_343 (O_343,N_9248,N_9206);
and UO_344 (O_344,N_9553,N_9570);
nor UO_345 (O_345,N_9981,N_9218);
and UO_346 (O_346,N_9668,N_9597);
or UO_347 (O_347,N_9246,N_9079);
or UO_348 (O_348,N_9352,N_9023);
and UO_349 (O_349,N_9063,N_9519);
nor UO_350 (O_350,N_9754,N_9386);
nand UO_351 (O_351,N_9501,N_9080);
or UO_352 (O_352,N_9502,N_9065);
nand UO_353 (O_353,N_9780,N_9791);
nor UO_354 (O_354,N_9041,N_9173);
nand UO_355 (O_355,N_9613,N_9406);
or UO_356 (O_356,N_9986,N_9105);
or UO_357 (O_357,N_9543,N_9451);
or UO_358 (O_358,N_9528,N_9741);
or UO_359 (O_359,N_9405,N_9108);
nor UO_360 (O_360,N_9138,N_9150);
nor UO_361 (O_361,N_9131,N_9899);
and UO_362 (O_362,N_9195,N_9339);
or UO_363 (O_363,N_9024,N_9127);
nor UO_364 (O_364,N_9040,N_9102);
xor UO_365 (O_365,N_9897,N_9048);
nand UO_366 (O_366,N_9955,N_9439);
or UO_367 (O_367,N_9224,N_9778);
nor UO_368 (O_368,N_9336,N_9466);
nand UO_369 (O_369,N_9152,N_9766);
nor UO_370 (O_370,N_9847,N_9947);
and UO_371 (O_371,N_9966,N_9545);
or UO_372 (O_372,N_9718,N_9175);
nand UO_373 (O_373,N_9470,N_9530);
and UO_374 (O_374,N_9192,N_9801);
nor UO_375 (O_375,N_9812,N_9715);
nor UO_376 (O_376,N_9575,N_9003);
nand UO_377 (O_377,N_9725,N_9031);
or UO_378 (O_378,N_9382,N_9596);
nor UO_379 (O_379,N_9085,N_9271);
and UO_380 (O_380,N_9488,N_9475);
xnor UO_381 (O_381,N_9043,N_9495);
nor UO_382 (O_382,N_9551,N_9961);
or UO_383 (O_383,N_9437,N_9641);
nor UO_384 (O_384,N_9819,N_9223);
nor UO_385 (O_385,N_9697,N_9092);
nand UO_386 (O_386,N_9667,N_9163);
nand UO_387 (O_387,N_9034,N_9751);
nand UO_388 (O_388,N_9126,N_9620);
xnor UO_389 (O_389,N_9086,N_9235);
or UO_390 (O_390,N_9254,N_9018);
and UO_391 (O_391,N_9415,N_9344);
nor UO_392 (O_392,N_9646,N_9375);
and UO_393 (O_393,N_9653,N_9317);
and UO_394 (O_394,N_9645,N_9237);
and UO_395 (O_395,N_9403,N_9227);
nor UO_396 (O_396,N_9541,N_9880);
and UO_397 (O_397,N_9648,N_9793);
nand UO_398 (O_398,N_9089,N_9936);
nand UO_399 (O_399,N_9276,N_9707);
nor UO_400 (O_400,N_9971,N_9265);
and UO_401 (O_401,N_9017,N_9099);
or UO_402 (O_402,N_9513,N_9413);
nor UO_403 (O_403,N_9672,N_9335);
and UO_404 (O_404,N_9390,N_9838);
and UO_405 (O_405,N_9356,N_9589);
nand UO_406 (O_406,N_9144,N_9816);
and UO_407 (O_407,N_9926,N_9186);
nand UO_408 (O_408,N_9429,N_9796);
nand UO_409 (O_409,N_9906,N_9368);
or UO_410 (O_410,N_9460,N_9200);
or UO_411 (O_411,N_9084,N_9400);
nand UO_412 (O_412,N_9490,N_9792);
nand UO_413 (O_413,N_9772,N_9614);
and UO_414 (O_414,N_9160,N_9061);
nor UO_415 (O_415,N_9071,N_9584);
or UO_416 (O_416,N_9446,N_9525);
nor UO_417 (O_417,N_9871,N_9133);
nor UO_418 (O_418,N_9608,N_9116);
and UO_419 (O_419,N_9510,N_9155);
nor UO_420 (O_420,N_9997,N_9208);
nor UO_421 (O_421,N_9734,N_9456);
nor UO_422 (O_422,N_9959,N_9930);
and UO_423 (O_423,N_9038,N_9711);
and UO_424 (O_424,N_9316,N_9002);
nand UO_425 (O_425,N_9913,N_9568);
nand UO_426 (O_426,N_9948,N_9544);
nand UO_427 (O_427,N_9154,N_9205);
or UO_428 (O_428,N_9231,N_9477);
and UO_429 (O_429,N_9963,N_9559);
or UO_430 (O_430,N_9967,N_9143);
nand UO_431 (O_431,N_9782,N_9303);
nand UO_432 (O_432,N_9578,N_9141);
and UO_433 (O_433,N_9087,N_9923);
nor UO_434 (O_434,N_9887,N_9827);
nor UO_435 (O_435,N_9949,N_9889);
nor UO_436 (O_436,N_9864,N_9937);
and UO_437 (O_437,N_9311,N_9442);
nor UO_438 (O_438,N_9062,N_9753);
or UO_439 (O_439,N_9262,N_9068);
or UO_440 (O_440,N_9634,N_9992);
and UO_441 (O_441,N_9685,N_9865);
or UO_442 (O_442,N_9939,N_9628);
nand UO_443 (O_443,N_9095,N_9665);
and UO_444 (O_444,N_9657,N_9030);
or UO_445 (O_445,N_9950,N_9821);
nor UO_446 (O_446,N_9196,N_9202);
nor UO_447 (O_447,N_9247,N_9664);
nor UO_448 (O_448,N_9423,N_9590);
nand UO_449 (O_449,N_9651,N_9393);
nand UO_450 (O_450,N_9710,N_9862);
nor UO_451 (O_451,N_9736,N_9298);
nand UO_452 (O_452,N_9012,N_9359);
xnor UO_453 (O_453,N_9193,N_9605);
nor UO_454 (O_454,N_9872,N_9014);
and UO_455 (O_455,N_9706,N_9328);
xor UO_456 (O_456,N_9497,N_9434);
nor UO_457 (O_457,N_9273,N_9463);
nor UO_458 (O_458,N_9496,N_9562);
or UO_459 (O_459,N_9554,N_9716);
and UO_460 (O_460,N_9059,N_9777);
or UO_461 (O_461,N_9517,N_9420);
nor UO_462 (O_462,N_9366,N_9425);
nor UO_463 (O_463,N_9407,N_9786);
and UO_464 (O_464,N_9656,N_9988);
and UO_465 (O_465,N_9066,N_9010);
nor UO_466 (O_466,N_9680,N_9441);
nand UO_467 (O_467,N_9264,N_9494);
nand UO_468 (O_468,N_9401,N_9908);
and UO_469 (O_469,N_9593,N_9122);
nand UO_470 (O_470,N_9029,N_9518);
or UO_471 (O_471,N_9286,N_9654);
nor UO_472 (O_472,N_9714,N_9504);
nand UO_473 (O_473,N_9168,N_9953);
nor UO_474 (O_474,N_9794,N_9527);
and UO_475 (O_475,N_9976,N_9747);
nand UO_476 (O_476,N_9647,N_9118);
or UO_477 (O_477,N_9292,N_9633);
nand UO_478 (O_478,N_9338,N_9693);
and UO_479 (O_479,N_9547,N_9779);
or UO_480 (O_480,N_9270,N_9914);
nand UO_481 (O_481,N_9067,N_9228);
nand UO_482 (O_482,N_9616,N_9267);
nand UO_483 (O_483,N_9432,N_9875);
or UO_484 (O_484,N_9484,N_9805);
or UO_485 (O_485,N_9083,N_9968);
or UO_486 (O_486,N_9006,N_9818);
and UO_487 (O_487,N_9073,N_9250);
and UO_488 (O_488,N_9673,N_9671);
or UO_489 (O_489,N_9774,N_9520);
nand UO_490 (O_490,N_9187,N_9744);
nand UO_491 (O_491,N_9498,N_9357);
or UO_492 (O_492,N_9094,N_9902);
nor UO_493 (O_493,N_9353,N_9020);
or UO_494 (O_494,N_9326,N_9692);
nor UO_495 (O_495,N_9209,N_9256);
nand UO_496 (O_496,N_9381,N_9474);
or UO_497 (O_497,N_9579,N_9319);
nor UO_498 (O_498,N_9729,N_9472);
nand UO_499 (O_499,N_9455,N_9615);
nor UO_500 (O_500,N_9206,N_9940);
nor UO_501 (O_501,N_9179,N_9386);
nor UO_502 (O_502,N_9117,N_9145);
or UO_503 (O_503,N_9932,N_9395);
or UO_504 (O_504,N_9205,N_9301);
nor UO_505 (O_505,N_9713,N_9522);
or UO_506 (O_506,N_9716,N_9479);
nand UO_507 (O_507,N_9666,N_9943);
nor UO_508 (O_508,N_9072,N_9105);
nand UO_509 (O_509,N_9296,N_9222);
or UO_510 (O_510,N_9764,N_9919);
or UO_511 (O_511,N_9915,N_9313);
and UO_512 (O_512,N_9075,N_9260);
and UO_513 (O_513,N_9071,N_9739);
or UO_514 (O_514,N_9967,N_9065);
and UO_515 (O_515,N_9651,N_9697);
nand UO_516 (O_516,N_9320,N_9318);
nor UO_517 (O_517,N_9960,N_9911);
and UO_518 (O_518,N_9827,N_9692);
and UO_519 (O_519,N_9520,N_9418);
or UO_520 (O_520,N_9678,N_9767);
or UO_521 (O_521,N_9494,N_9104);
or UO_522 (O_522,N_9248,N_9382);
or UO_523 (O_523,N_9817,N_9398);
nand UO_524 (O_524,N_9177,N_9434);
nand UO_525 (O_525,N_9965,N_9817);
and UO_526 (O_526,N_9578,N_9164);
nand UO_527 (O_527,N_9793,N_9236);
nor UO_528 (O_528,N_9150,N_9539);
and UO_529 (O_529,N_9748,N_9298);
nand UO_530 (O_530,N_9055,N_9494);
and UO_531 (O_531,N_9007,N_9077);
or UO_532 (O_532,N_9235,N_9106);
nor UO_533 (O_533,N_9180,N_9342);
and UO_534 (O_534,N_9876,N_9931);
or UO_535 (O_535,N_9012,N_9085);
or UO_536 (O_536,N_9564,N_9318);
nand UO_537 (O_537,N_9881,N_9180);
and UO_538 (O_538,N_9572,N_9825);
nor UO_539 (O_539,N_9366,N_9512);
nand UO_540 (O_540,N_9266,N_9762);
nor UO_541 (O_541,N_9513,N_9549);
or UO_542 (O_542,N_9691,N_9003);
nor UO_543 (O_543,N_9350,N_9935);
and UO_544 (O_544,N_9644,N_9440);
nor UO_545 (O_545,N_9236,N_9628);
and UO_546 (O_546,N_9710,N_9443);
or UO_547 (O_547,N_9335,N_9062);
and UO_548 (O_548,N_9833,N_9391);
or UO_549 (O_549,N_9446,N_9697);
and UO_550 (O_550,N_9294,N_9673);
and UO_551 (O_551,N_9567,N_9459);
and UO_552 (O_552,N_9501,N_9492);
or UO_553 (O_553,N_9673,N_9308);
and UO_554 (O_554,N_9049,N_9385);
and UO_555 (O_555,N_9083,N_9431);
nor UO_556 (O_556,N_9931,N_9918);
nor UO_557 (O_557,N_9607,N_9728);
nor UO_558 (O_558,N_9814,N_9172);
or UO_559 (O_559,N_9887,N_9578);
and UO_560 (O_560,N_9823,N_9922);
and UO_561 (O_561,N_9557,N_9507);
nor UO_562 (O_562,N_9415,N_9025);
or UO_563 (O_563,N_9126,N_9393);
nand UO_564 (O_564,N_9243,N_9062);
or UO_565 (O_565,N_9988,N_9148);
nor UO_566 (O_566,N_9721,N_9024);
nor UO_567 (O_567,N_9459,N_9264);
and UO_568 (O_568,N_9455,N_9003);
nor UO_569 (O_569,N_9495,N_9065);
xnor UO_570 (O_570,N_9441,N_9594);
and UO_571 (O_571,N_9883,N_9884);
nand UO_572 (O_572,N_9895,N_9222);
or UO_573 (O_573,N_9119,N_9557);
and UO_574 (O_574,N_9129,N_9345);
nand UO_575 (O_575,N_9759,N_9928);
or UO_576 (O_576,N_9692,N_9699);
nor UO_577 (O_577,N_9447,N_9946);
nand UO_578 (O_578,N_9716,N_9074);
nand UO_579 (O_579,N_9132,N_9914);
or UO_580 (O_580,N_9555,N_9040);
nand UO_581 (O_581,N_9425,N_9618);
and UO_582 (O_582,N_9782,N_9786);
nor UO_583 (O_583,N_9554,N_9732);
nand UO_584 (O_584,N_9425,N_9414);
nand UO_585 (O_585,N_9906,N_9949);
nor UO_586 (O_586,N_9232,N_9419);
nor UO_587 (O_587,N_9344,N_9135);
and UO_588 (O_588,N_9781,N_9317);
and UO_589 (O_589,N_9206,N_9156);
nor UO_590 (O_590,N_9403,N_9889);
nor UO_591 (O_591,N_9497,N_9069);
nand UO_592 (O_592,N_9633,N_9661);
nand UO_593 (O_593,N_9898,N_9087);
and UO_594 (O_594,N_9317,N_9039);
or UO_595 (O_595,N_9356,N_9716);
nand UO_596 (O_596,N_9199,N_9184);
or UO_597 (O_597,N_9845,N_9638);
nand UO_598 (O_598,N_9294,N_9586);
xor UO_599 (O_599,N_9108,N_9481);
or UO_600 (O_600,N_9595,N_9407);
or UO_601 (O_601,N_9474,N_9345);
and UO_602 (O_602,N_9486,N_9833);
nor UO_603 (O_603,N_9979,N_9930);
and UO_604 (O_604,N_9946,N_9178);
or UO_605 (O_605,N_9100,N_9706);
nor UO_606 (O_606,N_9163,N_9399);
nor UO_607 (O_607,N_9237,N_9933);
nand UO_608 (O_608,N_9707,N_9795);
nand UO_609 (O_609,N_9485,N_9078);
nand UO_610 (O_610,N_9143,N_9393);
or UO_611 (O_611,N_9463,N_9695);
or UO_612 (O_612,N_9858,N_9607);
and UO_613 (O_613,N_9163,N_9746);
or UO_614 (O_614,N_9280,N_9184);
and UO_615 (O_615,N_9414,N_9469);
nor UO_616 (O_616,N_9462,N_9278);
nand UO_617 (O_617,N_9493,N_9383);
nand UO_618 (O_618,N_9689,N_9505);
nand UO_619 (O_619,N_9079,N_9372);
or UO_620 (O_620,N_9053,N_9387);
and UO_621 (O_621,N_9428,N_9753);
nor UO_622 (O_622,N_9850,N_9761);
or UO_623 (O_623,N_9243,N_9659);
and UO_624 (O_624,N_9483,N_9897);
nand UO_625 (O_625,N_9150,N_9125);
nor UO_626 (O_626,N_9310,N_9567);
nand UO_627 (O_627,N_9812,N_9033);
nor UO_628 (O_628,N_9016,N_9218);
xor UO_629 (O_629,N_9780,N_9016);
nor UO_630 (O_630,N_9377,N_9473);
and UO_631 (O_631,N_9354,N_9691);
nand UO_632 (O_632,N_9262,N_9807);
nand UO_633 (O_633,N_9783,N_9911);
nor UO_634 (O_634,N_9216,N_9813);
nor UO_635 (O_635,N_9381,N_9460);
nand UO_636 (O_636,N_9337,N_9179);
and UO_637 (O_637,N_9413,N_9725);
or UO_638 (O_638,N_9242,N_9033);
xor UO_639 (O_639,N_9034,N_9463);
and UO_640 (O_640,N_9558,N_9088);
or UO_641 (O_641,N_9792,N_9675);
nand UO_642 (O_642,N_9235,N_9550);
or UO_643 (O_643,N_9723,N_9368);
nor UO_644 (O_644,N_9593,N_9248);
nor UO_645 (O_645,N_9435,N_9586);
or UO_646 (O_646,N_9599,N_9433);
nor UO_647 (O_647,N_9837,N_9378);
or UO_648 (O_648,N_9256,N_9051);
and UO_649 (O_649,N_9507,N_9091);
nand UO_650 (O_650,N_9899,N_9329);
nor UO_651 (O_651,N_9558,N_9768);
nor UO_652 (O_652,N_9883,N_9125);
and UO_653 (O_653,N_9027,N_9637);
and UO_654 (O_654,N_9776,N_9655);
nand UO_655 (O_655,N_9897,N_9363);
nand UO_656 (O_656,N_9536,N_9157);
or UO_657 (O_657,N_9580,N_9400);
and UO_658 (O_658,N_9913,N_9775);
or UO_659 (O_659,N_9630,N_9339);
or UO_660 (O_660,N_9396,N_9257);
nand UO_661 (O_661,N_9477,N_9881);
or UO_662 (O_662,N_9496,N_9461);
and UO_663 (O_663,N_9633,N_9736);
nor UO_664 (O_664,N_9922,N_9825);
and UO_665 (O_665,N_9527,N_9615);
and UO_666 (O_666,N_9401,N_9642);
nand UO_667 (O_667,N_9286,N_9167);
nor UO_668 (O_668,N_9665,N_9770);
nand UO_669 (O_669,N_9083,N_9469);
nand UO_670 (O_670,N_9453,N_9456);
nand UO_671 (O_671,N_9003,N_9942);
nand UO_672 (O_672,N_9419,N_9428);
or UO_673 (O_673,N_9596,N_9721);
nand UO_674 (O_674,N_9332,N_9894);
or UO_675 (O_675,N_9501,N_9099);
or UO_676 (O_676,N_9533,N_9927);
and UO_677 (O_677,N_9064,N_9745);
nand UO_678 (O_678,N_9963,N_9576);
or UO_679 (O_679,N_9981,N_9409);
and UO_680 (O_680,N_9753,N_9244);
and UO_681 (O_681,N_9372,N_9576);
nor UO_682 (O_682,N_9351,N_9082);
nor UO_683 (O_683,N_9371,N_9190);
or UO_684 (O_684,N_9206,N_9607);
xor UO_685 (O_685,N_9468,N_9100);
nor UO_686 (O_686,N_9279,N_9852);
and UO_687 (O_687,N_9129,N_9335);
and UO_688 (O_688,N_9928,N_9994);
nor UO_689 (O_689,N_9640,N_9607);
or UO_690 (O_690,N_9204,N_9127);
nor UO_691 (O_691,N_9175,N_9931);
nor UO_692 (O_692,N_9093,N_9484);
nand UO_693 (O_693,N_9451,N_9827);
and UO_694 (O_694,N_9462,N_9415);
nor UO_695 (O_695,N_9779,N_9402);
or UO_696 (O_696,N_9203,N_9270);
nand UO_697 (O_697,N_9135,N_9571);
or UO_698 (O_698,N_9878,N_9355);
nor UO_699 (O_699,N_9667,N_9428);
and UO_700 (O_700,N_9419,N_9425);
or UO_701 (O_701,N_9579,N_9889);
and UO_702 (O_702,N_9720,N_9870);
or UO_703 (O_703,N_9777,N_9545);
nor UO_704 (O_704,N_9339,N_9202);
or UO_705 (O_705,N_9310,N_9799);
or UO_706 (O_706,N_9675,N_9065);
nor UO_707 (O_707,N_9100,N_9834);
and UO_708 (O_708,N_9760,N_9467);
nor UO_709 (O_709,N_9281,N_9559);
nand UO_710 (O_710,N_9014,N_9619);
or UO_711 (O_711,N_9331,N_9027);
nand UO_712 (O_712,N_9380,N_9134);
or UO_713 (O_713,N_9740,N_9508);
or UO_714 (O_714,N_9459,N_9215);
nand UO_715 (O_715,N_9954,N_9446);
and UO_716 (O_716,N_9556,N_9914);
or UO_717 (O_717,N_9237,N_9876);
or UO_718 (O_718,N_9568,N_9377);
and UO_719 (O_719,N_9007,N_9110);
nor UO_720 (O_720,N_9314,N_9898);
nand UO_721 (O_721,N_9605,N_9427);
nand UO_722 (O_722,N_9429,N_9695);
or UO_723 (O_723,N_9841,N_9474);
or UO_724 (O_724,N_9620,N_9556);
nand UO_725 (O_725,N_9946,N_9097);
or UO_726 (O_726,N_9909,N_9841);
or UO_727 (O_727,N_9059,N_9816);
or UO_728 (O_728,N_9167,N_9324);
or UO_729 (O_729,N_9474,N_9450);
nand UO_730 (O_730,N_9049,N_9844);
and UO_731 (O_731,N_9706,N_9120);
or UO_732 (O_732,N_9329,N_9202);
or UO_733 (O_733,N_9055,N_9276);
or UO_734 (O_734,N_9452,N_9872);
nor UO_735 (O_735,N_9973,N_9458);
nand UO_736 (O_736,N_9563,N_9825);
or UO_737 (O_737,N_9608,N_9706);
nor UO_738 (O_738,N_9274,N_9060);
nand UO_739 (O_739,N_9788,N_9928);
and UO_740 (O_740,N_9643,N_9996);
nor UO_741 (O_741,N_9198,N_9254);
nor UO_742 (O_742,N_9566,N_9461);
and UO_743 (O_743,N_9897,N_9545);
and UO_744 (O_744,N_9983,N_9021);
and UO_745 (O_745,N_9126,N_9634);
nor UO_746 (O_746,N_9687,N_9037);
and UO_747 (O_747,N_9109,N_9625);
nor UO_748 (O_748,N_9015,N_9241);
nand UO_749 (O_749,N_9661,N_9395);
or UO_750 (O_750,N_9403,N_9331);
or UO_751 (O_751,N_9187,N_9867);
nor UO_752 (O_752,N_9879,N_9465);
or UO_753 (O_753,N_9847,N_9766);
nor UO_754 (O_754,N_9483,N_9228);
nor UO_755 (O_755,N_9317,N_9916);
and UO_756 (O_756,N_9204,N_9546);
nor UO_757 (O_757,N_9804,N_9775);
nor UO_758 (O_758,N_9657,N_9927);
nor UO_759 (O_759,N_9170,N_9635);
nor UO_760 (O_760,N_9084,N_9099);
nand UO_761 (O_761,N_9007,N_9621);
nand UO_762 (O_762,N_9878,N_9141);
nor UO_763 (O_763,N_9315,N_9337);
or UO_764 (O_764,N_9163,N_9747);
nor UO_765 (O_765,N_9590,N_9308);
nor UO_766 (O_766,N_9234,N_9961);
nor UO_767 (O_767,N_9743,N_9666);
nand UO_768 (O_768,N_9426,N_9079);
nand UO_769 (O_769,N_9468,N_9742);
nor UO_770 (O_770,N_9620,N_9047);
or UO_771 (O_771,N_9846,N_9455);
or UO_772 (O_772,N_9146,N_9406);
nor UO_773 (O_773,N_9456,N_9611);
nor UO_774 (O_774,N_9387,N_9419);
and UO_775 (O_775,N_9892,N_9426);
or UO_776 (O_776,N_9593,N_9888);
and UO_777 (O_777,N_9148,N_9929);
and UO_778 (O_778,N_9769,N_9432);
nor UO_779 (O_779,N_9180,N_9122);
or UO_780 (O_780,N_9259,N_9171);
and UO_781 (O_781,N_9153,N_9941);
or UO_782 (O_782,N_9503,N_9159);
nor UO_783 (O_783,N_9207,N_9543);
nand UO_784 (O_784,N_9599,N_9012);
nand UO_785 (O_785,N_9876,N_9199);
or UO_786 (O_786,N_9837,N_9579);
or UO_787 (O_787,N_9916,N_9041);
nor UO_788 (O_788,N_9072,N_9558);
and UO_789 (O_789,N_9836,N_9448);
nor UO_790 (O_790,N_9463,N_9812);
nand UO_791 (O_791,N_9456,N_9762);
nand UO_792 (O_792,N_9125,N_9872);
nor UO_793 (O_793,N_9468,N_9617);
and UO_794 (O_794,N_9228,N_9096);
and UO_795 (O_795,N_9994,N_9106);
nand UO_796 (O_796,N_9101,N_9436);
and UO_797 (O_797,N_9970,N_9203);
nor UO_798 (O_798,N_9229,N_9659);
nor UO_799 (O_799,N_9135,N_9086);
or UO_800 (O_800,N_9231,N_9908);
nor UO_801 (O_801,N_9252,N_9859);
or UO_802 (O_802,N_9425,N_9358);
nand UO_803 (O_803,N_9579,N_9412);
or UO_804 (O_804,N_9434,N_9893);
nand UO_805 (O_805,N_9500,N_9048);
and UO_806 (O_806,N_9394,N_9247);
nor UO_807 (O_807,N_9285,N_9602);
nand UO_808 (O_808,N_9281,N_9120);
and UO_809 (O_809,N_9477,N_9425);
or UO_810 (O_810,N_9215,N_9879);
or UO_811 (O_811,N_9640,N_9479);
or UO_812 (O_812,N_9259,N_9943);
or UO_813 (O_813,N_9385,N_9469);
nand UO_814 (O_814,N_9377,N_9756);
and UO_815 (O_815,N_9993,N_9919);
or UO_816 (O_816,N_9169,N_9016);
nand UO_817 (O_817,N_9570,N_9321);
and UO_818 (O_818,N_9904,N_9840);
and UO_819 (O_819,N_9330,N_9608);
and UO_820 (O_820,N_9584,N_9638);
or UO_821 (O_821,N_9150,N_9740);
nand UO_822 (O_822,N_9558,N_9817);
nor UO_823 (O_823,N_9533,N_9396);
nand UO_824 (O_824,N_9150,N_9056);
or UO_825 (O_825,N_9354,N_9985);
nor UO_826 (O_826,N_9139,N_9203);
or UO_827 (O_827,N_9750,N_9167);
and UO_828 (O_828,N_9453,N_9733);
and UO_829 (O_829,N_9362,N_9938);
nor UO_830 (O_830,N_9716,N_9821);
or UO_831 (O_831,N_9457,N_9956);
nand UO_832 (O_832,N_9387,N_9916);
or UO_833 (O_833,N_9281,N_9937);
nor UO_834 (O_834,N_9669,N_9831);
nand UO_835 (O_835,N_9136,N_9691);
and UO_836 (O_836,N_9170,N_9227);
or UO_837 (O_837,N_9395,N_9042);
or UO_838 (O_838,N_9329,N_9124);
nand UO_839 (O_839,N_9695,N_9754);
nand UO_840 (O_840,N_9336,N_9650);
or UO_841 (O_841,N_9072,N_9857);
nor UO_842 (O_842,N_9495,N_9765);
nand UO_843 (O_843,N_9001,N_9497);
xnor UO_844 (O_844,N_9366,N_9615);
nand UO_845 (O_845,N_9322,N_9425);
nor UO_846 (O_846,N_9645,N_9931);
and UO_847 (O_847,N_9258,N_9095);
and UO_848 (O_848,N_9886,N_9368);
nor UO_849 (O_849,N_9045,N_9202);
nor UO_850 (O_850,N_9734,N_9900);
and UO_851 (O_851,N_9756,N_9428);
nand UO_852 (O_852,N_9184,N_9257);
nor UO_853 (O_853,N_9650,N_9324);
nor UO_854 (O_854,N_9192,N_9364);
nand UO_855 (O_855,N_9014,N_9063);
and UO_856 (O_856,N_9712,N_9635);
and UO_857 (O_857,N_9826,N_9635);
xor UO_858 (O_858,N_9963,N_9434);
or UO_859 (O_859,N_9687,N_9405);
nor UO_860 (O_860,N_9528,N_9869);
nand UO_861 (O_861,N_9151,N_9507);
nor UO_862 (O_862,N_9943,N_9966);
and UO_863 (O_863,N_9733,N_9599);
and UO_864 (O_864,N_9304,N_9416);
or UO_865 (O_865,N_9336,N_9104);
or UO_866 (O_866,N_9195,N_9990);
and UO_867 (O_867,N_9568,N_9299);
or UO_868 (O_868,N_9713,N_9200);
or UO_869 (O_869,N_9065,N_9979);
or UO_870 (O_870,N_9914,N_9793);
or UO_871 (O_871,N_9966,N_9947);
nand UO_872 (O_872,N_9370,N_9580);
nor UO_873 (O_873,N_9953,N_9870);
nand UO_874 (O_874,N_9122,N_9860);
nor UO_875 (O_875,N_9014,N_9156);
nand UO_876 (O_876,N_9121,N_9861);
and UO_877 (O_877,N_9524,N_9940);
nor UO_878 (O_878,N_9901,N_9653);
and UO_879 (O_879,N_9862,N_9731);
nand UO_880 (O_880,N_9532,N_9922);
nand UO_881 (O_881,N_9636,N_9573);
and UO_882 (O_882,N_9791,N_9775);
nand UO_883 (O_883,N_9528,N_9391);
or UO_884 (O_884,N_9837,N_9122);
or UO_885 (O_885,N_9420,N_9767);
or UO_886 (O_886,N_9504,N_9330);
nand UO_887 (O_887,N_9488,N_9507);
nand UO_888 (O_888,N_9127,N_9323);
nand UO_889 (O_889,N_9001,N_9900);
or UO_890 (O_890,N_9966,N_9713);
and UO_891 (O_891,N_9976,N_9741);
nor UO_892 (O_892,N_9843,N_9473);
nor UO_893 (O_893,N_9017,N_9957);
xnor UO_894 (O_894,N_9104,N_9161);
nand UO_895 (O_895,N_9678,N_9317);
and UO_896 (O_896,N_9001,N_9467);
and UO_897 (O_897,N_9475,N_9916);
nand UO_898 (O_898,N_9784,N_9183);
nand UO_899 (O_899,N_9067,N_9743);
and UO_900 (O_900,N_9923,N_9105);
nand UO_901 (O_901,N_9815,N_9968);
nor UO_902 (O_902,N_9159,N_9331);
or UO_903 (O_903,N_9675,N_9285);
nand UO_904 (O_904,N_9261,N_9673);
or UO_905 (O_905,N_9064,N_9236);
nor UO_906 (O_906,N_9309,N_9374);
nor UO_907 (O_907,N_9002,N_9062);
or UO_908 (O_908,N_9666,N_9287);
and UO_909 (O_909,N_9126,N_9008);
and UO_910 (O_910,N_9123,N_9381);
and UO_911 (O_911,N_9279,N_9477);
and UO_912 (O_912,N_9254,N_9620);
nor UO_913 (O_913,N_9723,N_9343);
and UO_914 (O_914,N_9420,N_9433);
nand UO_915 (O_915,N_9969,N_9867);
nand UO_916 (O_916,N_9857,N_9376);
nor UO_917 (O_917,N_9211,N_9099);
and UO_918 (O_918,N_9102,N_9002);
nand UO_919 (O_919,N_9978,N_9657);
nor UO_920 (O_920,N_9743,N_9889);
or UO_921 (O_921,N_9211,N_9732);
and UO_922 (O_922,N_9166,N_9953);
and UO_923 (O_923,N_9985,N_9486);
nand UO_924 (O_924,N_9887,N_9435);
or UO_925 (O_925,N_9574,N_9722);
and UO_926 (O_926,N_9982,N_9659);
nand UO_927 (O_927,N_9038,N_9745);
nand UO_928 (O_928,N_9669,N_9997);
and UO_929 (O_929,N_9510,N_9478);
and UO_930 (O_930,N_9007,N_9808);
nor UO_931 (O_931,N_9304,N_9257);
nor UO_932 (O_932,N_9278,N_9445);
nor UO_933 (O_933,N_9405,N_9704);
nor UO_934 (O_934,N_9985,N_9461);
nor UO_935 (O_935,N_9778,N_9411);
and UO_936 (O_936,N_9152,N_9269);
nand UO_937 (O_937,N_9577,N_9470);
or UO_938 (O_938,N_9941,N_9948);
or UO_939 (O_939,N_9118,N_9228);
nand UO_940 (O_940,N_9777,N_9421);
nor UO_941 (O_941,N_9221,N_9466);
nor UO_942 (O_942,N_9039,N_9141);
or UO_943 (O_943,N_9286,N_9418);
or UO_944 (O_944,N_9661,N_9955);
or UO_945 (O_945,N_9881,N_9799);
nand UO_946 (O_946,N_9356,N_9785);
nor UO_947 (O_947,N_9529,N_9992);
nand UO_948 (O_948,N_9496,N_9853);
and UO_949 (O_949,N_9271,N_9586);
nor UO_950 (O_950,N_9493,N_9864);
and UO_951 (O_951,N_9394,N_9726);
nand UO_952 (O_952,N_9756,N_9118);
nand UO_953 (O_953,N_9957,N_9011);
and UO_954 (O_954,N_9028,N_9937);
or UO_955 (O_955,N_9142,N_9548);
and UO_956 (O_956,N_9031,N_9204);
or UO_957 (O_957,N_9952,N_9214);
nand UO_958 (O_958,N_9650,N_9762);
nor UO_959 (O_959,N_9070,N_9300);
or UO_960 (O_960,N_9811,N_9161);
nor UO_961 (O_961,N_9770,N_9569);
nand UO_962 (O_962,N_9613,N_9789);
nand UO_963 (O_963,N_9060,N_9496);
and UO_964 (O_964,N_9440,N_9030);
nand UO_965 (O_965,N_9574,N_9788);
nor UO_966 (O_966,N_9861,N_9006);
nand UO_967 (O_967,N_9446,N_9615);
nor UO_968 (O_968,N_9836,N_9102);
and UO_969 (O_969,N_9819,N_9340);
nand UO_970 (O_970,N_9856,N_9381);
nor UO_971 (O_971,N_9224,N_9122);
nand UO_972 (O_972,N_9193,N_9311);
nand UO_973 (O_973,N_9057,N_9826);
nor UO_974 (O_974,N_9829,N_9238);
or UO_975 (O_975,N_9107,N_9653);
and UO_976 (O_976,N_9615,N_9934);
nand UO_977 (O_977,N_9811,N_9366);
nand UO_978 (O_978,N_9674,N_9684);
nor UO_979 (O_979,N_9530,N_9553);
nor UO_980 (O_980,N_9342,N_9064);
or UO_981 (O_981,N_9134,N_9739);
or UO_982 (O_982,N_9510,N_9867);
nand UO_983 (O_983,N_9216,N_9939);
and UO_984 (O_984,N_9293,N_9216);
or UO_985 (O_985,N_9226,N_9152);
nor UO_986 (O_986,N_9221,N_9090);
nor UO_987 (O_987,N_9736,N_9758);
and UO_988 (O_988,N_9993,N_9538);
or UO_989 (O_989,N_9465,N_9050);
and UO_990 (O_990,N_9723,N_9810);
nand UO_991 (O_991,N_9747,N_9152);
and UO_992 (O_992,N_9167,N_9883);
nand UO_993 (O_993,N_9529,N_9963);
nand UO_994 (O_994,N_9403,N_9633);
nand UO_995 (O_995,N_9402,N_9309);
or UO_996 (O_996,N_9259,N_9807);
nand UO_997 (O_997,N_9751,N_9588);
or UO_998 (O_998,N_9199,N_9005);
and UO_999 (O_999,N_9331,N_9875);
or UO_1000 (O_1000,N_9580,N_9605);
and UO_1001 (O_1001,N_9211,N_9938);
nand UO_1002 (O_1002,N_9592,N_9786);
or UO_1003 (O_1003,N_9299,N_9077);
and UO_1004 (O_1004,N_9388,N_9956);
nand UO_1005 (O_1005,N_9745,N_9870);
nor UO_1006 (O_1006,N_9431,N_9821);
and UO_1007 (O_1007,N_9021,N_9744);
nor UO_1008 (O_1008,N_9964,N_9557);
and UO_1009 (O_1009,N_9482,N_9067);
nand UO_1010 (O_1010,N_9847,N_9197);
nand UO_1011 (O_1011,N_9136,N_9650);
or UO_1012 (O_1012,N_9414,N_9904);
nor UO_1013 (O_1013,N_9875,N_9170);
nand UO_1014 (O_1014,N_9333,N_9861);
nor UO_1015 (O_1015,N_9099,N_9837);
nor UO_1016 (O_1016,N_9453,N_9407);
nor UO_1017 (O_1017,N_9224,N_9766);
or UO_1018 (O_1018,N_9824,N_9245);
and UO_1019 (O_1019,N_9272,N_9682);
nand UO_1020 (O_1020,N_9958,N_9258);
nor UO_1021 (O_1021,N_9223,N_9455);
and UO_1022 (O_1022,N_9948,N_9784);
and UO_1023 (O_1023,N_9238,N_9735);
and UO_1024 (O_1024,N_9433,N_9656);
and UO_1025 (O_1025,N_9907,N_9915);
or UO_1026 (O_1026,N_9725,N_9895);
or UO_1027 (O_1027,N_9347,N_9663);
or UO_1028 (O_1028,N_9494,N_9990);
and UO_1029 (O_1029,N_9191,N_9825);
nor UO_1030 (O_1030,N_9632,N_9961);
nor UO_1031 (O_1031,N_9635,N_9396);
or UO_1032 (O_1032,N_9120,N_9803);
nand UO_1033 (O_1033,N_9072,N_9439);
nor UO_1034 (O_1034,N_9096,N_9603);
nor UO_1035 (O_1035,N_9088,N_9960);
or UO_1036 (O_1036,N_9028,N_9067);
nand UO_1037 (O_1037,N_9334,N_9394);
nor UO_1038 (O_1038,N_9132,N_9601);
nor UO_1039 (O_1039,N_9054,N_9393);
or UO_1040 (O_1040,N_9149,N_9937);
nand UO_1041 (O_1041,N_9663,N_9367);
or UO_1042 (O_1042,N_9283,N_9743);
and UO_1043 (O_1043,N_9022,N_9608);
nor UO_1044 (O_1044,N_9924,N_9870);
and UO_1045 (O_1045,N_9479,N_9466);
and UO_1046 (O_1046,N_9208,N_9702);
nor UO_1047 (O_1047,N_9059,N_9817);
nor UO_1048 (O_1048,N_9872,N_9995);
and UO_1049 (O_1049,N_9018,N_9047);
or UO_1050 (O_1050,N_9943,N_9072);
or UO_1051 (O_1051,N_9163,N_9239);
and UO_1052 (O_1052,N_9444,N_9303);
nand UO_1053 (O_1053,N_9339,N_9316);
and UO_1054 (O_1054,N_9904,N_9254);
and UO_1055 (O_1055,N_9718,N_9019);
nor UO_1056 (O_1056,N_9909,N_9962);
and UO_1057 (O_1057,N_9749,N_9636);
or UO_1058 (O_1058,N_9515,N_9958);
or UO_1059 (O_1059,N_9760,N_9912);
or UO_1060 (O_1060,N_9765,N_9216);
nor UO_1061 (O_1061,N_9784,N_9120);
nor UO_1062 (O_1062,N_9089,N_9898);
nor UO_1063 (O_1063,N_9350,N_9513);
or UO_1064 (O_1064,N_9443,N_9837);
and UO_1065 (O_1065,N_9209,N_9852);
and UO_1066 (O_1066,N_9664,N_9518);
and UO_1067 (O_1067,N_9802,N_9778);
nand UO_1068 (O_1068,N_9386,N_9567);
xor UO_1069 (O_1069,N_9440,N_9809);
nand UO_1070 (O_1070,N_9810,N_9561);
nand UO_1071 (O_1071,N_9186,N_9429);
or UO_1072 (O_1072,N_9664,N_9245);
and UO_1073 (O_1073,N_9616,N_9911);
nand UO_1074 (O_1074,N_9547,N_9347);
nand UO_1075 (O_1075,N_9979,N_9380);
and UO_1076 (O_1076,N_9473,N_9399);
nor UO_1077 (O_1077,N_9512,N_9854);
nor UO_1078 (O_1078,N_9650,N_9531);
and UO_1079 (O_1079,N_9021,N_9446);
nor UO_1080 (O_1080,N_9784,N_9012);
nor UO_1081 (O_1081,N_9396,N_9657);
nor UO_1082 (O_1082,N_9111,N_9768);
and UO_1083 (O_1083,N_9624,N_9931);
nor UO_1084 (O_1084,N_9004,N_9825);
and UO_1085 (O_1085,N_9597,N_9160);
or UO_1086 (O_1086,N_9620,N_9967);
and UO_1087 (O_1087,N_9643,N_9383);
nand UO_1088 (O_1088,N_9650,N_9546);
or UO_1089 (O_1089,N_9524,N_9027);
or UO_1090 (O_1090,N_9751,N_9526);
and UO_1091 (O_1091,N_9817,N_9510);
and UO_1092 (O_1092,N_9072,N_9829);
nor UO_1093 (O_1093,N_9566,N_9730);
nand UO_1094 (O_1094,N_9461,N_9319);
and UO_1095 (O_1095,N_9055,N_9974);
nor UO_1096 (O_1096,N_9447,N_9966);
nand UO_1097 (O_1097,N_9272,N_9950);
nand UO_1098 (O_1098,N_9284,N_9189);
and UO_1099 (O_1099,N_9186,N_9520);
or UO_1100 (O_1100,N_9276,N_9647);
and UO_1101 (O_1101,N_9848,N_9514);
nand UO_1102 (O_1102,N_9845,N_9433);
or UO_1103 (O_1103,N_9480,N_9899);
nand UO_1104 (O_1104,N_9157,N_9048);
nor UO_1105 (O_1105,N_9604,N_9219);
nor UO_1106 (O_1106,N_9711,N_9383);
nand UO_1107 (O_1107,N_9435,N_9022);
or UO_1108 (O_1108,N_9729,N_9933);
or UO_1109 (O_1109,N_9236,N_9631);
or UO_1110 (O_1110,N_9695,N_9010);
and UO_1111 (O_1111,N_9092,N_9230);
nand UO_1112 (O_1112,N_9279,N_9365);
or UO_1113 (O_1113,N_9563,N_9459);
and UO_1114 (O_1114,N_9128,N_9477);
or UO_1115 (O_1115,N_9750,N_9561);
and UO_1116 (O_1116,N_9141,N_9245);
nand UO_1117 (O_1117,N_9570,N_9700);
nor UO_1118 (O_1118,N_9953,N_9554);
nand UO_1119 (O_1119,N_9731,N_9406);
nor UO_1120 (O_1120,N_9520,N_9909);
nor UO_1121 (O_1121,N_9261,N_9458);
and UO_1122 (O_1122,N_9197,N_9422);
nand UO_1123 (O_1123,N_9323,N_9914);
nand UO_1124 (O_1124,N_9299,N_9223);
and UO_1125 (O_1125,N_9156,N_9308);
and UO_1126 (O_1126,N_9372,N_9235);
nand UO_1127 (O_1127,N_9559,N_9369);
and UO_1128 (O_1128,N_9023,N_9248);
or UO_1129 (O_1129,N_9786,N_9921);
or UO_1130 (O_1130,N_9650,N_9346);
nor UO_1131 (O_1131,N_9794,N_9614);
nor UO_1132 (O_1132,N_9269,N_9000);
nor UO_1133 (O_1133,N_9174,N_9116);
nand UO_1134 (O_1134,N_9010,N_9168);
and UO_1135 (O_1135,N_9524,N_9882);
and UO_1136 (O_1136,N_9080,N_9305);
nor UO_1137 (O_1137,N_9151,N_9411);
or UO_1138 (O_1138,N_9477,N_9451);
or UO_1139 (O_1139,N_9380,N_9138);
nand UO_1140 (O_1140,N_9356,N_9590);
or UO_1141 (O_1141,N_9787,N_9546);
or UO_1142 (O_1142,N_9986,N_9194);
nand UO_1143 (O_1143,N_9399,N_9757);
nor UO_1144 (O_1144,N_9344,N_9404);
and UO_1145 (O_1145,N_9000,N_9170);
and UO_1146 (O_1146,N_9557,N_9261);
nand UO_1147 (O_1147,N_9148,N_9034);
or UO_1148 (O_1148,N_9838,N_9559);
and UO_1149 (O_1149,N_9029,N_9495);
or UO_1150 (O_1150,N_9385,N_9387);
and UO_1151 (O_1151,N_9902,N_9212);
and UO_1152 (O_1152,N_9151,N_9536);
nor UO_1153 (O_1153,N_9549,N_9127);
nor UO_1154 (O_1154,N_9786,N_9866);
or UO_1155 (O_1155,N_9194,N_9391);
nor UO_1156 (O_1156,N_9321,N_9700);
nand UO_1157 (O_1157,N_9544,N_9957);
nor UO_1158 (O_1158,N_9834,N_9986);
nor UO_1159 (O_1159,N_9069,N_9080);
and UO_1160 (O_1160,N_9607,N_9847);
and UO_1161 (O_1161,N_9597,N_9379);
and UO_1162 (O_1162,N_9673,N_9341);
and UO_1163 (O_1163,N_9563,N_9395);
nand UO_1164 (O_1164,N_9818,N_9736);
nand UO_1165 (O_1165,N_9448,N_9692);
nor UO_1166 (O_1166,N_9028,N_9437);
nand UO_1167 (O_1167,N_9507,N_9323);
and UO_1168 (O_1168,N_9006,N_9908);
or UO_1169 (O_1169,N_9863,N_9765);
nor UO_1170 (O_1170,N_9170,N_9677);
nor UO_1171 (O_1171,N_9184,N_9065);
and UO_1172 (O_1172,N_9849,N_9093);
nand UO_1173 (O_1173,N_9819,N_9571);
nand UO_1174 (O_1174,N_9948,N_9171);
nand UO_1175 (O_1175,N_9984,N_9978);
nor UO_1176 (O_1176,N_9541,N_9887);
and UO_1177 (O_1177,N_9348,N_9362);
and UO_1178 (O_1178,N_9538,N_9479);
or UO_1179 (O_1179,N_9375,N_9907);
nor UO_1180 (O_1180,N_9186,N_9857);
nand UO_1181 (O_1181,N_9154,N_9536);
nand UO_1182 (O_1182,N_9240,N_9835);
or UO_1183 (O_1183,N_9964,N_9457);
nand UO_1184 (O_1184,N_9716,N_9296);
nand UO_1185 (O_1185,N_9319,N_9006);
nor UO_1186 (O_1186,N_9614,N_9955);
or UO_1187 (O_1187,N_9588,N_9585);
or UO_1188 (O_1188,N_9442,N_9761);
nor UO_1189 (O_1189,N_9805,N_9342);
nor UO_1190 (O_1190,N_9843,N_9936);
or UO_1191 (O_1191,N_9256,N_9769);
or UO_1192 (O_1192,N_9879,N_9035);
or UO_1193 (O_1193,N_9996,N_9653);
and UO_1194 (O_1194,N_9870,N_9381);
and UO_1195 (O_1195,N_9011,N_9086);
or UO_1196 (O_1196,N_9814,N_9957);
or UO_1197 (O_1197,N_9761,N_9931);
and UO_1198 (O_1198,N_9080,N_9456);
nor UO_1199 (O_1199,N_9309,N_9755);
nor UO_1200 (O_1200,N_9262,N_9081);
nand UO_1201 (O_1201,N_9588,N_9967);
nor UO_1202 (O_1202,N_9960,N_9350);
and UO_1203 (O_1203,N_9779,N_9131);
and UO_1204 (O_1204,N_9212,N_9645);
or UO_1205 (O_1205,N_9608,N_9467);
nor UO_1206 (O_1206,N_9290,N_9827);
nand UO_1207 (O_1207,N_9720,N_9839);
nand UO_1208 (O_1208,N_9396,N_9841);
and UO_1209 (O_1209,N_9350,N_9434);
and UO_1210 (O_1210,N_9854,N_9327);
or UO_1211 (O_1211,N_9465,N_9973);
and UO_1212 (O_1212,N_9044,N_9522);
nand UO_1213 (O_1213,N_9741,N_9004);
nand UO_1214 (O_1214,N_9667,N_9366);
and UO_1215 (O_1215,N_9177,N_9358);
and UO_1216 (O_1216,N_9944,N_9706);
nand UO_1217 (O_1217,N_9009,N_9396);
or UO_1218 (O_1218,N_9071,N_9613);
nor UO_1219 (O_1219,N_9281,N_9914);
and UO_1220 (O_1220,N_9107,N_9874);
nand UO_1221 (O_1221,N_9199,N_9745);
nor UO_1222 (O_1222,N_9611,N_9124);
nor UO_1223 (O_1223,N_9879,N_9958);
nand UO_1224 (O_1224,N_9235,N_9834);
nor UO_1225 (O_1225,N_9069,N_9707);
or UO_1226 (O_1226,N_9947,N_9138);
and UO_1227 (O_1227,N_9694,N_9233);
and UO_1228 (O_1228,N_9733,N_9506);
nor UO_1229 (O_1229,N_9263,N_9342);
or UO_1230 (O_1230,N_9408,N_9578);
nand UO_1231 (O_1231,N_9972,N_9919);
or UO_1232 (O_1232,N_9402,N_9056);
nand UO_1233 (O_1233,N_9447,N_9387);
nand UO_1234 (O_1234,N_9819,N_9943);
nor UO_1235 (O_1235,N_9527,N_9160);
nand UO_1236 (O_1236,N_9688,N_9868);
and UO_1237 (O_1237,N_9213,N_9304);
nor UO_1238 (O_1238,N_9716,N_9852);
nor UO_1239 (O_1239,N_9525,N_9364);
nand UO_1240 (O_1240,N_9801,N_9690);
or UO_1241 (O_1241,N_9953,N_9087);
and UO_1242 (O_1242,N_9711,N_9939);
and UO_1243 (O_1243,N_9381,N_9224);
or UO_1244 (O_1244,N_9326,N_9443);
nand UO_1245 (O_1245,N_9818,N_9046);
and UO_1246 (O_1246,N_9841,N_9676);
nor UO_1247 (O_1247,N_9205,N_9482);
or UO_1248 (O_1248,N_9402,N_9734);
and UO_1249 (O_1249,N_9073,N_9455);
nor UO_1250 (O_1250,N_9854,N_9304);
nor UO_1251 (O_1251,N_9833,N_9699);
or UO_1252 (O_1252,N_9452,N_9894);
or UO_1253 (O_1253,N_9945,N_9841);
nor UO_1254 (O_1254,N_9942,N_9950);
or UO_1255 (O_1255,N_9020,N_9825);
nor UO_1256 (O_1256,N_9411,N_9223);
or UO_1257 (O_1257,N_9222,N_9760);
nand UO_1258 (O_1258,N_9184,N_9515);
nand UO_1259 (O_1259,N_9821,N_9799);
nand UO_1260 (O_1260,N_9644,N_9211);
or UO_1261 (O_1261,N_9977,N_9765);
nand UO_1262 (O_1262,N_9134,N_9858);
or UO_1263 (O_1263,N_9833,N_9832);
nor UO_1264 (O_1264,N_9025,N_9747);
or UO_1265 (O_1265,N_9093,N_9198);
nand UO_1266 (O_1266,N_9220,N_9923);
nor UO_1267 (O_1267,N_9894,N_9604);
or UO_1268 (O_1268,N_9734,N_9682);
nand UO_1269 (O_1269,N_9589,N_9364);
and UO_1270 (O_1270,N_9274,N_9222);
nor UO_1271 (O_1271,N_9310,N_9688);
nor UO_1272 (O_1272,N_9594,N_9331);
nand UO_1273 (O_1273,N_9442,N_9990);
nor UO_1274 (O_1274,N_9439,N_9241);
or UO_1275 (O_1275,N_9835,N_9703);
or UO_1276 (O_1276,N_9449,N_9171);
nand UO_1277 (O_1277,N_9690,N_9209);
and UO_1278 (O_1278,N_9517,N_9396);
nand UO_1279 (O_1279,N_9571,N_9840);
or UO_1280 (O_1280,N_9007,N_9098);
nand UO_1281 (O_1281,N_9903,N_9166);
nor UO_1282 (O_1282,N_9017,N_9012);
or UO_1283 (O_1283,N_9591,N_9019);
nand UO_1284 (O_1284,N_9403,N_9118);
and UO_1285 (O_1285,N_9390,N_9168);
and UO_1286 (O_1286,N_9477,N_9355);
nand UO_1287 (O_1287,N_9546,N_9235);
nor UO_1288 (O_1288,N_9339,N_9405);
and UO_1289 (O_1289,N_9666,N_9150);
and UO_1290 (O_1290,N_9151,N_9352);
nand UO_1291 (O_1291,N_9277,N_9547);
nor UO_1292 (O_1292,N_9693,N_9533);
nor UO_1293 (O_1293,N_9104,N_9505);
and UO_1294 (O_1294,N_9895,N_9465);
nand UO_1295 (O_1295,N_9546,N_9318);
nor UO_1296 (O_1296,N_9078,N_9842);
nor UO_1297 (O_1297,N_9608,N_9300);
xor UO_1298 (O_1298,N_9366,N_9147);
nand UO_1299 (O_1299,N_9405,N_9332);
nand UO_1300 (O_1300,N_9658,N_9113);
and UO_1301 (O_1301,N_9335,N_9423);
nor UO_1302 (O_1302,N_9800,N_9835);
nand UO_1303 (O_1303,N_9677,N_9472);
nand UO_1304 (O_1304,N_9905,N_9351);
or UO_1305 (O_1305,N_9857,N_9441);
nand UO_1306 (O_1306,N_9783,N_9710);
nor UO_1307 (O_1307,N_9449,N_9718);
nand UO_1308 (O_1308,N_9565,N_9888);
nor UO_1309 (O_1309,N_9262,N_9783);
and UO_1310 (O_1310,N_9986,N_9488);
and UO_1311 (O_1311,N_9197,N_9285);
and UO_1312 (O_1312,N_9699,N_9223);
or UO_1313 (O_1313,N_9847,N_9791);
and UO_1314 (O_1314,N_9587,N_9963);
nand UO_1315 (O_1315,N_9222,N_9875);
nand UO_1316 (O_1316,N_9980,N_9519);
nand UO_1317 (O_1317,N_9550,N_9303);
nor UO_1318 (O_1318,N_9321,N_9571);
nand UO_1319 (O_1319,N_9896,N_9924);
and UO_1320 (O_1320,N_9506,N_9422);
nor UO_1321 (O_1321,N_9482,N_9245);
and UO_1322 (O_1322,N_9233,N_9598);
nor UO_1323 (O_1323,N_9863,N_9356);
or UO_1324 (O_1324,N_9984,N_9505);
or UO_1325 (O_1325,N_9708,N_9281);
or UO_1326 (O_1326,N_9529,N_9189);
or UO_1327 (O_1327,N_9658,N_9451);
nor UO_1328 (O_1328,N_9628,N_9728);
xnor UO_1329 (O_1329,N_9258,N_9489);
and UO_1330 (O_1330,N_9301,N_9056);
or UO_1331 (O_1331,N_9712,N_9271);
nor UO_1332 (O_1332,N_9718,N_9162);
nor UO_1333 (O_1333,N_9165,N_9519);
nor UO_1334 (O_1334,N_9047,N_9759);
or UO_1335 (O_1335,N_9210,N_9743);
nor UO_1336 (O_1336,N_9366,N_9581);
nand UO_1337 (O_1337,N_9405,N_9862);
and UO_1338 (O_1338,N_9808,N_9915);
or UO_1339 (O_1339,N_9022,N_9978);
nand UO_1340 (O_1340,N_9535,N_9824);
nand UO_1341 (O_1341,N_9796,N_9472);
nand UO_1342 (O_1342,N_9157,N_9850);
and UO_1343 (O_1343,N_9374,N_9020);
nor UO_1344 (O_1344,N_9713,N_9445);
and UO_1345 (O_1345,N_9091,N_9523);
and UO_1346 (O_1346,N_9529,N_9946);
or UO_1347 (O_1347,N_9827,N_9179);
or UO_1348 (O_1348,N_9186,N_9761);
nand UO_1349 (O_1349,N_9376,N_9096);
nor UO_1350 (O_1350,N_9909,N_9101);
or UO_1351 (O_1351,N_9512,N_9184);
nand UO_1352 (O_1352,N_9764,N_9247);
nand UO_1353 (O_1353,N_9375,N_9578);
or UO_1354 (O_1354,N_9788,N_9476);
nor UO_1355 (O_1355,N_9707,N_9744);
and UO_1356 (O_1356,N_9254,N_9315);
and UO_1357 (O_1357,N_9692,N_9362);
or UO_1358 (O_1358,N_9765,N_9956);
and UO_1359 (O_1359,N_9838,N_9920);
nor UO_1360 (O_1360,N_9845,N_9329);
nor UO_1361 (O_1361,N_9215,N_9164);
nor UO_1362 (O_1362,N_9872,N_9619);
nor UO_1363 (O_1363,N_9502,N_9217);
or UO_1364 (O_1364,N_9207,N_9477);
nor UO_1365 (O_1365,N_9428,N_9005);
nand UO_1366 (O_1366,N_9851,N_9110);
and UO_1367 (O_1367,N_9521,N_9317);
or UO_1368 (O_1368,N_9742,N_9474);
nand UO_1369 (O_1369,N_9934,N_9490);
nand UO_1370 (O_1370,N_9460,N_9532);
nand UO_1371 (O_1371,N_9040,N_9474);
nor UO_1372 (O_1372,N_9992,N_9195);
nor UO_1373 (O_1373,N_9778,N_9115);
nor UO_1374 (O_1374,N_9051,N_9429);
nand UO_1375 (O_1375,N_9697,N_9266);
nand UO_1376 (O_1376,N_9324,N_9383);
or UO_1377 (O_1377,N_9666,N_9938);
or UO_1378 (O_1378,N_9891,N_9395);
nand UO_1379 (O_1379,N_9412,N_9463);
nor UO_1380 (O_1380,N_9910,N_9895);
nand UO_1381 (O_1381,N_9329,N_9887);
or UO_1382 (O_1382,N_9220,N_9083);
and UO_1383 (O_1383,N_9743,N_9226);
and UO_1384 (O_1384,N_9974,N_9857);
and UO_1385 (O_1385,N_9652,N_9110);
and UO_1386 (O_1386,N_9683,N_9724);
nand UO_1387 (O_1387,N_9406,N_9322);
nor UO_1388 (O_1388,N_9849,N_9879);
nand UO_1389 (O_1389,N_9707,N_9633);
nor UO_1390 (O_1390,N_9073,N_9957);
nor UO_1391 (O_1391,N_9979,N_9463);
and UO_1392 (O_1392,N_9881,N_9577);
nor UO_1393 (O_1393,N_9382,N_9323);
or UO_1394 (O_1394,N_9896,N_9866);
nor UO_1395 (O_1395,N_9458,N_9590);
nand UO_1396 (O_1396,N_9207,N_9715);
or UO_1397 (O_1397,N_9963,N_9299);
nor UO_1398 (O_1398,N_9019,N_9558);
and UO_1399 (O_1399,N_9040,N_9434);
nor UO_1400 (O_1400,N_9371,N_9252);
and UO_1401 (O_1401,N_9202,N_9899);
nor UO_1402 (O_1402,N_9429,N_9304);
nand UO_1403 (O_1403,N_9796,N_9176);
nor UO_1404 (O_1404,N_9589,N_9448);
nor UO_1405 (O_1405,N_9126,N_9617);
and UO_1406 (O_1406,N_9866,N_9429);
nor UO_1407 (O_1407,N_9704,N_9759);
nand UO_1408 (O_1408,N_9359,N_9063);
and UO_1409 (O_1409,N_9399,N_9437);
or UO_1410 (O_1410,N_9915,N_9135);
and UO_1411 (O_1411,N_9477,N_9093);
and UO_1412 (O_1412,N_9242,N_9713);
nor UO_1413 (O_1413,N_9367,N_9833);
nor UO_1414 (O_1414,N_9954,N_9139);
nor UO_1415 (O_1415,N_9477,N_9247);
and UO_1416 (O_1416,N_9027,N_9091);
and UO_1417 (O_1417,N_9057,N_9357);
nor UO_1418 (O_1418,N_9822,N_9212);
nor UO_1419 (O_1419,N_9024,N_9695);
and UO_1420 (O_1420,N_9979,N_9538);
nor UO_1421 (O_1421,N_9967,N_9345);
and UO_1422 (O_1422,N_9439,N_9976);
or UO_1423 (O_1423,N_9492,N_9107);
or UO_1424 (O_1424,N_9577,N_9974);
nand UO_1425 (O_1425,N_9972,N_9724);
nor UO_1426 (O_1426,N_9869,N_9378);
and UO_1427 (O_1427,N_9835,N_9420);
xor UO_1428 (O_1428,N_9741,N_9726);
and UO_1429 (O_1429,N_9332,N_9908);
nor UO_1430 (O_1430,N_9211,N_9911);
or UO_1431 (O_1431,N_9617,N_9840);
or UO_1432 (O_1432,N_9831,N_9862);
or UO_1433 (O_1433,N_9943,N_9048);
nor UO_1434 (O_1434,N_9062,N_9487);
or UO_1435 (O_1435,N_9074,N_9324);
nor UO_1436 (O_1436,N_9334,N_9714);
nand UO_1437 (O_1437,N_9178,N_9655);
nand UO_1438 (O_1438,N_9430,N_9152);
nand UO_1439 (O_1439,N_9286,N_9226);
and UO_1440 (O_1440,N_9197,N_9449);
nor UO_1441 (O_1441,N_9590,N_9271);
or UO_1442 (O_1442,N_9979,N_9191);
and UO_1443 (O_1443,N_9447,N_9244);
and UO_1444 (O_1444,N_9463,N_9577);
nor UO_1445 (O_1445,N_9270,N_9640);
and UO_1446 (O_1446,N_9756,N_9057);
nand UO_1447 (O_1447,N_9293,N_9193);
and UO_1448 (O_1448,N_9153,N_9038);
nand UO_1449 (O_1449,N_9334,N_9059);
and UO_1450 (O_1450,N_9769,N_9713);
or UO_1451 (O_1451,N_9271,N_9787);
or UO_1452 (O_1452,N_9739,N_9879);
nor UO_1453 (O_1453,N_9048,N_9580);
and UO_1454 (O_1454,N_9344,N_9603);
or UO_1455 (O_1455,N_9201,N_9206);
and UO_1456 (O_1456,N_9085,N_9793);
nor UO_1457 (O_1457,N_9369,N_9575);
nor UO_1458 (O_1458,N_9869,N_9964);
or UO_1459 (O_1459,N_9648,N_9211);
or UO_1460 (O_1460,N_9772,N_9014);
nor UO_1461 (O_1461,N_9472,N_9660);
and UO_1462 (O_1462,N_9195,N_9217);
or UO_1463 (O_1463,N_9734,N_9203);
xor UO_1464 (O_1464,N_9640,N_9621);
or UO_1465 (O_1465,N_9064,N_9458);
and UO_1466 (O_1466,N_9342,N_9705);
nor UO_1467 (O_1467,N_9700,N_9722);
and UO_1468 (O_1468,N_9575,N_9283);
nor UO_1469 (O_1469,N_9231,N_9854);
xnor UO_1470 (O_1470,N_9969,N_9571);
or UO_1471 (O_1471,N_9841,N_9493);
nand UO_1472 (O_1472,N_9006,N_9397);
nor UO_1473 (O_1473,N_9959,N_9759);
and UO_1474 (O_1474,N_9196,N_9791);
or UO_1475 (O_1475,N_9624,N_9033);
nand UO_1476 (O_1476,N_9429,N_9817);
nor UO_1477 (O_1477,N_9970,N_9568);
nand UO_1478 (O_1478,N_9342,N_9445);
nand UO_1479 (O_1479,N_9221,N_9661);
and UO_1480 (O_1480,N_9018,N_9900);
nor UO_1481 (O_1481,N_9721,N_9547);
nor UO_1482 (O_1482,N_9849,N_9746);
nor UO_1483 (O_1483,N_9824,N_9609);
and UO_1484 (O_1484,N_9330,N_9104);
or UO_1485 (O_1485,N_9047,N_9704);
nor UO_1486 (O_1486,N_9026,N_9805);
or UO_1487 (O_1487,N_9778,N_9723);
or UO_1488 (O_1488,N_9266,N_9522);
nand UO_1489 (O_1489,N_9669,N_9370);
and UO_1490 (O_1490,N_9953,N_9413);
nand UO_1491 (O_1491,N_9944,N_9471);
nor UO_1492 (O_1492,N_9942,N_9422);
nand UO_1493 (O_1493,N_9107,N_9715);
and UO_1494 (O_1494,N_9051,N_9762);
nand UO_1495 (O_1495,N_9373,N_9293);
nand UO_1496 (O_1496,N_9670,N_9552);
and UO_1497 (O_1497,N_9190,N_9288);
nand UO_1498 (O_1498,N_9826,N_9150);
or UO_1499 (O_1499,N_9088,N_9617);
endmodule