module basic_1000_10000_1500_20_levels_2xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_711,In_880);
nand U1 (N_1,In_616,In_83);
nor U2 (N_2,In_434,In_498);
and U3 (N_3,In_984,In_840);
nand U4 (N_4,In_604,In_558);
and U5 (N_5,In_933,In_583);
or U6 (N_6,In_223,In_447);
and U7 (N_7,In_72,In_160);
nor U8 (N_8,In_932,In_352);
nor U9 (N_9,In_980,In_140);
and U10 (N_10,In_955,In_235);
or U11 (N_11,In_582,In_445);
nor U12 (N_12,In_326,In_358);
and U13 (N_13,In_146,In_284);
nor U14 (N_14,In_674,In_309);
nor U15 (N_15,In_5,In_288);
or U16 (N_16,In_972,In_945);
or U17 (N_17,In_49,In_580);
nand U18 (N_18,In_772,In_383);
or U19 (N_19,In_148,In_988);
and U20 (N_20,In_666,In_131);
nor U21 (N_21,In_490,In_466);
nor U22 (N_22,In_813,In_561);
nand U23 (N_23,In_322,In_659);
and U24 (N_24,In_225,In_707);
nand U25 (N_25,In_397,In_970);
or U26 (N_26,In_172,In_748);
and U27 (N_27,In_563,In_540);
nand U28 (N_28,In_479,In_536);
and U29 (N_29,In_66,In_30);
and U30 (N_30,In_423,In_306);
nand U31 (N_31,In_474,In_15);
nand U32 (N_32,In_769,In_862);
or U33 (N_33,In_814,In_570);
nor U34 (N_34,In_873,In_915);
or U35 (N_35,In_496,In_145);
nor U36 (N_36,In_463,In_168);
or U37 (N_37,In_400,In_133);
and U38 (N_38,In_559,In_130);
nor U39 (N_39,In_251,In_670);
nor U40 (N_40,In_820,In_743);
or U41 (N_41,In_230,In_893);
nor U42 (N_42,In_657,In_13);
nand U43 (N_43,In_105,In_281);
nand U44 (N_44,In_176,In_387);
nand U45 (N_45,In_506,In_6);
nand U46 (N_46,In_40,In_449);
nor U47 (N_47,In_417,In_297);
or U48 (N_48,In_751,In_854);
and U49 (N_49,In_804,In_994);
nand U50 (N_50,In_904,In_931);
or U51 (N_51,In_294,In_695);
or U52 (N_52,In_499,In_33);
and U53 (N_53,In_468,In_224);
and U54 (N_54,In_716,In_938);
and U55 (N_55,In_418,In_596);
or U56 (N_56,In_909,In_696);
nor U57 (N_57,In_245,In_532);
or U58 (N_58,In_649,In_942);
nand U59 (N_59,In_113,In_422);
or U60 (N_60,In_234,In_683);
nor U61 (N_61,In_947,In_275);
nand U62 (N_62,In_855,In_754);
nor U63 (N_63,In_812,In_43);
nor U64 (N_64,In_848,In_76);
xor U65 (N_65,In_411,In_246);
nor U66 (N_66,In_29,In_51);
or U67 (N_67,In_412,In_555);
nand U68 (N_68,In_456,In_719);
nor U69 (N_69,In_872,In_469);
nor U70 (N_70,In_316,In_512);
and U71 (N_71,In_776,In_180);
and U72 (N_72,In_109,In_263);
or U73 (N_73,In_860,In_591);
nor U74 (N_74,In_557,In_23);
nor U75 (N_75,In_857,In_442);
and U76 (N_76,In_686,In_92);
nor U77 (N_77,In_876,In_375);
nand U78 (N_78,In_733,In_356);
or U79 (N_79,In_808,In_757);
nor U80 (N_80,In_597,In_635);
nand U81 (N_81,In_386,In_321);
or U82 (N_82,In_729,In_702);
and U83 (N_83,In_210,In_953);
nand U84 (N_84,In_828,In_233);
nand U85 (N_85,In_727,In_773);
or U86 (N_86,In_486,In_287);
nand U87 (N_87,In_344,In_504);
nor U88 (N_88,In_925,In_421);
xor U89 (N_89,In_749,In_671);
nand U90 (N_90,In_553,In_487);
and U91 (N_91,In_542,In_771);
nand U92 (N_92,In_88,In_12);
nor U93 (N_93,In_983,In_373);
or U94 (N_94,In_443,In_259);
nor U95 (N_95,In_81,In_471);
and U96 (N_96,In_77,In_170);
and U97 (N_97,In_775,In_328);
nand U98 (N_98,In_856,In_903);
nand U99 (N_99,In_357,In_999);
or U100 (N_100,In_107,In_950);
or U101 (N_101,In_85,In_547);
and U102 (N_102,In_985,In_746);
and U103 (N_103,In_200,In_80);
or U104 (N_104,In_850,In_493);
nor U105 (N_105,In_936,In_835);
or U106 (N_106,In_91,In_323);
nand U107 (N_107,In_120,In_53);
and U108 (N_108,In_761,In_630);
nand U109 (N_109,In_98,In_788);
nor U110 (N_110,In_193,In_965);
nand U111 (N_111,In_615,In_261);
and U112 (N_112,In_881,In_18);
or U113 (N_113,In_207,In_292);
nand U114 (N_114,In_52,In_150);
or U115 (N_115,In_467,In_827);
or U116 (N_116,In_178,In_710);
nand U117 (N_117,In_361,In_668);
or U118 (N_118,In_681,In_173);
nor U119 (N_119,In_731,In_943);
nand U120 (N_120,In_723,In_930);
nand U121 (N_121,In_560,In_637);
and U122 (N_122,In_747,In_189);
or U123 (N_123,In_502,In_908);
nand U124 (N_124,In_527,In_651);
and U125 (N_125,In_278,In_825);
or U126 (N_126,In_379,In_673);
and U127 (N_127,In_58,In_16);
or U128 (N_128,In_161,In_260);
nor U129 (N_129,In_897,In_157);
nor U130 (N_130,In_481,In_521);
nor U131 (N_131,In_394,In_509);
nor U132 (N_132,In_73,In_97);
nand U133 (N_133,In_156,In_432);
and U134 (N_134,In_894,In_162);
and U135 (N_135,In_822,In_530);
or U136 (N_136,In_78,In_703);
or U137 (N_137,In_138,In_482);
and U138 (N_138,In_114,In_992);
nand U139 (N_139,In_842,In_214);
and U140 (N_140,In_354,In_304);
nand U141 (N_141,In_44,In_662);
and U142 (N_142,In_913,In_313);
xor U143 (N_143,In_149,In_778);
or U144 (N_144,In_353,In_401);
or U145 (N_145,In_998,In_462);
nor U146 (N_146,In_899,In_128);
nand U147 (N_147,In_895,In_69);
nor U148 (N_148,In_414,In_520);
and U149 (N_149,In_198,In_971);
or U150 (N_150,In_902,In_265);
nand U151 (N_151,In_295,In_568);
or U152 (N_152,In_376,In_704);
or U153 (N_153,In_937,In_519);
nor U154 (N_154,In_510,In_905);
nor U155 (N_155,In_575,In_917);
and U156 (N_156,In_679,In_99);
xor U157 (N_157,In_779,In_111);
and U158 (N_158,In_650,In_231);
and U159 (N_159,In_185,In_717);
nand U160 (N_160,In_874,In_351);
nor U161 (N_161,In_766,In_41);
xor U162 (N_162,In_55,In_632);
or U163 (N_163,In_979,In_392);
or U164 (N_164,In_991,In_851);
or U165 (N_165,In_452,In_8);
nor U166 (N_166,In_868,In_366);
nand U167 (N_167,In_664,In_964);
nand U168 (N_168,In_426,In_839);
or U169 (N_169,In_692,In_218);
or U170 (N_170,In_222,In_378);
or U171 (N_171,In_959,In_312);
and U172 (N_172,In_305,In_330);
nand U173 (N_173,In_941,In_640);
and U174 (N_174,In_694,In_255);
or U175 (N_175,In_182,In_884);
and U176 (N_176,In_45,In_684);
nand U177 (N_177,In_291,In_550);
and U178 (N_178,In_405,In_619);
and U179 (N_179,In_319,In_203);
or U180 (N_180,In_672,In_177);
and U181 (N_181,In_514,In_934);
or U182 (N_182,In_333,In_262);
nand U183 (N_183,In_789,In_602);
and U184 (N_184,In_861,In_617);
and U185 (N_185,In_923,In_551);
and U186 (N_186,In_477,In_976);
nor U187 (N_187,In_25,In_987);
or U188 (N_188,In_508,In_57);
or U189 (N_189,In_537,In_237);
nor U190 (N_190,In_996,In_989);
or U191 (N_191,In_35,In_787);
nand U192 (N_192,In_623,In_795);
nor U193 (N_193,In_712,In_646);
and U194 (N_194,In_564,In_365);
nor U195 (N_195,In_566,In_753);
or U196 (N_196,In_541,In_974);
and U197 (N_197,In_533,In_726);
nand U198 (N_198,In_398,In_791);
nor U199 (N_199,In_183,In_781);
nor U200 (N_200,In_380,In_293);
and U201 (N_201,In_495,In_194);
nor U202 (N_202,In_982,In_737);
nor U203 (N_203,In_458,In_377);
or U204 (N_204,In_382,In_491);
xor U205 (N_205,In_489,In_543);
nand U206 (N_206,In_949,In_720);
nand U207 (N_207,In_918,In_0);
nor U208 (N_208,In_658,In_75);
nor U209 (N_209,In_158,In_648);
nor U210 (N_210,In_28,In_192);
or U211 (N_211,In_800,In_634);
xor U212 (N_212,In_381,In_112);
nor U213 (N_213,In_317,In_141);
or U214 (N_214,In_732,In_954);
and U215 (N_215,In_2,In_137);
and U216 (N_216,In_79,In_308);
nand U217 (N_217,In_817,In_977);
and U218 (N_218,In_935,In_310);
and U219 (N_219,In_967,In_402);
nor U220 (N_220,In_699,In_132);
or U221 (N_221,In_724,In_71);
nor U222 (N_222,In_267,In_164);
or U223 (N_223,In_239,In_74);
or U224 (N_224,In_572,In_236);
xnor U225 (N_225,In_734,In_888);
or U226 (N_226,In_552,In_212);
nor U227 (N_227,In_687,In_348);
nand U228 (N_228,In_475,In_545);
and U229 (N_229,In_643,In_837);
nor U230 (N_230,In_957,In_363);
or U231 (N_231,In_494,In_359);
nor U232 (N_232,In_54,In_513);
nand U233 (N_233,In_253,In_863);
xor U234 (N_234,In_390,In_609);
nor U235 (N_235,In_129,In_593);
nor U236 (N_236,In_878,In_4);
or U237 (N_237,In_325,In_385);
nor U238 (N_238,In_393,In_735);
nand U239 (N_239,In_700,In_594);
nor U240 (N_240,In_782,In_592);
nand U241 (N_241,In_911,In_410);
and U242 (N_242,In_429,In_450);
nor U243 (N_243,In_1,In_206);
nand U244 (N_244,In_258,In_901);
nand U245 (N_245,In_832,In_388);
nand U246 (N_246,In_631,In_745);
xor U247 (N_247,In_14,In_315);
and U248 (N_248,In_415,In_143);
and U249 (N_249,In_755,In_836);
nand U250 (N_250,In_110,In_48);
nor U251 (N_251,In_829,In_229);
and U252 (N_252,In_618,In_473);
nand U253 (N_253,In_298,In_216);
or U254 (N_254,In_420,In_993);
or U255 (N_255,In_127,In_480);
or U256 (N_256,In_752,In_238);
nand U257 (N_257,In_436,In_562);
nor U258 (N_258,In_556,In_440);
and U259 (N_259,In_155,In_713);
nand U260 (N_260,In_497,In_303);
nand U261 (N_261,In_606,In_221);
nor U262 (N_262,In_360,In_774);
or U263 (N_263,In_730,In_535);
or U264 (N_264,In_685,In_603);
nand U265 (N_265,In_123,In_981);
nor U266 (N_266,In_846,In_197);
and U267 (N_267,In_264,In_20);
nand U268 (N_268,In_26,In_849);
or U269 (N_269,In_395,In_691);
or U270 (N_270,In_966,In_122);
nand U271 (N_271,In_929,In_944);
nand U272 (N_272,In_451,In_95);
nand U273 (N_273,In_756,In_518);
or U274 (N_274,In_907,In_86);
or U275 (N_275,In_100,In_341);
and U276 (N_276,In_830,In_384);
nand U277 (N_277,In_896,In_784);
nand U278 (N_278,In_84,In_34);
nor U279 (N_279,In_741,In_302);
or U280 (N_280,In_528,In_144);
and U281 (N_281,In_736,In_889);
or U282 (N_282,In_525,In_573);
and U283 (N_283,In_87,In_598);
nor U284 (N_284,In_777,In_995);
and U285 (N_285,In_94,In_318);
or U286 (N_286,In_910,In_10);
and U287 (N_287,In_522,In_147);
nand U288 (N_288,In_833,In_625);
nor U289 (N_289,In_60,In_369);
nor U290 (N_290,In_529,In_174);
nand U291 (N_291,In_589,In_346);
nor U292 (N_292,In_249,In_948);
or U293 (N_293,In_364,In_9);
and U294 (N_294,In_355,In_65);
nor U295 (N_295,In_3,In_399);
xor U296 (N_296,In_116,In_847);
or U297 (N_297,In_927,In_406);
nor U298 (N_298,In_920,In_990);
or U299 (N_299,In_652,In_136);
nor U300 (N_300,In_823,In_269);
and U301 (N_301,In_21,In_121);
nor U302 (N_302,In_644,In_581);
nor U303 (N_303,In_882,In_569);
nand U304 (N_304,In_476,In_454);
xnor U305 (N_305,In_254,In_424);
and U306 (N_306,In_534,In_419);
or U307 (N_307,In_343,In_19);
and U308 (N_308,In_952,In_963);
nand U309 (N_309,In_796,In_299);
nor U310 (N_310,In_311,In_142);
nor U311 (N_311,In_661,In_961);
nand U312 (N_312,In_571,In_916);
or U313 (N_313,In_653,In_892);
nor U314 (N_314,In_821,In_638);
or U315 (N_315,In_826,In_669);
and U316 (N_316,In_811,In_407);
or U317 (N_317,In_824,In_42);
or U318 (N_318,In_370,In_554);
nand U319 (N_319,In_750,In_336);
nand U320 (N_320,In_324,In_270);
nand U321 (N_321,In_960,In_912);
and U322 (N_322,In_331,In_362);
nor U323 (N_323,In_928,In_459);
or U324 (N_324,In_332,In_163);
and U325 (N_325,In_46,In_608);
nor U326 (N_326,In_578,In_134);
and U327 (N_327,In_574,In_204);
or U328 (N_328,In_119,In_645);
and U329 (N_329,In_226,In_431);
nor U330 (N_330,In_605,In_810);
or U331 (N_331,In_636,In_803);
nand U332 (N_332,In_831,In_539);
and U333 (N_333,In_389,In_647);
or U334 (N_334,In_61,In_63);
nand U335 (N_335,In_969,In_154);
nand U336 (N_336,In_588,In_629);
or U337 (N_337,In_864,In_838);
or U338 (N_338,In_866,In_867);
nor U339 (N_339,In_196,In_427);
nand U340 (N_340,In_641,In_108);
and U341 (N_341,In_654,In_472);
nor U342 (N_342,In_36,In_507);
and U343 (N_343,In_585,In_372);
or U344 (N_344,In_764,In_492);
and U345 (N_345,In_701,In_877);
or U346 (N_346,In_926,In_106);
or U347 (N_347,In_257,In_682);
or U348 (N_348,In_688,In_101);
or U349 (N_349,In_300,In_38);
nor U350 (N_350,In_601,In_549);
nor U351 (N_351,In_437,In_586);
nand U352 (N_352,In_806,In_279);
nand U353 (N_353,In_256,In_538);
nand U354 (N_354,In_900,In_760);
nand U355 (N_355,In_215,In_802);
and U356 (N_356,In_102,In_722);
and U357 (N_357,In_243,In_875);
nand U358 (N_358,In_633,In_62);
and U359 (N_359,In_289,In_922);
nand U360 (N_360,In_171,In_350);
nor U361 (N_361,In_272,In_962);
or U362 (N_362,In_416,In_767);
and U363 (N_363,In_501,In_188);
or U364 (N_364,In_577,In_448);
or U365 (N_365,In_798,In_600);
and U366 (N_366,In_655,In_816);
nor U367 (N_367,In_67,In_852);
and U368 (N_368,In_786,In_500);
nor U369 (N_369,In_792,In_186);
nor U370 (N_370,In_277,In_834);
or U371 (N_371,In_921,In_958);
nand U372 (N_372,In_347,In_391);
nor U373 (N_373,In_620,In_280);
nor U374 (N_374,In_339,In_978);
nor U375 (N_375,In_104,In_165);
nor U376 (N_376,In_622,In_470);
and U377 (N_377,In_587,In_709);
or U378 (N_378,In_898,In_511);
nand U379 (N_379,In_815,In_505);
xnor U380 (N_380,In_858,In_208);
nand U381 (N_381,In_125,In_329);
nand U382 (N_382,In_340,In_219);
and U383 (N_383,In_191,In_181);
nand U384 (N_384,In_24,In_624);
and U385 (N_385,In_17,In_408);
or U386 (N_386,In_166,In_296);
nand U387 (N_387,In_209,In_345);
nor U388 (N_388,In_956,In_153);
and U389 (N_389,In_190,In_22);
and U390 (N_390,In_349,In_268);
or U391 (N_391,In_217,In_282);
nand U392 (N_392,In_184,In_286);
and U393 (N_393,In_374,In_413);
or U394 (N_394,In_595,In_202);
or U395 (N_395,In_320,In_584);
nor U396 (N_396,In_783,In_517);
nor U397 (N_397,In_951,In_740);
nand U398 (N_398,In_59,In_516);
or U399 (N_399,In_338,In_56);
nand U400 (N_400,In_446,In_886);
nor U401 (N_401,In_973,In_244);
nand U402 (N_402,In_742,In_986);
or U403 (N_403,In_819,In_27);
nor U404 (N_404,In_285,In_887);
nand U405 (N_405,In_975,In_488);
nor U406 (N_406,In_367,In_579);
nand U407 (N_407,In_663,In_879);
and U408 (N_408,In_765,In_228);
nor U409 (N_409,In_453,In_461);
and U410 (N_410,In_118,In_396);
or U411 (N_411,In_871,In_247);
and U412 (N_412,In_807,In_68);
nand U413 (N_413,In_211,In_460);
and U414 (N_414,In_438,In_763);
nand U415 (N_415,In_37,In_744);
nor U416 (N_416,In_768,In_232);
and U417 (N_417,In_327,In_152);
and U418 (N_418,In_465,In_248);
or U419 (N_419,In_613,In_610);
and U420 (N_420,In_865,In_718);
nor U421 (N_421,In_576,In_117);
and U422 (N_422,In_678,In_611);
nand U423 (N_423,In_841,In_546);
nor U424 (N_424,In_82,In_780);
or U425 (N_425,In_175,In_714);
nor U426 (N_426,In_342,In_274);
xor U427 (N_427,In_503,In_271);
and U428 (N_428,In_859,In_607);
or U429 (N_429,In_103,In_169);
and U430 (N_430,In_612,In_199);
nand U431 (N_431,In_869,In_599);
nor U432 (N_432,In_124,In_428);
or U433 (N_433,In_337,In_485);
nand U434 (N_434,In_924,In_283);
nor U435 (N_435,In_441,In_276);
and U436 (N_436,In_50,In_241);
and U437 (N_437,In_220,In_266);
nor U438 (N_438,In_435,In_151);
nand U439 (N_439,In_368,In_409);
and U440 (N_440,In_32,In_252);
and U441 (N_441,In_785,In_371);
or U442 (N_442,In_891,In_845);
nand U443 (N_443,In_805,In_47);
or U444 (N_444,In_853,In_676);
or U445 (N_445,In_455,In_544);
and U446 (N_446,In_843,In_946);
nand U447 (N_447,In_213,In_250);
or U448 (N_448,In_526,In_939);
nand U449 (N_449,In_883,In_439);
nand U450 (N_450,In_201,In_759);
or U451 (N_451,In_793,In_801);
nand U452 (N_452,In_968,In_890);
and U453 (N_453,In_758,In_725);
nand U454 (N_454,In_693,In_7);
and U455 (N_455,In_457,In_89);
or U456 (N_456,In_273,In_690);
or U457 (N_457,In_790,In_334);
nand U458 (N_458,In_621,In_524);
nor U459 (N_459,In_187,In_227);
nor U460 (N_460,In_762,In_797);
nor U461 (N_461,In_627,In_167);
or U462 (N_462,In_205,In_706);
or U463 (N_463,In_708,In_404);
and U464 (N_464,In_590,In_667);
nand U465 (N_465,In_794,In_739);
and U466 (N_466,In_940,In_126);
or U467 (N_467,In_689,In_464);
nor U468 (N_468,In_567,In_799);
nor U469 (N_469,In_483,In_195);
and U470 (N_470,In_721,In_818);
and U471 (N_471,In_430,In_478);
and U472 (N_472,In_403,In_656);
and U473 (N_473,In_997,In_665);
nand U474 (N_474,In_809,In_70);
or U475 (N_475,In_639,In_301);
nand U476 (N_476,In_626,In_548);
or U477 (N_477,In_93,In_11);
nand U478 (N_478,In_844,In_433);
nand U479 (N_479,In_715,In_728);
and U480 (N_480,In_179,In_885);
nor U481 (N_481,In_770,In_870);
nand U482 (N_482,In_697,In_115);
or U483 (N_483,In_705,In_628);
or U484 (N_484,In_242,In_565);
or U485 (N_485,In_515,In_90);
nand U486 (N_486,In_307,In_314);
nand U487 (N_487,In_914,In_523);
and U488 (N_488,In_698,In_680);
and U489 (N_489,In_614,In_39);
or U490 (N_490,In_906,In_660);
or U491 (N_491,In_31,In_642);
xor U492 (N_492,In_531,In_240);
nor U493 (N_493,In_335,In_159);
and U494 (N_494,In_96,In_677);
nor U495 (N_495,In_738,In_919);
nor U496 (N_496,In_444,In_139);
or U497 (N_497,In_675,In_425);
or U498 (N_498,In_484,In_290);
or U499 (N_499,In_135,In_64);
and U500 (N_500,N_464,N_87);
nor U501 (N_501,N_264,N_387);
xor U502 (N_502,N_370,N_235);
nand U503 (N_503,N_32,N_498);
nor U504 (N_504,N_189,N_396);
nand U505 (N_505,N_180,N_65);
nor U506 (N_506,N_472,N_167);
and U507 (N_507,N_371,N_291);
and U508 (N_508,N_15,N_380);
nand U509 (N_509,N_321,N_406);
xnor U510 (N_510,N_94,N_285);
nor U511 (N_511,N_379,N_314);
xor U512 (N_512,N_299,N_302);
nor U513 (N_513,N_148,N_146);
or U514 (N_514,N_327,N_51);
nand U515 (N_515,N_211,N_57);
nand U516 (N_516,N_471,N_363);
and U517 (N_517,N_455,N_177);
nand U518 (N_518,N_53,N_295);
or U519 (N_519,N_277,N_438);
and U520 (N_520,N_384,N_428);
nand U521 (N_521,N_325,N_267);
and U522 (N_522,N_322,N_116);
or U523 (N_523,N_290,N_23);
or U524 (N_524,N_328,N_427);
xnor U525 (N_525,N_447,N_89);
nand U526 (N_526,N_304,N_75);
xnor U527 (N_527,N_296,N_147);
or U528 (N_528,N_338,N_160);
and U529 (N_529,N_181,N_8);
xnor U530 (N_530,N_303,N_256);
and U531 (N_531,N_491,N_381);
nand U532 (N_532,N_198,N_445);
nor U533 (N_533,N_400,N_193);
and U534 (N_534,N_376,N_190);
nor U535 (N_535,N_217,N_297);
or U536 (N_536,N_203,N_305);
and U537 (N_537,N_333,N_108);
xnor U538 (N_538,N_310,N_431);
and U539 (N_539,N_90,N_336);
nor U540 (N_540,N_154,N_174);
nand U541 (N_541,N_96,N_214);
and U542 (N_542,N_166,N_492);
and U543 (N_543,N_76,N_298);
and U544 (N_544,N_481,N_258);
or U545 (N_545,N_266,N_342);
nor U546 (N_546,N_330,N_262);
and U547 (N_547,N_42,N_357);
nor U548 (N_548,N_421,N_317);
and U549 (N_549,N_182,N_142);
nand U550 (N_550,N_286,N_229);
nand U551 (N_551,N_58,N_137);
nand U552 (N_552,N_369,N_412);
or U553 (N_553,N_268,N_62);
nor U554 (N_554,N_326,N_403);
nand U555 (N_555,N_165,N_402);
and U556 (N_556,N_139,N_3);
or U557 (N_557,N_239,N_155);
nand U558 (N_558,N_372,N_453);
nand U559 (N_559,N_91,N_483);
and U560 (N_560,N_360,N_233);
or U561 (N_561,N_176,N_64);
or U562 (N_562,N_104,N_365);
or U563 (N_563,N_207,N_458);
or U564 (N_564,N_63,N_187);
nor U565 (N_565,N_476,N_465);
and U566 (N_566,N_39,N_237);
nor U567 (N_567,N_88,N_16);
or U568 (N_568,N_440,N_47);
nand U569 (N_569,N_13,N_331);
nor U570 (N_570,N_417,N_113);
nand U571 (N_571,N_468,N_388);
or U572 (N_572,N_257,N_279);
and U573 (N_573,N_119,N_393);
nand U574 (N_574,N_287,N_289);
nor U575 (N_575,N_54,N_430);
and U576 (N_576,N_272,N_121);
nor U577 (N_577,N_485,N_419);
and U578 (N_578,N_78,N_347);
or U579 (N_579,N_115,N_294);
and U580 (N_580,N_143,N_474);
nand U581 (N_581,N_339,N_409);
nand U582 (N_582,N_101,N_212);
and U583 (N_583,N_43,N_374);
nor U584 (N_584,N_240,N_111);
or U585 (N_585,N_24,N_199);
and U586 (N_586,N_40,N_102);
and U587 (N_587,N_467,N_225);
nand U588 (N_588,N_110,N_126);
or U589 (N_589,N_79,N_263);
xor U590 (N_590,N_224,N_394);
or U591 (N_591,N_466,N_209);
nor U592 (N_592,N_316,N_29);
nand U593 (N_593,N_318,N_171);
or U594 (N_594,N_249,N_169);
and U595 (N_595,N_118,N_20);
and U596 (N_596,N_50,N_488);
nor U597 (N_597,N_486,N_25);
nand U598 (N_598,N_346,N_22);
nand U599 (N_599,N_80,N_105);
or U600 (N_600,N_140,N_103);
nor U601 (N_601,N_270,N_74);
and U602 (N_602,N_49,N_109);
nand U603 (N_603,N_276,N_202);
nor U604 (N_604,N_236,N_153);
and U605 (N_605,N_460,N_259);
nand U606 (N_606,N_30,N_292);
and U607 (N_607,N_238,N_86);
and U608 (N_608,N_136,N_200);
nor U609 (N_609,N_141,N_52);
and U610 (N_610,N_130,N_213);
nor U611 (N_611,N_68,N_344);
xor U612 (N_612,N_125,N_149);
or U613 (N_613,N_21,N_461);
or U614 (N_614,N_329,N_28);
nand U615 (N_615,N_332,N_245);
or U616 (N_616,N_367,N_73);
nor U617 (N_617,N_389,N_281);
or U618 (N_618,N_399,N_38);
nor U619 (N_619,N_271,N_422);
or U620 (N_620,N_114,N_34);
nor U621 (N_621,N_429,N_250);
and U622 (N_622,N_10,N_210);
and U623 (N_623,N_334,N_172);
nand U624 (N_624,N_248,N_366);
or U625 (N_625,N_46,N_437);
nor U626 (N_626,N_69,N_220);
and U627 (N_627,N_67,N_127);
nor U628 (N_628,N_82,N_335);
or U629 (N_629,N_255,N_66);
nor U630 (N_630,N_383,N_418);
nor U631 (N_631,N_1,N_478);
and U632 (N_632,N_443,N_72);
nand U633 (N_633,N_497,N_92);
nor U634 (N_634,N_283,N_247);
or U635 (N_635,N_222,N_494);
nor U636 (N_636,N_61,N_161);
or U637 (N_637,N_480,N_456);
nor U638 (N_638,N_19,N_435);
or U639 (N_639,N_164,N_37);
and U640 (N_640,N_473,N_133);
or U641 (N_641,N_151,N_162);
xor U642 (N_642,N_186,N_395);
and U643 (N_643,N_85,N_426);
and U644 (N_644,N_132,N_31);
nand U645 (N_645,N_231,N_373);
and U646 (N_646,N_392,N_244);
nand U647 (N_647,N_191,N_309);
nand U648 (N_648,N_470,N_420);
and U649 (N_649,N_463,N_205);
and U650 (N_650,N_232,N_44);
and U651 (N_651,N_386,N_274);
nand U652 (N_652,N_441,N_145);
nand U653 (N_653,N_451,N_343);
xnor U654 (N_654,N_36,N_14);
or U655 (N_655,N_269,N_156);
and U656 (N_656,N_359,N_265);
or U657 (N_657,N_356,N_196);
nand U658 (N_658,N_228,N_226);
or U659 (N_659,N_218,N_352);
and U660 (N_660,N_227,N_457);
and U661 (N_661,N_444,N_35);
or U662 (N_662,N_98,N_241);
and U663 (N_663,N_195,N_221);
and U664 (N_664,N_150,N_243);
nand U665 (N_665,N_452,N_183);
or U666 (N_666,N_158,N_407);
or U667 (N_667,N_7,N_157);
or U668 (N_668,N_475,N_434);
nor U669 (N_669,N_301,N_354);
or U670 (N_670,N_489,N_282);
nand U671 (N_671,N_254,N_311);
and U672 (N_672,N_436,N_280);
nor U673 (N_673,N_423,N_323);
nor U674 (N_674,N_405,N_48);
or U675 (N_675,N_391,N_112);
nand U676 (N_676,N_83,N_41);
nor U677 (N_677,N_242,N_275);
or U678 (N_678,N_482,N_230);
and U679 (N_679,N_253,N_93);
nand U680 (N_680,N_197,N_106);
and U681 (N_681,N_495,N_415);
xnor U682 (N_682,N_401,N_77);
and U683 (N_683,N_324,N_84);
and U684 (N_684,N_135,N_18);
nand U685 (N_685,N_144,N_454);
nor U686 (N_686,N_348,N_390);
nand U687 (N_687,N_284,N_95);
or U688 (N_688,N_413,N_0);
nand U689 (N_689,N_4,N_433);
and U690 (N_690,N_131,N_188);
nand U691 (N_691,N_355,N_364);
or U692 (N_692,N_138,N_99);
nor U693 (N_693,N_251,N_410);
nor U694 (N_694,N_117,N_12);
or U695 (N_695,N_351,N_416);
xnor U696 (N_696,N_496,N_273);
or U697 (N_697,N_378,N_362);
or U698 (N_698,N_184,N_17);
and U699 (N_699,N_60,N_201);
nor U700 (N_700,N_70,N_260);
nor U701 (N_701,N_134,N_120);
and U702 (N_702,N_340,N_385);
nand U703 (N_703,N_361,N_204);
and U704 (N_704,N_159,N_313);
or U705 (N_705,N_411,N_179);
and U706 (N_706,N_308,N_300);
nor U707 (N_707,N_246,N_377);
nor U708 (N_708,N_499,N_71);
xnor U709 (N_709,N_382,N_128);
nand U710 (N_710,N_493,N_55);
xnor U711 (N_711,N_448,N_307);
nand U712 (N_712,N_5,N_397);
nand U713 (N_713,N_206,N_219);
nand U714 (N_714,N_306,N_462);
and U715 (N_715,N_26,N_469);
and U716 (N_716,N_185,N_100);
or U717 (N_717,N_2,N_459);
nand U718 (N_718,N_168,N_353);
and U719 (N_719,N_442,N_358);
and U720 (N_720,N_124,N_450);
nand U721 (N_721,N_178,N_477);
nand U722 (N_722,N_261,N_192);
nand U723 (N_723,N_341,N_484);
and U724 (N_724,N_439,N_278);
nand U725 (N_725,N_216,N_170);
or U726 (N_726,N_208,N_408);
or U727 (N_727,N_375,N_425);
and U728 (N_728,N_123,N_312);
nor U729 (N_729,N_350,N_97);
and U730 (N_730,N_449,N_414);
nor U731 (N_731,N_479,N_6);
nand U732 (N_732,N_319,N_81);
nand U733 (N_733,N_59,N_11);
nor U734 (N_734,N_45,N_337);
nand U735 (N_735,N_368,N_315);
nand U736 (N_736,N_446,N_223);
nor U737 (N_737,N_215,N_252);
nand U738 (N_738,N_490,N_288);
nand U739 (N_739,N_424,N_9);
nand U740 (N_740,N_152,N_404);
nand U741 (N_741,N_345,N_27);
nor U742 (N_742,N_173,N_293);
nor U743 (N_743,N_33,N_487);
and U744 (N_744,N_163,N_194);
and U745 (N_745,N_175,N_320);
and U746 (N_746,N_56,N_122);
and U747 (N_747,N_432,N_129);
nor U748 (N_748,N_234,N_349);
or U749 (N_749,N_398,N_107);
or U750 (N_750,N_348,N_38);
and U751 (N_751,N_433,N_185);
and U752 (N_752,N_363,N_41);
or U753 (N_753,N_313,N_141);
and U754 (N_754,N_440,N_223);
or U755 (N_755,N_265,N_31);
or U756 (N_756,N_175,N_292);
or U757 (N_757,N_489,N_119);
nor U758 (N_758,N_248,N_35);
and U759 (N_759,N_12,N_419);
nor U760 (N_760,N_291,N_321);
and U761 (N_761,N_457,N_83);
nor U762 (N_762,N_313,N_250);
and U763 (N_763,N_108,N_372);
nand U764 (N_764,N_118,N_398);
nand U765 (N_765,N_250,N_271);
xnor U766 (N_766,N_296,N_175);
nand U767 (N_767,N_200,N_211);
nor U768 (N_768,N_477,N_160);
nor U769 (N_769,N_435,N_288);
nor U770 (N_770,N_211,N_257);
nand U771 (N_771,N_434,N_34);
xor U772 (N_772,N_259,N_343);
and U773 (N_773,N_287,N_273);
nand U774 (N_774,N_324,N_46);
and U775 (N_775,N_359,N_194);
and U776 (N_776,N_423,N_133);
and U777 (N_777,N_34,N_75);
or U778 (N_778,N_129,N_106);
xor U779 (N_779,N_428,N_203);
nor U780 (N_780,N_226,N_57);
nor U781 (N_781,N_33,N_347);
and U782 (N_782,N_250,N_305);
or U783 (N_783,N_75,N_477);
and U784 (N_784,N_425,N_361);
nand U785 (N_785,N_137,N_317);
or U786 (N_786,N_86,N_458);
and U787 (N_787,N_495,N_44);
nor U788 (N_788,N_205,N_374);
or U789 (N_789,N_117,N_390);
and U790 (N_790,N_359,N_240);
nor U791 (N_791,N_350,N_168);
nor U792 (N_792,N_325,N_419);
or U793 (N_793,N_419,N_229);
or U794 (N_794,N_463,N_424);
nor U795 (N_795,N_431,N_498);
and U796 (N_796,N_249,N_165);
or U797 (N_797,N_44,N_138);
nor U798 (N_798,N_53,N_374);
nand U799 (N_799,N_130,N_176);
xnor U800 (N_800,N_193,N_243);
and U801 (N_801,N_412,N_201);
or U802 (N_802,N_493,N_229);
nor U803 (N_803,N_396,N_284);
and U804 (N_804,N_147,N_100);
nand U805 (N_805,N_381,N_95);
nand U806 (N_806,N_472,N_259);
or U807 (N_807,N_83,N_447);
nor U808 (N_808,N_344,N_227);
nor U809 (N_809,N_324,N_315);
xnor U810 (N_810,N_14,N_270);
nand U811 (N_811,N_260,N_8);
nor U812 (N_812,N_197,N_460);
and U813 (N_813,N_320,N_163);
nand U814 (N_814,N_377,N_113);
nor U815 (N_815,N_171,N_226);
and U816 (N_816,N_319,N_310);
or U817 (N_817,N_462,N_209);
or U818 (N_818,N_322,N_111);
xor U819 (N_819,N_153,N_466);
nor U820 (N_820,N_29,N_471);
nor U821 (N_821,N_430,N_384);
and U822 (N_822,N_429,N_0);
or U823 (N_823,N_377,N_459);
and U824 (N_824,N_190,N_96);
or U825 (N_825,N_11,N_20);
and U826 (N_826,N_360,N_431);
or U827 (N_827,N_424,N_108);
nand U828 (N_828,N_442,N_225);
nor U829 (N_829,N_214,N_389);
and U830 (N_830,N_488,N_105);
nor U831 (N_831,N_173,N_33);
nor U832 (N_832,N_230,N_451);
nand U833 (N_833,N_184,N_213);
nand U834 (N_834,N_224,N_161);
and U835 (N_835,N_226,N_70);
nand U836 (N_836,N_464,N_128);
or U837 (N_837,N_469,N_81);
or U838 (N_838,N_471,N_183);
or U839 (N_839,N_40,N_344);
xnor U840 (N_840,N_482,N_476);
nand U841 (N_841,N_146,N_34);
and U842 (N_842,N_459,N_409);
or U843 (N_843,N_409,N_377);
and U844 (N_844,N_432,N_267);
nor U845 (N_845,N_430,N_180);
nand U846 (N_846,N_130,N_342);
nand U847 (N_847,N_405,N_357);
nor U848 (N_848,N_261,N_153);
and U849 (N_849,N_349,N_324);
or U850 (N_850,N_221,N_162);
nand U851 (N_851,N_316,N_124);
and U852 (N_852,N_14,N_256);
or U853 (N_853,N_433,N_403);
nand U854 (N_854,N_400,N_419);
and U855 (N_855,N_257,N_167);
xor U856 (N_856,N_304,N_37);
or U857 (N_857,N_329,N_481);
nor U858 (N_858,N_148,N_179);
nor U859 (N_859,N_45,N_307);
nor U860 (N_860,N_449,N_109);
and U861 (N_861,N_198,N_333);
or U862 (N_862,N_112,N_128);
or U863 (N_863,N_173,N_346);
or U864 (N_864,N_289,N_332);
and U865 (N_865,N_127,N_12);
and U866 (N_866,N_338,N_167);
and U867 (N_867,N_33,N_169);
and U868 (N_868,N_471,N_128);
xnor U869 (N_869,N_17,N_475);
or U870 (N_870,N_423,N_123);
or U871 (N_871,N_272,N_327);
nor U872 (N_872,N_60,N_84);
nand U873 (N_873,N_337,N_64);
nand U874 (N_874,N_177,N_330);
nor U875 (N_875,N_332,N_360);
or U876 (N_876,N_425,N_441);
nor U877 (N_877,N_224,N_105);
nor U878 (N_878,N_352,N_235);
or U879 (N_879,N_393,N_292);
nor U880 (N_880,N_433,N_20);
or U881 (N_881,N_406,N_2);
xor U882 (N_882,N_390,N_371);
nand U883 (N_883,N_172,N_395);
and U884 (N_884,N_74,N_160);
nor U885 (N_885,N_79,N_55);
nor U886 (N_886,N_68,N_256);
or U887 (N_887,N_301,N_391);
and U888 (N_888,N_352,N_345);
nand U889 (N_889,N_114,N_430);
or U890 (N_890,N_474,N_227);
nand U891 (N_891,N_75,N_254);
and U892 (N_892,N_51,N_298);
nor U893 (N_893,N_238,N_383);
or U894 (N_894,N_293,N_194);
or U895 (N_895,N_23,N_372);
nand U896 (N_896,N_323,N_442);
nand U897 (N_897,N_92,N_155);
and U898 (N_898,N_376,N_52);
or U899 (N_899,N_483,N_486);
nand U900 (N_900,N_206,N_282);
or U901 (N_901,N_446,N_335);
or U902 (N_902,N_203,N_31);
nor U903 (N_903,N_97,N_45);
nor U904 (N_904,N_297,N_235);
nor U905 (N_905,N_372,N_18);
or U906 (N_906,N_44,N_387);
nand U907 (N_907,N_161,N_28);
nor U908 (N_908,N_246,N_171);
nor U909 (N_909,N_355,N_383);
or U910 (N_910,N_260,N_164);
nand U911 (N_911,N_375,N_260);
and U912 (N_912,N_150,N_399);
and U913 (N_913,N_442,N_217);
xnor U914 (N_914,N_329,N_314);
or U915 (N_915,N_218,N_346);
and U916 (N_916,N_333,N_129);
and U917 (N_917,N_491,N_438);
xor U918 (N_918,N_474,N_150);
and U919 (N_919,N_258,N_314);
nand U920 (N_920,N_342,N_483);
and U921 (N_921,N_3,N_142);
and U922 (N_922,N_448,N_137);
and U923 (N_923,N_455,N_406);
or U924 (N_924,N_178,N_282);
and U925 (N_925,N_477,N_127);
nor U926 (N_926,N_196,N_345);
nor U927 (N_927,N_414,N_453);
nor U928 (N_928,N_417,N_206);
and U929 (N_929,N_384,N_396);
nand U930 (N_930,N_132,N_84);
nand U931 (N_931,N_129,N_37);
nor U932 (N_932,N_214,N_72);
or U933 (N_933,N_102,N_427);
and U934 (N_934,N_350,N_392);
xor U935 (N_935,N_296,N_269);
nor U936 (N_936,N_461,N_104);
and U937 (N_937,N_459,N_122);
nand U938 (N_938,N_40,N_121);
nand U939 (N_939,N_18,N_162);
nor U940 (N_940,N_20,N_453);
nor U941 (N_941,N_422,N_223);
and U942 (N_942,N_364,N_303);
nand U943 (N_943,N_241,N_217);
and U944 (N_944,N_213,N_86);
or U945 (N_945,N_297,N_246);
or U946 (N_946,N_332,N_482);
and U947 (N_947,N_377,N_481);
nor U948 (N_948,N_353,N_127);
nor U949 (N_949,N_111,N_282);
nand U950 (N_950,N_442,N_403);
nor U951 (N_951,N_24,N_191);
and U952 (N_952,N_406,N_46);
nor U953 (N_953,N_280,N_287);
nor U954 (N_954,N_438,N_222);
and U955 (N_955,N_183,N_122);
and U956 (N_956,N_63,N_229);
or U957 (N_957,N_54,N_409);
xnor U958 (N_958,N_456,N_148);
and U959 (N_959,N_333,N_229);
and U960 (N_960,N_154,N_463);
or U961 (N_961,N_139,N_230);
or U962 (N_962,N_389,N_279);
nor U963 (N_963,N_441,N_394);
nor U964 (N_964,N_175,N_0);
nor U965 (N_965,N_385,N_429);
or U966 (N_966,N_425,N_144);
nor U967 (N_967,N_71,N_397);
nand U968 (N_968,N_363,N_407);
and U969 (N_969,N_265,N_111);
and U970 (N_970,N_175,N_345);
nor U971 (N_971,N_105,N_186);
and U972 (N_972,N_196,N_341);
or U973 (N_973,N_268,N_53);
and U974 (N_974,N_65,N_366);
nor U975 (N_975,N_232,N_314);
nor U976 (N_976,N_255,N_242);
and U977 (N_977,N_100,N_403);
or U978 (N_978,N_302,N_269);
or U979 (N_979,N_218,N_397);
nand U980 (N_980,N_342,N_211);
or U981 (N_981,N_94,N_373);
nand U982 (N_982,N_19,N_268);
and U983 (N_983,N_326,N_42);
nor U984 (N_984,N_314,N_5);
nor U985 (N_985,N_343,N_445);
or U986 (N_986,N_142,N_72);
or U987 (N_987,N_50,N_442);
nor U988 (N_988,N_338,N_414);
nor U989 (N_989,N_464,N_191);
and U990 (N_990,N_165,N_294);
nor U991 (N_991,N_139,N_55);
nand U992 (N_992,N_255,N_307);
nor U993 (N_993,N_6,N_269);
and U994 (N_994,N_75,N_444);
nor U995 (N_995,N_362,N_44);
nor U996 (N_996,N_230,N_473);
or U997 (N_997,N_321,N_31);
or U998 (N_998,N_97,N_469);
nor U999 (N_999,N_348,N_141);
nor U1000 (N_1000,N_526,N_851);
nand U1001 (N_1001,N_621,N_798);
and U1002 (N_1002,N_728,N_883);
nand U1003 (N_1003,N_508,N_685);
nor U1004 (N_1004,N_680,N_555);
nand U1005 (N_1005,N_896,N_747);
and U1006 (N_1006,N_639,N_664);
nor U1007 (N_1007,N_834,N_749);
nand U1008 (N_1008,N_674,N_736);
nand U1009 (N_1009,N_960,N_886);
nand U1010 (N_1010,N_977,N_507);
nand U1011 (N_1011,N_585,N_676);
nor U1012 (N_1012,N_908,N_697);
nand U1013 (N_1013,N_796,N_524);
nand U1014 (N_1014,N_564,N_840);
nor U1015 (N_1015,N_945,N_907);
or U1016 (N_1016,N_829,N_916);
or U1017 (N_1017,N_765,N_751);
nand U1018 (N_1018,N_666,N_737);
nor U1019 (N_1019,N_876,N_503);
nor U1020 (N_1020,N_641,N_627);
or U1021 (N_1021,N_784,N_826);
or U1022 (N_1022,N_970,N_567);
nand U1023 (N_1023,N_578,N_910);
or U1024 (N_1024,N_689,N_677);
or U1025 (N_1025,N_501,N_645);
and U1026 (N_1026,N_963,N_912);
xnor U1027 (N_1027,N_763,N_861);
and U1028 (N_1028,N_904,N_981);
or U1029 (N_1029,N_563,N_922);
and U1030 (N_1030,N_815,N_832);
and U1031 (N_1031,N_619,N_636);
nor U1032 (N_1032,N_787,N_618);
and U1033 (N_1033,N_949,N_545);
nor U1034 (N_1034,N_573,N_661);
or U1035 (N_1035,N_571,N_761);
or U1036 (N_1036,N_790,N_983);
nand U1037 (N_1037,N_962,N_565);
or U1038 (N_1038,N_593,N_948);
nand U1039 (N_1039,N_748,N_616);
nor U1040 (N_1040,N_679,N_793);
or U1041 (N_1041,N_600,N_538);
and U1042 (N_1042,N_993,N_810);
or U1043 (N_1043,N_506,N_601);
nand U1044 (N_1044,N_668,N_724);
nor U1045 (N_1045,N_837,N_505);
nor U1046 (N_1046,N_959,N_732);
and U1047 (N_1047,N_591,N_660);
nand U1048 (N_1048,N_688,N_942);
nor U1049 (N_1049,N_541,N_650);
and U1050 (N_1050,N_930,N_788);
and U1051 (N_1051,N_821,N_580);
nor U1052 (N_1052,N_553,N_570);
nand U1053 (N_1053,N_917,N_850);
nand U1054 (N_1054,N_781,N_675);
nand U1055 (N_1055,N_903,N_870);
nor U1056 (N_1056,N_905,N_901);
or U1057 (N_1057,N_986,N_865);
and U1058 (N_1058,N_766,N_739);
or U1059 (N_1059,N_969,N_828);
and U1060 (N_1060,N_864,N_682);
or U1061 (N_1061,N_527,N_574);
and U1062 (N_1062,N_509,N_534);
xor U1063 (N_1063,N_672,N_562);
and U1064 (N_1064,N_590,N_695);
or U1065 (N_1065,N_568,N_950);
nand U1066 (N_1066,N_975,N_909);
or U1067 (N_1067,N_898,N_684);
nand U1068 (N_1068,N_806,N_956);
or U1069 (N_1069,N_757,N_596);
nand U1070 (N_1070,N_953,N_741);
and U1071 (N_1071,N_731,N_632);
and U1072 (N_1072,N_520,N_577);
and U1073 (N_1073,N_902,N_702);
and U1074 (N_1074,N_657,N_719);
or U1075 (N_1075,N_853,N_770);
nor U1076 (N_1076,N_549,N_722);
or U1077 (N_1077,N_807,N_831);
or U1078 (N_1078,N_725,N_536);
and U1079 (N_1079,N_974,N_889);
or U1080 (N_1080,N_811,N_566);
nor U1081 (N_1081,N_871,N_873);
and U1082 (N_1082,N_822,N_935);
nand U1083 (N_1083,N_671,N_995);
nand U1084 (N_1084,N_704,N_780);
and U1085 (N_1085,N_631,N_699);
nand U1086 (N_1086,N_880,N_537);
nor U1087 (N_1087,N_595,N_978);
nand U1088 (N_1088,N_965,N_718);
and U1089 (N_1089,N_510,N_630);
xnor U1090 (N_1090,N_643,N_698);
or U1091 (N_1091,N_654,N_827);
nand U1092 (N_1092,N_838,N_771);
and U1093 (N_1093,N_813,N_523);
xor U1094 (N_1094,N_852,N_554);
and U1095 (N_1095,N_769,N_795);
or U1096 (N_1096,N_745,N_786);
nor U1097 (N_1097,N_946,N_655);
nand U1098 (N_1098,N_777,N_597);
nor U1099 (N_1099,N_775,N_584);
or U1100 (N_1100,N_872,N_620);
nor U1101 (N_1101,N_622,N_874);
nor U1102 (N_1102,N_594,N_947);
nand U1103 (N_1103,N_516,N_605);
or U1104 (N_1104,N_670,N_586);
nand U1105 (N_1105,N_954,N_525);
and U1106 (N_1106,N_936,N_797);
and U1107 (N_1107,N_729,N_713);
and U1108 (N_1108,N_642,N_714);
and U1109 (N_1109,N_955,N_712);
nand U1110 (N_1110,N_692,N_881);
nand U1111 (N_1111,N_637,N_967);
or U1112 (N_1112,N_681,N_701);
and U1113 (N_1113,N_693,N_742);
or U1114 (N_1114,N_663,N_548);
and U1115 (N_1115,N_860,N_891);
nand U1116 (N_1116,N_502,N_721);
and U1117 (N_1117,N_938,N_653);
or U1118 (N_1118,N_820,N_706);
and U1119 (N_1119,N_530,N_603);
and U1120 (N_1120,N_613,N_550);
nand U1121 (N_1121,N_980,N_687);
and U1122 (N_1122,N_733,N_939);
or U1123 (N_1123,N_964,N_992);
and U1124 (N_1124,N_582,N_515);
nor U1125 (N_1125,N_934,N_919);
nor U1126 (N_1126,N_924,N_823);
nor U1127 (N_1127,N_707,N_705);
and U1128 (N_1128,N_996,N_500);
nor U1129 (N_1129,N_859,N_547);
nand U1130 (N_1130,N_615,N_740);
nand U1131 (N_1131,N_892,N_875);
nand U1132 (N_1132,N_858,N_669);
or U1133 (N_1133,N_957,N_890);
or U1134 (N_1134,N_849,N_678);
nand U1135 (N_1135,N_543,N_906);
or U1136 (N_1136,N_843,N_624);
xnor U1137 (N_1137,N_973,N_709);
nand U1138 (N_1138,N_762,N_990);
and U1139 (N_1139,N_521,N_800);
nand U1140 (N_1140,N_783,N_649);
nand U1141 (N_1141,N_551,N_504);
and U1142 (N_1142,N_928,N_931);
or U1143 (N_1143,N_626,N_517);
or U1144 (N_1144,N_589,N_855);
nor U1145 (N_1145,N_971,N_791);
nor U1146 (N_1146,N_529,N_801);
nor U1147 (N_1147,N_662,N_606);
and U1148 (N_1148,N_772,N_633);
or U1149 (N_1149,N_885,N_998);
nor U1150 (N_1150,N_544,N_799);
nor U1151 (N_1151,N_921,N_514);
nor U1152 (N_1152,N_560,N_532);
and U1153 (N_1153,N_968,N_617);
nand U1154 (N_1154,N_792,N_857);
and U1155 (N_1155,N_744,N_816);
and U1156 (N_1156,N_929,N_989);
or U1157 (N_1157,N_743,N_528);
nand U1158 (N_1158,N_734,N_542);
nor U1159 (N_1159,N_767,N_623);
xor U1160 (N_1160,N_839,N_652);
nor U1161 (N_1161,N_760,N_836);
nor U1162 (N_1162,N_863,N_943);
and U1163 (N_1163,N_915,N_647);
or U1164 (N_1164,N_588,N_776);
nor U1165 (N_1165,N_899,N_944);
nor U1166 (N_1166,N_690,N_941);
and U1167 (N_1167,N_835,N_561);
nor U1168 (N_1168,N_691,N_862);
or U1169 (N_1169,N_779,N_844);
and U1170 (N_1170,N_696,N_878);
nand U1171 (N_1171,N_976,N_609);
or U1172 (N_1172,N_940,N_755);
nor U1173 (N_1173,N_535,N_854);
nor U1174 (N_1174,N_894,N_985);
nand U1175 (N_1175,N_756,N_830);
nand U1176 (N_1176,N_966,N_531);
or U1177 (N_1177,N_644,N_819);
and U1178 (N_1178,N_809,N_559);
or U1179 (N_1179,N_884,N_753);
or U1180 (N_1180,N_614,N_808);
or U1181 (N_1181,N_758,N_764);
or U1182 (N_1182,N_727,N_683);
and U1183 (N_1183,N_867,N_895);
or U1184 (N_1184,N_557,N_982);
or U1185 (N_1185,N_932,N_686);
or U1186 (N_1186,N_552,N_715);
and U1187 (N_1187,N_846,N_768);
nor U1188 (N_1188,N_658,N_583);
or U1189 (N_1189,N_752,N_625);
nor U1190 (N_1190,N_694,N_711);
and U1191 (N_1191,N_994,N_735);
nor U1192 (N_1192,N_925,N_598);
nor U1193 (N_1193,N_716,N_911);
nor U1194 (N_1194,N_599,N_754);
or U1195 (N_1195,N_604,N_556);
xor U1196 (N_1196,N_634,N_611);
and U1197 (N_1197,N_511,N_888);
and U1198 (N_1198,N_825,N_856);
or U1199 (N_1199,N_628,N_656);
nand U1200 (N_1200,N_659,N_952);
and U1201 (N_1201,N_805,N_607);
and U1202 (N_1202,N_984,N_900);
or U1203 (N_1203,N_738,N_665);
nand U1204 (N_1204,N_866,N_927);
or U1205 (N_1205,N_773,N_778);
and U1206 (N_1206,N_845,N_958);
nand U1207 (N_1207,N_794,N_897);
nor U1208 (N_1208,N_882,N_914);
or U1209 (N_1209,N_804,N_602);
nand U1210 (N_1210,N_893,N_569);
nand U1211 (N_1211,N_723,N_629);
nor U1212 (N_1212,N_802,N_726);
nand U1213 (N_1213,N_592,N_841);
nand U1214 (N_1214,N_518,N_951);
and U1215 (N_1215,N_558,N_920);
nor U1216 (N_1216,N_869,N_812);
xor U1217 (N_1217,N_785,N_750);
nand U1218 (N_1218,N_847,N_774);
and U1219 (N_1219,N_879,N_887);
and U1220 (N_1220,N_933,N_710);
and U1221 (N_1221,N_972,N_638);
and U1222 (N_1222,N_646,N_987);
and U1223 (N_1223,N_519,N_817);
or U1224 (N_1224,N_640,N_575);
or U1225 (N_1225,N_540,N_824);
nor U1226 (N_1226,N_576,N_789);
and U1227 (N_1227,N_877,N_997);
nand U1228 (N_1228,N_546,N_923);
nand U1229 (N_1229,N_581,N_579);
and U1230 (N_1230,N_814,N_651);
nand U1231 (N_1231,N_759,N_610);
and U1232 (N_1232,N_673,N_926);
nor U1233 (N_1233,N_918,N_533);
nor U1234 (N_1234,N_842,N_868);
nor U1235 (N_1235,N_700,N_730);
xor U1236 (N_1236,N_539,N_913);
nor U1237 (N_1237,N_512,N_818);
nand U1238 (N_1238,N_937,N_988);
or U1239 (N_1239,N_991,N_572);
nand U1240 (N_1240,N_803,N_746);
nand U1241 (N_1241,N_708,N_635);
nor U1242 (N_1242,N_522,N_720);
nand U1243 (N_1243,N_648,N_608);
and U1244 (N_1244,N_961,N_833);
nor U1245 (N_1245,N_513,N_848);
nand U1246 (N_1246,N_782,N_717);
and U1247 (N_1247,N_667,N_587);
nand U1248 (N_1248,N_612,N_979);
nand U1249 (N_1249,N_999,N_703);
or U1250 (N_1250,N_572,N_832);
nand U1251 (N_1251,N_751,N_901);
and U1252 (N_1252,N_796,N_528);
nor U1253 (N_1253,N_879,N_748);
or U1254 (N_1254,N_966,N_741);
and U1255 (N_1255,N_544,N_719);
nand U1256 (N_1256,N_839,N_681);
xor U1257 (N_1257,N_517,N_989);
nor U1258 (N_1258,N_947,N_799);
nand U1259 (N_1259,N_891,N_796);
nand U1260 (N_1260,N_952,N_580);
and U1261 (N_1261,N_758,N_775);
nand U1262 (N_1262,N_860,N_714);
and U1263 (N_1263,N_928,N_500);
nor U1264 (N_1264,N_624,N_970);
nor U1265 (N_1265,N_895,N_555);
nor U1266 (N_1266,N_791,N_746);
or U1267 (N_1267,N_832,N_687);
nand U1268 (N_1268,N_841,N_908);
nand U1269 (N_1269,N_520,N_726);
nor U1270 (N_1270,N_902,N_653);
nor U1271 (N_1271,N_861,N_722);
nand U1272 (N_1272,N_599,N_706);
or U1273 (N_1273,N_623,N_649);
or U1274 (N_1274,N_701,N_791);
nor U1275 (N_1275,N_592,N_573);
or U1276 (N_1276,N_942,N_813);
nand U1277 (N_1277,N_853,N_656);
or U1278 (N_1278,N_559,N_902);
or U1279 (N_1279,N_612,N_813);
xor U1280 (N_1280,N_946,N_554);
nand U1281 (N_1281,N_514,N_612);
and U1282 (N_1282,N_997,N_939);
nor U1283 (N_1283,N_823,N_639);
nor U1284 (N_1284,N_693,N_641);
nor U1285 (N_1285,N_501,N_788);
or U1286 (N_1286,N_537,N_817);
xnor U1287 (N_1287,N_630,N_866);
xnor U1288 (N_1288,N_783,N_954);
xnor U1289 (N_1289,N_701,N_808);
or U1290 (N_1290,N_832,N_831);
or U1291 (N_1291,N_500,N_836);
xor U1292 (N_1292,N_736,N_508);
nor U1293 (N_1293,N_789,N_764);
nor U1294 (N_1294,N_704,N_805);
and U1295 (N_1295,N_685,N_910);
and U1296 (N_1296,N_700,N_981);
and U1297 (N_1297,N_624,N_694);
and U1298 (N_1298,N_979,N_864);
nand U1299 (N_1299,N_785,N_629);
xnor U1300 (N_1300,N_789,N_571);
or U1301 (N_1301,N_749,N_924);
nand U1302 (N_1302,N_787,N_509);
nor U1303 (N_1303,N_571,N_700);
or U1304 (N_1304,N_619,N_839);
or U1305 (N_1305,N_793,N_929);
and U1306 (N_1306,N_608,N_783);
nand U1307 (N_1307,N_738,N_675);
or U1308 (N_1308,N_938,N_822);
nand U1309 (N_1309,N_603,N_764);
and U1310 (N_1310,N_916,N_702);
or U1311 (N_1311,N_811,N_808);
or U1312 (N_1312,N_802,N_831);
nor U1313 (N_1313,N_770,N_637);
nand U1314 (N_1314,N_610,N_616);
and U1315 (N_1315,N_742,N_532);
or U1316 (N_1316,N_946,N_873);
nor U1317 (N_1317,N_807,N_549);
and U1318 (N_1318,N_863,N_591);
nand U1319 (N_1319,N_791,N_642);
nand U1320 (N_1320,N_671,N_860);
and U1321 (N_1321,N_648,N_674);
nand U1322 (N_1322,N_926,N_631);
xor U1323 (N_1323,N_552,N_813);
or U1324 (N_1324,N_783,N_901);
or U1325 (N_1325,N_918,N_950);
and U1326 (N_1326,N_545,N_623);
and U1327 (N_1327,N_806,N_845);
and U1328 (N_1328,N_801,N_616);
nor U1329 (N_1329,N_908,N_999);
or U1330 (N_1330,N_778,N_745);
and U1331 (N_1331,N_652,N_894);
and U1332 (N_1332,N_780,N_991);
nor U1333 (N_1333,N_824,N_783);
nand U1334 (N_1334,N_807,N_535);
nand U1335 (N_1335,N_688,N_558);
and U1336 (N_1336,N_665,N_951);
or U1337 (N_1337,N_995,N_628);
nor U1338 (N_1338,N_749,N_767);
or U1339 (N_1339,N_806,N_515);
or U1340 (N_1340,N_988,N_720);
nor U1341 (N_1341,N_612,N_540);
and U1342 (N_1342,N_830,N_949);
or U1343 (N_1343,N_940,N_880);
nor U1344 (N_1344,N_827,N_653);
nor U1345 (N_1345,N_787,N_727);
and U1346 (N_1346,N_596,N_553);
xor U1347 (N_1347,N_777,N_976);
nand U1348 (N_1348,N_723,N_925);
or U1349 (N_1349,N_591,N_815);
or U1350 (N_1350,N_564,N_543);
and U1351 (N_1351,N_842,N_755);
or U1352 (N_1352,N_600,N_557);
or U1353 (N_1353,N_565,N_993);
and U1354 (N_1354,N_778,N_908);
and U1355 (N_1355,N_702,N_552);
nand U1356 (N_1356,N_806,N_691);
nand U1357 (N_1357,N_926,N_902);
nand U1358 (N_1358,N_584,N_936);
nor U1359 (N_1359,N_679,N_633);
or U1360 (N_1360,N_709,N_671);
nor U1361 (N_1361,N_654,N_890);
nand U1362 (N_1362,N_862,N_521);
nor U1363 (N_1363,N_680,N_930);
nand U1364 (N_1364,N_693,N_858);
nand U1365 (N_1365,N_802,N_693);
or U1366 (N_1366,N_651,N_615);
xor U1367 (N_1367,N_819,N_888);
and U1368 (N_1368,N_833,N_883);
nand U1369 (N_1369,N_880,N_815);
and U1370 (N_1370,N_910,N_531);
nand U1371 (N_1371,N_670,N_575);
nor U1372 (N_1372,N_664,N_592);
and U1373 (N_1373,N_854,N_978);
or U1374 (N_1374,N_802,N_960);
or U1375 (N_1375,N_908,N_777);
or U1376 (N_1376,N_620,N_747);
nor U1377 (N_1377,N_531,N_522);
or U1378 (N_1378,N_823,N_764);
and U1379 (N_1379,N_709,N_712);
nor U1380 (N_1380,N_874,N_561);
or U1381 (N_1381,N_899,N_904);
and U1382 (N_1382,N_614,N_578);
xnor U1383 (N_1383,N_946,N_527);
nor U1384 (N_1384,N_780,N_759);
or U1385 (N_1385,N_592,N_788);
nand U1386 (N_1386,N_546,N_638);
or U1387 (N_1387,N_768,N_704);
nor U1388 (N_1388,N_705,N_979);
nand U1389 (N_1389,N_723,N_672);
and U1390 (N_1390,N_716,N_839);
or U1391 (N_1391,N_523,N_982);
nor U1392 (N_1392,N_620,N_733);
or U1393 (N_1393,N_651,N_593);
or U1394 (N_1394,N_784,N_593);
nor U1395 (N_1395,N_930,N_870);
or U1396 (N_1396,N_990,N_578);
nand U1397 (N_1397,N_854,N_638);
nor U1398 (N_1398,N_749,N_627);
and U1399 (N_1399,N_716,N_519);
or U1400 (N_1400,N_680,N_896);
nor U1401 (N_1401,N_795,N_629);
or U1402 (N_1402,N_759,N_529);
nor U1403 (N_1403,N_873,N_900);
nor U1404 (N_1404,N_887,N_898);
and U1405 (N_1405,N_721,N_914);
nand U1406 (N_1406,N_628,N_976);
and U1407 (N_1407,N_806,N_683);
xnor U1408 (N_1408,N_860,N_655);
and U1409 (N_1409,N_593,N_899);
nor U1410 (N_1410,N_631,N_528);
nand U1411 (N_1411,N_596,N_738);
and U1412 (N_1412,N_738,N_589);
nand U1413 (N_1413,N_906,N_965);
and U1414 (N_1414,N_632,N_598);
nand U1415 (N_1415,N_694,N_878);
and U1416 (N_1416,N_634,N_754);
and U1417 (N_1417,N_822,N_642);
nand U1418 (N_1418,N_979,N_515);
nand U1419 (N_1419,N_835,N_852);
and U1420 (N_1420,N_859,N_958);
xnor U1421 (N_1421,N_670,N_876);
and U1422 (N_1422,N_827,N_642);
and U1423 (N_1423,N_511,N_790);
and U1424 (N_1424,N_636,N_560);
nand U1425 (N_1425,N_695,N_837);
nor U1426 (N_1426,N_987,N_628);
nand U1427 (N_1427,N_735,N_865);
or U1428 (N_1428,N_779,N_564);
nand U1429 (N_1429,N_645,N_568);
and U1430 (N_1430,N_817,N_526);
or U1431 (N_1431,N_817,N_513);
or U1432 (N_1432,N_621,N_667);
nand U1433 (N_1433,N_586,N_949);
nor U1434 (N_1434,N_997,N_918);
nor U1435 (N_1435,N_628,N_849);
nor U1436 (N_1436,N_641,N_519);
nor U1437 (N_1437,N_766,N_622);
or U1438 (N_1438,N_516,N_515);
nand U1439 (N_1439,N_637,N_626);
nand U1440 (N_1440,N_947,N_751);
or U1441 (N_1441,N_535,N_812);
nor U1442 (N_1442,N_927,N_754);
or U1443 (N_1443,N_758,N_700);
nor U1444 (N_1444,N_664,N_509);
or U1445 (N_1445,N_723,N_977);
nand U1446 (N_1446,N_571,N_731);
or U1447 (N_1447,N_781,N_756);
nor U1448 (N_1448,N_925,N_670);
nand U1449 (N_1449,N_936,N_666);
xor U1450 (N_1450,N_532,N_575);
and U1451 (N_1451,N_679,N_532);
nor U1452 (N_1452,N_504,N_837);
nand U1453 (N_1453,N_857,N_858);
nor U1454 (N_1454,N_508,N_765);
nand U1455 (N_1455,N_843,N_678);
and U1456 (N_1456,N_581,N_684);
or U1457 (N_1457,N_675,N_518);
nor U1458 (N_1458,N_620,N_918);
and U1459 (N_1459,N_772,N_675);
and U1460 (N_1460,N_887,N_950);
and U1461 (N_1461,N_794,N_939);
and U1462 (N_1462,N_958,N_712);
nor U1463 (N_1463,N_566,N_718);
or U1464 (N_1464,N_915,N_949);
and U1465 (N_1465,N_861,N_710);
or U1466 (N_1466,N_978,N_575);
and U1467 (N_1467,N_847,N_981);
nor U1468 (N_1468,N_670,N_826);
and U1469 (N_1469,N_701,N_628);
nor U1470 (N_1470,N_541,N_935);
nor U1471 (N_1471,N_753,N_515);
or U1472 (N_1472,N_645,N_520);
nor U1473 (N_1473,N_877,N_657);
or U1474 (N_1474,N_914,N_927);
or U1475 (N_1475,N_878,N_911);
nor U1476 (N_1476,N_550,N_714);
nor U1477 (N_1477,N_516,N_644);
or U1478 (N_1478,N_785,N_953);
nand U1479 (N_1479,N_526,N_842);
and U1480 (N_1480,N_616,N_753);
and U1481 (N_1481,N_739,N_699);
and U1482 (N_1482,N_944,N_630);
and U1483 (N_1483,N_866,N_638);
nand U1484 (N_1484,N_684,N_811);
nor U1485 (N_1485,N_723,N_633);
and U1486 (N_1486,N_798,N_874);
or U1487 (N_1487,N_834,N_736);
and U1488 (N_1488,N_767,N_590);
nor U1489 (N_1489,N_683,N_500);
and U1490 (N_1490,N_696,N_839);
or U1491 (N_1491,N_980,N_991);
nand U1492 (N_1492,N_721,N_750);
and U1493 (N_1493,N_751,N_979);
nand U1494 (N_1494,N_938,N_869);
or U1495 (N_1495,N_704,N_682);
nor U1496 (N_1496,N_788,N_950);
or U1497 (N_1497,N_580,N_689);
or U1498 (N_1498,N_580,N_621);
and U1499 (N_1499,N_974,N_544);
or U1500 (N_1500,N_1267,N_1160);
nor U1501 (N_1501,N_1100,N_1050);
nor U1502 (N_1502,N_1398,N_1431);
and U1503 (N_1503,N_1009,N_1063);
or U1504 (N_1504,N_1279,N_1020);
nor U1505 (N_1505,N_1459,N_1270);
xor U1506 (N_1506,N_1414,N_1373);
nor U1507 (N_1507,N_1128,N_1147);
nor U1508 (N_1508,N_1011,N_1001);
nor U1509 (N_1509,N_1467,N_1276);
nand U1510 (N_1510,N_1040,N_1323);
and U1511 (N_1511,N_1164,N_1377);
or U1512 (N_1512,N_1318,N_1132);
or U1513 (N_1513,N_1089,N_1444);
or U1514 (N_1514,N_1358,N_1194);
nor U1515 (N_1515,N_1034,N_1419);
or U1516 (N_1516,N_1376,N_1299);
and U1517 (N_1517,N_1479,N_1405);
and U1518 (N_1518,N_1284,N_1145);
and U1519 (N_1519,N_1082,N_1366);
and U1520 (N_1520,N_1314,N_1226);
or U1521 (N_1521,N_1326,N_1411);
and U1522 (N_1522,N_1111,N_1189);
nor U1523 (N_1523,N_1028,N_1057);
or U1524 (N_1524,N_1384,N_1229);
nor U1525 (N_1525,N_1085,N_1105);
nor U1526 (N_1526,N_1409,N_1204);
nor U1527 (N_1527,N_1337,N_1148);
or U1528 (N_1528,N_1367,N_1150);
nor U1529 (N_1529,N_1039,N_1248);
nand U1530 (N_1530,N_1016,N_1492);
or U1531 (N_1531,N_1472,N_1300);
nand U1532 (N_1532,N_1247,N_1106);
and U1533 (N_1533,N_1303,N_1296);
nand U1534 (N_1534,N_1076,N_1362);
nor U1535 (N_1535,N_1493,N_1103);
nor U1536 (N_1536,N_1486,N_1173);
or U1537 (N_1537,N_1309,N_1401);
or U1538 (N_1538,N_1332,N_1192);
nor U1539 (N_1539,N_1213,N_1097);
and U1540 (N_1540,N_1458,N_1096);
nor U1541 (N_1541,N_1046,N_1269);
or U1542 (N_1542,N_1310,N_1048);
xor U1543 (N_1543,N_1363,N_1038);
nor U1544 (N_1544,N_1116,N_1179);
and U1545 (N_1545,N_1348,N_1017);
nand U1546 (N_1546,N_1448,N_1215);
nand U1547 (N_1547,N_1385,N_1455);
nor U1548 (N_1548,N_1088,N_1438);
nand U1549 (N_1549,N_1186,N_1168);
nor U1550 (N_1550,N_1412,N_1005);
xor U1551 (N_1551,N_1102,N_1292);
nor U1552 (N_1552,N_1255,N_1045);
or U1553 (N_1553,N_1465,N_1115);
nor U1554 (N_1554,N_1322,N_1211);
or U1555 (N_1555,N_1361,N_1484);
nand U1556 (N_1556,N_1118,N_1056);
and U1557 (N_1557,N_1101,N_1035);
nand U1558 (N_1558,N_1433,N_1415);
nor U1559 (N_1559,N_1262,N_1054);
nand U1560 (N_1560,N_1131,N_1325);
nand U1561 (N_1561,N_1002,N_1022);
nand U1562 (N_1562,N_1058,N_1202);
or U1563 (N_1563,N_1165,N_1487);
nor U1564 (N_1564,N_1007,N_1346);
or U1565 (N_1565,N_1357,N_1305);
nor U1566 (N_1566,N_1060,N_1268);
and U1567 (N_1567,N_1335,N_1133);
and U1568 (N_1568,N_1290,N_1067);
or U1569 (N_1569,N_1080,N_1266);
or U1570 (N_1570,N_1206,N_1077);
nand U1571 (N_1571,N_1381,N_1475);
nand U1572 (N_1572,N_1393,N_1280);
and U1573 (N_1573,N_1079,N_1339);
or U1574 (N_1574,N_1437,N_1336);
nand U1575 (N_1575,N_1108,N_1264);
nor U1576 (N_1576,N_1157,N_1029);
nor U1577 (N_1577,N_1151,N_1242);
nand U1578 (N_1578,N_1386,N_1081);
or U1579 (N_1579,N_1306,N_1181);
nand U1580 (N_1580,N_1090,N_1349);
and U1581 (N_1581,N_1452,N_1167);
nand U1582 (N_1582,N_1359,N_1187);
or U1583 (N_1583,N_1435,N_1134);
nor U1584 (N_1584,N_1170,N_1199);
or U1585 (N_1585,N_1093,N_1162);
and U1586 (N_1586,N_1117,N_1178);
or U1587 (N_1587,N_1291,N_1354);
and U1588 (N_1588,N_1389,N_1329);
or U1589 (N_1589,N_1338,N_1421);
or U1590 (N_1590,N_1425,N_1109);
and U1591 (N_1591,N_1485,N_1141);
nor U1592 (N_1592,N_1483,N_1169);
nor U1593 (N_1593,N_1104,N_1153);
nand U1594 (N_1594,N_1383,N_1078);
or U1595 (N_1595,N_1478,N_1183);
and U1596 (N_1596,N_1434,N_1087);
nand U1597 (N_1597,N_1480,N_1397);
or U1598 (N_1598,N_1289,N_1023);
nand U1599 (N_1599,N_1124,N_1392);
nand U1600 (N_1600,N_1238,N_1193);
or U1601 (N_1601,N_1466,N_1295);
nor U1602 (N_1602,N_1320,N_1417);
nand U1603 (N_1603,N_1272,N_1094);
nor U1604 (N_1604,N_1008,N_1454);
nor U1605 (N_1605,N_1344,N_1110);
nor U1606 (N_1606,N_1471,N_1043);
nand U1607 (N_1607,N_1227,N_1070);
nor U1608 (N_1608,N_1155,N_1321);
or U1609 (N_1609,N_1390,N_1298);
and U1610 (N_1610,N_1351,N_1368);
nand U1611 (N_1611,N_1031,N_1198);
or U1612 (N_1612,N_1190,N_1423);
nand U1613 (N_1613,N_1429,N_1490);
and U1614 (N_1614,N_1004,N_1473);
and U1615 (N_1615,N_1196,N_1271);
and U1616 (N_1616,N_1312,N_1330);
nor U1617 (N_1617,N_1166,N_1234);
nand U1618 (N_1618,N_1441,N_1136);
or U1619 (N_1619,N_1231,N_1184);
or U1620 (N_1620,N_1282,N_1146);
or U1621 (N_1621,N_1251,N_1180);
nand U1622 (N_1622,N_1442,N_1470);
or U1623 (N_1623,N_1259,N_1071);
or U1624 (N_1624,N_1462,N_1374);
and U1625 (N_1625,N_1388,N_1240);
and U1626 (N_1626,N_1304,N_1174);
and U1627 (N_1627,N_1288,N_1301);
nand U1628 (N_1628,N_1073,N_1083);
nor U1629 (N_1629,N_1084,N_1278);
xor U1630 (N_1630,N_1033,N_1237);
or U1631 (N_1631,N_1218,N_1369);
or U1632 (N_1632,N_1014,N_1225);
and U1633 (N_1633,N_1000,N_1222);
and U1634 (N_1634,N_1203,N_1208);
or U1635 (N_1635,N_1364,N_1175);
nand U1636 (N_1636,N_1123,N_1158);
nand U1637 (N_1637,N_1027,N_1404);
or U1638 (N_1638,N_1285,N_1356);
nor U1639 (N_1639,N_1026,N_1221);
and U1640 (N_1640,N_1399,N_1379);
or U1641 (N_1641,N_1069,N_1460);
or U1642 (N_1642,N_1126,N_1098);
or U1643 (N_1643,N_1313,N_1395);
and U1644 (N_1644,N_1341,N_1408);
and U1645 (N_1645,N_1340,N_1457);
and U1646 (N_1646,N_1129,N_1327);
nor U1647 (N_1647,N_1302,N_1403);
and U1648 (N_1648,N_1059,N_1154);
nor U1649 (N_1649,N_1261,N_1275);
nand U1650 (N_1650,N_1439,N_1396);
nand U1651 (N_1651,N_1443,N_1445);
xor U1652 (N_1652,N_1328,N_1024);
and U1653 (N_1653,N_1311,N_1308);
or U1654 (N_1654,N_1464,N_1477);
and U1655 (N_1655,N_1019,N_1394);
or U1656 (N_1656,N_1372,N_1496);
nor U1657 (N_1657,N_1143,N_1427);
nor U1658 (N_1658,N_1121,N_1049);
nand U1659 (N_1659,N_1201,N_1252);
nor U1660 (N_1660,N_1371,N_1297);
nand U1661 (N_1661,N_1254,N_1382);
nor U1662 (N_1662,N_1161,N_1125);
nand U1663 (N_1663,N_1257,N_1113);
and U1664 (N_1664,N_1307,N_1450);
and U1665 (N_1665,N_1274,N_1068);
or U1666 (N_1666,N_1072,N_1316);
nand U1667 (N_1667,N_1494,N_1406);
and U1668 (N_1668,N_1253,N_1461);
nand U1669 (N_1669,N_1426,N_1319);
nand U1670 (N_1670,N_1220,N_1209);
nand U1671 (N_1671,N_1239,N_1210);
or U1672 (N_1672,N_1378,N_1416);
nor U1673 (N_1673,N_1137,N_1243);
or U1674 (N_1674,N_1498,N_1424);
nor U1675 (N_1675,N_1236,N_1216);
or U1676 (N_1676,N_1065,N_1230);
nor U1677 (N_1677,N_1430,N_1420);
nor U1678 (N_1678,N_1402,N_1232);
and U1679 (N_1679,N_1176,N_1495);
nand U1680 (N_1680,N_1456,N_1256);
nand U1681 (N_1681,N_1013,N_1041);
or U1682 (N_1682,N_1224,N_1171);
nor U1683 (N_1683,N_1061,N_1387);
nand U1684 (N_1684,N_1212,N_1352);
nor U1685 (N_1685,N_1172,N_1112);
xnor U1686 (N_1686,N_1099,N_1315);
and U1687 (N_1687,N_1149,N_1030);
or U1688 (N_1688,N_1142,N_1263);
nand U1689 (N_1689,N_1380,N_1436);
nor U1690 (N_1690,N_1451,N_1066);
nor U1691 (N_1691,N_1249,N_1241);
and U1692 (N_1692,N_1428,N_1260);
or U1693 (N_1693,N_1422,N_1055);
nand U1694 (N_1694,N_1317,N_1407);
or U1695 (N_1695,N_1195,N_1053);
and U1696 (N_1696,N_1114,N_1233);
nor U1697 (N_1697,N_1446,N_1074);
xnor U1698 (N_1698,N_1086,N_1006);
nand U1699 (N_1699,N_1163,N_1036);
nand U1700 (N_1700,N_1075,N_1120);
nand U1701 (N_1701,N_1250,N_1021);
and U1702 (N_1702,N_1092,N_1245);
nor U1703 (N_1703,N_1391,N_1294);
nor U1704 (N_1704,N_1091,N_1499);
nand U1705 (N_1705,N_1122,N_1025);
nor U1706 (N_1706,N_1258,N_1197);
and U1707 (N_1707,N_1214,N_1355);
nor U1708 (N_1708,N_1432,N_1228);
and U1709 (N_1709,N_1334,N_1244);
or U1710 (N_1710,N_1453,N_1476);
and U1711 (N_1711,N_1342,N_1140);
and U1712 (N_1712,N_1156,N_1003);
and U1713 (N_1713,N_1447,N_1217);
nor U1714 (N_1714,N_1345,N_1152);
or U1715 (N_1715,N_1365,N_1144);
and U1716 (N_1716,N_1127,N_1488);
nand U1717 (N_1717,N_1287,N_1497);
and U1718 (N_1718,N_1139,N_1095);
and U1719 (N_1719,N_1463,N_1281);
xor U1720 (N_1720,N_1353,N_1235);
and U1721 (N_1721,N_1413,N_1481);
nand U1722 (N_1722,N_1047,N_1177);
nor U1723 (N_1723,N_1051,N_1469);
nand U1724 (N_1724,N_1037,N_1205);
or U1725 (N_1725,N_1015,N_1489);
nor U1726 (N_1726,N_1343,N_1491);
nor U1727 (N_1727,N_1062,N_1032);
and U1728 (N_1728,N_1277,N_1042);
or U1729 (N_1729,N_1200,N_1360);
and U1730 (N_1730,N_1273,N_1418);
or U1731 (N_1731,N_1350,N_1474);
or U1732 (N_1732,N_1286,N_1449);
nand U1733 (N_1733,N_1246,N_1107);
or U1734 (N_1734,N_1010,N_1468);
or U1735 (N_1735,N_1370,N_1223);
or U1736 (N_1736,N_1119,N_1265);
nand U1737 (N_1737,N_1052,N_1219);
and U1738 (N_1738,N_1410,N_1064);
or U1739 (N_1739,N_1207,N_1188);
and U1740 (N_1740,N_1135,N_1018);
nor U1741 (N_1741,N_1482,N_1331);
or U1742 (N_1742,N_1185,N_1130);
nand U1743 (N_1743,N_1044,N_1347);
and U1744 (N_1744,N_1191,N_1182);
nand U1745 (N_1745,N_1324,N_1283);
nand U1746 (N_1746,N_1138,N_1400);
and U1747 (N_1747,N_1293,N_1159);
or U1748 (N_1748,N_1440,N_1333);
and U1749 (N_1749,N_1012,N_1375);
nand U1750 (N_1750,N_1251,N_1204);
nand U1751 (N_1751,N_1034,N_1345);
xnor U1752 (N_1752,N_1382,N_1095);
and U1753 (N_1753,N_1054,N_1129);
xor U1754 (N_1754,N_1169,N_1136);
or U1755 (N_1755,N_1068,N_1189);
and U1756 (N_1756,N_1371,N_1272);
or U1757 (N_1757,N_1129,N_1275);
and U1758 (N_1758,N_1307,N_1262);
and U1759 (N_1759,N_1119,N_1313);
and U1760 (N_1760,N_1439,N_1422);
and U1761 (N_1761,N_1068,N_1186);
or U1762 (N_1762,N_1104,N_1052);
nand U1763 (N_1763,N_1313,N_1426);
nand U1764 (N_1764,N_1463,N_1197);
and U1765 (N_1765,N_1076,N_1468);
and U1766 (N_1766,N_1331,N_1299);
nor U1767 (N_1767,N_1038,N_1092);
nand U1768 (N_1768,N_1075,N_1233);
and U1769 (N_1769,N_1212,N_1126);
or U1770 (N_1770,N_1161,N_1185);
and U1771 (N_1771,N_1064,N_1205);
nand U1772 (N_1772,N_1149,N_1292);
and U1773 (N_1773,N_1086,N_1105);
nand U1774 (N_1774,N_1475,N_1179);
nor U1775 (N_1775,N_1450,N_1254);
or U1776 (N_1776,N_1483,N_1367);
and U1777 (N_1777,N_1333,N_1313);
nand U1778 (N_1778,N_1221,N_1421);
nor U1779 (N_1779,N_1478,N_1334);
nor U1780 (N_1780,N_1308,N_1062);
nor U1781 (N_1781,N_1278,N_1112);
nor U1782 (N_1782,N_1327,N_1358);
or U1783 (N_1783,N_1225,N_1415);
nor U1784 (N_1784,N_1004,N_1457);
and U1785 (N_1785,N_1286,N_1165);
nand U1786 (N_1786,N_1432,N_1192);
nand U1787 (N_1787,N_1392,N_1254);
nand U1788 (N_1788,N_1187,N_1049);
or U1789 (N_1789,N_1303,N_1480);
or U1790 (N_1790,N_1427,N_1132);
nand U1791 (N_1791,N_1439,N_1076);
nor U1792 (N_1792,N_1190,N_1194);
or U1793 (N_1793,N_1081,N_1178);
xor U1794 (N_1794,N_1303,N_1235);
or U1795 (N_1795,N_1068,N_1402);
or U1796 (N_1796,N_1398,N_1224);
xor U1797 (N_1797,N_1418,N_1082);
nor U1798 (N_1798,N_1486,N_1268);
or U1799 (N_1799,N_1350,N_1194);
nand U1800 (N_1800,N_1030,N_1377);
or U1801 (N_1801,N_1127,N_1039);
nor U1802 (N_1802,N_1394,N_1030);
xor U1803 (N_1803,N_1021,N_1125);
or U1804 (N_1804,N_1220,N_1128);
or U1805 (N_1805,N_1174,N_1295);
nor U1806 (N_1806,N_1198,N_1430);
and U1807 (N_1807,N_1207,N_1292);
or U1808 (N_1808,N_1041,N_1117);
nand U1809 (N_1809,N_1366,N_1123);
or U1810 (N_1810,N_1107,N_1393);
nand U1811 (N_1811,N_1218,N_1434);
nand U1812 (N_1812,N_1252,N_1392);
or U1813 (N_1813,N_1174,N_1231);
or U1814 (N_1814,N_1336,N_1188);
nor U1815 (N_1815,N_1495,N_1344);
or U1816 (N_1816,N_1462,N_1015);
xor U1817 (N_1817,N_1005,N_1309);
nor U1818 (N_1818,N_1169,N_1231);
or U1819 (N_1819,N_1457,N_1078);
nor U1820 (N_1820,N_1343,N_1087);
or U1821 (N_1821,N_1372,N_1134);
and U1822 (N_1822,N_1063,N_1118);
or U1823 (N_1823,N_1015,N_1292);
or U1824 (N_1824,N_1261,N_1076);
nor U1825 (N_1825,N_1303,N_1174);
nand U1826 (N_1826,N_1297,N_1130);
and U1827 (N_1827,N_1090,N_1084);
or U1828 (N_1828,N_1055,N_1125);
or U1829 (N_1829,N_1326,N_1116);
nor U1830 (N_1830,N_1034,N_1279);
or U1831 (N_1831,N_1446,N_1212);
nand U1832 (N_1832,N_1273,N_1258);
and U1833 (N_1833,N_1301,N_1233);
or U1834 (N_1834,N_1208,N_1058);
nand U1835 (N_1835,N_1228,N_1406);
or U1836 (N_1836,N_1279,N_1026);
nor U1837 (N_1837,N_1334,N_1177);
nor U1838 (N_1838,N_1340,N_1171);
and U1839 (N_1839,N_1487,N_1191);
nand U1840 (N_1840,N_1052,N_1176);
and U1841 (N_1841,N_1219,N_1499);
or U1842 (N_1842,N_1205,N_1326);
and U1843 (N_1843,N_1178,N_1015);
nor U1844 (N_1844,N_1431,N_1022);
nor U1845 (N_1845,N_1299,N_1272);
and U1846 (N_1846,N_1352,N_1277);
and U1847 (N_1847,N_1412,N_1041);
and U1848 (N_1848,N_1277,N_1349);
nor U1849 (N_1849,N_1298,N_1377);
nor U1850 (N_1850,N_1068,N_1282);
and U1851 (N_1851,N_1368,N_1360);
or U1852 (N_1852,N_1099,N_1000);
nand U1853 (N_1853,N_1364,N_1035);
nor U1854 (N_1854,N_1474,N_1170);
nor U1855 (N_1855,N_1077,N_1191);
nor U1856 (N_1856,N_1237,N_1310);
nor U1857 (N_1857,N_1405,N_1135);
nor U1858 (N_1858,N_1230,N_1382);
nor U1859 (N_1859,N_1220,N_1368);
and U1860 (N_1860,N_1173,N_1413);
or U1861 (N_1861,N_1445,N_1377);
nor U1862 (N_1862,N_1026,N_1042);
nor U1863 (N_1863,N_1329,N_1044);
and U1864 (N_1864,N_1444,N_1461);
nand U1865 (N_1865,N_1395,N_1079);
and U1866 (N_1866,N_1228,N_1167);
nor U1867 (N_1867,N_1150,N_1321);
and U1868 (N_1868,N_1247,N_1028);
nand U1869 (N_1869,N_1423,N_1477);
nor U1870 (N_1870,N_1058,N_1313);
and U1871 (N_1871,N_1262,N_1023);
nand U1872 (N_1872,N_1178,N_1310);
xnor U1873 (N_1873,N_1257,N_1186);
or U1874 (N_1874,N_1255,N_1446);
or U1875 (N_1875,N_1013,N_1047);
xor U1876 (N_1876,N_1298,N_1408);
nand U1877 (N_1877,N_1196,N_1337);
nand U1878 (N_1878,N_1182,N_1184);
and U1879 (N_1879,N_1207,N_1083);
nand U1880 (N_1880,N_1442,N_1014);
and U1881 (N_1881,N_1360,N_1492);
nor U1882 (N_1882,N_1463,N_1004);
nor U1883 (N_1883,N_1114,N_1401);
and U1884 (N_1884,N_1146,N_1039);
and U1885 (N_1885,N_1052,N_1334);
and U1886 (N_1886,N_1479,N_1155);
and U1887 (N_1887,N_1070,N_1100);
xnor U1888 (N_1888,N_1086,N_1429);
nor U1889 (N_1889,N_1480,N_1212);
or U1890 (N_1890,N_1298,N_1366);
or U1891 (N_1891,N_1150,N_1441);
or U1892 (N_1892,N_1313,N_1397);
nor U1893 (N_1893,N_1308,N_1342);
nand U1894 (N_1894,N_1116,N_1469);
and U1895 (N_1895,N_1351,N_1141);
or U1896 (N_1896,N_1281,N_1016);
nor U1897 (N_1897,N_1277,N_1106);
and U1898 (N_1898,N_1199,N_1077);
nand U1899 (N_1899,N_1104,N_1446);
xor U1900 (N_1900,N_1117,N_1060);
and U1901 (N_1901,N_1413,N_1039);
nor U1902 (N_1902,N_1051,N_1015);
nand U1903 (N_1903,N_1294,N_1224);
and U1904 (N_1904,N_1071,N_1411);
nand U1905 (N_1905,N_1219,N_1469);
and U1906 (N_1906,N_1031,N_1235);
or U1907 (N_1907,N_1061,N_1444);
and U1908 (N_1908,N_1026,N_1183);
or U1909 (N_1909,N_1318,N_1235);
and U1910 (N_1910,N_1249,N_1200);
or U1911 (N_1911,N_1464,N_1117);
nand U1912 (N_1912,N_1288,N_1429);
nand U1913 (N_1913,N_1332,N_1017);
and U1914 (N_1914,N_1434,N_1255);
or U1915 (N_1915,N_1474,N_1478);
nor U1916 (N_1916,N_1478,N_1139);
and U1917 (N_1917,N_1060,N_1288);
nor U1918 (N_1918,N_1290,N_1097);
and U1919 (N_1919,N_1182,N_1232);
nor U1920 (N_1920,N_1101,N_1048);
nor U1921 (N_1921,N_1457,N_1237);
nand U1922 (N_1922,N_1066,N_1043);
and U1923 (N_1923,N_1239,N_1195);
nor U1924 (N_1924,N_1178,N_1283);
or U1925 (N_1925,N_1382,N_1435);
or U1926 (N_1926,N_1466,N_1353);
or U1927 (N_1927,N_1026,N_1490);
nand U1928 (N_1928,N_1411,N_1291);
or U1929 (N_1929,N_1010,N_1153);
or U1930 (N_1930,N_1408,N_1380);
or U1931 (N_1931,N_1430,N_1403);
xnor U1932 (N_1932,N_1030,N_1427);
nand U1933 (N_1933,N_1374,N_1132);
and U1934 (N_1934,N_1096,N_1273);
nor U1935 (N_1935,N_1152,N_1008);
nand U1936 (N_1936,N_1136,N_1295);
and U1937 (N_1937,N_1482,N_1491);
nor U1938 (N_1938,N_1080,N_1465);
nand U1939 (N_1939,N_1232,N_1436);
nor U1940 (N_1940,N_1150,N_1247);
nor U1941 (N_1941,N_1493,N_1193);
nand U1942 (N_1942,N_1107,N_1102);
nand U1943 (N_1943,N_1489,N_1080);
or U1944 (N_1944,N_1477,N_1232);
or U1945 (N_1945,N_1418,N_1211);
nand U1946 (N_1946,N_1076,N_1096);
or U1947 (N_1947,N_1411,N_1226);
or U1948 (N_1948,N_1170,N_1488);
nand U1949 (N_1949,N_1035,N_1048);
nand U1950 (N_1950,N_1319,N_1272);
nor U1951 (N_1951,N_1313,N_1402);
nor U1952 (N_1952,N_1080,N_1066);
nor U1953 (N_1953,N_1205,N_1136);
nor U1954 (N_1954,N_1332,N_1173);
and U1955 (N_1955,N_1256,N_1434);
nor U1956 (N_1956,N_1035,N_1472);
nand U1957 (N_1957,N_1320,N_1159);
nand U1958 (N_1958,N_1296,N_1188);
nor U1959 (N_1959,N_1113,N_1473);
and U1960 (N_1960,N_1164,N_1121);
or U1961 (N_1961,N_1285,N_1203);
or U1962 (N_1962,N_1332,N_1244);
xor U1963 (N_1963,N_1368,N_1013);
nand U1964 (N_1964,N_1014,N_1171);
or U1965 (N_1965,N_1475,N_1291);
xnor U1966 (N_1966,N_1041,N_1406);
or U1967 (N_1967,N_1204,N_1126);
nor U1968 (N_1968,N_1270,N_1050);
or U1969 (N_1969,N_1304,N_1385);
and U1970 (N_1970,N_1076,N_1395);
nand U1971 (N_1971,N_1247,N_1135);
nor U1972 (N_1972,N_1270,N_1205);
and U1973 (N_1973,N_1206,N_1203);
nand U1974 (N_1974,N_1240,N_1013);
and U1975 (N_1975,N_1446,N_1078);
and U1976 (N_1976,N_1030,N_1433);
nor U1977 (N_1977,N_1313,N_1362);
or U1978 (N_1978,N_1396,N_1347);
nor U1979 (N_1979,N_1452,N_1109);
nor U1980 (N_1980,N_1061,N_1239);
and U1981 (N_1981,N_1220,N_1373);
and U1982 (N_1982,N_1160,N_1419);
and U1983 (N_1983,N_1440,N_1234);
xor U1984 (N_1984,N_1043,N_1287);
and U1985 (N_1985,N_1477,N_1009);
and U1986 (N_1986,N_1004,N_1461);
and U1987 (N_1987,N_1052,N_1108);
and U1988 (N_1988,N_1443,N_1075);
and U1989 (N_1989,N_1441,N_1113);
and U1990 (N_1990,N_1446,N_1109);
or U1991 (N_1991,N_1375,N_1286);
and U1992 (N_1992,N_1167,N_1030);
or U1993 (N_1993,N_1135,N_1146);
and U1994 (N_1994,N_1408,N_1129);
nand U1995 (N_1995,N_1016,N_1396);
and U1996 (N_1996,N_1407,N_1393);
nor U1997 (N_1997,N_1002,N_1392);
nand U1998 (N_1998,N_1149,N_1456);
nor U1999 (N_1999,N_1374,N_1003);
nor U2000 (N_2000,N_1971,N_1580);
and U2001 (N_2001,N_1575,N_1646);
or U2002 (N_2002,N_1810,N_1742);
and U2003 (N_2003,N_1788,N_1609);
or U2004 (N_2004,N_1531,N_1914);
and U2005 (N_2005,N_1639,N_1841);
and U2006 (N_2006,N_1756,N_1899);
or U2007 (N_2007,N_1940,N_1809);
nand U2008 (N_2008,N_1607,N_1709);
or U2009 (N_2009,N_1708,N_1731);
nand U2010 (N_2010,N_1791,N_1994);
or U2011 (N_2011,N_1564,N_1988);
or U2012 (N_2012,N_1986,N_1864);
nand U2013 (N_2013,N_1855,N_1659);
and U2014 (N_2014,N_1856,N_1908);
nand U2015 (N_2015,N_1683,N_1510);
nor U2016 (N_2016,N_1770,N_1904);
nand U2017 (N_2017,N_1823,N_1502);
or U2018 (N_2018,N_1910,N_1506);
nor U2019 (N_2019,N_1858,N_1740);
nand U2020 (N_2020,N_1789,N_1888);
or U2021 (N_2021,N_1640,N_1549);
or U2022 (N_2022,N_1625,N_1577);
nor U2023 (N_2023,N_1642,N_1633);
and U2024 (N_2024,N_1542,N_1630);
and U2025 (N_2025,N_1964,N_1569);
nand U2026 (N_2026,N_1634,N_1777);
nor U2027 (N_2027,N_1974,N_1931);
or U2028 (N_2028,N_1557,N_1952);
or U2029 (N_2029,N_1892,N_1738);
and U2030 (N_2030,N_1776,N_1728);
or U2031 (N_2031,N_1932,N_1887);
nand U2032 (N_2032,N_1690,N_1758);
and U2033 (N_2033,N_1675,N_1648);
or U2034 (N_2034,N_1890,N_1845);
xnor U2035 (N_2035,N_1806,N_1893);
and U2036 (N_2036,N_1949,N_1915);
or U2037 (N_2037,N_1583,N_1837);
nand U2038 (N_2038,N_1741,N_1539);
nor U2039 (N_2039,N_1563,N_1520);
and U2040 (N_2040,N_1925,N_1647);
xor U2041 (N_2041,N_1980,N_1627);
or U2042 (N_2042,N_1905,N_1840);
or U2043 (N_2043,N_1733,N_1500);
nand U2044 (N_2044,N_1853,N_1713);
nor U2045 (N_2045,N_1956,N_1702);
and U2046 (N_2046,N_1934,N_1787);
nor U2047 (N_2047,N_1727,N_1793);
and U2048 (N_2048,N_1821,N_1763);
and U2049 (N_2049,N_1796,N_1800);
nor U2050 (N_2050,N_1969,N_1595);
nor U2051 (N_2051,N_1803,N_1505);
nor U2052 (N_2052,N_1778,N_1814);
nor U2053 (N_2053,N_1857,N_1848);
or U2054 (N_2054,N_1521,N_1735);
nand U2055 (N_2055,N_1678,N_1963);
or U2056 (N_2056,N_1573,N_1541);
nor U2057 (N_2057,N_1977,N_1743);
nand U2058 (N_2058,N_1918,N_1732);
and U2059 (N_2059,N_1978,N_1873);
or U2060 (N_2060,N_1551,N_1571);
nor U2061 (N_2061,N_1818,N_1903);
and U2062 (N_2062,N_1984,N_1671);
or U2063 (N_2063,N_1779,N_1680);
or U2064 (N_2064,N_1698,N_1661);
or U2065 (N_2065,N_1783,N_1859);
nand U2066 (N_2066,N_1817,N_1773);
nand U2067 (N_2067,N_1649,N_1926);
and U2068 (N_2068,N_1975,N_1826);
and U2069 (N_2069,N_1699,N_1656);
nor U2070 (N_2070,N_1507,N_1920);
and U2071 (N_2071,N_1697,N_1704);
nor U2072 (N_2072,N_1979,N_1513);
nand U2073 (N_2073,N_1771,N_1517);
nor U2074 (N_2074,N_1759,N_1871);
and U2075 (N_2075,N_1812,N_1665);
or U2076 (N_2076,N_1679,N_1650);
nor U2077 (N_2077,N_1852,N_1916);
nor U2078 (N_2078,N_1691,N_1847);
nand U2079 (N_2079,N_1533,N_1881);
and U2080 (N_2080,N_1839,N_1987);
nor U2081 (N_2081,N_1538,N_1598);
nor U2082 (N_2082,N_1955,N_1559);
nand U2083 (N_2083,N_1842,N_1604);
nand U2084 (N_2084,N_1550,N_1958);
nor U2085 (N_2085,N_1961,N_1568);
and U2086 (N_2086,N_1667,N_1862);
or U2087 (N_2087,N_1938,N_1747);
nand U2088 (N_2088,N_1976,N_1991);
nand U2089 (N_2089,N_1902,N_1636);
and U2090 (N_2090,N_1626,N_1749);
and U2091 (N_2091,N_1898,N_1816);
and U2092 (N_2092,N_1947,N_1637);
and U2093 (N_2093,N_1957,N_1901);
nand U2094 (N_2094,N_1906,N_1614);
or U2095 (N_2095,N_1965,N_1825);
nand U2096 (N_2096,N_1596,N_1819);
or U2097 (N_2097,N_1951,N_1886);
or U2098 (N_2098,N_1681,N_1561);
xor U2099 (N_2099,N_1725,N_1673);
or U2100 (N_2100,N_1767,N_1772);
or U2101 (N_2101,N_1532,N_1616);
nand U2102 (N_2102,N_1919,N_1993);
nand U2103 (N_2103,N_1572,N_1566);
or U2104 (N_2104,N_1757,N_1959);
nor U2105 (N_2105,N_1827,N_1799);
and U2106 (N_2106,N_1754,N_1768);
or U2107 (N_2107,N_1913,N_1555);
or U2108 (N_2108,N_1643,N_1982);
nor U2109 (N_2109,N_1548,N_1843);
nand U2110 (N_2110,N_1526,N_1879);
or U2111 (N_2111,N_1654,N_1597);
and U2112 (N_2112,N_1820,N_1652);
and U2113 (N_2113,N_1950,N_1981);
or U2114 (N_2114,N_1589,N_1612);
nor U2115 (N_2115,N_1835,N_1894);
and U2116 (N_2116,N_1601,N_1792);
nor U2117 (N_2117,N_1524,N_1522);
or U2118 (N_2118,N_1953,N_1701);
or U2119 (N_2119,N_1501,N_1734);
and U2120 (N_2120,N_1752,N_1664);
nor U2121 (N_2121,N_1628,N_1782);
or U2122 (N_2122,N_1865,N_1882);
nand U2123 (N_2123,N_1594,N_1726);
and U2124 (N_2124,N_1765,N_1670);
nor U2125 (N_2125,N_1606,N_1874);
or U2126 (N_2126,N_1570,N_1605);
nand U2127 (N_2127,N_1935,N_1578);
or U2128 (N_2128,N_1795,N_1794);
nand U2129 (N_2129,N_1784,N_1813);
nand U2130 (N_2130,N_1895,N_1774);
nand U2131 (N_2131,N_1751,N_1515);
nand U2132 (N_2132,N_1942,N_1868);
nor U2133 (N_2133,N_1536,N_1860);
nand U2134 (N_2134,N_1719,N_1828);
nand U2135 (N_2135,N_1721,N_1884);
nand U2136 (N_2136,N_1831,N_1644);
and U2137 (N_2137,N_1534,N_1944);
or U2138 (N_2138,N_1824,N_1924);
or U2139 (N_2139,N_1775,N_1880);
nand U2140 (N_2140,N_1618,N_1875);
xnor U2141 (N_2141,N_1807,N_1599);
nor U2142 (N_2142,N_1585,N_1929);
nor U2143 (N_2143,N_1897,N_1834);
nor U2144 (N_2144,N_1836,N_1900);
or U2145 (N_2145,N_1543,N_1736);
or U2146 (N_2146,N_1685,N_1737);
and U2147 (N_2147,N_1877,N_1937);
xor U2148 (N_2148,N_1832,N_1863);
nand U2149 (N_2149,N_1870,N_1707);
nor U2150 (N_2150,N_1948,N_1540);
nor U2151 (N_2151,N_1554,N_1682);
or U2152 (N_2152,N_1686,N_1562);
nand U2153 (N_2153,N_1694,N_1503);
or U2154 (N_2154,N_1622,N_1602);
nor U2155 (N_2155,N_1655,N_1801);
and U2156 (N_2156,N_1593,N_1833);
nor U2157 (N_2157,N_1651,N_1808);
or U2158 (N_2158,N_1576,N_1907);
nand U2159 (N_2159,N_1624,N_1687);
nor U2160 (N_2160,N_1968,N_1781);
nor U2161 (N_2161,N_1802,N_1723);
or U2162 (N_2162,N_1769,N_1629);
and U2163 (N_2163,N_1545,N_1621);
nor U2164 (N_2164,N_1567,N_1527);
and U2165 (N_2165,N_1672,N_1590);
nor U2166 (N_2166,N_1844,N_1620);
nor U2167 (N_2167,N_1669,N_1973);
or U2168 (N_2168,N_1552,N_1512);
nand U2169 (N_2169,N_1983,N_1535);
and U2170 (N_2170,N_1525,N_1547);
nand U2171 (N_2171,N_1565,N_1850);
or U2172 (N_2172,N_1706,N_1668);
nand U2173 (N_2173,N_1941,N_1703);
nand U2174 (N_2174,N_1528,N_1511);
nand U2175 (N_2175,N_1936,N_1876);
nor U2176 (N_2176,N_1608,N_1861);
nand U2177 (N_2177,N_1967,N_1762);
or U2178 (N_2178,N_1786,N_1996);
or U2179 (N_2179,N_1730,N_1750);
nand U2180 (N_2180,N_1692,N_1746);
nor U2181 (N_2181,N_1954,N_1966);
nor U2182 (N_2182,N_1558,N_1574);
nand U2183 (N_2183,N_1815,N_1748);
nor U2184 (N_2184,N_1912,N_1544);
or U2185 (N_2185,N_1700,N_1927);
nand U2186 (N_2186,N_1523,N_1529);
nand U2187 (N_2187,N_1946,N_1600);
nand U2188 (N_2188,N_1998,N_1739);
nand U2189 (N_2189,N_1588,N_1645);
or U2190 (N_2190,N_1970,N_1923);
or U2191 (N_2191,N_1867,N_1885);
or U2192 (N_2192,N_1712,N_1695);
nor U2193 (N_2193,N_1849,N_1693);
and U2194 (N_2194,N_1560,N_1760);
or U2195 (N_2195,N_1761,N_1720);
nor U2196 (N_2196,N_1846,N_1917);
and U2197 (N_2197,N_1657,N_1689);
or U2198 (N_2198,N_1985,N_1744);
and U2199 (N_2199,N_1745,N_1660);
nand U2200 (N_2200,N_1790,N_1995);
or U2201 (N_2201,N_1688,N_1933);
nand U2202 (N_2202,N_1638,N_1530);
nor U2203 (N_2203,N_1753,N_1714);
nor U2204 (N_2204,N_1623,N_1546);
and U2205 (N_2205,N_1592,N_1990);
nor U2206 (N_2206,N_1891,N_1508);
or U2207 (N_2207,N_1684,N_1504);
and U2208 (N_2208,N_1921,N_1509);
nand U2209 (N_2209,N_1676,N_1653);
and U2210 (N_2210,N_1909,N_1711);
and U2211 (N_2211,N_1514,N_1872);
nand U2212 (N_2212,N_1613,N_1663);
nand U2213 (N_2213,N_1632,N_1716);
or U2214 (N_2214,N_1610,N_1537);
nor U2215 (N_2215,N_1989,N_1805);
nand U2216 (N_2216,N_1715,N_1724);
nand U2217 (N_2217,N_1960,N_1943);
xnor U2218 (N_2218,N_1635,N_1677);
nand U2219 (N_2219,N_1717,N_1641);
nor U2220 (N_2220,N_1718,N_1911);
nor U2221 (N_2221,N_1516,N_1556);
nor U2222 (N_2222,N_1586,N_1666);
nor U2223 (N_2223,N_1945,N_1822);
or U2224 (N_2224,N_1780,N_1587);
or U2225 (N_2225,N_1939,N_1785);
nor U2226 (N_2226,N_1851,N_1922);
nand U2227 (N_2227,N_1611,N_1928);
nand U2228 (N_2228,N_1518,N_1992);
and U2229 (N_2229,N_1705,N_1999);
and U2230 (N_2230,N_1658,N_1674);
nand U2231 (N_2231,N_1962,N_1617);
xnor U2232 (N_2232,N_1811,N_1755);
or U2233 (N_2233,N_1603,N_1883);
nand U2234 (N_2234,N_1866,N_1619);
nand U2235 (N_2235,N_1930,N_1729);
or U2236 (N_2236,N_1696,N_1582);
nand U2237 (N_2237,N_1889,N_1710);
nand U2238 (N_2238,N_1878,N_1764);
and U2239 (N_2239,N_1662,N_1579);
nor U2240 (N_2240,N_1972,N_1631);
nand U2241 (N_2241,N_1896,N_1798);
and U2242 (N_2242,N_1722,N_1581);
xnor U2243 (N_2243,N_1553,N_1854);
nand U2244 (N_2244,N_1829,N_1766);
or U2245 (N_2245,N_1519,N_1591);
or U2246 (N_2246,N_1584,N_1830);
nand U2247 (N_2247,N_1797,N_1838);
and U2248 (N_2248,N_1997,N_1804);
and U2249 (N_2249,N_1615,N_1869);
or U2250 (N_2250,N_1757,N_1756);
and U2251 (N_2251,N_1859,N_1748);
nand U2252 (N_2252,N_1866,N_1727);
and U2253 (N_2253,N_1894,N_1614);
nand U2254 (N_2254,N_1515,N_1976);
or U2255 (N_2255,N_1520,N_1571);
or U2256 (N_2256,N_1693,N_1923);
and U2257 (N_2257,N_1799,N_1592);
or U2258 (N_2258,N_1832,N_1536);
nand U2259 (N_2259,N_1841,N_1877);
xnor U2260 (N_2260,N_1643,N_1854);
nor U2261 (N_2261,N_1858,N_1668);
and U2262 (N_2262,N_1679,N_1670);
nand U2263 (N_2263,N_1596,N_1640);
nor U2264 (N_2264,N_1748,N_1864);
nor U2265 (N_2265,N_1821,N_1927);
and U2266 (N_2266,N_1655,N_1797);
nand U2267 (N_2267,N_1908,N_1793);
and U2268 (N_2268,N_1746,N_1585);
nor U2269 (N_2269,N_1654,N_1825);
nor U2270 (N_2270,N_1897,N_1850);
nor U2271 (N_2271,N_1755,N_1753);
nand U2272 (N_2272,N_1876,N_1955);
nand U2273 (N_2273,N_1948,N_1959);
nor U2274 (N_2274,N_1837,N_1812);
nand U2275 (N_2275,N_1806,N_1779);
and U2276 (N_2276,N_1958,N_1981);
or U2277 (N_2277,N_1520,N_1813);
nand U2278 (N_2278,N_1729,N_1867);
nand U2279 (N_2279,N_1702,N_1962);
nand U2280 (N_2280,N_1755,N_1946);
or U2281 (N_2281,N_1785,N_1642);
nand U2282 (N_2282,N_1975,N_1815);
and U2283 (N_2283,N_1711,N_1609);
and U2284 (N_2284,N_1635,N_1662);
and U2285 (N_2285,N_1962,N_1628);
or U2286 (N_2286,N_1723,N_1524);
and U2287 (N_2287,N_1826,N_1737);
or U2288 (N_2288,N_1744,N_1523);
or U2289 (N_2289,N_1643,N_1501);
or U2290 (N_2290,N_1541,N_1707);
and U2291 (N_2291,N_1735,N_1625);
and U2292 (N_2292,N_1703,N_1804);
and U2293 (N_2293,N_1563,N_1860);
or U2294 (N_2294,N_1924,N_1985);
nor U2295 (N_2295,N_1947,N_1677);
nor U2296 (N_2296,N_1570,N_1620);
or U2297 (N_2297,N_1784,N_1904);
nand U2298 (N_2298,N_1538,N_1629);
nand U2299 (N_2299,N_1815,N_1901);
and U2300 (N_2300,N_1744,N_1729);
and U2301 (N_2301,N_1545,N_1731);
or U2302 (N_2302,N_1953,N_1580);
nor U2303 (N_2303,N_1788,N_1913);
and U2304 (N_2304,N_1726,N_1761);
nor U2305 (N_2305,N_1546,N_1666);
and U2306 (N_2306,N_1814,N_1938);
nand U2307 (N_2307,N_1538,N_1924);
or U2308 (N_2308,N_1969,N_1779);
nor U2309 (N_2309,N_1831,N_1814);
nand U2310 (N_2310,N_1575,N_1584);
nor U2311 (N_2311,N_1885,N_1921);
nor U2312 (N_2312,N_1854,N_1674);
nand U2313 (N_2313,N_1566,N_1887);
nor U2314 (N_2314,N_1805,N_1591);
nand U2315 (N_2315,N_1984,N_1501);
or U2316 (N_2316,N_1991,N_1602);
nor U2317 (N_2317,N_1745,N_1967);
nor U2318 (N_2318,N_1878,N_1884);
nor U2319 (N_2319,N_1756,N_1683);
and U2320 (N_2320,N_1848,N_1546);
and U2321 (N_2321,N_1772,N_1953);
and U2322 (N_2322,N_1892,N_1599);
nand U2323 (N_2323,N_1751,N_1537);
and U2324 (N_2324,N_1594,N_1970);
xnor U2325 (N_2325,N_1792,N_1731);
nor U2326 (N_2326,N_1626,N_1964);
and U2327 (N_2327,N_1619,N_1983);
and U2328 (N_2328,N_1681,N_1565);
nand U2329 (N_2329,N_1849,N_1559);
or U2330 (N_2330,N_1521,N_1928);
and U2331 (N_2331,N_1539,N_1846);
nor U2332 (N_2332,N_1552,N_1694);
nor U2333 (N_2333,N_1524,N_1951);
and U2334 (N_2334,N_1697,N_1571);
and U2335 (N_2335,N_1770,N_1521);
or U2336 (N_2336,N_1519,N_1886);
nor U2337 (N_2337,N_1735,N_1645);
nand U2338 (N_2338,N_1725,N_1873);
or U2339 (N_2339,N_1929,N_1663);
nand U2340 (N_2340,N_1872,N_1679);
nor U2341 (N_2341,N_1610,N_1796);
nand U2342 (N_2342,N_1765,N_1961);
and U2343 (N_2343,N_1893,N_1540);
nand U2344 (N_2344,N_1612,N_1812);
or U2345 (N_2345,N_1699,N_1906);
nor U2346 (N_2346,N_1519,N_1806);
nand U2347 (N_2347,N_1564,N_1740);
and U2348 (N_2348,N_1572,N_1511);
and U2349 (N_2349,N_1937,N_1550);
or U2350 (N_2350,N_1501,N_1887);
or U2351 (N_2351,N_1572,N_1670);
nor U2352 (N_2352,N_1557,N_1731);
and U2353 (N_2353,N_1969,N_1986);
and U2354 (N_2354,N_1748,N_1871);
and U2355 (N_2355,N_1662,N_1861);
nand U2356 (N_2356,N_1908,N_1620);
nand U2357 (N_2357,N_1727,N_1578);
nand U2358 (N_2358,N_1960,N_1645);
or U2359 (N_2359,N_1608,N_1652);
nand U2360 (N_2360,N_1947,N_1706);
or U2361 (N_2361,N_1549,N_1987);
or U2362 (N_2362,N_1954,N_1684);
or U2363 (N_2363,N_1779,N_1717);
nand U2364 (N_2364,N_1913,N_1579);
nor U2365 (N_2365,N_1676,N_1717);
nand U2366 (N_2366,N_1818,N_1923);
nand U2367 (N_2367,N_1595,N_1697);
nor U2368 (N_2368,N_1538,N_1543);
nor U2369 (N_2369,N_1810,N_1632);
nand U2370 (N_2370,N_1814,N_1999);
and U2371 (N_2371,N_1785,N_1623);
or U2372 (N_2372,N_1785,N_1651);
nand U2373 (N_2373,N_1675,N_1532);
nor U2374 (N_2374,N_1602,N_1954);
or U2375 (N_2375,N_1744,N_1849);
nand U2376 (N_2376,N_1561,N_1626);
nor U2377 (N_2377,N_1780,N_1948);
nor U2378 (N_2378,N_1650,N_1652);
xor U2379 (N_2379,N_1876,N_1916);
and U2380 (N_2380,N_1859,N_1880);
and U2381 (N_2381,N_1670,N_1543);
nor U2382 (N_2382,N_1702,N_1723);
xor U2383 (N_2383,N_1953,N_1951);
nor U2384 (N_2384,N_1679,N_1850);
and U2385 (N_2385,N_1670,N_1618);
and U2386 (N_2386,N_1551,N_1635);
nand U2387 (N_2387,N_1946,N_1779);
or U2388 (N_2388,N_1986,N_1638);
nor U2389 (N_2389,N_1512,N_1568);
or U2390 (N_2390,N_1913,N_1848);
and U2391 (N_2391,N_1838,N_1643);
nor U2392 (N_2392,N_1559,N_1609);
nor U2393 (N_2393,N_1746,N_1661);
nor U2394 (N_2394,N_1586,N_1776);
nand U2395 (N_2395,N_1842,N_1613);
nand U2396 (N_2396,N_1700,N_1682);
and U2397 (N_2397,N_1888,N_1802);
nand U2398 (N_2398,N_1595,N_1668);
nand U2399 (N_2399,N_1852,N_1932);
or U2400 (N_2400,N_1580,N_1662);
and U2401 (N_2401,N_1923,N_1524);
or U2402 (N_2402,N_1632,N_1617);
and U2403 (N_2403,N_1654,N_1601);
or U2404 (N_2404,N_1590,N_1577);
or U2405 (N_2405,N_1802,N_1686);
nand U2406 (N_2406,N_1566,N_1917);
nand U2407 (N_2407,N_1520,N_1889);
nor U2408 (N_2408,N_1590,N_1549);
xnor U2409 (N_2409,N_1658,N_1511);
and U2410 (N_2410,N_1614,N_1895);
and U2411 (N_2411,N_1806,N_1822);
nor U2412 (N_2412,N_1702,N_1909);
nor U2413 (N_2413,N_1793,N_1910);
or U2414 (N_2414,N_1805,N_1847);
nor U2415 (N_2415,N_1678,N_1795);
or U2416 (N_2416,N_1570,N_1831);
and U2417 (N_2417,N_1949,N_1878);
nor U2418 (N_2418,N_1823,N_1730);
and U2419 (N_2419,N_1943,N_1887);
nand U2420 (N_2420,N_1895,N_1735);
or U2421 (N_2421,N_1633,N_1752);
and U2422 (N_2422,N_1931,N_1508);
nor U2423 (N_2423,N_1500,N_1912);
nor U2424 (N_2424,N_1584,N_1566);
or U2425 (N_2425,N_1657,N_1557);
nor U2426 (N_2426,N_1813,N_1818);
and U2427 (N_2427,N_1852,N_1649);
nor U2428 (N_2428,N_1928,N_1858);
nor U2429 (N_2429,N_1593,N_1944);
or U2430 (N_2430,N_1816,N_1786);
and U2431 (N_2431,N_1671,N_1580);
nor U2432 (N_2432,N_1582,N_1505);
nand U2433 (N_2433,N_1630,N_1693);
nor U2434 (N_2434,N_1601,N_1715);
nor U2435 (N_2435,N_1651,N_1813);
nor U2436 (N_2436,N_1515,N_1880);
xnor U2437 (N_2437,N_1610,N_1550);
nand U2438 (N_2438,N_1588,N_1838);
nor U2439 (N_2439,N_1686,N_1964);
and U2440 (N_2440,N_1913,N_1959);
or U2441 (N_2441,N_1754,N_1765);
or U2442 (N_2442,N_1916,N_1541);
xor U2443 (N_2443,N_1861,N_1738);
and U2444 (N_2444,N_1566,N_1862);
nand U2445 (N_2445,N_1554,N_1594);
nand U2446 (N_2446,N_1708,N_1517);
nor U2447 (N_2447,N_1600,N_1655);
nor U2448 (N_2448,N_1747,N_1695);
nand U2449 (N_2449,N_1511,N_1762);
or U2450 (N_2450,N_1729,N_1844);
and U2451 (N_2451,N_1922,N_1540);
nand U2452 (N_2452,N_1580,N_1526);
or U2453 (N_2453,N_1836,N_1558);
nand U2454 (N_2454,N_1647,N_1832);
or U2455 (N_2455,N_1642,N_1646);
and U2456 (N_2456,N_1740,N_1762);
nand U2457 (N_2457,N_1521,N_1844);
or U2458 (N_2458,N_1580,N_1831);
nand U2459 (N_2459,N_1755,N_1919);
or U2460 (N_2460,N_1878,N_1639);
and U2461 (N_2461,N_1551,N_1567);
xor U2462 (N_2462,N_1707,N_1974);
nand U2463 (N_2463,N_1506,N_1723);
and U2464 (N_2464,N_1902,N_1931);
and U2465 (N_2465,N_1760,N_1603);
nand U2466 (N_2466,N_1661,N_1976);
nor U2467 (N_2467,N_1563,N_1665);
and U2468 (N_2468,N_1635,N_1817);
and U2469 (N_2469,N_1740,N_1919);
nor U2470 (N_2470,N_1729,N_1570);
nor U2471 (N_2471,N_1521,N_1685);
nor U2472 (N_2472,N_1552,N_1744);
and U2473 (N_2473,N_1687,N_1672);
and U2474 (N_2474,N_1705,N_1514);
or U2475 (N_2475,N_1542,N_1953);
and U2476 (N_2476,N_1717,N_1947);
nor U2477 (N_2477,N_1835,N_1938);
and U2478 (N_2478,N_1556,N_1739);
or U2479 (N_2479,N_1744,N_1656);
nor U2480 (N_2480,N_1743,N_1740);
nor U2481 (N_2481,N_1905,N_1573);
or U2482 (N_2482,N_1938,N_1673);
or U2483 (N_2483,N_1680,N_1713);
nand U2484 (N_2484,N_1676,N_1558);
nand U2485 (N_2485,N_1550,N_1707);
or U2486 (N_2486,N_1544,N_1674);
and U2487 (N_2487,N_1591,N_1807);
and U2488 (N_2488,N_1723,N_1949);
nor U2489 (N_2489,N_1729,N_1733);
nor U2490 (N_2490,N_1861,N_1799);
and U2491 (N_2491,N_1574,N_1573);
xor U2492 (N_2492,N_1550,N_1603);
or U2493 (N_2493,N_1848,N_1751);
or U2494 (N_2494,N_1653,N_1980);
nand U2495 (N_2495,N_1831,N_1800);
nand U2496 (N_2496,N_1945,N_1641);
nor U2497 (N_2497,N_1742,N_1650);
and U2498 (N_2498,N_1721,N_1711);
or U2499 (N_2499,N_1600,N_1672);
or U2500 (N_2500,N_2383,N_2471);
nor U2501 (N_2501,N_2392,N_2277);
and U2502 (N_2502,N_2219,N_2474);
and U2503 (N_2503,N_2336,N_2415);
or U2504 (N_2504,N_2213,N_2438);
and U2505 (N_2505,N_2351,N_2171);
nand U2506 (N_2506,N_2429,N_2332);
nand U2507 (N_2507,N_2183,N_2265);
xor U2508 (N_2508,N_2456,N_2267);
or U2509 (N_2509,N_2387,N_2096);
nor U2510 (N_2510,N_2012,N_2036);
or U2511 (N_2511,N_2488,N_2376);
and U2512 (N_2512,N_2228,N_2168);
or U2513 (N_2513,N_2099,N_2320);
nor U2514 (N_2514,N_2367,N_2083);
and U2515 (N_2515,N_2377,N_2358);
and U2516 (N_2516,N_2234,N_2273);
and U2517 (N_2517,N_2087,N_2023);
and U2518 (N_2518,N_2208,N_2485);
nor U2519 (N_2519,N_2451,N_2431);
and U2520 (N_2520,N_2394,N_2495);
or U2521 (N_2521,N_2430,N_2340);
or U2522 (N_2522,N_2255,N_2078);
or U2523 (N_2523,N_2315,N_2209);
nor U2524 (N_2524,N_2420,N_2442);
and U2525 (N_2525,N_2380,N_2068);
nor U2526 (N_2526,N_2196,N_2236);
or U2527 (N_2527,N_2008,N_2066);
and U2528 (N_2528,N_2027,N_2342);
or U2529 (N_2529,N_2436,N_2417);
nor U2530 (N_2530,N_2090,N_2347);
nor U2531 (N_2531,N_2335,N_2092);
nand U2532 (N_2532,N_2085,N_2256);
nor U2533 (N_2533,N_2455,N_2278);
nor U2534 (N_2534,N_2356,N_2481);
and U2535 (N_2535,N_2125,N_2165);
nand U2536 (N_2536,N_2005,N_2077);
nor U2537 (N_2537,N_2251,N_2084);
nor U2538 (N_2538,N_2200,N_2112);
and U2539 (N_2539,N_2288,N_2206);
nand U2540 (N_2540,N_2454,N_2312);
nand U2541 (N_2541,N_2184,N_2137);
nand U2542 (N_2542,N_2047,N_2229);
or U2543 (N_2543,N_2182,N_2469);
nor U2544 (N_2544,N_2154,N_2432);
nand U2545 (N_2545,N_2447,N_2398);
or U2546 (N_2546,N_2143,N_2248);
nand U2547 (N_2547,N_2289,N_2249);
nor U2548 (N_2548,N_2250,N_2384);
or U2549 (N_2549,N_2227,N_2355);
nor U2550 (N_2550,N_2155,N_2339);
nand U2551 (N_2551,N_2461,N_2460);
nor U2552 (N_2552,N_2016,N_2327);
or U2553 (N_2553,N_2070,N_2475);
and U2554 (N_2554,N_2181,N_2310);
and U2555 (N_2555,N_2483,N_2296);
and U2556 (N_2556,N_2379,N_2161);
or U2557 (N_2557,N_2030,N_2011);
and U2558 (N_2558,N_2220,N_2202);
and U2559 (N_2559,N_2266,N_2478);
and U2560 (N_2560,N_2276,N_2364);
or U2561 (N_2561,N_2080,N_2319);
nor U2562 (N_2562,N_2362,N_2174);
and U2563 (N_2563,N_2424,N_2318);
and U2564 (N_2564,N_2348,N_2440);
and U2565 (N_2565,N_2166,N_2263);
or U2566 (N_2566,N_2437,N_2097);
nor U2567 (N_2567,N_2100,N_2217);
and U2568 (N_2568,N_2244,N_2138);
nor U2569 (N_2569,N_2374,N_2257);
and U2570 (N_2570,N_2314,N_2245);
and U2571 (N_2571,N_2486,N_2258);
nand U2572 (N_2572,N_2477,N_2410);
nand U2573 (N_2573,N_2283,N_2185);
nor U2574 (N_2574,N_2224,N_2121);
nand U2575 (N_2575,N_2282,N_2307);
and U2576 (N_2576,N_2223,N_2158);
and U2577 (N_2577,N_2313,N_2345);
and U2578 (N_2578,N_2007,N_2350);
or U2579 (N_2579,N_2239,N_2285);
nor U2580 (N_2580,N_2179,N_2371);
nand U2581 (N_2581,N_2104,N_2020);
or U2582 (N_2582,N_2082,N_2055);
nor U2583 (N_2583,N_2024,N_2006);
nand U2584 (N_2584,N_2026,N_2139);
and U2585 (N_2585,N_2443,N_2328);
nand U2586 (N_2586,N_2439,N_2069);
nand U2587 (N_2587,N_2091,N_2446);
nand U2588 (N_2588,N_2109,N_2052);
nor U2589 (N_2589,N_2299,N_2218);
nand U2590 (N_2590,N_2311,N_2041);
or U2591 (N_2591,N_2389,N_2043);
nor U2592 (N_2592,N_2441,N_2473);
and U2593 (N_2593,N_2357,N_2260);
or U2594 (N_2594,N_2094,N_2452);
nand U2595 (N_2595,N_2064,N_2366);
or U2596 (N_2596,N_2309,N_2130);
and U2597 (N_2597,N_2022,N_2042);
or U2598 (N_2598,N_2468,N_2416);
and U2599 (N_2599,N_2049,N_2129);
nand U2600 (N_2600,N_2406,N_2400);
nor U2601 (N_2601,N_2145,N_2017);
and U2602 (N_2602,N_2386,N_2038);
nand U2603 (N_2603,N_2075,N_2003);
nand U2604 (N_2604,N_2081,N_2458);
nor U2605 (N_2605,N_2186,N_2222);
nand U2606 (N_2606,N_2060,N_2190);
or U2607 (N_2607,N_2144,N_2086);
or U2608 (N_2608,N_2466,N_2302);
and U2609 (N_2609,N_2113,N_2467);
or U2610 (N_2610,N_2074,N_2173);
or U2611 (N_2611,N_2402,N_2063);
nor U2612 (N_2612,N_2395,N_2287);
or U2613 (N_2613,N_2304,N_2088);
and U2614 (N_2614,N_2300,N_2433);
nand U2615 (N_2615,N_2463,N_2344);
nand U2616 (N_2616,N_2157,N_2221);
nor U2617 (N_2617,N_2180,N_2116);
and U2618 (N_2618,N_2025,N_2034);
nor U2619 (N_2619,N_2105,N_2491);
nor U2620 (N_2620,N_2292,N_2413);
nand U2621 (N_2621,N_2427,N_2284);
or U2622 (N_2622,N_2151,N_2295);
and U2623 (N_2623,N_2059,N_2054);
and U2624 (N_2624,N_2131,N_2193);
or U2625 (N_2625,N_2408,N_2393);
and U2626 (N_2626,N_2153,N_2065);
or U2627 (N_2627,N_2388,N_2163);
nand U2628 (N_2628,N_2149,N_2423);
nor U2629 (N_2629,N_2498,N_2396);
or U2630 (N_2630,N_2124,N_2061);
and U2631 (N_2631,N_2462,N_2487);
nand U2632 (N_2632,N_2286,N_2192);
and U2633 (N_2633,N_2457,N_2210);
and U2634 (N_2634,N_2201,N_2253);
xor U2635 (N_2635,N_2194,N_2268);
nor U2636 (N_2636,N_2259,N_2051);
nand U2637 (N_2637,N_2419,N_2382);
xor U2638 (N_2638,N_2363,N_2341);
or U2639 (N_2639,N_2373,N_2290);
nor U2640 (N_2640,N_2493,N_2148);
or U2641 (N_2641,N_2127,N_2490);
and U2642 (N_2642,N_2411,N_2226);
nand U2643 (N_2643,N_2019,N_2412);
and U2644 (N_2644,N_2067,N_2294);
and U2645 (N_2645,N_2334,N_2031);
nand U2646 (N_2646,N_2470,N_2275);
or U2647 (N_2647,N_2141,N_2207);
or U2648 (N_2648,N_2204,N_2337);
and U2649 (N_2649,N_2496,N_2000);
nor U2650 (N_2650,N_2136,N_2164);
xnor U2651 (N_2651,N_2499,N_2274);
or U2652 (N_2652,N_2102,N_2106);
nor U2653 (N_2653,N_2238,N_2178);
nand U2654 (N_2654,N_2370,N_2492);
xnor U2655 (N_2655,N_2323,N_2089);
nand U2656 (N_2656,N_2128,N_2333);
nand U2657 (N_2657,N_2279,N_2150);
nor U2658 (N_2658,N_2444,N_2039);
and U2659 (N_2659,N_2421,N_2449);
or U2660 (N_2660,N_2252,N_2448);
and U2661 (N_2661,N_2142,N_2385);
and U2662 (N_2662,N_2009,N_2001);
or U2663 (N_2663,N_2346,N_2272);
and U2664 (N_2664,N_2293,N_2324);
or U2665 (N_2665,N_2303,N_2365);
nand U2666 (N_2666,N_2280,N_2464);
and U2667 (N_2667,N_2426,N_2317);
and U2668 (N_2668,N_2191,N_2115);
or U2669 (N_2669,N_2018,N_2240);
and U2670 (N_2670,N_2409,N_2322);
or U2671 (N_2671,N_2422,N_2349);
nand U2672 (N_2672,N_2435,N_2140);
nand U2673 (N_2673,N_2445,N_2414);
and U2674 (N_2674,N_2015,N_2407);
or U2675 (N_2675,N_2434,N_2212);
nand U2676 (N_2676,N_2241,N_2172);
nand U2677 (N_2677,N_2021,N_2391);
or U2678 (N_2678,N_2243,N_2134);
or U2679 (N_2679,N_2308,N_2372);
nand U2680 (N_2680,N_2399,N_2119);
nand U2681 (N_2681,N_2199,N_2135);
nor U2682 (N_2682,N_2198,N_2162);
nand U2683 (N_2683,N_2476,N_2029);
and U2684 (N_2684,N_2237,N_2111);
nor U2685 (N_2685,N_2484,N_2459);
nand U2686 (N_2686,N_2479,N_2298);
or U2687 (N_2687,N_2326,N_2152);
nor U2688 (N_2688,N_2305,N_2375);
nor U2689 (N_2689,N_2401,N_2261);
and U2690 (N_2690,N_2281,N_2133);
nand U2691 (N_2691,N_2247,N_2205);
nor U2692 (N_2692,N_2072,N_2403);
and U2693 (N_2693,N_2330,N_2120);
nand U2694 (N_2694,N_2167,N_2215);
nor U2695 (N_2695,N_2101,N_2354);
and U2696 (N_2696,N_2132,N_2233);
nand U2697 (N_2697,N_2044,N_2004);
and U2698 (N_2698,N_2405,N_2397);
nor U2699 (N_2699,N_2188,N_2361);
xnor U2700 (N_2700,N_2231,N_2013);
and U2701 (N_2701,N_2203,N_2033);
or U2702 (N_2702,N_2425,N_2331);
and U2703 (N_2703,N_2076,N_2062);
and U2704 (N_2704,N_2028,N_2262);
or U2705 (N_2705,N_2494,N_2108);
and U2706 (N_2706,N_2037,N_2325);
and U2707 (N_2707,N_2301,N_2291);
and U2708 (N_2708,N_2359,N_2368);
nor U2709 (N_2709,N_2254,N_2056);
and U2710 (N_2710,N_2214,N_2225);
and U2711 (N_2711,N_2271,N_2117);
and U2712 (N_2712,N_2306,N_2118);
and U2713 (N_2713,N_2032,N_2369);
nand U2714 (N_2714,N_2329,N_2235);
and U2715 (N_2715,N_2122,N_2014);
or U2716 (N_2716,N_2169,N_2418);
or U2717 (N_2717,N_2175,N_2058);
and U2718 (N_2718,N_2048,N_2126);
nand U2719 (N_2719,N_2453,N_2230);
and U2720 (N_2720,N_2079,N_2123);
or U2721 (N_2721,N_2045,N_2338);
and U2722 (N_2722,N_2146,N_2465);
nor U2723 (N_2723,N_2321,N_2093);
nor U2724 (N_2724,N_2316,N_2195);
nor U2725 (N_2725,N_2159,N_2489);
nand U2726 (N_2726,N_2264,N_2211);
nand U2727 (N_2727,N_2189,N_2232);
nand U2728 (N_2728,N_2095,N_2057);
nand U2729 (N_2729,N_2352,N_2472);
or U2730 (N_2730,N_2269,N_2098);
or U2731 (N_2731,N_2187,N_2160);
nand U2732 (N_2732,N_2378,N_2216);
or U2733 (N_2733,N_2242,N_2404);
nor U2734 (N_2734,N_2297,N_2156);
nor U2735 (N_2735,N_2197,N_2107);
and U2736 (N_2736,N_2390,N_2050);
nor U2737 (N_2737,N_2073,N_2170);
nand U2738 (N_2738,N_2040,N_2246);
nand U2739 (N_2739,N_2353,N_2270);
nand U2740 (N_2740,N_2114,N_2176);
and U2741 (N_2741,N_2497,N_2428);
and U2742 (N_2742,N_2071,N_2002);
or U2743 (N_2743,N_2482,N_2053);
or U2744 (N_2744,N_2110,N_2177);
or U2745 (N_2745,N_2103,N_2343);
or U2746 (N_2746,N_2360,N_2480);
nor U2747 (N_2747,N_2381,N_2147);
nand U2748 (N_2748,N_2450,N_2046);
and U2749 (N_2749,N_2035,N_2010);
or U2750 (N_2750,N_2001,N_2225);
or U2751 (N_2751,N_2411,N_2238);
nor U2752 (N_2752,N_2322,N_2117);
or U2753 (N_2753,N_2061,N_2146);
or U2754 (N_2754,N_2444,N_2275);
nor U2755 (N_2755,N_2000,N_2478);
nor U2756 (N_2756,N_2385,N_2177);
nor U2757 (N_2757,N_2009,N_2472);
or U2758 (N_2758,N_2341,N_2159);
or U2759 (N_2759,N_2126,N_2391);
and U2760 (N_2760,N_2235,N_2006);
nand U2761 (N_2761,N_2452,N_2209);
nor U2762 (N_2762,N_2292,N_2034);
nand U2763 (N_2763,N_2350,N_2477);
or U2764 (N_2764,N_2436,N_2187);
and U2765 (N_2765,N_2433,N_2292);
or U2766 (N_2766,N_2463,N_2270);
nor U2767 (N_2767,N_2202,N_2412);
or U2768 (N_2768,N_2499,N_2039);
or U2769 (N_2769,N_2369,N_2312);
nand U2770 (N_2770,N_2095,N_2058);
xor U2771 (N_2771,N_2050,N_2269);
or U2772 (N_2772,N_2491,N_2443);
xnor U2773 (N_2773,N_2391,N_2015);
nor U2774 (N_2774,N_2208,N_2447);
nor U2775 (N_2775,N_2041,N_2383);
nor U2776 (N_2776,N_2304,N_2287);
or U2777 (N_2777,N_2103,N_2357);
and U2778 (N_2778,N_2169,N_2450);
nand U2779 (N_2779,N_2469,N_2447);
and U2780 (N_2780,N_2408,N_2107);
nand U2781 (N_2781,N_2336,N_2467);
and U2782 (N_2782,N_2440,N_2133);
or U2783 (N_2783,N_2237,N_2372);
nand U2784 (N_2784,N_2317,N_2124);
or U2785 (N_2785,N_2471,N_2406);
and U2786 (N_2786,N_2271,N_2432);
and U2787 (N_2787,N_2122,N_2347);
nor U2788 (N_2788,N_2360,N_2211);
or U2789 (N_2789,N_2387,N_2271);
or U2790 (N_2790,N_2027,N_2054);
and U2791 (N_2791,N_2433,N_2430);
nor U2792 (N_2792,N_2165,N_2135);
nor U2793 (N_2793,N_2451,N_2487);
nand U2794 (N_2794,N_2245,N_2323);
nor U2795 (N_2795,N_2096,N_2318);
or U2796 (N_2796,N_2123,N_2057);
or U2797 (N_2797,N_2204,N_2127);
and U2798 (N_2798,N_2135,N_2325);
nor U2799 (N_2799,N_2090,N_2073);
nand U2800 (N_2800,N_2334,N_2485);
nand U2801 (N_2801,N_2275,N_2181);
and U2802 (N_2802,N_2451,N_2033);
and U2803 (N_2803,N_2273,N_2281);
and U2804 (N_2804,N_2279,N_2427);
xor U2805 (N_2805,N_2278,N_2154);
and U2806 (N_2806,N_2253,N_2150);
or U2807 (N_2807,N_2491,N_2104);
nand U2808 (N_2808,N_2145,N_2454);
nand U2809 (N_2809,N_2401,N_2259);
nor U2810 (N_2810,N_2094,N_2223);
nor U2811 (N_2811,N_2121,N_2088);
nand U2812 (N_2812,N_2140,N_2003);
and U2813 (N_2813,N_2414,N_2195);
xor U2814 (N_2814,N_2432,N_2046);
or U2815 (N_2815,N_2376,N_2209);
and U2816 (N_2816,N_2342,N_2022);
nand U2817 (N_2817,N_2384,N_2202);
nand U2818 (N_2818,N_2403,N_2029);
nor U2819 (N_2819,N_2014,N_2496);
and U2820 (N_2820,N_2080,N_2121);
nor U2821 (N_2821,N_2370,N_2121);
and U2822 (N_2822,N_2417,N_2491);
nand U2823 (N_2823,N_2148,N_2351);
and U2824 (N_2824,N_2134,N_2492);
nor U2825 (N_2825,N_2314,N_2247);
nor U2826 (N_2826,N_2139,N_2145);
nor U2827 (N_2827,N_2427,N_2181);
nor U2828 (N_2828,N_2055,N_2369);
or U2829 (N_2829,N_2223,N_2392);
and U2830 (N_2830,N_2311,N_2154);
and U2831 (N_2831,N_2279,N_2256);
nor U2832 (N_2832,N_2381,N_2457);
nor U2833 (N_2833,N_2051,N_2353);
and U2834 (N_2834,N_2163,N_2230);
nor U2835 (N_2835,N_2386,N_2308);
nor U2836 (N_2836,N_2397,N_2474);
or U2837 (N_2837,N_2193,N_2202);
nor U2838 (N_2838,N_2047,N_2168);
nand U2839 (N_2839,N_2399,N_2110);
nand U2840 (N_2840,N_2248,N_2370);
nand U2841 (N_2841,N_2085,N_2451);
or U2842 (N_2842,N_2326,N_2172);
and U2843 (N_2843,N_2339,N_2121);
nand U2844 (N_2844,N_2038,N_2399);
nor U2845 (N_2845,N_2158,N_2468);
nand U2846 (N_2846,N_2348,N_2138);
nand U2847 (N_2847,N_2309,N_2280);
xor U2848 (N_2848,N_2439,N_2007);
and U2849 (N_2849,N_2298,N_2324);
and U2850 (N_2850,N_2367,N_2455);
or U2851 (N_2851,N_2273,N_2474);
or U2852 (N_2852,N_2259,N_2285);
or U2853 (N_2853,N_2137,N_2012);
nor U2854 (N_2854,N_2351,N_2360);
and U2855 (N_2855,N_2457,N_2265);
nor U2856 (N_2856,N_2085,N_2308);
nand U2857 (N_2857,N_2038,N_2439);
or U2858 (N_2858,N_2261,N_2137);
nor U2859 (N_2859,N_2439,N_2193);
or U2860 (N_2860,N_2254,N_2478);
nand U2861 (N_2861,N_2282,N_2433);
or U2862 (N_2862,N_2245,N_2412);
or U2863 (N_2863,N_2069,N_2092);
nor U2864 (N_2864,N_2402,N_2219);
nand U2865 (N_2865,N_2140,N_2252);
nand U2866 (N_2866,N_2379,N_2003);
or U2867 (N_2867,N_2066,N_2422);
and U2868 (N_2868,N_2308,N_2383);
nor U2869 (N_2869,N_2294,N_2391);
nand U2870 (N_2870,N_2352,N_2217);
nand U2871 (N_2871,N_2192,N_2088);
and U2872 (N_2872,N_2257,N_2397);
nand U2873 (N_2873,N_2394,N_2048);
or U2874 (N_2874,N_2200,N_2366);
nor U2875 (N_2875,N_2499,N_2395);
nor U2876 (N_2876,N_2226,N_2220);
nor U2877 (N_2877,N_2212,N_2106);
nand U2878 (N_2878,N_2386,N_2297);
nand U2879 (N_2879,N_2369,N_2114);
and U2880 (N_2880,N_2055,N_2458);
nand U2881 (N_2881,N_2350,N_2144);
and U2882 (N_2882,N_2273,N_2165);
nand U2883 (N_2883,N_2274,N_2336);
nand U2884 (N_2884,N_2069,N_2462);
nor U2885 (N_2885,N_2118,N_2154);
and U2886 (N_2886,N_2258,N_2335);
nor U2887 (N_2887,N_2041,N_2487);
nor U2888 (N_2888,N_2312,N_2190);
or U2889 (N_2889,N_2269,N_2185);
and U2890 (N_2890,N_2326,N_2124);
nor U2891 (N_2891,N_2164,N_2435);
and U2892 (N_2892,N_2075,N_2272);
and U2893 (N_2893,N_2302,N_2090);
or U2894 (N_2894,N_2337,N_2113);
nand U2895 (N_2895,N_2110,N_2355);
or U2896 (N_2896,N_2144,N_2126);
and U2897 (N_2897,N_2269,N_2292);
or U2898 (N_2898,N_2073,N_2064);
nand U2899 (N_2899,N_2449,N_2240);
nand U2900 (N_2900,N_2425,N_2231);
nand U2901 (N_2901,N_2487,N_2084);
xnor U2902 (N_2902,N_2128,N_2462);
nor U2903 (N_2903,N_2459,N_2454);
nor U2904 (N_2904,N_2031,N_2181);
and U2905 (N_2905,N_2147,N_2499);
nand U2906 (N_2906,N_2030,N_2410);
or U2907 (N_2907,N_2129,N_2478);
and U2908 (N_2908,N_2461,N_2330);
nor U2909 (N_2909,N_2018,N_2085);
or U2910 (N_2910,N_2203,N_2350);
nor U2911 (N_2911,N_2287,N_2025);
or U2912 (N_2912,N_2066,N_2493);
and U2913 (N_2913,N_2148,N_2441);
nand U2914 (N_2914,N_2475,N_2199);
nor U2915 (N_2915,N_2437,N_2078);
and U2916 (N_2916,N_2254,N_2263);
and U2917 (N_2917,N_2309,N_2235);
nor U2918 (N_2918,N_2384,N_2240);
or U2919 (N_2919,N_2103,N_2433);
nand U2920 (N_2920,N_2265,N_2216);
and U2921 (N_2921,N_2064,N_2487);
nand U2922 (N_2922,N_2389,N_2387);
nor U2923 (N_2923,N_2122,N_2148);
nor U2924 (N_2924,N_2052,N_2409);
or U2925 (N_2925,N_2255,N_2286);
and U2926 (N_2926,N_2224,N_2141);
and U2927 (N_2927,N_2137,N_2161);
xor U2928 (N_2928,N_2068,N_2027);
and U2929 (N_2929,N_2415,N_2435);
nor U2930 (N_2930,N_2421,N_2222);
or U2931 (N_2931,N_2380,N_2073);
or U2932 (N_2932,N_2117,N_2205);
nor U2933 (N_2933,N_2044,N_2486);
nand U2934 (N_2934,N_2173,N_2336);
nor U2935 (N_2935,N_2233,N_2031);
or U2936 (N_2936,N_2254,N_2087);
nand U2937 (N_2937,N_2436,N_2202);
nor U2938 (N_2938,N_2384,N_2326);
or U2939 (N_2939,N_2076,N_2124);
nand U2940 (N_2940,N_2006,N_2368);
nand U2941 (N_2941,N_2125,N_2064);
and U2942 (N_2942,N_2196,N_2132);
and U2943 (N_2943,N_2331,N_2118);
and U2944 (N_2944,N_2019,N_2386);
nand U2945 (N_2945,N_2183,N_2227);
and U2946 (N_2946,N_2261,N_2494);
or U2947 (N_2947,N_2024,N_2367);
xnor U2948 (N_2948,N_2110,N_2420);
and U2949 (N_2949,N_2165,N_2128);
and U2950 (N_2950,N_2310,N_2036);
or U2951 (N_2951,N_2297,N_2081);
and U2952 (N_2952,N_2116,N_2351);
or U2953 (N_2953,N_2074,N_2082);
nand U2954 (N_2954,N_2444,N_2487);
nand U2955 (N_2955,N_2292,N_2264);
or U2956 (N_2956,N_2081,N_2174);
nor U2957 (N_2957,N_2113,N_2328);
xor U2958 (N_2958,N_2081,N_2137);
or U2959 (N_2959,N_2272,N_2070);
nor U2960 (N_2960,N_2492,N_2166);
nor U2961 (N_2961,N_2350,N_2236);
or U2962 (N_2962,N_2164,N_2474);
and U2963 (N_2963,N_2473,N_2337);
nand U2964 (N_2964,N_2066,N_2394);
nor U2965 (N_2965,N_2187,N_2346);
and U2966 (N_2966,N_2084,N_2129);
nand U2967 (N_2967,N_2168,N_2121);
nor U2968 (N_2968,N_2197,N_2461);
or U2969 (N_2969,N_2011,N_2084);
xor U2970 (N_2970,N_2242,N_2200);
and U2971 (N_2971,N_2061,N_2190);
xnor U2972 (N_2972,N_2333,N_2247);
and U2973 (N_2973,N_2069,N_2055);
nor U2974 (N_2974,N_2341,N_2044);
nand U2975 (N_2975,N_2361,N_2109);
nor U2976 (N_2976,N_2163,N_2384);
and U2977 (N_2977,N_2233,N_2455);
nor U2978 (N_2978,N_2484,N_2247);
nand U2979 (N_2979,N_2467,N_2449);
or U2980 (N_2980,N_2321,N_2346);
nor U2981 (N_2981,N_2443,N_2032);
and U2982 (N_2982,N_2003,N_2119);
nor U2983 (N_2983,N_2391,N_2488);
nor U2984 (N_2984,N_2028,N_2484);
nand U2985 (N_2985,N_2317,N_2422);
and U2986 (N_2986,N_2352,N_2120);
or U2987 (N_2987,N_2491,N_2051);
and U2988 (N_2988,N_2254,N_2173);
nor U2989 (N_2989,N_2066,N_2456);
and U2990 (N_2990,N_2317,N_2284);
or U2991 (N_2991,N_2242,N_2187);
nand U2992 (N_2992,N_2381,N_2342);
and U2993 (N_2993,N_2095,N_2190);
and U2994 (N_2994,N_2239,N_2495);
or U2995 (N_2995,N_2109,N_2334);
nand U2996 (N_2996,N_2001,N_2002);
or U2997 (N_2997,N_2212,N_2428);
nor U2998 (N_2998,N_2296,N_2442);
and U2999 (N_2999,N_2470,N_2389);
or U3000 (N_3000,N_2948,N_2946);
and U3001 (N_3001,N_2819,N_2715);
nor U3002 (N_3002,N_2924,N_2616);
nor U3003 (N_3003,N_2860,N_2568);
and U3004 (N_3004,N_2675,N_2713);
or U3005 (N_3005,N_2595,N_2662);
nor U3006 (N_3006,N_2575,N_2642);
and U3007 (N_3007,N_2983,N_2809);
and U3008 (N_3008,N_2889,N_2626);
nand U3009 (N_3009,N_2517,N_2979);
nand U3010 (N_3010,N_2947,N_2835);
nor U3011 (N_3011,N_2991,N_2898);
or U3012 (N_3012,N_2960,N_2927);
nor U3013 (N_3013,N_2623,N_2605);
or U3014 (N_3014,N_2895,N_2921);
or U3015 (N_3015,N_2756,N_2646);
nand U3016 (N_3016,N_2980,N_2825);
or U3017 (N_3017,N_2711,N_2741);
nand U3018 (N_3018,N_2964,N_2910);
and U3019 (N_3019,N_2743,N_2788);
nor U3020 (N_3020,N_2515,N_2665);
or U3021 (N_3021,N_2716,N_2841);
nand U3022 (N_3022,N_2651,N_2591);
or U3023 (N_3023,N_2552,N_2859);
nor U3024 (N_3024,N_2698,N_2962);
nor U3025 (N_3025,N_2978,N_2805);
nor U3026 (N_3026,N_2998,N_2974);
nor U3027 (N_3027,N_2613,N_2648);
nand U3028 (N_3028,N_2563,N_2858);
and U3029 (N_3029,N_2864,N_2754);
or U3030 (N_3030,N_2718,N_2580);
nor U3031 (N_3031,N_2888,N_2846);
and U3032 (N_3032,N_2932,N_2855);
nor U3033 (N_3033,N_2637,N_2644);
or U3034 (N_3034,N_2543,N_2993);
nor U3035 (N_3035,N_2759,N_2724);
xnor U3036 (N_3036,N_2597,N_2832);
or U3037 (N_3037,N_2972,N_2638);
nand U3038 (N_3038,N_2663,N_2919);
or U3039 (N_3039,N_2562,N_2996);
and U3040 (N_3040,N_2769,N_2565);
nand U3041 (N_3041,N_2952,N_2514);
and U3042 (N_3042,N_2857,N_2699);
nor U3043 (N_3043,N_2770,N_2607);
and U3044 (N_3044,N_2670,N_2882);
or U3045 (N_3045,N_2585,N_2886);
nand U3046 (N_3046,N_2781,N_2522);
nand U3047 (N_3047,N_2842,N_2686);
nand U3048 (N_3048,N_2837,N_2655);
nand U3049 (N_3049,N_2752,N_2577);
and U3050 (N_3050,N_2620,N_2868);
and U3051 (N_3051,N_2659,N_2934);
and U3052 (N_3052,N_2541,N_2918);
nor U3053 (N_3053,N_2973,N_2786);
nand U3054 (N_3054,N_2959,N_2624);
nor U3055 (N_3055,N_2679,N_2779);
nand U3056 (N_3056,N_2518,N_2869);
nand U3057 (N_3057,N_2981,N_2907);
and U3058 (N_3058,N_2750,N_2745);
and U3059 (N_3059,N_2672,N_2818);
nand U3060 (N_3060,N_2903,N_2574);
or U3061 (N_3061,N_2806,N_2787);
nor U3062 (N_3062,N_2717,N_2922);
nand U3063 (N_3063,N_2576,N_2969);
or U3064 (N_3064,N_2813,N_2951);
or U3065 (N_3065,N_2722,N_2684);
or U3066 (N_3066,N_2506,N_2906);
and U3067 (N_3067,N_2554,N_2821);
nor U3068 (N_3068,N_2594,N_2749);
nand U3069 (N_3069,N_2720,N_2949);
nor U3070 (N_3070,N_2505,N_2887);
nor U3071 (N_3071,N_2564,N_2984);
nand U3072 (N_3072,N_2997,N_2693);
nand U3073 (N_3073,N_2854,N_2782);
nand U3074 (N_3074,N_2671,N_2872);
nand U3075 (N_3075,N_2634,N_2789);
nor U3076 (N_3076,N_2765,N_2852);
nand U3077 (N_3077,N_2617,N_2762);
nor U3078 (N_3078,N_2673,N_2767);
and U3079 (N_3079,N_2798,N_2650);
and U3080 (N_3080,N_2739,N_2555);
and U3081 (N_3081,N_2967,N_2584);
and U3082 (N_3082,N_2917,N_2538);
or U3083 (N_3083,N_2810,N_2558);
nor U3084 (N_3084,N_2950,N_2795);
or U3085 (N_3085,N_2677,N_2500);
nand U3086 (N_3086,N_2849,N_2791);
nand U3087 (N_3087,N_2830,N_2838);
nor U3088 (N_3088,N_2590,N_2884);
nor U3089 (N_3089,N_2583,N_2897);
and U3090 (N_3090,N_2714,N_2687);
nand U3091 (N_3091,N_2916,N_2862);
and U3092 (N_3092,N_2531,N_2870);
nand U3093 (N_3093,N_2933,N_2744);
or U3094 (N_3094,N_2566,N_2645);
xor U3095 (N_3095,N_2804,N_2545);
or U3096 (N_3096,N_2828,N_2661);
or U3097 (N_3097,N_2847,N_2625);
nand U3098 (N_3098,N_2530,N_2502);
nand U3099 (N_3099,N_2635,N_2908);
nor U3100 (N_3100,N_2970,N_2920);
nor U3101 (N_3101,N_2523,N_2829);
xor U3102 (N_3102,N_2778,N_2676);
nor U3103 (N_3103,N_2682,N_2550);
nand U3104 (N_3104,N_2764,N_2723);
and U3105 (N_3105,N_2866,N_2956);
nand U3106 (N_3106,N_2525,N_2513);
nor U3107 (N_3107,N_2851,N_2811);
nand U3108 (N_3108,N_2939,N_2794);
nor U3109 (N_3109,N_2706,N_2877);
or U3110 (N_3110,N_2943,N_2905);
and U3111 (N_3111,N_2654,N_2975);
nand U3112 (N_3112,N_2742,N_2604);
or U3113 (N_3113,N_2596,N_2885);
or U3114 (N_3114,N_2509,N_2503);
nor U3115 (N_3115,N_2938,N_2823);
or U3116 (N_3116,N_2601,N_2957);
or U3117 (N_3117,N_2579,N_2527);
or U3118 (N_3118,N_2894,N_2628);
nand U3119 (N_3119,N_2982,N_2578);
and U3120 (N_3120,N_2871,N_2935);
nand U3121 (N_3121,N_2629,N_2844);
or U3122 (N_3122,N_2913,N_2704);
or U3123 (N_3123,N_2664,N_2833);
and U3124 (N_3124,N_2986,N_2912);
and U3125 (N_3125,N_2937,N_2930);
or U3126 (N_3126,N_2532,N_2740);
nand U3127 (N_3127,N_2533,N_2614);
nor U3128 (N_3128,N_2736,N_2529);
and U3129 (N_3129,N_2548,N_2603);
or U3130 (N_3130,N_2630,N_2599);
nor U3131 (N_3131,N_2755,N_2843);
and U3132 (N_3132,N_2690,N_2587);
and U3133 (N_3133,N_2547,N_2944);
nand U3134 (N_3134,N_2516,N_2734);
nor U3135 (N_3135,N_2612,N_2721);
nand U3136 (N_3136,N_2586,N_2669);
nand U3137 (N_3137,N_2685,N_2507);
xor U3138 (N_3138,N_2928,N_2971);
or U3139 (N_3139,N_2689,N_2892);
nor U3140 (N_3140,N_2621,N_2936);
and U3141 (N_3141,N_2761,N_2727);
and U3142 (N_3142,N_2876,N_2987);
xnor U3143 (N_3143,N_2940,N_2800);
nor U3144 (N_3144,N_2560,N_2836);
and U3145 (N_3145,N_2510,N_2840);
nand U3146 (N_3146,N_2707,N_2737);
nand U3147 (N_3147,N_2520,N_2783);
nand U3148 (N_3148,N_2549,N_2817);
or U3149 (N_3149,N_2536,N_2528);
and U3150 (N_3150,N_2521,N_2901);
and U3151 (N_3151,N_2942,N_2816);
nand U3152 (N_3152,N_2653,N_2559);
and U3153 (N_3153,N_2738,N_2799);
nand U3154 (N_3154,N_2881,N_2668);
nor U3155 (N_3155,N_2780,N_2691);
nand U3156 (N_3156,N_2988,N_2963);
xor U3157 (N_3157,N_2524,N_2702);
nand U3158 (N_3158,N_2611,N_2569);
nand U3159 (N_3159,N_2773,N_2619);
xnor U3160 (N_3160,N_2772,N_2923);
and U3161 (N_3161,N_2802,N_2891);
and U3162 (N_3162,N_2719,N_2931);
and U3163 (N_3163,N_2966,N_2863);
nand U3164 (N_3164,N_2695,N_2853);
or U3165 (N_3165,N_2504,N_2880);
or U3166 (N_3166,N_2641,N_2732);
and U3167 (N_3167,N_2639,N_2815);
or U3168 (N_3168,N_2501,N_2537);
nor U3169 (N_3169,N_2582,N_2519);
nand U3170 (N_3170,N_2588,N_2992);
or U3171 (N_3171,N_2774,N_2708);
and U3172 (N_3172,N_2725,N_2953);
or U3173 (N_3173,N_2995,N_2994);
nor U3174 (N_3174,N_2753,N_2955);
nor U3175 (N_3175,N_2649,N_2883);
nor U3176 (N_3176,N_2726,N_2561);
nor U3177 (N_3177,N_2848,N_2570);
nor U3178 (N_3178,N_2567,N_2729);
or U3179 (N_3179,N_2674,N_2989);
nand U3180 (N_3180,N_2961,N_2879);
and U3181 (N_3181,N_2571,N_2608);
nand U3182 (N_3182,N_2730,N_2683);
nor U3183 (N_3183,N_2822,N_2534);
or U3184 (N_3184,N_2904,N_2824);
nor U3185 (N_3185,N_2915,N_2508);
nand U3186 (N_3186,N_2766,N_2856);
or U3187 (N_3187,N_2540,N_2990);
nor U3188 (N_3188,N_2826,N_2965);
nand U3189 (N_3189,N_2705,N_2512);
and U3190 (N_3190,N_2968,N_2610);
or U3191 (N_3191,N_2697,N_2593);
nand U3192 (N_3192,N_2875,N_2784);
nor U3193 (N_3193,N_2977,N_2700);
or U3194 (N_3194,N_2573,N_2776);
nor U3195 (N_3195,N_2710,N_2909);
nand U3196 (N_3196,N_2874,N_2834);
xnor U3197 (N_3197,N_2688,N_2758);
or U3198 (N_3198,N_2839,N_2985);
nand U3199 (N_3199,N_2793,N_2666);
and U3200 (N_3200,N_2771,N_2797);
nor U3201 (N_3201,N_2615,N_2600);
nand U3202 (N_3202,N_2735,N_2899);
and U3203 (N_3203,N_2760,N_2694);
and U3204 (N_3204,N_2902,N_2785);
or U3205 (N_3205,N_2681,N_2556);
nor U3206 (N_3206,N_2790,N_2812);
nor U3207 (N_3207,N_2526,N_2632);
and U3208 (N_3208,N_2627,N_2551);
or U3209 (N_3209,N_2511,N_2636);
or U3210 (N_3210,N_2643,N_2618);
and U3211 (N_3211,N_2633,N_2660);
nor U3212 (N_3212,N_2808,N_2652);
or U3213 (N_3213,N_2999,N_2807);
nand U3214 (N_3214,N_2640,N_2602);
nor U3215 (N_3215,N_2680,N_2535);
or U3216 (N_3216,N_2746,N_2911);
nand U3217 (N_3217,N_2850,N_2747);
and U3218 (N_3218,N_2820,N_2598);
nor U3219 (N_3219,N_2542,N_2731);
or U3220 (N_3220,N_2831,N_2941);
nor U3221 (N_3221,N_2733,N_2926);
and U3222 (N_3222,N_2814,N_2757);
nand U3223 (N_3223,N_2748,N_2658);
or U3224 (N_3224,N_2945,N_2803);
nor U3225 (N_3225,N_2622,N_2701);
and U3226 (N_3226,N_2751,N_2544);
and U3227 (N_3227,N_2792,N_2925);
nand U3228 (N_3228,N_2929,N_2728);
nor U3229 (N_3229,N_2796,N_2976);
or U3230 (N_3230,N_2861,N_2631);
and U3231 (N_3231,N_2777,N_2678);
nand U3232 (N_3232,N_2572,N_2890);
nand U3233 (N_3233,N_2657,N_2763);
or U3234 (N_3234,N_2768,N_2845);
nand U3235 (N_3235,N_2867,N_2692);
nand U3236 (N_3236,N_2606,N_2553);
and U3237 (N_3237,N_2865,N_2656);
nand U3238 (N_3238,N_2873,N_2954);
nor U3239 (N_3239,N_2589,N_2539);
or U3240 (N_3240,N_2609,N_2712);
nor U3241 (N_3241,N_2557,N_2667);
or U3242 (N_3242,N_2703,N_2958);
nor U3243 (N_3243,N_2775,N_2592);
nand U3244 (N_3244,N_2900,N_2878);
and U3245 (N_3245,N_2647,N_2696);
nand U3246 (N_3246,N_2709,N_2896);
nand U3247 (N_3247,N_2546,N_2893);
nand U3248 (N_3248,N_2914,N_2801);
and U3249 (N_3249,N_2827,N_2581);
nor U3250 (N_3250,N_2737,N_2597);
and U3251 (N_3251,N_2805,N_2678);
or U3252 (N_3252,N_2827,N_2844);
nor U3253 (N_3253,N_2620,N_2538);
and U3254 (N_3254,N_2749,N_2705);
nor U3255 (N_3255,N_2933,N_2553);
nand U3256 (N_3256,N_2538,N_2909);
nand U3257 (N_3257,N_2792,N_2949);
nand U3258 (N_3258,N_2752,N_2993);
nand U3259 (N_3259,N_2877,N_2510);
or U3260 (N_3260,N_2729,N_2920);
or U3261 (N_3261,N_2872,N_2807);
nand U3262 (N_3262,N_2637,N_2688);
and U3263 (N_3263,N_2694,N_2601);
or U3264 (N_3264,N_2951,N_2703);
nor U3265 (N_3265,N_2654,N_2758);
nor U3266 (N_3266,N_2996,N_2645);
or U3267 (N_3267,N_2601,N_2739);
nor U3268 (N_3268,N_2778,N_2560);
nor U3269 (N_3269,N_2724,N_2569);
and U3270 (N_3270,N_2753,N_2534);
nand U3271 (N_3271,N_2696,N_2989);
or U3272 (N_3272,N_2897,N_2594);
nor U3273 (N_3273,N_2755,N_2663);
or U3274 (N_3274,N_2944,N_2732);
and U3275 (N_3275,N_2686,N_2772);
nand U3276 (N_3276,N_2883,N_2722);
and U3277 (N_3277,N_2590,N_2956);
nand U3278 (N_3278,N_2648,N_2535);
nand U3279 (N_3279,N_2854,N_2565);
nand U3280 (N_3280,N_2529,N_2842);
nor U3281 (N_3281,N_2663,N_2516);
nand U3282 (N_3282,N_2503,N_2832);
nor U3283 (N_3283,N_2824,N_2626);
nand U3284 (N_3284,N_2685,N_2830);
nand U3285 (N_3285,N_2584,N_2932);
nand U3286 (N_3286,N_2575,N_2705);
nand U3287 (N_3287,N_2806,N_2714);
nor U3288 (N_3288,N_2615,N_2648);
and U3289 (N_3289,N_2823,N_2907);
or U3290 (N_3290,N_2910,N_2683);
and U3291 (N_3291,N_2523,N_2822);
nor U3292 (N_3292,N_2536,N_2696);
or U3293 (N_3293,N_2661,N_2833);
or U3294 (N_3294,N_2576,N_2903);
nor U3295 (N_3295,N_2927,N_2564);
or U3296 (N_3296,N_2590,N_2651);
xnor U3297 (N_3297,N_2779,N_2552);
nand U3298 (N_3298,N_2710,N_2674);
nand U3299 (N_3299,N_2883,N_2522);
nand U3300 (N_3300,N_2915,N_2855);
or U3301 (N_3301,N_2764,N_2679);
nand U3302 (N_3302,N_2810,N_2651);
nand U3303 (N_3303,N_2940,N_2650);
nand U3304 (N_3304,N_2859,N_2609);
or U3305 (N_3305,N_2647,N_2995);
or U3306 (N_3306,N_2763,N_2642);
or U3307 (N_3307,N_2992,N_2804);
nand U3308 (N_3308,N_2927,N_2567);
and U3309 (N_3309,N_2677,N_2567);
and U3310 (N_3310,N_2826,N_2830);
nor U3311 (N_3311,N_2672,N_2620);
and U3312 (N_3312,N_2657,N_2642);
nand U3313 (N_3313,N_2522,N_2848);
nor U3314 (N_3314,N_2513,N_2697);
nand U3315 (N_3315,N_2653,N_2968);
or U3316 (N_3316,N_2596,N_2666);
or U3317 (N_3317,N_2574,N_2733);
nor U3318 (N_3318,N_2656,N_2726);
nor U3319 (N_3319,N_2604,N_2573);
and U3320 (N_3320,N_2757,N_2689);
and U3321 (N_3321,N_2841,N_2917);
or U3322 (N_3322,N_2635,N_2654);
nor U3323 (N_3323,N_2739,N_2988);
and U3324 (N_3324,N_2548,N_2955);
nand U3325 (N_3325,N_2621,N_2810);
and U3326 (N_3326,N_2707,N_2503);
or U3327 (N_3327,N_2525,N_2914);
or U3328 (N_3328,N_2596,N_2797);
nor U3329 (N_3329,N_2621,N_2793);
and U3330 (N_3330,N_2954,N_2784);
nor U3331 (N_3331,N_2574,N_2906);
and U3332 (N_3332,N_2503,N_2619);
or U3333 (N_3333,N_2743,N_2984);
nand U3334 (N_3334,N_2734,N_2701);
or U3335 (N_3335,N_2700,N_2939);
nand U3336 (N_3336,N_2802,N_2821);
and U3337 (N_3337,N_2922,N_2907);
nor U3338 (N_3338,N_2952,N_2807);
or U3339 (N_3339,N_2697,N_2574);
nand U3340 (N_3340,N_2977,N_2652);
and U3341 (N_3341,N_2892,N_2557);
and U3342 (N_3342,N_2885,N_2613);
nor U3343 (N_3343,N_2789,N_2958);
nand U3344 (N_3344,N_2731,N_2745);
and U3345 (N_3345,N_2690,N_2805);
nand U3346 (N_3346,N_2817,N_2974);
and U3347 (N_3347,N_2779,N_2777);
nor U3348 (N_3348,N_2739,N_2819);
and U3349 (N_3349,N_2913,N_2868);
nand U3350 (N_3350,N_2973,N_2649);
nor U3351 (N_3351,N_2971,N_2730);
nand U3352 (N_3352,N_2826,N_2997);
and U3353 (N_3353,N_2940,N_2960);
xor U3354 (N_3354,N_2702,N_2603);
and U3355 (N_3355,N_2729,N_2916);
or U3356 (N_3356,N_2774,N_2948);
nor U3357 (N_3357,N_2645,N_2701);
or U3358 (N_3358,N_2530,N_2834);
nand U3359 (N_3359,N_2866,N_2659);
nand U3360 (N_3360,N_2871,N_2905);
and U3361 (N_3361,N_2666,N_2891);
nand U3362 (N_3362,N_2585,N_2981);
and U3363 (N_3363,N_2674,N_2867);
nor U3364 (N_3364,N_2589,N_2648);
and U3365 (N_3365,N_2753,N_2948);
or U3366 (N_3366,N_2535,N_2994);
and U3367 (N_3367,N_2934,N_2930);
nand U3368 (N_3368,N_2850,N_2525);
or U3369 (N_3369,N_2874,N_2939);
and U3370 (N_3370,N_2577,N_2968);
or U3371 (N_3371,N_2859,N_2667);
and U3372 (N_3372,N_2978,N_2941);
nor U3373 (N_3373,N_2614,N_2804);
nor U3374 (N_3374,N_2810,N_2865);
and U3375 (N_3375,N_2675,N_2584);
nand U3376 (N_3376,N_2906,N_2684);
nand U3377 (N_3377,N_2853,N_2790);
and U3378 (N_3378,N_2692,N_2669);
nand U3379 (N_3379,N_2520,N_2588);
nor U3380 (N_3380,N_2621,N_2868);
nor U3381 (N_3381,N_2934,N_2580);
nor U3382 (N_3382,N_2844,N_2955);
nor U3383 (N_3383,N_2764,N_2864);
nand U3384 (N_3384,N_2550,N_2528);
and U3385 (N_3385,N_2841,N_2834);
xor U3386 (N_3386,N_2557,N_2622);
or U3387 (N_3387,N_2980,N_2945);
and U3388 (N_3388,N_2892,N_2532);
nand U3389 (N_3389,N_2963,N_2594);
and U3390 (N_3390,N_2903,N_2829);
and U3391 (N_3391,N_2703,N_2809);
and U3392 (N_3392,N_2758,N_2656);
nand U3393 (N_3393,N_2609,N_2795);
and U3394 (N_3394,N_2927,N_2537);
nor U3395 (N_3395,N_2711,N_2660);
and U3396 (N_3396,N_2561,N_2724);
and U3397 (N_3397,N_2725,N_2983);
nor U3398 (N_3398,N_2643,N_2833);
nand U3399 (N_3399,N_2697,N_2749);
and U3400 (N_3400,N_2649,N_2724);
nor U3401 (N_3401,N_2520,N_2954);
nor U3402 (N_3402,N_2939,N_2504);
xor U3403 (N_3403,N_2823,N_2688);
or U3404 (N_3404,N_2988,N_2547);
nor U3405 (N_3405,N_2555,N_2704);
or U3406 (N_3406,N_2820,N_2512);
and U3407 (N_3407,N_2625,N_2764);
nand U3408 (N_3408,N_2633,N_2538);
xor U3409 (N_3409,N_2873,N_2906);
or U3410 (N_3410,N_2931,N_2744);
or U3411 (N_3411,N_2814,N_2984);
and U3412 (N_3412,N_2694,N_2562);
nand U3413 (N_3413,N_2805,N_2731);
nor U3414 (N_3414,N_2921,N_2757);
and U3415 (N_3415,N_2645,N_2987);
or U3416 (N_3416,N_2534,N_2916);
nand U3417 (N_3417,N_2631,N_2666);
or U3418 (N_3418,N_2710,N_2939);
nor U3419 (N_3419,N_2763,N_2767);
and U3420 (N_3420,N_2556,N_2692);
xor U3421 (N_3421,N_2907,N_2635);
and U3422 (N_3422,N_2939,N_2801);
or U3423 (N_3423,N_2667,N_2611);
nor U3424 (N_3424,N_2542,N_2986);
and U3425 (N_3425,N_2692,N_2578);
nand U3426 (N_3426,N_2971,N_2791);
or U3427 (N_3427,N_2680,N_2881);
nor U3428 (N_3428,N_2953,N_2980);
nor U3429 (N_3429,N_2554,N_2505);
nor U3430 (N_3430,N_2659,N_2682);
or U3431 (N_3431,N_2846,N_2924);
or U3432 (N_3432,N_2727,N_2707);
nor U3433 (N_3433,N_2770,N_2568);
nand U3434 (N_3434,N_2732,N_2898);
nor U3435 (N_3435,N_2758,N_2796);
and U3436 (N_3436,N_2918,N_2687);
or U3437 (N_3437,N_2978,N_2781);
nor U3438 (N_3438,N_2535,N_2807);
nand U3439 (N_3439,N_2705,N_2755);
nand U3440 (N_3440,N_2646,N_2827);
nand U3441 (N_3441,N_2556,N_2770);
nand U3442 (N_3442,N_2726,N_2644);
or U3443 (N_3443,N_2975,N_2551);
xor U3444 (N_3444,N_2715,N_2776);
nor U3445 (N_3445,N_2661,N_2752);
or U3446 (N_3446,N_2839,N_2975);
nor U3447 (N_3447,N_2830,N_2601);
and U3448 (N_3448,N_2777,N_2756);
or U3449 (N_3449,N_2879,N_2767);
nor U3450 (N_3450,N_2671,N_2863);
nand U3451 (N_3451,N_2739,N_2958);
nand U3452 (N_3452,N_2767,N_2672);
and U3453 (N_3453,N_2995,N_2607);
nand U3454 (N_3454,N_2570,N_2732);
and U3455 (N_3455,N_2650,N_2527);
or U3456 (N_3456,N_2965,N_2696);
nand U3457 (N_3457,N_2980,N_2914);
xnor U3458 (N_3458,N_2500,N_2709);
and U3459 (N_3459,N_2685,N_2826);
and U3460 (N_3460,N_2925,N_2511);
and U3461 (N_3461,N_2695,N_2522);
nor U3462 (N_3462,N_2994,N_2630);
and U3463 (N_3463,N_2799,N_2898);
and U3464 (N_3464,N_2750,N_2581);
nor U3465 (N_3465,N_2976,N_2933);
or U3466 (N_3466,N_2643,N_2837);
nor U3467 (N_3467,N_2531,N_2953);
and U3468 (N_3468,N_2501,N_2594);
and U3469 (N_3469,N_2593,N_2749);
nand U3470 (N_3470,N_2833,N_2895);
and U3471 (N_3471,N_2972,N_2608);
nor U3472 (N_3472,N_2523,N_2999);
or U3473 (N_3473,N_2661,N_2836);
or U3474 (N_3474,N_2789,N_2592);
nand U3475 (N_3475,N_2930,N_2703);
or U3476 (N_3476,N_2561,N_2619);
and U3477 (N_3477,N_2770,N_2572);
and U3478 (N_3478,N_2545,N_2713);
or U3479 (N_3479,N_2748,N_2500);
nand U3480 (N_3480,N_2944,N_2990);
nand U3481 (N_3481,N_2702,N_2988);
nand U3482 (N_3482,N_2669,N_2974);
nor U3483 (N_3483,N_2519,N_2548);
and U3484 (N_3484,N_2961,N_2983);
or U3485 (N_3485,N_2738,N_2835);
and U3486 (N_3486,N_2823,N_2629);
and U3487 (N_3487,N_2986,N_2989);
nor U3488 (N_3488,N_2556,N_2848);
and U3489 (N_3489,N_2639,N_2822);
nor U3490 (N_3490,N_2546,N_2835);
nor U3491 (N_3491,N_2671,N_2715);
nand U3492 (N_3492,N_2967,N_2527);
nand U3493 (N_3493,N_2720,N_2872);
nand U3494 (N_3494,N_2560,N_2747);
nand U3495 (N_3495,N_2712,N_2998);
nand U3496 (N_3496,N_2590,N_2679);
nor U3497 (N_3497,N_2954,N_2662);
and U3498 (N_3498,N_2674,N_2754);
and U3499 (N_3499,N_2550,N_2963);
nand U3500 (N_3500,N_3013,N_3160);
and U3501 (N_3501,N_3217,N_3048);
nor U3502 (N_3502,N_3211,N_3359);
nand U3503 (N_3503,N_3427,N_3260);
nand U3504 (N_3504,N_3283,N_3207);
and U3505 (N_3505,N_3370,N_3313);
nand U3506 (N_3506,N_3125,N_3090);
and U3507 (N_3507,N_3096,N_3183);
nand U3508 (N_3508,N_3055,N_3018);
nand U3509 (N_3509,N_3146,N_3153);
or U3510 (N_3510,N_3488,N_3097);
and U3511 (N_3511,N_3155,N_3021);
or U3512 (N_3512,N_3367,N_3496);
and U3513 (N_3513,N_3280,N_3400);
nand U3514 (N_3514,N_3420,N_3466);
nand U3515 (N_3515,N_3034,N_3042);
nand U3516 (N_3516,N_3103,N_3452);
and U3517 (N_3517,N_3429,N_3343);
and U3518 (N_3518,N_3123,N_3324);
and U3519 (N_3519,N_3286,N_3059);
nand U3520 (N_3520,N_3356,N_3479);
nand U3521 (N_3521,N_3043,N_3263);
and U3522 (N_3522,N_3027,N_3381);
and U3523 (N_3523,N_3223,N_3349);
or U3524 (N_3524,N_3181,N_3205);
nor U3525 (N_3525,N_3032,N_3242);
and U3526 (N_3526,N_3285,N_3179);
or U3527 (N_3527,N_3212,N_3172);
or U3528 (N_3528,N_3082,N_3432);
or U3529 (N_3529,N_3053,N_3386);
nor U3530 (N_3530,N_3354,N_3317);
and U3531 (N_3531,N_3455,N_3133);
and U3532 (N_3532,N_3255,N_3341);
nand U3533 (N_3533,N_3041,N_3281);
nand U3534 (N_3534,N_3312,N_3063);
nand U3535 (N_3535,N_3150,N_3166);
or U3536 (N_3536,N_3065,N_3014);
xor U3537 (N_3537,N_3306,N_3143);
nor U3538 (N_3538,N_3029,N_3112);
nor U3539 (N_3539,N_3483,N_3372);
nor U3540 (N_3540,N_3373,N_3028);
or U3541 (N_3541,N_3089,N_3136);
and U3542 (N_3542,N_3377,N_3336);
or U3543 (N_3543,N_3406,N_3025);
nand U3544 (N_3544,N_3239,N_3450);
nor U3545 (N_3545,N_3363,N_3469);
nor U3546 (N_3546,N_3291,N_3492);
nand U3547 (N_3547,N_3338,N_3438);
nor U3548 (N_3548,N_3056,N_3031);
xnor U3549 (N_3549,N_3494,N_3320);
or U3550 (N_3550,N_3376,N_3011);
nand U3551 (N_3551,N_3099,N_3246);
and U3552 (N_3552,N_3221,N_3006);
and U3553 (N_3553,N_3075,N_3110);
nor U3554 (N_3554,N_3241,N_3010);
and U3555 (N_3555,N_3148,N_3319);
or U3556 (N_3556,N_3062,N_3094);
nor U3557 (N_3557,N_3194,N_3297);
and U3558 (N_3558,N_3098,N_3084);
and U3559 (N_3559,N_3325,N_3451);
nand U3560 (N_3560,N_3463,N_3487);
and U3561 (N_3561,N_3135,N_3300);
nand U3562 (N_3562,N_3039,N_3277);
nand U3563 (N_3563,N_3446,N_3137);
and U3564 (N_3564,N_3149,N_3460);
nand U3565 (N_3565,N_3269,N_3440);
nor U3566 (N_3566,N_3301,N_3220);
or U3567 (N_3567,N_3173,N_3392);
and U3568 (N_3568,N_3001,N_3276);
and U3569 (N_3569,N_3165,N_3379);
and U3570 (N_3570,N_3293,N_3215);
or U3571 (N_3571,N_3000,N_3424);
nand U3572 (N_3572,N_3201,N_3131);
and U3573 (N_3573,N_3154,N_3050);
or U3574 (N_3574,N_3468,N_3493);
nand U3575 (N_3575,N_3247,N_3298);
or U3576 (N_3576,N_3200,N_3401);
or U3577 (N_3577,N_3348,N_3362);
nand U3578 (N_3578,N_3433,N_3475);
and U3579 (N_3579,N_3045,N_3422);
or U3580 (N_3580,N_3250,N_3107);
nand U3581 (N_3581,N_3193,N_3345);
nand U3582 (N_3582,N_3169,N_3405);
nor U3583 (N_3583,N_3282,N_3270);
or U3584 (N_3584,N_3157,N_3161);
and U3585 (N_3585,N_3016,N_3295);
and U3586 (N_3586,N_3151,N_3278);
nand U3587 (N_3587,N_3156,N_3311);
or U3588 (N_3588,N_3419,N_3374);
and U3589 (N_3589,N_3403,N_3116);
or U3590 (N_3590,N_3275,N_3326);
nor U3591 (N_3591,N_3396,N_3478);
nor U3592 (N_3592,N_3369,N_3458);
nor U3593 (N_3593,N_3104,N_3252);
nand U3594 (N_3594,N_3497,N_3120);
nor U3595 (N_3595,N_3020,N_3476);
and U3596 (N_3596,N_3304,N_3289);
nor U3597 (N_3597,N_3368,N_3233);
and U3598 (N_3598,N_3329,N_3076);
and U3599 (N_3599,N_3393,N_3431);
nor U3600 (N_3600,N_3257,N_3002);
nand U3601 (N_3601,N_3078,N_3421);
nor U3602 (N_3602,N_3178,N_3414);
nand U3603 (N_3603,N_3266,N_3038);
nand U3604 (N_3604,N_3232,N_3184);
nand U3605 (N_3605,N_3117,N_3287);
nand U3606 (N_3606,N_3017,N_3391);
and U3607 (N_3607,N_3334,N_3108);
nor U3608 (N_3608,N_3327,N_3259);
nor U3609 (N_3609,N_3482,N_3077);
or U3610 (N_3610,N_3115,N_3477);
nor U3611 (N_3611,N_3256,N_3410);
nor U3612 (N_3612,N_3267,N_3088);
and U3613 (N_3613,N_3397,N_3404);
or U3614 (N_3614,N_3339,N_3170);
and U3615 (N_3615,N_3037,N_3079);
or U3616 (N_3616,N_3198,N_3457);
nand U3617 (N_3617,N_3331,N_3105);
nor U3618 (N_3618,N_3127,N_3132);
xnor U3619 (N_3619,N_3176,N_3484);
and U3620 (N_3620,N_3271,N_3413);
nand U3621 (N_3621,N_3360,N_3005);
or U3622 (N_3622,N_3191,N_3465);
or U3623 (N_3623,N_3353,N_3265);
nor U3624 (N_3624,N_3185,N_3129);
nand U3625 (N_3625,N_3204,N_3192);
or U3626 (N_3626,N_3399,N_3310);
nor U3627 (N_3627,N_3113,N_3385);
or U3628 (N_3628,N_3441,N_3294);
and U3629 (N_3629,N_3224,N_3321);
nand U3630 (N_3630,N_3187,N_3174);
and U3631 (N_3631,N_3245,N_3142);
nand U3632 (N_3632,N_3315,N_3425);
xnor U3633 (N_3633,N_3430,N_3415);
or U3634 (N_3634,N_3064,N_3305);
or U3635 (N_3635,N_3009,N_3340);
nand U3636 (N_3636,N_3019,N_3426);
or U3637 (N_3637,N_3122,N_3248);
and U3638 (N_3638,N_3357,N_3308);
nor U3639 (N_3639,N_3057,N_3251);
and U3640 (N_3640,N_3060,N_3051);
or U3641 (N_3641,N_3471,N_3109);
nor U3642 (N_3642,N_3118,N_3126);
or U3643 (N_3643,N_3024,N_3086);
and U3644 (N_3644,N_3499,N_3459);
nand U3645 (N_3645,N_3383,N_3302);
or U3646 (N_3646,N_3296,N_3012);
nand U3647 (N_3647,N_3054,N_3080);
or U3648 (N_3648,N_3180,N_3417);
nor U3649 (N_3649,N_3159,N_3008);
nor U3650 (N_3650,N_3238,N_3316);
nor U3651 (N_3651,N_3114,N_3299);
nor U3652 (N_3652,N_3490,N_3412);
or U3653 (N_3653,N_3498,N_3047);
nor U3654 (N_3654,N_3249,N_3030);
nand U3655 (N_3655,N_3456,N_3309);
nand U3656 (N_3656,N_3230,N_3070);
or U3657 (N_3657,N_3290,N_3095);
nor U3658 (N_3658,N_3167,N_3485);
or U3659 (N_3659,N_3163,N_3445);
and U3660 (N_3660,N_3144,N_3213);
nand U3661 (N_3661,N_3408,N_3342);
nor U3662 (N_3662,N_3140,N_3480);
nor U3663 (N_3663,N_3145,N_3330);
or U3664 (N_3664,N_3323,N_3371);
nor U3665 (N_3665,N_3168,N_3284);
nor U3666 (N_3666,N_3467,N_3052);
and U3667 (N_3667,N_3226,N_3219);
or U3668 (N_3668,N_3394,N_3346);
and U3669 (N_3669,N_3128,N_3272);
nand U3670 (N_3670,N_3350,N_3100);
nand U3671 (N_3671,N_3264,N_3073);
nand U3672 (N_3672,N_3022,N_3111);
nand U3673 (N_3673,N_3210,N_3378);
or U3674 (N_3674,N_3453,N_3489);
or U3675 (N_3675,N_3454,N_3069);
and U3676 (N_3676,N_3058,N_3402);
and U3677 (N_3677,N_3119,N_3152);
nor U3678 (N_3678,N_3328,N_3288);
and U3679 (N_3679,N_3365,N_3186);
and U3680 (N_3680,N_3416,N_3244);
nand U3681 (N_3681,N_3398,N_3081);
and U3682 (N_3682,N_3481,N_3189);
nand U3683 (N_3683,N_3225,N_3448);
and U3684 (N_3684,N_3007,N_3208);
or U3685 (N_3685,N_3472,N_3067);
nand U3686 (N_3686,N_3361,N_3102);
and U3687 (N_3687,N_3093,N_3202);
nand U3688 (N_3688,N_3380,N_3411);
or U3689 (N_3689,N_3423,N_3375);
and U3690 (N_3690,N_3307,N_3209);
nand U3691 (N_3691,N_3087,N_3407);
or U3692 (N_3692,N_3390,N_3382);
and U3693 (N_3693,N_3046,N_3439);
nand U3694 (N_3694,N_3253,N_3083);
or U3695 (N_3695,N_3214,N_3106);
or U3696 (N_3696,N_3072,N_3061);
nand U3697 (N_3697,N_3358,N_3437);
or U3698 (N_3698,N_3121,N_3033);
nor U3699 (N_3699,N_3387,N_3206);
nor U3700 (N_3700,N_3388,N_3227);
or U3701 (N_3701,N_3464,N_3395);
and U3702 (N_3702,N_3344,N_3162);
and U3703 (N_3703,N_3495,N_3332);
nor U3704 (N_3704,N_3337,N_3101);
nor U3705 (N_3705,N_3199,N_3234);
and U3706 (N_3706,N_3138,N_3442);
nand U3707 (N_3707,N_3462,N_3236);
nand U3708 (N_3708,N_3347,N_3074);
nand U3709 (N_3709,N_3436,N_3461);
and U3710 (N_3710,N_3351,N_3071);
nor U3711 (N_3711,N_3092,N_3218);
xor U3712 (N_3712,N_3085,N_3254);
and U3713 (N_3713,N_3040,N_3314);
nand U3714 (N_3714,N_3182,N_3164);
nor U3715 (N_3715,N_3262,N_3384);
nor U3716 (N_3716,N_3231,N_3486);
and U3717 (N_3717,N_3023,N_3261);
nand U3718 (N_3718,N_3222,N_3258);
nor U3719 (N_3719,N_3279,N_3273);
nand U3720 (N_3720,N_3229,N_3470);
and U3721 (N_3721,N_3243,N_3139);
and U3722 (N_3722,N_3196,N_3158);
nor U3723 (N_3723,N_3091,N_3364);
and U3724 (N_3724,N_3352,N_3333);
nor U3725 (N_3725,N_3292,N_3355);
or U3726 (N_3726,N_3235,N_3175);
or U3727 (N_3727,N_3274,N_3444);
nand U3728 (N_3728,N_3409,N_3068);
nand U3729 (N_3729,N_3268,N_3237);
nand U3730 (N_3730,N_3447,N_3335);
nor U3731 (N_3731,N_3443,N_3195);
and U3732 (N_3732,N_3171,N_3389);
nand U3733 (N_3733,N_3026,N_3228);
nor U3734 (N_3734,N_3015,N_3035);
nand U3735 (N_3735,N_3004,N_3190);
nand U3736 (N_3736,N_3418,N_3197);
nand U3737 (N_3737,N_3044,N_3318);
or U3738 (N_3738,N_3240,N_3434);
and U3739 (N_3739,N_3449,N_3066);
nand U3740 (N_3740,N_3036,N_3124);
nor U3741 (N_3741,N_3130,N_3177);
nand U3742 (N_3742,N_3147,N_3203);
or U3743 (N_3743,N_3473,N_3003);
and U3744 (N_3744,N_3474,N_3366);
nor U3745 (N_3745,N_3303,N_3428);
and U3746 (N_3746,N_3049,N_3216);
nor U3747 (N_3747,N_3134,N_3491);
or U3748 (N_3748,N_3322,N_3141);
nand U3749 (N_3749,N_3188,N_3435);
nor U3750 (N_3750,N_3461,N_3449);
and U3751 (N_3751,N_3340,N_3422);
and U3752 (N_3752,N_3212,N_3488);
nor U3753 (N_3753,N_3057,N_3030);
or U3754 (N_3754,N_3154,N_3301);
or U3755 (N_3755,N_3142,N_3193);
nand U3756 (N_3756,N_3324,N_3236);
xnor U3757 (N_3757,N_3491,N_3433);
nand U3758 (N_3758,N_3266,N_3042);
and U3759 (N_3759,N_3448,N_3199);
or U3760 (N_3760,N_3033,N_3254);
nor U3761 (N_3761,N_3431,N_3492);
nand U3762 (N_3762,N_3382,N_3020);
and U3763 (N_3763,N_3332,N_3117);
or U3764 (N_3764,N_3013,N_3067);
nand U3765 (N_3765,N_3056,N_3012);
and U3766 (N_3766,N_3295,N_3340);
xnor U3767 (N_3767,N_3433,N_3497);
and U3768 (N_3768,N_3401,N_3148);
and U3769 (N_3769,N_3406,N_3451);
nor U3770 (N_3770,N_3427,N_3097);
and U3771 (N_3771,N_3238,N_3272);
and U3772 (N_3772,N_3082,N_3335);
xnor U3773 (N_3773,N_3014,N_3079);
or U3774 (N_3774,N_3358,N_3309);
and U3775 (N_3775,N_3182,N_3279);
nand U3776 (N_3776,N_3161,N_3415);
or U3777 (N_3777,N_3016,N_3270);
nand U3778 (N_3778,N_3416,N_3449);
nand U3779 (N_3779,N_3383,N_3221);
nor U3780 (N_3780,N_3193,N_3127);
and U3781 (N_3781,N_3301,N_3358);
and U3782 (N_3782,N_3166,N_3106);
and U3783 (N_3783,N_3488,N_3166);
or U3784 (N_3784,N_3388,N_3312);
and U3785 (N_3785,N_3122,N_3428);
nor U3786 (N_3786,N_3053,N_3480);
or U3787 (N_3787,N_3305,N_3010);
and U3788 (N_3788,N_3340,N_3228);
nand U3789 (N_3789,N_3143,N_3426);
and U3790 (N_3790,N_3061,N_3273);
nand U3791 (N_3791,N_3386,N_3213);
nand U3792 (N_3792,N_3213,N_3348);
and U3793 (N_3793,N_3095,N_3000);
and U3794 (N_3794,N_3114,N_3034);
nor U3795 (N_3795,N_3021,N_3316);
or U3796 (N_3796,N_3347,N_3442);
and U3797 (N_3797,N_3034,N_3221);
or U3798 (N_3798,N_3439,N_3324);
or U3799 (N_3799,N_3396,N_3287);
and U3800 (N_3800,N_3441,N_3031);
and U3801 (N_3801,N_3440,N_3458);
and U3802 (N_3802,N_3402,N_3073);
and U3803 (N_3803,N_3183,N_3304);
or U3804 (N_3804,N_3386,N_3332);
nand U3805 (N_3805,N_3366,N_3240);
nor U3806 (N_3806,N_3199,N_3092);
nand U3807 (N_3807,N_3153,N_3221);
nor U3808 (N_3808,N_3210,N_3161);
nor U3809 (N_3809,N_3097,N_3319);
nor U3810 (N_3810,N_3287,N_3305);
or U3811 (N_3811,N_3345,N_3251);
nor U3812 (N_3812,N_3236,N_3310);
or U3813 (N_3813,N_3461,N_3432);
nor U3814 (N_3814,N_3231,N_3465);
nand U3815 (N_3815,N_3260,N_3113);
nor U3816 (N_3816,N_3378,N_3287);
nand U3817 (N_3817,N_3313,N_3401);
nand U3818 (N_3818,N_3048,N_3275);
nor U3819 (N_3819,N_3146,N_3366);
and U3820 (N_3820,N_3483,N_3039);
or U3821 (N_3821,N_3137,N_3376);
and U3822 (N_3822,N_3111,N_3278);
nand U3823 (N_3823,N_3151,N_3158);
and U3824 (N_3824,N_3488,N_3342);
nand U3825 (N_3825,N_3422,N_3451);
nor U3826 (N_3826,N_3452,N_3201);
nor U3827 (N_3827,N_3215,N_3091);
nor U3828 (N_3828,N_3414,N_3001);
nor U3829 (N_3829,N_3264,N_3236);
or U3830 (N_3830,N_3165,N_3181);
nand U3831 (N_3831,N_3107,N_3432);
nand U3832 (N_3832,N_3270,N_3303);
nor U3833 (N_3833,N_3459,N_3144);
or U3834 (N_3834,N_3109,N_3074);
nand U3835 (N_3835,N_3016,N_3172);
nor U3836 (N_3836,N_3232,N_3273);
nor U3837 (N_3837,N_3052,N_3134);
and U3838 (N_3838,N_3371,N_3004);
or U3839 (N_3839,N_3143,N_3065);
nand U3840 (N_3840,N_3109,N_3350);
nand U3841 (N_3841,N_3492,N_3459);
nor U3842 (N_3842,N_3072,N_3015);
nand U3843 (N_3843,N_3362,N_3364);
or U3844 (N_3844,N_3199,N_3271);
or U3845 (N_3845,N_3445,N_3437);
and U3846 (N_3846,N_3293,N_3431);
and U3847 (N_3847,N_3151,N_3456);
or U3848 (N_3848,N_3483,N_3115);
nor U3849 (N_3849,N_3357,N_3067);
nor U3850 (N_3850,N_3325,N_3195);
and U3851 (N_3851,N_3161,N_3356);
and U3852 (N_3852,N_3028,N_3361);
and U3853 (N_3853,N_3061,N_3036);
and U3854 (N_3854,N_3135,N_3086);
or U3855 (N_3855,N_3029,N_3391);
nand U3856 (N_3856,N_3170,N_3043);
and U3857 (N_3857,N_3499,N_3102);
or U3858 (N_3858,N_3487,N_3156);
nand U3859 (N_3859,N_3408,N_3112);
xnor U3860 (N_3860,N_3227,N_3133);
xnor U3861 (N_3861,N_3449,N_3374);
nand U3862 (N_3862,N_3054,N_3162);
and U3863 (N_3863,N_3177,N_3285);
nor U3864 (N_3864,N_3000,N_3208);
or U3865 (N_3865,N_3300,N_3241);
nor U3866 (N_3866,N_3380,N_3425);
and U3867 (N_3867,N_3167,N_3395);
or U3868 (N_3868,N_3142,N_3408);
and U3869 (N_3869,N_3087,N_3339);
nor U3870 (N_3870,N_3070,N_3013);
or U3871 (N_3871,N_3108,N_3075);
nand U3872 (N_3872,N_3442,N_3325);
nor U3873 (N_3873,N_3049,N_3232);
or U3874 (N_3874,N_3005,N_3453);
or U3875 (N_3875,N_3459,N_3057);
and U3876 (N_3876,N_3484,N_3048);
or U3877 (N_3877,N_3035,N_3095);
and U3878 (N_3878,N_3322,N_3369);
nor U3879 (N_3879,N_3182,N_3226);
or U3880 (N_3880,N_3397,N_3307);
and U3881 (N_3881,N_3169,N_3016);
nor U3882 (N_3882,N_3180,N_3317);
and U3883 (N_3883,N_3447,N_3196);
and U3884 (N_3884,N_3392,N_3270);
nand U3885 (N_3885,N_3278,N_3056);
or U3886 (N_3886,N_3240,N_3070);
nand U3887 (N_3887,N_3255,N_3301);
nor U3888 (N_3888,N_3414,N_3113);
nor U3889 (N_3889,N_3451,N_3315);
or U3890 (N_3890,N_3186,N_3333);
nand U3891 (N_3891,N_3451,N_3139);
nand U3892 (N_3892,N_3242,N_3485);
nand U3893 (N_3893,N_3138,N_3017);
or U3894 (N_3894,N_3459,N_3408);
or U3895 (N_3895,N_3059,N_3349);
nand U3896 (N_3896,N_3209,N_3180);
or U3897 (N_3897,N_3361,N_3081);
and U3898 (N_3898,N_3135,N_3472);
and U3899 (N_3899,N_3062,N_3449);
nor U3900 (N_3900,N_3021,N_3466);
or U3901 (N_3901,N_3047,N_3189);
nand U3902 (N_3902,N_3194,N_3025);
nor U3903 (N_3903,N_3476,N_3069);
nor U3904 (N_3904,N_3461,N_3396);
xnor U3905 (N_3905,N_3061,N_3264);
or U3906 (N_3906,N_3309,N_3327);
nor U3907 (N_3907,N_3007,N_3008);
nor U3908 (N_3908,N_3250,N_3468);
or U3909 (N_3909,N_3343,N_3000);
nand U3910 (N_3910,N_3181,N_3358);
nor U3911 (N_3911,N_3054,N_3241);
xnor U3912 (N_3912,N_3073,N_3437);
nor U3913 (N_3913,N_3389,N_3330);
nor U3914 (N_3914,N_3130,N_3337);
and U3915 (N_3915,N_3498,N_3259);
nor U3916 (N_3916,N_3190,N_3446);
nor U3917 (N_3917,N_3338,N_3065);
and U3918 (N_3918,N_3411,N_3014);
nor U3919 (N_3919,N_3444,N_3386);
nor U3920 (N_3920,N_3288,N_3253);
nor U3921 (N_3921,N_3114,N_3414);
or U3922 (N_3922,N_3297,N_3211);
nand U3923 (N_3923,N_3020,N_3477);
nor U3924 (N_3924,N_3479,N_3061);
and U3925 (N_3925,N_3068,N_3386);
nand U3926 (N_3926,N_3347,N_3336);
nand U3927 (N_3927,N_3040,N_3007);
nand U3928 (N_3928,N_3369,N_3491);
or U3929 (N_3929,N_3436,N_3391);
and U3930 (N_3930,N_3341,N_3265);
nor U3931 (N_3931,N_3370,N_3104);
nor U3932 (N_3932,N_3319,N_3005);
nand U3933 (N_3933,N_3404,N_3177);
nor U3934 (N_3934,N_3145,N_3110);
or U3935 (N_3935,N_3377,N_3059);
nand U3936 (N_3936,N_3159,N_3369);
or U3937 (N_3937,N_3004,N_3259);
or U3938 (N_3938,N_3446,N_3215);
and U3939 (N_3939,N_3306,N_3236);
nand U3940 (N_3940,N_3220,N_3038);
nand U3941 (N_3941,N_3443,N_3257);
nand U3942 (N_3942,N_3352,N_3047);
nor U3943 (N_3943,N_3141,N_3072);
nand U3944 (N_3944,N_3362,N_3049);
nor U3945 (N_3945,N_3387,N_3400);
and U3946 (N_3946,N_3485,N_3437);
nor U3947 (N_3947,N_3323,N_3359);
or U3948 (N_3948,N_3459,N_3138);
and U3949 (N_3949,N_3164,N_3018);
or U3950 (N_3950,N_3030,N_3293);
and U3951 (N_3951,N_3197,N_3226);
nor U3952 (N_3952,N_3127,N_3488);
xor U3953 (N_3953,N_3391,N_3056);
nor U3954 (N_3954,N_3115,N_3177);
or U3955 (N_3955,N_3243,N_3205);
nand U3956 (N_3956,N_3225,N_3406);
and U3957 (N_3957,N_3480,N_3079);
and U3958 (N_3958,N_3312,N_3036);
and U3959 (N_3959,N_3066,N_3128);
and U3960 (N_3960,N_3299,N_3444);
nor U3961 (N_3961,N_3496,N_3404);
or U3962 (N_3962,N_3386,N_3031);
nand U3963 (N_3963,N_3068,N_3012);
xnor U3964 (N_3964,N_3000,N_3193);
nor U3965 (N_3965,N_3239,N_3308);
or U3966 (N_3966,N_3387,N_3131);
or U3967 (N_3967,N_3323,N_3246);
and U3968 (N_3968,N_3166,N_3081);
and U3969 (N_3969,N_3229,N_3259);
nor U3970 (N_3970,N_3435,N_3295);
or U3971 (N_3971,N_3221,N_3487);
and U3972 (N_3972,N_3393,N_3252);
and U3973 (N_3973,N_3377,N_3468);
or U3974 (N_3974,N_3466,N_3105);
or U3975 (N_3975,N_3049,N_3361);
nand U3976 (N_3976,N_3197,N_3438);
and U3977 (N_3977,N_3022,N_3132);
nor U3978 (N_3978,N_3475,N_3350);
nand U3979 (N_3979,N_3027,N_3241);
and U3980 (N_3980,N_3353,N_3385);
nand U3981 (N_3981,N_3210,N_3470);
or U3982 (N_3982,N_3215,N_3348);
and U3983 (N_3983,N_3268,N_3376);
or U3984 (N_3984,N_3260,N_3404);
or U3985 (N_3985,N_3250,N_3375);
nand U3986 (N_3986,N_3075,N_3163);
or U3987 (N_3987,N_3479,N_3247);
nand U3988 (N_3988,N_3227,N_3219);
or U3989 (N_3989,N_3214,N_3125);
nor U3990 (N_3990,N_3381,N_3297);
or U3991 (N_3991,N_3457,N_3497);
or U3992 (N_3992,N_3175,N_3373);
nand U3993 (N_3993,N_3423,N_3316);
nand U3994 (N_3994,N_3189,N_3320);
or U3995 (N_3995,N_3116,N_3008);
nor U3996 (N_3996,N_3124,N_3112);
or U3997 (N_3997,N_3419,N_3325);
nand U3998 (N_3998,N_3452,N_3096);
nand U3999 (N_3999,N_3015,N_3391);
nor U4000 (N_4000,N_3928,N_3919);
and U4001 (N_4001,N_3963,N_3829);
and U4002 (N_4002,N_3708,N_3825);
nor U4003 (N_4003,N_3715,N_3733);
or U4004 (N_4004,N_3538,N_3965);
nor U4005 (N_4005,N_3700,N_3754);
and U4006 (N_4006,N_3648,N_3529);
and U4007 (N_4007,N_3939,N_3736);
nand U4008 (N_4008,N_3576,N_3892);
nand U4009 (N_4009,N_3775,N_3956);
or U4010 (N_4010,N_3973,N_3575);
and U4011 (N_4011,N_3502,N_3916);
and U4012 (N_4012,N_3975,N_3568);
and U4013 (N_4013,N_3804,N_3637);
nor U4014 (N_4014,N_3604,N_3967);
nor U4015 (N_4015,N_3812,N_3561);
nor U4016 (N_4016,N_3912,N_3657);
nand U4017 (N_4017,N_3946,N_3696);
nor U4018 (N_4018,N_3757,N_3945);
nor U4019 (N_4019,N_3814,N_3875);
and U4020 (N_4020,N_3920,N_3776);
or U4021 (N_4021,N_3552,N_3583);
nor U4022 (N_4022,N_3587,N_3745);
or U4023 (N_4023,N_3861,N_3905);
nor U4024 (N_4024,N_3666,N_3799);
nand U4025 (N_4025,N_3541,N_3857);
and U4026 (N_4026,N_3750,N_3959);
and U4027 (N_4027,N_3629,N_3990);
or U4028 (N_4028,N_3887,N_3810);
or U4029 (N_4029,N_3501,N_3893);
or U4030 (N_4030,N_3542,N_3738);
nor U4031 (N_4031,N_3773,N_3867);
or U4032 (N_4032,N_3524,N_3739);
and U4033 (N_4033,N_3950,N_3760);
and U4034 (N_4034,N_3543,N_3915);
or U4035 (N_4035,N_3823,N_3589);
nor U4036 (N_4036,N_3876,N_3765);
nor U4037 (N_4037,N_3870,N_3922);
nand U4038 (N_4038,N_3544,N_3880);
or U4039 (N_4039,N_3599,N_3507);
nor U4040 (N_4040,N_3882,N_3838);
nand U4041 (N_4041,N_3707,N_3550);
nor U4042 (N_4042,N_3753,N_3966);
and U4043 (N_4043,N_3660,N_3714);
or U4044 (N_4044,N_3659,N_3646);
nor U4045 (N_4045,N_3603,N_3743);
and U4046 (N_4046,N_3772,N_3549);
or U4047 (N_4047,N_3682,N_3938);
nor U4048 (N_4048,N_3904,N_3996);
and U4049 (N_4049,N_3645,N_3651);
nor U4050 (N_4050,N_3551,N_3989);
and U4051 (N_4051,N_3594,N_3795);
or U4052 (N_4052,N_3830,N_3514);
nor U4053 (N_4053,N_3617,N_3855);
nor U4054 (N_4054,N_3994,N_3506);
nand U4055 (N_4055,N_3656,N_3807);
and U4056 (N_4056,N_3547,N_3968);
nand U4057 (N_4057,N_3711,N_3530);
nor U4058 (N_4058,N_3789,N_3598);
nand U4059 (N_4059,N_3802,N_3792);
or U4060 (N_4060,N_3947,N_3525);
and U4061 (N_4061,N_3592,N_3889);
nor U4062 (N_4062,N_3567,N_3737);
nand U4063 (N_4063,N_3621,N_3722);
nor U4064 (N_4064,N_3957,N_3664);
and U4065 (N_4065,N_3570,N_3716);
nand U4066 (N_4066,N_3566,N_3510);
nor U4067 (N_4067,N_3782,N_3741);
nand U4068 (N_4068,N_3793,N_3719);
or U4069 (N_4069,N_3951,N_3937);
and U4070 (N_4070,N_3559,N_3586);
nor U4071 (N_4071,N_3631,N_3731);
and U4072 (N_4072,N_3798,N_3844);
and U4073 (N_4073,N_3866,N_3974);
or U4074 (N_4074,N_3518,N_3761);
or U4075 (N_4075,N_3560,N_3608);
and U4076 (N_4076,N_3819,N_3863);
nor U4077 (N_4077,N_3602,N_3862);
or U4078 (N_4078,N_3623,N_3585);
nor U4079 (N_4079,N_3704,N_3613);
nor U4080 (N_4080,N_3686,N_3509);
nor U4081 (N_4081,N_3703,N_3545);
and U4082 (N_4082,N_3747,N_3847);
nand U4083 (N_4083,N_3824,N_3500);
nand U4084 (N_4084,N_3991,N_3987);
and U4085 (N_4085,N_3885,N_3512);
nand U4086 (N_4086,N_3769,N_3619);
nand U4087 (N_4087,N_3597,N_3624);
or U4088 (N_4088,N_3532,N_3834);
or U4089 (N_4089,N_3988,N_3781);
and U4090 (N_4090,N_3751,N_3816);
or U4091 (N_4091,N_3744,N_3699);
nand U4092 (N_4092,N_3924,N_3684);
or U4093 (N_4093,N_3535,N_3685);
or U4094 (N_4094,N_3851,N_3569);
nor U4095 (N_4095,N_3677,N_3969);
nand U4096 (N_4096,N_3976,N_3890);
nor U4097 (N_4097,N_3874,N_3788);
or U4098 (N_4098,N_3521,N_3644);
or U4099 (N_4099,N_3815,N_3516);
and U4100 (N_4100,N_3571,N_3641);
or U4101 (N_4101,N_3710,N_3591);
nor U4102 (N_4102,N_3752,N_3794);
nand U4103 (N_4103,N_3590,N_3609);
nor U4104 (N_4104,N_3717,N_3790);
xor U4105 (N_4105,N_3681,N_3981);
or U4106 (N_4106,N_3971,N_3910);
or U4107 (N_4107,N_3800,N_3626);
or U4108 (N_4108,N_3577,N_3859);
xnor U4109 (N_4109,N_3649,N_3999);
nand U4110 (N_4110,N_3955,N_3786);
nor U4111 (N_4111,N_3513,N_3895);
or U4112 (N_4112,N_3809,N_3709);
nand U4113 (N_4113,N_3735,N_3909);
nand U4114 (N_4114,N_3826,N_3632);
and U4115 (N_4115,N_3522,N_3746);
or U4116 (N_4116,N_3980,N_3907);
nand U4117 (N_4117,N_3993,N_3953);
or U4118 (N_4118,N_3891,N_3929);
and U4119 (N_4119,N_3588,N_3596);
or U4120 (N_4120,N_3740,N_3948);
nor U4121 (N_4121,N_3785,N_3877);
and U4122 (N_4122,N_3846,N_3574);
and U4123 (N_4123,N_3845,N_3690);
and U4124 (N_4124,N_3694,N_3523);
and U4125 (N_4125,N_3713,N_3764);
nor U4126 (N_4126,N_3534,N_3768);
and U4127 (N_4127,N_3848,N_3520);
and U4128 (N_4128,N_3943,N_3540);
nand U4129 (N_4129,N_3777,N_3858);
or U4130 (N_4130,N_3970,N_3625);
nand U4131 (N_4131,N_3808,N_3932);
nand U4132 (N_4132,N_3505,N_3771);
or U4133 (N_4133,N_3977,N_3732);
or U4134 (N_4134,N_3584,N_3936);
nand U4135 (N_4135,N_3986,N_3558);
nor U4136 (N_4136,N_3724,N_3705);
and U4137 (N_4137,N_3511,N_3820);
or U4138 (N_4138,N_3533,N_3688);
nand U4139 (N_4139,N_3811,N_3640);
nand U4140 (N_4140,N_3580,N_3837);
or U4141 (N_4141,N_3553,N_3852);
or U4142 (N_4142,N_3658,N_3872);
nand U4143 (N_4143,N_3849,N_3949);
nor U4144 (N_4144,N_3519,N_3600);
nand U4145 (N_4145,N_3721,N_3898);
or U4146 (N_4146,N_3868,N_3998);
and U4147 (N_4147,N_3620,N_3923);
nor U4148 (N_4148,N_3564,N_3888);
nand U4149 (N_4149,N_3821,N_3818);
nor U4150 (N_4150,N_3997,N_3758);
xnor U4151 (N_4151,N_3762,N_3712);
nand U4152 (N_4152,N_3903,N_3652);
and U4153 (N_4153,N_3663,N_3831);
or U4154 (N_4154,N_3979,N_3899);
nor U4155 (N_4155,N_3667,N_3610);
and U4156 (N_4156,N_3805,N_3636);
nand U4157 (N_4157,N_3729,N_3940);
nand U4158 (N_4158,N_3985,N_3983);
xor U4159 (N_4159,N_3557,N_3555);
and U4160 (N_4160,N_3601,N_3668);
nand U4161 (N_4161,N_3770,N_3536);
nand U4162 (N_4162,N_3896,N_3650);
nor U4163 (N_4163,N_3748,N_3774);
nor U4164 (N_4164,N_3528,N_3615);
or U4165 (N_4165,N_3680,N_3972);
nand U4166 (N_4166,N_3642,N_3960);
nand U4167 (N_4167,N_3833,N_3606);
nand U4168 (N_4168,N_3803,N_3653);
and U4169 (N_4169,N_3673,N_3579);
or U4170 (N_4170,N_3548,N_3595);
nor U4171 (N_4171,N_3839,N_3720);
and U4172 (N_4172,N_3678,N_3931);
nand U4173 (N_4173,N_3995,N_3779);
nand U4174 (N_4174,N_3886,N_3871);
nor U4175 (N_4175,N_3727,N_3883);
and U4176 (N_4176,N_3639,N_3628);
and U4177 (N_4177,N_3702,N_3730);
or U4178 (N_4178,N_3783,N_3661);
and U4179 (N_4179,N_3836,N_3921);
nand U4180 (N_4180,N_3692,N_3546);
nor U4181 (N_4181,N_3539,N_3901);
nor U4182 (N_4182,N_3873,N_3726);
and U4183 (N_4183,N_3878,N_3647);
or U4184 (N_4184,N_3618,N_3695);
or U4185 (N_4185,N_3913,N_3643);
and U4186 (N_4186,N_3954,N_3778);
or U4187 (N_4187,N_3655,N_3578);
nor U4188 (N_4188,N_3728,N_3835);
and U4189 (N_4189,N_3843,N_3962);
nand U4190 (N_4190,N_3822,N_3897);
nand U4191 (N_4191,N_3934,N_3515);
nand U4192 (N_4192,N_3562,N_3503);
nand U4193 (N_4193,N_3734,N_3864);
and U4194 (N_4194,N_3508,N_3723);
or U4195 (N_4195,N_3926,N_3622);
nand U4196 (N_4196,N_3672,N_3669);
and U4197 (N_4197,N_3787,N_3791);
nor U4198 (N_4198,N_3832,N_3554);
nand U4199 (N_4199,N_3676,N_3627);
or U4200 (N_4200,N_3638,N_3693);
nand U4201 (N_4201,N_3817,N_3842);
and U4202 (N_4202,N_3813,N_3698);
nor U4203 (N_4203,N_3869,N_3796);
nor U4204 (N_4204,N_3942,N_3573);
nor U4205 (N_4205,N_3616,N_3806);
nand U4206 (N_4206,N_3840,N_3927);
nor U4207 (N_4207,N_3581,N_3982);
nand U4208 (N_4208,N_3925,N_3634);
and U4209 (N_4209,N_3675,N_3749);
or U4210 (N_4210,N_3854,N_3630);
or U4211 (N_4211,N_3902,N_3827);
nor U4212 (N_4212,N_3766,N_3689);
nor U4213 (N_4213,N_3908,N_3917);
nor U4214 (N_4214,N_3881,N_3900);
or U4215 (N_4215,N_3884,N_3952);
nand U4216 (N_4216,N_3984,N_3701);
nand U4217 (N_4217,N_3992,N_3911);
or U4218 (N_4218,N_3879,N_3865);
or U4219 (N_4219,N_3918,N_3767);
and U4220 (N_4220,N_3718,N_3933);
or U4221 (N_4221,N_3556,N_3565);
and U4222 (N_4222,N_3687,N_3662);
or U4223 (N_4223,N_3611,N_3784);
nor U4224 (N_4224,N_3856,N_3801);
nand U4225 (N_4225,N_3853,N_3860);
and U4226 (N_4226,N_3572,N_3964);
and U4227 (N_4227,N_3961,N_3605);
nor U4228 (N_4228,N_3582,N_3612);
xor U4229 (N_4229,N_3633,N_3828);
or U4230 (N_4230,N_3614,N_3531);
nor U4231 (N_4231,N_3665,N_3756);
and U4232 (N_4232,N_3563,N_3697);
nor U4233 (N_4233,N_3941,N_3763);
nor U4234 (N_4234,N_3683,N_3725);
or U4235 (N_4235,N_3635,N_3593);
and U4236 (N_4236,N_3679,N_3670);
and U4237 (N_4237,N_3517,N_3654);
nor U4238 (N_4238,N_3935,N_3894);
nor U4239 (N_4239,N_3691,N_3755);
nand U4240 (N_4240,N_3527,N_3759);
or U4241 (N_4241,N_3674,N_3914);
nor U4242 (N_4242,N_3850,N_3607);
nand U4243 (N_4243,N_3526,N_3797);
nand U4244 (N_4244,N_3978,N_3944);
or U4245 (N_4245,N_3742,N_3906);
and U4246 (N_4246,N_3671,N_3780);
or U4247 (N_4247,N_3841,N_3706);
nand U4248 (N_4248,N_3537,N_3958);
nor U4249 (N_4249,N_3930,N_3504);
nor U4250 (N_4250,N_3749,N_3909);
nand U4251 (N_4251,N_3724,N_3925);
and U4252 (N_4252,N_3599,N_3701);
nor U4253 (N_4253,N_3884,N_3512);
nand U4254 (N_4254,N_3990,N_3620);
nor U4255 (N_4255,N_3697,N_3787);
nor U4256 (N_4256,N_3921,N_3893);
and U4257 (N_4257,N_3800,N_3510);
nand U4258 (N_4258,N_3766,N_3931);
and U4259 (N_4259,N_3636,N_3848);
nor U4260 (N_4260,N_3682,N_3917);
nand U4261 (N_4261,N_3709,N_3562);
or U4262 (N_4262,N_3923,N_3617);
nand U4263 (N_4263,N_3866,N_3677);
xor U4264 (N_4264,N_3589,N_3717);
or U4265 (N_4265,N_3717,N_3998);
nand U4266 (N_4266,N_3727,N_3714);
nand U4267 (N_4267,N_3660,N_3564);
nand U4268 (N_4268,N_3831,N_3879);
or U4269 (N_4269,N_3646,N_3591);
or U4270 (N_4270,N_3713,N_3837);
nor U4271 (N_4271,N_3861,N_3835);
nand U4272 (N_4272,N_3952,N_3737);
or U4273 (N_4273,N_3985,N_3896);
nand U4274 (N_4274,N_3987,N_3774);
nor U4275 (N_4275,N_3628,N_3863);
and U4276 (N_4276,N_3929,N_3681);
or U4277 (N_4277,N_3612,N_3964);
and U4278 (N_4278,N_3777,N_3678);
nand U4279 (N_4279,N_3502,N_3586);
nand U4280 (N_4280,N_3768,N_3502);
nand U4281 (N_4281,N_3866,N_3938);
or U4282 (N_4282,N_3759,N_3564);
nor U4283 (N_4283,N_3804,N_3893);
or U4284 (N_4284,N_3525,N_3721);
nor U4285 (N_4285,N_3698,N_3679);
and U4286 (N_4286,N_3753,N_3552);
nor U4287 (N_4287,N_3748,N_3756);
nand U4288 (N_4288,N_3574,N_3894);
nand U4289 (N_4289,N_3742,N_3504);
and U4290 (N_4290,N_3585,N_3599);
nor U4291 (N_4291,N_3925,N_3626);
nand U4292 (N_4292,N_3742,N_3610);
nand U4293 (N_4293,N_3883,N_3522);
or U4294 (N_4294,N_3590,N_3716);
and U4295 (N_4295,N_3900,N_3840);
nor U4296 (N_4296,N_3953,N_3585);
and U4297 (N_4297,N_3746,N_3741);
xor U4298 (N_4298,N_3622,N_3890);
nand U4299 (N_4299,N_3721,N_3599);
or U4300 (N_4300,N_3564,N_3547);
nor U4301 (N_4301,N_3505,N_3666);
nor U4302 (N_4302,N_3536,N_3946);
nor U4303 (N_4303,N_3638,N_3727);
nand U4304 (N_4304,N_3826,N_3691);
nand U4305 (N_4305,N_3825,N_3839);
nand U4306 (N_4306,N_3682,N_3968);
and U4307 (N_4307,N_3909,N_3819);
nand U4308 (N_4308,N_3791,N_3645);
and U4309 (N_4309,N_3861,N_3660);
nand U4310 (N_4310,N_3792,N_3678);
nor U4311 (N_4311,N_3975,N_3974);
or U4312 (N_4312,N_3954,N_3640);
nor U4313 (N_4313,N_3658,N_3672);
nor U4314 (N_4314,N_3666,N_3959);
or U4315 (N_4315,N_3830,N_3616);
and U4316 (N_4316,N_3926,N_3859);
or U4317 (N_4317,N_3616,N_3949);
nand U4318 (N_4318,N_3817,N_3705);
nand U4319 (N_4319,N_3650,N_3522);
and U4320 (N_4320,N_3518,N_3746);
and U4321 (N_4321,N_3876,N_3664);
nor U4322 (N_4322,N_3927,N_3670);
nor U4323 (N_4323,N_3513,N_3589);
nand U4324 (N_4324,N_3604,N_3953);
or U4325 (N_4325,N_3753,N_3914);
and U4326 (N_4326,N_3906,N_3669);
nor U4327 (N_4327,N_3795,N_3534);
or U4328 (N_4328,N_3693,N_3553);
and U4329 (N_4329,N_3754,N_3532);
or U4330 (N_4330,N_3897,N_3606);
and U4331 (N_4331,N_3509,N_3734);
nor U4332 (N_4332,N_3528,N_3857);
nand U4333 (N_4333,N_3951,N_3765);
nand U4334 (N_4334,N_3883,N_3834);
or U4335 (N_4335,N_3725,N_3990);
and U4336 (N_4336,N_3859,N_3667);
and U4337 (N_4337,N_3553,N_3596);
or U4338 (N_4338,N_3542,N_3968);
nor U4339 (N_4339,N_3591,N_3901);
nor U4340 (N_4340,N_3838,N_3942);
nand U4341 (N_4341,N_3636,N_3645);
nor U4342 (N_4342,N_3745,N_3827);
or U4343 (N_4343,N_3550,N_3938);
or U4344 (N_4344,N_3861,N_3531);
nor U4345 (N_4345,N_3629,N_3789);
or U4346 (N_4346,N_3854,N_3829);
nand U4347 (N_4347,N_3774,N_3690);
xnor U4348 (N_4348,N_3918,N_3764);
or U4349 (N_4349,N_3631,N_3824);
or U4350 (N_4350,N_3560,N_3754);
nor U4351 (N_4351,N_3843,N_3939);
and U4352 (N_4352,N_3896,N_3990);
nor U4353 (N_4353,N_3882,N_3962);
nand U4354 (N_4354,N_3696,N_3587);
or U4355 (N_4355,N_3990,N_3885);
nor U4356 (N_4356,N_3642,N_3715);
nand U4357 (N_4357,N_3712,N_3660);
and U4358 (N_4358,N_3877,N_3591);
and U4359 (N_4359,N_3708,N_3814);
and U4360 (N_4360,N_3722,N_3940);
nand U4361 (N_4361,N_3640,N_3848);
nand U4362 (N_4362,N_3898,N_3606);
xnor U4363 (N_4363,N_3682,N_3764);
or U4364 (N_4364,N_3584,N_3575);
nand U4365 (N_4365,N_3585,N_3629);
nor U4366 (N_4366,N_3900,N_3860);
nand U4367 (N_4367,N_3924,N_3737);
nor U4368 (N_4368,N_3507,N_3538);
nor U4369 (N_4369,N_3570,N_3537);
nor U4370 (N_4370,N_3897,N_3927);
nand U4371 (N_4371,N_3967,N_3526);
nor U4372 (N_4372,N_3904,N_3573);
and U4373 (N_4373,N_3692,N_3570);
nor U4374 (N_4374,N_3860,N_3992);
and U4375 (N_4375,N_3880,N_3885);
or U4376 (N_4376,N_3784,N_3841);
and U4377 (N_4377,N_3912,N_3941);
and U4378 (N_4378,N_3701,N_3817);
nor U4379 (N_4379,N_3813,N_3581);
or U4380 (N_4380,N_3723,N_3877);
nor U4381 (N_4381,N_3565,N_3988);
and U4382 (N_4382,N_3984,N_3741);
nor U4383 (N_4383,N_3934,N_3848);
and U4384 (N_4384,N_3941,N_3767);
nand U4385 (N_4385,N_3678,N_3837);
and U4386 (N_4386,N_3916,N_3823);
or U4387 (N_4387,N_3905,N_3526);
nor U4388 (N_4388,N_3819,N_3851);
and U4389 (N_4389,N_3722,N_3958);
or U4390 (N_4390,N_3795,N_3549);
nand U4391 (N_4391,N_3643,N_3958);
nand U4392 (N_4392,N_3804,N_3761);
or U4393 (N_4393,N_3877,N_3886);
and U4394 (N_4394,N_3658,N_3601);
and U4395 (N_4395,N_3712,N_3996);
nand U4396 (N_4396,N_3806,N_3847);
and U4397 (N_4397,N_3621,N_3983);
nor U4398 (N_4398,N_3932,N_3627);
xor U4399 (N_4399,N_3617,N_3651);
and U4400 (N_4400,N_3917,N_3757);
or U4401 (N_4401,N_3968,N_3954);
nor U4402 (N_4402,N_3722,N_3556);
nand U4403 (N_4403,N_3537,N_3596);
or U4404 (N_4404,N_3701,N_3648);
or U4405 (N_4405,N_3938,N_3948);
and U4406 (N_4406,N_3730,N_3810);
or U4407 (N_4407,N_3720,N_3569);
and U4408 (N_4408,N_3929,N_3598);
nand U4409 (N_4409,N_3797,N_3904);
nor U4410 (N_4410,N_3951,N_3794);
nor U4411 (N_4411,N_3703,N_3951);
nor U4412 (N_4412,N_3910,N_3624);
or U4413 (N_4413,N_3510,N_3671);
and U4414 (N_4414,N_3600,N_3835);
nand U4415 (N_4415,N_3780,N_3758);
or U4416 (N_4416,N_3508,N_3951);
nor U4417 (N_4417,N_3711,N_3790);
or U4418 (N_4418,N_3981,N_3992);
or U4419 (N_4419,N_3815,N_3979);
nand U4420 (N_4420,N_3609,N_3575);
or U4421 (N_4421,N_3857,N_3925);
and U4422 (N_4422,N_3640,N_3675);
and U4423 (N_4423,N_3962,N_3776);
xnor U4424 (N_4424,N_3747,N_3692);
xor U4425 (N_4425,N_3900,N_3876);
nor U4426 (N_4426,N_3735,N_3663);
and U4427 (N_4427,N_3627,N_3897);
or U4428 (N_4428,N_3914,N_3946);
nor U4429 (N_4429,N_3998,N_3945);
xor U4430 (N_4430,N_3985,N_3945);
nor U4431 (N_4431,N_3557,N_3967);
xor U4432 (N_4432,N_3517,N_3777);
nand U4433 (N_4433,N_3584,N_3797);
nand U4434 (N_4434,N_3691,N_3612);
xnor U4435 (N_4435,N_3623,N_3928);
nand U4436 (N_4436,N_3940,N_3559);
nor U4437 (N_4437,N_3818,N_3938);
and U4438 (N_4438,N_3894,N_3938);
nand U4439 (N_4439,N_3704,N_3598);
or U4440 (N_4440,N_3833,N_3924);
nor U4441 (N_4441,N_3712,N_3944);
or U4442 (N_4442,N_3986,N_3970);
nand U4443 (N_4443,N_3924,N_3523);
and U4444 (N_4444,N_3988,N_3522);
and U4445 (N_4445,N_3999,N_3978);
nand U4446 (N_4446,N_3746,N_3701);
nand U4447 (N_4447,N_3652,N_3622);
nor U4448 (N_4448,N_3814,N_3730);
nand U4449 (N_4449,N_3706,N_3617);
and U4450 (N_4450,N_3598,N_3938);
nor U4451 (N_4451,N_3828,N_3809);
or U4452 (N_4452,N_3963,N_3714);
nor U4453 (N_4453,N_3665,N_3543);
nand U4454 (N_4454,N_3758,N_3982);
nand U4455 (N_4455,N_3538,N_3562);
and U4456 (N_4456,N_3722,N_3545);
nand U4457 (N_4457,N_3695,N_3764);
nor U4458 (N_4458,N_3837,N_3795);
and U4459 (N_4459,N_3797,N_3821);
nor U4460 (N_4460,N_3821,N_3640);
nor U4461 (N_4461,N_3564,N_3510);
or U4462 (N_4462,N_3538,N_3870);
nand U4463 (N_4463,N_3631,N_3774);
nand U4464 (N_4464,N_3504,N_3882);
or U4465 (N_4465,N_3804,N_3611);
or U4466 (N_4466,N_3860,N_3901);
and U4467 (N_4467,N_3896,N_3727);
or U4468 (N_4468,N_3609,N_3576);
or U4469 (N_4469,N_3688,N_3729);
or U4470 (N_4470,N_3950,N_3784);
or U4471 (N_4471,N_3587,N_3607);
or U4472 (N_4472,N_3778,N_3634);
and U4473 (N_4473,N_3650,N_3681);
and U4474 (N_4474,N_3836,N_3850);
or U4475 (N_4475,N_3522,N_3936);
or U4476 (N_4476,N_3518,N_3693);
nand U4477 (N_4477,N_3599,N_3516);
and U4478 (N_4478,N_3894,N_3540);
or U4479 (N_4479,N_3812,N_3906);
or U4480 (N_4480,N_3569,N_3622);
nor U4481 (N_4481,N_3970,N_3745);
or U4482 (N_4482,N_3775,N_3900);
and U4483 (N_4483,N_3772,N_3689);
nand U4484 (N_4484,N_3632,N_3870);
nor U4485 (N_4485,N_3951,N_3696);
nand U4486 (N_4486,N_3693,N_3596);
nor U4487 (N_4487,N_3823,N_3704);
or U4488 (N_4488,N_3871,N_3976);
and U4489 (N_4489,N_3816,N_3996);
nor U4490 (N_4490,N_3907,N_3589);
or U4491 (N_4491,N_3685,N_3620);
or U4492 (N_4492,N_3853,N_3835);
and U4493 (N_4493,N_3541,N_3540);
and U4494 (N_4494,N_3920,N_3698);
nand U4495 (N_4495,N_3821,N_3993);
and U4496 (N_4496,N_3897,N_3758);
nor U4497 (N_4497,N_3895,N_3651);
nor U4498 (N_4498,N_3568,N_3967);
and U4499 (N_4499,N_3778,N_3765);
and U4500 (N_4500,N_4067,N_4314);
nand U4501 (N_4501,N_4123,N_4162);
and U4502 (N_4502,N_4049,N_4471);
and U4503 (N_4503,N_4389,N_4379);
or U4504 (N_4504,N_4220,N_4409);
and U4505 (N_4505,N_4167,N_4369);
nor U4506 (N_4506,N_4420,N_4018);
nand U4507 (N_4507,N_4350,N_4164);
nor U4508 (N_4508,N_4107,N_4181);
or U4509 (N_4509,N_4457,N_4290);
nand U4510 (N_4510,N_4322,N_4077);
or U4511 (N_4511,N_4238,N_4171);
and U4512 (N_4512,N_4448,N_4361);
or U4513 (N_4513,N_4211,N_4044);
nand U4514 (N_4514,N_4278,N_4437);
nand U4515 (N_4515,N_4345,N_4154);
nand U4516 (N_4516,N_4255,N_4310);
nand U4517 (N_4517,N_4245,N_4493);
or U4518 (N_4518,N_4026,N_4359);
and U4519 (N_4519,N_4432,N_4249);
nor U4520 (N_4520,N_4479,N_4396);
or U4521 (N_4521,N_4126,N_4333);
nand U4522 (N_4522,N_4398,N_4120);
and U4523 (N_4523,N_4439,N_4159);
and U4524 (N_4524,N_4449,N_4052);
nand U4525 (N_4525,N_4299,N_4486);
and U4526 (N_4526,N_4055,N_4365);
nor U4527 (N_4527,N_4225,N_4112);
nor U4528 (N_4528,N_4308,N_4109);
nor U4529 (N_4529,N_4069,N_4202);
or U4530 (N_4530,N_4336,N_4467);
nand U4531 (N_4531,N_4499,N_4276);
nor U4532 (N_4532,N_4408,N_4246);
nor U4533 (N_4533,N_4149,N_4402);
and U4534 (N_4534,N_4051,N_4233);
and U4535 (N_4535,N_4101,N_4095);
or U4536 (N_4536,N_4039,N_4301);
or U4537 (N_4537,N_4262,N_4076);
and U4538 (N_4538,N_4491,N_4070);
and U4539 (N_4539,N_4043,N_4175);
nand U4540 (N_4540,N_4495,N_4334);
and U4541 (N_4541,N_4496,N_4190);
nand U4542 (N_4542,N_4300,N_4413);
nor U4543 (N_4543,N_4306,N_4232);
nand U4544 (N_4544,N_4279,N_4475);
and U4545 (N_4545,N_4141,N_4231);
nor U4546 (N_4546,N_4033,N_4074);
or U4547 (N_4547,N_4468,N_4323);
nand U4548 (N_4548,N_4316,N_4234);
nand U4549 (N_4549,N_4169,N_4286);
nand U4550 (N_4550,N_4161,N_4013);
nand U4551 (N_4551,N_4341,N_4046);
or U4552 (N_4552,N_4196,N_4452);
nand U4553 (N_4553,N_4269,N_4206);
or U4554 (N_4554,N_4360,N_4006);
and U4555 (N_4555,N_4143,N_4157);
nand U4556 (N_4556,N_4089,N_4405);
or U4557 (N_4557,N_4252,N_4460);
or U4558 (N_4558,N_4216,N_4108);
or U4559 (N_4559,N_4002,N_4118);
nor U4560 (N_4560,N_4168,N_4153);
or U4561 (N_4561,N_4094,N_4199);
and U4562 (N_4562,N_4366,N_4304);
and U4563 (N_4563,N_4391,N_4250);
and U4564 (N_4564,N_4145,N_4098);
nor U4565 (N_4565,N_4031,N_4434);
and U4566 (N_4566,N_4288,N_4458);
xnor U4567 (N_4567,N_4138,N_4223);
or U4568 (N_4568,N_4047,N_4326);
or U4569 (N_4569,N_4435,N_4390);
nand U4570 (N_4570,N_4189,N_4239);
nor U4571 (N_4571,N_4148,N_4351);
or U4572 (N_4572,N_4445,N_4251);
and U4573 (N_4573,N_4374,N_4419);
and U4574 (N_4574,N_4227,N_4003);
xnor U4575 (N_4575,N_4022,N_4183);
nor U4576 (N_4576,N_4103,N_4414);
and U4577 (N_4577,N_4447,N_4021);
or U4578 (N_4578,N_4335,N_4444);
nor U4579 (N_4579,N_4195,N_4241);
nand U4580 (N_4580,N_4462,N_4182);
or U4581 (N_4581,N_4348,N_4340);
or U4582 (N_4582,N_4338,N_4384);
and U4583 (N_4583,N_4265,N_4289);
nor U4584 (N_4584,N_4174,N_4260);
nor U4585 (N_4585,N_4240,N_4053);
and U4586 (N_4586,N_4235,N_4205);
or U4587 (N_4587,N_4424,N_4242);
or U4588 (N_4588,N_4372,N_4226);
nand U4589 (N_4589,N_4010,N_4482);
or U4590 (N_4590,N_4463,N_4000);
or U4591 (N_4591,N_4059,N_4364);
nand U4592 (N_4592,N_4179,N_4459);
nand U4593 (N_4593,N_4056,N_4040);
and U4594 (N_4594,N_4090,N_4100);
or U4595 (N_4595,N_4378,N_4110);
nand U4596 (N_4596,N_4099,N_4441);
nor U4597 (N_4597,N_4208,N_4011);
nand U4598 (N_4598,N_4236,N_4380);
and U4599 (N_4599,N_4488,N_4277);
or U4600 (N_4600,N_4080,N_4453);
nand U4601 (N_4601,N_4209,N_4283);
nor U4602 (N_4602,N_4025,N_4492);
nor U4603 (N_4603,N_4088,N_4274);
and U4604 (N_4604,N_4065,N_4433);
and U4605 (N_4605,N_4058,N_4229);
and U4606 (N_4606,N_4106,N_4176);
nand U4607 (N_4607,N_4117,N_4387);
nand U4608 (N_4608,N_4014,N_4184);
and U4609 (N_4609,N_4173,N_4004);
xor U4610 (N_4610,N_4130,N_4258);
nand U4611 (N_4611,N_4045,N_4124);
and U4612 (N_4612,N_4337,N_4429);
nand U4613 (N_4613,N_4219,N_4343);
and U4614 (N_4614,N_4354,N_4440);
or U4615 (N_4615,N_4375,N_4266);
and U4616 (N_4616,N_4007,N_4166);
nor U4617 (N_4617,N_4151,N_4020);
and U4618 (N_4618,N_4192,N_4297);
or U4619 (N_4619,N_4037,N_4019);
nor U4620 (N_4620,N_4293,N_4131);
and U4621 (N_4621,N_4093,N_4393);
or U4622 (N_4622,N_4105,N_4431);
nand U4623 (N_4623,N_4030,N_4498);
or U4624 (N_4624,N_4084,N_4358);
nor U4625 (N_4625,N_4066,N_4230);
nor U4626 (N_4626,N_4178,N_4349);
xnor U4627 (N_4627,N_4281,N_4024);
and U4628 (N_4628,N_4477,N_4042);
nand U4629 (N_4629,N_4275,N_4023);
nor U4630 (N_4630,N_4451,N_4285);
nand U4631 (N_4631,N_4152,N_4292);
nand U4632 (N_4632,N_4214,N_4356);
and U4633 (N_4633,N_4330,N_4446);
nand U4634 (N_4634,N_4305,N_4060);
xor U4635 (N_4635,N_4091,N_4422);
or U4636 (N_4636,N_4092,N_4368);
nor U4637 (N_4637,N_4137,N_4228);
or U4638 (N_4638,N_4421,N_4165);
nand U4639 (N_4639,N_4261,N_4050);
or U4640 (N_4640,N_4127,N_4303);
nand U4641 (N_4641,N_4357,N_4362);
nor U4642 (N_4642,N_4332,N_4038);
nor U4643 (N_4643,N_4036,N_4344);
or U4644 (N_4644,N_4342,N_4201);
nand U4645 (N_4645,N_4325,N_4385);
and U4646 (N_4646,N_4296,N_4312);
nand U4647 (N_4647,N_4193,N_4071);
nand U4648 (N_4648,N_4140,N_4207);
nand U4649 (N_4649,N_4407,N_4456);
or U4650 (N_4650,N_4347,N_4073);
or U4651 (N_4651,N_4324,N_4478);
nor U4652 (N_4652,N_4480,N_4061);
and U4653 (N_4653,N_4180,N_4489);
nor U4654 (N_4654,N_4054,N_4476);
or U4655 (N_4655,N_4156,N_4454);
nand U4656 (N_4656,N_4257,N_4243);
nand U4657 (N_4657,N_4404,N_4147);
nor U4658 (N_4658,N_4353,N_4273);
xnor U4659 (N_4659,N_4144,N_4016);
nand U4660 (N_4660,N_4346,N_4470);
and U4661 (N_4661,N_4086,N_4210);
or U4662 (N_4662,N_4102,N_4472);
and U4663 (N_4663,N_4097,N_4425);
or U4664 (N_4664,N_4150,N_4383);
or U4665 (N_4665,N_4373,N_4427);
or U4666 (N_4666,N_4442,N_4072);
nor U4667 (N_4667,N_4415,N_4485);
or U4668 (N_4668,N_4484,N_4388);
and U4669 (N_4669,N_4078,N_4139);
nand U4670 (N_4670,N_4291,N_4008);
or U4671 (N_4671,N_4009,N_4186);
nand U4672 (N_4672,N_4410,N_4247);
nand U4673 (N_4673,N_4001,N_4158);
nand U4674 (N_4674,N_4381,N_4237);
xor U4675 (N_4675,N_4370,N_4280);
and U4676 (N_4676,N_4027,N_4386);
nand U4677 (N_4677,N_4075,N_4048);
and U4678 (N_4678,N_4400,N_4494);
or U4679 (N_4679,N_4327,N_4417);
or U4680 (N_4680,N_4426,N_4155);
nor U4681 (N_4681,N_4443,N_4177);
or U4682 (N_4682,N_4244,N_4412);
and U4683 (N_4683,N_4087,N_4487);
or U4684 (N_4684,N_4318,N_4270);
nand U4685 (N_4685,N_4259,N_4397);
or U4686 (N_4686,N_4298,N_4194);
nor U4687 (N_4687,N_4085,N_4132);
nor U4688 (N_4688,N_4116,N_4197);
nor U4689 (N_4689,N_4371,N_4403);
nand U4690 (N_4690,N_4012,N_4215);
nand U4691 (N_4691,N_4253,N_4317);
and U4692 (N_4692,N_4015,N_4473);
and U4693 (N_4693,N_4315,N_4198);
nor U4694 (N_4694,N_4135,N_4163);
and U4695 (N_4695,N_4321,N_4302);
nor U4696 (N_4696,N_4081,N_4465);
nor U4697 (N_4697,N_4068,N_4083);
and U4698 (N_4698,N_4319,N_4328);
or U4699 (N_4699,N_4224,N_4146);
or U4700 (N_4700,N_4264,N_4170);
nand U4701 (N_4701,N_4490,N_4474);
or U4702 (N_4702,N_4111,N_4461);
nand U4703 (N_4703,N_4469,N_4200);
nand U4704 (N_4704,N_4436,N_4455);
nor U4705 (N_4705,N_4256,N_4423);
nor U4706 (N_4706,N_4204,N_4160);
nor U4707 (N_4707,N_4191,N_4221);
nor U4708 (N_4708,N_4079,N_4272);
or U4709 (N_4709,N_4411,N_4268);
nor U4710 (N_4710,N_4395,N_4082);
and U4711 (N_4711,N_4294,N_4497);
or U4712 (N_4712,N_4284,N_4129);
nand U4713 (N_4713,N_4331,N_4394);
nor U4714 (N_4714,N_4464,N_4483);
nor U4715 (N_4715,N_4134,N_4028);
or U4716 (N_4716,N_4254,N_4263);
or U4717 (N_4717,N_4136,N_4035);
nand U4718 (N_4718,N_4032,N_4438);
nor U4719 (N_4719,N_4119,N_4034);
or U4720 (N_4720,N_4248,N_4466);
nor U4721 (N_4721,N_4172,N_4185);
or U4722 (N_4722,N_4339,N_4271);
and U4723 (N_4723,N_4295,N_4311);
and U4724 (N_4724,N_4104,N_4188);
nand U4725 (N_4725,N_4005,N_4222);
and U4726 (N_4726,N_4367,N_4313);
or U4727 (N_4727,N_4213,N_4217);
and U4728 (N_4728,N_4376,N_4218);
and U4729 (N_4729,N_4041,N_4212);
nand U4730 (N_4730,N_4064,N_4063);
nand U4731 (N_4731,N_4377,N_4096);
or U4732 (N_4732,N_4017,N_4287);
nand U4733 (N_4733,N_4428,N_4309);
or U4734 (N_4734,N_4416,N_4307);
and U4735 (N_4735,N_4481,N_4392);
or U4736 (N_4736,N_4057,N_4113);
nand U4737 (N_4737,N_4128,N_4121);
or U4738 (N_4738,N_4320,N_4114);
nand U4739 (N_4739,N_4399,N_4203);
and U4740 (N_4740,N_4355,N_4401);
xor U4741 (N_4741,N_4406,N_4430);
nand U4742 (N_4742,N_4329,N_4122);
nor U4743 (N_4743,N_4382,N_4363);
or U4744 (N_4744,N_4142,N_4418);
and U4745 (N_4745,N_4133,N_4282);
nand U4746 (N_4746,N_4187,N_4352);
or U4747 (N_4747,N_4267,N_4125);
nor U4748 (N_4748,N_4062,N_4029);
or U4749 (N_4749,N_4115,N_4450);
xnor U4750 (N_4750,N_4237,N_4172);
or U4751 (N_4751,N_4462,N_4372);
nand U4752 (N_4752,N_4325,N_4073);
nand U4753 (N_4753,N_4073,N_4445);
or U4754 (N_4754,N_4008,N_4259);
nand U4755 (N_4755,N_4239,N_4300);
nor U4756 (N_4756,N_4406,N_4133);
or U4757 (N_4757,N_4332,N_4196);
nand U4758 (N_4758,N_4239,N_4213);
nor U4759 (N_4759,N_4242,N_4155);
and U4760 (N_4760,N_4265,N_4361);
nand U4761 (N_4761,N_4461,N_4473);
and U4762 (N_4762,N_4089,N_4252);
and U4763 (N_4763,N_4076,N_4431);
nor U4764 (N_4764,N_4160,N_4486);
xnor U4765 (N_4765,N_4101,N_4311);
nand U4766 (N_4766,N_4403,N_4119);
and U4767 (N_4767,N_4301,N_4375);
nand U4768 (N_4768,N_4163,N_4197);
or U4769 (N_4769,N_4303,N_4186);
or U4770 (N_4770,N_4128,N_4066);
nor U4771 (N_4771,N_4323,N_4067);
and U4772 (N_4772,N_4423,N_4006);
nand U4773 (N_4773,N_4294,N_4336);
nor U4774 (N_4774,N_4490,N_4124);
and U4775 (N_4775,N_4499,N_4145);
and U4776 (N_4776,N_4273,N_4276);
nand U4777 (N_4777,N_4006,N_4144);
nor U4778 (N_4778,N_4399,N_4298);
and U4779 (N_4779,N_4007,N_4056);
nor U4780 (N_4780,N_4185,N_4405);
nor U4781 (N_4781,N_4451,N_4358);
and U4782 (N_4782,N_4184,N_4239);
nor U4783 (N_4783,N_4062,N_4134);
nor U4784 (N_4784,N_4274,N_4334);
and U4785 (N_4785,N_4126,N_4072);
xnor U4786 (N_4786,N_4496,N_4090);
and U4787 (N_4787,N_4221,N_4443);
and U4788 (N_4788,N_4176,N_4205);
nand U4789 (N_4789,N_4331,N_4371);
or U4790 (N_4790,N_4429,N_4467);
nor U4791 (N_4791,N_4159,N_4161);
nand U4792 (N_4792,N_4400,N_4405);
nand U4793 (N_4793,N_4056,N_4084);
nand U4794 (N_4794,N_4115,N_4424);
nor U4795 (N_4795,N_4375,N_4229);
and U4796 (N_4796,N_4498,N_4044);
xor U4797 (N_4797,N_4038,N_4475);
and U4798 (N_4798,N_4090,N_4299);
and U4799 (N_4799,N_4431,N_4445);
or U4800 (N_4800,N_4476,N_4308);
nand U4801 (N_4801,N_4217,N_4096);
nand U4802 (N_4802,N_4041,N_4498);
nor U4803 (N_4803,N_4479,N_4047);
and U4804 (N_4804,N_4333,N_4388);
or U4805 (N_4805,N_4262,N_4422);
and U4806 (N_4806,N_4316,N_4151);
nand U4807 (N_4807,N_4224,N_4290);
and U4808 (N_4808,N_4028,N_4327);
or U4809 (N_4809,N_4118,N_4390);
nand U4810 (N_4810,N_4266,N_4059);
xnor U4811 (N_4811,N_4104,N_4371);
nand U4812 (N_4812,N_4348,N_4041);
and U4813 (N_4813,N_4301,N_4198);
nor U4814 (N_4814,N_4131,N_4111);
or U4815 (N_4815,N_4082,N_4135);
or U4816 (N_4816,N_4459,N_4121);
nand U4817 (N_4817,N_4001,N_4379);
and U4818 (N_4818,N_4238,N_4073);
nand U4819 (N_4819,N_4056,N_4265);
or U4820 (N_4820,N_4023,N_4293);
or U4821 (N_4821,N_4405,N_4309);
or U4822 (N_4822,N_4448,N_4189);
nand U4823 (N_4823,N_4025,N_4483);
and U4824 (N_4824,N_4097,N_4487);
nand U4825 (N_4825,N_4334,N_4228);
nor U4826 (N_4826,N_4277,N_4131);
nand U4827 (N_4827,N_4226,N_4141);
nor U4828 (N_4828,N_4057,N_4027);
nor U4829 (N_4829,N_4284,N_4388);
or U4830 (N_4830,N_4388,N_4189);
and U4831 (N_4831,N_4423,N_4417);
or U4832 (N_4832,N_4087,N_4036);
or U4833 (N_4833,N_4478,N_4430);
nand U4834 (N_4834,N_4359,N_4056);
nand U4835 (N_4835,N_4482,N_4475);
and U4836 (N_4836,N_4006,N_4129);
nand U4837 (N_4837,N_4002,N_4209);
or U4838 (N_4838,N_4274,N_4260);
nand U4839 (N_4839,N_4111,N_4291);
nor U4840 (N_4840,N_4096,N_4017);
or U4841 (N_4841,N_4365,N_4067);
nand U4842 (N_4842,N_4063,N_4174);
and U4843 (N_4843,N_4007,N_4494);
nor U4844 (N_4844,N_4211,N_4098);
and U4845 (N_4845,N_4365,N_4092);
nor U4846 (N_4846,N_4473,N_4421);
and U4847 (N_4847,N_4205,N_4381);
and U4848 (N_4848,N_4488,N_4493);
nand U4849 (N_4849,N_4058,N_4468);
or U4850 (N_4850,N_4087,N_4134);
nand U4851 (N_4851,N_4121,N_4388);
or U4852 (N_4852,N_4284,N_4401);
xnor U4853 (N_4853,N_4275,N_4378);
nand U4854 (N_4854,N_4155,N_4278);
nor U4855 (N_4855,N_4066,N_4494);
nor U4856 (N_4856,N_4162,N_4279);
or U4857 (N_4857,N_4182,N_4381);
nand U4858 (N_4858,N_4268,N_4392);
nand U4859 (N_4859,N_4294,N_4423);
nand U4860 (N_4860,N_4209,N_4109);
or U4861 (N_4861,N_4385,N_4044);
or U4862 (N_4862,N_4469,N_4063);
and U4863 (N_4863,N_4304,N_4127);
or U4864 (N_4864,N_4499,N_4074);
or U4865 (N_4865,N_4033,N_4216);
nor U4866 (N_4866,N_4234,N_4286);
nand U4867 (N_4867,N_4010,N_4393);
nor U4868 (N_4868,N_4355,N_4264);
or U4869 (N_4869,N_4226,N_4376);
nand U4870 (N_4870,N_4463,N_4227);
nand U4871 (N_4871,N_4448,N_4348);
nand U4872 (N_4872,N_4277,N_4168);
or U4873 (N_4873,N_4401,N_4178);
nor U4874 (N_4874,N_4075,N_4270);
nand U4875 (N_4875,N_4132,N_4350);
and U4876 (N_4876,N_4472,N_4202);
and U4877 (N_4877,N_4338,N_4003);
nor U4878 (N_4878,N_4302,N_4289);
and U4879 (N_4879,N_4333,N_4361);
nand U4880 (N_4880,N_4250,N_4111);
and U4881 (N_4881,N_4364,N_4445);
and U4882 (N_4882,N_4207,N_4238);
and U4883 (N_4883,N_4127,N_4087);
xor U4884 (N_4884,N_4232,N_4340);
nor U4885 (N_4885,N_4016,N_4356);
and U4886 (N_4886,N_4001,N_4245);
and U4887 (N_4887,N_4001,N_4372);
or U4888 (N_4888,N_4381,N_4494);
nand U4889 (N_4889,N_4346,N_4268);
and U4890 (N_4890,N_4356,N_4196);
or U4891 (N_4891,N_4079,N_4238);
or U4892 (N_4892,N_4114,N_4145);
nand U4893 (N_4893,N_4205,N_4370);
and U4894 (N_4894,N_4117,N_4259);
nor U4895 (N_4895,N_4449,N_4464);
and U4896 (N_4896,N_4379,N_4362);
nand U4897 (N_4897,N_4415,N_4406);
and U4898 (N_4898,N_4147,N_4463);
and U4899 (N_4899,N_4057,N_4269);
nor U4900 (N_4900,N_4499,N_4130);
nand U4901 (N_4901,N_4277,N_4442);
nand U4902 (N_4902,N_4412,N_4141);
or U4903 (N_4903,N_4202,N_4262);
nor U4904 (N_4904,N_4046,N_4235);
nor U4905 (N_4905,N_4452,N_4154);
nor U4906 (N_4906,N_4188,N_4306);
or U4907 (N_4907,N_4006,N_4150);
nor U4908 (N_4908,N_4363,N_4233);
or U4909 (N_4909,N_4405,N_4109);
and U4910 (N_4910,N_4289,N_4095);
or U4911 (N_4911,N_4071,N_4140);
nand U4912 (N_4912,N_4010,N_4218);
nand U4913 (N_4913,N_4072,N_4474);
nand U4914 (N_4914,N_4272,N_4146);
nor U4915 (N_4915,N_4187,N_4018);
nand U4916 (N_4916,N_4376,N_4309);
or U4917 (N_4917,N_4272,N_4477);
and U4918 (N_4918,N_4386,N_4438);
nand U4919 (N_4919,N_4242,N_4246);
and U4920 (N_4920,N_4215,N_4205);
nor U4921 (N_4921,N_4438,N_4156);
nand U4922 (N_4922,N_4346,N_4190);
or U4923 (N_4923,N_4091,N_4311);
nor U4924 (N_4924,N_4191,N_4286);
xnor U4925 (N_4925,N_4131,N_4326);
nand U4926 (N_4926,N_4483,N_4282);
nand U4927 (N_4927,N_4256,N_4414);
or U4928 (N_4928,N_4314,N_4099);
and U4929 (N_4929,N_4142,N_4303);
nor U4930 (N_4930,N_4454,N_4309);
nand U4931 (N_4931,N_4318,N_4351);
nor U4932 (N_4932,N_4442,N_4021);
and U4933 (N_4933,N_4129,N_4091);
nor U4934 (N_4934,N_4425,N_4207);
nor U4935 (N_4935,N_4483,N_4085);
nand U4936 (N_4936,N_4110,N_4306);
nand U4937 (N_4937,N_4456,N_4169);
and U4938 (N_4938,N_4105,N_4497);
or U4939 (N_4939,N_4059,N_4344);
nor U4940 (N_4940,N_4371,N_4006);
nor U4941 (N_4941,N_4109,N_4284);
nor U4942 (N_4942,N_4458,N_4016);
or U4943 (N_4943,N_4458,N_4100);
or U4944 (N_4944,N_4285,N_4496);
nand U4945 (N_4945,N_4229,N_4351);
nor U4946 (N_4946,N_4032,N_4315);
and U4947 (N_4947,N_4146,N_4023);
nor U4948 (N_4948,N_4407,N_4165);
nand U4949 (N_4949,N_4010,N_4428);
and U4950 (N_4950,N_4361,N_4150);
and U4951 (N_4951,N_4098,N_4183);
nand U4952 (N_4952,N_4297,N_4287);
or U4953 (N_4953,N_4021,N_4296);
nor U4954 (N_4954,N_4308,N_4446);
nor U4955 (N_4955,N_4202,N_4481);
nor U4956 (N_4956,N_4414,N_4059);
and U4957 (N_4957,N_4301,N_4022);
or U4958 (N_4958,N_4258,N_4460);
nor U4959 (N_4959,N_4260,N_4342);
nand U4960 (N_4960,N_4183,N_4069);
and U4961 (N_4961,N_4248,N_4310);
nor U4962 (N_4962,N_4013,N_4290);
xnor U4963 (N_4963,N_4395,N_4318);
or U4964 (N_4964,N_4440,N_4297);
nand U4965 (N_4965,N_4020,N_4317);
and U4966 (N_4966,N_4162,N_4494);
and U4967 (N_4967,N_4081,N_4417);
nand U4968 (N_4968,N_4476,N_4113);
or U4969 (N_4969,N_4037,N_4454);
nand U4970 (N_4970,N_4458,N_4419);
and U4971 (N_4971,N_4359,N_4060);
or U4972 (N_4972,N_4354,N_4495);
nand U4973 (N_4973,N_4052,N_4315);
nand U4974 (N_4974,N_4471,N_4234);
nand U4975 (N_4975,N_4144,N_4413);
and U4976 (N_4976,N_4200,N_4321);
or U4977 (N_4977,N_4076,N_4486);
nand U4978 (N_4978,N_4104,N_4083);
nor U4979 (N_4979,N_4107,N_4447);
nand U4980 (N_4980,N_4394,N_4476);
and U4981 (N_4981,N_4092,N_4475);
or U4982 (N_4982,N_4405,N_4356);
and U4983 (N_4983,N_4398,N_4210);
xnor U4984 (N_4984,N_4117,N_4019);
or U4985 (N_4985,N_4362,N_4271);
nor U4986 (N_4986,N_4289,N_4022);
nand U4987 (N_4987,N_4160,N_4338);
nor U4988 (N_4988,N_4214,N_4407);
or U4989 (N_4989,N_4334,N_4265);
and U4990 (N_4990,N_4354,N_4333);
xor U4991 (N_4991,N_4334,N_4052);
nor U4992 (N_4992,N_4207,N_4438);
nand U4993 (N_4993,N_4416,N_4215);
and U4994 (N_4994,N_4363,N_4490);
or U4995 (N_4995,N_4346,N_4015);
nor U4996 (N_4996,N_4365,N_4289);
and U4997 (N_4997,N_4327,N_4191);
nor U4998 (N_4998,N_4376,N_4034);
or U4999 (N_4999,N_4103,N_4056);
nor U5000 (N_5000,N_4696,N_4515);
nor U5001 (N_5001,N_4504,N_4763);
and U5002 (N_5002,N_4660,N_4945);
nor U5003 (N_5003,N_4645,N_4699);
or U5004 (N_5004,N_4835,N_4631);
or U5005 (N_5005,N_4843,N_4852);
nand U5006 (N_5006,N_4726,N_4767);
or U5007 (N_5007,N_4548,N_4685);
or U5008 (N_5008,N_4971,N_4926);
and U5009 (N_5009,N_4589,N_4951);
or U5010 (N_5010,N_4974,N_4879);
nor U5011 (N_5011,N_4571,N_4680);
nand U5012 (N_5012,N_4790,N_4523);
and U5013 (N_5013,N_4700,N_4941);
and U5014 (N_5014,N_4781,N_4987);
nor U5015 (N_5015,N_4908,N_4590);
or U5016 (N_5016,N_4716,N_4510);
or U5017 (N_5017,N_4818,N_4834);
and U5018 (N_5018,N_4770,N_4925);
nand U5019 (N_5019,N_4568,N_4842);
nand U5020 (N_5020,N_4506,N_4780);
nand U5021 (N_5021,N_4869,N_4562);
or U5022 (N_5022,N_4965,N_4611);
or U5023 (N_5023,N_4621,N_4964);
nand U5024 (N_5024,N_4988,N_4825);
nor U5025 (N_5025,N_4844,N_4764);
xnor U5026 (N_5026,N_4886,N_4737);
or U5027 (N_5027,N_4727,N_4858);
nand U5028 (N_5028,N_4778,N_4855);
nand U5029 (N_5029,N_4602,N_4677);
nor U5030 (N_5030,N_4918,N_4877);
or U5031 (N_5031,N_4829,N_4900);
or U5032 (N_5032,N_4675,N_4931);
and U5033 (N_5033,N_4681,N_4977);
and U5034 (N_5034,N_4513,N_4968);
or U5035 (N_5035,N_4898,N_4782);
and U5036 (N_5036,N_4522,N_4657);
and U5037 (N_5037,N_4676,N_4709);
or U5038 (N_5038,N_4610,N_4910);
or U5039 (N_5039,N_4623,N_4638);
nand U5040 (N_5040,N_4758,N_4644);
or U5041 (N_5041,N_4874,N_4996);
and U5042 (N_5042,N_4715,N_4574);
or U5043 (N_5043,N_4972,N_4804);
or U5044 (N_5044,N_4706,N_4719);
nand U5045 (N_5045,N_4628,N_4554);
and U5046 (N_5046,N_4615,N_4919);
and U5047 (N_5047,N_4836,N_4881);
nand U5048 (N_5048,N_4591,N_4538);
nor U5049 (N_5049,N_4608,N_4739);
nand U5050 (N_5050,N_4788,N_4952);
nor U5051 (N_5051,N_4928,N_4997);
and U5052 (N_5052,N_4800,N_4730);
or U5053 (N_5053,N_4728,N_4777);
or U5054 (N_5054,N_4774,N_4870);
or U5055 (N_5055,N_4885,N_4557);
or U5056 (N_5056,N_4786,N_4771);
or U5057 (N_5057,N_4775,N_4752);
nor U5058 (N_5058,N_4533,N_4979);
nor U5059 (N_5059,N_4731,N_4599);
or U5060 (N_5060,N_4514,N_4766);
and U5061 (N_5061,N_4937,N_4656);
and U5062 (N_5062,N_4635,N_4756);
nand U5063 (N_5063,N_4995,N_4856);
nand U5064 (N_5064,N_4601,N_4892);
nand U5065 (N_5065,N_4668,N_4641);
nand U5066 (N_5066,N_4605,N_4932);
and U5067 (N_5067,N_4787,N_4720);
nand U5068 (N_5068,N_4809,N_4849);
and U5069 (N_5069,N_4576,N_4950);
nor U5070 (N_5070,N_4582,N_4793);
nand U5071 (N_5071,N_4887,N_4954);
nor U5072 (N_5072,N_4876,N_4978);
nor U5073 (N_5073,N_4803,N_4519);
nor U5074 (N_5074,N_4906,N_4873);
and U5075 (N_5075,N_4986,N_4524);
nor U5076 (N_5076,N_4526,N_4822);
nand U5077 (N_5077,N_4587,N_4913);
or U5078 (N_5078,N_4646,N_4905);
nand U5079 (N_5079,N_4872,N_4802);
nor U5080 (N_5080,N_4903,N_4902);
nand U5081 (N_5081,N_4880,N_4757);
xor U5082 (N_5082,N_4542,N_4878);
and U5083 (N_5083,N_4652,N_4883);
and U5084 (N_5084,N_4831,N_4649);
and U5085 (N_5085,N_4759,N_4785);
nor U5086 (N_5086,N_4851,N_4684);
or U5087 (N_5087,N_4866,N_4961);
nor U5088 (N_5088,N_4629,N_4664);
or U5089 (N_5089,N_4654,N_4536);
nor U5090 (N_5090,N_4808,N_4982);
nor U5091 (N_5091,N_4584,N_4546);
or U5092 (N_5092,N_4854,N_4585);
or U5093 (N_5093,N_4695,N_4679);
nand U5094 (N_5094,N_4724,N_4946);
and U5095 (N_5095,N_4867,N_4537);
nand U5096 (N_5096,N_4606,N_4560);
nand U5097 (N_5097,N_4748,N_4967);
nor U5098 (N_5098,N_4772,N_4690);
or U5099 (N_5099,N_4922,N_4938);
nand U5100 (N_5100,N_4899,N_4505);
and U5101 (N_5101,N_4960,N_4865);
nor U5102 (N_5102,N_4799,N_4991);
nor U5103 (N_5103,N_4823,N_4632);
nand U5104 (N_5104,N_4847,N_4697);
nand U5105 (N_5105,N_4612,N_4503);
nor U5106 (N_5106,N_4934,N_4682);
nor U5107 (N_5107,N_4939,N_4705);
xnor U5108 (N_5108,N_4816,N_4776);
and U5109 (N_5109,N_4512,N_4710);
or U5110 (N_5110,N_4714,N_4572);
or U5111 (N_5111,N_4597,N_4529);
nor U5112 (N_5112,N_4738,N_4916);
nand U5113 (N_5113,N_4846,N_4807);
nand U5114 (N_5114,N_4920,N_4663);
or U5115 (N_5115,N_4559,N_4501);
and U5116 (N_5116,N_4973,N_4815);
and U5117 (N_5117,N_4666,N_4604);
or U5118 (N_5118,N_4754,N_4525);
and U5119 (N_5119,N_4915,N_4651);
or U5120 (N_5120,N_4897,N_4953);
nor U5121 (N_5121,N_4586,N_4662);
and U5122 (N_5122,N_4511,N_4875);
nand U5123 (N_5123,N_4600,N_4643);
and U5124 (N_5124,N_4634,N_4784);
and U5125 (N_5125,N_4698,N_4745);
nor U5126 (N_5126,N_4711,N_4821);
nor U5127 (N_5127,N_4575,N_4762);
or U5128 (N_5128,N_4647,N_4732);
nor U5129 (N_5129,N_4859,N_4544);
xor U5130 (N_5130,N_4796,N_4532);
nand U5131 (N_5131,N_4864,N_4595);
nand U5132 (N_5132,N_4528,N_4773);
or U5133 (N_5133,N_4890,N_4607);
and U5134 (N_5134,N_4751,N_4956);
and U5135 (N_5135,N_4653,N_4725);
and U5136 (N_5136,N_4923,N_4564);
and U5137 (N_5137,N_4545,N_4580);
or U5138 (N_5138,N_4627,N_4755);
nor U5139 (N_5139,N_4596,N_4520);
nor U5140 (N_5140,N_4556,N_4948);
nor U5141 (N_5141,N_4588,N_4712);
or U5142 (N_5142,N_4674,N_4517);
nand U5143 (N_5143,N_4530,N_4555);
and U5144 (N_5144,N_4686,N_4567);
nand U5145 (N_5145,N_4673,N_4783);
nand U5146 (N_5146,N_4630,N_4508);
or U5147 (N_5147,N_4765,N_4534);
or U5148 (N_5148,N_4990,N_4744);
nand U5149 (N_5149,N_4718,N_4687);
and U5150 (N_5150,N_4841,N_4701);
nand U5151 (N_5151,N_4994,N_4891);
nand U5152 (N_5152,N_4551,N_4579);
nand U5153 (N_5153,N_4549,N_4691);
or U5154 (N_5154,N_4717,N_4955);
nor U5155 (N_5155,N_4792,N_4861);
and U5156 (N_5156,N_4659,N_4863);
or U5157 (N_5157,N_4820,N_4985);
nor U5158 (N_5158,N_4502,N_4789);
nor U5159 (N_5159,N_4940,N_4936);
and U5160 (N_5160,N_4614,N_4998);
and U5161 (N_5161,N_4813,N_4578);
and U5162 (N_5162,N_4669,N_4637);
or U5163 (N_5163,N_4569,N_4707);
nand U5164 (N_5164,N_4500,N_4561);
nand U5165 (N_5165,N_4736,N_4570);
or U5166 (N_5166,N_4794,N_4671);
and U5167 (N_5167,N_4531,N_4661);
or U5168 (N_5168,N_4619,N_4640);
nor U5169 (N_5169,N_4577,N_4642);
nand U5170 (N_5170,N_4975,N_4907);
or U5171 (N_5171,N_4694,N_4672);
xnor U5172 (N_5172,N_4708,N_4558);
and U5173 (N_5173,N_4729,N_4678);
and U5174 (N_5174,N_4581,N_4895);
or U5175 (N_5175,N_4565,N_4983);
nand U5176 (N_5176,N_4911,N_4670);
or U5177 (N_5177,N_4924,N_4535);
and U5178 (N_5178,N_4942,N_4742);
nor U5179 (N_5179,N_4550,N_4617);
nand U5180 (N_5180,N_4958,N_4826);
and U5181 (N_5181,N_4845,N_4929);
nand U5182 (N_5182,N_4650,N_4658);
nor U5183 (N_5183,N_4655,N_4868);
and U5184 (N_5184,N_4566,N_4507);
nor U5185 (N_5185,N_4857,N_4624);
nand U5186 (N_5186,N_4840,N_4966);
xnor U5187 (N_5187,N_4917,N_4957);
or U5188 (N_5188,N_4594,N_4592);
or U5189 (N_5189,N_4693,N_4805);
or U5190 (N_5190,N_4980,N_4959);
or U5191 (N_5191,N_4944,N_4768);
nor U5192 (N_5192,N_4746,N_4509);
and U5193 (N_5193,N_4648,N_4893);
xnor U5194 (N_5194,N_4692,N_4824);
and U5195 (N_5195,N_4779,N_4633);
nand U5196 (N_5196,N_4688,N_4904);
or U5197 (N_5197,N_4993,N_4984);
and U5198 (N_5198,N_4833,N_4769);
nor U5199 (N_5199,N_4598,N_4909);
nor U5200 (N_5200,N_4828,N_4795);
or U5201 (N_5201,N_4989,N_4616);
and U5202 (N_5202,N_4702,N_4518);
nor U5203 (N_5203,N_4884,N_4713);
and U5204 (N_5204,N_4539,N_4827);
nand U5205 (N_5205,N_4626,N_4830);
nand U5206 (N_5206,N_4921,N_4552);
and U5207 (N_5207,N_4860,N_4583);
nand U5208 (N_5208,N_4721,N_4521);
nor U5209 (N_5209,N_4761,N_4889);
nand U5210 (N_5210,N_4733,N_4618);
nor U5211 (N_5211,N_4970,N_4806);
nand U5212 (N_5212,N_4896,N_4667);
or U5213 (N_5213,N_4563,N_4862);
nand U5214 (N_5214,N_4947,N_4704);
and U5215 (N_5215,N_4935,N_4992);
and U5216 (N_5216,N_4740,N_4969);
nand U5217 (N_5217,N_4837,N_4810);
or U5218 (N_5218,N_4943,N_4703);
or U5219 (N_5219,N_4553,N_4625);
xor U5220 (N_5220,N_4871,N_4593);
and U5221 (N_5221,N_4609,N_4817);
and U5222 (N_5222,N_4613,N_4540);
nor U5223 (N_5223,N_4927,N_4620);
or U5224 (N_5224,N_4798,N_4722);
or U5225 (N_5225,N_4622,N_4749);
and U5226 (N_5226,N_4527,N_4838);
nor U5227 (N_5227,N_4850,N_4930);
nand U5228 (N_5228,N_4812,N_4735);
and U5229 (N_5229,N_4914,N_4848);
and U5230 (N_5230,N_4797,N_4734);
xor U5231 (N_5231,N_4636,N_4888);
nor U5232 (N_5232,N_4603,N_4839);
nor U5233 (N_5233,N_4723,N_4747);
or U5234 (N_5234,N_4573,N_4543);
and U5235 (N_5235,N_4901,N_4811);
nand U5236 (N_5236,N_4981,N_4963);
nor U5237 (N_5237,N_4853,N_4976);
nand U5238 (N_5238,N_4832,N_4882);
and U5239 (N_5239,N_4516,N_4665);
nor U5240 (N_5240,N_4814,N_4801);
xnor U5241 (N_5241,N_4962,N_4894);
and U5242 (N_5242,N_4912,N_4933);
and U5243 (N_5243,N_4949,N_4819);
nor U5244 (N_5244,N_4760,N_4689);
nor U5245 (N_5245,N_4541,N_4741);
or U5246 (N_5246,N_4547,N_4683);
nor U5247 (N_5247,N_4753,N_4639);
or U5248 (N_5248,N_4791,N_4999);
nand U5249 (N_5249,N_4750,N_4743);
nand U5250 (N_5250,N_4880,N_4993);
and U5251 (N_5251,N_4637,N_4581);
nor U5252 (N_5252,N_4930,N_4774);
nor U5253 (N_5253,N_4522,N_4718);
nor U5254 (N_5254,N_4838,N_4600);
and U5255 (N_5255,N_4664,N_4984);
nor U5256 (N_5256,N_4819,N_4638);
nor U5257 (N_5257,N_4773,N_4971);
nor U5258 (N_5258,N_4602,N_4733);
nor U5259 (N_5259,N_4913,N_4616);
or U5260 (N_5260,N_4850,N_4991);
and U5261 (N_5261,N_4833,N_4788);
nand U5262 (N_5262,N_4993,N_4861);
nand U5263 (N_5263,N_4645,N_4636);
nor U5264 (N_5264,N_4633,N_4836);
nand U5265 (N_5265,N_4765,N_4523);
xnor U5266 (N_5266,N_4525,N_4510);
or U5267 (N_5267,N_4556,N_4544);
and U5268 (N_5268,N_4978,N_4579);
nor U5269 (N_5269,N_4717,N_4523);
or U5270 (N_5270,N_4867,N_4732);
or U5271 (N_5271,N_4717,N_4677);
nand U5272 (N_5272,N_4796,N_4530);
nor U5273 (N_5273,N_4704,N_4677);
or U5274 (N_5274,N_4957,N_4524);
or U5275 (N_5275,N_4791,N_4508);
nor U5276 (N_5276,N_4827,N_4990);
and U5277 (N_5277,N_4856,N_4645);
and U5278 (N_5278,N_4642,N_4835);
nor U5279 (N_5279,N_4651,N_4886);
xnor U5280 (N_5280,N_4577,N_4597);
and U5281 (N_5281,N_4613,N_4522);
nand U5282 (N_5282,N_4628,N_4539);
or U5283 (N_5283,N_4799,N_4854);
and U5284 (N_5284,N_4615,N_4854);
nand U5285 (N_5285,N_4795,N_4732);
nor U5286 (N_5286,N_4815,N_4972);
nor U5287 (N_5287,N_4656,N_4731);
nor U5288 (N_5288,N_4585,N_4887);
and U5289 (N_5289,N_4796,N_4916);
xnor U5290 (N_5290,N_4721,N_4559);
and U5291 (N_5291,N_4515,N_4526);
or U5292 (N_5292,N_4500,N_4999);
or U5293 (N_5293,N_4763,N_4637);
or U5294 (N_5294,N_4738,N_4936);
or U5295 (N_5295,N_4964,N_4581);
or U5296 (N_5296,N_4863,N_4646);
nor U5297 (N_5297,N_4959,N_4797);
and U5298 (N_5298,N_4855,N_4848);
nor U5299 (N_5299,N_4628,N_4704);
nand U5300 (N_5300,N_4710,N_4969);
nor U5301 (N_5301,N_4833,N_4749);
nor U5302 (N_5302,N_4917,N_4904);
or U5303 (N_5303,N_4619,N_4727);
nand U5304 (N_5304,N_4630,N_4955);
or U5305 (N_5305,N_4542,N_4728);
and U5306 (N_5306,N_4797,N_4617);
or U5307 (N_5307,N_4926,N_4585);
or U5308 (N_5308,N_4828,N_4953);
nor U5309 (N_5309,N_4604,N_4513);
nand U5310 (N_5310,N_4735,N_4620);
nand U5311 (N_5311,N_4514,N_4914);
or U5312 (N_5312,N_4793,N_4692);
or U5313 (N_5313,N_4693,N_4626);
nand U5314 (N_5314,N_4532,N_4934);
and U5315 (N_5315,N_4825,N_4894);
and U5316 (N_5316,N_4503,N_4946);
and U5317 (N_5317,N_4646,N_4781);
nand U5318 (N_5318,N_4911,N_4500);
nor U5319 (N_5319,N_4833,N_4837);
or U5320 (N_5320,N_4596,N_4957);
and U5321 (N_5321,N_4611,N_4806);
and U5322 (N_5322,N_4932,N_4907);
xnor U5323 (N_5323,N_4609,N_4851);
or U5324 (N_5324,N_4967,N_4584);
nor U5325 (N_5325,N_4801,N_4632);
and U5326 (N_5326,N_4872,N_4692);
nor U5327 (N_5327,N_4980,N_4798);
and U5328 (N_5328,N_4682,N_4610);
nand U5329 (N_5329,N_4733,N_4783);
and U5330 (N_5330,N_4535,N_4550);
or U5331 (N_5331,N_4604,N_4576);
or U5332 (N_5332,N_4642,N_4592);
nor U5333 (N_5333,N_4891,N_4698);
nand U5334 (N_5334,N_4916,N_4736);
nand U5335 (N_5335,N_4881,N_4655);
nand U5336 (N_5336,N_4858,N_4588);
and U5337 (N_5337,N_4901,N_4684);
and U5338 (N_5338,N_4609,N_4647);
and U5339 (N_5339,N_4952,N_4665);
and U5340 (N_5340,N_4639,N_4979);
and U5341 (N_5341,N_4945,N_4593);
nor U5342 (N_5342,N_4836,N_4842);
nand U5343 (N_5343,N_4763,N_4715);
or U5344 (N_5344,N_4502,N_4656);
and U5345 (N_5345,N_4858,N_4685);
or U5346 (N_5346,N_4760,N_4868);
and U5347 (N_5347,N_4530,N_4923);
and U5348 (N_5348,N_4871,N_4942);
and U5349 (N_5349,N_4904,N_4961);
nand U5350 (N_5350,N_4531,N_4569);
nor U5351 (N_5351,N_4849,N_4868);
and U5352 (N_5352,N_4866,N_4971);
nor U5353 (N_5353,N_4977,N_4511);
nand U5354 (N_5354,N_4561,N_4799);
and U5355 (N_5355,N_4731,N_4910);
or U5356 (N_5356,N_4527,N_4849);
nand U5357 (N_5357,N_4980,N_4552);
nor U5358 (N_5358,N_4945,N_4773);
nor U5359 (N_5359,N_4525,N_4514);
and U5360 (N_5360,N_4504,N_4883);
or U5361 (N_5361,N_4560,N_4787);
and U5362 (N_5362,N_4924,N_4657);
or U5363 (N_5363,N_4676,N_4664);
nor U5364 (N_5364,N_4944,N_4709);
nand U5365 (N_5365,N_4697,N_4513);
nand U5366 (N_5366,N_4603,N_4617);
nor U5367 (N_5367,N_4965,N_4586);
nor U5368 (N_5368,N_4665,N_4806);
or U5369 (N_5369,N_4923,N_4541);
or U5370 (N_5370,N_4676,N_4503);
nor U5371 (N_5371,N_4580,N_4625);
xor U5372 (N_5372,N_4967,N_4536);
or U5373 (N_5373,N_4509,N_4988);
nand U5374 (N_5374,N_4903,N_4828);
nand U5375 (N_5375,N_4645,N_4820);
nor U5376 (N_5376,N_4666,N_4691);
or U5377 (N_5377,N_4502,N_4713);
and U5378 (N_5378,N_4828,N_4911);
nor U5379 (N_5379,N_4718,N_4701);
and U5380 (N_5380,N_4813,N_4538);
nand U5381 (N_5381,N_4605,N_4963);
and U5382 (N_5382,N_4816,N_4714);
or U5383 (N_5383,N_4890,N_4990);
nand U5384 (N_5384,N_4832,N_4740);
nand U5385 (N_5385,N_4805,N_4868);
nor U5386 (N_5386,N_4860,N_4984);
or U5387 (N_5387,N_4784,N_4550);
nor U5388 (N_5388,N_4665,N_4595);
and U5389 (N_5389,N_4749,N_4898);
nand U5390 (N_5390,N_4951,N_4945);
or U5391 (N_5391,N_4693,N_4622);
nor U5392 (N_5392,N_4966,N_4825);
and U5393 (N_5393,N_4976,N_4720);
and U5394 (N_5394,N_4529,N_4516);
or U5395 (N_5395,N_4961,N_4667);
nand U5396 (N_5396,N_4792,N_4555);
and U5397 (N_5397,N_4776,N_4881);
or U5398 (N_5398,N_4547,N_4834);
or U5399 (N_5399,N_4679,N_4842);
nand U5400 (N_5400,N_4925,N_4816);
or U5401 (N_5401,N_4858,N_4676);
or U5402 (N_5402,N_4960,N_4916);
nor U5403 (N_5403,N_4825,N_4957);
and U5404 (N_5404,N_4822,N_4884);
or U5405 (N_5405,N_4844,N_4699);
nand U5406 (N_5406,N_4989,N_4966);
nor U5407 (N_5407,N_4767,N_4559);
nor U5408 (N_5408,N_4684,N_4862);
and U5409 (N_5409,N_4529,N_4719);
nor U5410 (N_5410,N_4559,N_4993);
nand U5411 (N_5411,N_4537,N_4926);
nor U5412 (N_5412,N_4913,N_4599);
nor U5413 (N_5413,N_4614,N_4504);
nor U5414 (N_5414,N_4929,N_4745);
xor U5415 (N_5415,N_4651,N_4669);
nor U5416 (N_5416,N_4676,N_4584);
nand U5417 (N_5417,N_4733,N_4511);
nand U5418 (N_5418,N_4655,N_4893);
and U5419 (N_5419,N_4861,N_4939);
and U5420 (N_5420,N_4551,N_4744);
nor U5421 (N_5421,N_4651,N_4905);
nand U5422 (N_5422,N_4509,N_4578);
nand U5423 (N_5423,N_4782,N_4730);
or U5424 (N_5424,N_4637,N_4562);
or U5425 (N_5425,N_4597,N_4820);
or U5426 (N_5426,N_4594,N_4739);
or U5427 (N_5427,N_4572,N_4783);
nand U5428 (N_5428,N_4502,N_4582);
nor U5429 (N_5429,N_4964,N_4996);
nor U5430 (N_5430,N_4525,N_4650);
nand U5431 (N_5431,N_4517,N_4892);
nand U5432 (N_5432,N_4684,N_4741);
nand U5433 (N_5433,N_4818,N_4696);
nor U5434 (N_5434,N_4885,N_4975);
nand U5435 (N_5435,N_4733,N_4610);
and U5436 (N_5436,N_4940,N_4610);
nor U5437 (N_5437,N_4804,N_4701);
nand U5438 (N_5438,N_4852,N_4601);
nor U5439 (N_5439,N_4776,N_4718);
and U5440 (N_5440,N_4754,N_4659);
and U5441 (N_5441,N_4603,N_4622);
nand U5442 (N_5442,N_4663,N_4743);
and U5443 (N_5443,N_4543,N_4959);
nor U5444 (N_5444,N_4757,N_4742);
and U5445 (N_5445,N_4829,N_4984);
nor U5446 (N_5446,N_4871,N_4865);
or U5447 (N_5447,N_4628,N_4808);
and U5448 (N_5448,N_4693,N_4802);
nor U5449 (N_5449,N_4964,N_4747);
and U5450 (N_5450,N_4775,N_4774);
or U5451 (N_5451,N_4771,N_4795);
or U5452 (N_5452,N_4749,N_4760);
nand U5453 (N_5453,N_4542,N_4889);
nor U5454 (N_5454,N_4540,N_4608);
xor U5455 (N_5455,N_4518,N_4690);
xor U5456 (N_5456,N_4792,N_4573);
nand U5457 (N_5457,N_4819,N_4683);
nor U5458 (N_5458,N_4967,N_4616);
nand U5459 (N_5459,N_4967,N_4657);
and U5460 (N_5460,N_4804,N_4846);
nor U5461 (N_5461,N_4564,N_4902);
nor U5462 (N_5462,N_4936,N_4865);
nand U5463 (N_5463,N_4981,N_4695);
and U5464 (N_5464,N_4758,N_4905);
nand U5465 (N_5465,N_4618,N_4622);
nor U5466 (N_5466,N_4843,N_4614);
nand U5467 (N_5467,N_4574,N_4551);
nor U5468 (N_5468,N_4650,N_4863);
or U5469 (N_5469,N_4765,N_4855);
nor U5470 (N_5470,N_4834,N_4832);
and U5471 (N_5471,N_4665,N_4898);
and U5472 (N_5472,N_4577,N_4855);
or U5473 (N_5473,N_4980,N_4740);
nor U5474 (N_5474,N_4670,N_4647);
nor U5475 (N_5475,N_4910,N_4558);
or U5476 (N_5476,N_4603,N_4914);
nand U5477 (N_5477,N_4805,N_4743);
nor U5478 (N_5478,N_4844,N_4599);
nand U5479 (N_5479,N_4934,N_4529);
nand U5480 (N_5480,N_4832,N_4826);
and U5481 (N_5481,N_4684,N_4559);
and U5482 (N_5482,N_4968,N_4824);
or U5483 (N_5483,N_4555,N_4727);
nor U5484 (N_5484,N_4803,N_4848);
nor U5485 (N_5485,N_4781,N_4841);
nand U5486 (N_5486,N_4550,N_4804);
nor U5487 (N_5487,N_4862,N_4926);
and U5488 (N_5488,N_4880,N_4552);
nand U5489 (N_5489,N_4655,N_4533);
and U5490 (N_5490,N_4783,N_4649);
nand U5491 (N_5491,N_4924,N_4512);
or U5492 (N_5492,N_4529,N_4605);
or U5493 (N_5493,N_4625,N_4952);
or U5494 (N_5494,N_4649,N_4788);
nand U5495 (N_5495,N_4885,N_4787);
and U5496 (N_5496,N_4989,N_4514);
and U5497 (N_5497,N_4689,N_4583);
nand U5498 (N_5498,N_4824,N_4623);
and U5499 (N_5499,N_4780,N_4750);
and U5500 (N_5500,N_5448,N_5327);
or U5501 (N_5501,N_5308,N_5183);
or U5502 (N_5502,N_5140,N_5335);
nor U5503 (N_5503,N_5251,N_5270);
and U5504 (N_5504,N_5344,N_5460);
nor U5505 (N_5505,N_5422,N_5434);
nand U5506 (N_5506,N_5386,N_5336);
nand U5507 (N_5507,N_5090,N_5383);
and U5508 (N_5508,N_5264,N_5026);
nand U5509 (N_5509,N_5033,N_5174);
nor U5510 (N_5510,N_5019,N_5471);
and U5511 (N_5511,N_5040,N_5388);
xor U5512 (N_5512,N_5363,N_5346);
and U5513 (N_5513,N_5061,N_5461);
nand U5514 (N_5514,N_5146,N_5405);
nand U5515 (N_5515,N_5170,N_5199);
nand U5516 (N_5516,N_5177,N_5182);
or U5517 (N_5517,N_5116,N_5057);
and U5518 (N_5518,N_5331,N_5167);
or U5519 (N_5519,N_5168,N_5348);
and U5520 (N_5520,N_5258,N_5157);
and U5521 (N_5521,N_5216,N_5124);
nor U5522 (N_5522,N_5400,N_5016);
or U5523 (N_5523,N_5161,N_5268);
nor U5524 (N_5524,N_5240,N_5282);
nor U5525 (N_5525,N_5111,N_5317);
xor U5526 (N_5526,N_5088,N_5401);
nand U5527 (N_5527,N_5103,N_5328);
and U5528 (N_5528,N_5145,N_5228);
and U5529 (N_5529,N_5466,N_5347);
or U5530 (N_5530,N_5244,N_5229);
and U5531 (N_5531,N_5274,N_5430);
or U5532 (N_5532,N_5000,N_5462);
and U5533 (N_5533,N_5293,N_5425);
or U5534 (N_5534,N_5214,N_5393);
xnor U5535 (N_5535,N_5360,N_5475);
or U5536 (N_5536,N_5075,N_5138);
or U5537 (N_5537,N_5028,N_5342);
or U5538 (N_5538,N_5097,N_5069);
nand U5539 (N_5539,N_5054,N_5439);
nand U5540 (N_5540,N_5421,N_5024);
nand U5541 (N_5541,N_5303,N_5417);
nor U5542 (N_5542,N_5094,N_5076);
nand U5543 (N_5543,N_5206,N_5458);
or U5544 (N_5544,N_5192,N_5144);
nor U5545 (N_5545,N_5212,N_5065);
and U5546 (N_5546,N_5048,N_5162);
or U5547 (N_5547,N_5198,N_5323);
nand U5548 (N_5548,N_5385,N_5106);
nor U5549 (N_5549,N_5012,N_5232);
nor U5550 (N_5550,N_5296,N_5053);
nor U5551 (N_5551,N_5397,N_5160);
or U5552 (N_5552,N_5486,N_5318);
nand U5553 (N_5553,N_5482,N_5469);
and U5554 (N_5554,N_5432,N_5487);
nand U5555 (N_5555,N_5431,N_5255);
or U5556 (N_5556,N_5427,N_5123);
nor U5557 (N_5557,N_5298,N_5250);
nand U5558 (N_5558,N_5237,N_5132);
or U5559 (N_5559,N_5442,N_5497);
nor U5560 (N_5560,N_5139,N_5239);
nor U5561 (N_5561,N_5299,N_5280);
or U5562 (N_5562,N_5234,N_5267);
nand U5563 (N_5563,N_5351,N_5355);
or U5564 (N_5564,N_5172,N_5188);
or U5565 (N_5565,N_5226,N_5257);
nand U5566 (N_5566,N_5339,N_5005);
or U5567 (N_5567,N_5474,N_5155);
or U5568 (N_5568,N_5231,N_5023);
and U5569 (N_5569,N_5450,N_5078);
or U5570 (N_5570,N_5100,N_5201);
and U5571 (N_5571,N_5429,N_5027);
nor U5572 (N_5572,N_5071,N_5008);
nor U5573 (N_5573,N_5083,N_5072);
nor U5574 (N_5574,N_5131,N_5241);
nand U5575 (N_5575,N_5227,N_5371);
nor U5576 (N_5576,N_5128,N_5249);
or U5577 (N_5577,N_5454,N_5309);
nor U5578 (N_5578,N_5295,N_5060);
nor U5579 (N_5579,N_5403,N_5269);
or U5580 (N_5580,N_5101,N_5007);
nor U5581 (N_5581,N_5366,N_5407);
nor U5582 (N_5582,N_5064,N_5437);
nand U5583 (N_5583,N_5014,N_5340);
nand U5584 (N_5584,N_5408,N_5025);
or U5585 (N_5585,N_5087,N_5030);
nand U5586 (N_5586,N_5452,N_5041);
or U5587 (N_5587,N_5010,N_5004);
nor U5588 (N_5588,N_5156,N_5082);
nor U5589 (N_5589,N_5306,N_5049);
or U5590 (N_5590,N_5294,N_5376);
and U5591 (N_5591,N_5017,N_5435);
or U5592 (N_5592,N_5052,N_5077);
and U5593 (N_5593,N_5080,N_5247);
nor U5594 (N_5594,N_5382,N_5099);
or U5595 (N_5595,N_5211,N_5176);
nor U5596 (N_5596,N_5266,N_5006);
nand U5597 (N_5597,N_5436,N_5219);
or U5598 (N_5598,N_5465,N_5029);
or U5599 (N_5599,N_5314,N_5130);
nand U5600 (N_5600,N_5324,N_5105);
nor U5601 (N_5601,N_5451,N_5472);
and U5602 (N_5602,N_5129,N_5457);
nor U5603 (N_5603,N_5112,N_5197);
nand U5604 (N_5604,N_5492,N_5301);
nor U5605 (N_5605,N_5118,N_5277);
nand U5606 (N_5606,N_5334,N_5022);
nor U5607 (N_5607,N_5428,N_5092);
or U5608 (N_5608,N_5217,N_5480);
nand U5609 (N_5609,N_5067,N_5345);
nor U5610 (N_5610,N_5391,N_5373);
nand U5611 (N_5611,N_5036,N_5402);
nor U5612 (N_5612,N_5134,N_5104);
nor U5613 (N_5613,N_5372,N_5142);
nor U5614 (N_5614,N_5137,N_5322);
nand U5615 (N_5615,N_5470,N_5350);
or U5616 (N_5616,N_5196,N_5001);
nor U5617 (N_5617,N_5009,N_5204);
nor U5618 (N_5618,N_5002,N_5395);
nand U5619 (N_5619,N_5473,N_5493);
xnor U5620 (N_5620,N_5389,N_5245);
nand U5621 (N_5621,N_5337,N_5369);
nand U5622 (N_5622,N_5265,N_5141);
or U5623 (N_5623,N_5352,N_5368);
nand U5624 (N_5624,N_5316,N_5343);
xnor U5625 (N_5625,N_5074,N_5085);
or U5626 (N_5626,N_5367,N_5494);
nand U5627 (N_5627,N_5433,N_5441);
nor U5628 (N_5628,N_5202,N_5370);
or U5629 (N_5629,N_5477,N_5164);
and U5630 (N_5630,N_5175,N_5222);
nor U5631 (N_5631,N_5374,N_5121);
nand U5632 (N_5632,N_5358,N_5096);
nor U5633 (N_5633,N_5114,N_5262);
nor U5634 (N_5634,N_5283,N_5221);
nor U5635 (N_5635,N_5377,N_5329);
or U5636 (N_5636,N_5396,N_5115);
and U5637 (N_5637,N_5305,N_5218);
nand U5638 (N_5638,N_5311,N_5254);
and U5639 (N_5639,N_5406,N_5070);
and U5640 (N_5640,N_5208,N_5120);
nor U5641 (N_5641,N_5320,N_5046);
nand U5642 (N_5642,N_5021,N_5260);
nand U5643 (N_5643,N_5276,N_5093);
nand U5644 (N_5644,N_5110,N_5468);
nand U5645 (N_5645,N_5261,N_5319);
or U5646 (N_5646,N_5349,N_5259);
nand U5647 (N_5647,N_5279,N_5039);
nor U5648 (N_5648,N_5278,N_5143);
nor U5649 (N_5649,N_5333,N_5499);
and U5650 (N_5650,N_5243,N_5387);
or U5651 (N_5651,N_5043,N_5271);
and U5652 (N_5652,N_5133,N_5483);
nor U5653 (N_5653,N_5292,N_5098);
and U5654 (N_5654,N_5476,N_5117);
nand U5655 (N_5655,N_5171,N_5200);
nor U5656 (N_5656,N_5426,N_5398);
nand U5657 (N_5657,N_5152,N_5286);
nand U5658 (N_5658,N_5220,N_5313);
or U5659 (N_5659,N_5399,N_5166);
nand U5660 (N_5660,N_5109,N_5419);
and U5661 (N_5661,N_5291,N_5089);
nand U5662 (N_5662,N_5119,N_5481);
and U5663 (N_5663,N_5125,N_5108);
or U5664 (N_5664,N_5489,N_5364);
nor U5665 (N_5665,N_5438,N_5068);
nand U5666 (N_5666,N_5095,N_5035);
nor U5667 (N_5667,N_5191,N_5047);
or U5668 (N_5668,N_5173,N_5365);
nor U5669 (N_5669,N_5302,N_5384);
nor U5670 (N_5670,N_5151,N_5420);
and U5671 (N_5671,N_5073,N_5058);
or U5672 (N_5672,N_5289,N_5378);
nand U5673 (N_5673,N_5307,N_5224);
and U5674 (N_5674,N_5037,N_5235);
and U5675 (N_5675,N_5409,N_5449);
nor U5676 (N_5676,N_5478,N_5424);
nor U5677 (N_5677,N_5136,N_5225);
or U5678 (N_5678,N_5189,N_5055);
nand U5679 (N_5679,N_5253,N_5163);
or U5680 (N_5680,N_5379,N_5248);
and U5681 (N_5681,N_5273,N_5392);
and U5682 (N_5682,N_5446,N_5184);
or U5683 (N_5683,N_5246,N_5193);
nor U5684 (N_5684,N_5252,N_5288);
and U5685 (N_5685,N_5223,N_5127);
nand U5686 (N_5686,N_5443,N_5045);
xor U5687 (N_5687,N_5051,N_5084);
or U5688 (N_5688,N_5086,N_5464);
nor U5689 (N_5689,N_5059,N_5038);
nor U5690 (N_5690,N_5107,N_5190);
nand U5691 (N_5691,N_5411,N_5159);
and U5692 (N_5692,N_5390,N_5375);
nand U5693 (N_5693,N_5381,N_5414);
and U5694 (N_5694,N_5495,N_5263);
and U5695 (N_5695,N_5415,N_5456);
xor U5696 (N_5696,N_5490,N_5185);
and U5697 (N_5697,N_5362,N_5126);
or U5698 (N_5698,N_5404,N_5326);
xnor U5699 (N_5699,N_5447,N_5300);
nand U5700 (N_5700,N_5050,N_5180);
nor U5701 (N_5701,N_5165,N_5091);
nand U5702 (N_5702,N_5325,N_5485);
and U5703 (N_5703,N_5013,N_5154);
nor U5704 (N_5704,N_5148,N_5297);
or U5705 (N_5705,N_5215,N_5459);
nand U5706 (N_5706,N_5209,N_5284);
nand U5707 (N_5707,N_5213,N_5236);
and U5708 (N_5708,N_5003,N_5275);
and U5709 (N_5709,N_5416,N_5187);
xnor U5710 (N_5710,N_5285,N_5062);
nor U5711 (N_5711,N_5498,N_5149);
or U5712 (N_5712,N_5338,N_5479);
and U5713 (N_5713,N_5147,N_5113);
nor U5714 (N_5714,N_5178,N_5020);
nand U5715 (N_5715,N_5042,N_5122);
and U5716 (N_5716,N_5354,N_5203);
nand U5717 (N_5717,N_5158,N_5356);
nand U5718 (N_5718,N_5195,N_5467);
nand U5719 (N_5719,N_5444,N_5423);
nor U5720 (N_5720,N_5491,N_5031);
nor U5721 (N_5721,N_5079,N_5287);
or U5722 (N_5722,N_5353,N_5413);
nor U5723 (N_5723,N_5361,N_5230);
or U5724 (N_5724,N_5321,N_5233);
nor U5725 (N_5725,N_5359,N_5181);
or U5726 (N_5726,N_5256,N_5018);
nand U5727 (N_5727,N_5210,N_5440);
or U5728 (N_5728,N_5304,N_5179);
and U5729 (N_5729,N_5066,N_5102);
nor U5730 (N_5730,N_5412,N_5194);
and U5731 (N_5731,N_5205,N_5238);
and U5732 (N_5732,N_5011,N_5186);
nand U5733 (N_5733,N_5044,N_5330);
and U5734 (N_5734,N_5380,N_5315);
and U5735 (N_5735,N_5150,N_5281);
nand U5736 (N_5736,N_5056,N_5312);
nor U5737 (N_5737,N_5169,N_5310);
and U5738 (N_5738,N_5081,N_5135);
and U5739 (N_5739,N_5207,N_5488);
nor U5740 (N_5740,N_5034,N_5418);
nor U5741 (N_5741,N_5445,N_5015);
nand U5742 (N_5742,N_5357,N_5032);
nand U5743 (N_5743,N_5453,N_5394);
nor U5744 (N_5744,N_5455,N_5290);
and U5745 (N_5745,N_5153,N_5341);
nor U5746 (N_5746,N_5272,N_5410);
or U5747 (N_5747,N_5496,N_5484);
nor U5748 (N_5748,N_5463,N_5332);
and U5749 (N_5749,N_5242,N_5063);
nor U5750 (N_5750,N_5015,N_5232);
nor U5751 (N_5751,N_5324,N_5215);
or U5752 (N_5752,N_5108,N_5415);
or U5753 (N_5753,N_5148,N_5449);
nand U5754 (N_5754,N_5056,N_5270);
and U5755 (N_5755,N_5122,N_5013);
nor U5756 (N_5756,N_5054,N_5095);
or U5757 (N_5757,N_5335,N_5162);
nor U5758 (N_5758,N_5266,N_5076);
or U5759 (N_5759,N_5341,N_5430);
nand U5760 (N_5760,N_5341,N_5298);
nor U5761 (N_5761,N_5015,N_5381);
nor U5762 (N_5762,N_5234,N_5458);
and U5763 (N_5763,N_5114,N_5467);
and U5764 (N_5764,N_5448,N_5050);
and U5765 (N_5765,N_5272,N_5232);
nor U5766 (N_5766,N_5251,N_5104);
nand U5767 (N_5767,N_5395,N_5378);
nor U5768 (N_5768,N_5446,N_5335);
nand U5769 (N_5769,N_5265,N_5435);
nor U5770 (N_5770,N_5187,N_5401);
or U5771 (N_5771,N_5021,N_5459);
and U5772 (N_5772,N_5312,N_5248);
nor U5773 (N_5773,N_5048,N_5045);
nor U5774 (N_5774,N_5420,N_5308);
and U5775 (N_5775,N_5473,N_5305);
or U5776 (N_5776,N_5262,N_5256);
and U5777 (N_5777,N_5493,N_5428);
nand U5778 (N_5778,N_5311,N_5457);
nand U5779 (N_5779,N_5197,N_5229);
or U5780 (N_5780,N_5460,N_5135);
and U5781 (N_5781,N_5167,N_5353);
and U5782 (N_5782,N_5290,N_5334);
nand U5783 (N_5783,N_5041,N_5433);
and U5784 (N_5784,N_5430,N_5484);
nor U5785 (N_5785,N_5161,N_5460);
nand U5786 (N_5786,N_5252,N_5022);
nand U5787 (N_5787,N_5322,N_5221);
nand U5788 (N_5788,N_5126,N_5470);
nor U5789 (N_5789,N_5191,N_5389);
or U5790 (N_5790,N_5411,N_5238);
and U5791 (N_5791,N_5263,N_5147);
nand U5792 (N_5792,N_5081,N_5401);
and U5793 (N_5793,N_5402,N_5072);
or U5794 (N_5794,N_5044,N_5262);
or U5795 (N_5795,N_5238,N_5057);
or U5796 (N_5796,N_5400,N_5172);
or U5797 (N_5797,N_5359,N_5438);
and U5798 (N_5798,N_5373,N_5154);
or U5799 (N_5799,N_5361,N_5055);
or U5800 (N_5800,N_5066,N_5263);
and U5801 (N_5801,N_5396,N_5117);
nand U5802 (N_5802,N_5167,N_5244);
nor U5803 (N_5803,N_5316,N_5165);
nor U5804 (N_5804,N_5033,N_5102);
and U5805 (N_5805,N_5342,N_5177);
nand U5806 (N_5806,N_5468,N_5415);
or U5807 (N_5807,N_5187,N_5179);
nor U5808 (N_5808,N_5145,N_5471);
or U5809 (N_5809,N_5304,N_5099);
or U5810 (N_5810,N_5196,N_5446);
nand U5811 (N_5811,N_5047,N_5307);
or U5812 (N_5812,N_5250,N_5460);
nor U5813 (N_5813,N_5225,N_5272);
nor U5814 (N_5814,N_5019,N_5380);
or U5815 (N_5815,N_5179,N_5220);
nor U5816 (N_5816,N_5175,N_5137);
or U5817 (N_5817,N_5313,N_5474);
or U5818 (N_5818,N_5057,N_5261);
or U5819 (N_5819,N_5017,N_5383);
and U5820 (N_5820,N_5363,N_5068);
nor U5821 (N_5821,N_5215,N_5412);
nand U5822 (N_5822,N_5469,N_5171);
nor U5823 (N_5823,N_5413,N_5247);
or U5824 (N_5824,N_5060,N_5284);
or U5825 (N_5825,N_5234,N_5413);
xor U5826 (N_5826,N_5278,N_5290);
and U5827 (N_5827,N_5112,N_5092);
nand U5828 (N_5828,N_5225,N_5054);
and U5829 (N_5829,N_5043,N_5481);
or U5830 (N_5830,N_5259,N_5034);
xor U5831 (N_5831,N_5191,N_5063);
nand U5832 (N_5832,N_5358,N_5427);
or U5833 (N_5833,N_5380,N_5166);
and U5834 (N_5834,N_5118,N_5296);
nor U5835 (N_5835,N_5425,N_5034);
and U5836 (N_5836,N_5295,N_5211);
or U5837 (N_5837,N_5193,N_5461);
and U5838 (N_5838,N_5044,N_5095);
and U5839 (N_5839,N_5022,N_5482);
nand U5840 (N_5840,N_5440,N_5341);
or U5841 (N_5841,N_5327,N_5322);
or U5842 (N_5842,N_5473,N_5471);
nor U5843 (N_5843,N_5462,N_5464);
or U5844 (N_5844,N_5271,N_5080);
and U5845 (N_5845,N_5274,N_5472);
nand U5846 (N_5846,N_5302,N_5150);
or U5847 (N_5847,N_5201,N_5189);
or U5848 (N_5848,N_5391,N_5372);
or U5849 (N_5849,N_5011,N_5249);
xnor U5850 (N_5850,N_5356,N_5497);
nor U5851 (N_5851,N_5201,N_5338);
nor U5852 (N_5852,N_5219,N_5169);
nor U5853 (N_5853,N_5338,N_5442);
xor U5854 (N_5854,N_5082,N_5187);
and U5855 (N_5855,N_5132,N_5352);
and U5856 (N_5856,N_5275,N_5122);
and U5857 (N_5857,N_5299,N_5226);
nor U5858 (N_5858,N_5177,N_5431);
and U5859 (N_5859,N_5410,N_5090);
nand U5860 (N_5860,N_5292,N_5401);
and U5861 (N_5861,N_5460,N_5196);
or U5862 (N_5862,N_5364,N_5279);
or U5863 (N_5863,N_5209,N_5238);
nand U5864 (N_5864,N_5018,N_5041);
nor U5865 (N_5865,N_5497,N_5343);
and U5866 (N_5866,N_5228,N_5338);
or U5867 (N_5867,N_5362,N_5423);
xor U5868 (N_5868,N_5159,N_5121);
nand U5869 (N_5869,N_5144,N_5063);
nand U5870 (N_5870,N_5246,N_5365);
nor U5871 (N_5871,N_5034,N_5217);
nor U5872 (N_5872,N_5021,N_5153);
nor U5873 (N_5873,N_5038,N_5024);
or U5874 (N_5874,N_5485,N_5382);
and U5875 (N_5875,N_5019,N_5058);
nand U5876 (N_5876,N_5432,N_5273);
nand U5877 (N_5877,N_5071,N_5483);
nor U5878 (N_5878,N_5075,N_5236);
or U5879 (N_5879,N_5205,N_5021);
nand U5880 (N_5880,N_5217,N_5164);
and U5881 (N_5881,N_5366,N_5082);
nor U5882 (N_5882,N_5275,N_5096);
or U5883 (N_5883,N_5494,N_5238);
nand U5884 (N_5884,N_5162,N_5015);
and U5885 (N_5885,N_5352,N_5448);
and U5886 (N_5886,N_5423,N_5174);
nand U5887 (N_5887,N_5116,N_5144);
and U5888 (N_5888,N_5146,N_5103);
nand U5889 (N_5889,N_5222,N_5300);
nor U5890 (N_5890,N_5300,N_5185);
or U5891 (N_5891,N_5493,N_5196);
nand U5892 (N_5892,N_5260,N_5355);
xnor U5893 (N_5893,N_5213,N_5063);
nand U5894 (N_5894,N_5298,N_5479);
or U5895 (N_5895,N_5220,N_5054);
xor U5896 (N_5896,N_5071,N_5010);
nand U5897 (N_5897,N_5135,N_5277);
and U5898 (N_5898,N_5088,N_5046);
and U5899 (N_5899,N_5054,N_5209);
nand U5900 (N_5900,N_5254,N_5379);
nand U5901 (N_5901,N_5310,N_5009);
or U5902 (N_5902,N_5287,N_5275);
nand U5903 (N_5903,N_5283,N_5119);
nor U5904 (N_5904,N_5002,N_5139);
nand U5905 (N_5905,N_5197,N_5000);
nor U5906 (N_5906,N_5106,N_5141);
and U5907 (N_5907,N_5350,N_5360);
or U5908 (N_5908,N_5283,N_5087);
nor U5909 (N_5909,N_5299,N_5006);
nor U5910 (N_5910,N_5247,N_5353);
and U5911 (N_5911,N_5401,N_5141);
nor U5912 (N_5912,N_5493,N_5335);
and U5913 (N_5913,N_5053,N_5441);
nor U5914 (N_5914,N_5422,N_5027);
nor U5915 (N_5915,N_5210,N_5018);
and U5916 (N_5916,N_5202,N_5135);
nor U5917 (N_5917,N_5423,N_5380);
nor U5918 (N_5918,N_5102,N_5401);
nor U5919 (N_5919,N_5121,N_5420);
nand U5920 (N_5920,N_5360,N_5247);
nand U5921 (N_5921,N_5412,N_5482);
nor U5922 (N_5922,N_5432,N_5231);
or U5923 (N_5923,N_5465,N_5052);
and U5924 (N_5924,N_5113,N_5246);
or U5925 (N_5925,N_5161,N_5136);
nor U5926 (N_5926,N_5358,N_5155);
nor U5927 (N_5927,N_5464,N_5411);
and U5928 (N_5928,N_5085,N_5173);
nor U5929 (N_5929,N_5341,N_5014);
nand U5930 (N_5930,N_5177,N_5375);
xor U5931 (N_5931,N_5421,N_5338);
nand U5932 (N_5932,N_5176,N_5237);
nor U5933 (N_5933,N_5173,N_5308);
and U5934 (N_5934,N_5206,N_5496);
nand U5935 (N_5935,N_5410,N_5412);
or U5936 (N_5936,N_5164,N_5459);
xor U5937 (N_5937,N_5087,N_5145);
or U5938 (N_5938,N_5027,N_5107);
and U5939 (N_5939,N_5194,N_5336);
or U5940 (N_5940,N_5025,N_5375);
nand U5941 (N_5941,N_5045,N_5028);
or U5942 (N_5942,N_5366,N_5190);
nand U5943 (N_5943,N_5300,N_5337);
nor U5944 (N_5944,N_5242,N_5178);
and U5945 (N_5945,N_5157,N_5399);
nor U5946 (N_5946,N_5138,N_5413);
or U5947 (N_5947,N_5425,N_5438);
and U5948 (N_5948,N_5436,N_5022);
nand U5949 (N_5949,N_5320,N_5462);
and U5950 (N_5950,N_5367,N_5380);
or U5951 (N_5951,N_5420,N_5040);
nor U5952 (N_5952,N_5126,N_5402);
nand U5953 (N_5953,N_5368,N_5323);
and U5954 (N_5954,N_5219,N_5279);
nor U5955 (N_5955,N_5077,N_5277);
and U5956 (N_5956,N_5410,N_5373);
nor U5957 (N_5957,N_5445,N_5332);
nor U5958 (N_5958,N_5248,N_5403);
nand U5959 (N_5959,N_5449,N_5269);
nand U5960 (N_5960,N_5437,N_5033);
nor U5961 (N_5961,N_5498,N_5354);
and U5962 (N_5962,N_5395,N_5242);
or U5963 (N_5963,N_5194,N_5118);
or U5964 (N_5964,N_5359,N_5131);
nor U5965 (N_5965,N_5106,N_5216);
nand U5966 (N_5966,N_5216,N_5253);
nor U5967 (N_5967,N_5235,N_5384);
or U5968 (N_5968,N_5374,N_5185);
or U5969 (N_5969,N_5424,N_5240);
nand U5970 (N_5970,N_5494,N_5406);
xnor U5971 (N_5971,N_5364,N_5092);
nand U5972 (N_5972,N_5138,N_5369);
nand U5973 (N_5973,N_5159,N_5074);
xnor U5974 (N_5974,N_5036,N_5175);
and U5975 (N_5975,N_5413,N_5113);
or U5976 (N_5976,N_5084,N_5106);
or U5977 (N_5977,N_5316,N_5496);
nor U5978 (N_5978,N_5378,N_5349);
or U5979 (N_5979,N_5106,N_5056);
and U5980 (N_5980,N_5094,N_5239);
nand U5981 (N_5981,N_5270,N_5409);
nand U5982 (N_5982,N_5338,N_5306);
nand U5983 (N_5983,N_5316,N_5047);
nand U5984 (N_5984,N_5072,N_5024);
and U5985 (N_5985,N_5357,N_5386);
nand U5986 (N_5986,N_5167,N_5074);
nand U5987 (N_5987,N_5117,N_5115);
nor U5988 (N_5988,N_5368,N_5250);
and U5989 (N_5989,N_5278,N_5044);
xor U5990 (N_5990,N_5330,N_5435);
or U5991 (N_5991,N_5078,N_5009);
and U5992 (N_5992,N_5334,N_5460);
or U5993 (N_5993,N_5289,N_5411);
nor U5994 (N_5994,N_5204,N_5259);
nand U5995 (N_5995,N_5223,N_5294);
nand U5996 (N_5996,N_5239,N_5276);
nand U5997 (N_5997,N_5367,N_5095);
and U5998 (N_5998,N_5321,N_5452);
or U5999 (N_5999,N_5206,N_5068);
nor U6000 (N_6000,N_5618,N_5982);
nor U6001 (N_6001,N_5698,N_5946);
and U6002 (N_6002,N_5539,N_5792);
nor U6003 (N_6003,N_5540,N_5641);
and U6004 (N_6004,N_5840,N_5744);
nor U6005 (N_6005,N_5870,N_5808);
or U6006 (N_6006,N_5644,N_5746);
nand U6007 (N_6007,N_5521,N_5750);
xnor U6008 (N_6008,N_5661,N_5938);
nor U6009 (N_6009,N_5510,N_5949);
xnor U6010 (N_6010,N_5724,N_5761);
or U6011 (N_6011,N_5885,N_5884);
nand U6012 (N_6012,N_5677,N_5914);
or U6013 (N_6013,N_5509,N_5570);
nand U6014 (N_6014,N_5787,N_5719);
nand U6015 (N_6015,N_5720,N_5821);
nand U6016 (N_6016,N_5906,N_5584);
nor U6017 (N_6017,N_5688,N_5924);
nand U6018 (N_6018,N_5827,N_5793);
or U6019 (N_6019,N_5846,N_5713);
nand U6020 (N_6020,N_5782,N_5554);
nand U6021 (N_6021,N_5614,N_5780);
or U6022 (N_6022,N_5843,N_5771);
and U6023 (N_6023,N_5933,N_5756);
nor U6024 (N_6024,N_5586,N_5910);
or U6025 (N_6025,N_5541,N_5980);
or U6026 (N_6026,N_5533,N_5805);
nand U6027 (N_6027,N_5546,N_5610);
nor U6028 (N_6028,N_5764,N_5944);
or U6029 (N_6029,N_5653,N_5684);
nor U6030 (N_6030,N_5623,N_5574);
nand U6031 (N_6031,N_5599,N_5550);
nand U6032 (N_6032,N_5703,N_5881);
and U6033 (N_6033,N_5536,N_5516);
nor U6034 (N_6034,N_5630,N_5887);
or U6035 (N_6035,N_5515,N_5812);
and U6036 (N_6036,N_5850,N_5851);
nor U6037 (N_6037,N_5833,N_5867);
and U6038 (N_6038,N_5942,N_5975);
or U6039 (N_6039,N_5642,N_5733);
or U6040 (N_6040,N_5935,N_5665);
nor U6041 (N_6041,N_5810,N_5525);
nand U6042 (N_6042,N_5549,N_5852);
and U6043 (N_6043,N_5594,N_5718);
nand U6044 (N_6044,N_5728,N_5693);
nand U6045 (N_6045,N_5514,N_5994);
and U6046 (N_6046,N_5662,N_5993);
and U6047 (N_6047,N_5847,N_5856);
nor U6048 (N_6048,N_5504,N_5936);
and U6049 (N_6049,N_5832,N_5822);
nor U6050 (N_6050,N_5760,N_5502);
and U6051 (N_6051,N_5562,N_5916);
and U6052 (N_6052,N_5894,N_5876);
or U6053 (N_6053,N_5537,N_5648);
xnor U6054 (N_6054,N_5604,N_5606);
and U6055 (N_6055,N_5730,N_5758);
nor U6056 (N_6056,N_5775,N_5889);
or U6057 (N_6057,N_5877,N_5818);
and U6058 (N_6058,N_5804,N_5528);
nand U6059 (N_6059,N_5700,N_5791);
nand U6060 (N_6060,N_5869,N_5951);
nor U6061 (N_6061,N_5954,N_5796);
nor U6062 (N_6062,N_5664,N_5666);
xor U6063 (N_6063,N_5825,N_5712);
nand U6064 (N_6064,N_5723,N_5786);
nor U6065 (N_6065,N_5826,N_5973);
or U6066 (N_6066,N_5567,N_5948);
or U6067 (N_6067,N_5895,N_5807);
or U6068 (N_6068,N_5683,N_5940);
or U6069 (N_6069,N_5842,N_5527);
nand U6070 (N_6070,N_5864,N_5689);
or U6071 (N_6071,N_5711,N_5830);
nand U6072 (N_6072,N_5501,N_5595);
or U6073 (N_6073,N_5937,N_5544);
nand U6074 (N_6074,N_5934,N_5592);
and U6075 (N_6075,N_5738,N_5809);
nand U6076 (N_6076,N_5646,N_5566);
nor U6077 (N_6077,N_5526,N_5617);
or U6078 (N_6078,N_5962,N_5878);
xor U6079 (N_6079,N_5841,N_5520);
nor U6080 (N_6080,N_5725,N_5800);
nor U6081 (N_6081,N_5619,N_5957);
xnor U6082 (N_6082,N_5687,N_5757);
or U6083 (N_6083,N_5972,N_5961);
and U6084 (N_6084,N_5577,N_5999);
nand U6085 (N_6085,N_5645,N_5849);
or U6086 (N_6086,N_5997,N_5890);
xnor U6087 (N_6087,N_5837,N_5500);
nor U6088 (N_6088,N_5919,N_5995);
nand U6089 (N_6089,N_5923,N_5695);
nand U6090 (N_6090,N_5788,N_5801);
or U6091 (N_6091,N_5569,N_5626);
and U6092 (N_6092,N_5838,N_5766);
and U6093 (N_6093,N_5704,N_5789);
and U6094 (N_6094,N_5803,N_5769);
nand U6095 (N_6095,N_5640,N_5605);
nand U6096 (N_6096,N_5799,N_5579);
nor U6097 (N_6097,N_5716,N_5779);
nor U6098 (N_6098,N_5759,N_5970);
nor U6099 (N_6099,N_5691,N_5522);
nor U6100 (N_6100,N_5545,N_5658);
and U6101 (N_6101,N_5968,N_5752);
nor U6102 (N_6102,N_5542,N_5998);
and U6103 (N_6103,N_5547,N_5920);
nand U6104 (N_6104,N_5952,N_5706);
nor U6105 (N_6105,N_5740,N_5503);
nand U6106 (N_6106,N_5941,N_5900);
or U6107 (N_6107,N_5866,N_5597);
nand U6108 (N_6108,N_5735,N_5573);
nand U6109 (N_6109,N_5848,N_5992);
or U6110 (N_6110,N_5690,N_5588);
or U6111 (N_6111,N_5722,N_5708);
and U6112 (N_6112,N_5663,N_5797);
or U6113 (N_6113,N_5902,N_5831);
nand U6114 (N_6114,N_5697,N_5839);
or U6115 (N_6115,N_5639,N_5603);
nand U6116 (N_6116,N_5580,N_5670);
nand U6117 (N_6117,N_5806,N_5679);
nor U6118 (N_6118,N_5748,N_5552);
and U6119 (N_6119,N_5873,N_5783);
or U6120 (N_6120,N_5702,N_5829);
and U6121 (N_6121,N_5753,N_5508);
nand U6122 (N_6122,N_5754,N_5671);
or U6123 (N_6123,N_5749,N_5958);
nand U6124 (N_6124,N_5581,N_5602);
nand U6125 (N_6125,N_5600,N_5907);
or U6126 (N_6126,N_5676,N_5633);
nand U6127 (N_6127,N_5932,N_5795);
nor U6128 (N_6128,N_5755,N_5621);
nor U6129 (N_6129,N_5917,N_5969);
nand U6130 (N_6130,N_5765,N_5731);
and U6131 (N_6131,N_5991,N_5798);
or U6132 (N_6132,N_5726,N_5925);
nor U6133 (N_6133,N_5741,N_5709);
or U6134 (N_6134,N_5669,N_5572);
and U6135 (N_6135,N_5911,N_5772);
or U6136 (N_6136,N_5901,N_5931);
or U6137 (N_6137,N_5548,N_5823);
and U6138 (N_6138,N_5861,N_5654);
and U6139 (N_6139,N_5612,N_5507);
nor U6140 (N_6140,N_5784,N_5745);
nor U6141 (N_6141,N_5737,N_5678);
and U6142 (N_6142,N_5715,N_5794);
nor U6143 (N_6143,N_5694,N_5979);
and U6144 (N_6144,N_5875,N_5717);
and U6145 (N_6145,N_5751,N_5622);
nand U6146 (N_6146,N_5627,N_5732);
or U6147 (N_6147,N_5816,N_5776);
or U6148 (N_6148,N_5930,N_5777);
nor U6149 (N_6149,N_5965,N_5986);
nand U6150 (N_6150,N_5845,N_5564);
nand U6151 (N_6151,N_5988,N_5710);
and U6152 (N_6152,N_5767,N_5611);
nand U6153 (N_6153,N_5616,N_5817);
or U6154 (N_6154,N_5506,N_5976);
nand U6155 (N_6155,N_5768,N_5868);
or U6156 (N_6156,N_5883,N_5747);
xnor U6157 (N_6157,N_5964,N_5535);
nand U6158 (N_6158,N_5774,N_5634);
nor U6159 (N_6159,N_5707,N_5859);
and U6160 (N_6160,N_5828,N_5729);
nor U6161 (N_6161,N_5559,N_5512);
nor U6162 (N_6162,N_5971,N_5686);
nand U6163 (N_6163,N_5929,N_5888);
and U6164 (N_6164,N_5680,N_5908);
nor U6165 (N_6165,N_5561,N_5519);
nor U6166 (N_6166,N_5762,N_5596);
nor U6167 (N_6167,N_5913,N_5682);
and U6168 (N_6168,N_5736,N_5672);
or U6169 (N_6169,N_5739,N_5956);
nand U6170 (N_6170,N_5989,N_5898);
nand U6171 (N_6171,N_5593,N_5770);
nand U6172 (N_6172,N_5523,N_5987);
nand U6173 (N_6173,N_5629,N_5624);
nand U6174 (N_6174,N_5854,N_5576);
or U6175 (N_6175,N_5657,N_5863);
nor U6176 (N_6176,N_5966,N_5696);
or U6177 (N_6177,N_5880,N_5601);
and U6178 (N_6178,N_5530,N_5977);
and U6179 (N_6179,N_5555,N_5638);
or U6180 (N_6180,N_5844,N_5862);
and U6181 (N_6181,N_5814,N_5763);
or U6182 (N_6182,N_5882,N_5699);
nand U6183 (N_6183,N_5967,N_5781);
and U6184 (N_6184,N_5921,N_5990);
nor U6185 (N_6185,N_5674,N_5532);
or U6186 (N_6186,N_5557,N_5636);
nor U6187 (N_6187,N_5587,N_5872);
or U6188 (N_6188,N_5649,N_5897);
or U6189 (N_6189,N_5529,N_5891);
and U6190 (N_6190,N_5834,N_5615);
or U6191 (N_6191,N_5815,N_5912);
and U6192 (N_6192,N_5893,N_5945);
and U6193 (N_6193,N_5865,N_5583);
or U6194 (N_6194,N_5556,N_5608);
and U6195 (N_6195,N_5551,N_5538);
or U6196 (N_6196,N_5860,N_5896);
or U6197 (N_6197,N_5668,N_5613);
and U6198 (N_6198,N_5978,N_5675);
nand U6199 (N_6199,N_5785,N_5534);
and U6200 (N_6200,N_5681,N_5558);
or U6201 (N_6201,N_5963,N_5820);
xnor U6202 (N_6202,N_5743,N_5959);
or U6203 (N_6203,N_5905,N_5926);
or U6204 (N_6204,N_5524,N_5589);
and U6205 (N_6205,N_5590,N_5582);
nand U6206 (N_6206,N_5655,N_5607);
nor U6207 (N_6207,N_5778,N_5628);
nand U6208 (N_6208,N_5563,N_5714);
nor U6209 (N_6209,N_5836,N_5631);
nand U6210 (N_6210,N_5651,N_5955);
and U6211 (N_6211,N_5568,N_5647);
nand U6212 (N_6212,N_5835,N_5996);
nor U6213 (N_6213,N_5802,N_5824);
or U6214 (N_6214,N_5518,N_5667);
or U6215 (N_6215,N_5575,N_5773);
nor U6216 (N_6216,N_5953,N_5909);
or U6217 (N_6217,N_5927,N_5673);
nand U6218 (N_6218,N_5635,N_5659);
or U6219 (N_6219,N_5981,N_5790);
or U6220 (N_6220,N_5734,N_5578);
nor U6221 (N_6221,N_5939,N_5625);
or U6222 (N_6222,N_5918,N_5650);
xnor U6223 (N_6223,N_5571,N_5560);
xnor U6224 (N_6224,N_5922,N_5643);
or U6225 (N_6225,N_5984,N_5513);
nand U6226 (N_6226,N_5853,N_5656);
nor U6227 (N_6227,N_5947,N_5637);
and U6228 (N_6228,N_5915,N_5685);
or U6229 (N_6229,N_5857,N_5813);
and U6230 (N_6230,N_5701,N_5705);
or U6231 (N_6231,N_5505,N_5886);
nand U6232 (N_6232,N_5543,N_5943);
nor U6233 (N_6233,N_5874,N_5858);
nor U6234 (N_6234,N_5928,N_5742);
nand U6235 (N_6235,N_5879,N_5531);
nor U6236 (N_6236,N_5511,N_5983);
xor U6237 (N_6237,N_5985,N_5904);
and U6238 (N_6238,N_5960,N_5811);
nor U6239 (N_6239,N_5652,N_5598);
or U6240 (N_6240,N_5632,N_5721);
xnor U6241 (N_6241,N_5899,N_5620);
nor U6242 (N_6242,N_5727,N_5692);
or U6243 (N_6243,N_5871,N_5892);
or U6244 (N_6244,N_5819,N_5855);
or U6245 (N_6245,N_5517,N_5553);
and U6246 (N_6246,N_5660,N_5591);
nand U6247 (N_6247,N_5585,N_5609);
nor U6248 (N_6248,N_5565,N_5903);
or U6249 (N_6249,N_5974,N_5950);
nand U6250 (N_6250,N_5937,N_5576);
and U6251 (N_6251,N_5714,N_5520);
and U6252 (N_6252,N_5885,N_5677);
nand U6253 (N_6253,N_5965,N_5623);
or U6254 (N_6254,N_5866,N_5698);
and U6255 (N_6255,N_5951,N_5699);
nor U6256 (N_6256,N_5595,N_5738);
and U6257 (N_6257,N_5939,N_5947);
or U6258 (N_6258,N_5630,N_5805);
nor U6259 (N_6259,N_5953,N_5820);
nor U6260 (N_6260,N_5945,N_5676);
nand U6261 (N_6261,N_5795,N_5676);
nor U6262 (N_6262,N_5760,N_5636);
or U6263 (N_6263,N_5584,N_5691);
xnor U6264 (N_6264,N_5545,N_5926);
or U6265 (N_6265,N_5986,N_5768);
or U6266 (N_6266,N_5883,N_5751);
or U6267 (N_6267,N_5837,N_5600);
and U6268 (N_6268,N_5514,N_5513);
or U6269 (N_6269,N_5648,N_5926);
nand U6270 (N_6270,N_5857,N_5613);
nand U6271 (N_6271,N_5695,N_5980);
and U6272 (N_6272,N_5961,N_5868);
nor U6273 (N_6273,N_5867,N_5550);
or U6274 (N_6274,N_5520,N_5897);
nand U6275 (N_6275,N_5910,N_5505);
or U6276 (N_6276,N_5832,N_5644);
nand U6277 (N_6277,N_5680,N_5512);
nand U6278 (N_6278,N_5525,N_5900);
nor U6279 (N_6279,N_5886,N_5750);
and U6280 (N_6280,N_5731,N_5992);
or U6281 (N_6281,N_5912,N_5593);
nand U6282 (N_6282,N_5868,N_5812);
and U6283 (N_6283,N_5756,N_5765);
nand U6284 (N_6284,N_5697,N_5689);
and U6285 (N_6285,N_5630,N_5855);
nand U6286 (N_6286,N_5650,N_5885);
nand U6287 (N_6287,N_5893,N_5521);
or U6288 (N_6288,N_5769,N_5940);
nor U6289 (N_6289,N_5984,N_5507);
nand U6290 (N_6290,N_5658,N_5976);
and U6291 (N_6291,N_5580,N_5718);
and U6292 (N_6292,N_5507,N_5633);
and U6293 (N_6293,N_5938,N_5833);
and U6294 (N_6294,N_5966,N_5709);
or U6295 (N_6295,N_5606,N_5791);
nor U6296 (N_6296,N_5882,N_5648);
nor U6297 (N_6297,N_5773,N_5935);
nand U6298 (N_6298,N_5614,N_5909);
or U6299 (N_6299,N_5884,N_5663);
nand U6300 (N_6300,N_5667,N_5777);
and U6301 (N_6301,N_5503,N_5915);
or U6302 (N_6302,N_5986,N_5757);
or U6303 (N_6303,N_5810,N_5807);
or U6304 (N_6304,N_5922,N_5812);
nor U6305 (N_6305,N_5923,N_5532);
and U6306 (N_6306,N_5954,N_5866);
nand U6307 (N_6307,N_5993,N_5599);
or U6308 (N_6308,N_5554,N_5995);
and U6309 (N_6309,N_5810,N_5969);
nand U6310 (N_6310,N_5706,N_5979);
or U6311 (N_6311,N_5657,N_5976);
nor U6312 (N_6312,N_5544,N_5526);
or U6313 (N_6313,N_5616,N_5632);
and U6314 (N_6314,N_5500,N_5708);
nor U6315 (N_6315,N_5849,N_5919);
or U6316 (N_6316,N_5535,N_5702);
or U6317 (N_6317,N_5620,N_5915);
nand U6318 (N_6318,N_5635,N_5926);
nand U6319 (N_6319,N_5825,N_5635);
or U6320 (N_6320,N_5717,N_5707);
nor U6321 (N_6321,N_5833,N_5905);
nor U6322 (N_6322,N_5756,N_5793);
nand U6323 (N_6323,N_5859,N_5655);
or U6324 (N_6324,N_5508,N_5679);
nand U6325 (N_6325,N_5803,N_5917);
nand U6326 (N_6326,N_5625,N_5936);
nand U6327 (N_6327,N_5576,N_5749);
and U6328 (N_6328,N_5915,N_5731);
nor U6329 (N_6329,N_5845,N_5824);
and U6330 (N_6330,N_5862,N_5535);
and U6331 (N_6331,N_5754,N_5692);
and U6332 (N_6332,N_5834,N_5653);
nand U6333 (N_6333,N_5693,N_5954);
or U6334 (N_6334,N_5514,N_5744);
and U6335 (N_6335,N_5520,N_5951);
or U6336 (N_6336,N_5635,N_5543);
nor U6337 (N_6337,N_5571,N_5513);
nor U6338 (N_6338,N_5509,N_5606);
nor U6339 (N_6339,N_5721,N_5985);
and U6340 (N_6340,N_5926,N_5663);
and U6341 (N_6341,N_5957,N_5567);
nor U6342 (N_6342,N_5827,N_5578);
or U6343 (N_6343,N_5914,N_5920);
nor U6344 (N_6344,N_5759,N_5920);
or U6345 (N_6345,N_5687,N_5732);
nand U6346 (N_6346,N_5923,N_5635);
and U6347 (N_6347,N_5674,N_5727);
or U6348 (N_6348,N_5771,N_5534);
or U6349 (N_6349,N_5622,N_5634);
nand U6350 (N_6350,N_5708,N_5677);
or U6351 (N_6351,N_5787,N_5995);
nand U6352 (N_6352,N_5581,N_5552);
and U6353 (N_6353,N_5681,N_5743);
and U6354 (N_6354,N_5627,N_5743);
nor U6355 (N_6355,N_5899,N_5532);
or U6356 (N_6356,N_5508,N_5550);
nand U6357 (N_6357,N_5599,N_5719);
nand U6358 (N_6358,N_5740,N_5774);
or U6359 (N_6359,N_5697,N_5869);
or U6360 (N_6360,N_5807,N_5913);
and U6361 (N_6361,N_5994,N_5883);
nand U6362 (N_6362,N_5578,N_5920);
nor U6363 (N_6363,N_5552,N_5796);
nor U6364 (N_6364,N_5851,N_5582);
nor U6365 (N_6365,N_5602,N_5961);
or U6366 (N_6366,N_5725,N_5528);
nand U6367 (N_6367,N_5885,N_5876);
nand U6368 (N_6368,N_5980,N_5830);
or U6369 (N_6369,N_5845,N_5504);
and U6370 (N_6370,N_5515,N_5677);
nor U6371 (N_6371,N_5814,N_5719);
or U6372 (N_6372,N_5724,N_5827);
nand U6373 (N_6373,N_5597,N_5875);
and U6374 (N_6374,N_5645,N_5949);
nor U6375 (N_6375,N_5715,N_5661);
nor U6376 (N_6376,N_5959,N_5989);
or U6377 (N_6377,N_5758,N_5785);
and U6378 (N_6378,N_5721,N_5663);
or U6379 (N_6379,N_5813,N_5567);
nor U6380 (N_6380,N_5537,N_5741);
and U6381 (N_6381,N_5589,N_5626);
and U6382 (N_6382,N_5540,N_5506);
nand U6383 (N_6383,N_5973,N_5748);
or U6384 (N_6384,N_5511,N_5502);
or U6385 (N_6385,N_5593,N_5804);
and U6386 (N_6386,N_5826,N_5582);
or U6387 (N_6387,N_5904,N_5628);
nand U6388 (N_6388,N_5875,N_5686);
xnor U6389 (N_6389,N_5973,N_5921);
and U6390 (N_6390,N_5876,N_5836);
nor U6391 (N_6391,N_5752,N_5536);
or U6392 (N_6392,N_5803,N_5510);
or U6393 (N_6393,N_5587,N_5971);
nor U6394 (N_6394,N_5742,N_5915);
and U6395 (N_6395,N_5768,N_5562);
and U6396 (N_6396,N_5597,N_5805);
and U6397 (N_6397,N_5899,N_5938);
and U6398 (N_6398,N_5968,N_5950);
or U6399 (N_6399,N_5896,N_5714);
nand U6400 (N_6400,N_5992,N_5755);
or U6401 (N_6401,N_5646,N_5550);
or U6402 (N_6402,N_5500,N_5592);
nand U6403 (N_6403,N_5877,N_5841);
or U6404 (N_6404,N_5694,N_5939);
nand U6405 (N_6405,N_5592,N_5693);
nand U6406 (N_6406,N_5786,N_5540);
nand U6407 (N_6407,N_5951,N_5873);
nor U6408 (N_6408,N_5807,N_5640);
nor U6409 (N_6409,N_5667,N_5632);
nor U6410 (N_6410,N_5598,N_5937);
or U6411 (N_6411,N_5925,N_5663);
nand U6412 (N_6412,N_5571,N_5761);
nand U6413 (N_6413,N_5767,N_5825);
nand U6414 (N_6414,N_5950,N_5713);
and U6415 (N_6415,N_5591,N_5645);
nand U6416 (N_6416,N_5602,N_5901);
nand U6417 (N_6417,N_5667,N_5666);
nor U6418 (N_6418,N_5729,N_5808);
or U6419 (N_6419,N_5611,N_5578);
and U6420 (N_6420,N_5864,N_5950);
nor U6421 (N_6421,N_5564,N_5591);
and U6422 (N_6422,N_5744,N_5565);
nand U6423 (N_6423,N_5986,N_5888);
nand U6424 (N_6424,N_5507,N_5953);
or U6425 (N_6425,N_5716,N_5840);
nand U6426 (N_6426,N_5595,N_5874);
or U6427 (N_6427,N_5949,N_5885);
nor U6428 (N_6428,N_5842,N_5534);
nand U6429 (N_6429,N_5978,N_5856);
nor U6430 (N_6430,N_5675,N_5740);
and U6431 (N_6431,N_5653,N_5935);
nor U6432 (N_6432,N_5998,N_5870);
or U6433 (N_6433,N_5821,N_5801);
nor U6434 (N_6434,N_5838,N_5723);
or U6435 (N_6435,N_5861,N_5506);
nor U6436 (N_6436,N_5553,N_5606);
and U6437 (N_6437,N_5885,N_5538);
nor U6438 (N_6438,N_5782,N_5558);
nand U6439 (N_6439,N_5607,N_5557);
and U6440 (N_6440,N_5992,N_5903);
or U6441 (N_6441,N_5999,N_5968);
nand U6442 (N_6442,N_5673,N_5761);
or U6443 (N_6443,N_5851,N_5620);
and U6444 (N_6444,N_5570,N_5849);
nor U6445 (N_6445,N_5975,N_5539);
nand U6446 (N_6446,N_5811,N_5729);
nand U6447 (N_6447,N_5899,N_5905);
or U6448 (N_6448,N_5790,N_5730);
nand U6449 (N_6449,N_5742,N_5998);
nor U6450 (N_6450,N_5729,N_5807);
and U6451 (N_6451,N_5878,N_5958);
and U6452 (N_6452,N_5571,N_5767);
nor U6453 (N_6453,N_5626,N_5622);
or U6454 (N_6454,N_5524,N_5698);
and U6455 (N_6455,N_5767,N_5618);
and U6456 (N_6456,N_5661,N_5882);
or U6457 (N_6457,N_5902,N_5791);
or U6458 (N_6458,N_5772,N_5646);
or U6459 (N_6459,N_5870,N_5510);
and U6460 (N_6460,N_5881,N_5947);
and U6461 (N_6461,N_5742,N_5892);
and U6462 (N_6462,N_5853,N_5841);
nand U6463 (N_6463,N_5539,N_5893);
nand U6464 (N_6464,N_5947,N_5996);
nor U6465 (N_6465,N_5663,N_5986);
or U6466 (N_6466,N_5761,N_5732);
or U6467 (N_6467,N_5533,N_5633);
xor U6468 (N_6468,N_5855,N_5687);
nand U6469 (N_6469,N_5663,N_5752);
and U6470 (N_6470,N_5645,N_5689);
nand U6471 (N_6471,N_5856,N_5840);
nor U6472 (N_6472,N_5981,N_5527);
nor U6473 (N_6473,N_5735,N_5542);
nand U6474 (N_6474,N_5581,N_5937);
or U6475 (N_6475,N_5561,N_5794);
and U6476 (N_6476,N_5821,N_5793);
nor U6477 (N_6477,N_5764,N_5956);
and U6478 (N_6478,N_5580,N_5898);
and U6479 (N_6479,N_5758,N_5560);
nand U6480 (N_6480,N_5942,N_5836);
or U6481 (N_6481,N_5707,N_5598);
or U6482 (N_6482,N_5805,N_5964);
nand U6483 (N_6483,N_5583,N_5629);
nand U6484 (N_6484,N_5984,N_5647);
nand U6485 (N_6485,N_5671,N_5513);
nor U6486 (N_6486,N_5542,N_5852);
nor U6487 (N_6487,N_5515,N_5656);
and U6488 (N_6488,N_5631,N_5857);
nor U6489 (N_6489,N_5998,N_5841);
and U6490 (N_6490,N_5719,N_5808);
nand U6491 (N_6491,N_5695,N_5538);
and U6492 (N_6492,N_5681,N_5567);
nand U6493 (N_6493,N_5971,N_5575);
nor U6494 (N_6494,N_5904,N_5507);
nor U6495 (N_6495,N_5615,N_5794);
nor U6496 (N_6496,N_5887,N_5676);
nand U6497 (N_6497,N_5640,N_5912);
and U6498 (N_6498,N_5659,N_5961);
nor U6499 (N_6499,N_5609,N_5590);
or U6500 (N_6500,N_6180,N_6450);
or U6501 (N_6501,N_6182,N_6032);
nor U6502 (N_6502,N_6200,N_6239);
nor U6503 (N_6503,N_6287,N_6465);
nor U6504 (N_6504,N_6463,N_6270);
or U6505 (N_6505,N_6135,N_6376);
and U6506 (N_6506,N_6486,N_6215);
and U6507 (N_6507,N_6003,N_6179);
nand U6508 (N_6508,N_6093,N_6153);
nand U6509 (N_6509,N_6046,N_6106);
nor U6510 (N_6510,N_6255,N_6475);
nor U6511 (N_6511,N_6053,N_6000);
nor U6512 (N_6512,N_6452,N_6407);
nand U6513 (N_6513,N_6216,N_6298);
xnor U6514 (N_6514,N_6131,N_6211);
nand U6515 (N_6515,N_6055,N_6394);
or U6516 (N_6516,N_6184,N_6326);
nor U6517 (N_6517,N_6063,N_6162);
nand U6518 (N_6518,N_6393,N_6345);
or U6519 (N_6519,N_6439,N_6022);
and U6520 (N_6520,N_6142,N_6299);
nand U6521 (N_6521,N_6488,N_6068);
nand U6522 (N_6522,N_6399,N_6444);
nor U6523 (N_6523,N_6476,N_6001);
nor U6524 (N_6524,N_6327,N_6372);
or U6525 (N_6525,N_6487,N_6420);
and U6526 (N_6526,N_6169,N_6462);
or U6527 (N_6527,N_6230,N_6227);
nand U6528 (N_6528,N_6258,N_6234);
xnor U6529 (N_6529,N_6176,N_6322);
and U6530 (N_6530,N_6181,N_6262);
nor U6531 (N_6531,N_6281,N_6132);
nand U6532 (N_6532,N_6099,N_6477);
nand U6533 (N_6533,N_6056,N_6336);
nor U6534 (N_6534,N_6461,N_6037);
nor U6535 (N_6535,N_6263,N_6449);
and U6536 (N_6536,N_6335,N_6124);
or U6537 (N_6537,N_6061,N_6283);
nor U6538 (N_6538,N_6458,N_6079);
nor U6539 (N_6539,N_6341,N_6256);
nor U6540 (N_6540,N_6286,N_6346);
nand U6541 (N_6541,N_6254,N_6233);
nor U6542 (N_6542,N_6279,N_6082);
or U6543 (N_6543,N_6014,N_6494);
nor U6544 (N_6544,N_6212,N_6221);
or U6545 (N_6545,N_6006,N_6315);
or U6546 (N_6546,N_6272,N_6409);
and U6547 (N_6547,N_6455,N_6277);
and U6548 (N_6548,N_6342,N_6267);
nor U6549 (N_6549,N_6284,N_6357);
or U6550 (N_6550,N_6163,N_6447);
or U6551 (N_6551,N_6320,N_6173);
nand U6552 (N_6552,N_6222,N_6060);
nor U6553 (N_6553,N_6021,N_6261);
or U6554 (N_6554,N_6490,N_6011);
nor U6555 (N_6555,N_6023,N_6199);
or U6556 (N_6556,N_6347,N_6107);
and U6557 (N_6557,N_6292,N_6363);
or U6558 (N_6558,N_6479,N_6004);
and U6559 (N_6559,N_6139,N_6090);
nand U6560 (N_6560,N_6058,N_6469);
nor U6561 (N_6561,N_6291,N_6094);
and U6562 (N_6562,N_6120,N_6325);
nor U6563 (N_6563,N_6097,N_6166);
or U6564 (N_6564,N_6430,N_6115);
nand U6565 (N_6565,N_6373,N_6196);
nand U6566 (N_6566,N_6008,N_6489);
nor U6567 (N_6567,N_6497,N_6240);
or U6568 (N_6568,N_6020,N_6382);
and U6569 (N_6569,N_6189,N_6413);
or U6570 (N_6570,N_6446,N_6377);
nand U6571 (N_6571,N_6312,N_6136);
nand U6572 (N_6572,N_6033,N_6116);
and U6573 (N_6573,N_6236,N_6086);
or U6574 (N_6574,N_6334,N_6105);
or U6575 (N_6575,N_6483,N_6380);
or U6576 (N_6576,N_6043,N_6297);
nor U6577 (N_6577,N_6433,N_6171);
nor U6578 (N_6578,N_6231,N_6057);
or U6579 (N_6579,N_6134,N_6353);
or U6580 (N_6580,N_6348,N_6493);
nand U6581 (N_6581,N_6137,N_6225);
nand U6582 (N_6582,N_6141,N_6203);
and U6583 (N_6583,N_6114,N_6138);
and U6584 (N_6584,N_6400,N_6030);
nand U6585 (N_6585,N_6146,N_6470);
nand U6586 (N_6586,N_6391,N_6285);
nand U6587 (N_6587,N_6226,N_6229);
or U6588 (N_6588,N_6083,N_6499);
and U6589 (N_6589,N_6340,N_6350);
or U6590 (N_6590,N_6319,N_6029);
xnor U6591 (N_6591,N_6157,N_6337);
or U6592 (N_6592,N_6034,N_6208);
and U6593 (N_6593,N_6054,N_6091);
nor U6594 (N_6594,N_6431,N_6425);
nand U6595 (N_6595,N_6388,N_6121);
nor U6596 (N_6596,N_6009,N_6456);
and U6597 (N_6597,N_6491,N_6117);
and U6598 (N_6598,N_6251,N_6355);
nor U6599 (N_6599,N_6126,N_6036);
or U6600 (N_6600,N_6160,N_6035);
or U6601 (N_6601,N_6156,N_6453);
nand U6602 (N_6602,N_6219,N_6265);
nor U6603 (N_6603,N_6062,N_6459);
nor U6604 (N_6604,N_6024,N_6412);
nand U6605 (N_6605,N_6218,N_6468);
or U6606 (N_6606,N_6178,N_6276);
or U6607 (N_6607,N_6111,N_6411);
or U6608 (N_6608,N_6358,N_6323);
nor U6609 (N_6609,N_6457,N_6300);
nor U6610 (N_6610,N_6419,N_6332);
or U6611 (N_6611,N_6275,N_6370);
nor U6612 (N_6612,N_6076,N_6213);
or U6613 (N_6613,N_6209,N_6371);
nor U6614 (N_6614,N_6460,N_6442);
nand U6615 (N_6615,N_6404,N_6390);
xnor U6616 (N_6616,N_6250,N_6129);
or U6617 (N_6617,N_6220,N_6038);
nor U6618 (N_6618,N_6144,N_6271);
xnor U6619 (N_6619,N_6402,N_6081);
nand U6620 (N_6620,N_6268,N_6017);
nand U6621 (N_6621,N_6464,N_6127);
and U6622 (N_6622,N_6059,N_6274);
nor U6623 (N_6623,N_6122,N_6387);
and U6624 (N_6624,N_6496,N_6428);
nand U6625 (N_6625,N_6405,N_6311);
nor U6626 (N_6626,N_6324,N_6410);
or U6627 (N_6627,N_6047,N_6290);
nand U6628 (N_6628,N_6302,N_6403);
and U6629 (N_6629,N_6232,N_6374);
and U6630 (N_6630,N_6167,N_6108);
xor U6631 (N_6631,N_6197,N_6080);
nor U6632 (N_6632,N_6188,N_6010);
and U6633 (N_6633,N_6352,N_6454);
nand U6634 (N_6634,N_6472,N_6308);
or U6635 (N_6635,N_6362,N_6165);
and U6636 (N_6636,N_6466,N_6205);
and U6637 (N_6637,N_6329,N_6448);
nand U6638 (N_6638,N_6128,N_6133);
or U6639 (N_6639,N_6422,N_6103);
nor U6640 (N_6640,N_6339,N_6273);
or U6641 (N_6641,N_6198,N_6088);
and U6642 (N_6642,N_6074,N_6481);
nor U6643 (N_6643,N_6228,N_6044);
and U6644 (N_6644,N_6386,N_6065);
nand U6645 (N_6645,N_6406,N_6306);
nor U6646 (N_6646,N_6257,N_6084);
and U6647 (N_6647,N_6396,N_6066);
nand U6648 (N_6648,N_6092,N_6241);
nand U6649 (N_6649,N_6395,N_6474);
or U6650 (N_6650,N_6143,N_6002);
nand U6651 (N_6651,N_6042,N_6045);
and U6652 (N_6652,N_6039,N_6366);
or U6653 (N_6653,N_6098,N_6201);
or U6654 (N_6654,N_6151,N_6304);
nand U6655 (N_6655,N_6295,N_6204);
or U6656 (N_6656,N_6480,N_6440);
and U6657 (N_6657,N_6492,N_6186);
or U6658 (N_6658,N_6244,N_6149);
or U6659 (N_6659,N_6025,N_6113);
nor U6660 (N_6660,N_6102,N_6170);
nor U6661 (N_6661,N_6223,N_6177);
or U6662 (N_6662,N_6217,N_6049);
or U6663 (N_6663,N_6018,N_6130);
and U6664 (N_6664,N_6161,N_6207);
and U6665 (N_6665,N_6148,N_6206);
nand U6666 (N_6666,N_6360,N_6417);
and U6667 (N_6667,N_6288,N_6005);
and U6668 (N_6668,N_6224,N_6289);
nor U6669 (N_6669,N_6147,N_6085);
nand U6670 (N_6670,N_6072,N_6125);
or U6671 (N_6671,N_6109,N_6193);
xnor U6672 (N_6672,N_6089,N_6351);
or U6673 (N_6673,N_6155,N_6026);
or U6674 (N_6674,N_6172,N_6112);
or U6675 (N_6675,N_6140,N_6443);
nand U6676 (N_6676,N_6194,N_6482);
xnor U6677 (N_6677,N_6359,N_6260);
nand U6678 (N_6678,N_6484,N_6445);
nor U6679 (N_6679,N_6012,N_6408);
nor U6680 (N_6680,N_6118,N_6451);
nand U6681 (N_6681,N_6389,N_6331);
nand U6682 (N_6682,N_6101,N_6152);
nand U6683 (N_6683,N_6145,N_6031);
and U6684 (N_6684,N_6243,N_6361);
or U6685 (N_6685,N_6249,N_6238);
nor U6686 (N_6686,N_6245,N_6296);
nor U6687 (N_6687,N_6191,N_6478);
nor U6688 (N_6688,N_6187,N_6168);
and U6689 (N_6689,N_6498,N_6075);
and U6690 (N_6690,N_6367,N_6242);
nand U6691 (N_6691,N_6195,N_6266);
or U6692 (N_6692,N_6154,N_6343);
nor U6693 (N_6693,N_6423,N_6473);
nor U6694 (N_6694,N_6383,N_6333);
or U6695 (N_6695,N_6307,N_6158);
nand U6696 (N_6696,N_6314,N_6190);
nor U6697 (N_6697,N_6071,N_6100);
nand U6698 (N_6698,N_6384,N_6040);
nand U6699 (N_6699,N_6070,N_6248);
or U6700 (N_6700,N_6150,N_6175);
and U6701 (N_6701,N_6310,N_6344);
nand U6702 (N_6702,N_6426,N_6379);
or U6703 (N_6703,N_6051,N_6278);
and U6704 (N_6704,N_6338,N_6305);
nand U6705 (N_6705,N_6415,N_6159);
nand U6706 (N_6706,N_6110,N_6210);
nor U6707 (N_6707,N_6164,N_6048);
nor U6708 (N_6708,N_6264,N_6015);
and U6709 (N_6709,N_6416,N_6364);
or U6710 (N_6710,N_6427,N_6356);
nand U6711 (N_6711,N_6368,N_6202);
or U6712 (N_6712,N_6016,N_6354);
nor U6713 (N_6713,N_6013,N_6471);
nand U6714 (N_6714,N_6027,N_6434);
and U6715 (N_6715,N_6375,N_6067);
or U6716 (N_6716,N_6050,N_6087);
nand U6717 (N_6717,N_6437,N_6328);
or U6718 (N_6718,N_6041,N_6019);
or U6719 (N_6719,N_6432,N_6252);
nand U6720 (N_6720,N_6282,N_6435);
and U6721 (N_6721,N_6247,N_6095);
nor U6722 (N_6722,N_6301,N_6414);
or U6723 (N_6723,N_6064,N_6069);
or U6724 (N_6724,N_6309,N_6418);
and U6725 (N_6725,N_6467,N_6269);
nor U6726 (N_6726,N_6381,N_6073);
or U6727 (N_6727,N_6318,N_6385);
and U6728 (N_6728,N_6495,N_6294);
nor U6729 (N_6729,N_6438,N_6235);
nand U6730 (N_6730,N_6007,N_6313);
nand U6731 (N_6731,N_6052,N_6123);
nor U6732 (N_6732,N_6185,N_6401);
nor U6733 (N_6733,N_6441,N_6096);
or U6734 (N_6734,N_6237,N_6316);
and U6735 (N_6735,N_6293,N_6392);
nor U6736 (N_6736,N_6421,N_6424);
or U6737 (N_6737,N_6317,N_6369);
nor U6738 (N_6738,N_6429,N_6246);
nand U6739 (N_6739,N_6397,N_6436);
or U6740 (N_6740,N_6214,N_6183);
and U6741 (N_6741,N_6485,N_6378);
nor U6742 (N_6742,N_6077,N_6303);
or U6743 (N_6743,N_6078,N_6330);
and U6744 (N_6744,N_6192,N_6365);
and U6745 (N_6745,N_6253,N_6119);
or U6746 (N_6746,N_6104,N_6028);
or U6747 (N_6747,N_6349,N_6398);
or U6748 (N_6748,N_6280,N_6321);
nand U6749 (N_6749,N_6259,N_6174);
and U6750 (N_6750,N_6216,N_6416);
nor U6751 (N_6751,N_6176,N_6162);
nand U6752 (N_6752,N_6324,N_6394);
and U6753 (N_6753,N_6355,N_6205);
or U6754 (N_6754,N_6449,N_6034);
and U6755 (N_6755,N_6240,N_6019);
nand U6756 (N_6756,N_6217,N_6224);
and U6757 (N_6757,N_6033,N_6410);
nand U6758 (N_6758,N_6486,N_6289);
nor U6759 (N_6759,N_6203,N_6463);
and U6760 (N_6760,N_6336,N_6314);
or U6761 (N_6761,N_6222,N_6432);
nor U6762 (N_6762,N_6085,N_6064);
or U6763 (N_6763,N_6003,N_6343);
and U6764 (N_6764,N_6057,N_6081);
nor U6765 (N_6765,N_6043,N_6362);
nand U6766 (N_6766,N_6088,N_6169);
nor U6767 (N_6767,N_6065,N_6281);
and U6768 (N_6768,N_6429,N_6187);
nor U6769 (N_6769,N_6194,N_6145);
nand U6770 (N_6770,N_6257,N_6163);
and U6771 (N_6771,N_6260,N_6159);
nor U6772 (N_6772,N_6435,N_6029);
nand U6773 (N_6773,N_6477,N_6350);
nor U6774 (N_6774,N_6010,N_6066);
nor U6775 (N_6775,N_6298,N_6027);
or U6776 (N_6776,N_6192,N_6220);
and U6777 (N_6777,N_6478,N_6178);
nand U6778 (N_6778,N_6234,N_6468);
nor U6779 (N_6779,N_6076,N_6455);
or U6780 (N_6780,N_6133,N_6056);
or U6781 (N_6781,N_6336,N_6148);
or U6782 (N_6782,N_6362,N_6162);
or U6783 (N_6783,N_6453,N_6395);
nand U6784 (N_6784,N_6469,N_6427);
and U6785 (N_6785,N_6146,N_6339);
nor U6786 (N_6786,N_6128,N_6199);
nand U6787 (N_6787,N_6172,N_6358);
and U6788 (N_6788,N_6362,N_6012);
nor U6789 (N_6789,N_6123,N_6027);
nor U6790 (N_6790,N_6338,N_6109);
or U6791 (N_6791,N_6181,N_6077);
nor U6792 (N_6792,N_6312,N_6260);
nor U6793 (N_6793,N_6257,N_6203);
or U6794 (N_6794,N_6127,N_6354);
and U6795 (N_6795,N_6425,N_6012);
nor U6796 (N_6796,N_6400,N_6161);
nand U6797 (N_6797,N_6058,N_6065);
and U6798 (N_6798,N_6461,N_6281);
and U6799 (N_6799,N_6149,N_6415);
or U6800 (N_6800,N_6499,N_6225);
and U6801 (N_6801,N_6452,N_6368);
and U6802 (N_6802,N_6059,N_6342);
and U6803 (N_6803,N_6451,N_6142);
or U6804 (N_6804,N_6396,N_6235);
or U6805 (N_6805,N_6399,N_6448);
nor U6806 (N_6806,N_6139,N_6483);
and U6807 (N_6807,N_6195,N_6307);
nor U6808 (N_6808,N_6482,N_6275);
nor U6809 (N_6809,N_6346,N_6312);
nand U6810 (N_6810,N_6468,N_6121);
and U6811 (N_6811,N_6459,N_6375);
or U6812 (N_6812,N_6439,N_6378);
nor U6813 (N_6813,N_6094,N_6382);
or U6814 (N_6814,N_6370,N_6272);
and U6815 (N_6815,N_6240,N_6094);
nand U6816 (N_6816,N_6371,N_6106);
nor U6817 (N_6817,N_6419,N_6123);
and U6818 (N_6818,N_6267,N_6151);
or U6819 (N_6819,N_6273,N_6422);
nand U6820 (N_6820,N_6456,N_6113);
and U6821 (N_6821,N_6399,N_6031);
and U6822 (N_6822,N_6314,N_6416);
or U6823 (N_6823,N_6487,N_6119);
and U6824 (N_6824,N_6131,N_6460);
or U6825 (N_6825,N_6487,N_6328);
or U6826 (N_6826,N_6415,N_6245);
nand U6827 (N_6827,N_6448,N_6133);
or U6828 (N_6828,N_6265,N_6433);
nor U6829 (N_6829,N_6144,N_6058);
or U6830 (N_6830,N_6013,N_6088);
or U6831 (N_6831,N_6385,N_6317);
or U6832 (N_6832,N_6427,N_6022);
nand U6833 (N_6833,N_6258,N_6229);
and U6834 (N_6834,N_6002,N_6174);
or U6835 (N_6835,N_6209,N_6113);
nand U6836 (N_6836,N_6439,N_6078);
nand U6837 (N_6837,N_6193,N_6406);
nor U6838 (N_6838,N_6389,N_6471);
nand U6839 (N_6839,N_6209,N_6420);
nor U6840 (N_6840,N_6359,N_6338);
or U6841 (N_6841,N_6280,N_6345);
nor U6842 (N_6842,N_6065,N_6294);
nor U6843 (N_6843,N_6254,N_6216);
and U6844 (N_6844,N_6406,N_6196);
and U6845 (N_6845,N_6177,N_6247);
nand U6846 (N_6846,N_6068,N_6263);
nand U6847 (N_6847,N_6437,N_6057);
nand U6848 (N_6848,N_6287,N_6011);
or U6849 (N_6849,N_6017,N_6266);
and U6850 (N_6850,N_6115,N_6455);
and U6851 (N_6851,N_6138,N_6080);
nand U6852 (N_6852,N_6107,N_6206);
or U6853 (N_6853,N_6167,N_6132);
nand U6854 (N_6854,N_6426,N_6316);
nor U6855 (N_6855,N_6347,N_6420);
nor U6856 (N_6856,N_6252,N_6140);
and U6857 (N_6857,N_6249,N_6049);
and U6858 (N_6858,N_6318,N_6252);
or U6859 (N_6859,N_6350,N_6370);
nand U6860 (N_6860,N_6062,N_6235);
and U6861 (N_6861,N_6387,N_6331);
and U6862 (N_6862,N_6414,N_6027);
and U6863 (N_6863,N_6063,N_6395);
or U6864 (N_6864,N_6490,N_6302);
or U6865 (N_6865,N_6372,N_6031);
and U6866 (N_6866,N_6117,N_6018);
or U6867 (N_6867,N_6054,N_6382);
or U6868 (N_6868,N_6044,N_6048);
nor U6869 (N_6869,N_6036,N_6184);
nand U6870 (N_6870,N_6497,N_6219);
nor U6871 (N_6871,N_6359,N_6185);
and U6872 (N_6872,N_6363,N_6220);
or U6873 (N_6873,N_6447,N_6104);
or U6874 (N_6874,N_6020,N_6356);
nand U6875 (N_6875,N_6310,N_6350);
nand U6876 (N_6876,N_6412,N_6064);
and U6877 (N_6877,N_6421,N_6354);
nand U6878 (N_6878,N_6140,N_6277);
and U6879 (N_6879,N_6447,N_6197);
nand U6880 (N_6880,N_6270,N_6378);
nor U6881 (N_6881,N_6437,N_6269);
nand U6882 (N_6882,N_6047,N_6311);
nand U6883 (N_6883,N_6087,N_6151);
nor U6884 (N_6884,N_6346,N_6238);
or U6885 (N_6885,N_6121,N_6159);
and U6886 (N_6886,N_6198,N_6476);
nor U6887 (N_6887,N_6424,N_6097);
nor U6888 (N_6888,N_6231,N_6244);
xnor U6889 (N_6889,N_6451,N_6495);
and U6890 (N_6890,N_6223,N_6285);
nand U6891 (N_6891,N_6115,N_6434);
nand U6892 (N_6892,N_6445,N_6296);
or U6893 (N_6893,N_6357,N_6178);
nand U6894 (N_6894,N_6271,N_6354);
and U6895 (N_6895,N_6345,N_6073);
and U6896 (N_6896,N_6376,N_6365);
and U6897 (N_6897,N_6454,N_6152);
and U6898 (N_6898,N_6359,N_6323);
or U6899 (N_6899,N_6467,N_6172);
nor U6900 (N_6900,N_6116,N_6214);
or U6901 (N_6901,N_6081,N_6084);
nor U6902 (N_6902,N_6416,N_6301);
or U6903 (N_6903,N_6453,N_6150);
or U6904 (N_6904,N_6109,N_6386);
nor U6905 (N_6905,N_6414,N_6133);
or U6906 (N_6906,N_6152,N_6274);
and U6907 (N_6907,N_6157,N_6331);
and U6908 (N_6908,N_6019,N_6183);
or U6909 (N_6909,N_6176,N_6151);
and U6910 (N_6910,N_6321,N_6167);
or U6911 (N_6911,N_6323,N_6235);
nand U6912 (N_6912,N_6296,N_6240);
nor U6913 (N_6913,N_6359,N_6043);
and U6914 (N_6914,N_6211,N_6496);
and U6915 (N_6915,N_6128,N_6118);
nor U6916 (N_6916,N_6193,N_6458);
nand U6917 (N_6917,N_6381,N_6472);
and U6918 (N_6918,N_6247,N_6468);
nand U6919 (N_6919,N_6334,N_6347);
and U6920 (N_6920,N_6296,N_6178);
nor U6921 (N_6921,N_6173,N_6393);
or U6922 (N_6922,N_6499,N_6179);
nand U6923 (N_6923,N_6040,N_6100);
and U6924 (N_6924,N_6001,N_6394);
nand U6925 (N_6925,N_6422,N_6155);
or U6926 (N_6926,N_6318,N_6448);
nor U6927 (N_6927,N_6134,N_6275);
nor U6928 (N_6928,N_6112,N_6240);
and U6929 (N_6929,N_6125,N_6195);
and U6930 (N_6930,N_6419,N_6204);
nor U6931 (N_6931,N_6491,N_6354);
xnor U6932 (N_6932,N_6336,N_6015);
nor U6933 (N_6933,N_6088,N_6463);
nor U6934 (N_6934,N_6336,N_6498);
nor U6935 (N_6935,N_6256,N_6426);
or U6936 (N_6936,N_6374,N_6433);
nor U6937 (N_6937,N_6363,N_6387);
and U6938 (N_6938,N_6165,N_6001);
or U6939 (N_6939,N_6013,N_6260);
nor U6940 (N_6940,N_6470,N_6259);
nor U6941 (N_6941,N_6434,N_6017);
nand U6942 (N_6942,N_6273,N_6377);
nand U6943 (N_6943,N_6053,N_6083);
nor U6944 (N_6944,N_6223,N_6369);
and U6945 (N_6945,N_6413,N_6074);
nor U6946 (N_6946,N_6188,N_6002);
nor U6947 (N_6947,N_6126,N_6449);
and U6948 (N_6948,N_6128,N_6358);
and U6949 (N_6949,N_6175,N_6260);
and U6950 (N_6950,N_6184,N_6261);
and U6951 (N_6951,N_6402,N_6131);
nor U6952 (N_6952,N_6071,N_6348);
or U6953 (N_6953,N_6214,N_6179);
nor U6954 (N_6954,N_6259,N_6274);
nor U6955 (N_6955,N_6087,N_6367);
or U6956 (N_6956,N_6052,N_6148);
nand U6957 (N_6957,N_6383,N_6018);
or U6958 (N_6958,N_6267,N_6087);
xor U6959 (N_6959,N_6373,N_6495);
or U6960 (N_6960,N_6499,N_6251);
nor U6961 (N_6961,N_6474,N_6390);
nor U6962 (N_6962,N_6051,N_6205);
xnor U6963 (N_6963,N_6128,N_6077);
nand U6964 (N_6964,N_6421,N_6241);
nor U6965 (N_6965,N_6048,N_6330);
and U6966 (N_6966,N_6231,N_6260);
and U6967 (N_6967,N_6383,N_6028);
nor U6968 (N_6968,N_6070,N_6129);
or U6969 (N_6969,N_6122,N_6026);
nor U6970 (N_6970,N_6367,N_6239);
nand U6971 (N_6971,N_6083,N_6450);
or U6972 (N_6972,N_6200,N_6421);
or U6973 (N_6973,N_6218,N_6499);
and U6974 (N_6974,N_6111,N_6017);
nor U6975 (N_6975,N_6460,N_6426);
nor U6976 (N_6976,N_6437,N_6039);
nand U6977 (N_6977,N_6100,N_6018);
nor U6978 (N_6978,N_6004,N_6236);
nand U6979 (N_6979,N_6448,N_6108);
or U6980 (N_6980,N_6411,N_6033);
nor U6981 (N_6981,N_6165,N_6337);
and U6982 (N_6982,N_6031,N_6094);
nor U6983 (N_6983,N_6048,N_6368);
or U6984 (N_6984,N_6399,N_6419);
or U6985 (N_6985,N_6094,N_6004);
or U6986 (N_6986,N_6081,N_6056);
and U6987 (N_6987,N_6334,N_6378);
and U6988 (N_6988,N_6035,N_6231);
and U6989 (N_6989,N_6035,N_6311);
or U6990 (N_6990,N_6096,N_6125);
and U6991 (N_6991,N_6123,N_6071);
or U6992 (N_6992,N_6276,N_6330);
nand U6993 (N_6993,N_6487,N_6163);
nor U6994 (N_6994,N_6294,N_6370);
nor U6995 (N_6995,N_6327,N_6441);
and U6996 (N_6996,N_6056,N_6228);
and U6997 (N_6997,N_6459,N_6159);
nand U6998 (N_6998,N_6187,N_6346);
xor U6999 (N_6999,N_6425,N_6190);
xnor U7000 (N_7000,N_6979,N_6832);
nor U7001 (N_7001,N_6947,N_6790);
nor U7002 (N_7002,N_6758,N_6848);
or U7003 (N_7003,N_6558,N_6925);
and U7004 (N_7004,N_6918,N_6683);
nand U7005 (N_7005,N_6567,N_6696);
and U7006 (N_7006,N_6762,N_6958);
or U7007 (N_7007,N_6616,N_6873);
nor U7008 (N_7008,N_6955,N_6736);
nand U7009 (N_7009,N_6662,N_6807);
or U7010 (N_7010,N_6936,N_6812);
nand U7011 (N_7011,N_6928,N_6811);
or U7012 (N_7012,N_6859,N_6634);
nand U7013 (N_7013,N_6959,N_6682);
nor U7014 (N_7014,N_6760,N_6954);
nand U7015 (N_7015,N_6734,N_6822);
and U7016 (N_7016,N_6923,N_6883);
nor U7017 (N_7017,N_6720,N_6524);
and U7018 (N_7018,N_6797,N_6861);
nor U7019 (N_7019,N_6920,N_6769);
or U7020 (N_7020,N_6863,N_6519);
nand U7021 (N_7021,N_6713,N_6772);
or U7022 (N_7022,N_6669,N_6689);
or U7023 (N_7023,N_6660,N_6602);
nor U7024 (N_7024,N_6818,N_6678);
or U7025 (N_7025,N_6628,N_6658);
or U7026 (N_7026,N_6515,N_6903);
and U7027 (N_7027,N_6949,N_6606);
nand U7028 (N_7028,N_6703,N_6901);
nand U7029 (N_7029,N_6562,N_6640);
and U7030 (N_7030,N_6874,N_6864);
and U7031 (N_7031,N_6555,N_6625);
nor U7032 (N_7032,N_6598,N_6526);
or U7033 (N_7033,N_6648,N_6950);
and U7034 (N_7034,N_6902,N_6897);
or U7035 (N_7035,N_6730,N_6907);
nor U7036 (N_7036,N_6846,N_6857);
or U7037 (N_7037,N_6610,N_6878);
and U7038 (N_7038,N_6595,N_6913);
nand U7039 (N_7039,N_6745,N_6800);
or U7040 (N_7040,N_6829,N_6547);
nor U7041 (N_7041,N_6666,N_6589);
and U7042 (N_7042,N_6796,N_6803);
nand U7043 (N_7043,N_6639,N_6718);
and U7044 (N_7044,N_6989,N_6621);
nand U7045 (N_7045,N_6935,N_6953);
or U7046 (N_7046,N_6617,N_6981);
nand U7047 (N_7047,N_6716,N_6728);
nand U7048 (N_7048,N_6768,N_6824);
or U7049 (N_7049,N_6850,N_6862);
nor U7050 (N_7050,N_6914,N_6688);
nand U7051 (N_7051,N_6732,N_6675);
or U7052 (N_7052,N_6929,N_6997);
and U7053 (N_7053,N_6564,N_6853);
nor U7054 (N_7054,N_6527,N_6536);
nor U7055 (N_7055,N_6637,N_6826);
or U7056 (N_7056,N_6709,N_6927);
or U7057 (N_7057,N_6744,N_6554);
and U7058 (N_7058,N_6847,N_6717);
and U7059 (N_7059,N_6712,N_6990);
nor U7060 (N_7060,N_6723,N_6851);
or U7061 (N_7061,N_6646,N_6512);
nor U7062 (N_7062,N_6719,N_6983);
nand U7063 (N_7063,N_6804,N_6722);
or U7064 (N_7064,N_6557,N_6521);
and U7065 (N_7065,N_6691,N_6529);
nor U7066 (N_7066,N_6692,N_6571);
nand U7067 (N_7067,N_6684,N_6892);
or U7068 (N_7068,N_6965,N_6600);
and U7069 (N_7069,N_6503,N_6507);
or U7070 (N_7070,N_6697,N_6568);
nand U7071 (N_7071,N_6542,N_6885);
nor U7072 (N_7072,N_6938,N_6500);
or U7073 (N_7073,N_6694,N_6566);
nor U7074 (N_7074,N_6619,N_6698);
or U7075 (N_7075,N_6548,N_6575);
and U7076 (N_7076,N_6932,N_6624);
and U7077 (N_7077,N_6517,N_6916);
and U7078 (N_7078,N_6887,N_6773);
nor U7079 (N_7079,N_6974,N_6771);
nand U7080 (N_7080,N_6942,N_6855);
nor U7081 (N_7081,N_6944,N_6594);
nor U7082 (N_7082,N_6502,N_6633);
or U7083 (N_7083,N_6978,N_6603);
nand U7084 (N_7084,N_6948,N_6565);
xor U7085 (N_7085,N_6592,N_6805);
or U7086 (N_7086,N_6614,N_6680);
and U7087 (N_7087,N_6879,N_6827);
or U7088 (N_7088,N_6733,N_6881);
and U7089 (N_7089,N_6747,N_6577);
nand U7090 (N_7090,N_6886,N_6963);
nand U7091 (N_7091,N_6560,N_6995);
and U7092 (N_7092,N_6875,N_6764);
nand U7093 (N_7093,N_6608,N_6842);
xnor U7094 (N_7094,N_6641,N_6952);
nor U7095 (N_7095,N_6817,N_6657);
or U7096 (N_7096,N_6534,N_6806);
or U7097 (N_7097,N_6638,N_6748);
and U7098 (N_7098,N_6630,N_6900);
and U7099 (N_7099,N_6582,N_6686);
and U7100 (N_7100,N_6996,N_6821);
or U7101 (N_7101,N_6854,N_6946);
nor U7102 (N_7102,N_6700,N_6998);
nor U7103 (N_7103,N_6843,N_6810);
or U7104 (N_7104,N_6750,N_6869);
or U7105 (N_7105,N_6945,N_6729);
or U7106 (N_7106,N_6917,N_6731);
or U7107 (N_7107,N_6553,N_6654);
and U7108 (N_7108,N_6931,N_6971);
nand U7109 (N_7109,N_6994,N_6967);
nand U7110 (N_7110,N_6735,N_6746);
nor U7111 (N_7111,N_6975,N_6535);
nand U7112 (N_7112,N_6739,N_6743);
nor U7113 (N_7113,N_6871,N_6708);
and U7114 (N_7114,N_6926,N_6834);
nor U7115 (N_7115,N_6627,N_6649);
xor U7116 (N_7116,N_6540,N_6710);
or U7117 (N_7117,N_6985,N_6973);
nand U7118 (N_7118,N_6636,N_6899);
and U7119 (N_7119,N_6752,N_6693);
nand U7120 (N_7120,N_6763,N_6702);
nand U7121 (N_7121,N_6581,N_6599);
nor U7122 (N_7122,N_6813,N_6960);
nor U7123 (N_7123,N_6652,N_6791);
and U7124 (N_7124,N_6650,N_6820);
nand U7125 (N_7125,N_6801,N_6623);
nand U7126 (N_7126,N_6551,N_6705);
nand U7127 (N_7127,N_6673,N_6992);
nand U7128 (N_7128,N_6586,N_6856);
nand U7129 (N_7129,N_6741,N_6968);
nor U7130 (N_7130,N_6596,N_6611);
nand U7131 (N_7131,N_6583,N_6844);
or U7132 (N_7132,N_6543,N_6756);
nand U7133 (N_7133,N_6877,N_6999);
or U7134 (N_7134,N_6780,N_6908);
nor U7135 (N_7135,N_6607,N_6792);
or U7136 (N_7136,N_6546,N_6837);
or U7137 (N_7137,N_6569,N_6742);
nor U7138 (N_7138,N_6645,N_6738);
and U7139 (N_7139,N_6831,N_6776);
or U7140 (N_7140,N_6852,N_6580);
nor U7141 (N_7141,N_6632,N_6839);
xnor U7142 (N_7142,N_6778,N_6563);
and U7143 (N_7143,N_6766,N_6940);
xor U7144 (N_7144,N_6685,N_6518);
nor U7145 (N_7145,N_6911,N_6905);
nor U7146 (N_7146,N_6721,N_6622);
and U7147 (N_7147,N_6891,N_6681);
nand U7148 (N_7148,N_6511,N_6514);
nand U7149 (N_7149,N_6751,N_6795);
nor U7150 (N_7150,N_6798,N_6501);
xnor U7151 (N_7151,N_6601,N_6819);
nor U7152 (N_7152,N_6690,N_6612);
and U7153 (N_7153,N_6987,N_6860);
and U7154 (N_7154,N_6777,N_6643);
or U7155 (N_7155,N_6814,N_6532);
nand U7156 (N_7156,N_6970,N_6591);
nand U7157 (N_7157,N_6510,N_6604);
nand U7158 (N_7158,N_6951,N_6865);
nand U7159 (N_7159,N_6613,N_6588);
or U7160 (N_7160,N_6525,N_6513);
nand U7161 (N_7161,N_6508,N_6921);
nand U7162 (N_7162,N_6695,N_6677);
nor U7163 (N_7163,N_6786,N_6833);
and U7164 (N_7164,N_6725,N_6784);
or U7165 (N_7165,N_6670,N_6785);
xor U7166 (N_7166,N_6753,N_6642);
nand U7167 (N_7167,N_6870,N_6964);
or U7168 (N_7168,N_6726,N_6969);
xor U7169 (N_7169,N_6934,N_6808);
or U7170 (N_7170,N_6727,N_6620);
and U7171 (N_7171,N_6664,N_6505);
nand U7172 (N_7172,N_6961,N_6896);
or U7173 (N_7173,N_6788,N_6941);
or U7174 (N_7174,N_6816,N_6815);
nor U7175 (N_7175,N_6782,N_6962);
or U7176 (N_7176,N_6523,N_6605);
nand U7177 (N_7177,N_6982,N_6561);
nor U7178 (N_7178,N_6520,N_6531);
nand U7179 (N_7179,N_6930,N_6674);
and U7180 (N_7180,N_6889,N_6779);
or U7181 (N_7181,N_6898,N_6794);
or U7182 (N_7182,N_6590,N_6706);
or U7183 (N_7183,N_6656,N_6754);
nand U7184 (N_7184,N_6858,N_6615);
and U7185 (N_7185,N_6574,N_6789);
nand U7186 (N_7186,N_6749,N_6597);
and U7187 (N_7187,N_6809,N_6910);
and U7188 (N_7188,N_6894,N_6919);
nand U7189 (N_7189,N_6825,N_6609);
nand U7190 (N_7190,N_6522,N_6665);
nand U7191 (N_7191,N_6909,N_6579);
nand U7192 (N_7192,N_6823,N_6872);
and U7193 (N_7193,N_6667,N_6631);
nand U7194 (N_7194,N_6537,N_6545);
nor U7195 (N_7195,N_6912,N_6986);
or U7196 (N_7196,N_6933,N_6701);
nor U7197 (N_7197,N_6552,N_6504);
or U7198 (N_7198,N_6761,N_6585);
and U7199 (N_7199,N_6679,N_6849);
and U7200 (N_7200,N_6573,N_6714);
or U7201 (N_7201,N_6802,N_6774);
and U7202 (N_7202,N_6980,N_6539);
and U7203 (N_7203,N_6939,N_6549);
or U7204 (N_7204,N_6893,N_6976);
nor U7205 (N_7205,N_6770,N_6687);
or U7206 (N_7206,N_6704,N_6880);
nand U7207 (N_7207,N_6966,N_6830);
nor U7208 (N_7208,N_6991,N_6924);
nor U7209 (N_7209,N_6836,N_6506);
and U7210 (N_7210,N_6676,N_6828);
nor U7211 (N_7211,N_6943,N_6626);
nand U7212 (N_7212,N_6559,N_6570);
nor U7213 (N_7213,N_6724,N_6867);
nand U7214 (N_7214,N_6841,N_6799);
nor U7215 (N_7215,N_6707,N_6882);
and U7216 (N_7216,N_6988,N_6644);
nor U7217 (N_7217,N_6765,N_6906);
or U7218 (N_7218,N_6576,N_6578);
and U7219 (N_7219,N_6544,N_6516);
nor U7220 (N_7220,N_6835,N_6671);
nand U7221 (N_7221,N_6651,N_6866);
nor U7222 (N_7222,N_6572,N_6584);
nand U7223 (N_7223,N_6533,N_6538);
and U7224 (N_7224,N_6775,N_6740);
or U7225 (N_7225,N_6647,N_6838);
or U7226 (N_7226,N_6618,N_6890);
xor U7227 (N_7227,N_6972,N_6840);
nor U7228 (N_7228,N_6783,N_6793);
nor U7229 (N_7229,N_6757,N_6876);
nor U7230 (N_7230,N_6755,N_6884);
or U7231 (N_7231,N_6629,N_6845);
xnor U7232 (N_7232,N_6984,N_6977);
and U7233 (N_7233,N_6668,N_6937);
or U7234 (N_7234,N_6956,N_6767);
and U7235 (N_7235,N_6655,N_6993);
nand U7236 (N_7236,N_6663,N_6895);
nand U7237 (N_7237,N_6787,N_6550);
nand U7238 (N_7238,N_6759,N_6593);
nand U7239 (N_7239,N_6672,N_6587);
nand U7240 (N_7240,N_6509,N_6556);
and U7241 (N_7241,N_6922,N_6737);
or U7242 (N_7242,N_6699,N_6868);
nor U7243 (N_7243,N_6781,N_6635);
nand U7244 (N_7244,N_6528,N_6653);
nor U7245 (N_7245,N_6530,N_6659);
nor U7246 (N_7246,N_6957,N_6711);
nor U7247 (N_7247,N_6915,N_6904);
or U7248 (N_7248,N_6661,N_6888);
nor U7249 (N_7249,N_6541,N_6715);
and U7250 (N_7250,N_6638,N_6829);
or U7251 (N_7251,N_6814,N_6889);
nor U7252 (N_7252,N_6676,N_6829);
and U7253 (N_7253,N_6884,N_6623);
nor U7254 (N_7254,N_6678,N_6789);
nand U7255 (N_7255,N_6900,N_6906);
and U7256 (N_7256,N_6865,N_6756);
nor U7257 (N_7257,N_6762,N_6765);
or U7258 (N_7258,N_6753,N_6532);
xnor U7259 (N_7259,N_6530,N_6700);
xor U7260 (N_7260,N_6500,N_6583);
nor U7261 (N_7261,N_6797,N_6780);
nand U7262 (N_7262,N_6938,N_6727);
and U7263 (N_7263,N_6515,N_6616);
nor U7264 (N_7264,N_6649,N_6994);
and U7265 (N_7265,N_6787,N_6577);
nor U7266 (N_7266,N_6524,N_6801);
nor U7267 (N_7267,N_6629,N_6729);
and U7268 (N_7268,N_6943,N_6717);
or U7269 (N_7269,N_6698,N_6571);
nand U7270 (N_7270,N_6637,N_6729);
and U7271 (N_7271,N_6842,N_6703);
or U7272 (N_7272,N_6771,N_6941);
nand U7273 (N_7273,N_6652,N_6742);
xor U7274 (N_7274,N_6807,N_6981);
and U7275 (N_7275,N_6720,N_6897);
nor U7276 (N_7276,N_6815,N_6568);
and U7277 (N_7277,N_6842,N_6668);
and U7278 (N_7278,N_6943,N_6990);
and U7279 (N_7279,N_6883,N_6954);
nand U7280 (N_7280,N_6509,N_6726);
nor U7281 (N_7281,N_6755,N_6885);
nor U7282 (N_7282,N_6820,N_6808);
and U7283 (N_7283,N_6973,N_6537);
or U7284 (N_7284,N_6952,N_6670);
nand U7285 (N_7285,N_6998,N_6564);
and U7286 (N_7286,N_6684,N_6592);
nor U7287 (N_7287,N_6860,N_6901);
or U7288 (N_7288,N_6537,N_6847);
nand U7289 (N_7289,N_6640,N_6661);
nand U7290 (N_7290,N_6895,N_6774);
nand U7291 (N_7291,N_6803,N_6833);
and U7292 (N_7292,N_6622,N_6586);
nor U7293 (N_7293,N_6835,N_6813);
and U7294 (N_7294,N_6808,N_6960);
nand U7295 (N_7295,N_6975,N_6902);
nor U7296 (N_7296,N_6555,N_6806);
nand U7297 (N_7297,N_6638,N_6605);
nor U7298 (N_7298,N_6540,N_6582);
or U7299 (N_7299,N_6592,N_6873);
nor U7300 (N_7300,N_6863,N_6853);
xor U7301 (N_7301,N_6738,N_6777);
nand U7302 (N_7302,N_6692,N_6687);
nor U7303 (N_7303,N_6552,N_6963);
nand U7304 (N_7304,N_6882,N_6504);
or U7305 (N_7305,N_6834,N_6745);
or U7306 (N_7306,N_6850,N_6776);
and U7307 (N_7307,N_6516,N_6865);
or U7308 (N_7308,N_6809,N_6770);
nor U7309 (N_7309,N_6791,N_6825);
or U7310 (N_7310,N_6812,N_6814);
or U7311 (N_7311,N_6862,N_6986);
or U7312 (N_7312,N_6964,N_6914);
nor U7313 (N_7313,N_6665,N_6687);
nand U7314 (N_7314,N_6701,N_6842);
nand U7315 (N_7315,N_6549,N_6742);
nand U7316 (N_7316,N_6569,N_6706);
nor U7317 (N_7317,N_6600,N_6817);
nand U7318 (N_7318,N_6725,N_6645);
nor U7319 (N_7319,N_6829,N_6533);
nand U7320 (N_7320,N_6800,N_6933);
and U7321 (N_7321,N_6563,N_6989);
xor U7322 (N_7322,N_6701,N_6814);
nand U7323 (N_7323,N_6956,N_6781);
or U7324 (N_7324,N_6615,N_6643);
xnor U7325 (N_7325,N_6990,N_6573);
and U7326 (N_7326,N_6931,N_6669);
nand U7327 (N_7327,N_6632,N_6515);
or U7328 (N_7328,N_6581,N_6537);
nor U7329 (N_7329,N_6654,N_6843);
and U7330 (N_7330,N_6742,N_6883);
and U7331 (N_7331,N_6670,N_6595);
xnor U7332 (N_7332,N_6505,N_6902);
and U7333 (N_7333,N_6770,N_6778);
and U7334 (N_7334,N_6831,N_6521);
nand U7335 (N_7335,N_6989,N_6513);
and U7336 (N_7336,N_6578,N_6638);
nand U7337 (N_7337,N_6911,N_6818);
and U7338 (N_7338,N_6717,N_6757);
and U7339 (N_7339,N_6698,N_6992);
and U7340 (N_7340,N_6999,N_6652);
nand U7341 (N_7341,N_6831,N_6993);
nand U7342 (N_7342,N_6799,N_6539);
nand U7343 (N_7343,N_6978,N_6901);
nand U7344 (N_7344,N_6606,N_6813);
nand U7345 (N_7345,N_6508,N_6981);
and U7346 (N_7346,N_6569,N_6841);
or U7347 (N_7347,N_6816,N_6869);
and U7348 (N_7348,N_6504,N_6836);
nand U7349 (N_7349,N_6774,N_6797);
xnor U7350 (N_7350,N_6762,N_6882);
nand U7351 (N_7351,N_6869,N_6878);
nor U7352 (N_7352,N_6578,N_6542);
or U7353 (N_7353,N_6642,N_6999);
and U7354 (N_7354,N_6543,N_6524);
and U7355 (N_7355,N_6794,N_6736);
nor U7356 (N_7356,N_6589,N_6625);
and U7357 (N_7357,N_6671,N_6946);
nand U7358 (N_7358,N_6874,N_6541);
or U7359 (N_7359,N_6511,N_6521);
nor U7360 (N_7360,N_6828,N_6885);
and U7361 (N_7361,N_6605,N_6573);
and U7362 (N_7362,N_6524,N_6530);
or U7363 (N_7363,N_6928,N_6800);
or U7364 (N_7364,N_6975,N_6642);
or U7365 (N_7365,N_6550,N_6726);
and U7366 (N_7366,N_6809,N_6564);
nor U7367 (N_7367,N_6727,N_6973);
and U7368 (N_7368,N_6551,N_6718);
nor U7369 (N_7369,N_6638,N_6903);
nand U7370 (N_7370,N_6865,N_6947);
nor U7371 (N_7371,N_6903,N_6588);
nand U7372 (N_7372,N_6786,N_6696);
nor U7373 (N_7373,N_6668,N_6899);
xnor U7374 (N_7374,N_6939,N_6999);
nor U7375 (N_7375,N_6569,N_6991);
and U7376 (N_7376,N_6667,N_6687);
nand U7377 (N_7377,N_6655,N_6748);
nor U7378 (N_7378,N_6778,N_6693);
or U7379 (N_7379,N_6857,N_6866);
nor U7380 (N_7380,N_6671,N_6821);
and U7381 (N_7381,N_6906,N_6595);
nor U7382 (N_7382,N_6584,N_6592);
or U7383 (N_7383,N_6978,N_6713);
nand U7384 (N_7384,N_6884,N_6998);
nor U7385 (N_7385,N_6885,N_6780);
and U7386 (N_7386,N_6986,N_6678);
and U7387 (N_7387,N_6703,N_6857);
or U7388 (N_7388,N_6628,N_6669);
or U7389 (N_7389,N_6635,N_6923);
and U7390 (N_7390,N_6996,N_6535);
or U7391 (N_7391,N_6937,N_6974);
nor U7392 (N_7392,N_6745,N_6824);
nand U7393 (N_7393,N_6738,N_6939);
nor U7394 (N_7394,N_6878,N_6786);
and U7395 (N_7395,N_6821,N_6550);
nand U7396 (N_7396,N_6769,N_6744);
or U7397 (N_7397,N_6754,N_6776);
and U7398 (N_7398,N_6561,N_6794);
nor U7399 (N_7399,N_6561,N_6886);
nand U7400 (N_7400,N_6622,N_6828);
and U7401 (N_7401,N_6934,N_6903);
or U7402 (N_7402,N_6632,N_6889);
nand U7403 (N_7403,N_6802,N_6922);
or U7404 (N_7404,N_6581,N_6937);
or U7405 (N_7405,N_6916,N_6774);
nor U7406 (N_7406,N_6984,N_6771);
and U7407 (N_7407,N_6554,N_6545);
nand U7408 (N_7408,N_6970,N_6837);
nand U7409 (N_7409,N_6931,N_6938);
and U7410 (N_7410,N_6836,N_6689);
or U7411 (N_7411,N_6852,N_6811);
nand U7412 (N_7412,N_6660,N_6649);
nand U7413 (N_7413,N_6560,N_6934);
and U7414 (N_7414,N_6590,N_6786);
or U7415 (N_7415,N_6663,N_6530);
nand U7416 (N_7416,N_6870,N_6875);
or U7417 (N_7417,N_6611,N_6913);
and U7418 (N_7418,N_6761,N_6764);
and U7419 (N_7419,N_6968,N_6936);
nand U7420 (N_7420,N_6737,N_6699);
nand U7421 (N_7421,N_6998,N_6864);
and U7422 (N_7422,N_6872,N_6819);
nor U7423 (N_7423,N_6969,N_6838);
nand U7424 (N_7424,N_6711,N_6632);
nand U7425 (N_7425,N_6562,N_6603);
or U7426 (N_7426,N_6523,N_6906);
and U7427 (N_7427,N_6645,N_6994);
or U7428 (N_7428,N_6608,N_6963);
nor U7429 (N_7429,N_6643,N_6560);
or U7430 (N_7430,N_6724,N_6984);
or U7431 (N_7431,N_6505,N_6731);
or U7432 (N_7432,N_6973,N_6524);
and U7433 (N_7433,N_6902,N_6827);
or U7434 (N_7434,N_6993,N_6551);
or U7435 (N_7435,N_6546,N_6988);
nand U7436 (N_7436,N_6679,N_6960);
or U7437 (N_7437,N_6691,N_6742);
nand U7438 (N_7438,N_6657,N_6722);
nand U7439 (N_7439,N_6941,N_6739);
or U7440 (N_7440,N_6851,N_6576);
nand U7441 (N_7441,N_6846,N_6580);
or U7442 (N_7442,N_6516,N_6810);
or U7443 (N_7443,N_6701,N_6557);
or U7444 (N_7444,N_6958,N_6766);
or U7445 (N_7445,N_6970,N_6923);
and U7446 (N_7446,N_6500,N_6630);
or U7447 (N_7447,N_6854,N_6515);
nor U7448 (N_7448,N_6836,N_6579);
nand U7449 (N_7449,N_6863,N_6897);
and U7450 (N_7450,N_6834,N_6596);
nand U7451 (N_7451,N_6734,N_6503);
and U7452 (N_7452,N_6968,N_6631);
nor U7453 (N_7453,N_6683,N_6604);
nand U7454 (N_7454,N_6519,N_6634);
and U7455 (N_7455,N_6538,N_6797);
or U7456 (N_7456,N_6614,N_6965);
or U7457 (N_7457,N_6811,N_6914);
nand U7458 (N_7458,N_6859,N_6947);
xor U7459 (N_7459,N_6732,N_6767);
nand U7460 (N_7460,N_6582,N_6861);
or U7461 (N_7461,N_6836,N_6745);
nor U7462 (N_7462,N_6777,N_6529);
and U7463 (N_7463,N_6861,N_6870);
nand U7464 (N_7464,N_6799,N_6631);
or U7465 (N_7465,N_6920,N_6529);
nor U7466 (N_7466,N_6553,N_6824);
nor U7467 (N_7467,N_6992,N_6665);
nand U7468 (N_7468,N_6565,N_6664);
and U7469 (N_7469,N_6528,N_6951);
or U7470 (N_7470,N_6857,N_6653);
xnor U7471 (N_7471,N_6769,N_6603);
or U7472 (N_7472,N_6937,N_6686);
or U7473 (N_7473,N_6929,N_6578);
and U7474 (N_7474,N_6773,N_6565);
or U7475 (N_7475,N_6821,N_6840);
nand U7476 (N_7476,N_6514,N_6640);
nand U7477 (N_7477,N_6709,N_6965);
nand U7478 (N_7478,N_6878,N_6887);
or U7479 (N_7479,N_6877,N_6685);
nand U7480 (N_7480,N_6892,N_6837);
nand U7481 (N_7481,N_6769,N_6655);
and U7482 (N_7482,N_6840,N_6841);
and U7483 (N_7483,N_6808,N_6857);
and U7484 (N_7484,N_6644,N_6791);
and U7485 (N_7485,N_6971,N_6930);
or U7486 (N_7486,N_6951,N_6568);
and U7487 (N_7487,N_6631,N_6875);
nand U7488 (N_7488,N_6606,N_6567);
and U7489 (N_7489,N_6628,N_6688);
nor U7490 (N_7490,N_6779,N_6950);
xnor U7491 (N_7491,N_6872,N_6616);
or U7492 (N_7492,N_6514,N_6510);
or U7493 (N_7493,N_6923,N_6638);
nor U7494 (N_7494,N_6892,N_6830);
nor U7495 (N_7495,N_6638,N_6960);
nand U7496 (N_7496,N_6907,N_6858);
nor U7497 (N_7497,N_6952,N_6844);
and U7498 (N_7498,N_6528,N_6650);
nand U7499 (N_7499,N_6656,N_6874);
and U7500 (N_7500,N_7329,N_7340);
or U7501 (N_7501,N_7062,N_7407);
nor U7502 (N_7502,N_7078,N_7045);
nor U7503 (N_7503,N_7082,N_7107);
nor U7504 (N_7504,N_7044,N_7497);
or U7505 (N_7505,N_7131,N_7008);
nor U7506 (N_7506,N_7305,N_7352);
nor U7507 (N_7507,N_7236,N_7475);
and U7508 (N_7508,N_7056,N_7255);
and U7509 (N_7509,N_7385,N_7128);
nor U7510 (N_7510,N_7126,N_7367);
and U7511 (N_7511,N_7054,N_7247);
or U7512 (N_7512,N_7351,N_7419);
nor U7513 (N_7513,N_7071,N_7046);
nand U7514 (N_7514,N_7271,N_7350);
nor U7515 (N_7515,N_7007,N_7444);
and U7516 (N_7516,N_7197,N_7389);
nand U7517 (N_7517,N_7499,N_7495);
or U7518 (N_7518,N_7343,N_7337);
and U7519 (N_7519,N_7482,N_7426);
nor U7520 (N_7520,N_7375,N_7339);
nor U7521 (N_7521,N_7153,N_7262);
nor U7522 (N_7522,N_7066,N_7167);
nor U7523 (N_7523,N_7098,N_7293);
or U7524 (N_7524,N_7383,N_7214);
nand U7525 (N_7525,N_7148,N_7109);
and U7526 (N_7526,N_7228,N_7021);
and U7527 (N_7527,N_7377,N_7278);
or U7528 (N_7528,N_7252,N_7015);
and U7529 (N_7529,N_7155,N_7381);
and U7530 (N_7530,N_7332,N_7422);
nand U7531 (N_7531,N_7326,N_7263);
or U7532 (N_7532,N_7286,N_7312);
or U7533 (N_7533,N_7276,N_7279);
or U7534 (N_7534,N_7466,N_7038);
or U7535 (N_7535,N_7403,N_7158);
or U7536 (N_7536,N_7074,N_7480);
or U7537 (N_7537,N_7069,N_7133);
nand U7538 (N_7538,N_7025,N_7485);
and U7539 (N_7539,N_7354,N_7244);
or U7540 (N_7540,N_7005,N_7017);
and U7541 (N_7541,N_7488,N_7462);
or U7542 (N_7542,N_7246,N_7171);
nor U7543 (N_7543,N_7111,N_7101);
nor U7544 (N_7544,N_7103,N_7321);
nor U7545 (N_7545,N_7446,N_7225);
and U7546 (N_7546,N_7392,N_7188);
and U7547 (N_7547,N_7484,N_7047);
xnor U7548 (N_7548,N_7260,N_7409);
and U7549 (N_7549,N_7489,N_7253);
or U7550 (N_7550,N_7130,N_7256);
or U7551 (N_7551,N_7215,N_7178);
and U7552 (N_7552,N_7308,N_7018);
nand U7553 (N_7553,N_7401,N_7478);
or U7554 (N_7554,N_7113,N_7006);
nor U7555 (N_7555,N_7146,N_7043);
nor U7556 (N_7556,N_7397,N_7053);
nor U7557 (N_7557,N_7134,N_7315);
or U7558 (N_7558,N_7299,N_7306);
nor U7559 (N_7559,N_7268,N_7145);
nand U7560 (N_7560,N_7075,N_7452);
nor U7561 (N_7561,N_7224,N_7487);
and U7562 (N_7562,N_7222,N_7122);
or U7563 (N_7563,N_7431,N_7492);
nor U7564 (N_7564,N_7233,N_7287);
nand U7565 (N_7565,N_7219,N_7050);
and U7566 (N_7566,N_7000,N_7420);
nor U7567 (N_7567,N_7079,N_7387);
nand U7568 (N_7568,N_7172,N_7259);
and U7569 (N_7569,N_7027,N_7105);
and U7570 (N_7570,N_7191,N_7211);
nand U7571 (N_7571,N_7437,N_7267);
and U7572 (N_7572,N_7194,N_7282);
and U7573 (N_7573,N_7302,N_7209);
nor U7574 (N_7574,N_7399,N_7176);
and U7575 (N_7575,N_7129,N_7090);
or U7576 (N_7576,N_7425,N_7288);
nor U7577 (N_7577,N_7196,N_7477);
xnor U7578 (N_7578,N_7037,N_7080);
or U7579 (N_7579,N_7363,N_7034);
nor U7580 (N_7580,N_7207,N_7342);
nor U7581 (N_7581,N_7471,N_7042);
nand U7582 (N_7582,N_7269,N_7456);
nand U7583 (N_7583,N_7041,N_7204);
or U7584 (N_7584,N_7097,N_7237);
and U7585 (N_7585,N_7216,N_7110);
nand U7586 (N_7586,N_7311,N_7138);
and U7587 (N_7587,N_7361,N_7055);
and U7588 (N_7588,N_7398,N_7447);
xnor U7589 (N_7589,N_7117,N_7203);
and U7590 (N_7590,N_7016,N_7151);
nand U7591 (N_7591,N_7160,N_7416);
or U7592 (N_7592,N_7099,N_7064);
nor U7593 (N_7593,N_7373,N_7430);
nand U7594 (N_7594,N_7402,N_7022);
nor U7595 (N_7595,N_7458,N_7081);
nor U7596 (N_7596,N_7077,N_7033);
nand U7597 (N_7597,N_7289,N_7379);
nand U7598 (N_7598,N_7031,N_7161);
nor U7599 (N_7599,N_7186,N_7322);
nor U7600 (N_7600,N_7028,N_7449);
nor U7601 (N_7601,N_7442,N_7212);
nand U7602 (N_7602,N_7073,N_7310);
nor U7603 (N_7603,N_7371,N_7063);
nand U7604 (N_7604,N_7229,N_7325);
or U7605 (N_7605,N_7460,N_7465);
or U7606 (N_7606,N_7159,N_7347);
or U7607 (N_7607,N_7116,N_7114);
nor U7608 (N_7608,N_7221,N_7448);
or U7609 (N_7609,N_7285,N_7149);
and U7610 (N_7610,N_7314,N_7438);
and U7611 (N_7611,N_7455,N_7365);
and U7612 (N_7612,N_7319,N_7275);
or U7613 (N_7613,N_7404,N_7170);
nand U7614 (N_7614,N_7357,N_7429);
nand U7615 (N_7615,N_7001,N_7147);
nor U7616 (N_7616,N_7234,N_7472);
and U7617 (N_7617,N_7434,N_7335);
nand U7618 (N_7618,N_7374,N_7010);
nor U7619 (N_7619,N_7024,N_7096);
nor U7620 (N_7620,N_7290,N_7210);
nand U7621 (N_7621,N_7092,N_7445);
or U7622 (N_7622,N_7089,N_7121);
nor U7623 (N_7623,N_7454,N_7245);
and U7624 (N_7624,N_7436,N_7423);
and U7625 (N_7625,N_7213,N_7336);
nor U7626 (N_7626,N_7164,N_7030);
nor U7627 (N_7627,N_7388,N_7384);
nand U7628 (N_7628,N_7185,N_7094);
or U7629 (N_7629,N_7360,N_7394);
nor U7630 (N_7630,N_7072,N_7184);
and U7631 (N_7631,N_7439,N_7156);
or U7632 (N_7632,N_7088,N_7441);
and U7633 (N_7633,N_7083,N_7205);
xor U7634 (N_7634,N_7093,N_7453);
or U7635 (N_7635,N_7320,N_7307);
and U7636 (N_7636,N_7264,N_7411);
nand U7637 (N_7637,N_7168,N_7070);
or U7638 (N_7638,N_7249,N_7218);
or U7639 (N_7639,N_7023,N_7345);
nand U7640 (N_7640,N_7303,N_7241);
nor U7641 (N_7641,N_7298,N_7065);
and U7642 (N_7642,N_7011,N_7450);
or U7643 (N_7643,N_7333,N_7272);
nor U7644 (N_7644,N_7468,N_7393);
nand U7645 (N_7645,N_7223,N_7199);
nand U7646 (N_7646,N_7144,N_7115);
or U7647 (N_7647,N_7193,N_7341);
nand U7648 (N_7648,N_7405,N_7364);
nand U7649 (N_7649,N_7162,N_7304);
and U7650 (N_7650,N_7330,N_7137);
and U7651 (N_7651,N_7087,N_7396);
or U7652 (N_7652,N_7201,N_7068);
or U7653 (N_7653,N_7474,N_7493);
or U7654 (N_7654,N_7135,N_7026);
nand U7655 (N_7655,N_7486,N_7032);
and U7656 (N_7656,N_7140,N_7318);
nor U7657 (N_7657,N_7494,N_7413);
nor U7658 (N_7658,N_7202,N_7481);
nor U7659 (N_7659,N_7418,N_7317);
or U7660 (N_7660,N_7012,N_7309);
nand U7661 (N_7661,N_7496,N_7100);
or U7662 (N_7662,N_7461,N_7119);
and U7663 (N_7663,N_7052,N_7150);
or U7664 (N_7664,N_7076,N_7334);
and U7665 (N_7665,N_7084,N_7220);
nor U7666 (N_7666,N_7283,N_7085);
nor U7667 (N_7667,N_7417,N_7242);
and U7668 (N_7668,N_7292,N_7057);
nor U7669 (N_7669,N_7198,N_7187);
and U7670 (N_7670,N_7226,N_7051);
or U7671 (N_7671,N_7157,N_7369);
nor U7672 (N_7672,N_7400,N_7459);
nand U7673 (N_7673,N_7136,N_7091);
or U7674 (N_7674,N_7395,N_7328);
nand U7675 (N_7675,N_7059,N_7370);
nor U7676 (N_7676,N_7344,N_7479);
or U7677 (N_7677,N_7443,N_7238);
xor U7678 (N_7678,N_7295,N_7118);
nor U7679 (N_7679,N_7410,N_7432);
and U7680 (N_7680,N_7208,N_7433);
nor U7681 (N_7681,N_7483,N_7274);
or U7682 (N_7682,N_7273,N_7476);
nor U7683 (N_7683,N_7378,N_7348);
nor U7684 (N_7684,N_7108,N_7391);
nand U7685 (N_7685,N_7166,N_7281);
or U7686 (N_7686,N_7424,N_7440);
or U7687 (N_7687,N_7102,N_7230);
nand U7688 (N_7688,N_7020,N_7316);
and U7689 (N_7689,N_7382,N_7251);
nand U7690 (N_7690,N_7291,N_7266);
nand U7691 (N_7691,N_7355,N_7386);
nor U7692 (N_7692,N_7296,N_7124);
nand U7693 (N_7693,N_7473,N_7175);
nor U7694 (N_7694,N_7313,N_7428);
or U7695 (N_7695,N_7060,N_7120);
and U7696 (N_7696,N_7143,N_7372);
and U7697 (N_7697,N_7067,N_7366);
and U7698 (N_7698,N_7227,N_7154);
nand U7699 (N_7699,N_7243,N_7190);
and U7700 (N_7700,N_7036,N_7013);
or U7701 (N_7701,N_7192,N_7095);
nor U7702 (N_7702,N_7415,N_7421);
nand U7703 (N_7703,N_7200,N_7412);
and U7704 (N_7704,N_7206,N_7270);
and U7705 (N_7705,N_7142,N_7451);
or U7706 (N_7706,N_7239,N_7284);
or U7707 (N_7707,N_7414,N_7174);
nand U7708 (N_7708,N_7235,N_7232);
and U7709 (N_7709,N_7004,N_7014);
nand U7710 (N_7710,N_7254,N_7331);
and U7711 (N_7711,N_7182,N_7301);
nor U7712 (N_7712,N_7323,N_7427);
and U7713 (N_7713,N_7240,N_7353);
and U7714 (N_7714,N_7173,N_7406);
or U7715 (N_7715,N_7390,N_7009);
nand U7716 (N_7716,N_7257,N_7324);
nor U7717 (N_7717,N_7127,N_7181);
and U7718 (N_7718,N_7368,N_7049);
or U7719 (N_7719,N_7338,N_7294);
and U7720 (N_7720,N_7058,N_7297);
nand U7721 (N_7721,N_7019,N_7469);
xnor U7722 (N_7722,N_7112,N_7359);
nand U7723 (N_7723,N_7217,N_7040);
or U7724 (N_7724,N_7470,N_7061);
nand U7725 (N_7725,N_7457,N_7376);
nor U7726 (N_7726,N_7163,N_7165);
nand U7727 (N_7727,N_7280,N_7177);
or U7728 (N_7728,N_7002,N_7106);
nor U7729 (N_7729,N_7195,N_7358);
or U7730 (N_7730,N_7356,N_7123);
nor U7731 (N_7731,N_7327,N_7261);
or U7732 (N_7732,N_7380,N_7003);
and U7733 (N_7733,N_7464,N_7248);
nand U7734 (N_7734,N_7132,N_7250);
and U7735 (N_7735,N_7104,N_7179);
nor U7736 (N_7736,N_7039,N_7189);
and U7737 (N_7737,N_7086,N_7048);
and U7738 (N_7738,N_7231,N_7408);
or U7739 (N_7739,N_7152,N_7035);
or U7740 (N_7740,N_7029,N_7277);
or U7741 (N_7741,N_7491,N_7362);
nor U7742 (N_7742,N_7258,N_7467);
or U7743 (N_7743,N_7346,N_7169);
nand U7744 (N_7744,N_7349,N_7300);
nand U7745 (N_7745,N_7183,N_7265);
and U7746 (N_7746,N_7498,N_7463);
or U7747 (N_7747,N_7180,N_7139);
nor U7748 (N_7748,N_7435,N_7490);
nand U7749 (N_7749,N_7141,N_7125);
or U7750 (N_7750,N_7455,N_7096);
nor U7751 (N_7751,N_7169,N_7003);
nor U7752 (N_7752,N_7000,N_7088);
and U7753 (N_7753,N_7017,N_7425);
and U7754 (N_7754,N_7299,N_7298);
nor U7755 (N_7755,N_7235,N_7250);
and U7756 (N_7756,N_7485,N_7003);
and U7757 (N_7757,N_7188,N_7418);
or U7758 (N_7758,N_7396,N_7315);
nand U7759 (N_7759,N_7222,N_7451);
nand U7760 (N_7760,N_7491,N_7431);
and U7761 (N_7761,N_7046,N_7189);
nand U7762 (N_7762,N_7268,N_7108);
nand U7763 (N_7763,N_7488,N_7473);
or U7764 (N_7764,N_7168,N_7182);
and U7765 (N_7765,N_7155,N_7077);
nor U7766 (N_7766,N_7220,N_7194);
or U7767 (N_7767,N_7446,N_7128);
nor U7768 (N_7768,N_7079,N_7389);
and U7769 (N_7769,N_7192,N_7269);
and U7770 (N_7770,N_7120,N_7240);
or U7771 (N_7771,N_7307,N_7354);
nor U7772 (N_7772,N_7280,N_7271);
or U7773 (N_7773,N_7469,N_7070);
nor U7774 (N_7774,N_7054,N_7118);
and U7775 (N_7775,N_7072,N_7486);
nor U7776 (N_7776,N_7406,N_7442);
or U7777 (N_7777,N_7028,N_7352);
or U7778 (N_7778,N_7433,N_7142);
and U7779 (N_7779,N_7228,N_7157);
or U7780 (N_7780,N_7239,N_7071);
or U7781 (N_7781,N_7025,N_7381);
and U7782 (N_7782,N_7339,N_7440);
and U7783 (N_7783,N_7401,N_7134);
and U7784 (N_7784,N_7199,N_7371);
or U7785 (N_7785,N_7370,N_7335);
or U7786 (N_7786,N_7222,N_7359);
or U7787 (N_7787,N_7422,N_7077);
nor U7788 (N_7788,N_7392,N_7357);
nand U7789 (N_7789,N_7113,N_7443);
nand U7790 (N_7790,N_7262,N_7375);
nor U7791 (N_7791,N_7132,N_7313);
or U7792 (N_7792,N_7262,N_7272);
or U7793 (N_7793,N_7237,N_7397);
and U7794 (N_7794,N_7129,N_7150);
and U7795 (N_7795,N_7044,N_7458);
nor U7796 (N_7796,N_7477,N_7315);
nand U7797 (N_7797,N_7332,N_7493);
and U7798 (N_7798,N_7057,N_7051);
nor U7799 (N_7799,N_7102,N_7068);
and U7800 (N_7800,N_7287,N_7072);
and U7801 (N_7801,N_7354,N_7191);
or U7802 (N_7802,N_7303,N_7106);
or U7803 (N_7803,N_7236,N_7350);
nand U7804 (N_7804,N_7421,N_7076);
nand U7805 (N_7805,N_7424,N_7415);
or U7806 (N_7806,N_7232,N_7376);
nand U7807 (N_7807,N_7450,N_7085);
and U7808 (N_7808,N_7383,N_7155);
nor U7809 (N_7809,N_7307,N_7431);
and U7810 (N_7810,N_7431,N_7306);
and U7811 (N_7811,N_7370,N_7069);
or U7812 (N_7812,N_7457,N_7201);
nand U7813 (N_7813,N_7164,N_7006);
and U7814 (N_7814,N_7337,N_7447);
nand U7815 (N_7815,N_7477,N_7216);
or U7816 (N_7816,N_7285,N_7017);
and U7817 (N_7817,N_7293,N_7348);
nor U7818 (N_7818,N_7407,N_7449);
or U7819 (N_7819,N_7359,N_7092);
and U7820 (N_7820,N_7377,N_7242);
and U7821 (N_7821,N_7177,N_7175);
or U7822 (N_7822,N_7106,N_7155);
nand U7823 (N_7823,N_7343,N_7137);
and U7824 (N_7824,N_7012,N_7166);
xor U7825 (N_7825,N_7474,N_7106);
and U7826 (N_7826,N_7212,N_7189);
and U7827 (N_7827,N_7486,N_7140);
nor U7828 (N_7828,N_7457,N_7053);
or U7829 (N_7829,N_7136,N_7078);
or U7830 (N_7830,N_7338,N_7175);
nor U7831 (N_7831,N_7289,N_7084);
or U7832 (N_7832,N_7283,N_7221);
nor U7833 (N_7833,N_7370,N_7297);
and U7834 (N_7834,N_7469,N_7341);
and U7835 (N_7835,N_7405,N_7471);
nand U7836 (N_7836,N_7265,N_7301);
and U7837 (N_7837,N_7431,N_7145);
nand U7838 (N_7838,N_7403,N_7473);
and U7839 (N_7839,N_7498,N_7194);
nor U7840 (N_7840,N_7470,N_7421);
nor U7841 (N_7841,N_7184,N_7337);
and U7842 (N_7842,N_7087,N_7479);
nor U7843 (N_7843,N_7408,N_7356);
nor U7844 (N_7844,N_7385,N_7245);
nand U7845 (N_7845,N_7153,N_7248);
nand U7846 (N_7846,N_7249,N_7316);
nand U7847 (N_7847,N_7176,N_7218);
nor U7848 (N_7848,N_7463,N_7305);
nor U7849 (N_7849,N_7132,N_7281);
nor U7850 (N_7850,N_7433,N_7003);
and U7851 (N_7851,N_7332,N_7141);
nor U7852 (N_7852,N_7155,N_7220);
or U7853 (N_7853,N_7238,N_7152);
nor U7854 (N_7854,N_7352,N_7194);
and U7855 (N_7855,N_7040,N_7189);
and U7856 (N_7856,N_7076,N_7136);
nor U7857 (N_7857,N_7396,N_7112);
or U7858 (N_7858,N_7418,N_7288);
or U7859 (N_7859,N_7282,N_7339);
nand U7860 (N_7860,N_7178,N_7389);
and U7861 (N_7861,N_7137,N_7405);
or U7862 (N_7862,N_7069,N_7420);
nor U7863 (N_7863,N_7332,N_7115);
nand U7864 (N_7864,N_7493,N_7018);
nand U7865 (N_7865,N_7256,N_7412);
and U7866 (N_7866,N_7490,N_7169);
nor U7867 (N_7867,N_7499,N_7316);
or U7868 (N_7868,N_7112,N_7160);
and U7869 (N_7869,N_7400,N_7263);
nand U7870 (N_7870,N_7458,N_7169);
xnor U7871 (N_7871,N_7439,N_7031);
or U7872 (N_7872,N_7128,N_7422);
or U7873 (N_7873,N_7266,N_7028);
or U7874 (N_7874,N_7011,N_7111);
or U7875 (N_7875,N_7135,N_7013);
and U7876 (N_7876,N_7140,N_7485);
nand U7877 (N_7877,N_7207,N_7014);
nor U7878 (N_7878,N_7126,N_7156);
xor U7879 (N_7879,N_7426,N_7009);
nor U7880 (N_7880,N_7351,N_7284);
nand U7881 (N_7881,N_7182,N_7395);
and U7882 (N_7882,N_7348,N_7004);
and U7883 (N_7883,N_7336,N_7449);
and U7884 (N_7884,N_7499,N_7227);
or U7885 (N_7885,N_7101,N_7310);
xor U7886 (N_7886,N_7032,N_7120);
nor U7887 (N_7887,N_7288,N_7228);
and U7888 (N_7888,N_7076,N_7468);
and U7889 (N_7889,N_7261,N_7099);
nor U7890 (N_7890,N_7397,N_7348);
or U7891 (N_7891,N_7081,N_7256);
nor U7892 (N_7892,N_7085,N_7499);
or U7893 (N_7893,N_7175,N_7230);
or U7894 (N_7894,N_7098,N_7274);
nor U7895 (N_7895,N_7420,N_7322);
and U7896 (N_7896,N_7145,N_7138);
or U7897 (N_7897,N_7473,N_7211);
and U7898 (N_7898,N_7421,N_7001);
nor U7899 (N_7899,N_7342,N_7078);
nand U7900 (N_7900,N_7487,N_7058);
or U7901 (N_7901,N_7187,N_7131);
nand U7902 (N_7902,N_7139,N_7384);
nand U7903 (N_7903,N_7192,N_7263);
and U7904 (N_7904,N_7370,N_7325);
or U7905 (N_7905,N_7152,N_7499);
and U7906 (N_7906,N_7128,N_7042);
or U7907 (N_7907,N_7294,N_7383);
or U7908 (N_7908,N_7056,N_7190);
nor U7909 (N_7909,N_7085,N_7016);
or U7910 (N_7910,N_7110,N_7163);
nand U7911 (N_7911,N_7344,N_7375);
and U7912 (N_7912,N_7093,N_7062);
nor U7913 (N_7913,N_7415,N_7391);
or U7914 (N_7914,N_7419,N_7339);
nor U7915 (N_7915,N_7035,N_7204);
nor U7916 (N_7916,N_7343,N_7247);
and U7917 (N_7917,N_7245,N_7105);
nor U7918 (N_7918,N_7093,N_7185);
nand U7919 (N_7919,N_7337,N_7057);
nor U7920 (N_7920,N_7100,N_7139);
nand U7921 (N_7921,N_7194,N_7135);
and U7922 (N_7922,N_7198,N_7057);
or U7923 (N_7923,N_7354,N_7363);
or U7924 (N_7924,N_7303,N_7483);
nor U7925 (N_7925,N_7285,N_7178);
nor U7926 (N_7926,N_7161,N_7330);
nand U7927 (N_7927,N_7188,N_7073);
and U7928 (N_7928,N_7434,N_7371);
and U7929 (N_7929,N_7438,N_7159);
nor U7930 (N_7930,N_7098,N_7373);
or U7931 (N_7931,N_7293,N_7309);
or U7932 (N_7932,N_7468,N_7153);
and U7933 (N_7933,N_7065,N_7051);
nand U7934 (N_7934,N_7406,N_7069);
nand U7935 (N_7935,N_7025,N_7017);
nor U7936 (N_7936,N_7419,N_7174);
nand U7937 (N_7937,N_7031,N_7442);
nand U7938 (N_7938,N_7487,N_7179);
nor U7939 (N_7939,N_7342,N_7447);
and U7940 (N_7940,N_7017,N_7210);
nand U7941 (N_7941,N_7354,N_7141);
nor U7942 (N_7942,N_7472,N_7073);
and U7943 (N_7943,N_7203,N_7415);
and U7944 (N_7944,N_7092,N_7180);
nor U7945 (N_7945,N_7097,N_7113);
and U7946 (N_7946,N_7229,N_7320);
nor U7947 (N_7947,N_7264,N_7435);
nor U7948 (N_7948,N_7003,N_7479);
and U7949 (N_7949,N_7243,N_7308);
nor U7950 (N_7950,N_7029,N_7387);
nor U7951 (N_7951,N_7171,N_7116);
and U7952 (N_7952,N_7341,N_7258);
nand U7953 (N_7953,N_7402,N_7136);
nor U7954 (N_7954,N_7008,N_7261);
nand U7955 (N_7955,N_7026,N_7120);
and U7956 (N_7956,N_7301,N_7293);
nand U7957 (N_7957,N_7371,N_7266);
or U7958 (N_7958,N_7206,N_7120);
and U7959 (N_7959,N_7375,N_7175);
and U7960 (N_7960,N_7022,N_7345);
and U7961 (N_7961,N_7257,N_7482);
and U7962 (N_7962,N_7276,N_7175);
or U7963 (N_7963,N_7138,N_7287);
and U7964 (N_7964,N_7400,N_7172);
and U7965 (N_7965,N_7094,N_7171);
or U7966 (N_7966,N_7292,N_7037);
xnor U7967 (N_7967,N_7221,N_7085);
nand U7968 (N_7968,N_7142,N_7015);
or U7969 (N_7969,N_7243,N_7424);
and U7970 (N_7970,N_7463,N_7047);
nor U7971 (N_7971,N_7421,N_7050);
nor U7972 (N_7972,N_7071,N_7132);
and U7973 (N_7973,N_7179,N_7433);
and U7974 (N_7974,N_7069,N_7088);
nor U7975 (N_7975,N_7434,N_7033);
and U7976 (N_7976,N_7166,N_7386);
or U7977 (N_7977,N_7433,N_7195);
nor U7978 (N_7978,N_7155,N_7192);
nand U7979 (N_7979,N_7029,N_7150);
nand U7980 (N_7980,N_7001,N_7311);
nand U7981 (N_7981,N_7467,N_7202);
and U7982 (N_7982,N_7106,N_7326);
or U7983 (N_7983,N_7283,N_7181);
nor U7984 (N_7984,N_7131,N_7204);
or U7985 (N_7985,N_7041,N_7468);
and U7986 (N_7986,N_7107,N_7020);
or U7987 (N_7987,N_7005,N_7161);
nor U7988 (N_7988,N_7282,N_7497);
and U7989 (N_7989,N_7398,N_7401);
and U7990 (N_7990,N_7384,N_7459);
nor U7991 (N_7991,N_7215,N_7234);
or U7992 (N_7992,N_7266,N_7185);
nand U7993 (N_7993,N_7269,N_7384);
nor U7994 (N_7994,N_7263,N_7489);
and U7995 (N_7995,N_7330,N_7194);
and U7996 (N_7996,N_7072,N_7114);
or U7997 (N_7997,N_7266,N_7166);
nor U7998 (N_7998,N_7135,N_7357);
nor U7999 (N_7999,N_7154,N_7204);
nor U8000 (N_8000,N_7937,N_7824);
nor U8001 (N_8001,N_7548,N_7953);
or U8002 (N_8002,N_7822,N_7729);
or U8003 (N_8003,N_7651,N_7900);
nand U8004 (N_8004,N_7679,N_7569);
and U8005 (N_8005,N_7701,N_7630);
and U8006 (N_8006,N_7888,N_7872);
or U8007 (N_8007,N_7594,N_7510);
or U8008 (N_8008,N_7547,N_7997);
or U8009 (N_8009,N_7757,N_7935);
nand U8010 (N_8010,N_7782,N_7852);
or U8011 (N_8011,N_7671,N_7948);
and U8012 (N_8012,N_7654,N_7882);
and U8013 (N_8013,N_7781,N_7850);
and U8014 (N_8014,N_7658,N_7620);
or U8015 (N_8015,N_7631,N_7675);
or U8016 (N_8016,N_7720,N_7921);
nand U8017 (N_8017,N_7592,N_7686);
xor U8018 (N_8018,N_7744,N_7881);
nand U8019 (N_8019,N_7857,N_7810);
nand U8020 (N_8020,N_7835,N_7732);
or U8021 (N_8021,N_7929,N_7940);
nor U8022 (N_8022,N_7661,N_7840);
nand U8023 (N_8023,N_7537,N_7821);
or U8024 (N_8024,N_7767,N_7559);
nand U8025 (N_8025,N_7933,N_7965);
and U8026 (N_8026,N_7946,N_7994);
nand U8027 (N_8027,N_7606,N_7819);
and U8028 (N_8028,N_7684,N_7804);
and U8029 (N_8029,N_7565,N_7632);
and U8030 (N_8030,N_7643,N_7977);
nand U8031 (N_8031,N_7723,N_7644);
or U8032 (N_8032,N_7750,N_7827);
or U8033 (N_8033,N_7902,N_7621);
or U8034 (N_8034,N_7527,N_7634);
and U8035 (N_8035,N_7628,N_7754);
and U8036 (N_8036,N_7982,N_7549);
nor U8037 (N_8037,N_7627,N_7554);
nand U8038 (N_8038,N_7942,N_7834);
nor U8039 (N_8039,N_7955,N_7867);
nand U8040 (N_8040,N_7746,N_7712);
and U8041 (N_8041,N_7980,N_7635);
nand U8042 (N_8042,N_7693,N_7597);
nor U8043 (N_8043,N_7970,N_7738);
nor U8044 (N_8044,N_7956,N_7832);
and U8045 (N_8045,N_7854,N_7960);
xor U8046 (N_8046,N_7568,N_7589);
or U8047 (N_8047,N_7562,N_7523);
or U8048 (N_8048,N_7696,N_7555);
nand U8049 (N_8049,N_7563,N_7914);
and U8050 (N_8050,N_7728,N_7919);
or U8051 (N_8051,N_7645,N_7864);
or U8052 (N_8052,N_7668,N_7927);
nor U8053 (N_8053,N_7969,N_7949);
and U8054 (N_8054,N_7616,N_7598);
and U8055 (N_8055,N_7709,N_7784);
and U8056 (N_8056,N_7747,N_7716);
nand U8057 (N_8057,N_7901,N_7637);
nand U8058 (N_8058,N_7930,N_7601);
and U8059 (N_8059,N_7939,N_7670);
and U8060 (N_8060,N_7604,N_7558);
or U8061 (N_8061,N_7531,N_7771);
or U8062 (N_8062,N_7653,N_7789);
xor U8063 (N_8063,N_7665,N_7599);
nor U8064 (N_8064,N_7695,N_7963);
nand U8065 (N_8065,N_7507,N_7988);
and U8066 (N_8066,N_7826,N_7780);
or U8067 (N_8067,N_7706,N_7806);
or U8068 (N_8068,N_7952,N_7813);
or U8069 (N_8069,N_7543,N_7557);
and U8070 (N_8070,N_7535,N_7736);
and U8071 (N_8071,N_7674,N_7760);
nand U8072 (N_8072,N_7950,N_7776);
or U8073 (N_8073,N_7801,N_7849);
and U8074 (N_8074,N_7719,N_7799);
nand U8075 (N_8075,N_7517,N_7505);
nand U8076 (N_8076,N_7739,N_7820);
nand U8077 (N_8077,N_7615,N_7646);
nand U8078 (N_8078,N_7979,N_7972);
nand U8079 (N_8079,N_7542,N_7957);
or U8080 (N_8080,N_7707,N_7509);
nand U8081 (N_8081,N_7540,N_7607);
nand U8082 (N_8082,N_7530,N_7725);
nand U8083 (N_8083,N_7690,N_7534);
or U8084 (N_8084,N_7873,N_7924);
and U8085 (N_8085,N_7842,N_7858);
or U8086 (N_8086,N_7923,N_7713);
nand U8087 (N_8087,N_7722,N_7614);
nand U8088 (N_8088,N_7875,N_7539);
nor U8089 (N_8089,N_7830,N_7947);
nand U8090 (N_8090,N_7501,N_7551);
nor U8091 (N_8091,N_7649,N_7681);
nor U8092 (N_8092,N_7828,N_7787);
nor U8093 (N_8093,N_7673,N_7639);
and U8094 (N_8094,N_7934,N_7998);
or U8095 (N_8095,N_7912,N_7847);
and U8096 (N_8096,N_7717,N_7591);
or U8097 (N_8097,N_7529,N_7610);
nor U8098 (N_8098,N_7660,N_7974);
nand U8099 (N_8099,N_7571,N_7803);
nor U8100 (N_8100,N_7567,N_7778);
or U8101 (N_8101,N_7506,N_7917);
or U8102 (N_8102,N_7552,N_7903);
nor U8103 (N_8103,N_7609,N_7731);
nor U8104 (N_8104,N_7996,N_7968);
nand U8105 (N_8105,N_7790,N_7544);
nand U8106 (N_8106,N_7655,N_7812);
and U8107 (N_8107,N_7876,N_7909);
nor U8108 (N_8108,N_7978,N_7848);
or U8109 (N_8109,N_7877,N_7667);
or U8110 (N_8110,N_7991,N_7920);
nand U8111 (N_8111,N_7522,N_7619);
nor U8112 (N_8112,N_7724,N_7663);
or U8113 (N_8113,N_7758,N_7593);
and U8114 (N_8114,N_7669,N_7737);
nor U8115 (N_8115,N_7865,N_7704);
or U8116 (N_8116,N_7556,N_7611);
and U8117 (N_8117,N_7536,N_7938);
or U8118 (N_8118,N_7676,N_7561);
nand U8119 (N_8119,N_7814,N_7577);
nand U8120 (N_8120,N_7648,N_7659);
nor U8121 (N_8121,N_7702,N_7697);
or U8122 (N_8122,N_7642,N_7795);
nor U8123 (N_8123,N_7786,N_7560);
nand U8124 (N_8124,N_7975,N_7762);
or U8125 (N_8125,N_7756,N_7613);
nor U8126 (N_8126,N_7764,N_7584);
or U8127 (N_8127,N_7809,N_7951);
and U8128 (N_8128,N_7656,N_7532);
nor U8129 (N_8129,N_7961,N_7871);
nor U8130 (N_8130,N_7817,N_7741);
nand U8131 (N_8131,N_7906,N_7726);
nor U8132 (N_8132,N_7973,N_7678);
nand U8133 (N_8133,N_7993,N_7868);
nor U8134 (N_8134,N_7735,N_7664);
nor U8135 (N_8135,N_7883,N_7805);
nor U8136 (N_8136,N_7926,N_7683);
and U8137 (N_8137,N_7662,N_7769);
and U8138 (N_8138,N_7859,N_7765);
or U8139 (N_8139,N_7770,N_7528);
and U8140 (N_8140,N_7845,N_7853);
nor U8141 (N_8141,N_7740,N_7525);
or U8142 (N_8142,N_7889,N_7582);
or U8143 (N_8143,N_7798,N_7541);
and U8144 (N_8144,N_7596,N_7886);
nand U8145 (N_8145,N_7892,N_7691);
and U8146 (N_8146,N_7841,N_7800);
and U8147 (N_8147,N_7692,N_7581);
or U8148 (N_8148,N_7755,N_7846);
nand U8149 (N_8149,N_7964,N_7761);
and U8150 (N_8150,N_7721,N_7989);
or U8151 (N_8151,N_7869,N_7793);
nand U8152 (N_8152,N_7703,N_7836);
or U8153 (N_8153,N_7500,N_7833);
nor U8154 (N_8154,N_7626,N_7700);
nand U8155 (N_8155,N_7585,N_7629);
nor U8156 (N_8156,N_7519,N_7575);
or U8157 (N_8157,N_7945,N_7579);
nand U8158 (N_8158,N_7516,N_7823);
nor U8159 (N_8159,N_7890,N_7520);
nand U8160 (N_8160,N_7602,N_7983);
and U8161 (N_8161,N_7860,N_7566);
or U8162 (N_8162,N_7502,N_7794);
and U8163 (N_8163,N_7941,N_7608);
or U8164 (N_8164,N_7698,N_7618);
nand U8165 (N_8165,N_7936,N_7672);
nand U8166 (N_8166,N_7636,N_7650);
and U8167 (N_8167,N_7897,N_7981);
nor U8168 (N_8168,N_7987,N_7887);
nor U8169 (N_8169,N_7788,N_7526);
and U8170 (N_8170,N_7647,N_7633);
nor U8171 (N_8171,N_7785,N_7796);
or U8172 (N_8172,N_7775,N_7570);
nor U8173 (N_8173,N_7811,N_7898);
nor U8174 (N_8174,N_7766,N_7962);
or U8175 (N_8175,N_7504,N_7727);
nand U8176 (N_8176,N_7880,N_7515);
or U8177 (N_8177,N_7751,N_7622);
and U8178 (N_8178,N_7710,N_7605);
nor U8179 (N_8179,N_7894,N_7885);
nand U8180 (N_8180,N_7773,N_7652);
nand U8181 (N_8181,N_7689,N_7954);
and U8182 (N_8182,N_7512,N_7878);
xnor U8183 (N_8183,N_7641,N_7791);
or U8184 (N_8184,N_7843,N_7545);
nor U8185 (N_8185,N_7931,N_7904);
nor U8186 (N_8186,N_7513,N_7907);
nor U8187 (N_8187,N_7518,N_7774);
or U8188 (N_8188,N_7600,N_7743);
or U8189 (N_8189,N_7682,N_7896);
nor U8190 (N_8190,N_7966,N_7984);
or U8191 (N_8191,N_7590,N_7863);
or U8192 (N_8192,N_7573,N_7752);
nor U8193 (N_8193,N_7851,N_7932);
nor U8194 (N_8194,N_7779,N_7734);
and U8195 (N_8195,N_7856,N_7546);
or U8196 (N_8196,N_7718,N_7943);
xor U8197 (N_8197,N_7638,N_7913);
nand U8198 (N_8198,N_7699,N_7874);
or U8199 (N_8199,N_7772,N_7837);
or U8200 (N_8200,N_7503,N_7749);
and U8201 (N_8201,N_7838,N_7657);
nand U8202 (N_8202,N_7999,N_7958);
nand U8203 (N_8203,N_7623,N_7587);
and U8204 (N_8204,N_7553,N_7915);
xor U8205 (N_8205,N_7730,N_7524);
and U8206 (N_8206,N_7944,N_7899);
nor U8207 (N_8207,N_7844,N_7550);
and U8208 (N_8208,N_7508,N_7574);
or U8209 (N_8209,N_7879,N_7688);
nor U8210 (N_8210,N_7768,N_7870);
nand U8211 (N_8211,N_7759,N_7715);
and U8212 (N_8212,N_7578,N_7891);
xor U8213 (N_8213,N_7792,N_7617);
and U8214 (N_8214,N_7777,N_7588);
and U8215 (N_8215,N_7797,N_7967);
or U8216 (N_8216,N_7910,N_7816);
nand U8217 (N_8217,N_7839,N_7884);
or U8218 (N_8218,N_7564,N_7831);
and U8219 (N_8219,N_7521,N_7916);
and U8220 (N_8220,N_7625,N_7708);
nor U8221 (N_8221,N_7818,N_7745);
and U8222 (N_8222,N_7925,N_7783);
nand U8223 (N_8223,N_7862,N_7538);
or U8224 (N_8224,N_7829,N_7624);
or U8225 (N_8225,N_7855,N_7705);
nand U8226 (N_8226,N_7576,N_7733);
nor U8227 (N_8227,N_7612,N_7990);
or U8228 (N_8228,N_7895,N_7687);
and U8229 (N_8229,N_7685,N_7511);
nor U8230 (N_8230,N_7911,N_7677);
and U8231 (N_8231,N_7866,N_7815);
nor U8232 (N_8232,N_7807,N_7918);
or U8233 (N_8233,N_7742,N_7959);
nand U8234 (N_8234,N_7583,N_7893);
or U8235 (N_8235,N_7533,N_7825);
nand U8236 (N_8236,N_7861,N_7595);
nor U8237 (N_8237,N_7666,N_7908);
nand U8238 (N_8238,N_7971,N_7763);
and U8239 (N_8239,N_7976,N_7748);
or U8240 (N_8240,N_7586,N_7711);
nand U8241 (N_8241,N_7640,N_7753);
and U8242 (N_8242,N_7922,N_7802);
nor U8243 (N_8243,N_7694,N_7714);
or U8244 (N_8244,N_7572,N_7603);
nand U8245 (N_8245,N_7995,N_7680);
nand U8246 (N_8246,N_7985,N_7992);
nor U8247 (N_8247,N_7514,N_7580);
or U8248 (N_8248,N_7928,N_7808);
and U8249 (N_8249,N_7905,N_7986);
nor U8250 (N_8250,N_7612,N_7513);
and U8251 (N_8251,N_7848,N_7924);
or U8252 (N_8252,N_7694,N_7784);
and U8253 (N_8253,N_7811,N_7889);
nand U8254 (N_8254,N_7578,N_7687);
or U8255 (N_8255,N_7714,N_7648);
or U8256 (N_8256,N_7545,N_7766);
and U8257 (N_8257,N_7848,N_7683);
or U8258 (N_8258,N_7953,N_7762);
nor U8259 (N_8259,N_7587,N_7552);
nand U8260 (N_8260,N_7630,N_7915);
nor U8261 (N_8261,N_7572,N_7685);
or U8262 (N_8262,N_7949,N_7674);
or U8263 (N_8263,N_7676,N_7847);
and U8264 (N_8264,N_7866,N_7967);
and U8265 (N_8265,N_7629,N_7891);
or U8266 (N_8266,N_7730,N_7970);
nand U8267 (N_8267,N_7709,N_7631);
nand U8268 (N_8268,N_7811,N_7843);
nor U8269 (N_8269,N_7808,N_7528);
nor U8270 (N_8270,N_7952,N_7948);
nor U8271 (N_8271,N_7859,N_7862);
or U8272 (N_8272,N_7514,N_7617);
nor U8273 (N_8273,N_7508,N_7578);
or U8274 (N_8274,N_7753,N_7901);
or U8275 (N_8275,N_7793,N_7990);
nor U8276 (N_8276,N_7700,N_7863);
nor U8277 (N_8277,N_7932,N_7903);
nor U8278 (N_8278,N_7962,N_7773);
and U8279 (N_8279,N_7758,N_7938);
and U8280 (N_8280,N_7559,N_7577);
nor U8281 (N_8281,N_7633,N_7604);
nand U8282 (N_8282,N_7806,N_7889);
or U8283 (N_8283,N_7559,N_7870);
or U8284 (N_8284,N_7735,N_7920);
nor U8285 (N_8285,N_7599,N_7794);
and U8286 (N_8286,N_7579,N_7788);
and U8287 (N_8287,N_7859,N_7683);
nor U8288 (N_8288,N_7784,N_7515);
nand U8289 (N_8289,N_7839,N_7770);
and U8290 (N_8290,N_7934,N_7677);
nor U8291 (N_8291,N_7841,N_7591);
nand U8292 (N_8292,N_7604,N_7661);
or U8293 (N_8293,N_7940,N_7938);
or U8294 (N_8294,N_7815,N_7683);
and U8295 (N_8295,N_7848,N_7750);
nand U8296 (N_8296,N_7675,N_7550);
or U8297 (N_8297,N_7609,N_7944);
nor U8298 (N_8298,N_7745,N_7619);
nor U8299 (N_8299,N_7771,N_7853);
nand U8300 (N_8300,N_7535,N_7553);
or U8301 (N_8301,N_7634,N_7546);
nor U8302 (N_8302,N_7527,N_7681);
nor U8303 (N_8303,N_7637,N_7954);
nor U8304 (N_8304,N_7736,N_7542);
and U8305 (N_8305,N_7861,N_7763);
nand U8306 (N_8306,N_7917,N_7920);
and U8307 (N_8307,N_7785,N_7846);
nor U8308 (N_8308,N_7985,N_7739);
and U8309 (N_8309,N_7509,N_7766);
and U8310 (N_8310,N_7582,N_7813);
or U8311 (N_8311,N_7770,N_7750);
nand U8312 (N_8312,N_7942,N_7759);
nand U8313 (N_8313,N_7520,N_7888);
nand U8314 (N_8314,N_7871,N_7648);
or U8315 (N_8315,N_7946,N_7532);
nand U8316 (N_8316,N_7574,N_7897);
nand U8317 (N_8317,N_7977,N_7964);
xnor U8318 (N_8318,N_7565,N_7766);
nor U8319 (N_8319,N_7785,N_7798);
nand U8320 (N_8320,N_7523,N_7779);
or U8321 (N_8321,N_7951,N_7823);
nand U8322 (N_8322,N_7745,N_7638);
nand U8323 (N_8323,N_7571,N_7742);
and U8324 (N_8324,N_7636,N_7628);
nor U8325 (N_8325,N_7736,N_7740);
and U8326 (N_8326,N_7794,N_7805);
nor U8327 (N_8327,N_7838,N_7610);
nand U8328 (N_8328,N_7894,N_7993);
nand U8329 (N_8329,N_7852,N_7945);
xor U8330 (N_8330,N_7680,N_7734);
or U8331 (N_8331,N_7870,N_7919);
nand U8332 (N_8332,N_7618,N_7931);
nor U8333 (N_8333,N_7606,N_7546);
nor U8334 (N_8334,N_7849,N_7807);
and U8335 (N_8335,N_7862,N_7969);
or U8336 (N_8336,N_7536,N_7798);
and U8337 (N_8337,N_7941,N_7992);
or U8338 (N_8338,N_7507,N_7532);
nand U8339 (N_8339,N_7961,N_7928);
and U8340 (N_8340,N_7990,N_7575);
nor U8341 (N_8341,N_7513,N_7867);
nor U8342 (N_8342,N_7781,N_7630);
nor U8343 (N_8343,N_7659,N_7926);
nand U8344 (N_8344,N_7667,N_7534);
nor U8345 (N_8345,N_7941,N_7688);
nor U8346 (N_8346,N_7786,N_7991);
nand U8347 (N_8347,N_7924,N_7611);
nor U8348 (N_8348,N_7544,N_7524);
or U8349 (N_8349,N_7734,N_7635);
nor U8350 (N_8350,N_7923,N_7681);
nor U8351 (N_8351,N_7543,N_7573);
and U8352 (N_8352,N_7770,N_7564);
and U8353 (N_8353,N_7909,N_7767);
nor U8354 (N_8354,N_7516,N_7637);
and U8355 (N_8355,N_7830,N_7587);
nor U8356 (N_8356,N_7802,N_7933);
nand U8357 (N_8357,N_7624,N_7793);
or U8358 (N_8358,N_7564,N_7833);
or U8359 (N_8359,N_7505,N_7538);
nand U8360 (N_8360,N_7954,N_7620);
nor U8361 (N_8361,N_7727,N_7647);
and U8362 (N_8362,N_7778,N_7712);
and U8363 (N_8363,N_7527,N_7798);
xnor U8364 (N_8364,N_7876,N_7646);
nand U8365 (N_8365,N_7697,N_7621);
nor U8366 (N_8366,N_7890,N_7887);
xor U8367 (N_8367,N_7949,N_7964);
nor U8368 (N_8368,N_7742,N_7971);
nor U8369 (N_8369,N_7617,N_7779);
nand U8370 (N_8370,N_7831,N_7615);
and U8371 (N_8371,N_7957,N_7974);
and U8372 (N_8372,N_7686,N_7727);
and U8373 (N_8373,N_7882,N_7526);
or U8374 (N_8374,N_7817,N_7562);
or U8375 (N_8375,N_7995,N_7661);
nor U8376 (N_8376,N_7987,N_7817);
nor U8377 (N_8377,N_7923,N_7695);
nand U8378 (N_8378,N_7733,N_7747);
or U8379 (N_8379,N_7811,N_7542);
and U8380 (N_8380,N_7510,N_7867);
nand U8381 (N_8381,N_7948,N_7722);
nand U8382 (N_8382,N_7684,N_7981);
nor U8383 (N_8383,N_7815,N_7958);
and U8384 (N_8384,N_7596,N_7565);
and U8385 (N_8385,N_7909,N_7963);
nand U8386 (N_8386,N_7584,N_7600);
or U8387 (N_8387,N_7538,N_7586);
nor U8388 (N_8388,N_7696,N_7785);
and U8389 (N_8389,N_7765,N_7508);
or U8390 (N_8390,N_7593,N_7715);
nor U8391 (N_8391,N_7741,N_7762);
or U8392 (N_8392,N_7919,N_7907);
nand U8393 (N_8393,N_7776,N_7793);
nor U8394 (N_8394,N_7742,N_7666);
nor U8395 (N_8395,N_7549,N_7608);
and U8396 (N_8396,N_7566,N_7996);
nor U8397 (N_8397,N_7977,N_7702);
and U8398 (N_8398,N_7974,N_7823);
or U8399 (N_8399,N_7975,N_7870);
or U8400 (N_8400,N_7943,N_7857);
nor U8401 (N_8401,N_7625,N_7720);
and U8402 (N_8402,N_7674,N_7560);
nand U8403 (N_8403,N_7897,N_7661);
nor U8404 (N_8404,N_7634,N_7577);
nand U8405 (N_8405,N_7513,N_7514);
or U8406 (N_8406,N_7751,N_7712);
or U8407 (N_8407,N_7526,N_7917);
nand U8408 (N_8408,N_7712,N_7768);
nor U8409 (N_8409,N_7957,N_7553);
or U8410 (N_8410,N_7636,N_7511);
and U8411 (N_8411,N_7842,N_7785);
or U8412 (N_8412,N_7529,N_7785);
and U8413 (N_8413,N_7509,N_7813);
nand U8414 (N_8414,N_7995,N_7694);
or U8415 (N_8415,N_7731,N_7550);
or U8416 (N_8416,N_7966,N_7996);
or U8417 (N_8417,N_7842,N_7541);
or U8418 (N_8418,N_7603,N_7501);
or U8419 (N_8419,N_7529,N_7962);
or U8420 (N_8420,N_7683,N_7804);
and U8421 (N_8421,N_7501,N_7744);
and U8422 (N_8422,N_7672,N_7675);
nor U8423 (N_8423,N_7879,N_7576);
xor U8424 (N_8424,N_7595,N_7955);
and U8425 (N_8425,N_7949,N_7582);
nor U8426 (N_8426,N_7717,N_7674);
and U8427 (N_8427,N_7520,N_7629);
or U8428 (N_8428,N_7947,N_7565);
nand U8429 (N_8429,N_7610,N_7914);
nor U8430 (N_8430,N_7569,N_7764);
or U8431 (N_8431,N_7949,N_7635);
or U8432 (N_8432,N_7783,N_7812);
or U8433 (N_8433,N_7586,N_7587);
and U8434 (N_8434,N_7923,N_7635);
and U8435 (N_8435,N_7712,N_7636);
or U8436 (N_8436,N_7961,N_7982);
and U8437 (N_8437,N_7549,N_7704);
or U8438 (N_8438,N_7783,N_7759);
or U8439 (N_8439,N_7561,N_7701);
nand U8440 (N_8440,N_7541,N_7888);
and U8441 (N_8441,N_7793,N_7625);
nand U8442 (N_8442,N_7933,N_7539);
or U8443 (N_8443,N_7550,N_7749);
and U8444 (N_8444,N_7633,N_7976);
nand U8445 (N_8445,N_7899,N_7839);
xor U8446 (N_8446,N_7515,N_7591);
nand U8447 (N_8447,N_7681,N_7949);
nand U8448 (N_8448,N_7777,N_7758);
nand U8449 (N_8449,N_7865,N_7711);
nand U8450 (N_8450,N_7747,N_7994);
nor U8451 (N_8451,N_7965,N_7820);
and U8452 (N_8452,N_7697,N_7643);
and U8453 (N_8453,N_7605,N_7740);
or U8454 (N_8454,N_7827,N_7885);
nand U8455 (N_8455,N_7547,N_7597);
nand U8456 (N_8456,N_7661,N_7674);
nor U8457 (N_8457,N_7791,N_7606);
and U8458 (N_8458,N_7631,N_7871);
nand U8459 (N_8459,N_7510,N_7516);
and U8460 (N_8460,N_7627,N_7846);
and U8461 (N_8461,N_7515,N_7843);
or U8462 (N_8462,N_7870,N_7638);
nand U8463 (N_8463,N_7670,N_7624);
nand U8464 (N_8464,N_7501,N_7576);
or U8465 (N_8465,N_7763,N_7707);
nand U8466 (N_8466,N_7609,N_7799);
or U8467 (N_8467,N_7577,N_7586);
nor U8468 (N_8468,N_7548,N_7877);
or U8469 (N_8469,N_7858,N_7577);
nand U8470 (N_8470,N_7976,N_7806);
and U8471 (N_8471,N_7769,N_7949);
nand U8472 (N_8472,N_7505,N_7780);
and U8473 (N_8473,N_7888,N_7633);
or U8474 (N_8474,N_7548,N_7898);
and U8475 (N_8475,N_7948,N_7552);
nor U8476 (N_8476,N_7660,N_7608);
nand U8477 (N_8477,N_7676,N_7833);
and U8478 (N_8478,N_7565,N_7675);
nor U8479 (N_8479,N_7898,N_7629);
or U8480 (N_8480,N_7892,N_7646);
or U8481 (N_8481,N_7629,N_7676);
nand U8482 (N_8482,N_7614,N_7814);
nor U8483 (N_8483,N_7762,N_7966);
or U8484 (N_8484,N_7660,N_7534);
nand U8485 (N_8485,N_7797,N_7578);
nand U8486 (N_8486,N_7566,N_7899);
nand U8487 (N_8487,N_7529,N_7767);
and U8488 (N_8488,N_7751,N_7606);
nand U8489 (N_8489,N_7622,N_7550);
nor U8490 (N_8490,N_7882,N_7860);
and U8491 (N_8491,N_7735,N_7520);
nand U8492 (N_8492,N_7980,N_7516);
and U8493 (N_8493,N_7880,N_7907);
and U8494 (N_8494,N_7879,N_7704);
nor U8495 (N_8495,N_7686,N_7689);
and U8496 (N_8496,N_7780,N_7645);
nand U8497 (N_8497,N_7985,N_7874);
or U8498 (N_8498,N_7756,N_7628);
nand U8499 (N_8499,N_7936,N_7786);
and U8500 (N_8500,N_8267,N_8495);
or U8501 (N_8501,N_8165,N_8381);
nor U8502 (N_8502,N_8323,N_8168);
nor U8503 (N_8503,N_8042,N_8390);
nor U8504 (N_8504,N_8286,N_8287);
and U8505 (N_8505,N_8280,N_8407);
nor U8506 (N_8506,N_8230,N_8318);
nand U8507 (N_8507,N_8021,N_8458);
and U8508 (N_8508,N_8160,N_8484);
or U8509 (N_8509,N_8462,N_8327);
and U8510 (N_8510,N_8232,N_8223);
or U8511 (N_8511,N_8054,N_8186);
or U8512 (N_8512,N_8245,N_8029);
or U8513 (N_8513,N_8356,N_8215);
nand U8514 (N_8514,N_8459,N_8337);
xnor U8515 (N_8515,N_8040,N_8308);
and U8516 (N_8516,N_8293,N_8285);
nor U8517 (N_8517,N_8465,N_8094);
or U8518 (N_8518,N_8480,N_8218);
xor U8519 (N_8519,N_8136,N_8005);
nor U8520 (N_8520,N_8247,N_8248);
xnor U8521 (N_8521,N_8176,N_8027);
and U8522 (N_8522,N_8310,N_8170);
and U8523 (N_8523,N_8262,N_8277);
and U8524 (N_8524,N_8139,N_8039);
xnor U8525 (N_8525,N_8055,N_8460);
or U8526 (N_8526,N_8350,N_8103);
nand U8527 (N_8527,N_8061,N_8034);
nand U8528 (N_8528,N_8111,N_8379);
and U8529 (N_8529,N_8288,N_8031);
nor U8530 (N_8530,N_8414,N_8433);
and U8531 (N_8531,N_8290,N_8071);
nand U8532 (N_8532,N_8208,N_8331);
and U8533 (N_8533,N_8131,N_8257);
nand U8534 (N_8534,N_8162,N_8332);
or U8535 (N_8535,N_8197,N_8043);
or U8536 (N_8536,N_8070,N_8169);
and U8537 (N_8537,N_8231,N_8254);
nand U8538 (N_8538,N_8341,N_8187);
nor U8539 (N_8539,N_8069,N_8454);
nor U8540 (N_8540,N_8493,N_8251);
nor U8541 (N_8541,N_8431,N_8423);
nor U8542 (N_8542,N_8046,N_8082);
and U8543 (N_8543,N_8296,N_8463);
nand U8544 (N_8544,N_8173,N_8372);
or U8545 (N_8545,N_8011,N_8305);
or U8546 (N_8546,N_8084,N_8199);
and U8547 (N_8547,N_8498,N_8491);
nand U8548 (N_8548,N_8122,N_8451);
or U8549 (N_8549,N_8348,N_8175);
nand U8550 (N_8550,N_8096,N_8393);
nor U8551 (N_8551,N_8126,N_8066);
nand U8552 (N_8552,N_8406,N_8338);
or U8553 (N_8553,N_8201,N_8079);
nor U8554 (N_8554,N_8319,N_8185);
and U8555 (N_8555,N_8353,N_8425);
or U8556 (N_8556,N_8018,N_8118);
or U8557 (N_8557,N_8456,N_8032);
and U8558 (N_8558,N_8282,N_8453);
nor U8559 (N_8559,N_8488,N_8291);
or U8560 (N_8560,N_8204,N_8249);
or U8561 (N_8561,N_8374,N_8067);
nand U8562 (N_8562,N_8107,N_8142);
or U8563 (N_8563,N_8345,N_8150);
xnor U8564 (N_8564,N_8256,N_8426);
xnor U8565 (N_8565,N_8057,N_8229);
or U8566 (N_8566,N_8302,N_8261);
and U8567 (N_8567,N_8134,N_8216);
or U8568 (N_8568,N_8238,N_8263);
nand U8569 (N_8569,N_8106,N_8252);
nor U8570 (N_8570,N_8387,N_8284);
nand U8571 (N_8571,N_8470,N_8474);
nor U8572 (N_8572,N_8236,N_8158);
nor U8573 (N_8573,N_8065,N_8340);
and U8574 (N_8574,N_8482,N_8146);
and U8575 (N_8575,N_8129,N_8472);
nor U8576 (N_8576,N_8152,N_8014);
nor U8577 (N_8577,N_8001,N_8481);
or U8578 (N_8578,N_8428,N_8127);
or U8579 (N_8579,N_8479,N_8396);
nand U8580 (N_8580,N_8113,N_8360);
nand U8581 (N_8581,N_8343,N_8050);
or U8582 (N_8582,N_8329,N_8378);
or U8583 (N_8583,N_8313,N_8270);
and U8584 (N_8584,N_8295,N_8279);
and U8585 (N_8585,N_8367,N_8221);
nor U8586 (N_8586,N_8172,N_8135);
nand U8587 (N_8587,N_8346,N_8240);
nand U8588 (N_8588,N_8321,N_8294);
xor U8589 (N_8589,N_8220,N_8180);
nor U8590 (N_8590,N_8022,N_8468);
nor U8591 (N_8591,N_8417,N_8427);
nand U8592 (N_8592,N_8016,N_8097);
or U8593 (N_8593,N_8044,N_8408);
and U8594 (N_8594,N_8085,N_8354);
nor U8595 (N_8595,N_8081,N_8355);
and U8596 (N_8596,N_8391,N_8405);
nor U8597 (N_8597,N_8063,N_8325);
nand U8598 (N_8598,N_8369,N_8148);
nor U8599 (N_8599,N_8342,N_8475);
nor U8600 (N_8600,N_8365,N_8086);
nand U8601 (N_8601,N_8492,N_8362);
and U8602 (N_8602,N_8322,N_8382);
nor U8603 (N_8603,N_8435,N_8411);
nand U8604 (N_8604,N_8429,N_8174);
or U8605 (N_8605,N_8078,N_8080);
and U8606 (N_8606,N_8226,N_8147);
xor U8607 (N_8607,N_8120,N_8141);
or U8608 (N_8608,N_8476,N_8398);
nand U8609 (N_8609,N_8415,N_8010);
or U8610 (N_8610,N_8167,N_8455);
or U8611 (N_8611,N_8289,N_8225);
and U8612 (N_8612,N_8181,N_8447);
nand U8613 (N_8613,N_8161,N_8105);
nand U8614 (N_8614,N_8190,N_8335);
nor U8615 (N_8615,N_8006,N_8183);
nor U8616 (N_8616,N_8166,N_8243);
nor U8617 (N_8617,N_8452,N_8219);
and U8618 (N_8618,N_8351,N_8145);
or U8619 (N_8619,N_8448,N_8009);
and U8620 (N_8620,N_8274,N_8269);
or U8621 (N_8621,N_8073,N_8133);
nor U8622 (N_8622,N_8485,N_8149);
xor U8623 (N_8623,N_8317,N_8089);
or U8624 (N_8624,N_8442,N_8138);
nand U8625 (N_8625,N_8487,N_8403);
or U8626 (N_8626,N_8059,N_8217);
nor U8627 (N_8627,N_8051,N_8316);
or U8628 (N_8628,N_8058,N_8047);
nor U8629 (N_8629,N_8164,N_8189);
nand U8630 (N_8630,N_8036,N_8401);
nor U8631 (N_8631,N_8400,N_8376);
and U8632 (N_8632,N_8191,N_8076);
nor U8633 (N_8633,N_8074,N_8203);
nand U8634 (N_8634,N_8037,N_8099);
nand U8635 (N_8635,N_8206,N_8483);
nand U8636 (N_8636,N_8281,N_8114);
and U8637 (N_8637,N_8330,N_8012);
or U8638 (N_8638,N_8392,N_8438);
and U8639 (N_8639,N_8091,N_8064);
nand U8640 (N_8640,N_8297,N_8366);
and U8641 (N_8641,N_8213,N_8024);
nand U8642 (N_8642,N_8496,N_8469);
or U8643 (N_8643,N_8449,N_8466);
nand U8644 (N_8644,N_8121,N_8163);
nand U8645 (N_8645,N_8422,N_8110);
nand U8646 (N_8646,N_8095,N_8464);
and U8647 (N_8647,N_8041,N_8389);
nand U8648 (N_8648,N_8184,N_8062);
and U8649 (N_8649,N_8312,N_8090);
nand U8650 (N_8650,N_8259,N_8368);
and U8651 (N_8651,N_8344,N_8255);
nand U8652 (N_8652,N_8273,N_8013);
nor U8653 (N_8653,N_8380,N_8478);
nand U8654 (N_8654,N_8373,N_8384);
and U8655 (N_8655,N_8371,N_8497);
nand U8656 (N_8656,N_8068,N_8052);
nor U8657 (N_8657,N_8446,N_8304);
nand U8658 (N_8658,N_8471,N_8177);
and U8659 (N_8659,N_8477,N_8056);
nor U8660 (N_8660,N_8420,N_8359);
nand U8661 (N_8661,N_8399,N_8241);
nand U8662 (N_8662,N_8019,N_8416);
and U8663 (N_8663,N_8233,N_8087);
nor U8664 (N_8664,N_8275,N_8404);
or U8665 (N_8665,N_8140,N_8198);
nand U8666 (N_8666,N_8048,N_8315);
and U8667 (N_8667,N_8212,N_8250);
nor U8668 (N_8668,N_8494,N_8123);
nand U8669 (N_8669,N_8002,N_8130);
nor U8670 (N_8670,N_8083,N_8156);
or U8671 (N_8671,N_8265,N_8410);
nand U8672 (N_8672,N_8104,N_8413);
or U8673 (N_8673,N_8260,N_8409);
or U8674 (N_8674,N_8457,N_8178);
xor U8675 (N_8675,N_8112,N_8195);
xor U8676 (N_8676,N_8473,N_8109);
nand U8677 (N_8677,N_8300,N_8108);
nand U8678 (N_8678,N_8124,N_8008);
or U8679 (N_8679,N_8128,N_8125);
and U8680 (N_8680,N_8347,N_8314);
and U8681 (N_8681,N_8276,N_8361);
and U8682 (N_8682,N_8102,N_8307);
nand U8683 (N_8683,N_8301,N_8182);
nand U8684 (N_8684,N_8100,N_8194);
or U8685 (N_8685,N_8437,N_8349);
nand U8686 (N_8686,N_8193,N_8264);
or U8687 (N_8687,N_8119,N_8222);
nor U8688 (N_8688,N_8358,N_8038);
and U8689 (N_8689,N_8278,N_8003);
nand U8690 (N_8690,N_8000,N_8271);
nor U8691 (N_8691,N_8299,N_8490);
and U8692 (N_8692,N_8434,N_8443);
and U8693 (N_8693,N_8244,N_8432);
and U8694 (N_8694,N_8210,N_8025);
or U8695 (N_8695,N_8283,N_8418);
and U8696 (N_8696,N_8385,N_8072);
nor U8697 (N_8697,N_8430,N_8336);
nand U8698 (N_8698,N_8035,N_8364);
nand U8699 (N_8699,N_8049,N_8098);
and U8700 (N_8700,N_8386,N_8309);
or U8701 (N_8701,N_8444,N_8157);
and U8702 (N_8702,N_8196,N_8214);
and U8703 (N_8703,N_8028,N_8151);
nor U8704 (N_8704,N_8440,N_8155);
nand U8705 (N_8705,N_8395,N_8394);
nor U8706 (N_8706,N_8154,N_8441);
and U8707 (N_8707,N_8397,N_8227);
nand U8708 (N_8708,N_8328,N_8333);
or U8709 (N_8709,N_8421,N_8235);
and U8710 (N_8710,N_8388,N_8357);
nor U8711 (N_8711,N_8377,N_8137);
and U8712 (N_8712,N_8311,N_8306);
and U8713 (N_8713,N_8334,N_8489);
and U8714 (N_8714,N_8298,N_8320);
nand U8715 (N_8715,N_8159,N_8412);
or U8716 (N_8716,N_8253,N_8060);
nor U8717 (N_8717,N_8188,N_8303);
or U8718 (N_8718,N_8339,N_8266);
nor U8719 (N_8719,N_8101,N_8026);
nand U8720 (N_8720,N_8211,N_8153);
nor U8721 (N_8721,N_8007,N_8326);
or U8722 (N_8722,N_8017,N_8023);
nor U8723 (N_8723,N_8205,N_8088);
and U8724 (N_8724,N_8207,N_8171);
nand U8725 (N_8725,N_8239,N_8092);
or U8726 (N_8726,N_8292,N_8116);
nor U8727 (N_8727,N_8436,N_8424);
nand U8728 (N_8728,N_8053,N_8192);
or U8729 (N_8729,N_8209,N_8499);
nand U8730 (N_8730,N_8237,N_8224);
or U8731 (N_8731,N_8445,N_8200);
and U8732 (N_8732,N_8370,N_8045);
nand U8733 (N_8733,N_8144,N_8461);
or U8734 (N_8734,N_8093,N_8077);
or U8735 (N_8735,N_8115,N_8033);
nand U8736 (N_8736,N_8202,N_8179);
and U8737 (N_8737,N_8228,N_8467);
nor U8738 (N_8738,N_8450,N_8004);
nand U8739 (N_8739,N_8132,N_8439);
and U8740 (N_8740,N_8246,N_8324);
and U8741 (N_8741,N_8020,N_8117);
or U8742 (N_8742,N_8242,N_8363);
nand U8743 (N_8743,N_8352,N_8383);
nand U8744 (N_8744,N_8402,N_8272);
or U8745 (N_8745,N_8486,N_8030);
nor U8746 (N_8746,N_8375,N_8419);
nand U8747 (N_8747,N_8143,N_8075);
nand U8748 (N_8748,N_8015,N_8234);
nor U8749 (N_8749,N_8258,N_8268);
and U8750 (N_8750,N_8365,N_8037);
nand U8751 (N_8751,N_8018,N_8023);
or U8752 (N_8752,N_8413,N_8406);
and U8753 (N_8753,N_8045,N_8005);
or U8754 (N_8754,N_8467,N_8226);
nand U8755 (N_8755,N_8264,N_8036);
nor U8756 (N_8756,N_8434,N_8202);
or U8757 (N_8757,N_8251,N_8358);
xnor U8758 (N_8758,N_8157,N_8064);
and U8759 (N_8759,N_8008,N_8062);
and U8760 (N_8760,N_8264,N_8173);
and U8761 (N_8761,N_8314,N_8208);
nand U8762 (N_8762,N_8349,N_8104);
or U8763 (N_8763,N_8378,N_8320);
nor U8764 (N_8764,N_8425,N_8209);
nand U8765 (N_8765,N_8181,N_8331);
and U8766 (N_8766,N_8003,N_8268);
nand U8767 (N_8767,N_8414,N_8439);
or U8768 (N_8768,N_8155,N_8397);
or U8769 (N_8769,N_8372,N_8415);
nor U8770 (N_8770,N_8457,N_8408);
and U8771 (N_8771,N_8225,N_8103);
nand U8772 (N_8772,N_8244,N_8347);
or U8773 (N_8773,N_8402,N_8354);
nor U8774 (N_8774,N_8427,N_8433);
and U8775 (N_8775,N_8021,N_8221);
xor U8776 (N_8776,N_8149,N_8318);
nor U8777 (N_8777,N_8197,N_8031);
nor U8778 (N_8778,N_8424,N_8016);
nand U8779 (N_8779,N_8083,N_8122);
xor U8780 (N_8780,N_8140,N_8404);
nand U8781 (N_8781,N_8461,N_8400);
nand U8782 (N_8782,N_8190,N_8379);
and U8783 (N_8783,N_8203,N_8447);
nand U8784 (N_8784,N_8362,N_8163);
and U8785 (N_8785,N_8267,N_8087);
and U8786 (N_8786,N_8407,N_8117);
and U8787 (N_8787,N_8451,N_8060);
nor U8788 (N_8788,N_8266,N_8085);
nand U8789 (N_8789,N_8168,N_8288);
nor U8790 (N_8790,N_8411,N_8015);
nor U8791 (N_8791,N_8276,N_8309);
nor U8792 (N_8792,N_8358,N_8227);
nand U8793 (N_8793,N_8409,N_8287);
nor U8794 (N_8794,N_8155,N_8308);
or U8795 (N_8795,N_8265,N_8420);
nand U8796 (N_8796,N_8231,N_8040);
and U8797 (N_8797,N_8305,N_8006);
nor U8798 (N_8798,N_8353,N_8287);
nor U8799 (N_8799,N_8078,N_8073);
and U8800 (N_8800,N_8233,N_8138);
or U8801 (N_8801,N_8468,N_8173);
nand U8802 (N_8802,N_8342,N_8307);
nand U8803 (N_8803,N_8083,N_8415);
nand U8804 (N_8804,N_8174,N_8004);
nand U8805 (N_8805,N_8094,N_8368);
nor U8806 (N_8806,N_8209,N_8136);
nand U8807 (N_8807,N_8458,N_8181);
nor U8808 (N_8808,N_8133,N_8070);
or U8809 (N_8809,N_8173,N_8459);
and U8810 (N_8810,N_8341,N_8318);
nor U8811 (N_8811,N_8021,N_8299);
or U8812 (N_8812,N_8120,N_8442);
nor U8813 (N_8813,N_8356,N_8261);
nand U8814 (N_8814,N_8080,N_8325);
nand U8815 (N_8815,N_8364,N_8204);
or U8816 (N_8816,N_8296,N_8491);
nand U8817 (N_8817,N_8198,N_8099);
nor U8818 (N_8818,N_8087,N_8265);
and U8819 (N_8819,N_8091,N_8214);
nand U8820 (N_8820,N_8159,N_8434);
nor U8821 (N_8821,N_8273,N_8203);
or U8822 (N_8822,N_8219,N_8062);
and U8823 (N_8823,N_8247,N_8237);
or U8824 (N_8824,N_8375,N_8217);
and U8825 (N_8825,N_8496,N_8079);
and U8826 (N_8826,N_8359,N_8102);
or U8827 (N_8827,N_8229,N_8393);
nor U8828 (N_8828,N_8025,N_8278);
and U8829 (N_8829,N_8010,N_8405);
nand U8830 (N_8830,N_8416,N_8470);
nand U8831 (N_8831,N_8127,N_8311);
nand U8832 (N_8832,N_8099,N_8174);
or U8833 (N_8833,N_8082,N_8391);
nand U8834 (N_8834,N_8335,N_8148);
or U8835 (N_8835,N_8365,N_8293);
nand U8836 (N_8836,N_8454,N_8403);
or U8837 (N_8837,N_8378,N_8274);
and U8838 (N_8838,N_8186,N_8242);
or U8839 (N_8839,N_8187,N_8205);
nand U8840 (N_8840,N_8404,N_8322);
or U8841 (N_8841,N_8278,N_8200);
nand U8842 (N_8842,N_8064,N_8376);
and U8843 (N_8843,N_8228,N_8143);
nand U8844 (N_8844,N_8490,N_8053);
or U8845 (N_8845,N_8400,N_8012);
or U8846 (N_8846,N_8084,N_8432);
nand U8847 (N_8847,N_8390,N_8148);
nor U8848 (N_8848,N_8368,N_8388);
nor U8849 (N_8849,N_8326,N_8064);
nor U8850 (N_8850,N_8382,N_8105);
nand U8851 (N_8851,N_8202,N_8306);
and U8852 (N_8852,N_8153,N_8471);
and U8853 (N_8853,N_8420,N_8181);
xor U8854 (N_8854,N_8495,N_8049);
and U8855 (N_8855,N_8191,N_8034);
nand U8856 (N_8856,N_8315,N_8058);
and U8857 (N_8857,N_8440,N_8495);
and U8858 (N_8858,N_8492,N_8132);
xnor U8859 (N_8859,N_8102,N_8430);
and U8860 (N_8860,N_8067,N_8336);
nor U8861 (N_8861,N_8166,N_8396);
and U8862 (N_8862,N_8276,N_8415);
nand U8863 (N_8863,N_8461,N_8342);
or U8864 (N_8864,N_8172,N_8187);
nand U8865 (N_8865,N_8400,N_8492);
nor U8866 (N_8866,N_8075,N_8299);
or U8867 (N_8867,N_8426,N_8295);
nor U8868 (N_8868,N_8163,N_8412);
nand U8869 (N_8869,N_8408,N_8497);
nand U8870 (N_8870,N_8159,N_8498);
nor U8871 (N_8871,N_8178,N_8485);
or U8872 (N_8872,N_8360,N_8464);
xor U8873 (N_8873,N_8055,N_8383);
nor U8874 (N_8874,N_8439,N_8297);
nor U8875 (N_8875,N_8238,N_8388);
or U8876 (N_8876,N_8353,N_8380);
and U8877 (N_8877,N_8083,N_8392);
nor U8878 (N_8878,N_8047,N_8368);
nand U8879 (N_8879,N_8064,N_8189);
nor U8880 (N_8880,N_8232,N_8070);
and U8881 (N_8881,N_8189,N_8469);
nand U8882 (N_8882,N_8401,N_8120);
nand U8883 (N_8883,N_8432,N_8144);
nand U8884 (N_8884,N_8155,N_8175);
nor U8885 (N_8885,N_8451,N_8004);
nand U8886 (N_8886,N_8016,N_8416);
or U8887 (N_8887,N_8364,N_8107);
nand U8888 (N_8888,N_8114,N_8001);
nor U8889 (N_8889,N_8459,N_8156);
and U8890 (N_8890,N_8088,N_8443);
nor U8891 (N_8891,N_8281,N_8003);
nor U8892 (N_8892,N_8457,N_8354);
nand U8893 (N_8893,N_8209,N_8140);
nand U8894 (N_8894,N_8096,N_8163);
and U8895 (N_8895,N_8013,N_8462);
and U8896 (N_8896,N_8486,N_8238);
and U8897 (N_8897,N_8495,N_8427);
or U8898 (N_8898,N_8158,N_8089);
and U8899 (N_8899,N_8343,N_8285);
nand U8900 (N_8900,N_8328,N_8019);
nor U8901 (N_8901,N_8493,N_8213);
nor U8902 (N_8902,N_8257,N_8340);
nand U8903 (N_8903,N_8499,N_8186);
and U8904 (N_8904,N_8350,N_8401);
nand U8905 (N_8905,N_8019,N_8471);
nor U8906 (N_8906,N_8130,N_8458);
nand U8907 (N_8907,N_8404,N_8095);
xor U8908 (N_8908,N_8388,N_8253);
nor U8909 (N_8909,N_8129,N_8268);
xor U8910 (N_8910,N_8166,N_8220);
or U8911 (N_8911,N_8370,N_8199);
and U8912 (N_8912,N_8263,N_8411);
nor U8913 (N_8913,N_8083,N_8151);
or U8914 (N_8914,N_8011,N_8185);
nor U8915 (N_8915,N_8038,N_8329);
nor U8916 (N_8916,N_8050,N_8280);
nor U8917 (N_8917,N_8297,N_8160);
nand U8918 (N_8918,N_8068,N_8256);
nor U8919 (N_8919,N_8259,N_8000);
or U8920 (N_8920,N_8126,N_8093);
nor U8921 (N_8921,N_8272,N_8106);
nor U8922 (N_8922,N_8277,N_8372);
and U8923 (N_8923,N_8282,N_8156);
nand U8924 (N_8924,N_8151,N_8173);
and U8925 (N_8925,N_8144,N_8189);
or U8926 (N_8926,N_8048,N_8217);
nor U8927 (N_8927,N_8004,N_8270);
xor U8928 (N_8928,N_8143,N_8312);
nor U8929 (N_8929,N_8363,N_8283);
or U8930 (N_8930,N_8431,N_8140);
nor U8931 (N_8931,N_8093,N_8413);
and U8932 (N_8932,N_8307,N_8365);
nand U8933 (N_8933,N_8088,N_8305);
nor U8934 (N_8934,N_8237,N_8104);
nor U8935 (N_8935,N_8300,N_8001);
or U8936 (N_8936,N_8103,N_8116);
nand U8937 (N_8937,N_8074,N_8235);
or U8938 (N_8938,N_8479,N_8254);
and U8939 (N_8939,N_8150,N_8297);
or U8940 (N_8940,N_8444,N_8320);
nor U8941 (N_8941,N_8342,N_8030);
or U8942 (N_8942,N_8488,N_8496);
and U8943 (N_8943,N_8400,N_8368);
nand U8944 (N_8944,N_8137,N_8132);
and U8945 (N_8945,N_8049,N_8063);
nand U8946 (N_8946,N_8146,N_8340);
nor U8947 (N_8947,N_8113,N_8425);
nor U8948 (N_8948,N_8353,N_8272);
and U8949 (N_8949,N_8227,N_8278);
and U8950 (N_8950,N_8285,N_8023);
and U8951 (N_8951,N_8337,N_8119);
nand U8952 (N_8952,N_8457,N_8058);
nor U8953 (N_8953,N_8134,N_8465);
or U8954 (N_8954,N_8160,N_8231);
nor U8955 (N_8955,N_8248,N_8438);
or U8956 (N_8956,N_8025,N_8452);
and U8957 (N_8957,N_8357,N_8249);
nor U8958 (N_8958,N_8171,N_8342);
and U8959 (N_8959,N_8005,N_8105);
or U8960 (N_8960,N_8128,N_8449);
and U8961 (N_8961,N_8248,N_8250);
nand U8962 (N_8962,N_8470,N_8349);
nand U8963 (N_8963,N_8379,N_8478);
and U8964 (N_8964,N_8433,N_8237);
and U8965 (N_8965,N_8260,N_8375);
or U8966 (N_8966,N_8064,N_8065);
or U8967 (N_8967,N_8294,N_8182);
nor U8968 (N_8968,N_8435,N_8231);
and U8969 (N_8969,N_8043,N_8497);
nor U8970 (N_8970,N_8127,N_8335);
or U8971 (N_8971,N_8407,N_8146);
or U8972 (N_8972,N_8131,N_8254);
or U8973 (N_8973,N_8052,N_8343);
or U8974 (N_8974,N_8109,N_8181);
nor U8975 (N_8975,N_8150,N_8018);
and U8976 (N_8976,N_8163,N_8465);
nand U8977 (N_8977,N_8136,N_8116);
or U8978 (N_8978,N_8075,N_8395);
nand U8979 (N_8979,N_8179,N_8379);
and U8980 (N_8980,N_8180,N_8436);
and U8981 (N_8981,N_8190,N_8226);
nor U8982 (N_8982,N_8232,N_8230);
or U8983 (N_8983,N_8097,N_8407);
and U8984 (N_8984,N_8153,N_8042);
nand U8985 (N_8985,N_8151,N_8348);
and U8986 (N_8986,N_8478,N_8262);
and U8987 (N_8987,N_8201,N_8388);
and U8988 (N_8988,N_8156,N_8197);
nand U8989 (N_8989,N_8277,N_8028);
nand U8990 (N_8990,N_8254,N_8347);
and U8991 (N_8991,N_8024,N_8090);
nor U8992 (N_8992,N_8083,N_8225);
nand U8993 (N_8993,N_8026,N_8134);
and U8994 (N_8994,N_8461,N_8281);
nor U8995 (N_8995,N_8495,N_8101);
and U8996 (N_8996,N_8160,N_8343);
and U8997 (N_8997,N_8469,N_8433);
nand U8998 (N_8998,N_8217,N_8433);
nand U8999 (N_8999,N_8344,N_8476);
or U9000 (N_9000,N_8585,N_8998);
and U9001 (N_9001,N_8602,N_8644);
nand U9002 (N_9002,N_8765,N_8774);
and U9003 (N_9003,N_8769,N_8626);
and U9004 (N_9004,N_8559,N_8944);
or U9005 (N_9005,N_8713,N_8825);
and U9006 (N_9006,N_8537,N_8505);
and U9007 (N_9007,N_8996,N_8962);
nand U9008 (N_9008,N_8588,N_8987);
xnor U9009 (N_9009,N_8797,N_8854);
or U9010 (N_9010,N_8690,N_8591);
nand U9011 (N_9011,N_8930,N_8880);
and U9012 (N_9012,N_8530,N_8587);
or U9013 (N_9013,N_8824,N_8540);
and U9014 (N_9014,N_8711,N_8871);
nand U9015 (N_9015,N_8958,N_8868);
nand U9016 (N_9016,N_8936,N_8803);
or U9017 (N_9017,N_8574,N_8771);
nand U9018 (N_9018,N_8781,N_8541);
nor U9019 (N_9019,N_8980,N_8667);
and U9020 (N_9020,N_8673,N_8934);
nor U9021 (N_9021,N_8633,N_8568);
and U9022 (N_9022,N_8580,N_8865);
and U9023 (N_9023,N_8560,N_8504);
and U9024 (N_9024,N_8828,N_8897);
and U9025 (N_9025,N_8977,N_8782);
or U9026 (N_9026,N_8992,N_8800);
nand U9027 (N_9027,N_8669,N_8903);
nand U9028 (N_9028,N_8918,N_8635);
nor U9029 (N_9029,N_8816,N_8881);
nand U9030 (N_9030,N_8570,N_8584);
or U9031 (N_9031,N_8773,N_8957);
or U9032 (N_9032,N_8755,N_8834);
nor U9033 (N_9033,N_8916,N_8524);
or U9034 (N_9034,N_8658,N_8567);
nor U9035 (N_9035,N_8843,N_8659);
and U9036 (N_9036,N_8613,N_8728);
or U9037 (N_9037,N_8627,N_8564);
or U9038 (N_9038,N_8717,N_8748);
nor U9039 (N_9039,N_8656,N_8666);
nand U9040 (N_9040,N_8820,N_8883);
nor U9041 (N_9041,N_8786,N_8718);
and U9042 (N_9042,N_8946,N_8842);
and U9043 (N_9043,N_8978,N_8510);
nor U9044 (N_9044,N_8573,N_8877);
nand U9045 (N_9045,N_8864,N_8698);
nor U9046 (N_9046,N_8508,N_8623);
and U9047 (N_9047,N_8988,N_8790);
and U9048 (N_9048,N_8625,N_8583);
nor U9049 (N_9049,N_8721,N_8604);
and U9050 (N_9050,N_8960,N_8549);
or U9051 (N_9051,N_8768,N_8831);
or U9052 (N_9052,N_8506,N_8931);
and U9053 (N_9053,N_8566,N_8575);
and U9054 (N_9054,N_8716,N_8735);
nor U9055 (N_9055,N_8527,N_8821);
nor U9056 (N_9056,N_8745,N_8503);
nor U9057 (N_9057,N_8684,N_8744);
and U9058 (N_9058,N_8961,N_8696);
and U9059 (N_9059,N_8724,N_8655);
nor U9060 (N_9060,N_8914,N_8875);
and U9061 (N_9061,N_8873,N_8789);
nand U9062 (N_9062,N_8902,N_8925);
or U9063 (N_9063,N_8979,N_8565);
or U9064 (N_9064,N_8787,N_8529);
or U9065 (N_9065,N_8911,N_8579);
nor U9066 (N_9066,N_8596,N_8830);
nor U9067 (N_9067,N_8929,N_8872);
and U9068 (N_9068,N_8521,N_8867);
xor U9069 (N_9069,N_8894,N_8976);
or U9070 (N_9070,N_8576,N_8533);
and U9071 (N_9071,N_8795,N_8829);
nand U9072 (N_9072,N_8994,N_8664);
nand U9073 (N_9073,N_8746,N_8532);
or U9074 (N_9074,N_8545,N_8837);
nor U9075 (N_9075,N_8599,N_8955);
nand U9076 (N_9076,N_8554,N_8823);
and U9077 (N_9077,N_8594,N_8523);
nand U9078 (N_9078,N_8600,N_8685);
and U9079 (N_9079,N_8766,N_8813);
or U9080 (N_9080,N_8704,N_8692);
or U9081 (N_9081,N_8542,N_8725);
nor U9082 (N_9082,N_8901,N_8762);
or U9083 (N_9083,N_8997,N_8796);
or U9084 (N_9084,N_8722,N_8593);
nor U9085 (N_9085,N_8513,N_8905);
or U9086 (N_9086,N_8663,N_8952);
and U9087 (N_9087,N_8848,N_8528);
and U9088 (N_9088,N_8779,N_8741);
nand U9089 (N_9089,N_8851,N_8544);
and U9090 (N_9090,N_8706,N_8642);
nor U9091 (N_9091,N_8743,N_8687);
or U9092 (N_9092,N_8967,N_8556);
or U9093 (N_9093,N_8707,N_8665);
and U9094 (N_9094,N_8647,N_8749);
nor U9095 (N_9095,N_8863,N_8753);
or U9096 (N_9096,N_8882,N_8720);
xor U9097 (N_9097,N_8712,N_8668);
nor U9098 (N_9098,N_8947,N_8640);
nand U9099 (N_9099,N_8595,N_8920);
or U9100 (N_9100,N_8900,N_8534);
nor U9101 (N_9101,N_8853,N_8557);
nor U9102 (N_9102,N_8605,N_8630);
nand U9103 (N_9103,N_8509,N_8689);
nor U9104 (N_9104,N_8592,N_8926);
nor U9105 (N_9105,N_8700,N_8709);
nand U9106 (N_9106,N_8857,N_8637);
nand U9107 (N_9107,N_8632,N_8995);
nor U9108 (N_9108,N_8798,N_8730);
or U9109 (N_9109,N_8971,N_8833);
or U9110 (N_9110,N_8518,N_8912);
and U9111 (N_9111,N_8699,N_8631);
nor U9112 (N_9112,N_8986,N_8535);
or U9113 (N_9113,N_8906,N_8758);
or U9114 (N_9114,N_8981,N_8909);
and U9115 (N_9115,N_8688,N_8806);
and U9116 (N_9116,N_8693,N_8571);
nand U9117 (N_9117,N_8661,N_8609);
nand U9118 (N_9118,N_8791,N_8512);
and U9119 (N_9119,N_8694,N_8740);
or U9120 (N_9120,N_8968,N_8859);
and U9121 (N_9121,N_8680,N_8569);
and U9122 (N_9122,N_8616,N_8650);
nand U9123 (N_9123,N_8678,N_8835);
nor U9124 (N_9124,N_8984,N_8836);
or U9125 (N_9125,N_8672,N_8641);
and U9126 (N_9126,N_8841,N_8671);
nor U9127 (N_9127,N_8899,N_8775);
or U9128 (N_9128,N_8818,N_8852);
or U9129 (N_9129,N_8840,N_8869);
nand U9130 (N_9130,N_8870,N_8783);
nand U9131 (N_9131,N_8990,N_8941);
nor U9132 (N_9132,N_8860,N_8621);
xor U9133 (N_9133,N_8683,N_8607);
or U9134 (N_9134,N_8586,N_8921);
nand U9135 (N_9135,N_8752,N_8951);
or U9136 (N_9136,N_8547,N_8638);
nor U9137 (N_9137,N_8785,N_8959);
and U9138 (N_9138,N_8674,N_8618);
nor U9139 (N_9139,N_8913,N_8691);
nand U9140 (N_9140,N_8731,N_8759);
nor U9141 (N_9141,N_8924,N_8653);
nor U9142 (N_9142,N_8582,N_8525);
nor U9143 (N_9143,N_8938,N_8855);
nor U9144 (N_9144,N_8892,N_8629);
nor U9145 (N_9145,N_8727,N_8969);
nand U9146 (N_9146,N_8636,N_8817);
nor U9147 (N_9147,N_8793,N_8608);
nand U9148 (N_9148,N_8945,N_8708);
or U9149 (N_9149,N_8612,N_8760);
or U9150 (N_9150,N_8670,N_8756);
and U9151 (N_9151,N_8891,N_8932);
nor U9152 (N_9152,N_8705,N_8732);
nand U9153 (N_9153,N_8888,N_8606);
nand U9154 (N_9154,N_8874,N_8948);
or U9155 (N_9155,N_8927,N_8526);
nor U9156 (N_9156,N_8826,N_8895);
or U9157 (N_9157,N_8839,N_8845);
nand U9158 (N_9158,N_8879,N_8832);
and U9159 (N_9159,N_8890,N_8770);
nor U9160 (N_9160,N_8729,N_8723);
or U9161 (N_9161,N_8738,N_8651);
or U9162 (N_9162,N_8907,N_8522);
xor U9163 (N_9163,N_8624,N_8531);
and U9164 (N_9164,N_8937,N_8622);
nand U9165 (N_9165,N_8514,N_8811);
nor U9166 (N_9166,N_8861,N_8778);
nor U9167 (N_9167,N_8776,N_8750);
and U9168 (N_9168,N_8819,N_8598);
nand U9169 (N_9169,N_8939,N_8703);
and U9170 (N_9170,N_8886,N_8849);
nor U9171 (N_9171,N_8767,N_8502);
nand U9172 (N_9172,N_8993,N_8884);
and U9173 (N_9173,N_8646,N_8772);
nand U9174 (N_9174,N_8763,N_8846);
nand U9175 (N_9175,N_8515,N_8517);
and U9176 (N_9176,N_8546,N_8808);
nor U9177 (N_9177,N_8619,N_8974);
nor U9178 (N_9178,N_8910,N_8536);
nand U9179 (N_9179,N_8949,N_8634);
and U9180 (N_9180,N_8966,N_8815);
nand U9181 (N_9181,N_8983,N_8652);
nand U9182 (N_9182,N_8539,N_8876);
and U9183 (N_9183,N_8553,N_8681);
nand U9184 (N_9184,N_8838,N_8964);
nand U9185 (N_9185,N_8590,N_8878);
and U9186 (N_9186,N_8558,N_8615);
or U9187 (N_9187,N_8885,N_8989);
or U9188 (N_9188,N_8581,N_8543);
and U9189 (N_9189,N_8904,N_8889);
nor U9190 (N_9190,N_8887,N_8552);
nand U9191 (N_9191,N_8784,N_8610);
and U9192 (N_9192,N_8617,N_8601);
and U9193 (N_9193,N_8548,N_8950);
nor U9194 (N_9194,N_8847,N_8827);
xnor U9195 (N_9195,N_8561,N_8734);
nor U9196 (N_9196,N_8963,N_8810);
nor U9197 (N_9197,N_8917,N_8919);
xor U9198 (N_9198,N_8614,N_8603);
and U9199 (N_9199,N_8679,N_8991);
and U9200 (N_9200,N_8893,N_8751);
or U9201 (N_9201,N_8942,N_8597);
and U9202 (N_9202,N_8715,N_8799);
nor U9203 (N_9203,N_8858,N_8501);
and U9204 (N_9204,N_8737,N_8923);
nand U9205 (N_9205,N_8620,N_8682);
xor U9206 (N_9206,N_8520,N_8922);
or U9207 (N_9207,N_8611,N_8982);
or U9208 (N_9208,N_8754,N_8896);
or U9209 (N_9209,N_8676,N_8805);
nand U9210 (N_9210,N_8714,N_8578);
and U9211 (N_9211,N_8649,N_8500);
xnor U9212 (N_9212,N_8965,N_8757);
nor U9213 (N_9213,N_8654,N_8710);
or U9214 (N_9214,N_8516,N_8777);
nand U9215 (N_9215,N_8742,N_8804);
and U9216 (N_9216,N_8985,N_8538);
nor U9217 (N_9217,N_8662,N_8563);
nand U9218 (N_9218,N_8643,N_8850);
or U9219 (N_9219,N_8577,N_8954);
and U9220 (N_9220,N_8761,N_8695);
and U9221 (N_9221,N_8589,N_8511);
and U9222 (N_9222,N_8807,N_8788);
nand U9223 (N_9223,N_8719,N_8628);
or U9224 (N_9224,N_8792,N_8822);
nor U9225 (N_9225,N_8507,N_8551);
and U9226 (N_9226,N_8908,N_8702);
xor U9227 (N_9227,N_8519,N_8972);
or U9228 (N_9228,N_8733,N_8736);
and U9229 (N_9229,N_8802,N_8956);
or U9230 (N_9230,N_8801,N_8677);
nor U9231 (N_9231,N_8856,N_8814);
or U9232 (N_9232,N_8898,N_8975);
nand U9233 (N_9233,N_8675,N_8747);
nor U9234 (N_9234,N_8726,N_8970);
and U9235 (N_9235,N_8697,N_8928);
nor U9236 (N_9236,N_8794,N_8555);
nor U9237 (N_9237,N_8648,N_8812);
xor U9238 (N_9238,N_8953,N_8562);
nor U9239 (N_9239,N_8645,N_8844);
or U9240 (N_9240,N_8639,N_8660);
nand U9241 (N_9241,N_8933,N_8943);
or U9242 (N_9242,N_8809,N_8657);
nor U9243 (N_9243,N_8686,N_8935);
nand U9244 (N_9244,N_8940,N_8866);
and U9245 (N_9245,N_8780,N_8915);
nand U9246 (N_9246,N_8550,N_8973);
or U9247 (N_9247,N_8739,N_8999);
nand U9248 (N_9248,N_8862,N_8764);
and U9249 (N_9249,N_8701,N_8572);
or U9250 (N_9250,N_8577,N_8568);
or U9251 (N_9251,N_8584,N_8589);
and U9252 (N_9252,N_8805,N_8518);
and U9253 (N_9253,N_8970,N_8641);
and U9254 (N_9254,N_8801,N_8949);
and U9255 (N_9255,N_8758,N_8820);
and U9256 (N_9256,N_8935,N_8884);
and U9257 (N_9257,N_8774,N_8869);
nand U9258 (N_9258,N_8953,N_8661);
nor U9259 (N_9259,N_8586,N_8666);
nand U9260 (N_9260,N_8998,N_8652);
or U9261 (N_9261,N_8816,N_8723);
nand U9262 (N_9262,N_8973,N_8853);
nand U9263 (N_9263,N_8874,N_8713);
or U9264 (N_9264,N_8948,N_8981);
nand U9265 (N_9265,N_8951,N_8648);
or U9266 (N_9266,N_8694,N_8519);
nor U9267 (N_9267,N_8869,N_8834);
nand U9268 (N_9268,N_8576,N_8813);
nand U9269 (N_9269,N_8947,N_8882);
or U9270 (N_9270,N_8608,N_8625);
nand U9271 (N_9271,N_8526,N_8895);
nor U9272 (N_9272,N_8694,N_8800);
or U9273 (N_9273,N_8686,N_8642);
and U9274 (N_9274,N_8785,N_8665);
nand U9275 (N_9275,N_8512,N_8864);
and U9276 (N_9276,N_8797,N_8910);
or U9277 (N_9277,N_8731,N_8623);
nand U9278 (N_9278,N_8514,N_8666);
and U9279 (N_9279,N_8594,N_8981);
and U9280 (N_9280,N_8887,N_8516);
nor U9281 (N_9281,N_8963,N_8610);
nand U9282 (N_9282,N_8636,N_8539);
or U9283 (N_9283,N_8564,N_8529);
or U9284 (N_9284,N_8701,N_8942);
nor U9285 (N_9285,N_8882,N_8546);
nand U9286 (N_9286,N_8694,N_8677);
nand U9287 (N_9287,N_8928,N_8748);
nor U9288 (N_9288,N_8546,N_8781);
and U9289 (N_9289,N_8594,N_8813);
nor U9290 (N_9290,N_8558,N_8985);
and U9291 (N_9291,N_8617,N_8918);
nand U9292 (N_9292,N_8526,N_8510);
and U9293 (N_9293,N_8744,N_8516);
nor U9294 (N_9294,N_8742,N_8625);
and U9295 (N_9295,N_8733,N_8577);
and U9296 (N_9296,N_8549,N_8801);
or U9297 (N_9297,N_8711,N_8685);
or U9298 (N_9298,N_8726,N_8730);
or U9299 (N_9299,N_8558,N_8832);
and U9300 (N_9300,N_8924,N_8692);
nor U9301 (N_9301,N_8933,N_8931);
or U9302 (N_9302,N_8982,N_8521);
nor U9303 (N_9303,N_8992,N_8753);
or U9304 (N_9304,N_8668,N_8733);
nand U9305 (N_9305,N_8996,N_8747);
or U9306 (N_9306,N_8527,N_8928);
and U9307 (N_9307,N_8652,N_8798);
nand U9308 (N_9308,N_8784,N_8749);
or U9309 (N_9309,N_8526,N_8634);
nor U9310 (N_9310,N_8890,N_8977);
nor U9311 (N_9311,N_8534,N_8915);
xnor U9312 (N_9312,N_8589,N_8644);
nand U9313 (N_9313,N_8737,N_8841);
nor U9314 (N_9314,N_8681,N_8705);
nand U9315 (N_9315,N_8965,N_8986);
nand U9316 (N_9316,N_8641,N_8546);
and U9317 (N_9317,N_8577,N_8929);
nand U9318 (N_9318,N_8817,N_8920);
nand U9319 (N_9319,N_8808,N_8681);
nand U9320 (N_9320,N_8792,N_8800);
nor U9321 (N_9321,N_8684,N_8839);
and U9322 (N_9322,N_8737,N_8624);
and U9323 (N_9323,N_8790,N_8861);
or U9324 (N_9324,N_8533,N_8831);
nand U9325 (N_9325,N_8530,N_8563);
nor U9326 (N_9326,N_8527,N_8856);
or U9327 (N_9327,N_8624,N_8943);
nand U9328 (N_9328,N_8727,N_8565);
nor U9329 (N_9329,N_8753,N_8903);
or U9330 (N_9330,N_8964,N_8646);
and U9331 (N_9331,N_8847,N_8944);
and U9332 (N_9332,N_8969,N_8627);
or U9333 (N_9333,N_8910,N_8858);
nor U9334 (N_9334,N_8937,N_8676);
or U9335 (N_9335,N_8974,N_8844);
and U9336 (N_9336,N_8805,N_8964);
and U9337 (N_9337,N_8619,N_8881);
nor U9338 (N_9338,N_8898,N_8873);
nand U9339 (N_9339,N_8806,N_8937);
and U9340 (N_9340,N_8723,N_8732);
nand U9341 (N_9341,N_8778,N_8993);
nor U9342 (N_9342,N_8918,N_8989);
or U9343 (N_9343,N_8659,N_8800);
and U9344 (N_9344,N_8587,N_8970);
nand U9345 (N_9345,N_8748,N_8653);
nor U9346 (N_9346,N_8889,N_8764);
nor U9347 (N_9347,N_8674,N_8876);
nor U9348 (N_9348,N_8610,N_8677);
nand U9349 (N_9349,N_8982,N_8518);
nor U9350 (N_9350,N_8986,N_8888);
nand U9351 (N_9351,N_8604,N_8968);
xnor U9352 (N_9352,N_8916,N_8743);
nand U9353 (N_9353,N_8522,N_8595);
nor U9354 (N_9354,N_8695,N_8555);
and U9355 (N_9355,N_8685,N_8799);
and U9356 (N_9356,N_8555,N_8885);
nand U9357 (N_9357,N_8680,N_8736);
or U9358 (N_9358,N_8686,N_8794);
or U9359 (N_9359,N_8984,N_8824);
and U9360 (N_9360,N_8608,N_8756);
and U9361 (N_9361,N_8848,N_8772);
or U9362 (N_9362,N_8512,N_8511);
nor U9363 (N_9363,N_8831,N_8794);
or U9364 (N_9364,N_8973,N_8582);
and U9365 (N_9365,N_8612,N_8871);
and U9366 (N_9366,N_8674,N_8991);
nand U9367 (N_9367,N_8528,N_8907);
nor U9368 (N_9368,N_8961,N_8634);
or U9369 (N_9369,N_8678,N_8946);
nor U9370 (N_9370,N_8899,N_8543);
and U9371 (N_9371,N_8665,N_8542);
and U9372 (N_9372,N_8520,N_8554);
nor U9373 (N_9373,N_8966,N_8670);
nand U9374 (N_9374,N_8930,N_8865);
and U9375 (N_9375,N_8578,N_8770);
and U9376 (N_9376,N_8753,N_8981);
nand U9377 (N_9377,N_8951,N_8631);
and U9378 (N_9378,N_8502,N_8935);
or U9379 (N_9379,N_8561,N_8546);
and U9380 (N_9380,N_8708,N_8764);
and U9381 (N_9381,N_8956,N_8877);
nor U9382 (N_9382,N_8803,N_8545);
nor U9383 (N_9383,N_8624,N_8557);
nor U9384 (N_9384,N_8836,N_8730);
and U9385 (N_9385,N_8696,N_8656);
nand U9386 (N_9386,N_8600,N_8815);
or U9387 (N_9387,N_8941,N_8821);
nor U9388 (N_9388,N_8685,N_8939);
and U9389 (N_9389,N_8960,N_8599);
or U9390 (N_9390,N_8605,N_8834);
and U9391 (N_9391,N_8575,N_8601);
nand U9392 (N_9392,N_8847,N_8739);
and U9393 (N_9393,N_8779,N_8660);
and U9394 (N_9394,N_8731,N_8514);
nand U9395 (N_9395,N_8653,N_8801);
nor U9396 (N_9396,N_8665,N_8768);
nand U9397 (N_9397,N_8852,N_8675);
nor U9398 (N_9398,N_8553,N_8505);
nor U9399 (N_9399,N_8769,N_8564);
and U9400 (N_9400,N_8553,N_8701);
nand U9401 (N_9401,N_8663,N_8546);
nor U9402 (N_9402,N_8919,N_8912);
and U9403 (N_9403,N_8774,N_8788);
or U9404 (N_9404,N_8928,N_8630);
and U9405 (N_9405,N_8862,N_8938);
nand U9406 (N_9406,N_8631,N_8736);
nand U9407 (N_9407,N_8619,N_8836);
and U9408 (N_9408,N_8719,N_8663);
and U9409 (N_9409,N_8880,N_8659);
nor U9410 (N_9410,N_8697,N_8593);
nor U9411 (N_9411,N_8771,N_8617);
and U9412 (N_9412,N_8591,N_8820);
and U9413 (N_9413,N_8838,N_8683);
or U9414 (N_9414,N_8805,N_8662);
nor U9415 (N_9415,N_8704,N_8753);
and U9416 (N_9416,N_8718,N_8957);
nor U9417 (N_9417,N_8531,N_8647);
and U9418 (N_9418,N_8786,N_8956);
nor U9419 (N_9419,N_8662,N_8886);
and U9420 (N_9420,N_8991,N_8970);
or U9421 (N_9421,N_8870,N_8954);
nor U9422 (N_9422,N_8806,N_8739);
nand U9423 (N_9423,N_8853,N_8948);
nor U9424 (N_9424,N_8605,N_8870);
or U9425 (N_9425,N_8603,N_8822);
and U9426 (N_9426,N_8547,N_8633);
nand U9427 (N_9427,N_8537,N_8722);
nor U9428 (N_9428,N_8529,N_8868);
nor U9429 (N_9429,N_8958,N_8659);
or U9430 (N_9430,N_8511,N_8770);
nor U9431 (N_9431,N_8717,N_8811);
xnor U9432 (N_9432,N_8659,N_8551);
and U9433 (N_9433,N_8882,N_8725);
nand U9434 (N_9434,N_8903,N_8714);
or U9435 (N_9435,N_8632,N_8670);
nor U9436 (N_9436,N_8751,N_8909);
and U9437 (N_9437,N_8746,N_8718);
or U9438 (N_9438,N_8584,N_8577);
or U9439 (N_9439,N_8761,N_8581);
and U9440 (N_9440,N_8871,N_8570);
nor U9441 (N_9441,N_8585,N_8822);
nand U9442 (N_9442,N_8985,N_8596);
nand U9443 (N_9443,N_8578,N_8911);
and U9444 (N_9444,N_8564,N_8947);
or U9445 (N_9445,N_8663,N_8875);
or U9446 (N_9446,N_8782,N_8687);
and U9447 (N_9447,N_8961,N_8542);
and U9448 (N_9448,N_8897,N_8636);
nand U9449 (N_9449,N_8957,N_8566);
nor U9450 (N_9450,N_8992,N_8944);
or U9451 (N_9451,N_8577,N_8519);
nor U9452 (N_9452,N_8679,N_8802);
and U9453 (N_9453,N_8534,N_8975);
and U9454 (N_9454,N_8754,N_8977);
nand U9455 (N_9455,N_8796,N_8760);
nand U9456 (N_9456,N_8937,N_8961);
nor U9457 (N_9457,N_8613,N_8554);
or U9458 (N_9458,N_8892,N_8855);
and U9459 (N_9459,N_8813,N_8633);
nand U9460 (N_9460,N_8884,N_8540);
nand U9461 (N_9461,N_8888,N_8926);
and U9462 (N_9462,N_8848,N_8992);
and U9463 (N_9463,N_8931,N_8950);
and U9464 (N_9464,N_8562,N_8522);
nand U9465 (N_9465,N_8874,N_8518);
and U9466 (N_9466,N_8962,N_8586);
or U9467 (N_9467,N_8536,N_8950);
or U9468 (N_9468,N_8862,N_8750);
nor U9469 (N_9469,N_8602,N_8964);
nand U9470 (N_9470,N_8555,N_8761);
and U9471 (N_9471,N_8888,N_8798);
nor U9472 (N_9472,N_8557,N_8546);
and U9473 (N_9473,N_8513,N_8720);
xnor U9474 (N_9474,N_8848,N_8939);
xnor U9475 (N_9475,N_8892,N_8891);
nand U9476 (N_9476,N_8691,N_8755);
and U9477 (N_9477,N_8702,N_8637);
or U9478 (N_9478,N_8861,N_8710);
nor U9479 (N_9479,N_8993,N_8550);
nand U9480 (N_9480,N_8583,N_8862);
nand U9481 (N_9481,N_8643,N_8707);
or U9482 (N_9482,N_8510,N_8940);
or U9483 (N_9483,N_8778,N_8832);
nand U9484 (N_9484,N_8524,N_8637);
nor U9485 (N_9485,N_8621,N_8892);
nand U9486 (N_9486,N_8951,N_8957);
nor U9487 (N_9487,N_8655,N_8641);
nor U9488 (N_9488,N_8903,N_8628);
nor U9489 (N_9489,N_8599,N_8941);
or U9490 (N_9490,N_8745,N_8690);
nor U9491 (N_9491,N_8946,N_8868);
or U9492 (N_9492,N_8878,N_8807);
nor U9493 (N_9493,N_8581,N_8606);
nand U9494 (N_9494,N_8838,N_8927);
nor U9495 (N_9495,N_8617,N_8800);
nand U9496 (N_9496,N_8857,N_8635);
and U9497 (N_9497,N_8964,N_8690);
and U9498 (N_9498,N_8788,N_8983);
or U9499 (N_9499,N_8641,N_8759);
nor U9500 (N_9500,N_9170,N_9099);
or U9501 (N_9501,N_9047,N_9145);
xnor U9502 (N_9502,N_9207,N_9000);
and U9503 (N_9503,N_9299,N_9013);
nor U9504 (N_9504,N_9187,N_9021);
nor U9505 (N_9505,N_9004,N_9141);
or U9506 (N_9506,N_9331,N_9418);
and U9507 (N_9507,N_9345,N_9442);
or U9508 (N_9508,N_9180,N_9045);
nand U9509 (N_9509,N_9341,N_9464);
nand U9510 (N_9510,N_9355,N_9243);
nor U9511 (N_9511,N_9071,N_9001);
nand U9512 (N_9512,N_9318,N_9356);
or U9513 (N_9513,N_9289,N_9194);
nand U9514 (N_9514,N_9451,N_9075);
nor U9515 (N_9515,N_9053,N_9157);
and U9516 (N_9516,N_9490,N_9192);
nor U9517 (N_9517,N_9292,N_9330);
and U9518 (N_9518,N_9465,N_9260);
nand U9519 (N_9519,N_9395,N_9242);
nand U9520 (N_9520,N_9279,N_9064);
nor U9521 (N_9521,N_9264,N_9386);
xnor U9522 (N_9522,N_9143,N_9486);
nor U9523 (N_9523,N_9156,N_9246);
nand U9524 (N_9524,N_9237,N_9044);
nor U9525 (N_9525,N_9029,N_9009);
nor U9526 (N_9526,N_9440,N_9425);
or U9527 (N_9527,N_9365,N_9480);
nand U9528 (N_9528,N_9074,N_9436);
nor U9529 (N_9529,N_9091,N_9140);
and U9530 (N_9530,N_9032,N_9148);
nand U9531 (N_9531,N_9107,N_9487);
or U9532 (N_9532,N_9063,N_9399);
or U9533 (N_9533,N_9234,N_9322);
nand U9534 (N_9534,N_9470,N_9460);
nand U9535 (N_9535,N_9108,N_9411);
nor U9536 (N_9536,N_9372,N_9041);
and U9537 (N_9537,N_9058,N_9094);
xnor U9538 (N_9538,N_9300,N_9153);
and U9539 (N_9539,N_9495,N_9446);
and U9540 (N_9540,N_9132,N_9133);
nor U9541 (N_9541,N_9334,N_9068);
or U9542 (N_9542,N_9188,N_9408);
nand U9543 (N_9543,N_9383,N_9097);
and U9544 (N_9544,N_9200,N_9251);
or U9545 (N_9545,N_9127,N_9118);
or U9546 (N_9546,N_9171,N_9422);
and U9547 (N_9547,N_9202,N_9239);
or U9548 (N_9548,N_9102,N_9311);
nor U9549 (N_9549,N_9271,N_9296);
nand U9550 (N_9550,N_9364,N_9326);
nand U9551 (N_9551,N_9429,N_9423);
nand U9552 (N_9552,N_9317,N_9381);
or U9553 (N_9553,N_9445,N_9070);
or U9554 (N_9554,N_9169,N_9481);
and U9555 (N_9555,N_9206,N_9201);
and U9556 (N_9556,N_9407,N_9252);
or U9557 (N_9557,N_9217,N_9349);
or U9558 (N_9558,N_9011,N_9024);
or U9559 (N_9559,N_9266,N_9054);
nor U9560 (N_9560,N_9461,N_9453);
nand U9561 (N_9561,N_9120,N_9427);
nand U9562 (N_9562,N_9276,N_9052);
and U9563 (N_9563,N_9337,N_9485);
or U9564 (N_9564,N_9366,N_9295);
or U9565 (N_9565,N_9125,N_9073);
and U9566 (N_9566,N_9240,N_9496);
nand U9567 (N_9567,N_9497,N_9190);
nand U9568 (N_9568,N_9413,N_9402);
nor U9569 (N_9569,N_9459,N_9406);
or U9570 (N_9570,N_9484,N_9473);
nor U9571 (N_9571,N_9443,N_9166);
or U9572 (N_9572,N_9403,N_9377);
nand U9573 (N_9573,N_9247,N_9104);
or U9574 (N_9574,N_9215,N_9475);
or U9575 (N_9575,N_9455,N_9163);
or U9576 (N_9576,N_9034,N_9335);
nor U9577 (N_9577,N_9297,N_9343);
nor U9578 (N_9578,N_9249,N_9112);
nor U9579 (N_9579,N_9250,N_9085);
or U9580 (N_9580,N_9288,N_9134);
nor U9581 (N_9581,N_9059,N_9286);
and U9582 (N_9582,N_9109,N_9439);
and U9583 (N_9583,N_9283,N_9208);
nand U9584 (N_9584,N_9030,N_9430);
nor U9585 (N_9585,N_9081,N_9493);
nor U9586 (N_9586,N_9361,N_9060);
and U9587 (N_9587,N_9352,N_9105);
nor U9588 (N_9588,N_9347,N_9437);
or U9589 (N_9589,N_9110,N_9261);
xor U9590 (N_9590,N_9198,N_9020);
nor U9591 (N_9591,N_9280,N_9274);
nand U9592 (N_9592,N_9348,N_9161);
or U9593 (N_9593,N_9150,N_9272);
nor U9594 (N_9594,N_9010,N_9390);
nor U9595 (N_9595,N_9375,N_9195);
and U9596 (N_9596,N_9137,N_9216);
and U9597 (N_9597,N_9253,N_9426);
and U9598 (N_9598,N_9088,N_9412);
nand U9599 (N_9599,N_9327,N_9328);
or U9600 (N_9600,N_9441,N_9444);
nor U9601 (N_9601,N_9373,N_9257);
nor U9602 (N_9602,N_9363,N_9244);
nor U9603 (N_9603,N_9062,N_9093);
nor U9604 (N_9604,N_9391,N_9087);
and U9605 (N_9605,N_9231,N_9040);
nand U9606 (N_9606,N_9357,N_9478);
xor U9607 (N_9607,N_9397,N_9432);
or U9608 (N_9608,N_9498,N_9165);
and U9609 (N_9609,N_9016,N_9258);
or U9610 (N_9610,N_9138,N_9056);
or U9611 (N_9611,N_9111,N_9065);
nand U9612 (N_9612,N_9154,N_9100);
and U9613 (N_9613,N_9398,N_9218);
or U9614 (N_9614,N_9126,N_9305);
and U9615 (N_9615,N_9462,N_9226);
and U9616 (N_9616,N_9387,N_9232);
or U9617 (N_9617,N_9342,N_9284);
nand U9618 (N_9618,N_9026,N_9124);
nor U9619 (N_9619,N_9416,N_9002);
and U9620 (N_9620,N_9324,N_9368);
or U9621 (N_9621,N_9128,N_9015);
nand U9622 (N_9622,N_9066,N_9410);
and U9623 (N_9623,N_9420,N_9076);
and U9624 (N_9624,N_9467,N_9101);
and U9625 (N_9625,N_9479,N_9259);
and U9626 (N_9626,N_9491,N_9433);
nand U9627 (N_9627,N_9483,N_9113);
nor U9628 (N_9628,N_9230,N_9119);
or U9629 (N_9629,N_9354,N_9472);
and U9630 (N_9630,N_9362,N_9293);
xor U9631 (N_9631,N_9008,N_9400);
nor U9632 (N_9632,N_9316,N_9499);
or U9633 (N_9633,N_9175,N_9277);
and U9634 (N_9634,N_9262,N_9417);
nand U9635 (N_9635,N_9458,N_9130);
or U9636 (N_9636,N_9454,N_9431);
nand U9637 (N_9637,N_9023,N_9067);
nand U9638 (N_9638,N_9248,N_9035);
and U9639 (N_9639,N_9199,N_9302);
or U9640 (N_9640,N_9312,N_9351);
nor U9641 (N_9641,N_9256,N_9409);
or U9642 (N_9642,N_9042,N_9307);
nand U9643 (N_9643,N_9007,N_9338);
nor U9644 (N_9644,N_9103,N_9254);
or U9645 (N_9645,N_9304,N_9350);
nand U9646 (N_9646,N_9382,N_9376);
nand U9647 (N_9647,N_9344,N_9469);
and U9648 (N_9648,N_9017,N_9235);
nor U9649 (N_9649,N_9203,N_9340);
nand U9650 (N_9650,N_9421,N_9384);
and U9651 (N_9651,N_9336,N_9168);
or U9652 (N_9652,N_9438,N_9268);
or U9653 (N_9653,N_9072,N_9018);
or U9654 (N_9654,N_9401,N_9329);
nor U9655 (N_9655,N_9178,N_9414);
nand U9656 (N_9656,N_9083,N_9313);
nor U9657 (N_9657,N_9255,N_9028);
and U9658 (N_9658,N_9014,N_9167);
nor U9659 (N_9659,N_9049,N_9131);
or U9660 (N_9660,N_9214,N_9039);
nand U9661 (N_9661,N_9385,N_9323);
nor U9662 (N_9662,N_9003,N_9048);
and U9663 (N_9663,N_9222,N_9419);
or U9664 (N_9664,N_9489,N_9238);
nor U9665 (N_9665,N_9358,N_9471);
or U9666 (N_9666,N_9077,N_9050);
nand U9667 (N_9667,N_9055,N_9123);
and U9668 (N_9668,N_9378,N_9424);
nand U9669 (N_9669,N_9474,N_9212);
nor U9670 (N_9670,N_9314,N_9122);
or U9671 (N_9671,N_9213,N_9449);
or U9672 (N_9672,N_9396,N_9078);
xor U9673 (N_9673,N_9183,N_9227);
and U9674 (N_9674,N_9172,N_9144);
nor U9675 (N_9675,N_9339,N_9151);
or U9676 (N_9676,N_9321,N_9281);
nand U9677 (N_9677,N_9448,N_9135);
or U9678 (N_9678,N_9309,N_9275);
nor U9679 (N_9679,N_9245,N_9006);
nor U9680 (N_9680,N_9388,N_9452);
and U9681 (N_9681,N_9147,N_9228);
nor U9682 (N_9682,N_9086,N_9415);
nor U9683 (N_9683,N_9179,N_9273);
or U9684 (N_9684,N_9174,N_9359);
nand U9685 (N_9685,N_9158,N_9369);
and U9686 (N_9686,N_9488,N_9038);
xor U9687 (N_9687,N_9160,N_9267);
nor U9688 (N_9688,N_9265,N_9193);
or U9689 (N_9689,N_9333,N_9456);
nand U9690 (N_9690,N_9374,N_9155);
xnor U9691 (N_9691,N_9176,N_9082);
or U9692 (N_9692,N_9114,N_9005);
nand U9693 (N_9693,N_9033,N_9080);
or U9694 (N_9694,N_9241,N_9450);
nor U9695 (N_9695,N_9301,N_9325);
and U9696 (N_9696,N_9173,N_9159);
and U9697 (N_9697,N_9142,N_9186);
nand U9698 (N_9698,N_9308,N_9098);
nand U9699 (N_9699,N_9084,N_9079);
nand U9700 (N_9700,N_9463,N_9146);
and U9701 (N_9701,N_9303,N_9294);
or U9702 (N_9702,N_9036,N_9221);
nand U9703 (N_9703,N_9298,N_9468);
and U9704 (N_9704,N_9181,N_9270);
nor U9705 (N_9705,N_9177,N_9057);
and U9706 (N_9706,N_9022,N_9404);
or U9707 (N_9707,N_9037,N_9184);
nor U9708 (N_9708,N_9428,N_9164);
nor U9709 (N_9709,N_9152,N_9319);
nand U9710 (N_9710,N_9116,N_9353);
nor U9711 (N_9711,N_9220,N_9457);
and U9712 (N_9712,N_9061,N_9019);
or U9713 (N_9713,N_9371,N_9482);
or U9714 (N_9714,N_9209,N_9129);
nor U9715 (N_9715,N_9043,N_9393);
or U9716 (N_9716,N_9466,N_9185);
nand U9717 (N_9717,N_9278,N_9405);
nand U9718 (N_9718,N_9106,N_9394);
nand U9719 (N_9719,N_9315,N_9392);
or U9720 (N_9720,N_9306,N_9204);
or U9721 (N_9721,N_9263,N_9370);
or U9722 (N_9722,N_9291,N_9379);
nand U9723 (N_9723,N_9096,N_9121);
and U9724 (N_9724,N_9477,N_9092);
nor U9725 (N_9725,N_9282,N_9090);
or U9726 (N_9726,N_9225,N_9117);
nand U9727 (N_9727,N_9290,N_9434);
nand U9728 (N_9728,N_9027,N_9389);
or U9729 (N_9729,N_9447,N_9360);
nor U9730 (N_9730,N_9051,N_9205);
nand U9731 (N_9731,N_9211,N_9189);
or U9732 (N_9732,N_9191,N_9162);
and U9733 (N_9733,N_9380,N_9223);
nor U9734 (N_9734,N_9285,N_9046);
and U9735 (N_9735,N_9139,N_9320);
and U9736 (N_9736,N_9115,N_9196);
or U9737 (N_9737,N_9224,N_9476);
or U9738 (N_9738,N_9089,N_9136);
nand U9739 (N_9739,N_9367,N_9149);
or U9740 (N_9740,N_9210,N_9492);
nand U9741 (N_9741,N_9269,N_9219);
nor U9742 (N_9742,N_9346,N_9332);
nor U9743 (N_9743,N_9031,N_9287);
or U9744 (N_9744,N_9310,N_9095);
nor U9745 (N_9745,N_9494,N_9229);
or U9746 (N_9746,N_9182,N_9069);
or U9747 (N_9747,N_9025,N_9197);
and U9748 (N_9748,N_9012,N_9233);
nor U9749 (N_9749,N_9435,N_9236);
nor U9750 (N_9750,N_9406,N_9219);
nor U9751 (N_9751,N_9237,N_9228);
and U9752 (N_9752,N_9478,N_9214);
nand U9753 (N_9753,N_9206,N_9451);
nand U9754 (N_9754,N_9121,N_9156);
nor U9755 (N_9755,N_9458,N_9411);
nand U9756 (N_9756,N_9086,N_9129);
or U9757 (N_9757,N_9288,N_9082);
and U9758 (N_9758,N_9157,N_9018);
nand U9759 (N_9759,N_9385,N_9465);
or U9760 (N_9760,N_9220,N_9476);
nor U9761 (N_9761,N_9043,N_9141);
nand U9762 (N_9762,N_9438,N_9144);
xor U9763 (N_9763,N_9038,N_9271);
nor U9764 (N_9764,N_9151,N_9280);
nand U9765 (N_9765,N_9055,N_9259);
nor U9766 (N_9766,N_9165,N_9236);
and U9767 (N_9767,N_9419,N_9390);
or U9768 (N_9768,N_9006,N_9162);
and U9769 (N_9769,N_9097,N_9046);
nor U9770 (N_9770,N_9222,N_9104);
and U9771 (N_9771,N_9001,N_9410);
and U9772 (N_9772,N_9006,N_9414);
nor U9773 (N_9773,N_9427,N_9124);
nand U9774 (N_9774,N_9470,N_9208);
nand U9775 (N_9775,N_9320,N_9238);
nor U9776 (N_9776,N_9066,N_9163);
or U9777 (N_9777,N_9133,N_9408);
or U9778 (N_9778,N_9355,N_9429);
nor U9779 (N_9779,N_9349,N_9073);
nand U9780 (N_9780,N_9189,N_9018);
nor U9781 (N_9781,N_9281,N_9140);
nand U9782 (N_9782,N_9009,N_9470);
xor U9783 (N_9783,N_9493,N_9242);
and U9784 (N_9784,N_9171,N_9457);
and U9785 (N_9785,N_9404,N_9080);
and U9786 (N_9786,N_9378,N_9333);
nor U9787 (N_9787,N_9439,N_9381);
or U9788 (N_9788,N_9481,N_9086);
and U9789 (N_9789,N_9368,N_9338);
or U9790 (N_9790,N_9194,N_9116);
nand U9791 (N_9791,N_9336,N_9466);
and U9792 (N_9792,N_9244,N_9364);
and U9793 (N_9793,N_9306,N_9130);
or U9794 (N_9794,N_9398,N_9028);
xnor U9795 (N_9795,N_9347,N_9244);
or U9796 (N_9796,N_9006,N_9032);
or U9797 (N_9797,N_9026,N_9497);
and U9798 (N_9798,N_9220,N_9165);
and U9799 (N_9799,N_9006,N_9163);
and U9800 (N_9800,N_9158,N_9040);
nor U9801 (N_9801,N_9400,N_9167);
and U9802 (N_9802,N_9196,N_9124);
and U9803 (N_9803,N_9438,N_9352);
or U9804 (N_9804,N_9192,N_9186);
nand U9805 (N_9805,N_9107,N_9242);
nand U9806 (N_9806,N_9432,N_9052);
nor U9807 (N_9807,N_9167,N_9298);
xor U9808 (N_9808,N_9375,N_9029);
nor U9809 (N_9809,N_9471,N_9082);
nor U9810 (N_9810,N_9180,N_9290);
nor U9811 (N_9811,N_9157,N_9411);
nor U9812 (N_9812,N_9234,N_9293);
or U9813 (N_9813,N_9206,N_9384);
xnor U9814 (N_9814,N_9005,N_9379);
and U9815 (N_9815,N_9085,N_9195);
and U9816 (N_9816,N_9315,N_9472);
or U9817 (N_9817,N_9140,N_9176);
nor U9818 (N_9818,N_9261,N_9150);
and U9819 (N_9819,N_9291,N_9342);
or U9820 (N_9820,N_9469,N_9108);
nor U9821 (N_9821,N_9016,N_9072);
and U9822 (N_9822,N_9340,N_9286);
and U9823 (N_9823,N_9158,N_9118);
or U9824 (N_9824,N_9175,N_9186);
or U9825 (N_9825,N_9388,N_9464);
nor U9826 (N_9826,N_9320,N_9031);
nor U9827 (N_9827,N_9053,N_9479);
or U9828 (N_9828,N_9005,N_9154);
and U9829 (N_9829,N_9312,N_9338);
and U9830 (N_9830,N_9327,N_9051);
and U9831 (N_9831,N_9177,N_9432);
or U9832 (N_9832,N_9486,N_9070);
nand U9833 (N_9833,N_9132,N_9490);
and U9834 (N_9834,N_9330,N_9428);
nor U9835 (N_9835,N_9356,N_9082);
nor U9836 (N_9836,N_9387,N_9386);
or U9837 (N_9837,N_9494,N_9283);
and U9838 (N_9838,N_9231,N_9335);
xor U9839 (N_9839,N_9350,N_9340);
nand U9840 (N_9840,N_9474,N_9258);
nor U9841 (N_9841,N_9206,N_9416);
nor U9842 (N_9842,N_9181,N_9429);
or U9843 (N_9843,N_9274,N_9141);
nor U9844 (N_9844,N_9022,N_9181);
nor U9845 (N_9845,N_9013,N_9380);
nor U9846 (N_9846,N_9256,N_9178);
nor U9847 (N_9847,N_9359,N_9059);
xnor U9848 (N_9848,N_9214,N_9344);
and U9849 (N_9849,N_9385,N_9414);
xor U9850 (N_9850,N_9147,N_9127);
or U9851 (N_9851,N_9357,N_9326);
and U9852 (N_9852,N_9141,N_9241);
nor U9853 (N_9853,N_9404,N_9150);
or U9854 (N_9854,N_9371,N_9305);
and U9855 (N_9855,N_9462,N_9280);
nand U9856 (N_9856,N_9344,N_9167);
or U9857 (N_9857,N_9128,N_9078);
and U9858 (N_9858,N_9228,N_9495);
and U9859 (N_9859,N_9152,N_9358);
nor U9860 (N_9860,N_9021,N_9470);
and U9861 (N_9861,N_9496,N_9459);
nand U9862 (N_9862,N_9383,N_9495);
nor U9863 (N_9863,N_9204,N_9150);
or U9864 (N_9864,N_9334,N_9091);
and U9865 (N_9865,N_9342,N_9316);
or U9866 (N_9866,N_9260,N_9258);
and U9867 (N_9867,N_9102,N_9072);
nand U9868 (N_9868,N_9081,N_9004);
or U9869 (N_9869,N_9418,N_9291);
or U9870 (N_9870,N_9212,N_9224);
nand U9871 (N_9871,N_9494,N_9188);
nor U9872 (N_9872,N_9317,N_9485);
or U9873 (N_9873,N_9243,N_9284);
or U9874 (N_9874,N_9487,N_9393);
nand U9875 (N_9875,N_9348,N_9397);
and U9876 (N_9876,N_9470,N_9330);
or U9877 (N_9877,N_9260,N_9449);
or U9878 (N_9878,N_9095,N_9181);
and U9879 (N_9879,N_9053,N_9111);
nor U9880 (N_9880,N_9181,N_9290);
nor U9881 (N_9881,N_9020,N_9154);
nor U9882 (N_9882,N_9118,N_9354);
and U9883 (N_9883,N_9455,N_9202);
and U9884 (N_9884,N_9243,N_9408);
nor U9885 (N_9885,N_9481,N_9020);
nor U9886 (N_9886,N_9397,N_9453);
and U9887 (N_9887,N_9184,N_9253);
nand U9888 (N_9888,N_9189,N_9325);
nand U9889 (N_9889,N_9367,N_9433);
nand U9890 (N_9890,N_9025,N_9392);
nand U9891 (N_9891,N_9026,N_9498);
or U9892 (N_9892,N_9462,N_9497);
and U9893 (N_9893,N_9120,N_9360);
nand U9894 (N_9894,N_9345,N_9287);
nor U9895 (N_9895,N_9488,N_9349);
nor U9896 (N_9896,N_9112,N_9493);
nand U9897 (N_9897,N_9257,N_9322);
nor U9898 (N_9898,N_9150,N_9361);
nor U9899 (N_9899,N_9491,N_9471);
nor U9900 (N_9900,N_9310,N_9460);
nor U9901 (N_9901,N_9369,N_9236);
nor U9902 (N_9902,N_9001,N_9201);
nand U9903 (N_9903,N_9040,N_9451);
nand U9904 (N_9904,N_9023,N_9224);
nand U9905 (N_9905,N_9171,N_9046);
nand U9906 (N_9906,N_9078,N_9065);
or U9907 (N_9907,N_9060,N_9167);
or U9908 (N_9908,N_9090,N_9144);
nand U9909 (N_9909,N_9025,N_9451);
nand U9910 (N_9910,N_9143,N_9116);
nand U9911 (N_9911,N_9220,N_9453);
nor U9912 (N_9912,N_9150,N_9326);
and U9913 (N_9913,N_9291,N_9127);
or U9914 (N_9914,N_9076,N_9277);
or U9915 (N_9915,N_9311,N_9189);
or U9916 (N_9916,N_9105,N_9263);
nor U9917 (N_9917,N_9453,N_9150);
nor U9918 (N_9918,N_9393,N_9297);
and U9919 (N_9919,N_9490,N_9319);
nand U9920 (N_9920,N_9191,N_9491);
nor U9921 (N_9921,N_9323,N_9307);
xor U9922 (N_9922,N_9374,N_9287);
nor U9923 (N_9923,N_9408,N_9067);
and U9924 (N_9924,N_9020,N_9223);
nand U9925 (N_9925,N_9108,N_9160);
and U9926 (N_9926,N_9252,N_9317);
nor U9927 (N_9927,N_9315,N_9385);
nand U9928 (N_9928,N_9352,N_9351);
nand U9929 (N_9929,N_9348,N_9449);
or U9930 (N_9930,N_9167,N_9284);
nor U9931 (N_9931,N_9142,N_9333);
nor U9932 (N_9932,N_9366,N_9012);
nand U9933 (N_9933,N_9455,N_9407);
nor U9934 (N_9934,N_9211,N_9421);
and U9935 (N_9935,N_9024,N_9356);
nand U9936 (N_9936,N_9145,N_9323);
and U9937 (N_9937,N_9404,N_9219);
or U9938 (N_9938,N_9087,N_9054);
nor U9939 (N_9939,N_9305,N_9143);
nor U9940 (N_9940,N_9450,N_9429);
nand U9941 (N_9941,N_9338,N_9343);
and U9942 (N_9942,N_9427,N_9332);
xnor U9943 (N_9943,N_9211,N_9031);
and U9944 (N_9944,N_9245,N_9062);
or U9945 (N_9945,N_9058,N_9494);
or U9946 (N_9946,N_9400,N_9295);
or U9947 (N_9947,N_9389,N_9397);
nand U9948 (N_9948,N_9312,N_9383);
or U9949 (N_9949,N_9138,N_9076);
and U9950 (N_9950,N_9241,N_9457);
and U9951 (N_9951,N_9247,N_9093);
nor U9952 (N_9952,N_9056,N_9454);
and U9953 (N_9953,N_9038,N_9243);
nand U9954 (N_9954,N_9130,N_9250);
nor U9955 (N_9955,N_9305,N_9081);
nand U9956 (N_9956,N_9492,N_9382);
and U9957 (N_9957,N_9169,N_9488);
nor U9958 (N_9958,N_9178,N_9014);
and U9959 (N_9959,N_9407,N_9088);
or U9960 (N_9960,N_9104,N_9170);
and U9961 (N_9961,N_9074,N_9261);
or U9962 (N_9962,N_9236,N_9163);
and U9963 (N_9963,N_9427,N_9157);
and U9964 (N_9964,N_9159,N_9224);
nor U9965 (N_9965,N_9026,N_9102);
and U9966 (N_9966,N_9060,N_9140);
nand U9967 (N_9967,N_9435,N_9474);
or U9968 (N_9968,N_9096,N_9267);
nor U9969 (N_9969,N_9400,N_9415);
nand U9970 (N_9970,N_9431,N_9102);
nand U9971 (N_9971,N_9464,N_9151);
or U9972 (N_9972,N_9297,N_9421);
or U9973 (N_9973,N_9291,N_9498);
and U9974 (N_9974,N_9496,N_9405);
or U9975 (N_9975,N_9200,N_9005);
and U9976 (N_9976,N_9272,N_9421);
and U9977 (N_9977,N_9114,N_9249);
and U9978 (N_9978,N_9031,N_9355);
nor U9979 (N_9979,N_9429,N_9125);
and U9980 (N_9980,N_9066,N_9299);
nor U9981 (N_9981,N_9335,N_9341);
xnor U9982 (N_9982,N_9444,N_9254);
or U9983 (N_9983,N_9390,N_9245);
and U9984 (N_9984,N_9275,N_9058);
nand U9985 (N_9985,N_9301,N_9140);
or U9986 (N_9986,N_9495,N_9461);
or U9987 (N_9987,N_9326,N_9081);
or U9988 (N_9988,N_9408,N_9077);
and U9989 (N_9989,N_9111,N_9228);
nor U9990 (N_9990,N_9444,N_9329);
or U9991 (N_9991,N_9009,N_9363);
or U9992 (N_9992,N_9280,N_9095);
nor U9993 (N_9993,N_9461,N_9460);
or U9994 (N_9994,N_9470,N_9035);
xnor U9995 (N_9995,N_9224,N_9005);
and U9996 (N_9996,N_9222,N_9267);
or U9997 (N_9997,N_9211,N_9011);
and U9998 (N_9998,N_9315,N_9418);
nor U9999 (N_9999,N_9360,N_9374);
and UO_0 (O_0,N_9609,N_9738);
nor UO_1 (O_1,N_9503,N_9612);
nor UO_2 (O_2,N_9945,N_9814);
and UO_3 (O_3,N_9960,N_9566);
xor UO_4 (O_4,N_9500,N_9598);
nor UO_5 (O_5,N_9619,N_9560);
or UO_6 (O_6,N_9915,N_9854);
nand UO_7 (O_7,N_9985,N_9839);
or UO_8 (O_8,N_9684,N_9623);
nor UO_9 (O_9,N_9645,N_9521);
nor UO_10 (O_10,N_9724,N_9949);
and UO_11 (O_11,N_9876,N_9926);
nor UO_12 (O_12,N_9508,N_9614);
or UO_13 (O_13,N_9996,N_9697);
nor UO_14 (O_14,N_9563,N_9950);
or UO_15 (O_15,N_9865,N_9747);
or UO_16 (O_16,N_9687,N_9533);
and UO_17 (O_17,N_9820,N_9823);
nand UO_18 (O_18,N_9727,N_9930);
nand UO_19 (O_19,N_9547,N_9743);
nor UO_20 (O_20,N_9590,N_9794);
or UO_21 (O_21,N_9752,N_9783);
or UO_22 (O_22,N_9657,N_9759);
nor UO_23 (O_23,N_9711,N_9755);
nand UO_24 (O_24,N_9976,N_9613);
and UO_25 (O_25,N_9692,N_9758);
nand UO_26 (O_26,N_9553,N_9673);
or UO_27 (O_27,N_9941,N_9957);
and UO_28 (O_28,N_9763,N_9534);
or UO_29 (O_29,N_9848,N_9837);
nor UO_30 (O_30,N_9526,N_9542);
and UO_31 (O_31,N_9603,N_9520);
and UO_32 (O_32,N_9982,N_9821);
or UO_33 (O_33,N_9658,N_9608);
nand UO_34 (O_34,N_9695,N_9517);
nor UO_35 (O_35,N_9929,N_9951);
nand UO_36 (O_36,N_9781,N_9977);
or UO_37 (O_37,N_9966,N_9723);
nand UO_38 (O_38,N_9942,N_9531);
and UO_39 (O_39,N_9884,N_9539);
nand UO_40 (O_40,N_9591,N_9923);
nand UO_41 (O_41,N_9897,N_9771);
and UO_42 (O_42,N_9796,N_9616);
or UO_43 (O_43,N_9660,N_9728);
or UO_44 (O_44,N_9548,N_9638);
nor UO_45 (O_45,N_9509,N_9979);
nor UO_46 (O_46,N_9557,N_9737);
or UO_47 (O_47,N_9644,N_9801);
or UO_48 (O_48,N_9572,N_9640);
nor UO_49 (O_49,N_9524,N_9766);
nand UO_50 (O_50,N_9819,N_9606);
nor UO_51 (O_51,N_9767,N_9733);
nand UO_52 (O_52,N_9652,N_9858);
nor UO_53 (O_53,N_9919,N_9588);
nand UO_54 (O_54,N_9883,N_9681);
and UO_55 (O_55,N_9601,N_9584);
or UO_56 (O_56,N_9561,N_9967);
nor UO_57 (O_57,N_9850,N_9842);
or UO_58 (O_58,N_9760,N_9896);
nor UO_59 (O_59,N_9739,N_9798);
and UO_60 (O_60,N_9899,N_9649);
nand UO_61 (O_61,N_9633,N_9831);
or UO_62 (O_62,N_9694,N_9643);
or UO_63 (O_63,N_9607,N_9556);
or UO_64 (O_64,N_9959,N_9732);
or UO_65 (O_65,N_9832,N_9514);
and UO_66 (O_66,N_9726,N_9902);
xnor UO_67 (O_67,N_9595,N_9834);
or UO_68 (O_68,N_9749,N_9862);
nand UO_69 (O_69,N_9506,N_9574);
or UO_70 (O_70,N_9881,N_9671);
nor UO_71 (O_71,N_9653,N_9688);
nor UO_72 (O_72,N_9800,N_9845);
xnor UO_73 (O_73,N_9825,N_9610);
or UO_74 (O_74,N_9594,N_9523);
nand UO_75 (O_75,N_9734,N_9879);
or UO_76 (O_76,N_9667,N_9946);
and UO_77 (O_77,N_9632,N_9529);
and UO_78 (O_78,N_9502,N_9750);
or UO_79 (O_79,N_9778,N_9817);
nor UO_80 (O_80,N_9700,N_9813);
nor UO_81 (O_81,N_9570,N_9736);
nor UO_82 (O_82,N_9708,N_9663);
or UO_83 (O_83,N_9824,N_9659);
nor UO_84 (O_84,N_9860,N_9559);
and UO_85 (O_85,N_9581,N_9611);
nor UO_86 (O_86,N_9804,N_9707);
or UO_87 (O_87,N_9620,N_9989);
and UO_88 (O_88,N_9628,N_9516);
and UO_89 (O_89,N_9838,N_9818);
and UO_90 (O_90,N_9893,N_9751);
nor UO_91 (O_91,N_9689,N_9669);
xor UO_92 (O_92,N_9690,N_9885);
or UO_93 (O_93,N_9940,N_9575);
or UO_94 (O_94,N_9849,N_9900);
nand UO_95 (O_95,N_9742,N_9762);
or UO_96 (O_96,N_9973,N_9605);
nand UO_97 (O_97,N_9784,N_9504);
or UO_98 (O_98,N_9868,N_9744);
nand UO_99 (O_99,N_9797,N_9933);
nor UO_100 (O_100,N_9910,N_9903);
and UO_101 (O_101,N_9599,N_9757);
nor UO_102 (O_102,N_9722,N_9866);
or UO_103 (O_103,N_9906,N_9958);
and UO_104 (O_104,N_9997,N_9725);
or UO_105 (O_105,N_9512,N_9682);
nor UO_106 (O_106,N_9835,N_9827);
and UO_107 (O_107,N_9550,N_9892);
or UO_108 (O_108,N_9585,N_9709);
nand UO_109 (O_109,N_9852,N_9920);
and UO_110 (O_110,N_9631,N_9731);
or UO_111 (O_111,N_9696,N_9676);
xnor UO_112 (O_112,N_9710,N_9537);
nor UO_113 (O_113,N_9856,N_9679);
or UO_114 (O_114,N_9935,N_9922);
and UO_115 (O_115,N_9851,N_9770);
nor UO_116 (O_116,N_9924,N_9712);
or UO_117 (O_117,N_9573,N_9768);
nor UO_118 (O_118,N_9592,N_9882);
nor UO_119 (O_119,N_9990,N_9785);
nor UO_120 (O_120,N_9639,N_9586);
or UO_121 (O_121,N_9562,N_9870);
or UO_122 (O_122,N_9986,N_9878);
or UO_123 (O_123,N_9981,N_9780);
nor UO_124 (O_124,N_9654,N_9911);
nand UO_125 (O_125,N_9863,N_9748);
or UO_126 (O_126,N_9918,N_9558);
xor UO_127 (O_127,N_9507,N_9932);
nand UO_128 (O_128,N_9543,N_9756);
nor UO_129 (O_129,N_9810,N_9861);
or UO_130 (O_130,N_9939,N_9948);
and UO_131 (O_131,N_9604,N_9706);
and UO_132 (O_132,N_9968,N_9971);
xor UO_133 (O_133,N_9917,N_9921);
or UO_134 (O_134,N_9895,N_9774);
nor UO_135 (O_135,N_9587,N_9799);
nand UO_136 (O_136,N_9955,N_9764);
and UO_137 (O_137,N_9909,N_9577);
and UO_138 (O_138,N_9872,N_9702);
and UO_139 (O_139,N_9809,N_9787);
nand UO_140 (O_140,N_9811,N_9816);
and UO_141 (O_141,N_9826,N_9907);
nand UO_142 (O_142,N_9943,N_9729);
nor UO_143 (O_143,N_9934,N_9925);
nor UO_144 (O_144,N_9735,N_9889);
nand UO_145 (O_145,N_9630,N_9532);
and UO_146 (O_146,N_9662,N_9988);
or UO_147 (O_147,N_9874,N_9969);
nand UO_148 (O_148,N_9666,N_9602);
and UO_149 (O_149,N_9741,N_9853);
nand UO_150 (O_150,N_9775,N_9754);
and UO_151 (O_151,N_9701,N_9956);
nand UO_152 (O_152,N_9627,N_9615);
and UO_153 (O_153,N_9721,N_9555);
nand UO_154 (O_154,N_9786,N_9908);
nor UO_155 (O_155,N_9991,N_9937);
and UO_156 (O_156,N_9888,N_9898);
and UO_157 (O_157,N_9664,N_9730);
nor UO_158 (O_158,N_9518,N_9536);
xor UO_159 (O_159,N_9670,N_9618);
or UO_160 (O_160,N_9546,N_9855);
or UO_161 (O_161,N_9650,N_9716);
and UO_162 (O_162,N_9843,N_9505);
nor UO_163 (O_163,N_9675,N_9719);
and UO_164 (O_164,N_9656,N_9699);
nand UO_165 (O_165,N_9636,N_9715);
and UO_166 (O_166,N_9857,N_9538);
nor UO_167 (O_167,N_9703,N_9642);
or UO_168 (O_168,N_9600,N_9978);
or UO_169 (O_169,N_9944,N_9564);
and UO_170 (O_170,N_9576,N_9962);
nand UO_171 (O_171,N_9789,N_9772);
or UO_172 (O_172,N_9873,N_9965);
or UO_173 (O_173,N_9793,N_9963);
and UO_174 (O_174,N_9720,N_9936);
and UO_175 (O_175,N_9905,N_9624);
nor UO_176 (O_176,N_9802,N_9891);
or UO_177 (O_177,N_9629,N_9769);
nor UO_178 (O_178,N_9938,N_9864);
xnor UO_179 (O_179,N_9999,N_9954);
nor UO_180 (O_180,N_9844,N_9693);
and UO_181 (O_181,N_9867,N_9931);
and UO_182 (O_182,N_9647,N_9829);
nor UO_183 (O_183,N_9880,N_9972);
and UO_184 (O_184,N_9571,N_9668);
and UO_185 (O_185,N_9519,N_9677);
nor UO_186 (O_186,N_9515,N_9705);
nand UO_187 (O_187,N_9625,N_9691);
and UO_188 (O_188,N_9527,N_9580);
and UO_189 (O_189,N_9840,N_9961);
and UO_190 (O_190,N_9953,N_9678);
and UO_191 (O_191,N_9578,N_9777);
or UO_192 (O_192,N_9554,N_9648);
nand UO_193 (O_193,N_9672,N_9589);
nand UO_194 (O_194,N_9593,N_9815);
or UO_195 (O_195,N_9745,N_9983);
nand UO_196 (O_196,N_9803,N_9773);
or UO_197 (O_197,N_9622,N_9927);
nor UO_198 (O_198,N_9788,N_9830);
nor UO_199 (O_199,N_9806,N_9822);
nand UO_200 (O_200,N_9655,N_9549);
and UO_201 (O_201,N_9782,N_9812);
nor UO_202 (O_202,N_9974,N_9987);
nor UO_203 (O_203,N_9597,N_9928);
nand UO_204 (O_204,N_9501,N_9540);
nor UO_205 (O_205,N_9952,N_9913);
nor UO_206 (O_206,N_9833,N_9565);
nor UO_207 (O_207,N_9626,N_9717);
and UO_208 (O_208,N_9846,N_9513);
and UO_209 (O_209,N_9993,N_9530);
nor UO_210 (O_210,N_9992,N_9836);
and UO_211 (O_211,N_9582,N_9621);
nor UO_212 (O_212,N_9579,N_9776);
nor UO_213 (O_213,N_9904,N_9890);
nor UO_214 (O_214,N_9901,N_9646);
and UO_215 (O_215,N_9807,N_9980);
and UO_216 (O_216,N_9552,N_9887);
and UO_217 (O_217,N_9665,N_9859);
xnor UO_218 (O_218,N_9567,N_9635);
or UO_219 (O_219,N_9686,N_9947);
and UO_220 (O_220,N_9698,N_9651);
or UO_221 (O_221,N_9975,N_9522);
or UO_222 (O_222,N_9661,N_9914);
or UO_223 (O_223,N_9994,N_9641);
nor UO_224 (O_224,N_9765,N_9718);
or UO_225 (O_225,N_9790,N_9525);
and UO_226 (O_226,N_9740,N_9791);
and UO_227 (O_227,N_9841,N_9746);
and UO_228 (O_228,N_9912,N_9637);
nor UO_229 (O_229,N_9674,N_9568);
and UO_230 (O_230,N_9528,N_9805);
and UO_231 (O_231,N_9541,N_9984);
nand UO_232 (O_232,N_9875,N_9871);
nand UO_233 (O_233,N_9869,N_9685);
nor UO_234 (O_234,N_9808,N_9535);
nand UO_235 (O_235,N_9779,N_9596);
nor UO_236 (O_236,N_9761,N_9964);
or UO_237 (O_237,N_9511,N_9970);
and UO_238 (O_238,N_9713,N_9704);
or UO_239 (O_239,N_9795,N_9998);
or UO_240 (O_240,N_9792,N_9714);
or UO_241 (O_241,N_9545,N_9894);
nor UO_242 (O_242,N_9544,N_9569);
xnor UO_243 (O_243,N_9847,N_9753);
and UO_244 (O_244,N_9683,N_9634);
nand UO_245 (O_245,N_9583,N_9510);
nand UO_246 (O_246,N_9995,N_9916);
nor UO_247 (O_247,N_9877,N_9617);
nand UO_248 (O_248,N_9886,N_9828);
and UO_249 (O_249,N_9551,N_9680);
or UO_250 (O_250,N_9743,N_9560);
and UO_251 (O_251,N_9842,N_9580);
nor UO_252 (O_252,N_9919,N_9784);
and UO_253 (O_253,N_9679,N_9960);
or UO_254 (O_254,N_9952,N_9889);
and UO_255 (O_255,N_9898,N_9523);
nor UO_256 (O_256,N_9610,N_9646);
nand UO_257 (O_257,N_9664,N_9827);
xor UO_258 (O_258,N_9830,N_9699);
and UO_259 (O_259,N_9701,N_9545);
xor UO_260 (O_260,N_9750,N_9835);
nor UO_261 (O_261,N_9859,N_9987);
and UO_262 (O_262,N_9912,N_9884);
and UO_263 (O_263,N_9986,N_9741);
nand UO_264 (O_264,N_9542,N_9633);
and UO_265 (O_265,N_9870,N_9883);
nand UO_266 (O_266,N_9658,N_9810);
and UO_267 (O_267,N_9595,N_9585);
nor UO_268 (O_268,N_9544,N_9944);
nor UO_269 (O_269,N_9676,N_9596);
nor UO_270 (O_270,N_9926,N_9733);
nor UO_271 (O_271,N_9863,N_9798);
and UO_272 (O_272,N_9973,N_9799);
nor UO_273 (O_273,N_9949,N_9929);
nor UO_274 (O_274,N_9970,N_9841);
nor UO_275 (O_275,N_9579,N_9958);
nor UO_276 (O_276,N_9998,N_9808);
nand UO_277 (O_277,N_9882,N_9841);
nand UO_278 (O_278,N_9980,N_9997);
and UO_279 (O_279,N_9752,N_9823);
nor UO_280 (O_280,N_9947,N_9807);
or UO_281 (O_281,N_9625,N_9775);
nand UO_282 (O_282,N_9983,N_9738);
or UO_283 (O_283,N_9888,N_9529);
nor UO_284 (O_284,N_9820,N_9646);
and UO_285 (O_285,N_9763,N_9722);
nor UO_286 (O_286,N_9528,N_9967);
or UO_287 (O_287,N_9753,N_9598);
nor UO_288 (O_288,N_9627,N_9745);
nand UO_289 (O_289,N_9609,N_9700);
nor UO_290 (O_290,N_9685,N_9884);
nor UO_291 (O_291,N_9928,N_9866);
and UO_292 (O_292,N_9810,N_9924);
nand UO_293 (O_293,N_9536,N_9624);
nand UO_294 (O_294,N_9800,N_9656);
or UO_295 (O_295,N_9799,N_9608);
nor UO_296 (O_296,N_9720,N_9785);
nor UO_297 (O_297,N_9695,N_9743);
nor UO_298 (O_298,N_9605,N_9615);
and UO_299 (O_299,N_9669,N_9983);
nand UO_300 (O_300,N_9894,N_9718);
nor UO_301 (O_301,N_9878,N_9592);
and UO_302 (O_302,N_9611,N_9610);
or UO_303 (O_303,N_9507,N_9592);
and UO_304 (O_304,N_9689,N_9717);
or UO_305 (O_305,N_9651,N_9981);
nor UO_306 (O_306,N_9622,N_9752);
xnor UO_307 (O_307,N_9687,N_9803);
or UO_308 (O_308,N_9918,N_9601);
nand UO_309 (O_309,N_9553,N_9512);
or UO_310 (O_310,N_9560,N_9910);
nor UO_311 (O_311,N_9834,N_9627);
and UO_312 (O_312,N_9604,N_9739);
nor UO_313 (O_313,N_9810,N_9700);
or UO_314 (O_314,N_9794,N_9629);
nand UO_315 (O_315,N_9908,N_9780);
and UO_316 (O_316,N_9575,N_9866);
or UO_317 (O_317,N_9852,N_9801);
nand UO_318 (O_318,N_9825,N_9675);
or UO_319 (O_319,N_9698,N_9726);
and UO_320 (O_320,N_9979,N_9871);
and UO_321 (O_321,N_9831,N_9961);
nand UO_322 (O_322,N_9871,N_9592);
nor UO_323 (O_323,N_9611,N_9566);
nand UO_324 (O_324,N_9591,N_9783);
or UO_325 (O_325,N_9730,N_9630);
nand UO_326 (O_326,N_9848,N_9816);
xor UO_327 (O_327,N_9977,N_9711);
or UO_328 (O_328,N_9808,N_9755);
or UO_329 (O_329,N_9808,N_9942);
nor UO_330 (O_330,N_9568,N_9714);
nand UO_331 (O_331,N_9660,N_9810);
and UO_332 (O_332,N_9863,N_9501);
and UO_333 (O_333,N_9926,N_9961);
nand UO_334 (O_334,N_9992,N_9668);
or UO_335 (O_335,N_9882,N_9711);
xor UO_336 (O_336,N_9918,N_9821);
and UO_337 (O_337,N_9960,N_9628);
nor UO_338 (O_338,N_9899,N_9768);
nor UO_339 (O_339,N_9934,N_9922);
or UO_340 (O_340,N_9616,N_9643);
nand UO_341 (O_341,N_9510,N_9710);
and UO_342 (O_342,N_9599,N_9658);
and UO_343 (O_343,N_9854,N_9855);
nor UO_344 (O_344,N_9914,N_9530);
nand UO_345 (O_345,N_9573,N_9699);
nand UO_346 (O_346,N_9556,N_9612);
and UO_347 (O_347,N_9518,N_9778);
nand UO_348 (O_348,N_9993,N_9652);
nor UO_349 (O_349,N_9660,N_9822);
or UO_350 (O_350,N_9972,N_9698);
or UO_351 (O_351,N_9594,N_9977);
nor UO_352 (O_352,N_9627,N_9628);
or UO_353 (O_353,N_9653,N_9724);
nor UO_354 (O_354,N_9781,N_9725);
or UO_355 (O_355,N_9696,N_9970);
nor UO_356 (O_356,N_9683,N_9932);
xnor UO_357 (O_357,N_9741,N_9666);
or UO_358 (O_358,N_9564,N_9638);
and UO_359 (O_359,N_9766,N_9692);
or UO_360 (O_360,N_9921,N_9725);
or UO_361 (O_361,N_9899,N_9711);
nor UO_362 (O_362,N_9651,N_9586);
or UO_363 (O_363,N_9715,N_9635);
nand UO_364 (O_364,N_9527,N_9695);
nand UO_365 (O_365,N_9681,N_9513);
or UO_366 (O_366,N_9721,N_9787);
nor UO_367 (O_367,N_9724,N_9841);
nor UO_368 (O_368,N_9976,N_9698);
or UO_369 (O_369,N_9933,N_9895);
nand UO_370 (O_370,N_9960,N_9896);
and UO_371 (O_371,N_9733,N_9552);
nand UO_372 (O_372,N_9983,N_9591);
and UO_373 (O_373,N_9714,N_9987);
nand UO_374 (O_374,N_9735,N_9981);
xnor UO_375 (O_375,N_9551,N_9729);
nor UO_376 (O_376,N_9872,N_9822);
nand UO_377 (O_377,N_9923,N_9859);
nor UO_378 (O_378,N_9681,N_9746);
and UO_379 (O_379,N_9504,N_9703);
nor UO_380 (O_380,N_9979,N_9726);
or UO_381 (O_381,N_9606,N_9749);
and UO_382 (O_382,N_9699,N_9589);
or UO_383 (O_383,N_9755,N_9911);
nand UO_384 (O_384,N_9617,N_9904);
xnor UO_385 (O_385,N_9580,N_9820);
and UO_386 (O_386,N_9564,N_9734);
and UO_387 (O_387,N_9971,N_9920);
or UO_388 (O_388,N_9602,N_9653);
nand UO_389 (O_389,N_9754,N_9635);
nor UO_390 (O_390,N_9809,N_9710);
nand UO_391 (O_391,N_9698,N_9603);
and UO_392 (O_392,N_9996,N_9877);
nor UO_393 (O_393,N_9942,N_9827);
nor UO_394 (O_394,N_9579,N_9680);
nor UO_395 (O_395,N_9867,N_9556);
or UO_396 (O_396,N_9787,N_9805);
nor UO_397 (O_397,N_9593,N_9631);
nor UO_398 (O_398,N_9623,N_9629);
and UO_399 (O_399,N_9869,N_9800);
and UO_400 (O_400,N_9913,N_9644);
xnor UO_401 (O_401,N_9798,N_9855);
nand UO_402 (O_402,N_9822,N_9755);
nand UO_403 (O_403,N_9679,N_9564);
or UO_404 (O_404,N_9792,N_9608);
nor UO_405 (O_405,N_9612,N_9789);
or UO_406 (O_406,N_9521,N_9979);
nand UO_407 (O_407,N_9890,N_9806);
and UO_408 (O_408,N_9790,N_9743);
and UO_409 (O_409,N_9749,N_9661);
and UO_410 (O_410,N_9747,N_9879);
nor UO_411 (O_411,N_9701,N_9825);
nor UO_412 (O_412,N_9751,N_9642);
or UO_413 (O_413,N_9509,N_9871);
and UO_414 (O_414,N_9826,N_9698);
or UO_415 (O_415,N_9604,N_9524);
nand UO_416 (O_416,N_9627,N_9942);
nand UO_417 (O_417,N_9812,N_9884);
or UO_418 (O_418,N_9883,N_9839);
and UO_419 (O_419,N_9537,N_9740);
or UO_420 (O_420,N_9735,N_9958);
and UO_421 (O_421,N_9694,N_9926);
nor UO_422 (O_422,N_9571,N_9583);
nand UO_423 (O_423,N_9991,N_9780);
and UO_424 (O_424,N_9561,N_9838);
nor UO_425 (O_425,N_9511,N_9776);
nor UO_426 (O_426,N_9949,N_9584);
nor UO_427 (O_427,N_9915,N_9656);
nand UO_428 (O_428,N_9760,N_9829);
or UO_429 (O_429,N_9507,N_9570);
or UO_430 (O_430,N_9917,N_9701);
nand UO_431 (O_431,N_9592,N_9894);
and UO_432 (O_432,N_9556,N_9889);
nand UO_433 (O_433,N_9877,N_9691);
nand UO_434 (O_434,N_9639,N_9676);
nand UO_435 (O_435,N_9655,N_9944);
nor UO_436 (O_436,N_9996,N_9742);
and UO_437 (O_437,N_9945,N_9799);
or UO_438 (O_438,N_9506,N_9915);
nand UO_439 (O_439,N_9639,N_9829);
nand UO_440 (O_440,N_9634,N_9903);
xor UO_441 (O_441,N_9751,N_9662);
or UO_442 (O_442,N_9767,N_9871);
nor UO_443 (O_443,N_9840,N_9958);
and UO_444 (O_444,N_9869,N_9746);
or UO_445 (O_445,N_9512,N_9604);
or UO_446 (O_446,N_9990,N_9585);
and UO_447 (O_447,N_9632,N_9838);
nor UO_448 (O_448,N_9698,N_9554);
and UO_449 (O_449,N_9577,N_9717);
nand UO_450 (O_450,N_9786,N_9849);
or UO_451 (O_451,N_9522,N_9927);
nand UO_452 (O_452,N_9693,N_9937);
nor UO_453 (O_453,N_9679,N_9712);
and UO_454 (O_454,N_9779,N_9518);
and UO_455 (O_455,N_9567,N_9746);
nand UO_456 (O_456,N_9931,N_9866);
nand UO_457 (O_457,N_9933,N_9899);
nand UO_458 (O_458,N_9809,N_9921);
nor UO_459 (O_459,N_9668,N_9946);
nand UO_460 (O_460,N_9766,N_9636);
and UO_461 (O_461,N_9546,N_9561);
or UO_462 (O_462,N_9579,N_9904);
or UO_463 (O_463,N_9732,N_9523);
nor UO_464 (O_464,N_9946,N_9991);
or UO_465 (O_465,N_9926,N_9984);
or UO_466 (O_466,N_9905,N_9623);
nand UO_467 (O_467,N_9948,N_9690);
and UO_468 (O_468,N_9945,N_9652);
and UO_469 (O_469,N_9681,N_9608);
nor UO_470 (O_470,N_9809,N_9669);
nand UO_471 (O_471,N_9563,N_9970);
nor UO_472 (O_472,N_9621,N_9910);
nor UO_473 (O_473,N_9579,N_9846);
nand UO_474 (O_474,N_9562,N_9949);
and UO_475 (O_475,N_9714,N_9950);
nand UO_476 (O_476,N_9828,N_9813);
nor UO_477 (O_477,N_9505,N_9726);
nor UO_478 (O_478,N_9775,N_9568);
or UO_479 (O_479,N_9952,N_9713);
and UO_480 (O_480,N_9616,N_9538);
nor UO_481 (O_481,N_9812,N_9643);
or UO_482 (O_482,N_9860,N_9896);
nand UO_483 (O_483,N_9675,N_9786);
nand UO_484 (O_484,N_9771,N_9673);
nor UO_485 (O_485,N_9776,N_9644);
and UO_486 (O_486,N_9893,N_9721);
nor UO_487 (O_487,N_9965,N_9761);
nand UO_488 (O_488,N_9710,N_9835);
nand UO_489 (O_489,N_9941,N_9855);
xnor UO_490 (O_490,N_9905,N_9714);
nor UO_491 (O_491,N_9545,N_9551);
nand UO_492 (O_492,N_9895,N_9985);
nand UO_493 (O_493,N_9784,N_9546);
and UO_494 (O_494,N_9620,N_9982);
nand UO_495 (O_495,N_9752,N_9896);
and UO_496 (O_496,N_9869,N_9708);
nor UO_497 (O_497,N_9526,N_9660);
or UO_498 (O_498,N_9758,N_9986);
xnor UO_499 (O_499,N_9560,N_9914);
xor UO_500 (O_500,N_9617,N_9963);
nor UO_501 (O_501,N_9907,N_9573);
and UO_502 (O_502,N_9850,N_9784);
nand UO_503 (O_503,N_9553,N_9578);
and UO_504 (O_504,N_9724,N_9795);
and UO_505 (O_505,N_9724,N_9820);
nor UO_506 (O_506,N_9524,N_9644);
nor UO_507 (O_507,N_9873,N_9915);
nor UO_508 (O_508,N_9859,N_9574);
or UO_509 (O_509,N_9878,N_9631);
and UO_510 (O_510,N_9737,N_9678);
and UO_511 (O_511,N_9573,N_9864);
or UO_512 (O_512,N_9653,N_9597);
nand UO_513 (O_513,N_9894,N_9822);
and UO_514 (O_514,N_9958,N_9544);
and UO_515 (O_515,N_9694,N_9729);
or UO_516 (O_516,N_9806,N_9683);
nand UO_517 (O_517,N_9755,N_9662);
nand UO_518 (O_518,N_9678,N_9910);
or UO_519 (O_519,N_9758,N_9818);
nor UO_520 (O_520,N_9789,N_9948);
and UO_521 (O_521,N_9747,N_9744);
nor UO_522 (O_522,N_9599,N_9770);
nand UO_523 (O_523,N_9832,N_9937);
nand UO_524 (O_524,N_9835,N_9839);
nor UO_525 (O_525,N_9577,N_9894);
nand UO_526 (O_526,N_9739,N_9640);
or UO_527 (O_527,N_9755,N_9799);
and UO_528 (O_528,N_9981,N_9989);
and UO_529 (O_529,N_9922,N_9793);
xor UO_530 (O_530,N_9883,N_9802);
or UO_531 (O_531,N_9746,N_9954);
nor UO_532 (O_532,N_9745,N_9533);
and UO_533 (O_533,N_9567,N_9987);
and UO_534 (O_534,N_9886,N_9641);
nor UO_535 (O_535,N_9885,N_9529);
or UO_536 (O_536,N_9527,N_9504);
nor UO_537 (O_537,N_9624,N_9717);
nand UO_538 (O_538,N_9926,N_9870);
or UO_539 (O_539,N_9747,N_9996);
nor UO_540 (O_540,N_9722,N_9651);
or UO_541 (O_541,N_9848,N_9822);
or UO_542 (O_542,N_9971,N_9503);
and UO_543 (O_543,N_9512,N_9710);
and UO_544 (O_544,N_9941,N_9799);
nor UO_545 (O_545,N_9857,N_9948);
and UO_546 (O_546,N_9736,N_9631);
nor UO_547 (O_547,N_9740,N_9564);
xnor UO_548 (O_548,N_9611,N_9848);
nand UO_549 (O_549,N_9559,N_9813);
and UO_550 (O_550,N_9532,N_9876);
and UO_551 (O_551,N_9515,N_9570);
and UO_552 (O_552,N_9582,N_9610);
or UO_553 (O_553,N_9799,N_9834);
nand UO_554 (O_554,N_9921,N_9635);
nor UO_555 (O_555,N_9806,N_9920);
or UO_556 (O_556,N_9565,N_9788);
or UO_557 (O_557,N_9784,N_9543);
nand UO_558 (O_558,N_9843,N_9938);
or UO_559 (O_559,N_9671,N_9541);
or UO_560 (O_560,N_9596,N_9649);
or UO_561 (O_561,N_9544,N_9895);
nand UO_562 (O_562,N_9634,N_9901);
nand UO_563 (O_563,N_9797,N_9523);
or UO_564 (O_564,N_9587,N_9962);
nand UO_565 (O_565,N_9779,N_9781);
nor UO_566 (O_566,N_9531,N_9783);
xnor UO_567 (O_567,N_9904,N_9728);
or UO_568 (O_568,N_9690,N_9812);
or UO_569 (O_569,N_9651,N_9950);
xnor UO_570 (O_570,N_9722,N_9937);
and UO_571 (O_571,N_9643,N_9762);
nand UO_572 (O_572,N_9911,N_9980);
or UO_573 (O_573,N_9870,N_9858);
nor UO_574 (O_574,N_9873,N_9725);
or UO_575 (O_575,N_9970,N_9805);
nand UO_576 (O_576,N_9716,N_9988);
nand UO_577 (O_577,N_9982,N_9795);
nor UO_578 (O_578,N_9952,N_9511);
nor UO_579 (O_579,N_9978,N_9513);
nand UO_580 (O_580,N_9750,N_9996);
and UO_581 (O_581,N_9562,N_9779);
or UO_582 (O_582,N_9754,N_9723);
or UO_583 (O_583,N_9777,N_9831);
nor UO_584 (O_584,N_9518,N_9537);
and UO_585 (O_585,N_9945,N_9550);
and UO_586 (O_586,N_9761,N_9786);
and UO_587 (O_587,N_9589,N_9639);
and UO_588 (O_588,N_9834,N_9986);
and UO_589 (O_589,N_9895,N_9700);
or UO_590 (O_590,N_9918,N_9572);
and UO_591 (O_591,N_9970,N_9940);
and UO_592 (O_592,N_9753,N_9580);
nand UO_593 (O_593,N_9555,N_9625);
or UO_594 (O_594,N_9654,N_9598);
and UO_595 (O_595,N_9760,N_9808);
nand UO_596 (O_596,N_9632,N_9502);
nor UO_597 (O_597,N_9531,N_9631);
nand UO_598 (O_598,N_9945,N_9693);
or UO_599 (O_599,N_9729,N_9589);
nor UO_600 (O_600,N_9698,N_9757);
and UO_601 (O_601,N_9846,N_9550);
or UO_602 (O_602,N_9821,N_9662);
and UO_603 (O_603,N_9852,N_9502);
and UO_604 (O_604,N_9515,N_9629);
or UO_605 (O_605,N_9946,N_9961);
or UO_606 (O_606,N_9815,N_9732);
and UO_607 (O_607,N_9718,N_9645);
nand UO_608 (O_608,N_9538,N_9796);
nor UO_609 (O_609,N_9999,N_9831);
and UO_610 (O_610,N_9953,N_9990);
or UO_611 (O_611,N_9696,N_9693);
nand UO_612 (O_612,N_9597,N_9872);
xor UO_613 (O_613,N_9626,N_9960);
or UO_614 (O_614,N_9529,N_9814);
nand UO_615 (O_615,N_9979,N_9595);
nand UO_616 (O_616,N_9817,N_9920);
nand UO_617 (O_617,N_9926,N_9900);
nor UO_618 (O_618,N_9863,N_9552);
or UO_619 (O_619,N_9605,N_9748);
and UO_620 (O_620,N_9631,N_9952);
and UO_621 (O_621,N_9885,N_9903);
and UO_622 (O_622,N_9921,N_9952);
nand UO_623 (O_623,N_9639,N_9872);
and UO_624 (O_624,N_9942,N_9568);
or UO_625 (O_625,N_9989,N_9842);
nand UO_626 (O_626,N_9792,N_9878);
and UO_627 (O_627,N_9798,N_9908);
nand UO_628 (O_628,N_9861,N_9975);
and UO_629 (O_629,N_9836,N_9752);
and UO_630 (O_630,N_9591,N_9875);
and UO_631 (O_631,N_9940,N_9868);
nand UO_632 (O_632,N_9509,N_9748);
or UO_633 (O_633,N_9754,N_9876);
nand UO_634 (O_634,N_9586,N_9980);
nand UO_635 (O_635,N_9641,N_9968);
or UO_636 (O_636,N_9516,N_9589);
or UO_637 (O_637,N_9530,N_9773);
or UO_638 (O_638,N_9609,N_9775);
nand UO_639 (O_639,N_9736,N_9563);
nand UO_640 (O_640,N_9812,N_9789);
nand UO_641 (O_641,N_9871,N_9990);
nor UO_642 (O_642,N_9842,N_9877);
or UO_643 (O_643,N_9725,N_9628);
or UO_644 (O_644,N_9990,N_9644);
nor UO_645 (O_645,N_9570,N_9581);
nand UO_646 (O_646,N_9610,N_9824);
or UO_647 (O_647,N_9681,N_9869);
and UO_648 (O_648,N_9942,N_9599);
nand UO_649 (O_649,N_9974,N_9939);
nor UO_650 (O_650,N_9972,N_9522);
nor UO_651 (O_651,N_9968,N_9606);
and UO_652 (O_652,N_9904,N_9864);
nor UO_653 (O_653,N_9901,N_9740);
xor UO_654 (O_654,N_9713,N_9602);
nor UO_655 (O_655,N_9657,N_9659);
and UO_656 (O_656,N_9834,N_9981);
or UO_657 (O_657,N_9947,N_9740);
and UO_658 (O_658,N_9597,N_9777);
and UO_659 (O_659,N_9998,N_9909);
nand UO_660 (O_660,N_9703,N_9880);
nor UO_661 (O_661,N_9695,N_9553);
and UO_662 (O_662,N_9512,N_9922);
or UO_663 (O_663,N_9761,N_9523);
or UO_664 (O_664,N_9611,N_9723);
nand UO_665 (O_665,N_9844,N_9788);
or UO_666 (O_666,N_9598,N_9907);
nand UO_667 (O_667,N_9631,N_9618);
and UO_668 (O_668,N_9539,N_9695);
nor UO_669 (O_669,N_9530,N_9963);
or UO_670 (O_670,N_9510,N_9626);
or UO_671 (O_671,N_9685,N_9812);
or UO_672 (O_672,N_9889,N_9512);
and UO_673 (O_673,N_9866,N_9667);
nand UO_674 (O_674,N_9848,N_9576);
or UO_675 (O_675,N_9590,N_9950);
or UO_676 (O_676,N_9736,N_9630);
and UO_677 (O_677,N_9965,N_9868);
xor UO_678 (O_678,N_9727,N_9893);
and UO_679 (O_679,N_9830,N_9844);
xor UO_680 (O_680,N_9774,N_9602);
nor UO_681 (O_681,N_9550,N_9713);
or UO_682 (O_682,N_9709,N_9735);
nor UO_683 (O_683,N_9865,N_9776);
or UO_684 (O_684,N_9936,N_9646);
nand UO_685 (O_685,N_9605,N_9956);
nand UO_686 (O_686,N_9922,N_9854);
and UO_687 (O_687,N_9922,N_9509);
nand UO_688 (O_688,N_9857,N_9893);
nand UO_689 (O_689,N_9680,N_9964);
nand UO_690 (O_690,N_9589,N_9667);
nor UO_691 (O_691,N_9516,N_9501);
nand UO_692 (O_692,N_9864,N_9902);
nor UO_693 (O_693,N_9839,N_9915);
and UO_694 (O_694,N_9640,N_9773);
nor UO_695 (O_695,N_9782,N_9697);
nor UO_696 (O_696,N_9659,N_9530);
nor UO_697 (O_697,N_9965,N_9772);
nand UO_698 (O_698,N_9699,N_9736);
nor UO_699 (O_699,N_9548,N_9511);
and UO_700 (O_700,N_9509,N_9911);
nand UO_701 (O_701,N_9912,N_9504);
or UO_702 (O_702,N_9851,N_9942);
and UO_703 (O_703,N_9876,N_9835);
or UO_704 (O_704,N_9702,N_9912);
or UO_705 (O_705,N_9826,N_9518);
nor UO_706 (O_706,N_9798,N_9620);
and UO_707 (O_707,N_9729,N_9879);
or UO_708 (O_708,N_9988,N_9528);
nand UO_709 (O_709,N_9561,N_9886);
nor UO_710 (O_710,N_9812,N_9848);
nand UO_711 (O_711,N_9640,N_9795);
nor UO_712 (O_712,N_9618,N_9513);
or UO_713 (O_713,N_9500,N_9986);
nand UO_714 (O_714,N_9931,N_9674);
nor UO_715 (O_715,N_9922,N_9852);
nand UO_716 (O_716,N_9576,N_9982);
nand UO_717 (O_717,N_9835,N_9658);
and UO_718 (O_718,N_9865,N_9864);
nand UO_719 (O_719,N_9748,N_9923);
and UO_720 (O_720,N_9953,N_9621);
and UO_721 (O_721,N_9794,N_9882);
or UO_722 (O_722,N_9651,N_9568);
nor UO_723 (O_723,N_9773,N_9981);
or UO_724 (O_724,N_9571,N_9746);
nand UO_725 (O_725,N_9669,N_9686);
nor UO_726 (O_726,N_9742,N_9972);
nor UO_727 (O_727,N_9871,N_9547);
nand UO_728 (O_728,N_9856,N_9554);
nand UO_729 (O_729,N_9898,N_9933);
and UO_730 (O_730,N_9970,N_9875);
nor UO_731 (O_731,N_9814,N_9636);
and UO_732 (O_732,N_9714,N_9619);
and UO_733 (O_733,N_9910,N_9666);
and UO_734 (O_734,N_9851,N_9974);
or UO_735 (O_735,N_9939,N_9716);
and UO_736 (O_736,N_9564,N_9639);
nor UO_737 (O_737,N_9972,N_9663);
and UO_738 (O_738,N_9702,N_9718);
nand UO_739 (O_739,N_9692,N_9906);
or UO_740 (O_740,N_9763,N_9639);
nand UO_741 (O_741,N_9680,N_9608);
or UO_742 (O_742,N_9878,N_9856);
nor UO_743 (O_743,N_9587,N_9611);
or UO_744 (O_744,N_9715,N_9537);
or UO_745 (O_745,N_9586,N_9503);
nand UO_746 (O_746,N_9878,N_9983);
nand UO_747 (O_747,N_9707,N_9592);
or UO_748 (O_748,N_9631,N_9722);
or UO_749 (O_749,N_9740,N_9513);
and UO_750 (O_750,N_9805,N_9890);
and UO_751 (O_751,N_9712,N_9651);
nand UO_752 (O_752,N_9798,N_9515);
and UO_753 (O_753,N_9810,N_9829);
nor UO_754 (O_754,N_9550,N_9943);
and UO_755 (O_755,N_9664,N_9641);
nor UO_756 (O_756,N_9669,N_9527);
nand UO_757 (O_757,N_9886,N_9591);
or UO_758 (O_758,N_9649,N_9997);
and UO_759 (O_759,N_9724,N_9689);
nand UO_760 (O_760,N_9650,N_9753);
nand UO_761 (O_761,N_9750,N_9855);
or UO_762 (O_762,N_9973,N_9690);
nand UO_763 (O_763,N_9605,N_9842);
xnor UO_764 (O_764,N_9709,N_9582);
nor UO_765 (O_765,N_9621,N_9889);
nor UO_766 (O_766,N_9859,N_9932);
nand UO_767 (O_767,N_9840,N_9762);
nor UO_768 (O_768,N_9875,N_9984);
or UO_769 (O_769,N_9715,N_9782);
nand UO_770 (O_770,N_9670,N_9842);
nand UO_771 (O_771,N_9746,N_9517);
nand UO_772 (O_772,N_9756,N_9619);
or UO_773 (O_773,N_9557,N_9764);
nor UO_774 (O_774,N_9662,N_9705);
or UO_775 (O_775,N_9684,N_9627);
nand UO_776 (O_776,N_9974,N_9897);
nor UO_777 (O_777,N_9504,N_9755);
and UO_778 (O_778,N_9811,N_9517);
nor UO_779 (O_779,N_9958,N_9617);
and UO_780 (O_780,N_9585,N_9614);
and UO_781 (O_781,N_9933,N_9968);
or UO_782 (O_782,N_9701,N_9966);
and UO_783 (O_783,N_9763,N_9929);
and UO_784 (O_784,N_9594,N_9985);
nand UO_785 (O_785,N_9996,N_9905);
or UO_786 (O_786,N_9808,N_9996);
and UO_787 (O_787,N_9595,N_9514);
nand UO_788 (O_788,N_9785,N_9839);
nor UO_789 (O_789,N_9867,N_9875);
or UO_790 (O_790,N_9899,N_9563);
nor UO_791 (O_791,N_9568,N_9987);
and UO_792 (O_792,N_9610,N_9781);
nor UO_793 (O_793,N_9503,N_9630);
nand UO_794 (O_794,N_9848,N_9976);
or UO_795 (O_795,N_9704,N_9666);
or UO_796 (O_796,N_9659,N_9508);
nor UO_797 (O_797,N_9543,N_9793);
and UO_798 (O_798,N_9979,N_9836);
and UO_799 (O_799,N_9631,N_9971);
or UO_800 (O_800,N_9735,N_9918);
and UO_801 (O_801,N_9616,N_9695);
and UO_802 (O_802,N_9834,N_9704);
xor UO_803 (O_803,N_9800,N_9895);
and UO_804 (O_804,N_9698,N_9506);
or UO_805 (O_805,N_9958,N_9720);
nor UO_806 (O_806,N_9954,N_9508);
or UO_807 (O_807,N_9754,N_9840);
xnor UO_808 (O_808,N_9653,N_9932);
nand UO_809 (O_809,N_9946,N_9819);
and UO_810 (O_810,N_9764,N_9606);
nand UO_811 (O_811,N_9730,N_9503);
nor UO_812 (O_812,N_9565,N_9636);
xnor UO_813 (O_813,N_9842,N_9744);
or UO_814 (O_814,N_9604,N_9682);
and UO_815 (O_815,N_9668,N_9971);
and UO_816 (O_816,N_9999,N_9779);
and UO_817 (O_817,N_9718,N_9971);
nor UO_818 (O_818,N_9744,N_9674);
nand UO_819 (O_819,N_9679,N_9693);
or UO_820 (O_820,N_9942,N_9921);
nor UO_821 (O_821,N_9540,N_9797);
nor UO_822 (O_822,N_9575,N_9680);
and UO_823 (O_823,N_9590,N_9549);
nor UO_824 (O_824,N_9751,N_9648);
and UO_825 (O_825,N_9749,N_9605);
or UO_826 (O_826,N_9605,N_9970);
or UO_827 (O_827,N_9581,N_9636);
or UO_828 (O_828,N_9555,N_9745);
and UO_829 (O_829,N_9968,N_9994);
nor UO_830 (O_830,N_9922,N_9810);
and UO_831 (O_831,N_9922,N_9652);
or UO_832 (O_832,N_9600,N_9819);
nand UO_833 (O_833,N_9811,N_9898);
and UO_834 (O_834,N_9802,N_9854);
nor UO_835 (O_835,N_9669,N_9587);
or UO_836 (O_836,N_9661,N_9698);
nand UO_837 (O_837,N_9836,N_9852);
nand UO_838 (O_838,N_9876,N_9949);
and UO_839 (O_839,N_9918,N_9560);
nand UO_840 (O_840,N_9987,N_9634);
nor UO_841 (O_841,N_9601,N_9525);
or UO_842 (O_842,N_9830,N_9559);
or UO_843 (O_843,N_9976,N_9562);
and UO_844 (O_844,N_9639,N_9953);
and UO_845 (O_845,N_9911,N_9580);
or UO_846 (O_846,N_9884,N_9509);
xor UO_847 (O_847,N_9840,N_9520);
nand UO_848 (O_848,N_9918,N_9559);
nand UO_849 (O_849,N_9714,N_9931);
or UO_850 (O_850,N_9669,N_9670);
or UO_851 (O_851,N_9724,N_9731);
and UO_852 (O_852,N_9990,N_9799);
and UO_853 (O_853,N_9563,N_9870);
and UO_854 (O_854,N_9876,N_9983);
nand UO_855 (O_855,N_9640,N_9573);
nor UO_856 (O_856,N_9531,N_9790);
and UO_857 (O_857,N_9727,N_9848);
and UO_858 (O_858,N_9711,N_9598);
nor UO_859 (O_859,N_9503,N_9874);
and UO_860 (O_860,N_9979,N_9735);
nor UO_861 (O_861,N_9717,N_9569);
and UO_862 (O_862,N_9541,N_9515);
nor UO_863 (O_863,N_9695,N_9525);
and UO_864 (O_864,N_9518,N_9991);
nand UO_865 (O_865,N_9672,N_9850);
or UO_866 (O_866,N_9633,N_9675);
and UO_867 (O_867,N_9834,N_9832);
and UO_868 (O_868,N_9795,N_9888);
and UO_869 (O_869,N_9806,N_9865);
nor UO_870 (O_870,N_9832,N_9654);
nand UO_871 (O_871,N_9970,N_9557);
nand UO_872 (O_872,N_9785,N_9915);
and UO_873 (O_873,N_9775,N_9683);
nor UO_874 (O_874,N_9832,N_9895);
nor UO_875 (O_875,N_9780,N_9636);
and UO_876 (O_876,N_9621,N_9740);
and UO_877 (O_877,N_9800,N_9788);
nand UO_878 (O_878,N_9627,N_9522);
nand UO_879 (O_879,N_9603,N_9837);
nand UO_880 (O_880,N_9770,N_9587);
or UO_881 (O_881,N_9978,N_9897);
or UO_882 (O_882,N_9756,N_9772);
and UO_883 (O_883,N_9990,N_9579);
and UO_884 (O_884,N_9712,N_9934);
or UO_885 (O_885,N_9923,N_9587);
nor UO_886 (O_886,N_9609,N_9746);
or UO_887 (O_887,N_9938,N_9891);
or UO_888 (O_888,N_9859,N_9846);
nand UO_889 (O_889,N_9757,N_9553);
or UO_890 (O_890,N_9902,N_9850);
nor UO_891 (O_891,N_9523,N_9728);
nor UO_892 (O_892,N_9995,N_9780);
and UO_893 (O_893,N_9592,N_9562);
nand UO_894 (O_894,N_9631,N_9759);
or UO_895 (O_895,N_9734,N_9890);
or UO_896 (O_896,N_9813,N_9628);
nor UO_897 (O_897,N_9947,N_9853);
and UO_898 (O_898,N_9696,N_9727);
and UO_899 (O_899,N_9956,N_9588);
nor UO_900 (O_900,N_9719,N_9916);
and UO_901 (O_901,N_9537,N_9751);
and UO_902 (O_902,N_9867,N_9883);
or UO_903 (O_903,N_9590,N_9548);
nand UO_904 (O_904,N_9982,N_9770);
nand UO_905 (O_905,N_9505,N_9732);
and UO_906 (O_906,N_9897,N_9504);
nand UO_907 (O_907,N_9601,N_9769);
nand UO_908 (O_908,N_9575,N_9819);
nand UO_909 (O_909,N_9682,N_9985);
and UO_910 (O_910,N_9593,N_9622);
nor UO_911 (O_911,N_9708,N_9588);
or UO_912 (O_912,N_9770,N_9944);
nand UO_913 (O_913,N_9840,N_9765);
nand UO_914 (O_914,N_9820,N_9919);
nand UO_915 (O_915,N_9645,N_9668);
or UO_916 (O_916,N_9742,N_9590);
and UO_917 (O_917,N_9728,N_9531);
and UO_918 (O_918,N_9660,N_9744);
nand UO_919 (O_919,N_9953,N_9725);
or UO_920 (O_920,N_9649,N_9685);
nor UO_921 (O_921,N_9875,N_9667);
xnor UO_922 (O_922,N_9777,N_9712);
or UO_923 (O_923,N_9911,N_9920);
nand UO_924 (O_924,N_9640,N_9982);
and UO_925 (O_925,N_9934,N_9588);
or UO_926 (O_926,N_9945,N_9931);
and UO_927 (O_927,N_9545,N_9926);
nand UO_928 (O_928,N_9605,N_9701);
and UO_929 (O_929,N_9743,N_9889);
or UO_930 (O_930,N_9516,N_9753);
or UO_931 (O_931,N_9776,N_9643);
or UO_932 (O_932,N_9621,N_9731);
nor UO_933 (O_933,N_9755,N_9971);
and UO_934 (O_934,N_9990,N_9971);
nand UO_935 (O_935,N_9652,N_9995);
and UO_936 (O_936,N_9576,N_9816);
nand UO_937 (O_937,N_9690,N_9714);
or UO_938 (O_938,N_9924,N_9657);
or UO_939 (O_939,N_9712,N_9597);
nor UO_940 (O_940,N_9694,N_9936);
and UO_941 (O_941,N_9562,N_9571);
xor UO_942 (O_942,N_9685,N_9853);
xnor UO_943 (O_943,N_9731,N_9835);
and UO_944 (O_944,N_9690,N_9736);
nand UO_945 (O_945,N_9904,N_9556);
and UO_946 (O_946,N_9821,N_9807);
or UO_947 (O_947,N_9959,N_9634);
nand UO_948 (O_948,N_9679,N_9831);
and UO_949 (O_949,N_9724,N_9664);
or UO_950 (O_950,N_9642,N_9775);
nor UO_951 (O_951,N_9853,N_9911);
nor UO_952 (O_952,N_9935,N_9738);
nor UO_953 (O_953,N_9552,N_9860);
or UO_954 (O_954,N_9815,N_9591);
nand UO_955 (O_955,N_9926,N_9973);
or UO_956 (O_956,N_9631,N_9814);
nor UO_957 (O_957,N_9939,N_9633);
or UO_958 (O_958,N_9651,N_9968);
and UO_959 (O_959,N_9761,N_9704);
nand UO_960 (O_960,N_9647,N_9582);
nand UO_961 (O_961,N_9826,N_9936);
nor UO_962 (O_962,N_9513,N_9716);
and UO_963 (O_963,N_9663,N_9852);
and UO_964 (O_964,N_9529,N_9865);
xor UO_965 (O_965,N_9790,N_9811);
and UO_966 (O_966,N_9987,N_9635);
and UO_967 (O_967,N_9902,N_9833);
nor UO_968 (O_968,N_9674,N_9765);
or UO_969 (O_969,N_9501,N_9836);
and UO_970 (O_970,N_9622,N_9824);
nand UO_971 (O_971,N_9886,N_9512);
nand UO_972 (O_972,N_9651,N_9537);
nand UO_973 (O_973,N_9979,N_9504);
nand UO_974 (O_974,N_9597,N_9814);
and UO_975 (O_975,N_9965,N_9912);
and UO_976 (O_976,N_9897,N_9878);
nor UO_977 (O_977,N_9679,N_9533);
nand UO_978 (O_978,N_9738,N_9851);
or UO_979 (O_979,N_9988,N_9790);
nand UO_980 (O_980,N_9658,N_9503);
and UO_981 (O_981,N_9821,N_9993);
nand UO_982 (O_982,N_9587,N_9591);
or UO_983 (O_983,N_9664,N_9775);
nor UO_984 (O_984,N_9889,N_9977);
and UO_985 (O_985,N_9839,N_9615);
and UO_986 (O_986,N_9776,N_9546);
nor UO_987 (O_987,N_9793,N_9841);
nor UO_988 (O_988,N_9790,N_9831);
nor UO_989 (O_989,N_9624,N_9674);
or UO_990 (O_990,N_9958,N_9894);
nor UO_991 (O_991,N_9716,N_9859);
nand UO_992 (O_992,N_9940,N_9881);
and UO_993 (O_993,N_9678,N_9906);
nand UO_994 (O_994,N_9545,N_9689);
or UO_995 (O_995,N_9510,N_9723);
nand UO_996 (O_996,N_9679,N_9503);
and UO_997 (O_997,N_9600,N_9763);
or UO_998 (O_998,N_9916,N_9587);
nand UO_999 (O_999,N_9788,N_9750);
nand UO_1000 (O_1000,N_9573,N_9615);
nor UO_1001 (O_1001,N_9974,N_9907);
xor UO_1002 (O_1002,N_9612,N_9961);
nor UO_1003 (O_1003,N_9982,N_9638);
nand UO_1004 (O_1004,N_9813,N_9602);
nand UO_1005 (O_1005,N_9511,N_9539);
xnor UO_1006 (O_1006,N_9757,N_9976);
nand UO_1007 (O_1007,N_9676,N_9945);
and UO_1008 (O_1008,N_9739,N_9812);
nand UO_1009 (O_1009,N_9750,N_9864);
nand UO_1010 (O_1010,N_9756,N_9843);
or UO_1011 (O_1011,N_9599,N_9775);
or UO_1012 (O_1012,N_9938,N_9934);
nor UO_1013 (O_1013,N_9938,N_9900);
or UO_1014 (O_1014,N_9852,N_9925);
nor UO_1015 (O_1015,N_9706,N_9869);
nor UO_1016 (O_1016,N_9679,N_9725);
or UO_1017 (O_1017,N_9678,N_9956);
and UO_1018 (O_1018,N_9847,N_9672);
or UO_1019 (O_1019,N_9699,N_9909);
and UO_1020 (O_1020,N_9861,N_9790);
and UO_1021 (O_1021,N_9766,N_9966);
nor UO_1022 (O_1022,N_9534,N_9683);
nor UO_1023 (O_1023,N_9961,N_9755);
nand UO_1024 (O_1024,N_9654,N_9868);
nand UO_1025 (O_1025,N_9665,N_9902);
nand UO_1026 (O_1026,N_9563,N_9880);
nand UO_1027 (O_1027,N_9597,N_9630);
and UO_1028 (O_1028,N_9676,N_9807);
and UO_1029 (O_1029,N_9528,N_9608);
and UO_1030 (O_1030,N_9508,N_9676);
and UO_1031 (O_1031,N_9729,N_9587);
nand UO_1032 (O_1032,N_9659,N_9837);
xnor UO_1033 (O_1033,N_9831,N_9901);
nand UO_1034 (O_1034,N_9919,N_9961);
and UO_1035 (O_1035,N_9541,N_9853);
nand UO_1036 (O_1036,N_9956,N_9606);
nand UO_1037 (O_1037,N_9998,N_9635);
nand UO_1038 (O_1038,N_9936,N_9769);
xnor UO_1039 (O_1039,N_9590,N_9919);
and UO_1040 (O_1040,N_9541,N_9742);
and UO_1041 (O_1041,N_9734,N_9904);
nor UO_1042 (O_1042,N_9656,N_9605);
and UO_1043 (O_1043,N_9795,N_9516);
and UO_1044 (O_1044,N_9590,N_9502);
nor UO_1045 (O_1045,N_9570,N_9719);
nand UO_1046 (O_1046,N_9637,N_9562);
and UO_1047 (O_1047,N_9910,N_9857);
or UO_1048 (O_1048,N_9651,N_9584);
nand UO_1049 (O_1049,N_9883,N_9798);
and UO_1050 (O_1050,N_9678,N_9895);
and UO_1051 (O_1051,N_9729,N_9680);
and UO_1052 (O_1052,N_9771,N_9677);
nor UO_1053 (O_1053,N_9891,N_9817);
nor UO_1054 (O_1054,N_9507,N_9580);
or UO_1055 (O_1055,N_9852,N_9830);
nor UO_1056 (O_1056,N_9636,N_9964);
and UO_1057 (O_1057,N_9712,N_9721);
nand UO_1058 (O_1058,N_9669,N_9760);
nor UO_1059 (O_1059,N_9926,N_9972);
nand UO_1060 (O_1060,N_9719,N_9738);
and UO_1061 (O_1061,N_9510,N_9990);
and UO_1062 (O_1062,N_9578,N_9785);
and UO_1063 (O_1063,N_9777,N_9819);
nand UO_1064 (O_1064,N_9684,N_9597);
and UO_1065 (O_1065,N_9584,N_9991);
and UO_1066 (O_1066,N_9770,N_9878);
and UO_1067 (O_1067,N_9785,N_9722);
nor UO_1068 (O_1068,N_9621,N_9792);
or UO_1069 (O_1069,N_9717,N_9992);
nand UO_1070 (O_1070,N_9880,N_9716);
or UO_1071 (O_1071,N_9579,N_9770);
nand UO_1072 (O_1072,N_9645,N_9999);
nor UO_1073 (O_1073,N_9903,N_9551);
or UO_1074 (O_1074,N_9852,N_9911);
nor UO_1075 (O_1075,N_9651,N_9582);
nand UO_1076 (O_1076,N_9914,N_9529);
or UO_1077 (O_1077,N_9959,N_9598);
or UO_1078 (O_1078,N_9673,N_9536);
and UO_1079 (O_1079,N_9822,N_9808);
or UO_1080 (O_1080,N_9908,N_9808);
or UO_1081 (O_1081,N_9668,N_9685);
nor UO_1082 (O_1082,N_9632,N_9500);
nor UO_1083 (O_1083,N_9578,N_9556);
nand UO_1084 (O_1084,N_9731,N_9747);
nor UO_1085 (O_1085,N_9912,N_9573);
nand UO_1086 (O_1086,N_9652,N_9649);
and UO_1087 (O_1087,N_9929,N_9739);
nor UO_1088 (O_1088,N_9724,N_9520);
nand UO_1089 (O_1089,N_9963,N_9894);
nand UO_1090 (O_1090,N_9960,N_9529);
and UO_1091 (O_1091,N_9592,N_9945);
nand UO_1092 (O_1092,N_9788,N_9720);
or UO_1093 (O_1093,N_9659,N_9843);
nand UO_1094 (O_1094,N_9917,N_9978);
nand UO_1095 (O_1095,N_9824,N_9961);
and UO_1096 (O_1096,N_9643,N_9626);
and UO_1097 (O_1097,N_9997,N_9711);
nor UO_1098 (O_1098,N_9630,N_9543);
nand UO_1099 (O_1099,N_9999,N_9568);
nor UO_1100 (O_1100,N_9847,N_9912);
or UO_1101 (O_1101,N_9945,N_9892);
nor UO_1102 (O_1102,N_9744,N_9891);
nand UO_1103 (O_1103,N_9881,N_9650);
nand UO_1104 (O_1104,N_9899,N_9570);
or UO_1105 (O_1105,N_9761,N_9987);
nand UO_1106 (O_1106,N_9782,N_9576);
and UO_1107 (O_1107,N_9634,N_9732);
nand UO_1108 (O_1108,N_9531,N_9925);
or UO_1109 (O_1109,N_9786,N_9540);
and UO_1110 (O_1110,N_9779,N_9598);
and UO_1111 (O_1111,N_9934,N_9935);
nor UO_1112 (O_1112,N_9578,N_9809);
xnor UO_1113 (O_1113,N_9778,N_9571);
nand UO_1114 (O_1114,N_9520,N_9940);
xnor UO_1115 (O_1115,N_9915,N_9508);
or UO_1116 (O_1116,N_9907,N_9895);
or UO_1117 (O_1117,N_9946,N_9751);
or UO_1118 (O_1118,N_9756,N_9993);
and UO_1119 (O_1119,N_9630,N_9863);
or UO_1120 (O_1120,N_9688,N_9750);
nor UO_1121 (O_1121,N_9848,N_9700);
nand UO_1122 (O_1122,N_9810,N_9747);
xor UO_1123 (O_1123,N_9600,N_9597);
and UO_1124 (O_1124,N_9529,N_9776);
and UO_1125 (O_1125,N_9846,N_9571);
and UO_1126 (O_1126,N_9903,N_9975);
and UO_1127 (O_1127,N_9740,N_9910);
and UO_1128 (O_1128,N_9540,N_9860);
and UO_1129 (O_1129,N_9823,N_9731);
xor UO_1130 (O_1130,N_9887,N_9534);
or UO_1131 (O_1131,N_9785,N_9829);
and UO_1132 (O_1132,N_9642,N_9783);
nand UO_1133 (O_1133,N_9837,N_9644);
nor UO_1134 (O_1134,N_9755,N_9919);
nand UO_1135 (O_1135,N_9771,N_9850);
nand UO_1136 (O_1136,N_9975,N_9911);
xnor UO_1137 (O_1137,N_9727,N_9743);
and UO_1138 (O_1138,N_9722,N_9961);
nor UO_1139 (O_1139,N_9849,N_9893);
nor UO_1140 (O_1140,N_9744,N_9844);
and UO_1141 (O_1141,N_9777,N_9729);
or UO_1142 (O_1142,N_9661,N_9999);
nor UO_1143 (O_1143,N_9573,N_9657);
and UO_1144 (O_1144,N_9598,N_9918);
and UO_1145 (O_1145,N_9599,N_9530);
nor UO_1146 (O_1146,N_9954,N_9837);
nor UO_1147 (O_1147,N_9538,N_9977);
nand UO_1148 (O_1148,N_9600,N_9810);
nor UO_1149 (O_1149,N_9524,N_9980);
xnor UO_1150 (O_1150,N_9537,N_9585);
and UO_1151 (O_1151,N_9543,N_9992);
nor UO_1152 (O_1152,N_9821,N_9745);
nand UO_1153 (O_1153,N_9919,N_9967);
nand UO_1154 (O_1154,N_9708,N_9562);
and UO_1155 (O_1155,N_9520,N_9845);
nor UO_1156 (O_1156,N_9798,N_9822);
nand UO_1157 (O_1157,N_9736,N_9924);
nand UO_1158 (O_1158,N_9830,N_9687);
or UO_1159 (O_1159,N_9724,N_9991);
or UO_1160 (O_1160,N_9813,N_9657);
nand UO_1161 (O_1161,N_9529,N_9528);
nor UO_1162 (O_1162,N_9892,N_9582);
or UO_1163 (O_1163,N_9721,N_9886);
nor UO_1164 (O_1164,N_9906,N_9879);
nand UO_1165 (O_1165,N_9671,N_9560);
nand UO_1166 (O_1166,N_9538,N_9724);
and UO_1167 (O_1167,N_9721,N_9911);
nand UO_1168 (O_1168,N_9665,N_9821);
nor UO_1169 (O_1169,N_9622,N_9787);
nand UO_1170 (O_1170,N_9791,N_9880);
xor UO_1171 (O_1171,N_9566,N_9965);
or UO_1172 (O_1172,N_9892,N_9980);
and UO_1173 (O_1173,N_9703,N_9538);
and UO_1174 (O_1174,N_9631,N_9543);
or UO_1175 (O_1175,N_9723,N_9717);
nor UO_1176 (O_1176,N_9867,N_9848);
nor UO_1177 (O_1177,N_9966,N_9830);
xor UO_1178 (O_1178,N_9612,N_9957);
and UO_1179 (O_1179,N_9748,N_9755);
nor UO_1180 (O_1180,N_9671,N_9865);
and UO_1181 (O_1181,N_9539,N_9610);
and UO_1182 (O_1182,N_9634,N_9774);
and UO_1183 (O_1183,N_9672,N_9750);
nand UO_1184 (O_1184,N_9977,N_9849);
nand UO_1185 (O_1185,N_9944,N_9991);
and UO_1186 (O_1186,N_9943,N_9618);
nand UO_1187 (O_1187,N_9699,N_9531);
nand UO_1188 (O_1188,N_9568,N_9659);
xor UO_1189 (O_1189,N_9781,N_9696);
xor UO_1190 (O_1190,N_9640,N_9871);
and UO_1191 (O_1191,N_9642,N_9860);
nand UO_1192 (O_1192,N_9795,N_9937);
and UO_1193 (O_1193,N_9638,N_9520);
and UO_1194 (O_1194,N_9715,N_9745);
and UO_1195 (O_1195,N_9669,N_9635);
nand UO_1196 (O_1196,N_9775,N_9751);
nand UO_1197 (O_1197,N_9880,N_9530);
and UO_1198 (O_1198,N_9995,N_9963);
nand UO_1199 (O_1199,N_9732,N_9778);
nor UO_1200 (O_1200,N_9936,N_9701);
and UO_1201 (O_1201,N_9923,N_9976);
or UO_1202 (O_1202,N_9569,N_9530);
nand UO_1203 (O_1203,N_9753,N_9743);
and UO_1204 (O_1204,N_9965,N_9826);
or UO_1205 (O_1205,N_9907,N_9672);
or UO_1206 (O_1206,N_9798,N_9969);
and UO_1207 (O_1207,N_9651,N_9762);
nor UO_1208 (O_1208,N_9955,N_9860);
nor UO_1209 (O_1209,N_9731,N_9532);
and UO_1210 (O_1210,N_9964,N_9827);
or UO_1211 (O_1211,N_9580,N_9974);
nand UO_1212 (O_1212,N_9882,N_9529);
and UO_1213 (O_1213,N_9830,N_9670);
and UO_1214 (O_1214,N_9605,N_9780);
nand UO_1215 (O_1215,N_9656,N_9703);
or UO_1216 (O_1216,N_9849,N_9655);
nor UO_1217 (O_1217,N_9904,N_9830);
and UO_1218 (O_1218,N_9672,N_9503);
and UO_1219 (O_1219,N_9764,N_9727);
or UO_1220 (O_1220,N_9819,N_9996);
or UO_1221 (O_1221,N_9794,N_9836);
and UO_1222 (O_1222,N_9899,N_9910);
and UO_1223 (O_1223,N_9801,N_9522);
nand UO_1224 (O_1224,N_9609,N_9520);
or UO_1225 (O_1225,N_9979,N_9507);
nor UO_1226 (O_1226,N_9612,N_9606);
and UO_1227 (O_1227,N_9509,N_9751);
nor UO_1228 (O_1228,N_9950,N_9695);
nor UO_1229 (O_1229,N_9695,N_9655);
nor UO_1230 (O_1230,N_9738,N_9748);
nor UO_1231 (O_1231,N_9796,N_9515);
or UO_1232 (O_1232,N_9860,N_9942);
and UO_1233 (O_1233,N_9953,N_9923);
nor UO_1234 (O_1234,N_9526,N_9623);
nor UO_1235 (O_1235,N_9881,N_9943);
nor UO_1236 (O_1236,N_9833,N_9905);
nor UO_1237 (O_1237,N_9938,N_9895);
nor UO_1238 (O_1238,N_9560,N_9744);
nor UO_1239 (O_1239,N_9609,N_9954);
nor UO_1240 (O_1240,N_9829,N_9981);
or UO_1241 (O_1241,N_9507,N_9910);
nor UO_1242 (O_1242,N_9765,N_9945);
and UO_1243 (O_1243,N_9587,N_9815);
nand UO_1244 (O_1244,N_9968,N_9661);
nor UO_1245 (O_1245,N_9772,N_9589);
nand UO_1246 (O_1246,N_9832,N_9916);
nor UO_1247 (O_1247,N_9620,N_9510);
or UO_1248 (O_1248,N_9777,N_9988);
or UO_1249 (O_1249,N_9900,N_9542);
nor UO_1250 (O_1250,N_9609,N_9834);
nand UO_1251 (O_1251,N_9902,N_9648);
or UO_1252 (O_1252,N_9879,N_9875);
nand UO_1253 (O_1253,N_9985,N_9891);
or UO_1254 (O_1254,N_9747,N_9939);
and UO_1255 (O_1255,N_9849,N_9540);
nand UO_1256 (O_1256,N_9868,N_9835);
and UO_1257 (O_1257,N_9636,N_9663);
or UO_1258 (O_1258,N_9856,N_9540);
and UO_1259 (O_1259,N_9762,N_9746);
xor UO_1260 (O_1260,N_9986,N_9728);
nand UO_1261 (O_1261,N_9825,N_9972);
nor UO_1262 (O_1262,N_9762,N_9816);
and UO_1263 (O_1263,N_9531,N_9638);
nand UO_1264 (O_1264,N_9903,N_9864);
nand UO_1265 (O_1265,N_9610,N_9607);
nand UO_1266 (O_1266,N_9512,N_9841);
nor UO_1267 (O_1267,N_9896,N_9907);
or UO_1268 (O_1268,N_9715,N_9911);
or UO_1269 (O_1269,N_9874,N_9991);
or UO_1270 (O_1270,N_9754,N_9888);
or UO_1271 (O_1271,N_9515,N_9600);
nand UO_1272 (O_1272,N_9551,N_9628);
and UO_1273 (O_1273,N_9663,N_9895);
and UO_1274 (O_1274,N_9757,N_9642);
and UO_1275 (O_1275,N_9977,N_9547);
or UO_1276 (O_1276,N_9946,N_9759);
xor UO_1277 (O_1277,N_9795,N_9846);
or UO_1278 (O_1278,N_9926,N_9947);
nand UO_1279 (O_1279,N_9710,N_9789);
nor UO_1280 (O_1280,N_9550,N_9797);
or UO_1281 (O_1281,N_9868,N_9784);
nand UO_1282 (O_1282,N_9549,N_9727);
nor UO_1283 (O_1283,N_9532,N_9637);
and UO_1284 (O_1284,N_9999,N_9639);
nand UO_1285 (O_1285,N_9788,N_9998);
nand UO_1286 (O_1286,N_9532,N_9506);
nor UO_1287 (O_1287,N_9911,N_9780);
and UO_1288 (O_1288,N_9564,N_9938);
nor UO_1289 (O_1289,N_9806,N_9500);
xnor UO_1290 (O_1290,N_9853,N_9992);
nor UO_1291 (O_1291,N_9976,N_9658);
or UO_1292 (O_1292,N_9586,N_9716);
or UO_1293 (O_1293,N_9962,N_9902);
and UO_1294 (O_1294,N_9970,N_9715);
or UO_1295 (O_1295,N_9550,N_9666);
nor UO_1296 (O_1296,N_9695,N_9548);
and UO_1297 (O_1297,N_9994,N_9830);
nand UO_1298 (O_1298,N_9850,N_9949);
or UO_1299 (O_1299,N_9691,N_9602);
nand UO_1300 (O_1300,N_9825,N_9990);
and UO_1301 (O_1301,N_9654,N_9565);
nor UO_1302 (O_1302,N_9884,N_9789);
nand UO_1303 (O_1303,N_9857,N_9976);
and UO_1304 (O_1304,N_9905,N_9765);
or UO_1305 (O_1305,N_9520,N_9521);
nor UO_1306 (O_1306,N_9914,N_9585);
or UO_1307 (O_1307,N_9842,N_9940);
nand UO_1308 (O_1308,N_9843,N_9675);
nand UO_1309 (O_1309,N_9908,N_9757);
or UO_1310 (O_1310,N_9783,N_9973);
and UO_1311 (O_1311,N_9558,N_9971);
nor UO_1312 (O_1312,N_9929,N_9913);
or UO_1313 (O_1313,N_9708,N_9956);
nand UO_1314 (O_1314,N_9552,N_9884);
and UO_1315 (O_1315,N_9751,N_9788);
nor UO_1316 (O_1316,N_9678,N_9557);
nor UO_1317 (O_1317,N_9675,N_9946);
nand UO_1318 (O_1318,N_9943,N_9687);
xor UO_1319 (O_1319,N_9922,N_9579);
or UO_1320 (O_1320,N_9701,N_9881);
and UO_1321 (O_1321,N_9595,N_9552);
nand UO_1322 (O_1322,N_9538,N_9725);
nand UO_1323 (O_1323,N_9731,N_9687);
or UO_1324 (O_1324,N_9854,N_9881);
or UO_1325 (O_1325,N_9903,N_9956);
and UO_1326 (O_1326,N_9870,N_9992);
or UO_1327 (O_1327,N_9631,N_9664);
nor UO_1328 (O_1328,N_9692,N_9940);
and UO_1329 (O_1329,N_9509,N_9802);
or UO_1330 (O_1330,N_9977,N_9533);
and UO_1331 (O_1331,N_9791,N_9920);
and UO_1332 (O_1332,N_9598,N_9565);
nor UO_1333 (O_1333,N_9701,N_9590);
or UO_1334 (O_1334,N_9568,N_9579);
nand UO_1335 (O_1335,N_9638,N_9523);
or UO_1336 (O_1336,N_9651,N_9531);
and UO_1337 (O_1337,N_9949,N_9852);
nand UO_1338 (O_1338,N_9858,N_9914);
nand UO_1339 (O_1339,N_9536,N_9716);
nor UO_1340 (O_1340,N_9789,N_9656);
or UO_1341 (O_1341,N_9634,N_9807);
nor UO_1342 (O_1342,N_9847,N_9794);
nor UO_1343 (O_1343,N_9555,N_9920);
nand UO_1344 (O_1344,N_9718,N_9913);
nor UO_1345 (O_1345,N_9898,N_9822);
nor UO_1346 (O_1346,N_9582,N_9683);
nor UO_1347 (O_1347,N_9503,N_9582);
nand UO_1348 (O_1348,N_9926,N_9760);
or UO_1349 (O_1349,N_9675,N_9724);
and UO_1350 (O_1350,N_9648,N_9690);
or UO_1351 (O_1351,N_9805,N_9723);
and UO_1352 (O_1352,N_9712,N_9655);
or UO_1353 (O_1353,N_9695,N_9981);
nor UO_1354 (O_1354,N_9773,N_9679);
and UO_1355 (O_1355,N_9650,N_9910);
or UO_1356 (O_1356,N_9870,N_9843);
nand UO_1357 (O_1357,N_9612,N_9962);
or UO_1358 (O_1358,N_9981,N_9728);
nor UO_1359 (O_1359,N_9625,N_9983);
nor UO_1360 (O_1360,N_9679,N_9561);
nor UO_1361 (O_1361,N_9822,N_9957);
or UO_1362 (O_1362,N_9585,N_9520);
and UO_1363 (O_1363,N_9950,N_9554);
nor UO_1364 (O_1364,N_9560,N_9740);
nor UO_1365 (O_1365,N_9948,N_9607);
nor UO_1366 (O_1366,N_9638,N_9894);
nand UO_1367 (O_1367,N_9511,N_9599);
and UO_1368 (O_1368,N_9599,N_9787);
nand UO_1369 (O_1369,N_9695,N_9516);
nor UO_1370 (O_1370,N_9597,N_9754);
or UO_1371 (O_1371,N_9786,N_9815);
and UO_1372 (O_1372,N_9966,N_9674);
nor UO_1373 (O_1373,N_9587,N_9781);
nor UO_1374 (O_1374,N_9939,N_9987);
or UO_1375 (O_1375,N_9896,N_9716);
or UO_1376 (O_1376,N_9984,N_9514);
nor UO_1377 (O_1377,N_9898,N_9562);
and UO_1378 (O_1378,N_9802,N_9567);
or UO_1379 (O_1379,N_9947,N_9786);
and UO_1380 (O_1380,N_9903,N_9902);
nand UO_1381 (O_1381,N_9645,N_9784);
nand UO_1382 (O_1382,N_9808,N_9636);
or UO_1383 (O_1383,N_9520,N_9613);
nand UO_1384 (O_1384,N_9509,N_9560);
and UO_1385 (O_1385,N_9849,N_9948);
and UO_1386 (O_1386,N_9933,N_9850);
xnor UO_1387 (O_1387,N_9649,N_9885);
or UO_1388 (O_1388,N_9805,N_9560);
nand UO_1389 (O_1389,N_9671,N_9538);
nand UO_1390 (O_1390,N_9845,N_9504);
nor UO_1391 (O_1391,N_9996,N_9922);
nand UO_1392 (O_1392,N_9993,N_9678);
nor UO_1393 (O_1393,N_9917,N_9711);
and UO_1394 (O_1394,N_9708,N_9836);
nand UO_1395 (O_1395,N_9636,N_9847);
nand UO_1396 (O_1396,N_9854,N_9838);
nor UO_1397 (O_1397,N_9998,N_9881);
nor UO_1398 (O_1398,N_9844,N_9769);
and UO_1399 (O_1399,N_9901,N_9749);
or UO_1400 (O_1400,N_9622,N_9613);
nand UO_1401 (O_1401,N_9534,N_9506);
and UO_1402 (O_1402,N_9918,N_9628);
and UO_1403 (O_1403,N_9642,N_9519);
nand UO_1404 (O_1404,N_9823,N_9578);
or UO_1405 (O_1405,N_9763,N_9909);
and UO_1406 (O_1406,N_9815,N_9759);
and UO_1407 (O_1407,N_9565,N_9816);
nand UO_1408 (O_1408,N_9725,N_9858);
nor UO_1409 (O_1409,N_9923,N_9769);
nor UO_1410 (O_1410,N_9503,N_9859);
or UO_1411 (O_1411,N_9938,N_9569);
or UO_1412 (O_1412,N_9599,N_9975);
nand UO_1413 (O_1413,N_9685,N_9605);
nand UO_1414 (O_1414,N_9534,N_9556);
nor UO_1415 (O_1415,N_9637,N_9749);
nor UO_1416 (O_1416,N_9713,N_9510);
nand UO_1417 (O_1417,N_9671,N_9701);
or UO_1418 (O_1418,N_9595,N_9870);
or UO_1419 (O_1419,N_9513,N_9734);
nor UO_1420 (O_1420,N_9758,N_9809);
or UO_1421 (O_1421,N_9841,N_9815);
nand UO_1422 (O_1422,N_9972,N_9507);
or UO_1423 (O_1423,N_9565,N_9691);
and UO_1424 (O_1424,N_9840,N_9931);
nand UO_1425 (O_1425,N_9729,N_9825);
nor UO_1426 (O_1426,N_9960,N_9681);
nand UO_1427 (O_1427,N_9694,N_9863);
or UO_1428 (O_1428,N_9651,N_9778);
and UO_1429 (O_1429,N_9893,N_9733);
nand UO_1430 (O_1430,N_9710,N_9583);
xnor UO_1431 (O_1431,N_9504,N_9573);
nand UO_1432 (O_1432,N_9682,N_9872);
nor UO_1433 (O_1433,N_9686,N_9738);
nor UO_1434 (O_1434,N_9600,N_9647);
or UO_1435 (O_1435,N_9773,N_9545);
and UO_1436 (O_1436,N_9848,N_9978);
and UO_1437 (O_1437,N_9824,N_9876);
nand UO_1438 (O_1438,N_9553,N_9667);
and UO_1439 (O_1439,N_9896,N_9556);
and UO_1440 (O_1440,N_9895,N_9903);
xnor UO_1441 (O_1441,N_9824,N_9943);
or UO_1442 (O_1442,N_9708,N_9586);
nand UO_1443 (O_1443,N_9584,N_9626);
nor UO_1444 (O_1444,N_9736,N_9746);
xor UO_1445 (O_1445,N_9522,N_9683);
nand UO_1446 (O_1446,N_9570,N_9502);
nor UO_1447 (O_1447,N_9645,N_9847);
or UO_1448 (O_1448,N_9667,N_9671);
or UO_1449 (O_1449,N_9544,N_9667);
and UO_1450 (O_1450,N_9685,N_9672);
and UO_1451 (O_1451,N_9529,N_9797);
nor UO_1452 (O_1452,N_9790,N_9621);
and UO_1453 (O_1453,N_9666,N_9680);
or UO_1454 (O_1454,N_9826,N_9887);
nand UO_1455 (O_1455,N_9855,N_9880);
nor UO_1456 (O_1456,N_9705,N_9864);
nor UO_1457 (O_1457,N_9519,N_9916);
nand UO_1458 (O_1458,N_9654,N_9706);
nand UO_1459 (O_1459,N_9645,N_9531);
nor UO_1460 (O_1460,N_9881,N_9566);
nand UO_1461 (O_1461,N_9583,N_9781);
xor UO_1462 (O_1462,N_9868,N_9701);
or UO_1463 (O_1463,N_9635,N_9845);
or UO_1464 (O_1464,N_9584,N_9833);
nor UO_1465 (O_1465,N_9625,N_9689);
nor UO_1466 (O_1466,N_9572,N_9829);
and UO_1467 (O_1467,N_9824,N_9639);
nor UO_1468 (O_1468,N_9707,N_9785);
nand UO_1469 (O_1469,N_9896,N_9728);
or UO_1470 (O_1470,N_9750,N_9861);
xor UO_1471 (O_1471,N_9946,N_9515);
and UO_1472 (O_1472,N_9799,N_9716);
and UO_1473 (O_1473,N_9709,N_9925);
nor UO_1474 (O_1474,N_9704,N_9718);
nor UO_1475 (O_1475,N_9811,N_9827);
or UO_1476 (O_1476,N_9775,N_9826);
and UO_1477 (O_1477,N_9718,N_9662);
nor UO_1478 (O_1478,N_9608,N_9533);
nor UO_1479 (O_1479,N_9661,N_9882);
xor UO_1480 (O_1480,N_9942,N_9707);
and UO_1481 (O_1481,N_9869,N_9580);
and UO_1482 (O_1482,N_9931,N_9735);
nor UO_1483 (O_1483,N_9889,N_9783);
and UO_1484 (O_1484,N_9568,N_9573);
or UO_1485 (O_1485,N_9924,N_9808);
and UO_1486 (O_1486,N_9814,N_9906);
nor UO_1487 (O_1487,N_9822,N_9541);
and UO_1488 (O_1488,N_9597,N_9724);
or UO_1489 (O_1489,N_9549,N_9555);
xnor UO_1490 (O_1490,N_9621,N_9964);
or UO_1491 (O_1491,N_9526,N_9842);
nor UO_1492 (O_1492,N_9992,N_9828);
nor UO_1493 (O_1493,N_9964,N_9978);
and UO_1494 (O_1494,N_9526,N_9573);
xnor UO_1495 (O_1495,N_9651,N_9614);
and UO_1496 (O_1496,N_9808,N_9846);
nand UO_1497 (O_1497,N_9706,N_9824);
nand UO_1498 (O_1498,N_9819,N_9920);
nor UO_1499 (O_1499,N_9543,N_9880);
endmodule