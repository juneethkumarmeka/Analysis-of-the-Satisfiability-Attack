module basic_1000_10000_1500_50_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
xor U0 (N_0,In_699,In_929);
and U1 (N_1,In_571,In_847);
and U2 (N_2,In_229,In_4);
xor U3 (N_3,In_899,In_761);
nand U4 (N_4,In_428,In_215);
nand U5 (N_5,In_327,In_9);
or U6 (N_6,In_454,In_719);
nand U7 (N_7,In_968,In_722);
nand U8 (N_8,In_592,In_599);
xnor U9 (N_9,In_377,In_160);
or U10 (N_10,In_708,In_411);
nand U11 (N_11,In_101,In_283);
or U12 (N_12,In_629,In_568);
nor U13 (N_13,In_560,In_725);
xnor U14 (N_14,In_831,In_365);
and U15 (N_15,In_903,In_881);
and U16 (N_16,In_689,In_777);
nand U17 (N_17,In_432,In_256);
nand U18 (N_18,In_973,In_760);
and U19 (N_19,In_298,In_805);
xor U20 (N_20,In_88,In_322);
xor U21 (N_21,In_29,In_75);
nand U22 (N_22,In_729,In_124);
nand U23 (N_23,In_112,In_195);
nand U24 (N_24,In_506,In_44);
nor U25 (N_25,In_300,In_717);
nor U26 (N_26,In_301,In_208);
and U27 (N_27,In_214,In_996);
nor U28 (N_28,In_196,In_133);
xor U29 (N_29,In_334,In_100);
and U30 (N_30,In_255,In_467);
and U31 (N_31,In_625,In_447);
nand U32 (N_32,In_343,In_634);
and U33 (N_33,In_509,In_995);
and U34 (N_34,In_466,In_745);
and U35 (N_35,In_993,In_740);
and U36 (N_36,In_217,In_249);
nor U37 (N_37,In_615,In_886);
nor U38 (N_38,In_767,In_547);
nand U39 (N_39,In_892,In_86);
xor U40 (N_40,In_230,In_170);
or U41 (N_41,In_700,In_320);
nand U42 (N_42,In_176,In_856);
and U43 (N_43,In_731,In_724);
nand U44 (N_44,In_905,In_434);
or U45 (N_45,In_34,In_464);
or U46 (N_46,In_51,In_122);
or U47 (N_47,In_969,In_280);
nor U48 (N_48,In_129,In_706);
or U49 (N_49,In_356,In_790);
nand U50 (N_50,In_89,In_656);
and U51 (N_51,In_505,In_750);
and U52 (N_52,In_303,In_335);
nor U53 (N_53,In_998,In_585);
and U54 (N_54,In_458,In_739);
nor U55 (N_55,In_74,In_928);
or U56 (N_56,In_999,In_545);
nor U57 (N_57,In_792,In_671);
nor U58 (N_58,In_940,In_429);
and U59 (N_59,In_288,In_476);
nand U60 (N_60,In_286,In_667);
nor U61 (N_61,In_198,In_223);
nor U62 (N_62,In_936,In_31);
or U63 (N_63,In_960,In_561);
nand U64 (N_64,In_226,In_801);
nor U65 (N_65,In_983,In_636);
nor U66 (N_66,In_380,In_147);
xor U67 (N_67,In_73,In_420);
and U68 (N_68,In_949,In_498);
xor U69 (N_69,In_497,In_493);
nand U70 (N_70,In_788,In_457);
or U71 (N_71,In_108,In_979);
nand U72 (N_72,In_342,In_179);
nor U73 (N_73,In_162,In_981);
or U74 (N_74,In_473,In_682);
or U75 (N_75,In_184,In_536);
nand U76 (N_76,In_621,In_985);
and U77 (N_77,In_810,In_190);
or U78 (N_78,In_475,In_237);
or U79 (N_79,In_837,In_694);
and U80 (N_80,In_394,In_10);
xor U81 (N_81,In_811,In_60);
xor U82 (N_82,In_462,In_838);
and U83 (N_83,In_988,In_382);
nand U84 (N_84,In_539,In_550);
nand U85 (N_85,In_309,In_486);
or U86 (N_86,In_879,In_62);
nor U87 (N_87,In_491,In_633);
nand U88 (N_88,In_832,In_850);
nand U89 (N_89,In_353,In_390);
or U90 (N_90,In_372,In_143);
and U91 (N_91,In_645,In_818);
nand U92 (N_92,In_35,In_480);
nand U93 (N_93,In_69,In_630);
xnor U94 (N_94,In_665,In_514);
or U95 (N_95,In_271,In_520);
nor U96 (N_96,In_889,In_576);
nor U97 (N_97,In_922,In_172);
nand U98 (N_98,In_180,In_772);
and U99 (N_99,In_906,In_734);
xnor U100 (N_100,In_310,In_670);
nor U101 (N_101,In_116,In_209);
xnor U102 (N_102,In_105,In_71);
and U103 (N_103,In_530,In_118);
or U104 (N_104,In_293,In_167);
or U105 (N_105,In_183,In_130);
nand U106 (N_106,In_613,In_808);
and U107 (N_107,In_225,In_367);
or U108 (N_108,In_527,In_938);
nand U109 (N_109,In_165,In_7);
or U110 (N_110,In_726,In_859);
or U111 (N_111,In_845,In_588);
and U112 (N_112,In_925,In_674);
nor U113 (N_113,In_851,In_931);
nor U114 (N_114,In_533,In_94);
nand U115 (N_115,In_142,In_554);
or U116 (N_116,In_774,In_933);
or U117 (N_117,In_265,In_581);
and U118 (N_118,In_274,In_809);
nor U119 (N_119,In_824,In_948);
or U120 (N_120,In_41,In_417);
and U121 (N_121,In_295,In_250);
and U122 (N_122,In_471,In_867);
or U123 (N_123,In_840,In_970);
and U124 (N_124,In_148,In_125);
or U125 (N_125,In_376,In_266);
nor U126 (N_126,In_556,In_854);
nor U127 (N_127,In_291,In_104);
nand U128 (N_128,In_600,In_747);
nor U129 (N_129,In_84,In_954);
or U130 (N_130,In_984,In_543);
or U131 (N_131,In_333,In_437);
xor U132 (N_132,In_934,In_238);
or U133 (N_133,In_595,In_780);
nand U134 (N_134,In_953,In_644);
or U135 (N_135,In_451,In_399);
nand U136 (N_136,In_405,In_641);
xor U137 (N_137,In_32,In_696);
nand U138 (N_138,In_139,In_529);
and U139 (N_139,In_594,In_83);
or U140 (N_140,In_684,In_381);
or U141 (N_141,In_623,In_446);
and U142 (N_142,In_308,In_589);
xor U143 (N_143,In_95,In_64);
or U144 (N_144,In_487,In_431);
nor U145 (N_145,In_526,In_285);
and U146 (N_146,In_566,In_637);
nor U147 (N_147,In_445,In_393);
nor U148 (N_148,In_721,In_324);
and U149 (N_149,In_593,In_81);
and U150 (N_150,In_779,In_501);
nor U151 (N_151,In_224,In_140);
or U152 (N_152,In_676,In_26);
nor U153 (N_153,In_338,In_268);
nand U154 (N_154,In_314,In_197);
nand U155 (N_155,In_369,In_806);
or U156 (N_156,In_153,In_789);
nand U157 (N_157,In_289,In_874);
and U158 (N_158,In_281,In_987);
nor U159 (N_159,In_956,In_478);
nor U160 (N_160,In_307,In_751);
nor U161 (N_161,In_37,In_80);
or U162 (N_162,In_695,In_609);
nand U163 (N_163,In_680,In_489);
nor U164 (N_164,In_681,In_963);
nor U165 (N_165,In_959,In_330);
or U166 (N_166,In_650,In_756);
nor U167 (N_167,In_952,In_614);
nand U168 (N_168,In_549,In_632);
and U169 (N_169,In_598,In_540);
nand U170 (N_170,In_188,In_785);
and U171 (N_171,In_241,In_628);
nor U172 (N_172,In_50,In_297);
nor U173 (N_173,In_397,In_880);
xor U174 (N_174,In_482,In_242);
nand U175 (N_175,In_575,In_231);
or U176 (N_176,In_765,In_299);
nor U177 (N_177,In_586,In_173);
and U178 (N_178,In_485,In_422);
or U179 (N_179,In_220,In_61);
or U180 (N_180,In_456,In_317);
nor U181 (N_181,In_145,In_775);
xor U182 (N_182,In_396,In_384);
and U183 (N_183,In_150,In_19);
or U184 (N_184,In_587,In_111);
nand U185 (N_185,In_77,In_76);
and U186 (N_186,In_305,In_164);
nand U187 (N_187,In_292,In_776);
or U188 (N_188,In_862,In_559);
and U189 (N_189,In_541,In_759);
or U190 (N_190,In_660,In_358);
and U191 (N_191,In_608,In_710);
or U192 (N_192,In_52,In_245);
nor U193 (N_193,In_98,In_407);
and U194 (N_194,In_276,In_516);
nor U195 (N_195,In_33,In_815);
and U196 (N_196,In_804,In_882);
nand U197 (N_197,In_821,In_638);
or U198 (N_198,In_647,In_402);
or U199 (N_199,In_414,In_0);
nand U200 (N_200,In_677,In_657);
xnor U201 (N_201,In_70,In_38);
or U202 (N_202,In_40,In_182);
nand U203 (N_203,In_222,N_144);
and U204 (N_204,In_323,In_313);
nand U205 (N_205,In_945,In_930);
or U206 (N_206,In_835,N_26);
xnor U207 (N_207,In_639,In_221);
nand U208 (N_208,N_154,N_189);
xor U209 (N_209,In_799,In_107);
and U210 (N_210,In_528,In_749);
nand U211 (N_211,In_311,N_89);
nand U212 (N_212,N_93,In_131);
nor U213 (N_213,N_59,In_897);
and U214 (N_214,In_386,In_513);
nand U215 (N_215,In_891,N_90);
nand U216 (N_216,N_188,In_387);
nor U217 (N_217,In_843,N_17);
or U218 (N_218,In_36,In_758);
nand U219 (N_219,In_186,In_730);
and U220 (N_220,In_910,In_860);
or U221 (N_221,N_56,In_814);
or U222 (N_222,In_273,In_79);
nor U223 (N_223,In_490,In_427);
and U224 (N_224,In_768,In_918);
xnor U225 (N_225,In_328,In_290);
nand U226 (N_226,N_3,N_57);
nor U227 (N_227,In_654,In_355);
or U228 (N_228,In_55,In_865);
nor U229 (N_229,In_715,N_11);
and U230 (N_230,In_379,In_612);
or U231 (N_231,N_39,In_714);
nor U232 (N_232,In_904,In_635);
nor U233 (N_233,In_213,In_319);
nand U234 (N_234,In_601,In_793);
nand U235 (N_235,In_460,N_162);
or U236 (N_236,In_784,In_169);
nor U237 (N_237,In_53,In_24);
nor U238 (N_238,N_49,In_896);
nand U239 (N_239,In_911,In_735);
or U240 (N_240,In_3,In_495);
nand U241 (N_241,In_45,N_178);
nand U242 (N_242,In_248,In_653);
and U243 (N_243,In_522,In_339);
nor U244 (N_244,In_701,In_120);
nor U245 (N_245,In_117,In_275);
or U246 (N_246,In_425,In_866);
nor U247 (N_247,In_158,In_114);
nor U248 (N_248,In_590,N_190);
nand U249 (N_249,In_22,In_483);
nand U250 (N_250,N_160,N_199);
nor U251 (N_251,In_385,In_174);
or U252 (N_252,In_395,In_375);
nand U253 (N_253,In_371,In_263);
or U254 (N_254,In_737,N_66);
nor U255 (N_255,In_240,In_618);
nand U256 (N_256,In_49,In_762);
nand U257 (N_257,In_119,N_121);
nor U258 (N_258,In_449,N_73);
nor U259 (N_259,N_136,In_869);
nand U260 (N_260,In_398,N_191);
nor U261 (N_261,N_142,In_78);
and U262 (N_262,N_132,In_67);
nand U263 (N_263,N_183,In_191);
or U264 (N_264,In_610,In_361);
or U265 (N_265,In_259,In_573);
nand U266 (N_266,In_894,In_461);
or U267 (N_267,In_484,In_193);
or U268 (N_268,N_38,N_64);
nor U269 (N_269,N_75,In_577);
and U270 (N_270,N_14,In_606);
or U271 (N_271,In_1,N_29);
or U272 (N_272,In_68,N_130);
or U273 (N_273,In_964,In_678);
and U274 (N_274,In_252,N_45);
or U275 (N_275,In_698,In_803);
and U276 (N_276,In_262,In_450);
nor U277 (N_277,In_110,In_63);
xor U278 (N_278,In_878,In_885);
nor U279 (N_279,N_194,In_771);
nor U280 (N_280,N_177,N_71);
xor U281 (N_281,In_781,In_651);
or U282 (N_282,In_65,In_820);
nor U283 (N_283,In_852,N_69);
or U284 (N_284,In_604,In_423);
xnor U285 (N_285,In_965,In_261);
nor U286 (N_286,In_919,In_42);
and U287 (N_287,In_349,N_184);
nor U288 (N_288,In_134,In_341);
nor U289 (N_289,In_738,In_519);
nor U290 (N_290,In_154,In_284);
and U291 (N_291,In_421,N_131);
nor U292 (N_292,In_424,N_88);
nor U293 (N_293,In_302,In_216);
or U294 (N_294,In_849,In_18);
or U295 (N_295,In_400,In_942);
nand U296 (N_296,In_469,In_544);
or U297 (N_297,In_702,In_754);
or U298 (N_298,In_875,In_151);
nand U299 (N_299,In_916,In_87);
and U300 (N_300,In_603,In_825);
nand U301 (N_301,N_13,In_944);
and U302 (N_302,In_254,In_138);
or U303 (N_303,In_212,N_161);
nand U304 (N_304,In_488,In_870);
and U305 (N_305,In_17,In_580);
or U306 (N_306,In_927,In_524);
nand U307 (N_307,In_496,N_117);
xor U308 (N_308,In_796,In_202);
or U309 (N_309,In_523,In_102);
and U310 (N_310,In_971,In_504);
or U311 (N_311,In_872,N_134);
nor U312 (N_312,In_640,In_807);
nand U313 (N_313,In_842,In_378);
xnor U314 (N_314,In_345,In_572);
or U315 (N_315,N_33,N_129);
or U316 (N_316,In_937,In_786);
or U317 (N_317,In_900,N_21);
and U318 (N_318,In_157,In_136);
or U319 (N_319,In_43,In_989);
or U320 (N_320,In_672,N_163);
nor U321 (N_321,N_139,In_200);
nand U322 (N_322,In_746,In_362);
or U323 (N_323,In_797,In_13);
nand U324 (N_324,N_67,N_197);
xnor U325 (N_325,In_769,In_264);
nor U326 (N_326,In_713,In_459);
nand U327 (N_327,In_902,N_78);
nand U328 (N_328,In_72,N_76);
nor U329 (N_329,In_673,In_711);
nor U330 (N_330,In_823,N_138);
and U331 (N_331,In_113,In_23);
or U332 (N_332,In_166,In_864);
and U333 (N_333,In_558,In_413);
and U334 (N_334,In_410,In_913);
nor U335 (N_335,In_247,In_373);
nor U336 (N_336,In_690,In_631);
or U337 (N_337,In_201,In_535);
nor U338 (N_338,In_939,In_648);
and U339 (N_339,N_62,In_419);
nand U340 (N_340,In_602,N_51);
and U341 (N_341,In_359,In_439);
nor U342 (N_342,In_861,In_794);
nor U343 (N_343,N_115,In_619);
nor U344 (N_344,N_149,In_346);
and U345 (N_345,In_622,In_697);
and U346 (N_346,In_551,In_115);
nor U347 (N_347,In_763,In_350);
nor U348 (N_348,In_525,In_463);
or U349 (N_349,In_178,In_582);
or U350 (N_350,N_152,N_173);
and U351 (N_351,In_752,N_135);
or U352 (N_352,In_584,In_203);
nand U353 (N_353,In_364,In_663);
and U354 (N_354,N_146,N_148);
nor U355 (N_355,In_884,In_227);
and U356 (N_356,In_474,In_20);
or U357 (N_357,In_12,N_106);
nand U358 (N_358,In_720,In_627);
and U359 (N_359,N_53,In_958);
nor U360 (N_360,In_507,In_967);
nand U361 (N_361,In_253,In_277);
or U362 (N_362,In_950,N_27);
or U363 (N_363,In_211,In_348);
nand U364 (N_364,In_974,N_99);
nor U365 (N_365,In_830,In_5);
or U366 (N_366,In_25,In_982);
or U367 (N_367,In_783,In_992);
xnor U368 (N_368,In_883,In_552);
xor U369 (N_369,N_179,In_659);
or U370 (N_370,In_909,In_972);
or U371 (N_371,In_205,In_438);
and U372 (N_372,In_146,In_827);
nor U373 (N_373,N_150,N_84);
nand U374 (N_374,In_453,In_961);
xnor U375 (N_375,In_742,In_66);
nor U376 (N_376,In_517,In_591);
and U377 (N_377,In_718,In_58);
and U378 (N_378,In_733,In_579);
nor U379 (N_379,In_537,N_116);
nor U380 (N_380,N_123,In_468);
nor U381 (N_381,In_39,In_403);
or U382 (N_382,N_68,In_819);
nor U383 (N_383,In_887,In_683);
xor U384 (N_384,In_531,In_748);
xnor U385 (N_385,In_626,In_351);
and U386 (N_386,N_113,In_272);
and U387 (N_387,In_546,In_6);
or U388 (N_388,In_914,In_16);
nor U389 (N_389,In_855,In_773);
and U390 (N_390,In_744,N_1);
nor U391 (N_391,In_316,N_185);
nor U392 (N_392,In_315,N_155);
nand U393 (N_393,In_137,In_688);
nand U394 (N_394,In_340,In_947);
xor U395 (N_395,In_616,In_121);
nand U396 (N_396,In_374,In_207);
or U397 (N_397,In_723,In_416);
and U398 (N_398,In_267,In_28);
or U399 (N_399,N_153,N_37);
nand U400 (N_400,In_443,In_787);
and U401 (N_401,In_318,In_123);
nand U402 (N_402,In_181,N_256);
or U403 (N_403,In_452,In_563);
and U404 (N_404,In_703,In_596);
nand U405 (N_405,In_898,N_377);
and U406 (N_406,N_362,In_56);
nand U407 (N_407,N_25,N_207);
nor U408 (N_408,N_320,In_912);
nand U409 (N_409,In_848,In_442);
and U410 (N_410,N_237,N_107);
nor U411 (N_411,N_329,In_778);
xnor U412 (N_412,N_128,N_4);
nand U413 (N_413,N_32,In_357);
or U414 (N_414,N_7,N_280);
or U415 (N_415,N_55,N_205);
and U416 (N_416,In_177,In_477);
or U417 (N_417,N_60,N_100);
and U418 (N_418,In_126,In_620);
or U419 (N_419,In_347,In_567);
or U420 (N_420,In_415,In_92);
nor U421 (N_421,N_327,In_834);
or U422 (N_422,In_664,N_42);
and U423 (N_423,In_857,N_345);
nor U424 (N_424,N_311,In_921);
nand U425 (N_425,N_157,N_200);
or U426 (N_426,N_286,N_18);
and U427 (N_427,In_234,In_243);
or U428 (N_428,In_926,In_500);
nor U429 (N_429,In_135,N_367);
or U430 (N_430,N_247,In_175);
and U431 (N_431,In_93,N_373);
and U432 (N_432,N_364,N_334);
nor U433 (N_433,In_409,N_211);
nand U434 (N_434,N_250,In_236);
and U435 (N_435,N_398,N_341);
nand U436 (N_436,N_277,N_394);
xor U437 (N_437,In_646,In_85);
nand U438 (N_438,In_941,In_669);
nand U439 (N_439,N_231,In_728);
or U440 (N_440,N_103,In_279);
nand U441 (N_441,N_166,In_901);
and U442 (N_442,N_360,In_149);
and U443 (N_443,N_215,N_314);
or U444 (N_444,In_757,In_990);
nor U445 (N_445,N_272,N_384);
xor U446 (N_446,In_344,N_225);
nor U447 (N_447,N_343,In_455);
nand U448 (N_448,In_235,N_118);
nand U449 (N_449,In_753,In_643);
nand U450 (N_450,N_101,N_288);
nand U451 (N_451,In_232,N_259);
nor U452 (N_452,N_257,N_318);
or U453 (N_453,N_98,In_841);
nand U454 (N_454,In_705,In_888);
nand U455 (N_455,N_383,In_920);
and U456 (N_456,N_16,N_19);
nand U457 (N_457,In_408,N_358);
nand U458 (N_458,N_213,In_185);
and U459 (N_459,N_43,N_308);
nor U460 (N_460,N_326,In_336);
nand U461 (N_461,N_251,N_285);
and U462 (N_462,N_376,N_380);
and U463 (N_463,N_241,N_397);
and U464 (N_464,In_510,N_63);
or U465 (N_465,N_47,N_340);
nor U466 (N_466,N_175,In_957);
nand U467 (N_467,N_87,N_104);
xor U468 (N_468,N_263,N_143);
nand U469 (N_469,In_997,N_206);
nand U470 (N_470,In_388,N_307);
or U471 (N_471,N_70,N_208);
and U472 (N_472,In_481,In_538);
and U473 (N_473,In_441,In_2);
and U474 (N_474,In_57,In_795);
nor U475 (N_475,N_344,In_189);
or U476 (N_476,In_233,N_141);
and U477 (N_477,N_281,N_95);
nor U478 (N_478,In_194,N_391);
nand U479 (N_479,N_319,In_278);
nor U480 (N_480,In_955,N_172);
and U481 (N_481,N_258,In_569);
xor U482 (N_482,N_393,In_833);
or U483 (N_483,In_144,N_105);
or U484 (N_484,In_48,N_292);
and U485 (N_485,In_534,N_357);
and U486 (N_486,In_470,In_27);
and U487 (N_487,N_266,In_99);
nor U488 (N_488,In_868,N_289);
and U489 (N_489,N_15,N_369);
and U490 (N_490,In_210,In_15);
nor U491 (N_491,N_366,In_691);
nor U492 (N_492,N_333,N_174);
nor U493 (N_493,N_375,N_214);
and U494 (N_494,In_935,In_521);
or U495 (N_495,N_24,In_152);
and U496 (N_496,N_268,N_198);
and U497 (N_497,In_515,N_79);
or U498 (N_498,In_30,N_94);
nor U499 (N_499,In_11,N_176);
nor U500 (N_500,In_564,In_966);
and U501 (N_501,In_943,N_335);
nor U502 (N_502,In_917,N_270);
nand U503 (N_503,In_976,In_326);
or U504 (N_504,In_331,In_923);
and U505 (N_505,N_159,N_296);
or U506 (N_506,N_316,In_611);
and U507 (N_507,N_192,N_5);
or U508 (N_508,In_132,N_92);
nor U509 (N_509,N_267,N_204);
nand U510 (N_510,N_242,N_388);
or U511 (N_511,In_685,In_895);
and U512 (N_512,In_97,In_363);
and U513 (N_513,In_876,In_192);
xnor U514 (N_514,In_816,In_389);
or U515 (N_515,N_252,N_239);
nor U516 (N_516,N_244,N_127);
nand U517 (N_517,In_562,In_46);
nor U518 (N_518,N_8,N_58);
or U519 (N_519,N_120,In_658);
and U520 (N_520,N_226,N_309);
and U521 (N_521,In_155,N_303);
nor U522 (N_522,In_736,N_86);
or U523 (N_523,N_186,N_193);
nand U524 (N_524,In_479,In_828);
nor U525 (N_525,N_390,N_392);
nor U526 (N_526,N_119,N_342);
nand U527 (N_527,N_321,In_583);
nand U528 (N_528,N_140,In_649);
nand U529 (N_529,In_716,N_238);
nor U530 (N_530,In_401,N_167);
or U531 (N_531,In_444,In_542);
nand U532 (N_532,In_607,N_352);
and U533 (N_533,In_82,N_379);
and U534 (N_534,N_269,N_182);
and U535 (N_535,N_96,In_21);
nor U536 (N_536,N_228,In_103);
or U537 (N_537,In_839,In_709);
or U538 (N_538,N_54,In_962);
nand U539 (N_539,N_112,N_355);
nand U540 (N_540,In_652,N_295);
or U541 (N_541,In_47,In_829);
or U542 (N_542,N_304,In_127);
nor U543 (N_543,In_741,In_624);
nor U544 (N_544,N_254,N_363);
xor U545 (N_545,In_570,In_666);
and U546 (N_546,N_298,In_448);
or U547 (N_547,N_31,N_34);
nor U548 (N_548,N_108,In_418);
and U549 (N_549,In_873,N_300);
or U550 (N_550,In_846,In_802);
or U551 (N_551,N_168,In_404);
and U552 (N_552,In_204,N_378);
and U553 (N_553,N_253,N_137);
and U554 (N_554,N_399,In_433);
nor U555 (N_555,In_218,In_858);
nor U556 (N_556,N_354,N_156);
nor U557 (N_557,N_293,In_109);
or U558 (N_558,In_260,N_349);
xor U559 (N_559,N_328,In_662);
or U560 (N_560,In_156,N_124);
nand U561 (N_561,In_332,N_243);
xor U562 (N_562,In_508,In_743);
or U563 (N_563,In_863,N_28);
nor U564 (N_564,In_270,N_82);
nand U565 (N_565,N_312,In_435);
or U566 (N_566,N_227,N_386);
xor U567 (N_567,In_893,In_383);
nand U568 (N_568,In_368,In_391);
and U569 (N_569,N_332,N_249);
nor U570 (N_570,N_10,In_54);
or U571 (N_571,In_686,N_35);
and U572 (N_572,N_387,In_986);
or U573 (N_573,In_755,In_246);
and U574 (N_574,In_426,In_732);
and U575 (N_575,In_96,In_791);
and U576 (N_576,N_271,In_915);
and U577 (N_577,N_232,In_321);
nor U578 (N_578,N_283,In_159);
or U579 (N_579,N_158,In_548);
nor U580 (N_580,N_222,In_472);
and U581 (N_581,N_246,In_555);
and U582 (N_582,In_171,In_199);
or U583 (N_583,N_170,N_210);
or U584 (N_584,In_727,N_126);
nand U585 (N_585,N_9,N_306);
nand U586 (N_586,N_236,In_430);
nor U587 (N_587,In_932,N_61);
nor U588 (N_588,In_91,N_290);
and U589 (N_589,N_336,N_111);
nor U590 (N_590,In_128,N_133);
and U591 (N_591,N_353,N_77);
xor U592 (N_592,N_125,N_151);
xnor U593 (N_593,N_181,N_284);
nand U594 (N_594,N_164,N_248);
nor U595 (N_595,N_324,In_853);
nand U596 (N_596,In_813,N_356);
and U597 (N_597,N_233,N_169);
or U598 (N_598,In_844,In_597);
nand U599 (N_599,In_502,In_675);
nand U600 (N_600,In_800,N_570);
and U601 (N_601,N_432,In_578);
or U602 (N_602,N_553,N_580);
or U603 (N_603,In_518,N_408);
nor U604 (N_604,N_2,In_392);
or U605 (N_605,In_494,N_419);
and U606 (N_606,N_548,In_239);
nor U607 (N_607,N_550,N_368);
nand U608 (N_608,N_540,N_109);
and U609 (N_609,In_782,N_401);
and U610 (N_610,N_509,N_374);
xor U611 (N_611,N_382,N_371);
nand U612 (N_612,N_485,N_209);
nand U613 (N_613,N_547,N_424);
nor U614 (N_614,In_257,N_171);
xnor U615 (N_615,In_354,N_585);
nand U616 (N_616,N_522,In_465);
and U617 (N_617,N_537,In_163);
and U618 (N_618,N_274,N_464);
and U619 (N_619,In_994,In_106);
and U620 (N_620,N_582,In_924);
or U621 (N_621,N_219,N_499);
or U622 (N_622,N_531,N_91);
and U623 (N_623,N_240,N_450);
xnor U624 (N_624,N_512,N_552);
nor U625 (N_625,N_317,In_492);
and U626 (N_626,N_483,In_282);
or U627 (N_627,N_110,N_560);
nor U628 (N_628,N_6,N_489);
or U629 (N_629,N_437,In_168);
or U630 (N_630,In_141,N_347);
and U631 (N_631,N_313,N_261);
or U632 (N_632,N_404,N_504);
nor U633 (N_633,N_491,In_704);
nor U634 (N_634,N_574,N_438);
or U635 (N_635,N_97,N_557);
and U636 (N_636,N_330,In_977);
and U637 (N_637,N_264,In_978);
or U638 (N_638,N_513,N_425);
nand U639 (N_639,N_440,N_466);
or U640 (N_640,N_488,N_279);
or U641 (N_641,N_229,In_565);
nand U642 (N_642,N_403,In_436);
nor U643 (N_643,In_412,N_455);
xnor U644 (N_644,N_331,N_433);
nand U645 (N_645,N_589,N_577);
and U646 (N_646,N_381,N_508);
nor U647 (N_647,N_402,N_396);
nor U648 (N_648,In_269,N_559);
or U649 (N_649,N_551,N_83);
nor U650 (N_650,N_365,In_287);
nand U651 (N_651,In_161,N_224);
nor U652 (N_652,N_569,N_370);
xor U653 (N_653,In_766,In_764);
or U654 (N_654,N_202,N_555);
or U655 (N_655,N_417,N_596);
and U656 (N_656,N_72,N_262);
or U657 (N_657,N_481,N_544);
nor U658 (N_658,N_418,In_532);
xor U659 (N_659,N_12,In_366);
nand U660 (N_660,N_278,N_497);
nand U661 (N_661,N_102,N_50);
nand U662 (N_662,N_505,N_460);
or U663 (N_663,In_337,In_14);
and U664 (N_664,N_275,N_452);
or U665 (N_665,N_471,N_30);
or U666 (N_666,N_546,N_468);
and U667 (N_667,N_543,N_498);
or U668 (N_668,N_315,In_975);
or U669 (N_669,N_525,N_434);
and U670 (N_670,N_573,N_385);
nand U671 (N_671,N_482,N_422);
nand U672 (N_672,N_457,N_479);
and U673 (N_673,In_770,N_36);
or U674 (N_674,In_244,N_415);
nand U675 (N_675,In_642,N_530);
or U676 (N_676,N_597,In_826);
and U677 (N_677,N_542,N_445);
or U678 (N_678,N_245,N_411);
nor U679 (N_679,N_421,N_494);
or U680 (N_680,N_591,N_523);
or U681 (N_681,N_359,N_446);
and U682 (N_682,N_564,N_412);
or U683 (N_683,In_219,N_431);
or U684 (N_684,N_495,N_65);
nor U685 (N_685,In_306,N_114);
nor U686 (N_686,N_212,N_443);
xor U687 (N_687,N_590,N_429);
nand U688 (N_688,N_350,N_456);
nand U689 (N_689,N_500,N_515);
nor U690 (N_690,N_348,N_592);
or U691 (N_691,N_441,N_524);
nor U692 (N_692,N_463,N_389);
nand U693 (N_693,N_294,N_430);
nand U694 (N_694,In_352,In_679);
nor U695 (N_695,N_510,N_444);
or U696 (N_696,N_218,N_486);
nor U697 (N_697,In_228,In_655);
and U698 (N_698,N_147,In_187);
or U699 (N_699,N_493,In_499);
or U700 (N_700,N_310,N_223);
and U701 (N_701,N_536,In_8);
xor U702 (N_702,In_707,N_521);
nand U703 (N_703,In_511,N_302);
or U704 (N_704,N_563,N_351);
nand U705 (N_705,N_565,N_195);
xor U706 (N_706,N_187,N_492);
or U707 (N_707,N_416,N_587);
xor U708 (N_708,N_46,In_687);
xor U709 (N_709,N_273,N_576);
or U710 (N_710,In_991,N_322);
nand U711 (N_711,N_282,N_230);
nand U712 (N_712,N_473,N_407);
or U713 (N_713,N_23,N_556);
nand U714 (N_714,N_538,N_52);
nor U715 (N_715,N_80,N_567);
and U716 (N_716,In_258,N_413);
and U717 (N_717,N_299,N_516);
or U718 (N_718,In_693,N_474);
or U719 (N_719,N_490,N_406);
or U720 (N_720,In_817,In_692);
xnor U721 (N_721,N_532,N_453);
or U722 (N_722,N_235,N_287);
nand U723 (N_723,In_574,N_558);
or U724 (N_724,In_503,N_517);
nor U725 (N_725,N_581,In_557);
nor U726 (N_726,N_511,N_451);
nand U727 (N_727,N_442,N_599);
nand U728 (N_728,N_484,N_507);
nor U729 (N_729,In_908,N_48);
and U730 (N_730,In_370,In_296);
nand U731 (N_731,N_276,N_220);
xor U732 (N_732,N_514,N_420);
and U733 (N_733,In_877,In_294);
or U734 (N_734,N_44,N_426);
and U735 (N_735,N_568,In_605);
and U736 (N_736,In_325,N_575);
nor U737 (N_737,N_122,In_206);
or U738 (N_738,N_461,In_661);
nor U739 (N_739,N_260,In_406);
nor U740 (N_740,N_454,N_462);
and U741 (N_741,N_400,N_584);
nor U742 (N_742,N_337,In_304);
nand U743 (N_743,N_323,In_360);
or U744 (N_744,N_165,N_566);
and U745 (N_745,N_554,N_447);
and U746 (N_746,N_561,N_203);
nand U747 (N_747,In_712,N_467);
or U748 (N_748,N_361,N_541);
nor U749 (N_749,N_503,N_217);
nand U750 (N_750,In_90,N_519);
and U751 (N_751,N_562,N_586);
nor U752 (N_752,N_325,N_305);
nand U753 (N_753,N_534,N_529);
or U754 (N_754,N_145,N_472);
and U755 (N_755,N_85,N_265);
nand U756 (N_756,In_871,N_0);
and U757 (N_757,N_469,In_512);
or U758 (N_758,N_234,N_439);
nor U759 (N_759,N_539,In_251);
nor U760 (N_760,N_449,N_81);
or U761 (N_761,N_496,N_527);
nand U762 (N_762,N_40,N_571);
nor U763 (N_763,N_410,N_572);
nor U764 (N_764,N_477,N_475);
and U765 (N_765,N_520,N_409);
and U766 (N_766,In_668,N_346);
nor U767 (N_767,In_553,N_518);
or U768 (N_768,In_812,N_338);
or U769 (N_769,In_951,N_395);
xnor U770 (N_770,N_526,In_980);
or U771 (N_771,In_312,N_423);
nand U772 (N_772,N_428,N_549);
xnor U773 (N_773,N_405,N_372);
or U774 (N_774,N_427,N_578);
nand U775 (N_775,N_20,N_476);
nor U776 (N_776,N_448,N_594);
and U777 (N_777,In_822,In_907);
nand U778 (N_778,N_22,N_291);
or U779 (N_779,N_502,N_435);
nor U780 (N_780,In_798,N_583);
nand U781 (N_781,N_339,N_588);
nor U782 (N_782,In_329,N_528);
and U783 (N_783,N_593,N_579);
nor U784 (N_784,N_458,N_480);
nand U785 (N_785,In_946,N_74);
xnor U786 (N_786,N_255,N_201);
or U787 (N_787,N_535,N_506);
nor U788 (N_788,N_414,N_41);
or U789 (N_789,N_465,N_221);
nor U790 (N_790,N_598,N_180);
nor U791 (N_791,N_196,N_545);
nor U792 (N_792,N_216,In_836);
nor U793 (N_793,N_459,N_595);
nor U794 (N_794,N_297,N_436);
nand U795 (N_795,N_301,In_440);
nor U796 (N_796,N_470,In_890);
nor U797 (N_797,N_478,N_487);
nand U798 (N_798,N_533,N_501);
and U799 (N_799,In_59,In_617);
or U800 (N_800,N_771,N_689);
nand U801 (N_801,N_617,N_731);
and U802 (N_802,N_740,N_652);
nand U803 (N_803,N_751,N_753);
nand U804 (N_804,N_668,N_749);
nand U805 (N_805,N_685,N_793);
nand U806 (N_806,N_755,N_759);
or U807 (N_807,N_664,N_710);
or U808 (N_808,N_775,N_687);
nand U809 (N_809,N_741,N_767);
or U810 (N_810,N_641,N_762);
or U811 (N_811,N_728,N_746);
xnor U812 (N_812,N_774,N_736);
nor U813 (N_813,N_661,N_783);
or U814 (N_814,N_708,N_795);
nor U815 (N_815,N_672,N_675);
or U816 (N_816,N_602,N_693);
nand U817 (N_817,N_765,N_626);
nand U818 (N_818,N_628,N_779);
nor U819 (N_819,N_622,N_797);
and U820 (N_820,N_657,N_656);
nand U821 (N_821,N_629,N_787);
and U822 (N_822,N_607,N_704);
nand U823 (N_823,N_663,N_676);
or U824 (N_824,N_703,N_620);
or U825 (N_825,N_729,N_630);
and U826 (N_826,N_651,N_621);
or U827 (N_827,N_606,N_719);
nand U828 (N_828,N_730,N_711);
and U829 (N_829,N_723,N_792);
nand U830 (N_830,N_667,N_677);
and U831 (N_831,N_690,N_776);
and U832 (N_832,N_697,N_724);
or U833 (N_833,N_758,N_642);
or U834 (N_834,N_698,N_678);
nand U835 (N_835,N_768,N_600);
or U836 (N_836,N_782,N_739);
xnor U837 (N_837,N_613,N_713);
and U838 (N_838,N_737,N_682);
and U839 (N_839,N_674,N_718);
xor U840 (N_840,N_785,N_650);
nand U841 (N_841,N_794,N_754);
nor U842 (N_842,N_761,N_684);
or U843 (N_843,N_618,N_688);
or U844 (N_844,N_743,N_638);
or U845 (N_845,N_766,N_700);
nand U846 (N_846,N_624,N_614);
or U847 (N_847,N_694,N_679);
nand U848 (N_848,N_760,N_757);
or U849 (N_849,N_778,N_715);
nor U850 (N_850,N_721,N_712);
nor U851 (N_851,N_786,N_605);
nor U852 (N_852,N_633,N_784);
and U853 (N_853,N_640,N_735);
or U854 (N_854,N_662,N_714);
and U855 (N_855,N_699,N_601);
xnor U856 (N_856,N_645,N_635);
and U857 (N_857,N_763,N_658);
or U858 (N_858,N_649,N_732);
nand U859 (N_859,N_655,N_643);
nand U860 (N_860,N_752,N_709);
nand U861 (N_861,N_799,N_659);
or U862 (N_862,N_734,N_727);
nand U863 (N_863,N_673,N_632);
xnor U864 (N_864,N_634,N_750);
or U865 (N_865,N_608,N_702);
or U866 (N_866,N_791,N_637);
nand U867 (N_867,N_660,N_773);
or U868 (N_868,N_669,N_747);
or U869 (N_869,N_625,N_716);
xnor U870 (N_870,N_627,N_619);
nand U871 (N_871,N_646,N_665);
or U872 (N_872,N_722,N_604);
nor U873 (N_873,N_733,N_680);
nor U874 (N_874,N_796,N_720);
nand U875 (N_875,N_612,N_744);
and U876 (N_876,N_648,N_790);
nor U877 (N_877,N_725,N_742);
or U878 (N_878,N_798,N_777);
nand U879 (N_879,N_696,N_789);
or U880 (N_880,N_683,N_707);
and U881 (N_881,N_701,N_653);
nor U882 (N_882,N_644,N_738);
or U883 (N_883,N_616,N_654);
and U884 (N_884,N_781,N_686);
xor U885 (N_885,N_636,N_615);
nor U886 (N_886,N_610,N_706);
and U887 (N_887,N_671,N_745);
or U888 (N_888,N_772,N_695);
or U889 (N_889,N_691,N_631);
or U890 (N_890,N_769,N_623);
nand U891 (N_891,N_764,N_647);
nor U892 (N_892,N_603,N_666);
nand U893 (N_893,N_681,N_756);
nand U894 (N_894,N_717,N_639);
xnor U895 (N_895,N_780,N_726);
xnor U896 (N_896,N_609,N_692);
nor U897 (N_897,N_705,N_770);
xor U898 (N_898,N_748,N_788);
nor U899 (N_899,N_670,N_611);
nor U900 (N_900,N_703,N_762);
nor U901 (N_901,N_728,N_708);
or U902 (N_902,N_663,N_787);
and U903 (N_903,N_600,N_710);
or U904 (N_904,N_681,N_679);
or U905 (N_905,N_699,N_788);
and U906 (N_906,N_696,N_678);
and U907 (N_907,N_757,N_613);
nor U908 (N_908,N_741,N_705);
xnor U909 (N_909,N_620,N_640);
or U910 (N_910,N_713,N_743);
and U911 (N_911,N_775,N_769);
and U912 (N_912,N_782,N_794);
nand U913 (N_913,N_793,N_725);
and U914 (N_914,N_674,N_620);
nand U915 (N_915,N_643,N_759);
xor U916 (N_916,N_785,N_704);
nand U917 (N_917,N_710,N_603);
and U918 (N_918,N_748,N_660);
and U919 (N_919,N_628,N_790);
nor U920 (N_920,N_651,N_712);
and U921 (N_921,N_696,N_773);
or U922 (N_922,N_738,N_799);
nor U923 (N_923,N_784,N_623);
xor U924 (N_924,N_780,N_605);
nor U925 (N_925,N_719,N_723);
nand U926 (N_926,N_687,N_752);
or U927 (N_927,N_693,N_617);
nor U928 (N_928,N_701,N_627);
nor U929 (N_929,N_715,N_635);
nand U930 (N_930,N_719,N_644);
nor U931 (N_931,N_772,N_614);
nand U932 (N_932,N_777,N_662);
xnor U933 (N_933,N_720,N_750);
nor U934 (N_934,N_674,N_787);
nand U935 (N_935,N_763,N_641);
xor U936 (N_936,N_625,N_600);
nand U937 (N_937,N_792,N_786);
nand U938 (N_938,N_725,N_731);
nand U939 (N_939,N_797,N_600);
nand U940 (N_940,N_717,N_749);
and U941 (N_941,N_689,N_716);
nor U942 (N_942,N_612,N_607);
nand U943 (N_943,N_775,N_737);
and U944 (N_944,N_746,N_783);
and U945 (N_945,N_653,N_740);
nand U946 (N_946,N_637,N_673);
and U947 (N_947,N_697,N_660);
and U948 (N_948,N_797,N_645);
or U949 (N_949,N_627,N_787);
nor U950 (N_950,N_660,N_669);
or U951 (N_951,N_715,N_705);
xnor U952 (N_952,N_769,N_709);
nor U953 (N_953,N_619,N_704);
or U954 (N_954,N_792,N_657);
or U955 (N_955,N_699,N_748);
or U956 (N_956,N_744,N_707);
and U957 (N_957,N_685,N_644);
or U958 (N_958,N_654,N_650);
nor U959 (N_959,N_745,N_694);
and U960 (N_960,N_715,N_736);
nand U961 (N_961,N_659,N_719);
xnor U962 (N_962,N_680,N_785);
nor U963 (N_963,N_681,N_778);
or U964 (N_964,N_617,N_609);
nor U965 (N_965,N_742,N_720);
or U966 (N_966,N_701,N_724);
nand U967 (N_967,N_664,N_633);
or U968 (N_968,N_738,N_688);
or U969 (N_969,N_669,N_706);
or U970 (N_970,N_682,N_710);
or U971 (N_971,N_697,N_677);
and U972 (N_972,N_648,N_680);
nand U973 (N_973,N_610,N_612);
and U974 (N_974,N_766,N_774);
nor U975 (N_975,N_736,N_693);
or U976 (N_976,N_745,N_747);
nand U977 (N_977,N_703,N_741);
nor U978 (N_978,N_649,N_725);
or U979 (N_979,N_616,N_615);
nand U980 (N_980,N_742,N_635);
nand U981 (N_981,N_736,N_682);
and U982 (N_982,N_742,N_784);
or U983 (N_983,N_602,N_764);
nor U984 (N_984,N_719,N_736);
and U985 (N_985,N_730,N_739);
and U986 (N_986,N_601,N_786);
nor U987 (N_987,N_767,N_698);
xor U988 (N_988,N_672,N_719);
and U989 (N_989,N_672,N_713);
nand U990 (N_990,N_782,N_710);
nand U991 (N_991,N_776,N_671);
xnor U992 (N_992,N_793,N_676);
and U993 (N_993,N_777,N_684);
nand U994 (N_994,N_638,N_632);
xor U995 (N_995,N_720,N_708);
or U996 (N_996,N_607,N_646);
nor U997 (N_997,N_757,N_603);
and U998 (N_998,N_747,N_606);
nand U999 (N_999,N_760,N_776);
or U1000 (N_1000,N_832,N_869);
nand U1001 (N_1001,N_939,N_895);
or U1002 (N_1002,N_828,N_920);
nor U1003 (N_1003,N_944,N_838);
or U1004 (N_1004,N_931,N_877);
and U1005 (N_1005,N_922,N_867);
or U1006 (N_1006,N_926,N_996);
and U1007 (N_1007,N_824,N_839);
or U1008 (N_1008,N_883,N_863);
or U1009 (N_1009,N_943,N_881);
nor U1010 (N_1010,N_882,N_803);
and U1011 (N_1011,N_983,N_800);
nand U1012 (N_1012,N_880,N_802);
and U1013 (N_1013,N_970,N_988);
nor U1014 (N_1014,N_887,N_974);
nand U1015 (N_1015,N_874,N_999);
nand U1016 (N_1016,N_907,N_950);
and U1017 (N_1017,N_915,N_989);
or U1018 (N_1018,N_963,N_976);
xor U1019 (N_1019,N_973,N_866);
and U1020 (N_1020,N_918,N_891);
nor U1021 (N_1021,N_959,N_987);
or U1022 (N_1022,N_940,N_985);
xnor U1023 (N_1023,N_814,N_945);
nor U1024 (N_1024,N_840,N_825);
and U1025 (N_1025,N_892,N_933);
nand U1026 (N_1026,N_835,N_914);
or U1027 (N_1027,N_951,N_902);
and U1028 (N_1028,N_911,N_893);
nand U1029 (N_1029,N_859,N_809);
nor U1030 (N_1030,N_971,N_962);
nand U1031 (N_1031,N_896,N_878);
nor U1032 (N_1032,N_956,N_995);
or U1033 (N_1033,N_879,N_831);
nor U1034 (N_1034,N_834,N_975);
nand U1035 (N_1035,N_868,N_948);
and U1036 (N_1036,N_848,N_849);
or U1037 (N_1037,N_827,N_936);
or U1038 (N_1038,N_841,N_934);
or U1039 (N_1039,N_826,N_829);
or U1040 (N_1040,N_861,N_870);
and U1041 (N_1041,N_818,N_901);
or U1042 (N_1042,N_855,N_935);
or U1043 (N_1043,N_967,N_949);
and U1044 (N_1044,N_994,N_919);
or U1045 (N_1045,N_952,N_913);
and U1046 (N_1046,N_889,N_972);
or U1047 (N_1047,N_924,N_958);
and U1048 (N_1048,N_860,N_847);
and U1049 (N_1049,N_925,N_890);
nand U1050 (N_1050,N_853,N_982);
and U1051 (N_1051,N_977,N_888);
and U1052 (N_1052,N_937,N_816);
nor U1053 (N_1053,N_897,N_843);
or U1054 (N_1054,N_928,N_905);
nand U1055 (N_1055,N_822,N_852);
nor U1056 (N_1056,N_904,N_986);
and U1057 (N_1057,N_961,N_854);
and U1058 (N_1058,N_871,N_929);
xor U1059 (N_1059,N_965,N_885);
and U1060 (N_1060,N_865,N_836);
and U1061 (N_1061,N_993,N_968);
and U1062 (N_1062,N_906,N_991);
or U1063 (N_1063,N_923,N_953);
nand U1064 (N_1064,N_805,N_947);
xor U1065 (N_1065,N_984,N_856);
nand U1066 (N_1066,N_864,N_842);
or U1067 (N_1067,N_980,N_857);
nor U1068 (N_1068,N_899,N_804);
nand U1069 (N_1069,N_812,N_969);
nor U1070 (N_1070,N_844,N_938);
xor U1071 (N_1071,N_964,N_921);
nor U1072 (N_1072,N_978,N_917);
or U1073 (N_1073,N_815,N_801);
and U1074 (N_1074,N_916,N_872);
nand U1075 (N_1075,N_846,N_908);
nand U1076 (N_1076,N_912,N_900);
nand U1077 (N_1077,N_817,N_910);
and U1078 (N_1078,N_909,N_941);
or U1079 (N_1079,N_990,N_837);
or U1080 (N_1080,N_946,N_979);
nand U1081 (N_1081,N_873,N_807);
nor U1082 (N_1082,N_875,N_955);
nor U1083 (N_1083,N_813,N_820);
or U1084 (N_1084,N_957,N_806);
nand U1085 (N_1085,N_862,N_992);
nor U1086 (N_1086,N_927,N_894);
or U1087 (N_1087,N_960,N_932);
xnor U1088 (N_1088,N_903,N_954);
and U1089 (N_1089,N_808,N_898);
xnor U1090 (N_1090,N_930,N_886);
nor U1091 (N_1091,N_810,N_819);
nor U1092 (N_1092,N_884,N_845);
or U1093 (N_1093,N_830,N_833);
nor U1094 (N_1094,N_850,N_966);
nor U1095 (N_1095,N_997,N_942);
and U1096 (N_1096,N_858,N_811);
and U1097 (N_1097,N_821,N_876);
and U1098 (N_1098,N_823,N_998);
nand U1099 (N_1099,N_851,N_981);
or U1100 (N_1100,N_881,N_946);
or U1101 (N_1101,N_809,N_989);
xor U1102 (N_1102,N_951,N_980);
or U1103 (N_1103,N_982,N_905);
and U1104 (N_1104,N_843,N_834);
nor U1105 (N_1105,N_885,N_820);
and U1106 (N_1106,N_987,N_991);
nor U1107 (N_1107,N_872,N_999);
nand U1108 (N_1108,N_865,N_924);
nand U1109 (N_1109,N_955,N_879);
or U1110 (N_1110,N_853,N_842);
or U1111 (N_1111,N_995,N_949);
or U1112 (N_1112,N_934,N_853);
and U1113 (N_1113,N_887,N_848);
and U1114 (N_1114,N_801,N_990);
nand U1115 (N_1115,N_901,N_914);
or U1116 (N_1116,N_924,N_976);
or U1117 (N_1117,N_851,N_826);
nor U1118 (N_1118,N_927,N_950);
and U1119 (N_1119,N_974,N_962);
xor U1120 (N_1120,N_966,N_864);
nand U1121 (N_1121,N_871,N_901);
xor U1122 (N_1122,N_971,N_819);
nor U1123 (N_1123,N_894,N_823);
or U1124 (N_1124,N_954,N_930);
or U1125 (N_1125,N_865,N_892);
xor U1126 (N_1126,N_919,N_921);
and U1127 (N_1127,N_859,N_990);
and U1128 (N_1128,N_942,N_900);
nand U1129 (N_1129,N_949,N_894);
nor U1130 (N_1130,N_820,N_974);
nand U1131 (N_1131,N_894,N_832);
nor U1132 (N_1132,N_977,N_865);
nand U1133 (N_1133,N_803,N_852);
nor U1134 (N_1134,N_922,N_914);
nor U1135 (N_1135,N_801,N_997);
xnor U1136 (N_1136,N_849,N_898);
nor U1137 (N_1137,N_934,N_918);
or U1138 (N_1138,N_824,N_807);
or U1139 (N_1139,N_807,N_988);
and U1140 (N_1140,N_974,N_904);
xor U1141 (N_1141,N_921,N_935);
and U1142 (N_1142,N_966,N_888);
or U1143 (N_1143,N_931,N_851);
nor U1144 (N_1144,N_812,N_852);
nor U1145 (N_1145,N_859,N_985);
xnor U1146 (N_1146,N_881,N_815);
nand U1147 (N_1147,N_945,N_863);
and U1148 (N_1148,N_905,N_901);
or U1149 (N_1149,N_917,N_921);
xor U1150 (N_1150,N_889,N_953);
xnor U1151 (N_1151,N_868,N_835);
or U1152 (N_1152,N_951,N_906);
nor U1153 (N_1153,N_990,N_806);
and U1154 (N_1154,N_861,N_865);
nor U1155 (N_1155,N_896,N_974);
nand U1156 (N_1156,N_912,N_993);
or U1157 (N_1157,N_840,N_810);
and U1158 (N_1158,N_935,N_818);
nand U1159 (N_1159,N_960,N_890);
and U1160 (N_1160,N_931,N_808);
nand U1161 (N_1161,N_932,N_878);
nor U1162 (N_1162,N_838,N_901);
xnor U1163 (N_1163,N_847,N_983);
and U1164 (N_1164,N_941,N_842);
and U1165 (N_1165,N_826,N_941);
nor U1166 (N_1166,N_914,N_879);
nor U1167 (N_1167,N_958,N_949);
nand U1168 (N_1168,N_950,N_976);
and U1169 (N_1169,N_821,N_975);
or U1170 (N_1170,N_961,N_800);
and U1171 (N_1171,N_815,N_940);
or U1172 (N_1172,N_949,N_916);
and U1173 (N_1173,N_886,N_996);
or U1174 (N_1174,N_856,N_803);
and U1175 (N_1175,N_903,N_981);
xnor U1176 (N_1176,N_842,N_800);
nor U1177 (N_1177,N_948,N_837);
nand U1178 (N_1178,N_931,N_827);
or U1179 (N_1179,N_844,N_995);
nor U1180 (N_1180,N_837,N_812);
and U1181 (N_1181,N_930,N_924);
or U1182 (N_1182,N_878,N_852);
nor U1183 (N_1183,N_960,N_813);
or U1184 (N_1184,N_839,N_846);
nand U1185 (N_1185,N_834,N_938);
nor U1186 (N_1186,N_990,N_863);
nor U1187 (N_1187,N_807,N_902);
nand U1188 (N_1188,N_880,N_849);
nor U1189 (N_1189,N_818,N_807);
or U1190 (N_1190,N_977,N_972);
nand U1191 (N_1191,N_857,N_816);
nand U1192 (N_1192,N_924,N_949);
nand U1193 (N_1193,N_874,N_855);
nor U1194 (N_1194,N_887,N_944);
nand U1195 (N_1195,N_967,N_812);
nand U1196 (N_1196,N_891,N_831);
nand U1197 (N_1197,N_849,N_870);
and U1198 (N_1198,N_860,N_806);
or U1199 (N_1199,N_961,N_919);
or U1200 (N_1200,N_1109,N_1028);
and U1201 (N_1201,N_1130,N_1129);
nand U1202 (N_1202,N_1018,N_1146);
or U1203 (N_1203,N_1140,N_1196);
or U1204 (N_1204,N_1041,N_1147);
nand U1205 (N_1205,N_1004,N_1183);
or U1206 (N_1206,N_1088,N_1185);
nor U1207 (N_1207,N_1163,N_1046);
nand U1208 (N_1208,N_1173,N_1000);
or U1209 (N_1209,N_1091,N_1067);
xnor U1210 (N_1210,N_1022,N_1124);
nand U1211 (N_1211,N_1081,N_1118);
nor U1212 (N_1212,N_1195,N_1178);
nor U1213 (N_1213,N_1034,N_1103);
and U1214 (N_1214,N_1056,N_1058);
nand U1215 (N_1215,N_1112,N_1015);
xnor U1216 (N_1216,N_1110,N_1136);
nand U1217 (N_1217,N_1098,N_1092);
nor U1218 (N_1218,N_1125,N_1165);
and U1219 (N_1219,N_1024,N_1199);
xor U1220 (N_1220,N_1038,N_1187);
and U1221 (N_1221,N_1055,N_1079);
and U1222 (N_1222,N_1037,N_1114);
and U1223 (N_1223,N_1005,N_1174);
nor U1224 (N_1224,N_1138,N_1181);
nand U1225 (N_1225,N_1193,N_1194);
or U1226 (N_1226,N_1019,N_1083);
nor U1227 (N_1227,N_1189,N_1116);
nand U1228 (N_1228,N_1117,N_1197);
xnor U1229 (N_1229,N_1107,N_1061);
and U1230 (N_1230,N_1084,N_1052);
or U1231 (N_1231,N_1074,N_1105);
xnor U1232 (N_1232,N_1035,N_1011);
and U1233 (N_1233,N_1069,N_1085);
nand U1234 (N_1234,N_1127,N_1065);
nand U1235 (N_1235,N_1198,N_1106);
and U1236 (N_1236,N_1145,N_1134);
nor U1237 (N_1237,N_1190,N_1184);
nand U1238 (N_1238,N_1104,N_1167);
and U1239 (N_1239,N_1172,N_1021);
or U1240 (N_1240,N_1076,N_1119);
or U1241 (N_1241,N_1009,N_1144);
nor U1242 (N_1242,N_1168,N_1157);
or U1243 (N_1243,N_1100,N_1066);
nor U1244 (N_1244,N_1156,N_1006);
and U1245 (N_1245,N_1108,N_1096);
xor U1246 (N_1246,N_1082,N_1169);
and U1247 (N_1247,N_1139,N_1036);
or U1248 (N_1248,N_1072,N_1075);
nand U1249 (N_1249,N_1008,N_1095);
nand U1250 (N_1250,N_1164,N_1120);
or U1251 (N_1251,N_1048,N_1045);
nand U1252 (N_1252,N_1151,N_1152);
or U1253 (N_1253,N_1161,N_1182);
nor U1254 (N_1254,N_1115,N_1097);
and U1255 (N_1255,N_1070,N_1054);
or U1256 (N_1256,N_1063,N_1012);
nand U1257 (N_1257,N_1122,N_1123);
xor U1258 (N_1258,N_1062,N_1071);
nand U1259 (N_1259,N_1007,N_1044);
or U1260 (N_1260,N_1162,N_1064);
nor U1261 (N_1261,N_1078,N_1020);
or U1262 (N_1262,N_1059,N_1040);
nor U1263 (N_1263,N_1025,N_1027);
nand U1264 (N_1264,N_1073,N_1188);
or U1265 (N_1265,N_1159,N_1090);
and U1266 (N_1266,N_1013,N_1016);
or U1267 (N_1267,N_1039,N_1179);
and U1268 (N_1268,N_1155,N_1128);
nor U1269 (N_1269,N_1029,N_1014);
and U1270 (N_1270,N_1137,N_1002);
and U1271 (N_1271,N_1031,N_1099);
nor U1272 (N_1272,N_1017,N_1087);
or U1273 (N_1273,N_1121,N_1033);
nand U1274 (N_1274,N_1160,N_1135);
or U1275 (N_1275,N_1047,N_1166);
and U1276 (N_1276,N_1143,N_1043);
nor U1277 (N_1277,N_1171,N_1060);
or U1278 (N_1278,N_1089,N_1026);
and U1279 (N_1279,N_1094,N_1113);
and U1280 (N_1280,N_1175,N_1042);
nand U1281 (N_1281,N_1053,N_1102);
nor U1282 (N_1282,N_1186,N_1050);
or U1283 (N_1283,N_1051,N_1003);
and U1284 (N_1284,N_1142,N_1176);
nand U1285 (N_1285,N_1149,N_1154);
nand U1286 (N_1286,N_1023,N_1158);
nor U1287 (N_1287,N_1030,N_1057);
nor U1288 (N_1288,N_1068,N_1192);
nand U1289 (N_1289,N_1170,N_1133);
nand U1290 (N_1290,N_1126,N_1141);
or U1291 (N_1291,N_1080,N_1180);
and U1292 (N_1292,N_1150,N_1049);
xnor U1293 (N_1293,N_1032,N_1077);
nand U1294 (N_1294,N_1111,N_1001);
xnor U1295 (N_1295,N_1132,N_1177);
nor U1296 (N_1296,N_1086,N_1093);
nand U1297 (N_1297,N_1191,N_1153);
nor U1298 (N_1298,N_1101,N_1131);
or U1299 (N_1299,N_1148,N_1010);
nand U1300 (N_1300,N_1023,N_1170);
or U1301 (N_1301,N_1096,N_1069);
and U1302 (N_1302,N_1076,N_1107);
nor U1303 (N_1303,N_1027,N_1042);
and U1304 (N_1304,N_1181,N_1001);
nand U1305 (N_1305,N_1056,N_1006);
xor U1306 (N_1306,N_1186,N_1030);
nor U1307 (N_1307,N_1126,N_1165);
nor U1308 (N_1308,N_1095,N_1117);
or U1309 (N_1309,N_1149,N_1148);
nand U1310 (N_1310,N_1162,N_1012);
or U1311 (N_1311,N_1079,N_1148);
xor U1312 (N_1312,N_1015,N_1133);
and U1313 (N_1313,N_1125,N_1134);
xnor U1314 (N_1314,N_1133,N_1162);
nor U1315 (N_1315,N_1160,N_1106);
nor U1316 (N_1316,N_1066,N_1048);
nand U1317 (N_1317,N_1024,N_1033);
nor U1318 (N_1318,N_1066,N_1185);
xor U1319 (N_1319,N_1112,N_1145);
or U1320 (N_1320,N_1038,N_1181);
nor U1321 (N_1321,N_1044,N_1113);
and U1322 (N_1322,N_1046,N_1174);
nor U1323 (N_1323,N_1052,N_1170);
nor U1324 (N_1324,N_1019,N_1180);
nor U1325 (N_1325,N_1055,N_1086);
or U1326 (N_1326,N_1176,N_1144);
or U1327 (N_1327,N_1169,N_1006);
or U1328 (N_1328,N_1069,N_1145);
or U1329 (N_1329,N_1146,N_1088);
and U1330 (N_1330,N_1044,N_1171);
nand U1331 (N_1331,N_1154,N_1081);
nand U1332 (N_1332,N_1086,N_1021);
or U1333 (N_1333,N_1000,N_1163);
nand U1334 (N_1334,N_1123,N_1019);
nor U1335 (N_1335,N_1167,N_1138);
nand U1336 (N_1336,N_1045,N_1097);
and U1337 (N_1337,N_1152,N_1192);
xor U1338 (N_1338,N_1195,N_1133);
or U1339 (N_1339,N_1078,N_1127);
xor U1340 (N_1340,N_1199,N_1046);
and U1341 (N_1341,N_1058,N_1046);
nor U1342 (N_1342,N_1090,N_1197);
xnor U1343 (N_1343,N_1172,N_1002);
or U1344 (N_1344,N_1128,N_1182);
and U1345 (N_1345,N_1002,N_1187);
nor U1346 (N_1346,N_1077,N_1047);
or U1347 (N_1347,N_1022,N_1106);
and U1348 (N_1348,N_1116,N_1156);
and U1349 (N_1349,N_1070,N_1020);
nand U1350 (N_1350,N_1031,N_1159);
or U1351 (N_1351,N_1093,N_1047);
nor U1352 (N_1352,N_1142,N_1167);
xor U1353 (N_1353,N_1150,N_1047);
nor U1354 (N_1354,N_1087,N_1161);
nor U1355 (N_1355,N_1052,N_1185);
or U1356 (N_1356,N_1106,N_1116);
and U1357 (N_1357,N_1058,N_1159);
and U1358 (N_1358,N_1018,N_1191);
nor U1359 (N_1359,N_1077,N_1001);
nand U1360 (N_1360,N_1197,N_1135);
and U1361 (N_1361,N_1037,N_1008);
nor U1362 (N_1362,N_1116,N_1147);
or U1363 (N_1363,N_1094,N_1008);
or U1364 (N_1364,N_1088,N_1123);
or U1365 (N_1365,N_1050,N_1096);
xnor U1366 (N_1366,N_1160,N_1133);
nor U1367 (N_1367,N_1046,N_1180);
nand U1368 (N_1368,N_1027,N_1034);
nand U1369 (N_1369,N_1051,N_1164);
nor U1370 (N_1370,N_1079,N_1038);
or U1371 (N_1371,N_1143,N_1121);
and U1372 (N_1372,N_1025,N_1195);
or U1373 (N_1373,N_1004,N_1184);
nand U1374 (N_1374,N_1094,N_1046);
nor U1375 (N_1375,N_1101,N_1070);
nand U1376 (N_1376,N_1149,N_1130);
nand U1377 (N_1377,N_1188,N_1082);
and U1378 (N_1378,N_1116,N_1079);
and U1379 (N_1379,N_1098,N_1108);
or U1380 (N_1380,N_1164,N_1098);
or U1381 (N_1381,N_1187,N_1026);
nand U1382 (N_1382,N_1150,N_1132);
xnor U1383 (N_1383,N_1020,N_1186);
xor U1384 (N_1384,N_1038,N_1062);
xnor U1385 (N_1385,N_1048,N_1178);
xnor U1386 (N_1386,N_1035,N_1032);
or U1387 (N_1387,N_1105,N_1184);
nor U1388 (N_1388,N_1023,N_1157);
nand U1389 (N_1389,N_1179,N_1098);
or U1390 (N_1390,N_1072,N_1043);
xnor U1391 (N_1391,N_1037,N_1123);
xnor U1392 (N_1392,N_1050,N_1150);
and U1393 (N_1393,N_1194,N_1022);
or U1394 (N_1394,N_1115,N_1122);
and U1395 (N_1395,N_1116,N_1001);
nor U1396 (N_1396,N_1058,N_1041);
and U1397 (N_1397,N_1031,N_1094);
and U1398 (N_1398,N_1162,N_1122);
and U1399 (N_1399,N_1037,N_1086);
nor U1400 (N_1400,N_1286,N_1389);
and U1401 (N_1401,N_1233,N_1330);
and U1402 (N_1402,N_1375,N_1265);
nand U1403 (N_1403,N_1316,N_1287);
and U1404 (N_1404,N_1300,N_1271);
nor U1405 (N_1405,N_1367,N_1256);
nand U1406 (N_1406,N_1273,N_1344);
or U1407 (N_1407,N_1246,N_1338);
and U1408 (N_1408,N_1226,N_1294);
xnor U1409 (N_1409,N_1295,N_1398);
or U1410 (N_1410,N_1228,N_1278);
nand U1411 (N_1411,N_1329,N_1229);
nand U1412 (N_1412,N_1303,N_1289);
or U1413 (N_1413,N_1393,N_1317);
and U1414 (N_1414,N_1282,N_1349);
and U1415 (N_1415,N_1326,N_1371);
nand U1416 (N_1416,N_1325,N_1203);
or U1417 (N_1417,N_1205,N_1202);
and U1418 (N_1418,N_1230,N_1381);
nor U1419 (N_1419,N_1264,N_1257);
and U1420 (N_1420,N_1245,N_1284);
nand U1421 (N_1421,N_1321,N_1372);
nor U1422 (N_1422,N_1259,N_1396);
nor U1423 (N_1423,N_1388,N_1281);
or U1424 (N_1424,N_1235,N_1336);
or U1425 (N_1425,N_1288,N_1204);
or U1426 (N_1426,N_1234,N_1251);
nor U1427 (N_1427,N_1266,N_1213);
nor U1428 (N_1428,N_1346,N_1353);
or U1429 (N_1429,N_1285,N_1399);
xnor U1430 (N_1430,N_1258,N_1253);
nand U1431 (N_1431,N_1387,N_1374);
or U1432 (N_1432,N_1331,N_1242);
nand U1433 (N_1433,N_1313,N_1248);
nand U1434 (N_1434,N_1223,N_1217);
nor U1435 (N_1435,N_1274,N_1267);
and U1436 (N_1436,N_1236,N_1312);
nand U1437 (N_1437,N_1322,N_1254);
or U1438 (N_1438,N_1276,N_1394);
nand U1439 (N_1439,N_1209,N_1255);
nor U1440 (N_1440,N_1260,N_1382);
nor U1441 (N_1441,N_1279,N_1351);
nand U1442 (N_1442,N_1320,N_1211);
xor U1443 (N_1443,N_1305,N_1385);
or U1444 (N_1444,N_1206,N_1333);
xnor U1445 (N_1445,N_1347,N_1306);
and U1446 (N_1446,N_1244,N_1283);
and U1447 (N_1447,N_1296,N_1359);
nor U1448 (N_1448,N_1324,N_1318);
nor U1449 (N_1449,N_1216,N_1247);
xnor U1450 (N_1450,N_1210,N_1309);
or U1451 (N_1451,N_1376,N_1231);
nand U1452 (N_1452,N_1323,N_1268);
nand U1453 (N_1453,N_1362,N_1290);
or U1454 (N_1454,N_1379,N_1249);
and U1455 (N_1455,N_1342,N_1291);
and U1456 (N_1456,N_1252,N_1332);
and U1457 (N_1457,N_1241,N_1357);
nor U1458 (N_1458,N_1315,N_1270);
nor U1459 (N_1459,N_1239,N_1299);
or U1460 (N_1460,N_1224,N_1361);
and U1461 (N_1461,N_1212,N_1201);
nor U1462 (N_1462,N_1302,N_1383);
or U1463 (N_1463,N_1238,N_1307);
nand U1464 (N_1464,N_1328,N_1352);
nor U1465 (N_1465,N_1275,N_1355);
or U1466 (N_1466,N_1222,N_1386);
or U1467 (N_1467,N_1363,N_1207);
nand U1468 (N_1468,N_1280,N_1377);
and U1469 (N_1469,N_1227,N_1218);
or U1470 (N_1470,N_1341,N_1219);
nor U1471 (N_1471,N_1215,N_1358);
nor U1472 (N_1472,N_1364,N_1380);
nor U1473 (N_1473,N_1373,N_1360);
xnor U1474 (N_1474,N_1390,N_1301);
or U1475 (N_1475,N_1269,N_1221);
nor U1476 (N_1476,N_1378,N_1277);
nand U1477 (N_1477,N_1370,N_1397);
or U1478 (N_1478,N_1337,N_1340);
nor U1479 (N_1479,N_1297,N_1308);
or U1480 (N_1480,N_1225,N_1368);
or U1481 (N_1481,N_1200,N_1237);
nand U1482 (N_1482,N_1310,N_1214);
nor U1483 (N_1483,N_1314,N_1366);
and U1484 (N_1484,N_1348,N_1369);
nor U1485 (N_1485,N_1232,N_1240);
or U1486 (N_1486,N_1384,N_1392);
and U1487 (N_1487,N_1339,N_1261);
nand U1488 (N_1488,N_1395,N_1243);
and U1489 (N_1489,N_1350,N_1293);
or U1490 (N_1490,N_1298,N_1391);
and U1491 (N_1491,N_1335,N_1311);
or U1492 (N_1492,N_1334,N_1356);
xnor U1493 (N_1493,N_1345,N_1262);
or U1494 (N_1494,N_1365,N_1272);
nor U1495 (N_1495,N_1343,N_1208);
and U1496 (N_1496,N_1292,N_1327);
nand U1497 (N_1497,N_1304,N_1354);
or U1498 (N_1498,N_1263,N_1319);
and U1499 (N_1499,N_1220,N_1250);
or U1500 (N_1500,N_1397,N_1227);
and U1501 (N_1501,N_1348,N_1218);
nor U1502 (N_1502,N_1347,N_1302);
or U1503 (N_1503,N_1355,N_1334);
or U1504 (N_1504,N_1324,N_1288);
xnor U1505 (N_1505,N_1249,N_1384);
or U1506 (N_1506,N_1299,N_1287);
and U1507 (N_1507,N_1312,N_1262);
or U1508 (N_1508,N_1202,N_1367);
nor U1509 (N_1509,N_1288,N_1265);
xnor U1510 (N_1510,N_1200,N_1229);
nand U1511 (N_1511,N_1294,N_1372);
and U1512 (N_1512,N_1244,N_1258);
nor U1513 (N_1513,N_1231,N_1285);
or U1514 (N_1514,N_1369,N_1337);
nand U1515 (N_1515,N_1336,N_1375);
nor U1516 (N_1516,N_1280,N_1317);
xor U1517 (N_1517,N_1330,N_1220);
or U1518 (N_1518,N_1331,N_1324);
nand U1519 (N_1519,N_1397,N_1304);
or U1520 (N_1520,N_1369,N_1390);
and U1521 (N_1521,N_1356,N_1254);
and U1522 (N_1522,N_1207,N_1389);
and U1523 (N_1523,N_1224,N_1366);
and U1524 (N_1524,N_1357,N_1269);
and U1525 (N_1525,N_1372,N_1267);
nand U1526 (N_1526,N_1225,N_1377);
nand U1527 (N_1527,N_1283,N_1201);
and U1528 (N_1528,N_1277,N_1252);
and U1529 (N_1529,N_1287,N_1204);
or U1530 (N_1530,N_1366,N_1277);
and U1531 (N_1531,N_1359,N_1310);
xor U1532 (N_1532,N_1255,N_1314);
and U1533 (N_1533,N_1323,N_1273);
xor U1534 (N_1534,N_1380,N_1202);
nor U1535 (N_1535,N_1326,N_1399);
and U1536 (N_1536,N_1209,N_1329);
nor U1537 (N_1537,N_1369,N_1382);
nand U1538 (N_1538,N_1216,N_1221);
and U1539 (N_1539,N_1294,N_1379);
and U1540 (N_1540,N_1242,N_1384);
xnor U1541 (N_1541,N_1374,N_1322);
and U1542 (N_1542,N_1361,N_1335);
nand U1543 (N_1543,N_1204,N_1386);
xor U1544 (N_1544,N_1373,N_1248);
and U1545 (N_1545,N_1371,N_1217);
and U1546 (N_1546,N_1347,N_1250);
and U1547 (N_1547,N_1217,N_1366);
or U1548 (N_1548,N_1213,N_1382);
and U1549 (N_1549,N_1388,N_1346);
or U1550 (N_1550,N_1297,N_1325);
nand U1551 (N_1551,N_1297,N_1291);
xnor U1552 (N_1552,N_1389,N_1382);
or U1553 (N_1553,N_1248,N_1255);
nor U1554 (N_1554,N_1250,N_1320);
xor U1555 (N_1555,N_1291,N_1302);
or U1556 (N_1556,N_1258,N_1228);
and U1557 (N_1557,N_1337,N_1254);
and U1558 (N_1558,N_1394,N_1214);
xnor U1559 (N_1559,N_1240,N_1331);
xnor U1560 (N_1560,N_1233,N_1312);
nand U1561 (N_1561,N_1253,N_1307);
nand U1562 (N_1562,N_1303,N_1291);
or U1563 (N_1563,N_1390,N_1312);
and U1564 (N_1564,N_1324,N_1310);
or U1565 (N_1565,N_1202,N_1276);
nand U1566 (N_1566,N_1230,N_1294);
nand U1567 (N_1567,N_1278,N_1239);
or U1568 (N_1568,N_1206,N_1359);
xnor U1569 (N_1569,N_1221,N_1260);
and U1570 (N_1570,N_1349,N_1352);
or U1571 (N_1571,N_1278,N_1254);
or U1572 (N_1572,N_1327,N_1268);
nand U1573 (N_1573,N_1324,N_1302);
and U1574 (N_1574,N_1371,N_1264);
nand U1575 (N_1575,N_1236,N_1396);
or U1576 (N_1576,N_1206,N_1258);
and U1577 (N_1577,N_1209,N_1261);
or U1578 (N_1578,N_1367,N_1304);
and U1579 (N_1579,N_1298,N_1354);
or U1580 (N_1580,N_1296,N_1256);
nand U1581 (N_1581,N_1245,N_1267);
and U1582 (N_1582,N_1348,N_1338);
nand U1583 (N_1583,N_1314,N_1301);
and U1584 (N_1584,N_1297,N_1272);
or U1585 (N_1585,N_1277,N_1211);
nand U1586 (N_1586,N_1231,N_1357);
nor U1587 (N_1587,N_1270,N_1250);
nor U1588 (N_1588,N_1368,N_1378);
nor U1589 (N_1589,N_1396,N_1300);
nor U1590 (N_1590,N_1251,N_1322);
and U1591 (N_1591,N_1318,N_1228);
nand U1592 (N_1592,N_1324,N_1322);
and U1593 (N_1593,N_1276,N_1228);
or U1594 (N_1594,N_1354,N_1277);
and U1595 (N_1595,N_1387,N_1247);
nand U1596 (N_1596,N_1229,N_1225);
nor U1597 (N_1597,N_1356,N_1328);
nand U1598 (N_1598,N_1342,N_1204);
nor U1599 (N_1599,N_1255,N_1219);
nor U1600 (N_1600,N_1544,N_1537);
and U1601 (N_1601,N_1578,N_1592);
nand U1602 (N_1602,N_1402,N_1561);
and U1603 (N_1603,N_1482,N_1575);
or U1604 (N_1604,N_1552,N_1485);
and U1605 (N_1605,N_1590,N_1582);
nor U1606 (N_1606,N_1464,N_1474);
or U1607 (N_1607,N_1576,N_1551);
xor U1608 (N_1608,N_1511,N_1593);
nand U1609 (N_1609,N_1441,N_1495);
and U1610 (N_1610,N_1571,N_1524);
and U1611 (N_1611,N_1505,N_1568);
xor U1612 (N_1612,N_1407,N_1420);
and U1613 (N_1613,N_1463,N_1523);
or U1614 (N_1614,N_1528,N_1480);
nand U1615 (N_1615,N_1522,N_1569);
nor U1616 (N_1616,N_1471,N_1547);
nand U1617 (N_1617,N_1581,N_1570);
nand U1618 (N_1618,N_1492,N_1428);
or U1619 (N_1619,N_1521,N_1494);
xor U1620 (N_1620,N_1510,N_1540);
or U1621 (N_1621,N_1577,N_1516);
nand U1622 (N_1622,N_1555,N_1475);
and U1623 (N_1623,N_1594,N_1451);
xor U1624 (N_1624,N_1439,N_1527);
or U1625 (N_1625,N_1560,N_1497);
nand U1626 (N_1626,N_1591,N_1586);
xnor U1627 (N_1627,N_1595,N_1583);
nand U1628 (N_1628,N_1514,N_1539);
or U1629 (N_1629,N_1449,N_1490);
nor U1630 (N_1630,N_1456,N_1409);
nor U1631 (N_1631,N_1580,N_1546);
and U1632 (N_1632,N_1432,N_1588);
or U1633 (N_1633,N_1448,N_1507);
or U1634 (N_1634,N_1424,N_1433);
nand U1635 (N_1635,N_1542,N_1419);
nand U1636 (N_1636,N_1421,N_1425);
or U1637 (N_1637,N_1440,N_1509);
nor U1638 (N_1638,N_1496,N_1556);
or U1639 (N_1639,N_1550,N_1417);
nor U1640 (N_1640,N_1403,N_1465);
nand U1641 (N_1641,N_1401,N_1435);
xnor U1642 (N_1642,N_1416,N_1526);
and U1643 (N_1643,N_1585,N_1579);
or U1644 (N_1644,N_1531,N_1442);
nor U1645 (N_1645,N_1430,N_1478);
or U1646 (N_1646,N_1541,N_1503);
nand U1647 (N_1647,N_1574,N_1437);
nor U1648 (N_1648,N_1587,N_1499);
nand U1649 (N_1649,N_1525,N_1455);
or U1650 (N_1650,N_1553,N_1512);
and U1651 (N_1651,N_1477,N_1469);
or U1652 (N_1652,N_1468,N_1484);
and U1653 (N_1653,N_1513,N_1508);
nand U1654 (N_1654,N_1502,N_1446);
and U1655 (N_1655,N_1558,N_1548);
nor U1656 (N_1656,N_1422,N_1567);
or U1657 (N_1657,N_1431,N_1452);
or U1658 (N_1658,N_1414,N_1459);
or U1659 (N_1659,N_1564,N_1434);
nand U1660 (N_1660,N_1483,N_1443);
nor U1661 (N_1661,N_1566,N_1412);
or U1662 (N_1662,N_1517,N_1519);
nor U1663 (N_1663,N_1563,N_1423);
and U1664 (N_1664,N_1534,N_1493);
and U1665 (N_1665,N_1472,N_1436);
and U1666 (N_1666,N_1445,N_1438);
and U1667 (N_1667,N_1457,N_1506);
nor U1668 (N_1668,N_1533,N_1557);
or U1669 (N_1669,N_1498,N_1406);
or U1670 (N_1670,N_1444,N_1554);
nand U1671 (N_1671,N_1460,N_1429);
nand U1672 (N_1672,N_1481,N_1486);
nor U1673 (N_1673,N_1565,N_1584);
nand U1674 (N_1674,N_1447,N_1427);
nand U1675 (N_1675,N_1411,N_1413);
and U1676 (N_1676,N_1545,N_1415);
nor U1677 (N_1677,N_1596,N_1461);
and U1678 (N_1678,N_1549,N_1562);
xor U1679 (N_1679,N_1462,N_1529);
and U1680 (N_1680,N_1426,N_1599);
and U1681 (N_1681,N_1572,N_1559);
nand U1682 (N_1682,N_1473,N_1504);
xnor U1683 (N_1683,N_1489,N_1500);
nand U1684 (N_1684,N_1598,N_1536);
nor U1685 (N_1685,N_1589,N_1501);
and U1686 (N_1686,N_1400,N_1476);
nand U1687 (N_1687,N_1543,N_1467);
nor U1688 (N_1688,N_1418,N_1532);
nor U1689 (N_1689,N_1466,N_1487);
nand U1690 (N_1690,N_1573,N_1404);
and U1691 (N_1691,N_1470,N_1408);
xnor U1692 (N_1692,N_1530,N_1518);
or U1693 (N_1693,N_1491,N_1458);
and U1694 (N_1694,N_1515,N_1453);
nand U1695 (N_1695,N_1488,N_1538);
or U1696 (N_1696,N_1597,N_1405);
and U1697 (N_1697,N_1479,N_1520);
xor U1698 (N_1698,N_1454,N_1535);
and U1699 (N_1699,N_1410,N_1450);
or U1700 (N_1700,N_1531,N_1475);
nand U1701 (N_1701,N_1580,N_1408);
and U1702 (N_1702,N_1544,N_1412);
nand U1703 (N_1703,N_1551,N_1415);
xor U1704 (N_1704,N_1475,N_1554);
xor U1705 (N_1705,N_1594,N_1471);
nor U1706 (N_1706,N_1537,N_1520);
nor U1707 (N_1707,N_1507,N_1540);
xnor U1708 (N_1708,N_1493,N_1549);
and U1709 (N_1709,N_1507,N_1579);
xor U1710 (N_1710,N_1420,N_1537);
or U1711 (N_1711,N_1449,N_1580);
nor U1712 (N_1712,N_1490,N_1451);
nor U1713 (N_1713,N_1505,N_1441);
xor U1714 (N_1714,N_1483,N_1542);
and U1715 (N_1715,N_1449,N_1486);
nand U1716 (N_1716,N_1478,N_1592);
nor U1717 (N_1717,N_1512,N_1418);
and U1718 (N_1718,N_1509,N_1463);
or U1719 (N_1719,N_1438,N_1479);
nor U1720 (N_1720,N_1456,N_1534);
nor U1721 (N_1721,N_1554,N_1495);
nand U1722 (N_1722,N_1425,N_1596);
nand U1723 (N_1723,N_1569,N_1558);
xnor U1724 (N_1724,N_1462,N_1505);
nand U1725 (N_1725,N_1567,N_1400);
nand U1726 (N_1726,N_1433,N_1469);
xnor U1727 (N_1727,N_1437,N_1533);
or U1728 (N_1728,N_1482,N_1501);
nor U1729 (N_1729,N_1474,N_1538);
nor U1730 (N_1730,N_1499,N_1562);
nand U1731 (N_1731,N_1502,N_1557);
nor U1732 (N_1732,N_1437,N_1541);
or U1733 (N_1733,N_1504,N_1514);
nor U1734 (N_1734,N_1448,N_1489);
and U1735 (N_1735,N_1555,N_1529);
and U1736 (N_1736,N_1409,N_1592);
or U1737 (N_1737,N_1554,N_1432);
nand U1738 (N_1738,N_1561,N_1509);
and U1739 (N_1739,N_1551,N_1424);
nor U1740 (N_1740,N_1542,N_1551);
and U1741 (N_1741,N_1584,N_1432);
and U1742 (N_1742,N_1460,N_1570);
nand U1743 (N_1743,N_1446,N_1596);
or U1744 (N_1744,N_1450,N_1417);
nand U1745 (N_1745,N_1487,N_1589);
nor U1746 (N_1746,N_1449,N_1561);
nand U1747 (N_1747,N_1419,N_1508);
or U1748 (N_1748,N_1480,N_1466);
nand U1749 (N_1749,N_1435,N_1441);
nor U1750 (N_1750,N_1421,N_1441);
nor U1751 (N_1751,N_1531,N_1408);
nor U1752 (N_1752,N_1429,N_1535);
xnor U1753 (N_1753,N_1442,N_1403);
nor U1754 (N_1754,N_1523,N_1508);
nand U1755 (N_1755,N_1461,N_1454);
nand U1756 (N_1756,N_1421,N_1593);
or U1757 (N_1757,N_1407,N_1584);
nand U1758 (N_1758,N_1568,N_1540);
xor U1759 (N_1759,N_1482,N_1417);
xor U1760 (N_1760,N_1423,N_1501);
xor U1761 (N_1761,N_1575,N_1577);
nor U1762 (N_1762,N_1513,N_1419);
nand U1763 (N_1763,N_1472,N_1414);
xor U1764 (N_1764,N_1407,N_1468);
nand U1765 (N_1765,N_1435,N_1565);
xor U1766 (N_1766,N_1535,N_1501);
or U1767 (N_1767,N_1412,N_1597);
nor U1768 (N_1768,N_1432,N_1537);
nand U1769 (N_1769,N_1426,N_1518);
and U1770 (N_1770,N_1419,N_1446);
and U1771 (N_1771,N_1470,N_1564);
or U1772 (N_1772,N_1572,N_1438);
or U1773 (N_1773,N_1423,N_1504);
nor U1774 (N_1774,N_1407,N_1463);
nand U1775 (N_1775,N_1516,N_1450);
xor U1776 (N_1776,N_1561,N_1549);
xnor U1777 (N_1777,N_1520,N_1477);
xor U1778 (N_1778,N_1438,N_1444);
or U1779 (N_1779,N_1452,N_1460);
or U1780 (N_1780,N_1596,N_1480);
or U1781 (N_1781,N_1587,N_1557);
or U1782 (N_1782,N_1452,N_1582);
and U1783 (N_1783,N_1498,N_1451);
or U1784 (N_1784,N_1494,N_1446);
or U1785 (N_1785,N_1471,N_1417);
and U1786 (N_1786,N_1428,N_1425);
xnor U1787 (N_1787,N_1572,N_1410);
nand U1788 (N_1788,N_1507,N_1525);
and U1789 (N_1789,N_1426,N_1477);
or U1790 (N_1790,N_1506,N_1562);
or U1791 (N_1791,N_1544,N_1507);
xor U1792 (N_1792,N_1511,N_1505);
nor U1793 (N_1793,N_1405,N_1479);
nor U1794 (N_1794,N_1408,N_1585);
or U1795 (N_1795,N_1417,N_1528);
xnor U1796 (N_1796,N_1455,N_1535);
or U1797 (N_1797,N_1527,N_1577);
and U1798 (N_1798,N_1428,N_1452);
and U1799 (N_1799,N_1597,N_1510);
and U1800 (N_1800,N_1738,N_1620);
xor U1801 (N_1801,N_1633,N_1629);
nand U1802 (N_1802,N_1721,N_1610);
or U1803 (N_1803,N_1762,N_1699);
nand U1804 (N_1804,N_1767,N_1730);
or U1805 (N_1805,N_1640,N_1717);
and U1806 (N_1806,N_1719,N_1679);
nand U1807 (N_1807,N_1630,N_1674);
nor U1808 (N_1808,N_1625,N_1771);
nand U1809 (N_1809,N_1728,N_1665);
nor U1810 (N_1810,N_1736,N_1684);
nor U1811 (N_1811,N_1723,N_1673);
nand U1812 (N_1812,N_1716,N_1713);
and U1813 (N_1813,N_1678,N_1731);
nor U1814 (N_1814,N_1754,N_1669);
or U1815 (N_1815,N_1793,N_1666);
and U1816 (N_1816,N_1656,N_1613);
and U1817 (N_1817,N_1733,N_1792);
and U1818 (N_1818,N_1745,N_1659);
nor U1819 (N_1819,N_1752,N_1744);
and U1820 (N_1820,N_1616,N_1720);
nor U1821 (N_1821,N_1794,N_1785);
nand U1822 (N_1822,N_1648,N_1769);
nor U1823 (N_1823,N_1690,N_1668);
xnor U1824 (N_1824,N_1756,N_1722);
or U1825 (N_1825,N_1710,N_1676);
nor U1826 (N_1826,N_1689,N_1761);
nand U1827 (N_1827,N_1646,N_1615);
or U1828 (N_1828,N_1639,N_1609);
or U1829 (N_1829,N_1604,N_1645);
xnor U1830 (N_1830,N_1667,N_1787);
and U1831 (N_1831,N_1628,N_1603);
nor U1832 (N_1832,N_1798,N_1724);
or U1833 (N_1833,N_1796,N_1680);
nor U1834 (N_1834,N_1618,N_1704);
or U1835 (N_1835,N_1677,N_1624);
nor U1836 (N_1836,N_1662,N_1660);
nor U1837 (N_1837,N_1619,N_1635);
nand U1838 (N_1838,N_1652,N_1779);
xor U1839 (N_1839,N_1746,N_1768);
or U1840 (N_1840,N_1750,N_1601);
nand U1841 (N_1841,N_1755,N_1627);
nor U1842 (N_1842,N_1748,N_1605);
nand U1843 (N_1843,N_1696,N_1612);
nor U1844 (N_1844,N_1644,N_1776);
and U1845 (N_1845,N_1735,N_1682);
and U1846 (N_1846,N_1760,N_1694);
or U1847 (N_1847,N_1636,N_1691);
or U1848 (N_1848,N_1751,N_1687);
xnor U1849 (N_1849,N_1661,N_1600);
nand U1850 (N_1850,N_1688,N_1715);
nor U1851 (N_1851,N_1778,N_1775);
nor U1852 (N_1852,N_1663,N_1734);
xor U1853 (N_1853,N_1718,N_1763);
nand U1854 (N_1854,N_1643,N_1693);
nor U1855 (N_1855,N_1786,N_1739);
nand U1856 (N_1856,N_1608,N_1743);
nand U1857 (N_1857,N_1758,N_1737);
nand U1858 (N_1858,N_1732,N_1714);
or U1859 (N_1859,N_1697,N_1703);
nor U1860 (N_1860,N_1607,N_1651);
nor U1861 (N_1861,N_1709,N_1638);
or U1862 (N_1862,N_1702,N_1757);
nor U1863 (N_1863,N_1654,N_1670);
xor U1864 (N_1864,N_1774,N_1614);
nor U1865 (N_1865,N_1708,N_1658);
and U1866 (N_1866,N_1695,N_1725);
or U1867 (N_1867,N_1729,N_1683);
nor U1868 (N_1868,N_1777,N_1741);
nand U1869 (N_1869,N_1780,N_1664);
and U1870 (N_1870,N_1606,N_1621);
nand U1871 (N_1871,N_1772,N_1781);
nor U1872 (N_1872,N_1782,N_1642);
nand U1873 (N_1873,N_1753,N_1602);
or U1874 (N_1874,N_1647,N_1740);
xnor U1875 (N_1875,N_1726,N_1707);
xor U1876 (N_1876,N_1742,N_1790);
nand U1877 (N_1877,N_1712,N_1773);
xnor U1878 (N_1878,N_1685,N_1770);
or U1879 (N_1879,N_1784,N_1637);
or U1880 (N_1880,N_1705,N_1765);
and U1881 (N_1881,N_1672,N_1783);
nor U1882 (N_1882,N_1655,N_1649);
xnor U1883 (N_1883,N_1611,N_1795);
nor U1884 (N_1884,N_1749,N_1692);
nor U1885 (N_1885,N_1650,N_1799);
and U1886 (N_1886,N_1622,N_1657);
or U1887 (N_1887,N_1797,N_1791);
or U1888 (N_1888,N_1759,N_1632);
and U1889 (N_1889,N_1706,N_1634);
or U1890 (N_1890,N_1698,N_1686);
nor U1891 (N_1891,N_1675,N_1711);
and U1892 (N_1892,N_1747,N_1617);
nor U1893 (N_1893,N_1626,N_1700);
and U1894 (N_1894,N_1789,N_1788);
or U1895 (N_1895,N_1681,N_1671);
and U1896 (N_1896,N_1727,N_1631);
nor U1897 (N_1897,N_1764,N_1623);
and U1898 (N_1898,N_1766,N_1641);
or U1899 (N_1899,N_1701,N_1653);
nand U1900 (N_1900,N_1702,N_1630);
and U1901 (N_1901,N_1661,N_1757);
or U1902 (N_1902,N_1664,N_1673);
nand U1903 (N_1903,N_1695,N_1745);
or U1904 (N_1904,N_1795,N_1741);
or U1905 (N_1905,N_1778,N_1766);
nor U1906 (N_1906,N_1684,N_1780);
xnor U1907 (N_1907,N_1741,N_1764);
or U1908 (N_1908,N_1620,N_1754);
and U1909 (N_1909,N_1776,N_1681);
or U1910 (N_1910,N_1712,N_1782);
and U1911 (N_1911,N_1702,N_1664);
or U1912 (N_1912,N_1720,N_1615);
nand U1913 (N_1913,N_1647,N_1672);
nor U1914 (N_1914,N_1768,N_1796);
or U1915 (N_1915,N_1691,N_1659);
nor U1916 (N_1916,N_1790,N_1710);
or U1917 (N_1917,N_1729,N_1778);
nor U1918 (N_1918,N_1698,N_1743);
or U1919 (N_1919,N_1774,N_1612);
xor U1920 (N_1920,N_1615,N_1694);
xnor U1921 (N_1921,N_1780,N_1706);
nor U1922 (N_1922,N_1773,N_1728);
nand U1923 (N_1923,N_1671,N_1612);
nor U1924 (N_1924,N_1671,N_1644);
nor U1925 (N_1925,N_1774,N_1627);
nand U1926 (N_1926,N_1771,N_1689);
nor U1927 (N_1927,N_1711,N_1643);
or U1928 (N_1928,N_1672,N_1797);
nor U1929 (N_1929,N_1749,N_1610);
or U1930 (N_1930,N_1721,N_1769);
nand U1931 (N_1931,N_1752,N_1783);
nand U1932 (N_1932,N_1660,N_1785);
nor U1933 (N_1933,N_1628,N_1699);
xnor U1934 (N_1934,N_1689,N_1616);
or U1935 (N_1935,N_1643,N_1652);
and U1936 (N_1936,N_1612,N_1698);
or U1937 (N_1937,N_1689,N_1785);
and U1938 (N_1938,N_1743,N_1709);
nor U1939 (N_1939,N_1628,N_1614);
nor U1940 (N_1940,N_1748,N_1628);
and U1941 (N_1941,N_1750,N_1790);
nand U1942 (N_1942,N_1750,N_1782);
or U1943 (N_1943,N_1755,N_1712);
nor U1944 (N_1944,N_1766,N_1722);
or U1945 (N_1945,N_1668,N_1608);
xnor U1946 (N_1946,N_1696,N_1796);
nand U1947 (N_1947,N_1785,N_1633);
and U1948 (N_1948,N_1782,N_1739);
nor U1949 (N_1949,N_1739,N_1624);
xor U1950 (N_1950,N_1718,N_1704);
and U1951 (N_1951,N_1617,N_1706);
and U1952 (N_1952,N_1751,N_1641);
or U1953 (N_1953,N_1700,N_1755);
nand U1954 (N_1954,N_1764,N_1621);
nand U1955 (N_1955,N_1612,N_1609);
nor U1956 (N_1956,N_1756,N_1654);
nor U1957 (N_1957,N_1628,N_1752);
nand U1958 (N_1958,N_1733,N_1639);
or U1959 (N_1959,N_1690,N_1616);
nor U1960 (N_1960,N_1729,N_1637);
or U1961 (N_1961,N_1607,N_1738);
nor U1962 (N_1962,N_1657,N_1620);
xor U1963 (N_1963,N_1608,N_1720);
and U1964 (N_1964,N_1759,N_1704);
and U1965 (N_1965,N_1734,N_1639);
nor U1966 (N_1966,N_1626,N_1745);
nand U1967 (N_1967,N_1663,N_1726);
xnor U1968 (N_1968,N_1782,N_1603);
nand U1969 (N_1969,N_1718,N_1610);
xnor U1970 (N_1970,N_1602,N_1752);
nand U1971 (N_1971,N_1745,N_1601);
or U1972 (N_1972,N_1795,N_1793);
nand U1973 (N_1973,N_1605,N_1799);
and U1974 (N_1974,N_1612,N_1633);
nor U1975 (N_1975,N_1721,N_1653);
nor U1976 (N_1976,N_1708,N_1744);
or U1977 (N_1977,N_1720,N_1672);
or U1978 (N_1978,N_1793,N_1654);
nand U1979 (N_1979,N_1789,N_1640);
nand U1980 (N_1980,N_1797,N_1692);
nand U1981 (N_1981,N_1666,N_1604);
xor U1982 (N_1982,N_1744,N_1612);
or U1983 (N_1983,N_1751,N_1709);
xor U1984 (N_1984,N_1601,N_1650);
nor U1985 (N_1985,N_1672,N_1605);
nand U1986 (N_1986,N_1777,N_1726);
or U1987 (N_1987,N_1709,N_1726);
nor U1988 (N_1988,N_1733,N_1782);
and U1989 (N_1989,N_1703,N_1651);
nor U1990 (N_1990,N_1640,N_1665);
nor U1991 (N_1991,N_1615,N_1737);
nor U1992 (N_1992,N_1600,N_1797);
nor U1993 (N_1993,N_1672,N_1794);
nor U1994 (N_1994,N_1757,N_1754);
nand U1995 (N_1995,N_1743,N_1722);
or U1996 (N_1996,N_1655,N_1724);
nor U1997 (N_1997,N_1631,N_1707);
nor U1998 (N_1998,N_1763,N_1624);
nand U1999 (N_1999,N_1681,N_1791);
nand U2000 (N_2000,N_1887,N_1875);
nor U2001 (N_2001,N_1939,N_1929);
nand U2002 (N_2002,N_1995,N_1973);
and U2003 (N_2003,N_1994,N_1872);
and U2004 (N_2004,N_1970,N_1867);
nand U2005 (N_2005,N_1981,N_1873);
and U2006 (N_2006,N_1903,N_1848);
or U2007 (N_2007,N_1951,N_1891);
xnor U2008 (N_2008,N_1888,N_1952);
or U2009 (N_2009,N_1895,N_1866);
and U2010 (N_2010,N_1874,N_1963);
or U2011 (N_2011,N_1828,N_1832);
or U2012 (N_2012,N_1945,N_1960);
or U2013 (N_2013,N_1871,N_1842);
xnor U2014 (N_2014,N_1984,N_1800);
or U2015 (N_2015,N_1819,N_1980);
and U2016 (N_2016,N_1930,N_1912);
xnor U2017 (N_2017,N_1997,N_1851);
xnor U2018 (N_2018,N_1830,N_1834);
nand U2019 (N_2019,N_1835,N_1999);
nor U2020 (N_2020,N_1885,N_1838);
nand U2021 (N_2021,N_1869,N_1979);
and U2022 (N_2022,N_1890,N_1804);
or U2023 (N_2023,N_1964,N_1863);
xor U2024 (N_2024,N_1827,N_1913);
nand U2025 (N_2025,N_1884,N_1957);
and U2026 (N_2026,N_1801,N_1852);
and U2027 (N_2027,N_1990,N_1946);
nor U2028 (N_2028,N_1932,N_1879);
and U2029 (N_2029,N_1868,N_1841);
nand U2030 (N_2030,N_1976,N_1893);
nor U2031 (N_2031,N_1808,N_1958);
or U2032 (N_2032,N_1983,N_1914);
or U2033 (N_2033,N_1961,N_1996);
xor U2034 (N_2034,N_1829,N_1940);
or U2035 (N_2035,N_1949,N_1825);
nand U2036 (N_2036,N_1998,N_1818);
and U2037 (N_2037,N_1921,N_1947);
xor U2038 (N_2038,N_1991,N_1924);
or U2039 (N_2039,N_1836,N_1977);
or U2040 (N_2040,N_1942,N_1986);
nor U2041 (N_2041,N_1959,N_1982);
or U2042 (N_2042,N_1896,N_1978);
or U2043 (N_2043,N_1811,N_1824);
and U2044 (N_2044,N_1908,N_1925);
or U2045 (N_2045,N_1826,N_1815);
nand U2046 (N_2046,N_1870,N_1931);
or U2047 (N_2047,N_1894,N_1943);
nand U2048 (N_2048,N_1992,N_1915);
nor U2049 (N_2049,N_1857,N_1989);
nor U2050 (N_2050,N_1966,N_1855);
and U2051 (N_2051,N_1840,N_1858);
nor U2052 (N_2052,N_1916,N_1993);
or U2053 (N_2053,N_1864,N_1882);
nand U2054 (N_2054,N_1962,N_1955);
nand U2055 (N_2055,N_1910,N_1805);
or U2056 (N_2056,N_1941,N_1967);
xnor U2057 (N_2057,N_1822,N_1904);
or U2058 (N_2058,N_1944,N_1837);
nor U2059 (N_2059,N_1909,N_1933);
and U2060 (N_2060,N_1965,N_1859);
or U2061 (N_2061,N_1860,N_1985);
or U2062 (N_2062,N_1820,N_1865);
or U2063 (N_2063,N_1843,N_1856);
or U2064 (N_2064,N_1936,N_1806);
nand U2065 (N_2065,N_1972,N_1813);
nor U2066 (N_2066,N_1954,N_1937);
nand U2067 (N_2067,N_1802,N_1918);
nor U2068 (N_2068,N_1809,N_1907);
nor U2069 (N_2069,N_1892,N_1934);
nand U2070 (N_2070,N_1917,N_1846);
and U2071 (N_2071,N_1878,N_1817);
or U2072 (N_2072,N_1987,N_1839);
xnor U2073 (N_2073,N_1911,N_1876);
nor U2074 (N_2074,N_1968,N_1900);
or U2075 (N_2075,N_1886,N_1928);
nand U2076 (N_2076,N_1898,N_1812);
or U2077 (N_2077,N_1862,N_1831);
and U2078 (N_2078,N_1877,N_1899);
nand U2079 (N_2079,N_1971,N_1844);
and U2080 (N_2080,N_1927,N_1901);
xnor U2081 (N_2081,N_1902,N_1803);
nand U2082 (N_2082,N_1953,N_1950);
xnor U2083 (N_2083,N_1956,N_1850);
and U2084 (N_2084,N_1923,N_1854);
xnor U2085 (N_2085,N_1922,N_1810);
xor U2086 (N_2086,N_1821,N_1816);
nand U2087 (N_2087,N_1814,N_1906);
xor U2088 (N_2088,N_1948,N_1935);
and U2089 (N_2089,N_1849,N_1883);
xnor U2090 (N_2090,N_1823,N_1853);
xor U2091 (N_2091,N_1920,N_1880);
nor U2092 (N_2092,N_1881,N_1897);
nor U2093 (N_2093,N_1905,N_1969);
nand U2094 (N_2094,N_1926,N_1847);
and U2095 (N_2095,N_1938,N_1974);
nor U2096 (N_2096,N_1861,N_1975);
nand U2097 (N_2097,N_1807,N_1833);
and U2098 (N_2098,N_1845,N_1988);
nor U2099 (N_2099,N_1889,N_1919);
and U2100 (N_2100,N_1918,N_1815);
or U2101 (N_2101,N_1984,N_1856);
or U2102 (N_2102,N_1848,N_1824);
xnor U2103 (N_2103,N_1872,N_1862);
and U2104 (N_2104,N_1879,N_1910);
and U2105 (N_2105,N_1854,N_1955);
xor U2106 (N_2106,N_1965,N_1921);
nand U2107 (N_2107,N_1917,N_1958);
nand U2108 (N_2108,N_1822,N_1971);
or U2109 (N_2109,N_1973,N_1844);
and U2110 (N_2110,N_1801,N_1993);
nand U2111 (N_2111,N_1801,N_1999);
and U2112 (N_2112,N_1825,N_1823);
and U2113 (N_2113,N_1943,N_1952);
and U2114 (N_2114,N_1916,N_1960);
or U2115 (N_2115,N_1859,N_1908);
or U2116 (N_2116,N_1915,N_1962);
nand U2117 (N_2117,N_1828,N_1860);
and U2118 (N_2118,N_1801,N_1844);
nor U2119 (N_2119,N_1935,N_1878);
xor U2120 (N_2120,N_1945,N_1953);
and U2121 (N_2121,N_1860,N_1893);
nor U2122 (N_2122,N_1971,N_1917);
or U2123 (N_2123,N_1859,N_1816);
xnor U2124 (N_2124,N_1816,N_1871);
nand U2125 (N_2125,N_1984,N_1911);
nand U2126 (N_2126,N_1945,N_1814);
nand U2127 (N_2127,N_1874,N_1959);
nand U2128 (N_2128,N_1851,N_1883);
nand U2129 (N_2129,N_1809,N_1967);
nand U2130 (N_2130,N_1888,N_1847);
nor U2131 (N_2131,N_1971,N_1923);
nand U2132 (N_2132,N_1876,N_1980);
xnor U2133 (N_2133,N_1892,N_1894);
nand U2134 (N_2134,N_1865,N_1944);
or U2135 (N_2135,N_1849,N_1985);
and U2136 (N_2136,N_1813,N_1825);
nor U2137 (N_2137,N_1998,N_1969);
nor U2138 (N_2138,N_1922,N_1848);
and U2139 (N_2139,N_1985,N_1991);
nand U2140 (N_2140,N_1942,N_1897);
or U2141 (N_2141,N_1810,N_1817);
nor U2142 (N_2142,N_1928,N_1949);
nor U2143 (N_2143,N_1863,N_1990);
nor U2144 (N_2144,N_1904,N_1999);
nor U2145 (N_2145,N_1849,N_1895);
and U2146 (N_2146,N_1881,N_1812);
nor U2147 (N_2147,N_1973,N_1832);
or U2148 (N_2148,N_1835,N_1853);
nand U2149 (N_2149,N_1894,N_1804);
nand U2150 (N_2150,N_1897,N_1911);
nand U2151 (N_2151,N_1836,N_1832);
nor U2152 (N_2152,N_1904,N_1828);
xnor U2153 (N_2153,N_1930,N_1909);
xor U2154 (N_2154,N_1940,N_1857);
nor U2155 (N_2155,N_1814,N_1887);
nor U2156 (N_2156,N_1932,N_1822);
nor U2157 (N_2157,N_1819,N_1913);
nor U2158 (N_2158,N_1975,N_1958);
and U2159 (N_2159,N_1948,N_1974);
or U2160 (N_2160,N_1942,N_1819);
xnor U2161 (N_2161,N_1802,N_1821);
nor U2162 (N_2162,N_1892,N_1862);
nand U2163 (N_2163,N_1809,N_1915);
and U2164 (N_2164,N_1817,N_1974);
and U2165 (N_2165,N_1919,N_1902);
or U2166 (N_2166,N_1920,N_1849);
nand U2167 (N_2167,N_1868,N_1910);
nand U2168 (N_2168,N_1816,N_1947);
or U2169 (N_2169,N_1840,N_1937);
or U2170 (N_2170,N_1857,N_1965);
nand U2171 (N_2171,N_1934,N_1967);
or U2172 (N_2172,N_1957,N_1805);
nand U2173 (N_2173,N_1813,N_1966);
and U2174 (N_2174,N_1902,N_1888);
nor U2175 (N_2175,N_1863,N_1982);
nand U2176 (N_2176,N_1851,N_1925);
xnor U2177 (N_2177,N_1903,N_1900);
nand U2178 (N_2178,N_1968,N_1923);
nand U2179 (N_2179,N_1841,N_1879);
and U2180 (N_2180,N_1855,N_1937);
nand U2181 (N_2181,N_1814,N_1994);
and U2182 (N_2182,N_1865,N_1972);
and U2183 (N_2183,N_1817,N_1957);
nand U2184 (N_2184,N_1940,N_1968);
nand U2185 (N_2185,N_1996,N_1993);
xnor U2186 (N_2186,N_1968,N_1852);
and U2187 (N_2187,N_1861,N_1984);
or U2188 (N_2188,N_1975,N_1909);
and U2189 (N_2189,N_1918,N_1939);
or U2190 (N_2190,N_1827,N_1997);
or U2191 (N_2191,N_1891,N_1834);
nor U2192 (N_2192,N_1968,N_1975);
and U2193 (N_2193,N_1867,N_1982);
and U2194 (N_2194,N_1838,N_1951);
xnor U2195 (N_2195,N_1828,N_1886);
and U2196 (N_2196,N_1881,N_1805);
or U2197 (N_2197,N_1810,N_1864);
and U2198 (N_2198,N_1890,N_1953);
or U2199 (N_2199,N_1815,N_1887);
nor U2200 (N_2200,N_2020,N_2093);
or U2201 (N_2201,N_2194,N_2089);
nor U2202 (N_2202,N_2003,N_2199);
or U2203 (N_2203,N_2082,N_2061);
nor U2204 (N_2204,N_2044,N_2091);
or U2205 (N_2205,N_2053,N_2198);
nand U2206 (N_2206,N_2103,N_2175);
nor U2207 (N_2207,N_2078,N_2111);
and U2208 (N_2208,N_2121,N_2150);
or U2209 (N_2209,N_2173,N_2149);
nand U2210 (N_2210,N_2163,N_2137);
or U2211 (N_2211,N_2130,N_2188);
or U2212 (N_2212,N_2054,N_2158);
and U2213 (N_2213,N_2098,N_2174);
nand U2214 (N_2214,N_2114,N_2104);
nor U2215 (N_2215,N_2110,N_2051);
nand U2216 (N_2216,N_2063,N_2105);
and U2217 (N_2217,N_2196,N_2142);
nand U2218 (N_2218,N_2145,N_2073);
nand U2219 (N_2219,N_2179,N_2008);
nand U2220 (N_2220,N_2007,N_2019);
and U2221 (N_2221,N_2124,N_2147);
or U2222 (N_2222,N_2046,N_2070);
and U2223 (N_2223,N_2165,N_2167);
and U2224 (N_2224,N_2172,N_2135);
and U2225 (N_2225,N_2009,N_2000);
and U2226 (N_2226,N_2056,N_2021);
or U2227 (N_2227,N_2086,N_2060);
nor U2228 (N_2228,N_2025,N_2031);
nor U2229 (N_2229,N_2189,N_2016);
or U2230 (N_2230,N_2144,N_2151);
nand U2231 (N_2231,N_2195,N_2171);
nor U2232 (N_2232,N_2100,N_2096);
and U2233 (N_2233,N_2115,N_2045);
and U2234 (N_2234,N_2097,N_2048);
or U2235 (N_2235,N_2084,N_2012);
xor U2236 (N_2236,N_2011,N_2052);
xnor U2237 (N_2237,N_2156,N_2160);
nand U2238 (N_2238,N_2029,N_2076);
or U2239 (N_2239,N_2183,N_2162);
xor U2240 (N_2240,N_2108,N_2069);
nor U2241 (N_2241,N_2032,N_2106);
or U2242 (N_2242,N_2143,N_2122);
nand U2243 (N_2243,N_2087,N_2065);
or U2244 (N_2244,N_2184,N_2131);
nand U2245 (N_2245,N_2140,N_2169);
or U2246 (N_2246,N_2191,N_2197);
xor U2247 (N_2247,N_2141,N_2180);
xor U2248 (N_2248,N_2107,N_2154);
and U2249 (N_2249,N_2068,N_2182);
and U2250 (N_2250,N_2112,N_2043);
nand U2251 (N_2251,N_2080,N_2133);
nand U2252 (N_2252,N_2037,N_2039);
xor U2253 (N_2253,N_2134,N_2005);
and U2254 (N_2254,N_2090,N_2139);
nor U2255 (N_2255,N_2146,N_2040);
nor U2256 (N_2256,N_2109,N_2153);
nor U2257 (N_2257,N_2035,N_2117);
and U2258 (N_2258,N_2041,N_2177);
xnor U2259 (N_2259,N_2138,N_2077);
nor U2260 (N_2260,N_2042,N_2120);
nor U2261 (N_2261,N_2058,N_2074);
nor U2262 (N_2262,N_2038,N_2193);
or U2263 (N_2263,N_2001,N_2034);
nand U2264 (N_2264,N_2059,N_2166);
nor U2265 (N_2265,N_2081,N_2102);
nand U2266 (N_2266,N_2088,N_2132);
and U2267 (N_2267,N_2079,N_2192);
nand U2268 (N_2268,N_2187,N_2123);
nor U2269 (N_2269,N_2085,N_2157);
nor U2270 (N_2270,N_2067,N_2075);
nor U2271 (N_2271,N_2047,N_2168);
xor U2272 (N_2272,N_2148,N_2185);
nand U2273 (N_2273,N_2015,N_2101);
nor U2274 (N_2274,N_2186,N_2055);
and U2275 (N_2275,N_2155,N_2064);
nor U2276 (N_2276,N_2125,N_2126);
nand U2277 (N_2277,N_2050,N_2028);
nand U2278 (N_2278,N_2022,N_2002);
nand U2279 (N_2279,N_2099,N_2062);
nand U2280 (N_2280,N_2026,N_2071);
and U2281 (N_2281,N_2004,N_2030);
and U2282 (N_2282,N_2057,N_2159);
and U2283 (N_2283,N_2033,N_2119);
or U2284 (N_2284,N_2095,N_2136);
nor U2285 (N_2285,N_2178,N_2014);
or U2286 (N_2286,N_2164,N_2024);
nand U2287 (N_2287,N_2152,N_2010);
nand U2288 (N_2288,N_2023,N_2094);
nor U2289 (N_2289,N_2036,N_2018);
or U2290 (N_2290,N_2017,N_2113);
xor U2291 (N_2291,N_2181,N_2128);
nand U2292 (N_2292,N_2176,N_2006);
or U2293 (N_2293,N_2170,N_2118);
nor U2294 (N_2294,N_2066,N_2092);
and U2295 (N_2295,N_2013,N_2027);
xnor U2296 (N_2296,N_2190,N_2083);
nand U2297 (N_2297,N_2049,N_2116);
nor U2298 (N_2298,N_2129,N_2161);
or U2299 (N_2299,N_2127,N_2072);
and U2300 (N_2300,N_2101,N_2154);
nor U2301 (N_2301,N_2173,N_2112);
nand U2302 (N_2302,N_2192,N_2038);
nor U2303 (N_2303,N_2165,N_2104);
and U2304 (N_2304,N_2061,N_2032);
nand U2305 (N_2305,N_2144,N_2020);
nand U2306 (N_2306,N_2014,N_2168);
xnor U2307 (N_2307,N_2124,N_2119);
xnor U2308 (N_2308,N_2006,N_2171);
and U2309 (N_2309,N_2070,N_2057);
nand U2310 (N_2310,N_2188,N_2034);
or U2311 (N_2311,N_2048,N_2154);
or U2312 (N_2312,N_2159,N_2143);
or U2313 (N_2313,N_2000,N_2034);
xnor U2314 (N_2314,N_2112,N_2133);
nand U2315 (N_2315,N_2030,N_2128);
nand U2316 (N_2316,N_2198,N_2104);
nor U2317 (N_2317,N_2126,N_2085);
xor U2318 (N_2318,N_2128,N_2148);
and U2319 (N_2319,N_2197,N_2123);
nand U2320 (N_2320,N_2101,N_2006);
xnor U2321 (N_2321,N_2081,N_2163);
nand U2322 (N_2322,N_2050,N_2136);
xor U2323 (N_2323,N_2093,N_2120);
nor U2324 (N_2324,N_2118,N_2157);
or U2325 (N_2325,N_2021,N_2028);
nand U2326 (N_2326,N_2191,N_2148);
nand U2327 (N_2327,N_2014,N_2190);
and U2328 (N_2328,N_2081,N_2170);
or U2329 (N_2329,N_2070,N_2098);
nor U2330 (N_2330,N_2110,N_2038);
nor U2331 (N_2331,N_2046,N_2079);
and U2332 (N_2332,N_2043,N_2151);
or U2333 (N_2333,N_2165,N_2072);
or U2334 (N_2334,N_2015,N_2125);
or U2335 (N_2335,N_2134,N_2073);
xnor U2336 (N_2336,N_2093,N_2107);
or U2337 (N_2337,N_2022,N_2072);
nand U2338 (N_2338,N_2061,N_2011);
nor U2339 (N_2339,N_2050,N_2056);
nor U2340 (N_2340,N_2077,N_2147);
and U2341 (N_2341,N_2049,N_2111);
nor U2342 (N_2342,N_2021,N_2022);
nand U2343 (N_2343,N_2167,N_2112);
nor U2344 (N_2344,N_2059,N_2022);
and U2345 (N_2345,N_2093,N_2114);
or U2346 (N_2346,N_2131,N_2093);
nor U2347 (N_2347,N_2195,N_2035);
and U2348 (N_2348,N_2067,N_2069);
xnor U2349 (N_2349,N_2103,N_2123);
nand U2350 (N_2350,N_2068,N_2145);
nand U2351 (N_2351,N_2121,N_2000);
or U2352 (N_2352,N_2172,N_2021);
nand U2353 (N_2353,N_2065,N_2192);
or U2354 (N_2354,N_2024,N_2084);
nor U2355 (N_2355,N_2042,N_2082);
nand U2356 (N_2356,N_2072,N_2123);
and U2357 (N_2357,N_2075,N_2085);
and U2358 (N_2358,N_2155,N_2077);
and U2359 (N_2359,N_2069,N_2169);
or U2360 (N_2360,N_2016,N_2005);
nor U2361 (N_2361,N_2089,N_2084);
or U2362 (N_2362,N_2042,N_2150);
and U2363 (N_2363,N_2126,N_2137);
xnor U2364 (N_2364,N_2000,N_2048);
xnor U2365 (N_2365,N_2191,N_2020);
nor U2366 (N_2366,N_2166,N_2119);
nor U2367 (N_2367,N_2134,N_2148);
or U2368 (N_2368,N_2185,N_2006);
or U2369 (N_2369,N_2070,N_2026);
nor U2370 (N_2370,N_2082,N_2035);
nor U2371 (N_2371,N_2089,N_2171);
or U2372 (N_2372,N_2125,N_2060);
nor U2373 (N_2373,N_2127,N_2165);
xor U2374 (N_2374,N_2122,N_2107);
nand U2375 (N_2375,N_2198,N_2070);
nor U2376 (N_2376,N_2048,N_2021);
or U2377 (N_2377,N_2069,N_2083);
and U2378 (N_2378,N_2020,N_2186);
or U2379 (N_2379,N_2056,N_2036);
nand U2380 (N_2380,N_2007,N_2065);
nor U2381 (N_2381,N_2032,N_2091);
nand U2382 (N_2382,N_2004,N_2013);
and U2383 (N_2383,N_2003,N_2133);
or U2384 (N_2384,N_2112,N_2098);
and U2385 (N_2385,N_2177,N_2024);
and U2386 (N_2386,N_2193,N_2092);
and U2387 (N_2387,N_2007,N_2027);
or U2388 (N_2388,N_2004,N_2190);
xnor U2389 (N_2389,N_2084,N_2065);
nand U2390 (N_2390,N_2171,N_2096);
and U2391 (N_2391,N_2104,N_2001);
nand U2392 (N_2392,N_2189,N_2197);
nand U2393 (N_2393,N_2183,N_2114);
or U2394 (N_2394,N_2194,N_2063);
nor U2395 (N_2395,N_2006,N_2082);
and U2396 (N_2396,N_2086,N_2108);
and U2397 (N_2397,N_2077,N_2190);
or U2398 (N_2398,N_2122,N_2130);
xnor U2399 (N_2399,N_2076,N_2004);
and U2400 (N_2400,N_2336,N_2237);
and U2401 (N_2401,N_2226,N_2369);
and U2402 (N_2402,N_2345,N_2353);
or U2403 (N_2403,N_2216,N_2257);
nor U2404 (N_2404,N_2269,N_2214);
nor U2405 (N_2405,N_2385,N_2334);
nor U2406 (N_2406,N_2220,N_2333);
nor U2407 (N_2407,N_2258,N_2380);
xor U2408 (N_2408,N_2329,N_2350);
nor U2409 (N_2409,N_2371,N_2358);
nand U2410 (N_2410,N_2359,N_2328);
or U2411 (N_2411,N_2312,N_2344);
or U2412 (N_2412,N_2305,N_2293);
nor U2413 (N_2413,N_2367,N_2215);
nand U2414 (N_2414,N_2292,N_2253);
or U2415 (N_2415,N_2354,N_2375);
or U2416 (N_2416,N_2379,N_2318);
nor U2417 (N_2417,N_2266,N_2223);
nand U2418 (N_2418,N_2327,N_2207);
xor U2419 (N_2419,N_2286,N_2213);
nor U2420 (N_2420,N_2386,N_2326);
nor U2421 (N_2421,N_2346,N_2339);
and U2422 (N_2422,N_2323,N_2316);
and U2423 (N_2423,N_2382,N_2370);
nor U2424 (N_2424,N_2325,N_2303);
nand U2425 (N_2425,N_2310,N_2397);
nand U2426 (N_2426,N_2264,N_2268);
or U2427 (N_2427,N_2224,N_2271);
nor U2428 (N_2428,N_2265,N_2285);
or U2429 (N_2429,N_2281,N_2311);
or U2430 (N_2430,N_2201,N_2372);
nand U2431 (N_2431,N_2277,N_2330);
or U2432 (N_2432,N_2282,N_2300);
or U2433 (N_2433,N_2217,N_2284);
and U2434 (N_2434,N_2396,N_2274);
nor U2435 (N_2435,N_2309,N_2221);
nor U2436 (N_2436,N_2381,N_2234);
nand U2437 (N_2437,N_2383,N_2204);
or U2438 (N_2438,N_2242,N_2315);
nand U2439 (N_2439,N_2211,N_2230);
and U2440 (N_2440,N_2262,N_2395);
or U2441 (N_2441,N_2297,N_2236);
nand U2442 (N_2442,N_2273,N_2392);
or U2443 (N_2443,N_2319,N_2390);
xor U2444 (N_2444,N_2294,N_2260);
and U2445 (N_2445,N_2299,N_2256);
or U2446 (N_2446,N_2366,N_2343);
nor U2447 (N_2447,N_2302,N_2296);
nand U2448 (N_2448,N_2252,N_2384);
or U2449 (N_2449,N_2317,N_2357);
or U2450 (N_2450,N_2363,N_2276);
nor U2451 (N_2451,N_2225,N_2391);
nand U2452 (N_2452,N_2368,N_2244);
or U2453 (N_2453,N_2321,N_2347);
nor U2454 (N_2454,N_2324,N_2241);
and U2455 (N_2455,N_2374,N_2348);
nand U2456 (N_2456,N_2218,N_2340);
nand U2457 (N_2457,N_2275,N_2261);
nand U2458 (N_2458,N_2206,N_2247);
nand U2459 (N_2459,N_2259,N_2356);
or U2460 (N_2460,N_2280,N_2306);
nand U2461 (N_2461,N_2243,N_2362);
and U2462 (N_2462,N_2228,N_2227);
xor U2463 (N_2463,N_2361,N_2222);
nand U2464 (N_2464,N_2210,N_2377);
and U2465 (N_2465,N_2376,N_2394);
nand U2466 (N_2466,N_2245,N_2239);
or U2467 (N_2467,N_2248,N_2202);
nand U2468 (N_2468,N_2322,N_2212);
and U2469 (N_2469,N_2229,N_2263);
xnor U2470 (N_2470,N_2298,N_2205);
and U2471 (N_2471,N_2200,N_2373);
or U2472 (N_2472,N_2314,N_2304);
or U2473 (N_2473,N_2320,N_2278);
and U2474 (N_2474,N_2355,N_2332);
xor U2475 (N_2475,N_2351,N_2335);
nor U2476 (N_2476,N_2233,N_2341);
nor U2477 (N_2477,N_2398,N_2364);
and U2478 (N_2478,N_2308,N_2288);
and U2479 (N_2479,N_2208,N_2389);
nand U2480 (N_2480,N_2255,N_2399);
or U2481 (N_2481,N_2287,N_2240);
nor U2482 (N_2482,N_2290,N_2360);
nand U2483 (N_2483,N_2238,N_2283);
and U2484 (N_2484,N_2279,N_2331);
nor U2485 (N_2485,N_2272,N_2291);
or U2486 (N_2486,N_2235,N_2209);
xor U2487 (N_2487,N_2254,N_2313);
or U2488 (N_2488,N_2289,N_2352);
xnor U2489 (N_2489,N_2203,N_2307);
or U2490 (N_2490,N_2270,N_2337);
nor U2491 (N_2491,N_2378,N_2301);
nand U2492 (N_2492,N_2387,N_2232);
or U2493 (N_2493,N_2231,N_2246);
or U2494 (N_2494,N_2267,N_2249);
and U2495 (N_2495,N_2388,N_2393);
or U2496 (N_2496,N_2342,N_2251);
nor U2497 (N_2497,N_2365,N_2219);
or U2498 (N_2498,N_2250,N_2349);
xor U2499 (N_2499,N_2295,N_2338);
or U2500 (N_2500,N_2334,N_2203);
or U2501 (N_2501,N_2333,N_2338);
nand U2502 (N_2502,N_2258,N_2333);
and U2503 (N_2503,N_2227,N_2201);
or U2504 (N_2504,N_2304,N_2208);
nand U2505 (N_2505,N_2299,N_2279);
and U2506 (N_2506,N_2329,N_2241);
and U2507 (N_2507,N_2398,N_2239);
or U2508 (N_2508,N_2204,N_2396);
or U2509 (N_2509,N_2305,N_2296);
and U2510 (N_2510,N_2231,N_2239);
and U2511 (N_2511,N_2331,N_2327);
nor U2512 (N_2512,N_2232,N_2295);
and U2513 (N_2513,N_2350,N_2261);
nor U2514 (N_2514,N_2383,N_2214);
xor U2515 (N_2515,N_2399,N_2206);
nand U2516 (N_2516,N_2274,N_2321);
nor U2517 (N_2517,N_2331,N_2244);
nand U2518 (N_2518,N_2200,N_2299);
nand U2519 (N_2519,N_2273,N_2378);
xnor U2520 (N_2520,N_2256,N_2335);
nand U2521 (N_2521,N_2228,N_2358);
nand U2522 (N_2522,N_2382,N_2246);
or U2523 (N_2523,N_2272,N_2306);
or U2524 (N_2524,N_2349,N_2275);
nand U2525 (N_2525,N_2215,N_2376);
xnor U2526 (N_2526,N_2243,N_2277);
xnor U2527 (N_2527,N_2351,N_2309);
and U2528 (N_2528,N_2382,N_2210);
nor U2529 (N_2529,N_2278,N_2312);
and U2530 (N_2530,N_2335,N_2392);
or U2531 (N_2531,N_2302,N_2214);
or U2532 (N_2532,N_2357,N_2385);
or U2533 (N_2533,N_2267,N_2330);
and U2534 (N_2534,N_2344,N_2328);
nor U2535 (N_2535,N_2375,N_2246);
nor U2536 (N_2536,N_2278,N_2277);
or U2537 (N_2537,N_2206,N_2394);
and U2538 (N_2538,N_2300,N_2244);
or U2539 (N_2539,N_2249,N_2228);
nand U2540 (N_2540,N_2318,N_2286);
xnor U2541 (N_2541,N_2255,N_2396);
nand U2542 (N_2542,N_2215,N_2211);
nand U2543 (N_2543,N_2215,N_2365);
and U2544 (N_2544,N_2205,N_2270);
xnor U2545 (N_2545,N_2391,N_2263);
nand U2546 (N_2546,N_2307,N_2257);
xnor U2547 (N_2547,N_2363,N_2299);
and U2548 (N_2548,N_2268,N_2313);
and U2549 (N_2549,N_2245,N_2318);
xnor U2550 (N_2550,N_2366,N_2242);
and U2551 (N_2551,N_2306,N_2323);
nand U2552 (N_2552,N_2258,N_2362);
or U2553 (N_2553,N_2240,N_2228);
nand U2554 (N_2554,N_2339,N_2229);
nor U2555 (N_2555,N_2379,N_2359);
nor U2556 (N_2556,N_2222,N_2238);
or U2557 (N_2557,N_2350,N_2394);
or U2558 (N_2558,N_2345,N_2332);
or U2559 (N_2559,N_2223,N_2345);
and U2560 (N_2560,N_2359,N_2395);
xnor U2561 (N_2561,N_2258,N_2391);
nand U2562 (N_2562,N_2296,N_2345);
nor U2563 (N_2563,N_2381,N_2393);
and U2564 (N_2564,N_2301,N_2217);
nor U2565 (N_2565,N_2305,N_2229);
or U2566 (N_2566,N_2336,N_2270);
nor U2567 (N_2567,N_2311,N_2278);
nor U2568 (N_2568,N_2368,N_2261);
nand U2569 (N_2569,N_2266,N_2301);
or U2570 (N_2570,N_2297,N_2273);
nor U2571 (N_2571,N_2227,N_2316);
nand U2572 (N_2572,N_2223,N_2307);
and U2573 (N_2573,N_2238,N_2385);
nor U2574 (N_2574,N_2388,N_2353);
nor U2575 (N_2575,N_2326,N_2268);
nor U2576 (N_2576,N_2375,N_2341);
nor U2577 (N_2577,N_2237,N_2305);
xnor U2578 (N_2578,N_2298,N_2289);
and U2579 (N_2579,N_2265,N_2391);
xor U2580 (N_2580,N_2350,N_2241);
nor U2581 (N_2581,N_2385,N_2292);
nor U2582 (N_2582,N_2361,N_2237);
nand U2583 (N_2583,N_2237,N_2232);
or U2584 (N_2584,N_2240,N_2229);
nor U2585 (N_2585,N_2399,N_2353);
nand U2586 (N_2586,N_2224,N_2329);
or U2587 (N_2587,N_2225,N_2355);
nor U2588 (N_2588,N_2388,N_2227);
or U2589 (N_2589,N_2326,N_2258);
nand U2590 (N_2590,N_2285,N_2217);
and U2591 (N_2591,N_2258,N_2389);
nand U2592 (N_2592,N_2351,N_2391);
nor U2593 (N_2593,N_2238,N_2227);
and U2594 (N_2594,N_2351,N_2206);
nand U2595 (N_2595,N_2283,N_2398);
nor U2596 (N_2596,N_2267,N_2357);
nor U2597 (N_2597,N_2260,N_2243);
xnor U2598 (N_2598,N_2371,N_2246);
or U2599 (N_2599,N_2236,N_2379);
and U2600 (N_2600,N_2481,N_2419);
nand U2601 (N_2601,N_2503,N_2477);
nor U2602 (N_2602,N_2573,N_2489);
nand U2603 (N_2603,N_2455,N_2548);
nor U2604 (N_2604,N_2545,N_2567);
nor U2605 (N_2605,N_2591,N_2575);
nor U2606 (N_2606,N_2407,N_2518);
or U2607 (N_2607,N_2589,N_2426);
nand U2608 (N_2608,N_2541,N_2499);
nor U2609 (N_2609,N_2469,N_2462);
xnor U2610 (N_2610,N_2590,N_2552);
nand U2611 (N_2611,N_2453,N_2409);
and U2612 (N_2612,N_2470,N_2562);
and U2613 (N_2613,N_2584,N_2547);
nor U2614 (N_2614,N_2558,N_2523);
nand U2615 (N_2615,N_2557,N_2555);
nor U2616 (N_2616,N_2417,N_2411);
or U2617 (N_2617,N_2597,N_2526);
or U2618 (N_2618,N_2519,N_2479);
nor U2619 (N_2619,N_2485,N_2450);
nand U2620 (N_2620,N_2429,N_2421);
nand U2621 (N_2621,N_2566,N_2515);
and U2622 (N_2622,N_2480,N_2451);
and U2623 (N_2623,N_2415,N_2520);
nand U2624 (N_2624,N_2529,N_2482);
nor U2625 (N_2625,N_2452,N_2550);
xnor U2626 (N_2626,N_2507,N_2554);
nor U2627 (N_2627,N_2546,N_2588);
or U2628 (N_2628,N_2471,N_2516);
or U2629 (N_2629,N_2410,N_2561);
xor U2630 (N_2630,N_2449,N_2468);
and U2631 (N_2631,N_2543,N_2528);
or U2632 (N_2632,N_2506,N_2565);
or U2633 (N_2633,N_2512,N_2495);
or U2634 (N_2634,N_2427,N_2522);
nand U2635 (N_2635,N_2420,N_2563);
xor U2636 (N_2636,N_2438,N_2599);
and U2637 (N_2637,N_2444,N_2542);
or U2638 (N_2638,N_2502,N_2556);
xor U2639 (N_2639,N_2577,N_2459);
nand U2640 (N_2640,N_2536,N_2490);
xor U2641 (N_2641,N_2423,N_2574);
or U2642 (N_2642,N_2447,N_2576);
nand U2643 (N_2643,N_2464,N_2486);
nand U2644 (N_2644,N_2494,N_2434);
nand U2645 (N_2645,N_2416,N_2592);
nand U2646 (N_2646,N_2514,N_2572);
and U2647 (N_2647,N_2484,N_2463);
nand U2648 (N_2648,N_2433,N_2568);
or U2649 (N_2649,N_2504,N_2517);
nor U2650 (N_2650,N_2532,N_2578);
and U2651 (N_2651,N_2446,N_2585);
and U2652 (N_2652,N_2445,N_2488);
nand U2653 (N_2653,N_2587,N_2594);
nand U2654 (N_2654,N_2475,N_2413);
nand U2655 (N_2655,N_2403,N_2460);
xnor U2656 (N_2656,N_2465,N_2593);
and U2657 (N_2657,N_2513,N_2598);
nand U2658 (N_2658,N_2527,N_2540);
nand U2659 (N_2659,N_2424,N_2472);
nand U2660 (N_2660,N_2509,N_2406);
and U2661 (N_2661,N_2442,N_2571);
nor U2662 (N_2662,N_2483,N_2428);
xnor U2663 (N_2663,N_2511,N_2430);
nor U2664 (N_2664,N_2414,N_2505);
or U2665 (N_2665,N_2501,N_2461);
xor U2666 (N_2666,N_2440,N_2498);
or U2667 (N_2667,N_2425,N_2458);
xor U2668 (N_2668,N_2492,N_2454);
nor U2669 (N_2669,N_2466,N_2583);
and U2670 (N_2670,N_2443,N_2435);
nand U2671 (N_2671,N_2569,N_2500);
nand U2672 (N_2672,N_2595,N_2570);
or U2673 (N_2673,N_2437,N_2582);
nand U2674 (N_2674,N_2580,N_2412);
nand U2675 (N_2675,N_2478,N_2400);
nand U2676 (N_2676,N_2448,N_2524);
nor U2677 (N_2677,N_2497,N_2467);
xor U2678 (N_2678,N_2560,N_2534);
or U2679 (N_2679,N_2544,N_2586);
or U2680 (N_2680,N_2539,N_2422);
or U2681 (N_2681,N_2456,N_2537);
and U2682 (N_2682,N_2418,N_2564);
or U2683 (N_2683,N_2510,N_2432);
and U2684 (N_2684,N_2493,N_2538);
xnor U2685 (N_2685,N_2533,N_2405);
nand U2686 (N_2686,N_2436,N_2551);
or U2687 (N_2687,N_2439,N_2579);
xor U2688 (N_2688,N_2401,N_2525);
nor U2689 (N_2689,N_2402,N_2408);
nor U2690 (N_2690,N_2431,N_2559);
nand U2691 (N_2691,N_2553,N_2530);
or U2692 (N_2692,N_2476,N_2531);
nand U2693 (N_2693,N_2535,N_2496);
or U2694 (N_2694,N_2581,N_2491);
or U2695 (N_2695,N_2457,N_2596);
nor U2696 (N_2696,N_2474,N_2549);
nand U2697 (N_2697,N_2508,N_2473);
or U2698 (N_2698,N_2404,N_2521);
nand U2699 (N_2699,N_2441,N_2487);
xnor U2700 (N_2700,N_2579,N_2566);
nand U2701 (N_2701,N_2445,N_2515);
nand U2702 (N_2702,N_2559,N_2585);
or U2703 (N_2703,N_2537,N_2449);
nor U2704 (N_2704,N_2500,N_2596);
nor U2705 (N_2705,N_2589,N_2487);
nor U2706 (N_2706,N_2432,N_2430);
and U2707 (N_2707,N_2557,N_2544);
nor U2708 (N_2708,N_2489,N_2528);
and U2709 (N_2709,N_2518,N_2552);
nor U2710 (N_2710,N_2472,N_2576);
xnor U2711 (N_2711,N_2527,N_2562);
nor U2712 (N_2712,N_2519,N_2571);
nand U2713 (N_2713,N_2585,N_2588);
xnor U2714 (N_2714,N_2571,N_2523);
or U2715 (N_2715,N_2410,N_2594);
nor U2716 (N_2716,N_2476,N_2406);
nand U2717 (N_2717,N_2594,N_2590);
nand U2718 (N_2718,N_2430,N_2472);
and U2719 (N_2719,N_2552,N_2546);
and U2720 (N_2720,N_2413,N_2441);
nand U2721 (N_2721,N_2533,N_2489);
or U2722 (N_2722,N_2439,N_2549);
and U2723 (N_2723,N_2402,N_2496);
and U2724 (N_2724,N_2539,N_2557);
nand U2725 (N_2725,N_2587,N_2493);
xnor U2726 (N_2726,N_2423,N_2447);
and U2727 (N_2727,N_2484,N_2506);
xnor U2728 (N_2728,N_2514,N_2519);
and U2729 (N_2729,N_2540,N_2409);
or U2730 (N_2730,N_2581,N_2488);
xnor U2731 (N_2731,N_2417,N_2408);
or U2732 (N_2732,N_2587,N_2546);
xnor U2733 (N_2733,N_2526,N_2537);
or U2734 (N_2734,N_2442,N_2546);
nand U2735 (N_2735,N_2426,N_2510);
nand U2736 (N_2736,N_2436,N_2410);
xnor U2737 (N_2737,N_2595,N_2493);
and U2738 (N_2738,N_2567,N_2460);
nor U2739 (N_2739,N_2416,N_2599);
or U2740 (N_2740,N_2480,N_2417);
nand U2741 (N_2741,N_2572,N_2478);
or U2742 (N_2742,N_2503,N_2565);
xor U2743 (N_2743,N_2414,N_2575);
and U2744 (N_2744,N_2460,N_2401);
and U2745 (N_2745,N_2545,N_2473);
nor U2746 (N_2746,N_2486,N_2465);
nor U2747 (N_2747,N_2534,N_2433);
xor U2748 (N_2748,N_2493,N_2422);
nand U2749 (N_2749,N_2476,N_2485);
or U2750 (N_2750,N_2460,N_2542);
and U2751 (N_2751,N_2465,N_2508);
nand U2752 (N_2752,N_2457,N_2498);
and U2753 (N_2753,N_2505,N_2485);
or U2754 (N_2754,N_2483,N_2449);
and U2755 (N_2755,N_2542,N_2493);
xor U2756 (N_2756,N_2479,N_2426);
xnor U2757 (N_2757,N_2435,N_2472);
xor U2758 (N_2758,N_2464,N_2455);
xnor U2759 (N_2759,N_2578,N_2573);
nand U2760 (N_2760,N_2477,N_2556);
and U2761 (N_2761,N_2458,N_2403);
xnor U2762 (N_2762,N_2490,N_2409);
and U2763 (N_2763,N_2497,N_2530);
nand U2764 (N_2764,N_2588,N_2523);
nor U2765 (N_2765,N_2464,N_2536);
and U2766 (N_2766,N_2559,N_2446);
and U2767 (N_2767,N_2453,N_2437);
nor U2768 (N_2768,N_2575,N_2584);
and U2769 (N_2769,N_2567,N_2451);
or U2770 (N_2770,N_2442,N_2537);
nand U2771 (N_2771,N_2452,N_2485);
and U2772 (N_2772,N_2495,N_2463);
nand U2773 (N_2773,N_2503,N_2547);
and U2774 (N_2774,N_2430,N_2479);
nand U2775 (N_2775,N_2585,N_2495);
nor U2776 (N_2776,N_2548,N_2521);
nand U2777 (N_2777,N_2581,N_2453);
xor U2778 (N_2778,N_2592,N_2561);
and U2779 (N_2779,N_2575,N_2598);
and U2780 (N_2780,N_2542,N_2525);
and U2781 (N_2781,N_2567,N_2598);
nand U2782 (N_2782,N_2456,N_2533);
or U2783 (N_2783,N_2472,N_2491);
and U2784 (N_2784,N_2465,N_2529);
nor U2785 (N_2785,N_2598,N_2579);
and U2786 (N_2786,N_2583,N_2588);
or U2787 (N_2787,N_2467,N_2473);
xnor U2788 (N_2788,N_2594,N_2588);
nand U2789 (N_2789,N_2485,N_2546);
or U2790 (N_2790,N_2422,N_2405);
nor U2791 (N_2791,N_2475,N_2429);
nor U2792 (N_2792,N_2573,N_2445);
nand U2793 (N_2793,N_2422,N_2515);
and U2794 (N_2794,N_2468,N_2460);
or U2795 (N_2795,N_2592,N_2454);
or U2796 (N_2796,N_2575,N_2490);
nand U2797 (N_2797,N_2400,N_2482);
or U2798 (N_2798,N_2405,N_2576);
nand U2799 (N_2799,N_2489,N_2483);
nor U2800 (N_2800,N_2770,N_2786);
and U2801 (N_2801,N_2642,N_2635);
or U2802 (N_2802,N_2617,N_2760);
nand U2803 (N_2803,N_2781,N_2679);
xor U2804 (N_2804,N_2676,N_2647);
nor U2805 (N_2805,N_2717,N_2790);
and U2806 (N_2806,N_2791,N_2604);
nand U2807 (N_2807,N_2723,N_2733);
nor U2808 (N_2808,N_2780,N_2784);
nand U2809 (N_2809,N_2616,N_2605);
and U2810 (N_2810,N_2757,N_2670);
nand U2811 (N_2811,N_2662,N_2600);
and U2812 (N_2812,N_2799,N_2615);
nor U2813 (N_2813,N_2603,N_2744);
nor U2814 (N_2814,N_2658,N_2764);
and U2815 (N_2815,N_2612,N_2697);
nor U2816 (N_2816,N_2671,N_2722);
nand U2817 (N_2817,N_2798,N_2636);
nand U2818 (N_2818,N_2724,N_2705);
xnor U2819 (N_2819,N_2735,N_2629);
or U2820 (N_2820,N_2749,N_2729);
or U2821 (N_2821,N_2755,N_2690);
and U2822 (N_2822,N_2795,N_2742);
nor U2823 (N_2823,N_2644,N_2631);
nand U2824 (N_2824,N_2687,N_2683);
nand U2825 (N_2825,N_2708,N_2653);
nor U2826 (N_2826,N_2718,N_2634);
and U2827 (N_2827,N_2787,N_2660);
nor U2828 (N_2828,N_2638,N_2637);
nor U2829 (N_2829,N_2624,N_2639);
nor U2830 (N_2830,N_2652,N_2665);
or U2831 (N_2831,N_2689,N_2711);
nor U2832 (N_2832,N_2661,N_2753);
nor U2833 (N_2833,N_2677,N_2756);
nor U2834 (N_2834,N_2626,N_2720);
or U2835 (N_2835,N_2649,N_2684);
and U2836 (N_2836,N_2759,N_2772);
nor U2837 (N_2837,N_2748,N_2669);
and U2838 (N_2838,N_2686,N_2719);
and U2839 (N_2839,N_2736,N_2695);
and U2840 (N_2840,N_2758,N_2655);
and U2841 (N_2841,N_2610,N_2675);
nand U2842 (N_2842,N_2743,N_2674);
nand U2843 (N_2843,N_2651,N_2673);
or U2844 (N_2844,N_2630,N_2727);
or U2845 (N_2845,N_2663,N_2707);
and U2846 (N_2846,N_2704,N_2712);
nand U2847 (N_2847,N_2678,N_2775);
and U2848 (N_2848,N_2646,N_2782);
xnor U2849 (N_2849,N_2609,N_2715);
nor U2850 (N_2850,N_2633,N_2613);
or U2851 (N_2851,N_2607,N_2606);
nand U2852 (N_2852,N_2783,N_2696);
nand U2853 (N_2853,N_2767,N_2738);
nand U2854 (N_2854,N_2728,N_2702);
nor U2855 (N_2855,N_2645,N_2721);
nand U2856 (N_2856,N_2648,N_2625);
or U2857 (N_2857,N_2794,N_2732);
and U2858 (N_2858,N_2619,N_2608);
nor U2859 (N_2859,N_2699,N_2725);
or U2860 (N_2860,N_2771,N_2627);
nor U2861 (N_2861,N_2730,N_2685);
or U2862 (N_2862,N_2698,N_2643);
or U2863 (N_2863,N_2710,N_2703);
and U2864 (N_2864,N_2693,N_2793);
and U2865 (N_2865,N_2611,N_2650);
xor U2866 (N_2866,N_2691,N_2734);
nand U2867 (N_2867,N_2682,N_2632);
xor U2868 (N_2868,N_2763,N_2785);
nor U2869 (N_2869,N_2623,N_2754);
and U2870 (N_2870,N_2680,N_2614);
or U2871 (N_2871,N_2766,N_2694);
and U2872 (N_2872,N_2773,N_2737);
xor U2873 (N_2873,N_2672,N_2765);
or U2874 (N_2874,N_2774,N_2796);
nand U2875 (N_2875,N_2731,N_2777);
and U2876 (N_2876,N_2792,N_2640);
nor U2877 (N_2877,N_2797,N_2701);
xor U2878 (N_2878,N_2745,N_2769);
nand U2879 (N_2879,N_2641,N_2788);
nor U2880 (N_2880,N_2681,N_2618);
xnor U2881 (N_2881,N_2700,N_2620);
or U2882 (N_2882,N_2746,N_2706);
and U2883 (N_2883,N_2622,N_2741);
or U2884 (N_2884,N_2664,N_2601);
nor U2885 (N_2885,N_2776,N_2656);
or U2886 (N_2886,N_2716,N_2750);
nor U2887 (N_2887,N_2714,N_2751);
nor U2888 (N_2888,N_2668,N_2768);
nand U2889 (N_2889,N_2739,N_2688);
and U2890 (N_2890,N_2692,N_2726);
or U2891 (N_2891,N_2778,N_2666);
nor U2892 (N_2892,N_2602,N_2659);
nand U2893 (N_2893,N_2667,N_2628);
nand U2894 (N_2894,N_2709,N_2621);
and U2895 (N_2895,N_2747,N_2761);
and U2896 (N_2896,N_2752,N_2779);
and U2897 (N_2897,N_2657,N_2762);
nor U2898 (N_2898,N_2713,N_2789);
and U2899 (N_2899,N_2740,N_2654);
or U2900 (N_2900,N_2609,N_2677);
nor U2901 (N_2901,N_2650,N_2751);
nand U2902 (N_2902,N_2680,N_2745);
or U2903 (N_2903,N_2711,N_2762);
nor U2904 (N_2904,N_2692,N_2633);
nand U2905 (N_2905,N_2674,N_2765);
nor U2906 (N_2906,N_2712,N_2767);
or U2907 (N_2907,N_2736,N_2648);
xor U2908 (N_2908,N_2793,N_2672);
or U2909 (N_2909,N_2645,N_2726);
nor U2910 (N_2910,N_2711,N_2676);
and U2911 (N_2911,N_2619,N_2628);
nor U2912 (N_2912,N_2729,N_2797);
nand U2913 (N_2913,N_2735,N_2723);
xnor U2914 (N_2914,N_2688,N_2644);
and U2915 (N_2915,N_2752,N_2670);
and U2916 (N_2916,N_2726,N_2653);
or U2917 (N_2917,N_2700,N_2609);
nor U2918 (N_2918,N_2713,N_2752);
and U2919 (N_2919,N_2786,N_2646);
nand U2920 (N_2920,N_2743,N_2681);
or U2921 (N_2921,N_2740,N_2668);
and U2922 (N_2922,N_2629,N_2784);
nor U2923 (N_2923,N_2702,N_2642);
and U2924 (N_2924,N_2663,N_2787);
or U2925 (N_2925,N_2777,N_2798);
nor U2926 (N_2926,N_2735,N_2607);
nor U2927 (N_2927,N_2620,N_2605);
and U2928 (N_2928,N_2683,N_2668);
nor U2929 (N_2929,N_2796,N_2647);
nor U2930 (N_2930,N_2746,N_2683);
and U2931 (N_2931,N_2653,N_2734);
or U2932 (N_2932,N_2752,N_2776);
nor U2933 (N_2933,N_2761,N_2723);
nand U2934 (N_2934,N_2607,N_2670);
or U2935 (N_2935,N_2638,N_2601);
xor U2936 (N_2936,N_2651,N_2796);
and U2937 (N_2937,N_2655,N_2654);
or U2938 (N_2938,N_2602,N_2643);
or U2939 (N_2939,N_2651,N_2707);
or U2940 (N_2940,N_2727,N_2629);
and U2941 (N_2941,N_2718,N_2776);
nor U2942 (N_2942,N_2771,N_2650);
xor U2943 (N_2943,N_2667,N_2768);
nand U2944 (N_2944,N_2720,N_2779);
and U2945 (N_2945,N_2654,N_2644);
and U2946 (N_2946,N_2760,N_2702);
or U2947 (N_2947,N_2604,N_2761);
nand U2948 (N_2948,N_2621,N_2769);
and U2949 (N_2949,N_2684,N_2614);
xnor U2950 (N_2950,N_2768,N_2644);
or U2951 (N_2951,N_2711,N_2655);
and U2952 (N_2952,N_2681,N_2741);
and U2953 (N_2953,N_2645,N_2652);
or U2954 (N_2954,N_2604,N_2679);
nor U2955 (N_2955,N_2762,N_2608);
or U2956 (N_2956,N_2775,N_2652);
nand U2957 (N_2957,N_2713,N_2744);
nand U2958 (N_2958,N_2720,N_2659);
and U2959 (N_2959,N_2778,N_2628);
or U2960 (N_2960,N_2779,N_2638);
nor U2961 (N_2961,N_2666,N_2708);
or U2962 (N_2962,N_2795,N_2649);
nand U2963 (N_2963,N_2636,N_2687);
nand U2964 (N_2964,N_2744,N_2779);
or U2965 (N_2965,N_2604,N_2680);
xnor U2966 (N_2966,N_2736,N_2696);
or U2967 (N_2967,N_2683,N_2711);
and U2968 (N_2968,N_2767,N_2793);
and U2969 (N_2969,N_2601,N_2602);
or U2970 (N_2970,N_2628,N_2662);
nand U2971 (N_2971,N_2787,N_2729);
nand U2972 (N_2972,N_2785,N_2619);
and U2973 (N_2973,N_2612,N_2744);
and U2974 (N_2974,N_2768,N_2745);
nand U2975 (N_2975,N_2724,N_2676);
or U2976 (N_2976,N_2713,N_2648);
nor U2977 (N_2977,N_2729,N_2722);
nor U2978 (N_2978,N_2642,N_2698);
and U2979 (N_2979,N_2796,N_2755);
nand U2980 (N_2980,N_2605,N_2745);
or U2981 (N_2981,N_2661,N_2762);
nor U2982 (N_2982,N_2709,N_2794);
and U2983 (N_2983,N_2707,N_2621);
or U2984 (N_2984,N_2677,N_2671);
nand U2985 (N_2985,N_2752,N_2794);
nor U2986 (N_2986,N_2747,N_2609);
nand U2987 (N_2987,N_2737,N_2609);
nand U2988 (N_2988,N_2712,N_2773);
nand U2989 (N_2989,N_2743,N_2675);
nand U2990 (N_2990,N_2677,N_2797);
nand U2991 (N_2991,N_2744,N_2646);
or U2992 (N_2992,N_2752,N_2631);
and U2993 (N_2993,N_2656,N_2747);
nand U2994 (N_2994,N_2628,N_2717);
nor U2995 (N_2995,N_2691,N_2604);
nor U2996 (N_2996,N_2626,N_2758);
nand U2997 (N_2997,N_2663,N_2743);
and U2998 (N_2998,N_2642,N_2633);
nand U2999 (N_2999,N_2753,N_2600);
and U3000 (N_3000,N_2862,N_2860);
xor U3001 (N_3001,N_2983,N_2923);
xnor U3002 (N_3002,N_2909,N_2900);
nand U3003 (N_3003,N_2999,N_2954);
nor U3004 (N_3004,N_2882,N_2885);
and U3005 (N_3005,N_2963,N_2852);
or U3006 (N_3006,N_2917,N_2830);
and U3007 (N_3007,N_2906,N_2896);
nor U3008 (N_3008,N_2823,N_2971);
xor U3009 (N_3009,N_2807,N_2974);
or U3010 (N_3010,N_2848,N_2969);
or U3011 (N_3011,N_2955,N_2874);
nor U3012 (N_3012,N_2832,N_2812);
nor U3013 (N_3013,N_2944,N_2957);
nor U3014 (N_3014,N_2869,N_2806);
nand U3015 (N_3015,N_2820,N_2819);
xor U3016 (N_3016,N_2849,N_2895);
and U3017 (N_3017,N_2984,N_2972);
nor U3018 (N_3018,N_2910,N_2867);
nor U3019 (N_3019,N_2991,N_2854);
nand U3020 (N_3020,N_2996,N_2843);
nand U3021 (N_3021,N_2824,N_2901);
nor U3022 (N_3022,N_2858,N_2877);
and U3023 (N_3023,N_2836,N_2912);
and U3024 (N_3024,N_2893,N_2907);
or U3025 (N_3025,N_2903,N_2811);
nand U3026 (N_3026,N_2902,N_2987);
and U3027 (N_3027,N_2816,N_2931);
or U3028 (N_3028,N_2829,N_2941);
nor U3029 (N_3029,N_2932,N_2894);
nor U3030 (N_3030,N_2985,N_2865);
nand U3031 (N_3031,N_2962,N_2851);
nand U3032 (N_3032,N_2929,N_2908);
nor U3033 (N_3033,N_2828,N_2964);
nand U3034 (N_3034,N_2891,N_2922);
or U3035 (N_3035,N_2815,N_2868);
xnor U3036 (N_3036,N_2925,N_2943);
and U3037 (N_3037,N_2935,N_2886);
nor U3038 (N_3038,N_2839,N_2937);
or U3039 (N_3039,N_2855,N_2966);
nand U3040 (N_3040,N_2838,N_2995);
or U3041 (N_3041,N_2881,N_2879);
xnor U3042 (N_3042,N_2800,N_2992);
nor U3043 (N_3043,N_2842,N_2953);
and U3044 (N_3044,N_2809,N_2977);
or U3045 (N_3045,N_2890,N_2945);
nand U3046 (N_3046,N_2927,N_2920);
nand U3047 (N_3047,N_2872,N_2870);
or U3048 (N_3048,N_2835,N_2880);
nand U3049 (N_3049,N_2915,N_2837);
xor U3050 (N_3050,N_2919,N_2949);
nor U3051 (N_3051,N_2850,N_2986);
nor U3052 (N_3052,N_2803,N_2804);
or U3053 (N_3053,N_2892,N_2965);
nor U3054 (N_3054,N_2846,N_2875);
nor U3055 (N_3055,N_2834,N_2951);
nor U3056 (N_3056,N_2805,N_2933);
or U3057 (N_3057,N_2960,N_2940);
xnor U3058 (N_3058,N_2831,N_2878);
nor U3059 (N_3059,N_2921,N_2844);
and U3060 (N_3060,N_2801,N_2889);
nand U3061 (N_3061,N_2887,N_2827);
nor U3062 (N_3062,N_2980,N_2866);
nand U3063 (N_3063,N_2864,N_2961);
and U3064 (N_3064,N_2939,N_2973);
nand U3065 (N_3065,N_2993,N_2873);
nor U3066 (N_3066,N_2817,N_2950);
xor U3067 (N_3067,N_2840,N_2863);
or U3068 (N_3068,N_2841,N_2959);
nand U3069 (N_3069,N_2978,N_2818);
and U3070 (N_3070,N_2904,N_2861);
and U3071 (N_3071,N_2926,N_2975);
nand U3072 (N_3072,N_2814,N_2916);
nor U3073 (N_3073,N_2876,N_2967);
nand U3074 (N_3074,N_2897,N_2845);
and U3075 (N_3075,N_2979,N_2952);
nor U3076 (N_3076,N_2822,N_2856);
and U3077 (N_3077,N_2976,N_2913);
nor U3078 (N_3078,N_2898,N_2928);
nor U3079 (N_3079,N_2813,N_2899);
or U3080 (N_3080,N_2934,N_2826);
xor U3081 (N_3081,N_2888,N_2936);
xnor U3082 (N_3082,N_2847,N_2833);
or U3083 (N_3083,N_2989,N_2958);
or U3084 (N_3084,N_2948,N_2911);
nand U3085 (N_3085,N_2853,N_2990);
nor U3086 (N_3086,N_2871,N_2998);
nor U3087 (N_3087,N_2884,N_2988);
nor U3088 (N_3088,N_2968,N_2810);
nand U3089 (N_3089,N_2942,N_2981);
nand U3090 (N_3090,N_2970,N_2956);
or U3091 (N_3091,N_2883,N_2947);
or U3092 (N_3092,N_2930,N_2914);
or U3093 (N_3093,N_2808,N_2821);
and U3094 (N_3094,N_2857,N_2946);
or U3095 (N_3095,N_2994,N_2918);
nand U3096 (N_3096,N_2997,N_2825);
and U3097 (N_3097,N_2982,N_2924);
or U3098 (N_3098,N_2938,N_2905);
nand U3099 (N_3099,N_2802,N_2859);
nand U3100 (N_3100,N_2996,N_2822);
and U3101 (N_3101,N_2999,N_2995);
nor U3102 (N_3102,N_2923,N_2948);
and U3103 (N_3103,N_2864,N_2989);
nor U3104 (N_3104,N_2820,N_2811);
nand U3105 (N_3105,N_2844,N_2813);
and U3106 (N_3106,N_2857,N_2950);
nor U3107 (N_3107,N_2825,N_2836);
or U3108 (N_3108,N_2919,N_2979);
or U3109 (N_3109,N_2915,N_2878);
nor U3110 (N_3110,N_2928,N_2803);
and U3111 (N_3111,N_2883,N_2953);
nand U3112 (N_3112,N_2911,N_2925);
nand U3113 (N_3113,N_2932,N_2865);
nor U3114 (N_3114,N_2916,N_2891);
nand U3115 (N_3115,N_2803,N_2850);
nor U3116 (N_3116,N_2877,N_2919);
nand U3117 (N_3117,N_2973,N_2868);
nor U3118 (N_3118,N_2857,N_2981);
nand U3119 (N_3119,N_2926,N_2810);
nor U3120 (N_3120,N_2847,N_2928);
xor U3121 (N_3121,N_2963,N_2999);
xnor U3122 (N_3122,N_2835,N_2972);
and U3123 (N_3123,N_2838,N_2929);
nor U3124 (N_3124,N_2986,N_2962);
nand U3125 (N_3125,N_2855,N_2987);
and U3126 (N_3126,N_2937,N_2921);
and U3127 (N_3127,N_2826,N_2847);
or U3128 (N_3128,N_2948,N_2855);
and U3129 (N_3129,N_2823,N_2889);
xor U3130 (N_3130,N_2817,N_2852);
nand U3131 (N_3131,N_2985,N_2975);
nor U3132 (N_3132,N_2962,N_2883);
nor U3133 (N_3133,N_2956,N_2843);
or U3134 (N_3134,N_2828,N_2818);
and U3135 (N_3135,N_2924,N_2988);
nor U3136 (N_3136,N_2926,N_2985);
nor U3137 (N_3137,N_2802,N_2929);
nor U3138 (N_3138,N_2903,N_2885);
or U3139 (N_3139,N_2976,N_2920);
xor U3140 (N_3140,N_2858,N_2835);
or U3141 (N_3141,N_2987,N_2890);
and U3142 (N_3142,N_2916,N_2811);
and U3143 (N_3143,N_2959,N_2822);
nand U3144 (N_3144,N_2971,N_2812);
or U3145 (N_3145,N_2821,N_2801);
xnor U3146 (N_3146,N_2842,N_2946);
and U3147 (N_3147,N_2887,N_2834);
xor U3148 (N_3148,N_2952,N_2862);
or U3149 (N_3149,N_2838,N_2905);
or U3150 (N_3150,N_2928,N_2856);
nor U3151 (N_3151,N_2889,N_2993);
xnor U3152 (N_3152,N_2818,N_2940);
and U3153 (N_3153,N_2906,N_2826);
and U3154 (N_3154,N_2994,N_2947);
and U3155 (N_3155,N_2886,N_2892);
and U3156 (N_3156,N_2993,N_2983);
or U3157 (N_3157,N_2901,N_2894);
nand U3158 (N_3158,N_2906,N_2824);
xnor U3159 (N_3159,N_2990,N_2883);
xor U3160 (N_3160,N_2995,N_2925);
and U3161 (N_3161,N_2976,N_2943);
and U3162 (N_3162,N_2839,N_2867);
xnor U3163 (N_3163,N_2800,N_2857);
nor U3164 (N_3164,N_2876,N_2971);
xnor U3165 (N_3165,N_2823,N_2822);
or U3166 (N_3166,N_2940,N_2832);
xnor U3167 (N_3167,N_2893,N_2976);
and U3168 (N_3168,N_2988,N_2875);
nor U3169 (N_3169,N_2844,N_2867);
nor U3170 (N_3170,N_2886,N_2885);
xnor U3171 (N_3171,N_2871,N_2825);
nand U3172 (N_3172,N_2930,N_2881);
and U3173 (N_3173,N_2860,N_2851);
nand U3174 (N_3174,N_2826,N_2890);
xor U3175 (N_3175,N_2967,N_2964);
and U3176 (N_3176,N_2860,N_2870);
nor U3177 (N_3177,N_2831,N_2986);
xor U3178 (N_3178,N_2880,N_2902);
xor U3179 (N_3179,N_2833,N_2944);
xor U3180 (N_3180,N_2925,N_2933);
nand U3181 (N_3181,N_2809,N_2837);
and U3182 (N_3182,N_2849,N_2885);
and U3183 (N_3183,N_2835,N_2818);
xnor U3184 (N_3184,N_2957,N_2874);
or U3185 (N_3185,N_2885,N_2963);
and U3186 (N_3186,N_2975,N_2837);
nand U3187 (N_3187,N_2840,N_2916);
nor U3188 (N_3188,N_2889,N_2894);
nor U3189 (N_3189,N_2816,N_2827);
and U3190 (N_3190,N_2830,N_2805);
or U3191 (N_3191,N_2867,N_2958);
nand U3192 (N_3192,N_2962,N_2823);
nand U3193 (N_3193,N_2982,N_2945);
nand U3194 (N_3194,N_2886,N_2962);
or U3195 (N_3195,N_2872,N_2970);
or U3196 (N_3196,N_2800,N_2833);
or U3197 (N_3197,N_2887,N_2918);
xor U3198 (N_3198,N_2827,N_2926);
and U3199 (N_3199,N_2859,N_2808);
nand U3200 (N_3200,N_3112,N_3048);
or U3201 (N_3201,N_3083,N_3117);
nand U3202 (N_3202,N_3064,N_3143);
nor U3203 (N_3203,N_3169,N_3002);
nand U3204 (N_3204,N_3059,N_3095);
and U3205 (N_3205,N_3029,N_3009);
or U3206 (N_3206,N_3045,N_3137);
nand U3207 (N_3207,N_3135,N_3104);
nand U3208 (N_3208,N_3172,N_3094);
or U3209 (N_3209,N_3134,N_3055);
xor U3210 (N_3210,N_3141,N_3115);
nand U3211 (N_3211,N_3056,N_3182);
nor U3212 (N_3212,N_3046,N_3071);
nand U3213 (N_3213,N_3007,N_3020);
xor U3214 (N_3214,N_3054,N_3139);
nor U3215 (N_3215,N_3121,N_3119);
nor U3216 (N_3216,N_3100,N_3049);
and U3217 (N_3217,N_3197,N_3025);
nor U3218 (N_3218,N_3185,N_3017);
or U3219 (N_3219,N_3107,N_3144);
and U3220 (N_3220,N_3090,N_3158);
nor U3221 (N_3221,N_3075,N_3173);
or U3222 (N_3222,N_3155,N_3034);
nand U3223 (N_3223,N_3022,N_3138);
and U3224 (N_3224,N_3163,N_3146);
or U3225 (N_3225,N_3092,N_3111);
or U3226 (N_3226,N_3194,N_3113);
nand U3227 (N_3227,N_3023,N_3057);
and U3228 (N_3228,N_3188,N_3140);
or U3229 (N_3229,N_3162,N_3067);
nor U3230 (N_3230,N_3050,N_3072);
and U3231 (N_3231,N_3177,N_3198);
nand U3232 (N_3232,N_3103,N_3041);
nand U3233 (N_3233,N_3058,N_3142);
nand U3234 (N_3234,N_3152,N_3091);
nor U3235 (N_3235,N_3108,N_3043);
nand U3236 (N_3236,N_3008,N_3062);
or U3237 (N_3237,N_3042,N_3066);
and U3238 (N_3238,N_3130,N_3039);
or U3239 (N_3239,N_3176,N_3080);
or U3240 (N_3240,N_3124,N_3000);
nand U3241 (N_3241,N_3109,N_3068);
or U3242 (N_3242,N_3166,N_3097);
and U3243 (N_3243,N_3175,N_3086);
nor U3244 (N_3244,N_3148,N_3150);
nand U3245 (N_3245,N_3195,N_3099);
and U3246 (N_3246,N_3074,N_3085);
nor U3247 (N_3247,N_3170,N_3191);
nand U3248 (N_3248,N_3035,N_3005);
and U3249 (N_3249,N_3053,N_3171);
nor U3250 (N_3250,N_3151,N_3164);
and U3251 (N_3251,N_3089,N_3019);
nand U3252 (N_3252,N_3013,N_3178);
or U3253 (N_3253,N_3168,N_3192);
nand U3254 (N_3254,N_3070,N_3156);
nor U3255 (N_3255,N_3021,N_3165);
or U3256 (N_3256,N_3106,N_3014);
xnor U3257 (N_3257,N_3036,N_3160);
nand U3258 (N_3258,N_3101,N_3073);
and U3259 (N_3259,N_3018,N_3174);
and U3260 (N_3260,N_3190,N_3187);
nand U3261 (N_3261,N_3102,N_3105);
and U3262 (N_3262,N_3180,N_3001);
nand U3263 (N_3263,N_3127,N_3044);
or U3264 (N_3264,N_3037,N_3015);
nor U3265 (N_3265,N_3193,N_3145);
nand U3266 (N_3266,N_3031,N_3006);
nand U3267 (N_3267,N_3125,N_3133);
nand U3268 (N_3268,N_3016,N_3051);
xnor U3269 (N_3269,N_3030,N_3012);
and U3270 (N_3270,N_3161,N_3033);
nor U3271 (N_3271,N_3153,N_3154);
and U3272 (N_3272,N_3081,N_3118);
nand U3273 (N_3273,N_3183,N_3069);
or U3274 (N_3274,N_3114,N_3128);
nand U3275 (N_3275,N_3010,N_3026);
or U3276 (N_3276,N_3040,N_3061);
xor U3277 (N_3277,N_3157,N_3186);
and U3278 (N_3278,N_3196,N_3126);
and U3279 (N_3279,N_3129,N_3047);
xor U3280 (N_3280,N_3123,N_3093);
xor U3281 (N_3281,N_3131,N_3110);
or U3282 (N_3282,N_3132,N_3179);
nor U3283 (N_3283,N_3098,N_3159);
nand U3284 (N_3284,N_3003,N_3122);
and U3285 (N_3285,N_3189,N_3065);
nand U3286 (N_3286,N_3060,N_3052);
xnor U3287 (N_3287,N_3079,N_3087);
xor U3288 (N_3288,N_3032,N_3181);
xnor U3289 (N_3289,N_3167,N_3028);
and U3290 (N_3290,N_3096,N_3011);
or U3291 (N_3291,N_3027,N_3004);
nand U3292 (N_3292,N_3120,N_3147);
nand U3293 (N_3293,N_3116,N_3136);
and U3294 (N_3294,N_3038,N_3084);
and U3295 (N_3295,N_3063,N_3024);
and U3296 (N_3296,N_3149,N_3184);
nand U3297 (N_3297,N_3077,N_3078);
nand U3298 (N_3298,N_3088,N_3199);
or U3299 (N_3299,N_3082,N_3076);
or U3300 (N_3300,N_3159,N_3100);
xor U3301 (N_3301,N_3114,N_3013);
nand U3302 (N_3302,N_3101,N_3025);
nor U3303 (N_3303,N_3122,N_3160);
nand U3304 (N_3304,N_3043,N_3048);
and U3305 (N_3305,N_3156,N_3034);
nand U3306 (N_3306,N_3143,N_3060);
and U3307 (N_3307,N_3097,N_3158);
xor U3308 (N_3308,N_3143,N_3022);
and U3309 (N_3309,N_3115,N_3084);
nand U3310 (N_3310,N_3073,N_3090);
nand U3311 (N_3311,N_3037,N_3135);
or U3312 (N_3312,N_3195,N_3118);
xor U3313 (N_3313,N_3089,N_3050);
or U3314 (N_3314,N_3164,N_3161);
nor U3315 (N_3315,N_3188,N_3157);
nor U3316 (N_3316,N_3189,N_3145);
nor U3317 (N_3317,N_3059,N_3180);
nand U3318 (N_3318,N_3069,N_3087);
nor U3319 (N_3319,N_3124,N_3159);
and U3320 (N_3320,N_3191,N_3146);
nor U3321 (N_3321,N_3125,N_3086);
and U3322 (N_3322,N_3087,N_3182);
or U3323 (N_3323,N_3156,N_3172);
and U3324 (N_3324,N_3034,N_3164);
and U3325 (N_3325,N_3077,N_3076);
and U3326 (N_3326,N_3079,N_3020);
and U3327 (N_3327,N_3141,N_3103);
nor U3328 (N_3328,N_3187,N_3152);
and U3329 (N_3329,N_3073,N_3020);
nand U3330 (N_3330,N_3178,N_3147);
and U3331 (N_3331,N_3040,N_3033);
and U3332 (N_3332,N_3166,N_3115);
nor U3333 (N_3333,N_3152,N_3101);
nand U3334 (N_3334,N_3083,N_3100);
nor U3335 (N_3335,N_3059,N_3092);
nand U3336 (N_3336,N_3030,N_3093);
or U3337 (N_3337,N_3045,N_3066);
and U3338 (N_3338,N_3023,N_3010);
or U3339 (N_3339,N_3027,N_3141);
and U3340 (N_3340,N_3120,N_3006);
nand U3341 (N_3341,N_3074,N_3061);
nor U3342 (N_3342,N_3152,N_3136);
or U3343 (N_3343,N_3018,N_3124);
and U3344 (N_3344,N_3159,N_3037);
nor U3345 (N_3345,N_3150,N_3068);
nand U3346 (N_3346,N_3138,N_3158);
nor U3347 (N_3347,N_3192,N_3039);
nor U3348 (N_3348,N_3098,N_3155);
and U3349 (N_3349,N_3071,N_3175);
and U3350 (N_3350,N_3191,N_3140);
nor U3351 (N_3351,N_3199,N_3165);
nand U3352 (N_3352,N_3105,N_3109);
nor U3353 (N_3353,N_3068,N_3137);
nand U3354 (N_3354,N_3058,N_3166);
nor U3355 (N_3355,N_3087,N_3029);
nand U3356 (N_3356,N_3198,N_3131);
or U3357 (N_3357,N_3019,N_3166);
nor U3358 (N_3358,N_3079,N_3003);
or U3359 (N_3359,N_3062,N_3052);
xor U3360 (N_3360,N_3170,N_3067);
and U3361 (N_3361,N_3023,N_3076);
and U3362 (N_3362,N_3007,N_3196);
and U3363 (N_3363,N_3192,N_3032);
xor U3364 (N_3364,N_3137,N_3063);
or U3365 (N_3365,N_3109,N_3027);
nor U3366 (N_3366,N_3079,N_3149);
nor U3367 (N_3367,N_3111,N_3162);
nor U3368 (N_3368,N_3180,N_3002);
nand U3369 (N_3369,N_3074,N_3024);
and U3370 (N_3370,N_3034,N_3072);
or U3371 (N_3371,N_3108,N_3196);
or U3372 (N_3372,N_3148,N_3035);
and U3373 (N_3373,N_3055,N_3065);
or U3374 (N_3374,N_3011,N_3117);
nor U3375 (N_3375,N_3100,N_3171);
nand U3376 (N_3376,N_3135,N_3122);
and U3377 (N_3377,N_3145,N_3185);
or U3378 (N_3378,N_3018,N_3195);
and U3379 (N_3379,N_3140,N_3021);
nor U3380 (N_3380,N_3132,N_3093);
or U3381 (N_3381,N_3010,N_3143);
or U3382 (N_3382,N_3108,N_3140);
or U3383 (N_3383,N_3078,N_3190);
nor U3384 (N_3384,N_3013,N_3091);
nor U3385 (N_3385,N_3021,N_3125);
xnor U3386 (N_3386,N_3145,N_3180);
or U3387 (N_3387,N_3041,N_3024);
nand U3388 (N_3388,N_3020,N_3000);
and U3389 (N_3389,N_3150,N_3049);
nand U3390 (N_3390,N_3005,N_3012);
and U3391 (N_3391,N_3064,N_3070);
or U3392 (N_3392,N_3176,N_3014);
or U3393 (N_3393,N_3130,N_3087);
nor U3394 (N_3394,N_3012,N_3022);
nand U3395 (N_3395,N_3141,N_3032);
or U3396 (N_3396,N_3062,N_3006);
xor U3397 (N_3397,N_3088,N_3005);
or U3398 (N_3398,N_3008,N_3179);
nor U3399 (N_3399,N_3166,N_3066);
nor U3400 (N_3400,N_3323,N_3285);
and U3401 (N_3401,N_3328,N_3232);
and U3402 (N_3402,N_3394,N_3380);
and U3403 (N_3403,N_3200,N_3353);
and U3404 (N_3404,N_3346,N_3365);
and U3405 (N_3405,N_3211,N_3276);
nand U3406 (N_3406,N_3343,N_3220);
or U3407 (N_3407,N_3273,N_3396);
or U3408 (N_3408,N_3361,N_3329);
nor U3409 (N_3409,N_3263,N_3397);
and U3410 (N_3410,N_3334,N_3384);
nor U3411 (N_3411,N_3298,N_3244);
and U3412 (N_3412,N_3216,N_3309);
nor U3413 (N_3413,N_3350,N_3387);
and U3414 (N_3414,N_3360,N_3283);
and U3415 (N_3415,N_3213,N_3234);
and U3416 (N_3416,N_3371,N_3310);
nand U3417 (N_3417,N_3293,N_3383);
xor U3418 (N_3418,N_3331,N_3245);
xnor U3419 (N_3419,N_3214,N_3377);
xor U3420 (N_3420,N_3363,N_3347);
xnor U3421 (N_3421,N_3327,N_3239);
or U3422 (N_3422,N_3289,N_3300);
or U3423 (N_3423,N_3307,N_3274);
nor U3424 (N_3424,N_3357,N_3338);
nand U3425 (N_3425,N_3287,N_3341);
or U3426 (N_3426,N_3279,N_3260);
nand U3427 (N_3427,N_3366,N_3324);
and U3428 (N_3428,N_3246,N_3372);
and U3429 (N_3429,N_3337,N_3325);
or U3430 (N_3430,N_3226,N_3284);
nor U3431 (N_3431,N_3288,N_3208);
nor U3432 (N_3432,N_3336,N_3215);
nor U3433 (N_3433,N_3322,N_3359);
and U3434 (N_3434,N_3332,N_3286);
or U3435 (N_3435,N_3294,N_3306);
and U3436 (N_3436,N_3296,N_3261);
nand U3437 (N_3437,N_3355,N_3352);
or U3438 (N_3438,N_3259,N_3262);
nand U3439 (N_3439,N_3367,N_3302);
nor U3440 (N_3440,N_3277,N_3201);
xor U3441 (N_3441,N_3326,N_3266);
and U3442 (N_3442,N_3392,N_3237);
nand U3443 (N_3443,N_3342,N_3399);
or U3444 (N_3444,N_3206,N_3388);
nor U3445 (N_3445,N_3268,N_3256);
xor U3446 (N_3446,N_3292,N_3319);
nor U3447 (N_3447,N_3345,N_3311);
nand U3448 (N_3448,N_3225,N_3252);
xnor U3449 (N_3449,N_3382,N_3335);
and U3450 (N_3450,N_3398,N_3330);
nand U3451 (N_3451,N_3265,N_3391);
or U3452 (N_3452,N_3351,N_3291);
nand U3453 (N_3453,N_3354,N_3210);
nor U3454 (N_3454,N_3235,N_3203);
nor U3455 (N_3455,N_3258,N_3317);
or U3456 (N_3456,N_3202,N_3281);
nor U3457 (N_3457,N_3305,N_3212);
or U3458 (N_3458,N_3224,N_3381);
nor U3459 (N_3459,N_3340,N_3221);
or U3460 (N_3460,N_3264,N_3242);
nand U3461 (N_3461,N_3315,N_3297);
or U3462 (N_3462,N_3364,N_3217);
nor U3463 (N_3463,N_3385,N_3267);
nor U3464 (N_3464,N_3393,N_3247);
nand U3465 (N_3465,N_3228,N_3278);
nor U3466 (N_3466,N_3241,N_3229);
or U3467 (N_3467,N_3218,N_3379);
nor U3468 (N_3468,N_3270,N_3227);
nand U3469 (N_3469,N_3378,N_3390);
or U3470 (N_3470,N_3250,N_3344);
nor U3471 (N_3471,N_3304,N_3376);
or U3472 (N_3472,N_3230,N_3370);
nor U3473 (N_3473,N_3282,N_3231);
or U3474 (N_3474,N_3362,N_3356);
xnor U3475 (N_3475,N_3312,N_3375);
nor U3476 (N_3476,N_3272,N_3255);
or U3477 (N_3477,N_3358,N_3290);
nor U3478 (N_3478,N_3233,N_3368);
and U3479 (N_3479,N_3318,N_3209);
nand U3480 (N_3480,N_3223,N_3389);
nor U3481 (N_3481,N_3205,N_3219);
nor U3482 (N_3482,N_3249,N_3308);
and U3483 (N_3483,N_3275,N_3374);
xor U3484 (N_3484,N_3240,N_3303);
and U3485 (N_3485,N_3369,N_3280);
xor U3486 (N_3486,N_3386,N_3301);
or U3487 (N_3487,N_3257,N_3299);
nor U3488 (N_3488,N_3236,N_3204);
and U3489 (N_3489,N_3321,N_3316);
nor U3490 (N_3490,N_3395,N_3222);
or U3491 (N_3491,N_3339,N_3295);
nor U3492 (N_3492,N_3320,N_3238);
or U3493 (N_3493,N_3243,N_3254);
or U3494 (N_3494,N_3373,N_3248);
nand U3495 (N_3495,N_3333,N_3251);
and U3496 (N_3496,N_3349,N_3271);
nor U3497 (N_3497,N_3348,N_3314);
xnor U3498 (N_3498,N_3207,N_3313);
nand U3499 (N_3499,N_3253,N_3269);
or U3500 (N_3500,N_3393,N_3310);
and U3501 (N_3501,N_3302,N_3207);
and U3502 (N_3502,N_3278,N_3299);
xor U3503 (N_3503,N_3348,N_3235);
xnor U3504 (N_3504,N_3397,N_3386);
nor U3505 (N_3505,N_3327,N_3249);
nor U3506 (N_3506,N_3352,N_3246);
and U3507 (N_3507,N_3209,N_3267);
and U3508 (N_3508,N_3371,N_3280);
nor U3509 (N_3509,N_3245,N_3344);
nor U3510 (N_3510,N_3205,N_3329);
nor U3511 (N_3511,N_3286,N_3207);
or U3512 (N_3512,N_3274,N_3366);
xor U3513 (N_3513,N_3206,N_3367);
and U3514 (N_3514,N_3267,N_3360);
nor U3515 (N_3515,N_3291,N_3217);
nor U3516 (N_3516,N_3280,N_3253);
xnor U3517 (N_3517,N_3325,N_3251);
nor U3518 (N_3518,N_3365,N_3222);
and U3519 (N_3519,N_3351,N_3320);
and U3520 (N_3520,N_3314,N_3250);
and U3521 (N_3521,N_3391,N_3294);
and U3522 (N_3522,N_3305,N_3283);
and U3523 (N_3523,N_3214,N_3298);
nand U3524 (N_3524,N_3224,N_3211);
and U3525 (N_3525,N_3348,N_3288);
nand U3526 (N_3526,N_3205,N_3328);
nor U3527 (N_3527,N_3372,N_3227);
nor U3528 (N_3528,N_3336,N_3277);
and U3529 (N_3529,N_3294,N_3283);
nor U3530 (N_3530,N_3325,N_3341);
xnor U3531 (N_3531,N_3225,N_3300);
and U3532 (N_3532,N_3204,N_3348);
or U3533 (N_3533,N_3389,N_3243);
xnor U3534 (N_3534,N_3397,N_3293);
or U3535 (N_3535,N_3259,N_3377);
and U3536 (N_3536,N_3208,N_3224);
xnor U3537 (N_3537,N_3331,N_3233);
xor U3538 (N_3538,N_3304,N_3363);
or U3539 (N_3539,N_3247,N_3209);
nand U3540 (N_3540,N_3289,N_3310);
and U3541 (N_3541,N_3274,N_3389);
nand U3542 (N_3542,N_3222,N_3339);
nor U3543 (N_3543,N_3328,N_3297);
xor U3544 (N_3544,N_3348,N_3380);
nand U3545 (N_3545,N_3284,N_3255);
nand U3546 (N_3546,N_3200,N_3220);
nor U3547 (N_3547,N_3398,N_3238);
xor U3548 (N_3548,N_3250,N_3370);
nand U3549 (N_3549,N_3300,N_3381);
and U3550 (N_3550,N_3387,N_3331);
nand U3551 (N_3551,N_3272,N_3240);
or U3552 (N_3552,N_3288,N_3248);
and U3553 (N_3553,N_3319,N_3258);
and U3554 (N_3554,N_3226,N_3318);
or U3555 (N_3555,N_3248,N_3263);
xor U3556 (N_3556,N_3266,N_3275);
nor U3557 (N_3557,N_3317,N_3222);
nor U3558 (N_3558,N_3266,N_3280);
or U3559 (N_3559,N_3259,N_3363);
and U3560 (N_3560,N_3241,N_3285);
nor U3561 (N_3561,N_3303,N_3278);
or U3562 (N_3562,N_3337,N_3310);
or U3563 (N_3563,N_3319,N_3306);
nand U3564 (N_3564,N_3318,N_3240);
or U3565 (N_3565,N_3232,N_3291);
nor U3566 (N_3566,N_3319,N_3342);
nand U3567 (N_3567,N_3267,N_3261);
nor U3568 (N_3568,N_3269,N_3229);
and U3569 (N_3569,N_3271,N_3372);
nand U3570 (N_3570,N_3307,N_3277);
nor U3571 (N_3571,N_3398,N_3307);
or U3572 (N_3572,N_3299,N_3267);
nor U3573 (N_3573,N_3358,N_3252);
nand U3574 (N_3574,N_3264,N_3265);
nor U3575 (N_3575,N_3286,N_3337);
and U3576 (N_3576,N_3305,N_3297);
and U3577 (N_3577,N_3324,N_3294);
or U3578 (N_3578,N_3325,N_3257);
or U3579 (N_3579,N_3226,N_3381);
nor U3580 (N_3580,N_3390,N_3200);
or U3581 (N_3581,N_3347,N_3381);
nand U3582 (N_3582,N_3314,N_3322);
nor U3583 (N_3583,N_3254,N_3270);
nand U3584 (N_3584,N_3313,N_3319);
nor U3585 (N_3585,N_3364,N_3394);
or U3586 (N_3586,N_3396,N_3381);
or U3587 (N_3587,N_3229,N_3202);
or U3588 (N_3588,N_3211,N_3282);
xor U3589 (N_3589,N_3205,N_3256);
xor U3590 (N_3590,N_3302,N_3220);
and U3591 (N_3591,N_3241,N_3364);
nand U3592 (N_3592,N_3313,N_3281);
nand U3593 (N_3593,N_3294,N_3263);
nand U3594 (N_3594,N_3216,N_3208);
nand U3595 (N_3595,N_3313,N_3303);
xnor U3596 (N_3596,N_3242,N_3250);
or U3597 (N_3597,N_3353,N_3226);
nor U3598 (N_3598,N_3382,N_3208);
xor U3599 (N_3599,N_3203,N_3333);
nand U3600 (N_3600,N_3586,N_3411);
nor U3601 (N_3601,N_3524,N_3408);
xor U3602 (N_3602,N_3588,N_3530);
nor U3603 (N_3603,N_3507,N_3457);
nand U3604 (N_3604,N_3535,N_3517);
and U3605 (N_3605,N_3481,N_3403);
nor U3606 (N_3606,N_3594,N_3518);
or U3607 (N_3607,N_3485,N_3545);
nor U3608 (N_3608,N_3423,N_3451);
and U3609 (N_3609,N_3592,N_3565);
or U3610 (N_3610,N_3538,N_3554);
or U3611 (N_3611,N_3448,N_3491);
and U3612 (N_3612,N_3543,N_3424);
or U3613 (N_3613,N_3504,N_3487);
nand U3614 (N_3614,N_3444,N_3443);
or U3615 (N_3615,N_3500,N_3573);
nor U3616 (N_3616,N_3537,N_3480);
and U3617 (N_3617,N_3402,N_3516);
nor U3618 (N_3618,N_3495,N_3497);
or U3619 (N_3619,N_3471,N_3439);
nand U3620 (N_3620,N_3461,N_3540);
nand U3621 (N_3621,N_3434,N_3429);
nand U3622 (N_3622,N_3599,N_3442);
nand U3623 (N_3623,N_3568,N_3532);
and U3624 (N_3624,N_3521,N_3478);
or U3625 (N_3625,N_3428,N_3553);
and U3626 (N_3626,N_3502,N_3463);
nor U3627 (N_3627,N_3595,N_3406);
and U3628 (N_3628,N_3559,N_3440);
nand U3629 (N_3629,N_3467,N_3483);
nand U3630 (N_3630,N_3556,N_3598);
nor U3631 (N_3631,N_3527,N_3528);
and U3632 (N_3632,N_3416,N_3409);
and U3633 (N_3633,N_3587,N_3513);
and U3634 (N_3634,N_3549,N_3561);
nand U3635 (N_3635,N_3430,N_3414);
nor U3636 (N_3636,N_3570,N_3453);
nor U3637 (N_3637,N_3454,N_3546);
or U3638 (N_3638,N_3571,N_3407);
nand U3639 (N_3639,N_3590,N_3476);
or U3640 (N_3640,N_3548,N_3466);
nand U3641 (N_3641,N_3575,N_3426);
nand U3642 (N_3642,N_3584,N_3474);
and U3643 (N_3643,N_3508,N_3415);
and U3644 (N_3644,N_3572,N_3400);
nand U3645 (N_3645,N_3550,N_3431);
or U3646 (N_3646,N_3404,N_3418);
or U3647 (N_3647,N_3462,N_3580);
nand U3648 (N_3648,N_3421,N_3526);
and U3649 (N_3649,N_3558,N_3493);
and U3650 (N_3650,N_3468,N_3512);
nor U3651 (N_3651,N_3456,N_3470);
nand U3652 (N_3652,N_3560,N_3432);
xor U3653 (N_3653,N_3464,N_3417);
nand U3654 (N_3654,N_3412,N_3551);
nand U3655 (N_3655,N_3482,N_3447);
or U3656 (N_3656,N_3501,N_3492);
or U3657 (N_3657,N_3479,N_3578);
or U3658 (N_3658,N_3583,N_3405);
and U3659 (N_3659,N_3539,N_3445);
and U3660 (N_3660,N_3593,N_3510);
nor U3661 (N_3661,N_3579,N_3452);
or U3662 (N_3662,N_3564,N_3438);
or U3663 (N_3663,N_3505,N_3503);
or U3664 (N_3664,N_3459,N_3514);
and U3665 (N_3665,N_3544,N_3520);
nand U3666 (N_3666,N_3486,N_3425);
nand U3667 (N_3667,N_3413,N_3475);
nand U3668 (N_3668,N_3509,N_3562);
nor U3669 (N_3669,N_3455,N_3472);
nor U3670 (N_3670,N_3494,N_3427);
nor U3671 (N_3671,N_3555,N_3460);
and U3672 (N_3672,N_3581,N_3511);
or U3673 (N_3673,N_3519,N_3536);
and U3674 (N_3674,N_3496,N_3566);
nor U3675 (N_3675,N_3582,N_3541);
xnor U3676 (N_3676,N_3534,N_3499);
or U3677 (N_3677,N_3465,N_3591);
or U3678 (N_3678,N_3490,N_3533);
nand U3679 (N_3679,N_3515,N_3506);
or U3680 (N_3680,N_3420,N_3585);
and U3681 (N_3681,N_3422,N_3433);
nand U3682 (N_3682,N_3589,N_3489);
nand U3683 (N_3683,N_3525,N_3410);
nor U3684 (N_3684,N_3437,N_3469);
xnor U3685 (N_3685,N_3435,N_3450);
and U3686 (N_3686,N_3557,N_3597);
nor U3687 (N_3687,N_3477,N_3574);
nor U3688 (N_3688,N_3441,N_3563);
xnor U3689 (N_3689,N_3523,N_3522);
and U3690 (N_3690,N_3576,N_3458);
nand U3691 (N_3691,N_3542,N_3577);
or U3692 (N_3692,N_3529,N_3567);
xnor U3693 (N_3693,N_3484,N_3531);
nor U3694 (N_3694,N_3449,N_3401);
xor U3695 (N_3695,N_3547,N_3419);
and U3696 (N_3696,N_3436,N_3596);
or U3697 (N_3697,N_3473,N_3498);
or U3698 (N_3698,N_3552,N_3569);
nor U3699 (N_3699,N_3488,N_3446);
nand U3700 (N_3700,N_3466,N_3471);
nor U3701 (N_3701,N_3470,N_3546);
xor U3702 (N_3702,N_3400,N_3554);
nor U3703 (N_3703,N_3554,N_3477);
nor U3704 (N_3704,N_3529,N_3516);
or U3705 (N_3705,N_3410,N_3518);
nand U3706 (N_3706,N_3448,N_3568);
nor U3707 (N_3707,N_3491,N_3413);
or U3708 (N_3708,N_3479,N_3523);
nor U3709 (N_3709,N_3439,N_3599);
or U3710 (N_3710,N_3531,N_3509);
nand U3711 (N_3711,N_3491,N_3457);
and U3712 (N_3712,N_3568,N_3438);
or U3713 (N_3713,N_3548,N_3400);
and U3714 (N_3714,N_3491,N_3582);
xnor U3715 (N_3715,N_3456,N_3492);
or U3716 (N_3716,N_3498,N_3430);
nor U3717 (N_3717,N_3583,N_3469);
nor U3718 (N_3718,N_3443,N_3569);
or U3719 (N_3719,N_3478,N_3449);
or U3720 (N_3720,N_3521,N_3593);
nand U3721 (N_3721,N_3577,N_3428);
or U3722 (N_3722,N_3424,N_3542);
and U3723 (N_3723,N_3490,N_3463);
nand U3724 (N_3724,N_3461,N_3527);
nand U3725 (N_3725,N_3568,N_3504);
nor U3726 (N_3726,N_3474,N_3407);
and U3727 (N_3727,N_3510,N_3445);
nand U3728 (N_3728,N_3515,N_3466);
nor U3729 (N_3729,N_3535,N_3456);
and U3730 (N_3730,N_3499,N_3472);
nor U3731 (N_3731,N_3432,N_3558);
and U3732 (N_3732,N_3464,N_3572);
nor U3733 (N_3733,N_3440,N_3557);
or U3734 (N_3734,N_3566,N_3430);
nand U3735 (N_3735,N_3525,N_3541);
xor U3736 (N_3736,N_3431,N_3466);
nand U3737 (N_3737,N_3578,N_3528);
nor U3738 (N_3738,N_3483,N_3525);
and U3739 (N_3739,N_3434,N_3431);
nand U3740 (N_3740,N_3524,N_3444);
nor U3741 (N_3741,N_3446,N_3470);
nor U3742 (N_3742,N_3413,N_3548);
nor U3743 (N_3743,N_3458,N_3420);
nor U3744 (N_3744,N_3581,N_3448);
nor U3745 (N_3745,N_3579,N_3510);
or U3746 (N_3746,N_3528,N_3465);
nor U3747 (N_3747,N_3437,N_3454);
nand U3748 (N_3748,N_3565,N_3550);
xnor U3749 (N_3749,N_3468,N_3411);
and U3750 (N_3750,N_3585,N_3445);
or U3751 (N_3751,N_3595,N_3566);
nand U3752 (N_3752,N_3544,N_3473);
nor U3753 (N_3753,N_3581,N_3480);
and U3754 (N_3754,N_3421,N_3577);
xnor U3755 (N_3755,N_3550,N_3407);
nor U3756 (N_3756,N_3545,N_3501);
xor U3757 (N_3757,N_3540,N_3598);
and U3758 (N_3758,N_3484,N_3410);
nand U3759 (N_3759,N_3559,N_3452);
or U3760 (N_3760,N_3475,N_3483);
and U3761 (N_3761,N_3411,N_3588);
xnor U3762 (N_3762,N_3534,N_3508);
nor U3763 (N_3763,N_3573,N_3403);
nand U3764 (N_3764,N_3456,N_3495);
nand U3765 (N_3765,N_3513,N_3530);
and U3766 (N_3766,N_3558,N_3553);
and U3767 (N_3767,N_3504,N_3517);
nand U3768 (N_3768,N_3467,N_3412);
nor U3769 (N_3769,N_3468,N_3530);
and U3770 (N_3770,N_3474,N_3481);
or U3771 (N_3771,N_3526,N_3444);
xnor U3772 (N_3772,N_3499,N_3545);
or U3773 (N_3773,N_3525,N_3553);
nor U3774 (N_3774,N_3547,N_3448);
xor U3775 (N_3775,N_3418,N_3494);
or U3776 (N_3776,N_3568,N_3470);
and U3777 (N_3777,N_3467,N_3567);
nand U3778 (N_3778,N_3437,N_3557);
nor U3779 (N_3779,N_3456,N_3486);
nor U3780 (N_3780,N_3536,N_3461);
nor U3781 (N_3781,N_3487,N_3479);
and U3782 (N_3782,N_3586,N_3595);
or U3783 (N_3783,N_3506,N_3478);
or U3784 (N_3784,N_3445,N_3423);
nor U3785 (N_3785,N_3400,N_3458);
or U3786 (N_3786,N_3418,N_3466);
nor U3787 (N_3787,N_3571,N_3549);
or U3788 (N_3788,N_3421,N_3571);
nand U3789 (N_3789,N_3586,N_3521);
xnor U3790 (N_3790,N_3537,N_3558);
or U3791 (N_3791,N_3471,N_3537);
xor U3792 (N_3792,N_3483,N_3555);
nor U3793 (N_3793,N_3490,N_3549);
nand U3794 (N_3794,N_3594,N_3402);
nor U3795 (N_3795,N_3582,N_3406);
and U3796 (N_3796,N_3438,N_3525);
nor U3797 (N_3797,N_3510,N_3478);
or U3798 (N_3798,N_3580,N_3550);
and U3799 (N_3799,N_3515,N_3429);
nor U3800 (N_3800,N_3677,N_3708);
and U3801 (N_3801,N_3676,N_3692);
nor U3802 (N_3802,N_3796,N_3613);
or U3803 (N_3803,N_3721,N_3643);
and U3804 (N_3804,N_3665,N_3647);
nand U3805 (N_3805,N_3789,N_3634);
or U3806 (N_3806,N_3663,N_3642);
nor U3807 (N_3807,N_3793,N_3654);
and U3808 (N_3808,N_3726,N_3610);
nand U3809 (N_3809,N_3618,N_3783);
nand U3810 (N_3810,N_3740,N_3601);
xor U3811 (N_3811,N_3703,N_3752);
and U3812 (N_3812,N_3735,N_3685);
nand U3813 (N_3813,N_3699,N_3668);
nor U3814 (N_3814,N_3653,N_3764);
or U3815 (N_3815,N_3736,N_3652);
or U3816 (N_3816,N_3636,N_3655);
nand U3817 (N_3817,N_3730,N_3689);
or U3818 (N_3818,N_3724,N_3725);
nand U3819 (N_3819,N_3619,N_3609);
or U3820 (N_3820,N_3630,N_3626);
nor U3821 (N_3821,N_3649,N_3629);
nand U3822 (N_3822,N_3628,N_3633);
or U3823 (N_3823,N_3678,N_3760);
nand U3824 (N_3824,N_3682,N_3656);
or U3825 (N_3825,N_3651,N_3615);
nand U3826 (N_3826,N_3694,N_3777);
nor U3827 (N_3827,N_3635,N_3738);
or U3828 (N_3828,N_3706,N_3639);
nand U3829 (N_3829,N_3746,N_3720);
and U3830 (N_3830,N_3604,N_3704);
or U3831 (N_3831,N_3687,N_3693);
nand U3832 (N_3832,N_3748,N_3780);
nor U3833 (N_3833,N_3718,N_3658);
nor U3834 (N_3834,N_3648,N_3614);
and U3835 (N_3835,N_3785,N_3782);
nor U3836 (N_3836,N_3681,N_3739);
xor U3837 (N_3837,N_3766,N_3640);
nand U3838 (N_3838,N_3625,N_3744);
and U3839 (N_3839,N_3666,N_3702);
xnor U3840 (N_3840,N_3715,N_3605);
xor U3841 (N_3841,N_3747,N_3672);
xor U3842 (N_3842,N_3788,N_3617);
and U3843 (N_3843,N_3751,N_3686);
and U3844 (N_3844,N_3797,N_3753);
and U3845 (N_3845,N_3621,N_3795);
nand U3846 (N_3846,N_3798,N_3731);
or U3847 (N_3847,N_3786,N_3770);
nor U3848 (N_3848,N_3771,N_3745);
nand U3849 (N_3849,N_3632,N_3637);
nor U3850 (N_3850,N_3723,N_3659);
nor U3851 (N_3851,N_3711,N_3749);
or U3852 (N_3852,N_3719,N_3624);
nor U3853 (N_3853,N_3674,N_3696);
nor U3854 (N_3854,N_3741,N_3716);
nand U3855 (N_3855,N_3733,N_3611);
nor U3856 (N_3856,N_3644,N_3743);
or U3857 (N_3857,N_3650,N_3606);
and U3858 (N_3858,N_3622,N_3774);
or U3859 (N_3859,N_3779,N_3631);
or U3860 (N_3860,N_3729,N_3707);
and U3861 (N_3861,N_3688,N_3600);
and U3862 (N_3862,N_3742,N_3710);
and U3863 (N_3863,N_3714,N_3680);
or U3864 (N_3864,N_3683,N_3792);
or U3865 (N_3865,N_3776,N_3698);
nand U3866 (N_3866,N_3664,N_3728);
or U3867 (N_3867,N_3662,N_3709);
and U3868 (N_3868,N_3645,N_3727);
xor U3869 (N_3869,N_3608,N_3768);
and U3870 (N_3870,N_3646,N_3761);
nand U3871 (N_3871,N_3657,N_3750);
nand U3872 (N_3872,N_3756,N_3762);
nand U3873 (N_3873,N_3765,N_3775);
nor U3874 (N_3874,N_3671,N_3612);
xnor U3875 (N_3875,N_3773,N_3759);
nand U3876 (N_3876,N_3794,N_3616);
xor U3877 (N_3877,N_3763,N_3667);
nor U3878 (N_3878,N_3627,N_3670);
nand U3879 (N_3879,N_3757,N_3669);
nand U3880 (N_3880,N_3754,N_3787);
or U3881 (N_3881,N_3737,N_3673);
and U3882 (N_3882,N_3660,N_3758);
nand U3883 (N_3883,N_3712,N_3641);
xnor U3884 (N_3884,N_3701,N_3769);
nor U3885 (N_3885,N_3623,N_3691);
nor U3886 (N_3886,N_3732,N_3791);
nor U3887 (N_3887,N_3700,N_3755);
and U3888 (N_3888,N_3684,N_3638);
nor U3889 (N_3889,N_3675,N_3767);
nand U3890 (N_3890,N_3799,N_3695);
nor U3891 (N_3891,N_3661,N_3679);
nand U3892 (N_3892,N_3790,N_3603);
nand U3893 (N_3893,N_3722,N_3734);
nor U3894 (N_3894,N_3784,N_3713);
nand U3895 (N_3895,N_3781,N_3778);
nor U3896 (N_3896,N_3705,N_3717);
or U3897 (N_3897,N_3772,N_3620);
nand U3898 (N_3898,N_3690,N_3602);
nor U3899 (N_3899,N_3697,N_3607);
nor U3900 (N_3900,N_3621,N_3626);
and U3901 (N_3901,N_3716,N_3684);
and U3902 (N_3902,N_3627,N_3610);
xor U3903 (N_3903,N_3717,N_3740);
or U3904 (N_3904,N_3700,N_3637);
and U3905 (N_3905,N_3762,N_3678);
and U3906 (N_3906,N_3629,N_3690);
or U3907 (N_3907,N_3631,N_3687);
nand U3908 (N_3908,N_3600,N_3717);
nand U3909 (N_3909,N_3610,N_3672);
and U3910 (N_3910,N_3794,N_3795);
nand U3911 (N_3911,N_3611,N_3796);
nand U3912 (N_3912,N_3736,N_3715);
nand U3913 (N_3913,N_3657,N_3653);
or U3914 (N_3914,N_3628,N_3758);
nor U3915 (N_3915,N_3767,N_3772);
nor U3916 (N_3916,N_3711,N_3689);
or U3917 (N_3917,N_3687,N_3700);
or U3918 (N_3918,N_3766,N_3672);
nor U3919 (N_3919,N_3656,N_3687);
or U3920 (N_3920,N_3737,N_3601);
nand U3921 (N_3921,N_3747,N_3743);
or U3922 (N_3922,N_3728,N_3740);
or U3923 (N_3923,N_3680,N_3633);
nor U3924 (N_3924,N_3783,N_3796);
nand U3925 (N_3925,N_3627,N_3630);
nand U3926 (N_3926,N_3763,N_3703);
nand U3927 (N_3927,N_3648,N_3606);
xnor U3928 (N_3928,N_3611,N_3755);
or U3929 (N_3929,N_3776,N_3707);
nand U3930 (N_3930,N_3741,N_3687);
nand U3931 (N_3931,N_3718,N_3707);
or U3932 (N_3932,N_3733,N_3763);
or U3933 (N_3933,N_3790,N_3619);
or U3934 (N_3934,N_3720,N_3641);
nor U3935 (N_3935,N_3609,N_3798);
and U3936 (N_3936,N_3696,N_3780);
xor U3937 (N_3937,N_3635,N_3621);
and U3938 (N_3938,N_3615,N_3605);
nand U3939 (N_3939,N_3749,N_3676);
or U3940 (N_3940,N_3618,N_3769);
and U3941 (N_3941,N_3781,N_3627);
or U3942 (N_3942,N_3792,N_3741);
or U3943 (N_3943,N_3762,N_3655);
and U3944 (N_3944,N_3634,N_3607);
xnor U3945 (N_3945,N_3689,N_3713);
xor U3946 (N_3946,N_3795,N_3797);
or U3947 (N_3947,N_3715,N_3799);
nor U3948 (N_3948,N_3790,N_3604);
and U3949 (N_3949,N_3687,N_3719);
nor U3950 (N_3950,N_3713,N_3736);
nor U3951 (N_3951,N_3640,N_3722);
nand U3952 (N_3952,N_3637,N_3781);
nor U3953 (N_3953,N_3748,N_3746);
or U3954 (N_3954,N_3741,N_3720);
and U3955 (N_3955,N_3622,N_3711);
and U3956 (N_3956,N_3765,N_3616);
nand U3957 (N_3957,N_3661,N_3738);
nand U3958 (N_3958,N_3680,N_3775);
nand U3959 (N_3959,N_3658,N_3620);
or U3960 (N_3960,N_3647,N_3655);
xnor U3961 (N_3961,N_3781,N_3737);
and U3962 (N_3962,N_3619,N_3690);
nand U3963 (N_3963,N_3787,N_3743);
or U3964 (N_3964,N_3627,N_3717);
and U3965 (N_3965,N_3752,N_3706);
nand U3966 (N_3966,N_3753,N_3685);
nor U3967 (N_3967,N_3783,N_3625);
or U3968 (N_3968,N_3713,N_3686);
xor U3969 (N_3969,N_3796,N_3602);
xor U3970 (N_3970,N_3638,N_3628);
nor U3971 (N_3971,N_3709,N_3616);
or U3972 (N_3972,N_3681,N_3651);
nor U3973 (N_3973,N_3608,N_3757);
nand U3974 (N_3974,N_3706,N_3756);
nor U3975 (N_3975,N_3645,N_3644);
or U3976 (N_3976,N_3706,N_3739);
or U3977 (N_3977,N_3739,N_3717);
nand U3978 (N_3978,N_3607,N_3631);
nand U3979 (N_3979,N_3771,N_3655);
nor U3980 (N_3980,N_3708,N_3608);
nor U3981 (N_3981,N_3601,N_3758);
and U3982 (N_3982,N_3726,N_3688);
and U3983 (N_3983,N_3757,N_3602);
and U3984 (N_3984,N_3657,N_3740);
nor U3985 (N_3985,N_3687,N_3641);
nand U3986 (N_3986,N_3607,N_3794);
and U3987 (N_3987,N_3605,N_3731);
nand U3988 (N_3988,N_3786,N_3679);
nand U3989 (N_3989,N_3678,N_3738);
nand U3990 (N_3990,N_3646,N_3736);
and U3991 (N_3991,N_3613,N_3698);
nand U3992 (N_3992,N_3707,N_3723);
nor U3993 (N_3993,N_3643,N_3682);
or U3994 (N_3994,N_3729,N_3740);
and U3995 (N_3995,N_3791,N_3656);
nor U3996 (N_3996,N_3678,N_3624);
and U3997 (N_3997,N_3674,N_3734);
nand U3998 (N_3998,N_3625,N_3610);
and U3999 (N_3999,N_3777,N_3794);
and U4000 (N_4000,N_3853,N_3802);
xor U4001 (N_4001,N_3957,N_3966);
nor U4002 (N_4002,N_3890,N_3922);
xnor U4003 (N_4003,N_3836,N_3964);
nand U4004 (N_4004,N_3867,N_3872);
nor U4005 (N_4005,N_3975,N_3842);
and U4006 (N_4006,N_3807,N_3998);
or U4007 (N_4007,N_3988,N_3960);
or U4008 (N_4008,N_3892,N_3967);
xnor U4009 (N_4009,N_3951,N_3990);
or U4010 (N_4010,N_3977,N_3875);
and U4011 (N_4011,N_3815,N_3818);
and U4012 (N_4012,N_3930,N_3936);
and U4013 (N_4013,N_3885,N_3856);
and U4014 (N_4014,N_3895,N_3898);
and U4015 (N_4015,N_3834,N_3912);
nand U4016 (N_4016,N_3906,N_3968);
nand U4017 (N_4017,N_3883,N_3983);
or U4018 (N_4018,N_3826,N_3909);
nand U4019 (N_4019,N_3854,N_3910);
and U4020 (N_4020,N_3938,N_3863);
and U4021 (N_4021,N_3986,N_3978);
nand U4022 (N_4022,N_3955,N_3846);
nand U4023 (N_4023,N_3933,N_3916);
nor U4024 (N_4024,N_3991,N_3982);
or U4025 (N_4025,N_3851,N_3946);
xnor U4026 (N_4026,N_3811,N_3821);
nand U4027 (N_4027,N_3928,N_3924);
xnor U4028 (N_4028,N_3932,N_3989);
and U4029 (N_4029,N_3864,N_3993);
xnor U4030 (N_4030,N_3862,N_3943);
and U4031 (N_4031,N_3812,N_3905);
and U4032 (N_4032,N_3891,N_3958);
or U4033 (N_4033,N_3859,N_3833);
and U4034 (N_4034,N_3900,N_3825);
or U4035 (N_4035,N_3979,N_3874);
nor U4036 (N_4036,N_3828,N_3866);
and U4037 (N_4037,N_3908,N_3817);
nand U4038 (N_4038,N_3848,N_3803);
nor U4039 (N_4039,N_3861,N_3913);
nand U4040 (N_4040,N_3871,N_3839);
nor U4041 (N_4041,N_3995,N_3956);
and U4042 (N_4042,N_3844,N_3838);
nor U4043 (N_4043,N_3920,N_3927);
nor U4044 (N_4044,N_3944,N_3923);
or U4045 (N_4045,N_3840,N_3820);
or U4046 (N_4046,N_3881,N_3852);
nand U4047 (N_4047,N_3823,N_3969);
or U4048 (N_4048,N_3919,N_3873);
nand U4049 (N_4049,N_3949,N_3918);
or U4050 (N_4050,N_3808,N_3810);
and U4051 (N_4051,N_3830,N_3987);
nand U4052 (N_4052,N_3819,N_3947);
xor U4053 (N_4053,N_3915,N_3952);
or U4054 (N_4054,N_3917,N_3901);
or U4055 (N_4055,N_3880,N_3902);
nor U4056 (N_4056,N_3970,N_3876);
xor U4057 (N_4057,N_3985,N_3896);
and U4058 (N_4058,N_3904,N_3903);
nor U4059 (N_4059,N_3824,N_3835);
nor U4060 (N_4060,N_3929,N_3907);
nor U4061 (N_4061,N_3940,N_3847);
xor U4062 (N_4062,N_3996,N_3837);
and U4063 (N_4063,N_3961,N_3972);
or U4064 (N_4064,N_3877,N_3963);
or U4065 (N_4065,N_3926,N_3935);
or U4066 (N_4066,N_3804,N_3857);
nand U4067 (N_4067,N_3845,N_3860);
nand U4068 (N_4068,N_3934,N_3953);
nand U4069 (N_4069,N_3843,N_3945);
or U4070 (N_4070,N_3813,N_3822);
or U4071 (N_4071,N_3931,N_3974);
nor U4072 (N_4072,N_3981,N_3899);
and U4073 (N_4073,N_3941,N_3816);
or U4074 (N_4074,N_3962,N_3965);
nor U4075 (N_4075,N_3976,N_3894);
or U4076 (N_4076,N_3831,N_3800);
nand U4077 (N_4077,N_3994,N_3855);
nor U4078 (N_4078,N_3950,N_3911);
or U4079 (N_4079,N_3868,N_3865);
or U4080 (N_4080,N_3897,N_3999);
and U4081 (N_4081,N_3973,N_3886);
or U4082 (N_4082,N_3887,N_3849);
xor U4083 (N_4083,N_3889,N_3869);
or U4084 (N_4084,N_3942,N_3925);
nor U4085 (N_4085,N_3992,N_3878);
nor U4086 (N_4086,N_3829,N_3888);
nand U4087 (N_4087,N_3939,N_3921);
and U4088 (N_4088,N_3997,N_3884);
or U4089 (N_4089,N_3959,N_3805);
nor U4090 (N_4090,N_3870,N_3954);
or U4091 (N_4091,N_3971,N_3893);
or U4092 (N_4092,N_3914,N_3827);
and U4093 (N_4093,N_3801,N_3858);
xor U4094 (N_4094,N_3948,N_3882);
xor U4095 (N_4095,N_3984,N_3841);
nand U4096 (N_4096,N_3980,N_3879);
and U4097 (N_4097,N_3806,N_3809);
or U4098 (N_4098,N_3850,N_3814);
and U4099 (N_4099,N_3832,N_3937);
nand U4100 (N_4100,N_3885,N_3858);
and U4101 (N_4101,N_3866,N_3972);
nand U4102 (N_4102,N_3930,N_3849);
or U4103 (N_4103,N_3800,N_3815);
or U4104 (N_4104,N_3830,N_3800);
xnor U4105 (N_4105,N_3876,N_3868);
nand U4106 (N_4106,N_3940,N_3930);
nand U4107 (N_4107,N_3861,N_3895);
nand U4108 (N_4108,N_3913,N_3998);
and U4109 (N_4109,N_3926,N_3884);
nor U4110 (N_4110,N_3983,N_3821);
and U4111 (N_4111,N_3965,N_3916);
nand U4112 (N_4112,N_3878,N_3887);
or U4113 (N_4113,N_3962,N_3903);
nor U4114 (N_4114,N_3881,N_3890);
nor U4115 (N_4115,N_3966,N_3882);
and U4116 (N_4116,N_3864,N_3810);
or U4117 (N_4117,N_3891,N_3890);
nor U4118 (N_4118,N_3972,N_3917);
nand U4119 (N_4119,N_3889,N_3860);
nor U4120 (N_4120,N_3811,N_3838);
and U4121 (N_4121,N_3906,N_3869);
nor U4122 (N_4122,N_3912,N_3800);
nand U4123 (N_4123,N_3902,N_3800);
or U4124 (N_4124,N_3982,N_3890);
nand U4125 (N_4125,N_3825,N_3875);
or U4126 (N_4126,N_3858,N_3965);
or U4127 (N_4127,N_3932,N_3987);
and U4128 (N_4128,N_3864,N_3936);
or U4129 (N_4129,N_3803,N_3912);
nand U4130 (N_4130,N_3869,N_3988);
nand U4131 (N_4131,N_3862,N_3861);
or U4132 (N_4132,N_3982,N_3854);
and U4133 (N_4133,N_3913,N_3894);
and U4134 (N_4134,N_3847,N_3987);
xor U4135 (N_4135,N_3874,N_3986);
nand U4136 (N_4136,N_3997,N_3855);
nand U4137 (N_4137,N_3822,N_3964);
or U4138 (N_4138,N_3839,N_3898);
nand U4139 (N_4139,N_3961,N_3855);
nand U4140 (N_4140,N_3994,N_3838);
xor U4141 (N_4141,N_3859,N_3935);
and U4142 (N_4142,N_3906,N_3942);
nor U4143 (N_4143,N_3985,N_3993);
nor U4144 (N_4144,N_3947,N_3877);
nor U4145 (N_4145,N_3936,N_3807);
nand U4146 (N_4146,N_3843,N_3963);
xor U4147 (N_4147,N_3925,N_3970);
or U4148 (N_4148,N_3937,N_3826);
xor U4149 (N_4149,N_3813,N_3809);
and U4150 (N_4150,N_3975,N_3977);
and U4151 (N_4151,N_3890,N_3825);
and U4152 (N_4152,N_3808,N_3912);
nand U4153 (N_4153,N_3814,N_3952);
or U4154 (N_4154,N_3812,N_3882);
nor U4155 (N_4155,N_3967,N_3983);
nand U4156 (N_4156,N_3999,N_3830);
nor U4157 (N_4157,N_3985,N_3850);
or U4158 (N_4158,N_3888,N_3846);
and U4159 (N_4159,N_3864,N_3872);
nor U4160 (N_4160,N_3812,N_3926);
xor U4161 (N_4161,N_3957,N_3973);
nor U4162 (N_4162,N_3864,N_3998);
and U4163 (N_4163,N_3937,N_3839);
or U4164 (N_4164,N_3923,N_3935);
nand U4165 (N_4165,N_3941,N_3822);
or U4166 (N_4166,N_3863,N_3934);
or U4167 (N_4167,N_3860,N_3943);
nand U4168 (N_4168,N_3920,N_3997);
or U4169 (N_4169,N_3945,N_3912);
xnor U4170 (N_4170,N_3938,N_3960);
nor U4171 (N_4171,N_3857,N_3991);
or U4172 (N_4172,N_3871,N_3954);
and U4173 (N_4173,N_3846,N_3830);
and U4174 (N_4174,N_3812,N_3977);
xor U4175 (N_4175,N_3989,N_3895);
nor U4176 (N_4176,N_3855,N_3931);
nand U4177 (N_4177,N_3985,N_3860);
and U4178 (N_4178,N_3802,N_3805);
nand U4179 (N_4179,N_3894,N_3955);
and U4180 (N_4180,N_3903,N_3837);
xor U4181 (N_4181,N_3995,N_3988);
nor U4182 (N_4182,N_3850,N_3840);
or U4183 (N_4183,N_3894,N_3964);
or U4184 (N_4184,N_3909,N_3803);
and U4185 (N_4185,N_3826,N_3830);
or U4186 (N_4186,N_3923,N_3995);
nand U4187 (N_4187,N_3869,N_3876);
xnor U4188 (N_4188,N_3983,N_3990);
nor U4189 (N_4189,N_3855,N_3962);
and U4190 (N_4190,N_3985,N_3962);
nand U4191 (N_4191,N_3856,N_3835);
nor U4192 (N_4192,N_3939,N_3854);
or U4193 (N_4193,N_3864,N_3848);
or U4194 (N_4194,N_3809,N_3955);
nand U4195 (N_4195,N_3851,N_3803);
or U4196 (N_4196,N_3965,N_3912);
nor U4197 (N_4197,N_3830,N_3934);
nor U4198 (N_4198,N_3981,N_3894);
nand U4199 (N_4199,N_3939,N_3870);
nor U4200 (N_4200,N_4167,N_4157);
nand U4201 (N_4201,N_4185,N_4050);
xnor U4202 (N_4202,N_4021,N_4132);
xor U4203 (N_4203,N_4096,N_4063);
nand U4204 (N_4204,N_4009,N_4124);
or U4205 (N_4205,N_4092,N_4115);
or U4206 (N_4206,N_4056,N_4077);
nor U4207 (N_4207,N_4064,N_4154);
nor U4208 (N_4208,N_4072,N_4094);
nor U4209 (N_4209,N_4129,N_4186);
nor U4210 (N_4210,N_4147,N_4106);
nand U4211 (N_4211,N_4125,N_4017);
and U4212 (N_4212,N_4062,N_4198);
or U4213 (N_4213,N_4095,N_4194);
nand U4214 (N_4214,N_4116,N_4054);
nor U4215 (N_4215,N_4078,N_4135);
or U4216 (N_4216,N_4105,N_4032);
nor U4217 (N_4217,N_4034,N_4087);
xor U4218 (N_4218,N_4173,N_4057);
and U4219 (N_4219,N_4030,N_4025);
nand U4220 (N_4220,N_4199,N_4086);
or U4221 (N_4221,N_4182,N_4191);
or U4222 (N_4222,N_4049,N_4097);
nor U4223 (N_4223,N_4101,N_4177);
or U4224 (N_4224,N_4073,N_4022);
or U4225 (N_4225,N_4148,N_4037);
nor U4226 (N_4226,N_4012,N_4184);
nand U4227 (N_4227,N_4142,N_4175);
and U4228 (N_4228,N_4151,N_4016);
or U4229 (N_4229,N_4102,N_4163);
nor U4230 (N_4230,N_4113,N_4122);
or U4231 (N_4231,N_4059,N_4023);
nand U4232 (N_4232,N_4112,N_4061);
nor U4233 (N_4233,N_4024,N_4162);
nor U4234 (N_4234,N_4174,N_4196);
nand U4235 (N_4235,N_4153,N_4080);
nor U4236 (N_4236,N_4110,N_4014);
and U4237 (N_4237,N_4139,N_4187);
nand U4238 (N_4238,N_4130,N_4001);
xor U4239 (N_4239,N_4195,N_4085);
xor U4240 (N_4240,N_4103,N_4192);
nor U4241 (N_4241,N_4165,N_4169);
or U4242 (N_4242,N_4104,N_4107);
or U4243 (N_4243,N_4019,N_4143);
or U4244 (N_4244,N_4166,N_4045);
nand U4245 (N_4245,N_4091,N_4046);
and U4246 (N_4246,N_4099,N_4028);
nand U4247 (N_4247,N_4069,N_4141);
xnor U4248 (N_4248,N_4183,N_4120);
nor U4249 (N_4249,N_4026,N_4137);
nor U4250 (N_4250,N_4041,N_4161);
or U4251 (N_4251,N_4060,N_4089);
or U4252 (N_4252,N_4053,N_4000);
or U4253 (N_4253,N_4052,N_4190);
or U4254 (N_4254,N_4121,N_4084);
or U4255 (N_4255,N_4168,N_4181);
nor U4256 (N_4256,N_4127,N_4006);
and U4257 (N_4257,N_4179,N_4180);
and U4258 (N_4258,N_4033,N_4011);
or U4259 (N_4259,N_4070,N_4079);
or U4260 (N_4260,N_4150,N_4068);
nand U4261 (N_4261,N_4109,N_4036);
and U4262 (N_4262,N_4118,N_4083);
or U4263 (N_4263,N_4039,N_4042);
nor U4264 (N_4264,N_4015,N_4058);
xnor U4265 (N_4265,N_4020,N_4149);
nand U4266 (N_4266,N_4055,N_4136);
nor U4267 (N_4267,N_4008,N_4076);
or U4268 (N_4268,N_4065,N_4005);
nand U4269 (N_4269,N_4171,N_4040);
and U4270 (N_4270,N_4027,N_4090);
nor U4271 (N_4271,N_4035,N_4133);
nand U4272 (N_4272,N_4188,N_4164);
nand U4273 (N_4273,N_4131,N_4146);
xnor U4274 (N_4274,N_4123,N_4178);
nand U4275 (N_4275,N_4126,N_4082);
or U4276 (N_4276,N_4152,N_4100);
or U4277 (N_4277,N_4197,N_4176);
and U4278 (N_4278,N_4155,N_4158);
xnor U4279 (N_4279,N_4145,N_4159);
nand U4280 (N_4280,N_4043,N_4067);
nand U4281 (N_4281,N_4108,N_4004);
or U4282 (N_4282,N_4018,N_4074);
nor U4283 (N_4283,N_4144,N_4013);
and U4284 (N_4284,N_4007,N_4031);
nand U4285 (N_4285,N_4140,N_4114);
or U4286 (N_4286,N_4010,N_4002);
nor U4287 (N_4287,N_4156,N_4047);
nand U4288 (N_4288,N_4189,N_4003);
or U4289 (N_4289,N_4071,N_4172);
nor U4290 (N_4290,N_4193,N_4066);
nor U4291 (N_4291,N_4048,N_4170);
and U4292 (N_4292,N_4134,N_4138);
xor U4293 (N_4293,N_4038,N_4160);
and U4294 (N_4294,N_4051,N_4044);
nand U4295 (N_4295,N_4119,N_4111);
and U4296 (N_4296,N_4128,N_4075);
nand U4297 (N_4297,N_4117,N_4029);
nand U4298 (N_4298,N_4098,N_4088);
and U4299 (N_4299,N_4081,N_4093);
and U4300 (N_4300,N_4005,N_4077);
nor U4301 (N_4301,N_4057,N_4107);
nor U4302 (N_4302,N_4009,N_4139);
and U4303 (N_4303,N_4005,N_4119);
nand U4304 (N_4304,N_4062,N_4032);
or U4305 (N_4305,N_4132,N_4057);
or U4306 (N_4306,N_4192,N_4195);
and U4307 (N_4307,N_4192,N_4129);
xor U4308 (N_4308,N_4022,N_4069);
and U4309 (N_4309,N_4136,N_4052);
and U4310 (N_4310,N_4158,N_4091);
nor U4311 (N_4311,N_4143,N_4053);
nor U4312 (N_4312,N_4027,N_4097);
nand U4313 (N_4313,N_4168,N_4016);
and U4314 (N_4314,N_4180,N_4046);
and U4315 (N_4315,N_4133,N_4197);
nor U4316 (N_4316,N_4144,N_4122);
or U4317 (N_4317,N_4030,N_4054);
or U4318 (N_4318,N_4014,N_4167);
and U4319 (N_4319,N_4151,N_4003);
or U4320 (N_4320,N_4192,N_4114);
nand U4321 (N_4321,N_4027,N_4174);
or U4322 (N_4322,N_4025,N_4113);
xnor U4323 (N_4323,N_4167,N_4089);
nor U4324 (N_4324,N_4165,N_4011);
or U4325 (N_4325,N_4077,N_4144);
or U4326 (N_4326,N_4012,N_4013);
nand U4327 (N_4327,N_4026,N_4112);
nor U4328 (N_4328,N_4170,N_4080);
xor U4329 (N_4329,N_4102,N_4085);
or U4330 (N_4330,N_4184,N_4158);
nand U4331 (N_4331,N_4185,N_4194);
nand U4332 (N_4332,N_4033,N_4030);
nor U4333 (N_4333,N_4165,N_4062);
nor U4334 (N_4334,N_4140,N_4080);
or U4335 (N_4335,N_4097,N_4186);
or U4336 (N_4336,N_4161,N_4153);
or U4337 (N_4337,N_4132,N_4122);
nor U4338 (N_4338,N_4179,N_4103);
nand U4339 (N_4339,N_4050,N_4106);
nand U4340 (N_4340,N_4154,N_4027);
and U4341 (N_4341,N_4154,N_4151);
or U4342 (N_4342,N_4135,N_4042);
nand U4343 (N_4343,N_4050,N_4031);
xnor U4344 (N_4344,N_4178,N_4149);
and U4345 (N_4345,N_4143,N_4156);
and U4346 (N_4346,N_4103,N_4146);
xnor U4347 (N_4347,N_4100,N_4118);
and U4348 (N_4348,N_4178,N_4055);
nand U4349 (N_4349,N_4194,N_4104);
and U4350 (N_4350,N_4039,N_4143);
and U4351 (N_4351,N_4075,N_4085);
and U4352 (N_4352,N_4102,N_4095);
or U4353 (N_4353,N_4185,N_4045);
and U4354 (N_4354,N_4025,N_4126);
and U4355 (N_4355,N_4124,N_4199);
or U4356 (N_4356,N_4198,N_4079);
or U4357 (N_4357,N_4191,N_4111);
and U4358 (N_4358,N_4108,N_4151);
nand U4359 (N_4359,N_4066,N_4058);
or U4360 (N_4360,N_4167,N_4174);
xnor U4361 (N_4361,N_4090,N_4016);
or U4362 (N_4362,N_4059,N_4169);
nor U4363 (N_4363,N_4015,N_4174);
nor U4364 (N_4364,N_4096,N_4034);
and U4365 (N_4365,N_4096,N_4067);
and U4366 (N_4366,N_4016,N_4014);
xor U4367 (N_4367,N_4145,N_4005);
and U4368 (N_4368,N_4116,N_4091);
nor U4369 (N_4369,N_4136,N_4157);
and U4370 (N_4370,N_4065,N_4152);
and U4371 (N_4371,N_4027,N_4142);
or U4372 (N_4372,N_4023,N_4113);
or U4373 (N_4373,N_4117,N_4033);
and U4374 (N_4374,N_4170,N_4026);
or U4375 (N_4375,N_4113,N_4156);
nor U4376 (N_4376,N_4026,N_4081);
xor U4377 (N_4377,N_4197,N_4084);
nand U4378 (N_4378,N_4026,N_4079);
nor U4379 (N_4379,N_4131,N_4042);
and U4380 (N_4380,N_4049,N_4182);
and U4381 (N_4381,N_4159,N_4010);
or U4382 (N_4382,N_4087,N_4183);
and U4383 (N_4383,N_4168,N_4185);
and U4384 (N_4384,N_4063,N_4162);
nor U4385 (N_4385,N_4006,N_4172);
and U4386 (N_4386,N_4026,N_4017);
and U4387 (N_4387,N_4086,N_4119);
or U4388 (N_4388,N_4063,N_4172);
nand U4389 (N_4389,N_4145,N_4011);
or U4390 (N_4390,N_4057,N_4056);
nand U4391 (N_4391,N_4179,N_4049);
nor U4392 (N_4392,N_4031,N_4115);
nand U4393 (N_4393,N_4192,N_4123);
and U4394 (N_4394,N_4127,N_4115);
xnor U4395 (N_4395,N_4104,N_4140);
nand U4396 (N_4396,N_4155,N_4133);
or U4397 (N_4397,N_4172,N_4027);
nand U4398 (N_4398,N_4143,N_4042);
nand U4399 (N_4399,N_4042,N_4050);
nand U4400 (N_4400,N_4201,N_4243);
nand U4401 (N_4401,N_4350,N_4258);
nor U4402 (N_4402,N_4333,N_4331);
nor U4403 (N_4403,N_4394,N_4286);
nor U4404 (N_4404,N_4227,N_4299);
nand U4405 (N_4405,N_4317,N_4265);
and U4406 (N_4406,N_4282,N_4386);
and U4407 (N_4407,N_4215,N_4303);
xnor U4408 (N_4408,N_4336,N_4373);
xor U4409 (N_4409,N_4345,N_4232);
and U4410 (N_4410,N_4272,N_4398);
or U4411 (N_4411,N_4221,N_4237);
and U4412 (N_4412,N_4295,N_4359);
xnor U4413 (N_4413,N_4250,N_4294);
or U4414 (N_4414,N_4288,N_4206);
xnor U4415 (N_4415,N_4363,N_4252);
xor U4416 (N_4416,N_4287,N_4328);
or U4417 (N_4417,N_4263,N_4271);
or U4418 (N_4418,N_4311,N_4378);
nand U4419 (N_4419,N_4259,N_4315);
nand U4420 (N_4420,N_4372,N_4285);
and U4421 (N_4421,N_4329,N_4321);
nor U4422 (N_4422,N_4360,N_4326);
nor U4423 (N_4423,N_4205,N_4224);
and U4424 (N_4424,N_4323,N_4383);
nand U4425 (N_4425,N_4318,N_4377);
nor U4426 (N_4426,N_4268,N_4313);
nor U4427 (N_4427,N_4385,N_4381);
or U4428 (N_4428,N_4247,N_4393);
or U4429 (N_4429,N_4217,N_4353);
or U4430 (N_4430,N_4355,N_4369);
nand U4431 (N_4431,N_4364,N_4256);
and U4432 (N_4432,N_4273,N_4362);
nand U4433 (N_4433,N_4339,N_4248);
nor U4434 (N_4434,N_4375,N_4255);
nand U4435 (N_4435,N_4361,N_4260);
nor U4436 (N_4436,N_4220,N_4396);
and U4437 (N_4437,N_4274,N_4322);
or U4438 (N_4438,N_4334,N_4305);
xor U4439 (N_4439,N_4214,N_4204);
nor U4440 (N_4440,N_4240,N_4283);
nand U4441 (N_4441,N_4209,N_4236);
nor U4442 (N_4442,N_4207,N_4325);
nor U4443 (N_4443,N_4357,N_4332);
xor U4444 (N_4444,N_4292,N_4289);
and U4445 (N_4445,N_4314,N_4370);
nand U4446 (N_4446,N_4399,N_4269);
nor U4447 (N_4447,N_4242,N_4379);
xor U4448 (N_4448,N_4210,N_4275);
or U4449 (N_4449,N_4284,N_4277);
and U4450 (N_4450,N_4307,N_4281);
nand U4451 (N_4451,N_4278,N_4327);
nor U4452 (N_4452,N_4293,N_4230);
nand U4453 (N_4453,N_4366,N_4392);
xor U4454 (N_4454,N_4342,N_4262);
nor U4455 (N_4455,N_4238,N_4397);
or U4456 (N_4456,N_4212,N_4233);
or U4457 (N_4457,N_4390,N_4337);
xor U4458 (N_4458,N_4382,N_4291);
or U4459 (N_4459,N_4203,N_4229);
xnor U4460 (N_4460,N_4228,N_4312);
and U4461 (N_4461,N_4267,N_4225);
xor U4462 (N_4462,N_4343,N_4202);
and U4463 (N_4463,N_4388,N_4344);
nor U4464 (N_4464,N_4304,N_4368);
and U4465 (N_4465,N_4223,N_4395);
and U4466 (N_4466,N_4219,N_4308);
or U4467 (N_4467,N_4348,N_4310);
xnor U4468 (N_4468,N_4371,N_4244);
nor U4469 (N_4469,N_4261,N_4222);
xor U4470 (N_4470,N_4249,N_4264);
nor U4471 (N_4471,N_4276,N_4320);
or U4472 (N_4472,N_4356,N_4266);
nor U4473 (N_4473,N_4352,N_4316);
nor U4474 (N_4474,N_4226,N_4241);
or U4475 (N_4475,N_4257,N_4367);
nand U4476 (N_4476,N_4380,N_4374);
nand U4477 (N_4477,N_4306,N_4302);
nor U4478 (N_4478,N_4200,N_4330);
or U4479 (N_4479,N_4349,N_4246);
and U4480 (N_4480,N_4384,N_4376);
or U4481 (N_4481,N_4235,N_4338);
or U4482 (N_4482,N_4347,N_4279);
nand U4483 (N_4483,N_4245,N_4253);
and U4484 (N_4484,N_4213,N_4296);
nand U4485 (N_4485,N_4254,N_4324);
nor U4486 (N_4486,N_4319,N_4351);
nand U4487 (N_4487,N_4309,N_4365);
nor U4488 (N_4488,N_4298,N_4297);
and U4489 (N_4489,N_4234,N_4335);
nand U4490 (N_4490,N_4218,N_4300);
nor U4491 (N_4491,N_4251,N_4270);
or U4492 (N_4492,N_4208,N_4389);
nor U4493 (N_4493,N_4216,N_4290);
or U4494 (N_4494,N_4387,N_4358);
xor U4495 (N_4495,N_4354,N_4391);
or U4496 (N_4496,N_4340,N_4280);
and U4497 (N_4497,N_4346,N_4341);
nor U4498 (N_4498,N_4301,N_4239);
or U4499 (N_4499,N_4211,N_4231);
or U4500 (N_4500,N_4265,N_4288);
xnor U4501 (N_4501,N_4281,N_4241);
nand U4502 (N_4502,N_4278,N_4268);
or U4503 (N_4503,N_4382,N_4203);
or U4504 (N_4504,N_4261,N_4351);
nand U4505 (N_4505,N_4354,N_4292);
nor U4506 (N_4506,N_4379,N_4287);
or U4507 (N_4507,N_4320,N_4313);
nor U4508 (N_4508,N_4349,N_4379);
xor U4509 (N_4509,N_4233,N_4386);
nand U4510 (N_4510,N_4267,N_4355);
nor U4511 (N_4511,N_4251,N_4235);
nor U4512 (N_4512,N_4359,N_4337);
nand U4513 (N_4513,N_4268,N_4210);
xor U4514 (N_4514,N_4267,N_4335);
or U4515 (N_4515,N_4296,N_4200);
or U4516 (N_4516,N_4382,N_4370);
or U4517 (N_4517,N_4271,N_4250);
nor U4518 (N_4518,N_4351,N_4201);
and U4519 (N_4519,N_4352,N_4203);
or U4520 (N_4520,N_4397,N_4247);
nand U4521 (N_4521,N_4218,N_4274);
or U4522 (N_4522,N_4249,N_4324);
nor U4523 (N_4523,N_4359,N_4347);
nand U4524 (N_4524,N_4230,N_4328);
and U4525 (N_4525,N_4321,N_4299);
nand U4526 (N_4526,N_4331,N_4388);
or U4527 (N_4527,N_4369,N_4214);
nand U4528 (N_4528,N_4302,N_4380);
and U4529 (N_4529,N_4307,N_4343);
xnor U4530 (N_4530,N_4279,N_4271);
nand U4531 (N_4531,N_4233,N_4352);
nand U4532 (N_4532,N_4228,N_4337);
or U4533 (N_4533,N_4284,N_4332);
xnor U4534 (N_4534,N_4281,N_4236);
and U4535 (N_4535,N_4304,N_4318);
xnor U4536 (N_4536,N_4272,N_4371);
or U4537 (N_4537,N_4368,N_4301);
or U4538 (N_4538,N_4382,N_4297);
nor U4539 (N_4539,N_4246,N_4341);
nand U4540 (N_4540,N_4319,N_4219);
and U4541 (N_4541,N_4205,N_4213);
nor U4542 (N_4542,N_4281,N_4352);
nor U4543 (N_4543,N_4292,N_4238);
or U4544 (N_4544,N_4220,N_4274);
and U4545 (N_4545,N_4290,N_4322);
or U4546 (N_4546,N_4379,N_4300);
xor U4547 (N_4547,N_4352,N_4334);
nor U4548 (N_4548,N_4207,N_4322);
and U4549 (N_4549,N_4341,N_4335);
or U4550 (N_4550,N_4213,N_4347);
xor U4551 (N_4551,N_4336,N_4309);
nand U4552 (N_4552,N_4381,N_4323);
nand U4553 (N_4553,N_4271,N_4318);
or U4554 (N_4554,N_4215,N_4332);
or U4555 (N_4555,N_4332,N_4254);
or U4556 (N_4556,N_4340,N_4208);
nand U4557 (N_4557,N_4204,N_4350);
xnor U4558 (N_4558,N_4253,N_4380);
or U4559 (N_4559,N_4382,N_4296);
nor U4560 (N_4560,N_4302,N_4287);
nand U4561 (N_4561,N_4273,N_4219);
xor U4562 (N_4562,N_4386,N_4385);
nor U4563 (N_4563,N_4262,N_4354);
and U4564 (N_4564,N_4243,N_4209);
and U4565 (N_4565,N_4355,N_4337);
nand U4566 (N_4566,N_4227,N_4272);
nand U4567 (N_4567,N_4209,N_4294);
nor U4568 (N_4568,N_4239,N_4235);
nand U4569 (N_4569,N_4263,N_4350);
and U4570 (N_4570,N_4372,N_4366);
or U4571 (N_4571,N_4351,N_4356);
nor U4572 (N_4572,N_4335,N_4206);
nand U4573 (N_4573,N_4262,N_4335);
nand U4574 (N_4574,N_4339,N_4367);
xnor U4575 (N_4575,N_4382,N_4237);
and U4576 (N_4576,N_4356,N_4204);
xnor U4577 (N_4577,N_4382,N_4396);
and U4578 (N_4578,N_4265,N_4202);
nand U4579 (N_4579,N_4227,N_4208);
and U4580 (N_4580,N_4374,N_4255);
and U4581 (N_4581,N_4394,N_4372);
nor U4582 (N_4582,N_4346,N_4359);
or U4583 (N_4583,N_4285,N_4393);
and U4584 (N_4584,N_4212,N_4290);
nor U4585 (N_4585,N_4308,N_4206);
nand U4586 (N_4586,N_4340,N_4368);
and U4587 (N_4587,N_4281,N_4379);
and U4588 (N_4588,N_4253,N_4220);
nor U4589 (N_4589,N_4322,N_4295);
or U4590 (N_4590,N_4295,N_4273);
or U4591 (N_4591,N_4225,N_4266);
nand U4592 (N_4592,N_4238,N_4293);
or U4593 (N_4593,N_4273,N_4216);
and U4594 (N_4594,N_4352,N_4306);
nor U4595 (N_4595,N_4395,N_4379);
nor U4596 (N_4596,N_4364,N_4354);
xor U4597 (N_4597,N_4317,N_4348);
nor U4598 (N_4598,N_4229,N_4319);
nand U4599 (N_4599,N_4307,N_4396);
nor U4600 (N_4600,N_4564,N_4562);
nor U4601 (N_4601,N_4588,N_4563);
xnor U4602 (N_4602,N_4423,N_4528);
nor U4603 (N_4603,N_4538,N_4558);
and U4604 (N_4604,N_4576,N_4452);
or U4605 (N_4605,N_4550,N_4505);
and U4606 (N_4606,N_4593,N_4549);
and U4607 (N_4607,N_4532,N_4465);
nand U4608 (N_4608,N_4531,N_4421);
and U4609 (N_4609,N_4493,N_4574);
and U4610 (N_4610,N_4568,N_4419);
nor U4611 (N_4611,N_4518,N_4583);
or U4612 (N_4612,N_4506,N_4468);
xor U4613 (N_4613,N_4447,N_4542);
nand U4614 (N_4614,N_4485,N_4488);
and U4615 (N_4615,N_4402,N_4596);
nor U4616 (N_4616,N_4536,N_4424);
and U4617 (N_4617,N_4586,N_4409);
xnor U4618 (N_4618,N_4579,N_4438);
or U4619 (N_4619,N_4565,N_4541);
nand U4620 (N_4620,N_4498,N_4557);
and U4621 (N_4621,N_4415,N_4501);
or U4622 (N_4622,N_4495,N_4537);
nor U4623 (N_4623,N_4560,N_4472);
nor U4624 (N_4624,N_4418,N_4570);
nor U4625 (N_4625,N_4470,N_4426);
xor U4626 (N_4626,N_4522,N_4578);
or U4627 (N_4627,N_4546,N_4408);
and U4628 (N_4628,N_4496,N_4575);
nand U4629 (N_4629,N_4484,N_4510);
and U4630 (N_4630,N_4569,N_4490);
xor U4631 (N_4631,N_4425,N_4428);
and U4632 (N_4632,N_4430,N_4526);
nor U4633 (N_4633,N_4442,N_4435);
nor U4634 (N_4634,N_4405,N_4420);
and U4635 (N_4635,N_4450,N_4494);
nor U4636 (N_4636,N_4486,N_4535);
or U4637 (N_4637,N_4410,N_4417);
nor U4638 (N_4638,N_4487,N_4509);
and U4639 (N_4639,N_4571,N_4585);
nor U4640 (N_4640,N_4414,N_4521);
nor U4641 (N_4641,N_4413,N_4553);
and U4642 (N_4642,N_4483,N_4469);
and U4643 (N_4643,N_4590,N_4489);
nor U4644 (N_4644,N_4540,N_4556);
and U4645 (N_4645,N_4457,N_4476);
nand U4646 (N_4646,N_4534,N_4459);
and U4647 (N_4647,N_4561,N_4401);
nand U4648 (N_4648,N_4422,N_4491);
nor U4649 (N_4649,N_4589,N_4427);
and U4650 (N_4650,N_4448,N_4530);
nor U4651 (N_4651,N_4591,N_4584);
or U4652 (N_4652,N_4441,N_4503);
and U4653 (N_4653,N_4524,N_4406);
nand U4654 (N_4654,N_4523,N_4411);
nor U4655 (N_4655,N_4434,N_4543);
and U4656 (N_4656,N_4516,N_4467);
or U4657 (N_4657,N_4461,N_4512);
nor U4658 (N_4658,N_4429,N_4592);
and U4659 (N_4659,N_4480,N_4548);
nor U4660 (N_4660,N_4481,N_4527);
or U4661 (N_4661,N_4400,N_4455);
nor U4662 (N_4662,N_4594,N_4407);
xnor U4663 (N_4663,N_4511,N_4499);
or U4664 (N_4664,N_4500,N_4513);
and U4665 (N_4665,N_4597,N_4595);
xor U4666 (N_4666,N_4525,N_4433);
xnor U4667 (N_4667,N_4566,N_4559);
nand U4668 (N_4668,N_4432,N_4473);
nand U4669 (N_4669,N_4577,N_4464);
nand U4670 (N_4670,N_4547,N_4479);
nand U4671 (N_4671,N_4555,N_4443);
nor U4672 (N_4672,N_4462,N_4474);
nor U4673 (N_4673,N_4504,N_4475);
nand U4674 (N_4674,N_4519,N_4412);
nor U4675 (N_4675,N_4444,N_4431);
nor U4676 (N_4676,N_4508,N_4437);
nor U4677 (N_4677,N_4544,N_4436);
nand U4678 (N_4678,N_4445,N_4582);
or U4679 (N_4679,N_4599,N_4458);
nor U4680 (N_4680,N_4454,N_4533);
nand U4681 (N_4681,N_4416,N_4439);
or U4682 (N_4682,N_4554,N_4545);
nor U4683 (N_4683,N_4460,N_4449);
nor U4684 (N_4684,N_4463,N_4580);
or U4685 (N_4685,N_4466,N_4529);
nor U4686 (N_4686,N_4572,N_4477);
and U4687 (N_4687,N_4471,N_4517);
or U4688 (N_4688,N_4581,N_4492);
or U4689 (N_4689,N_4404,N_4456);
xor U4690 (N_4690,N_4567,N_4478);
nand U4691 (N_4691,N_4587,N_4446);
nor U4692 (N_4692,N_4573,N_4482);
and U4693 (N_4693,N_4598,N_4552);
nand U4694 (N_4694,N_4520,N_4507);
nand U4695 (N_4695,N_4497,N_4451);
nor U4696 (N_4696,N_4514,N_4515);
nor U4697 (N_4697,N_4539,N_4453);
nor U4698 (N_4698,N_4403,N_4502);
or U4699 (N_4699,N_4440,N_4551);
and U4700 (N_4700,N_4452,N_4526);
nor U4701 (N_4701,N_4493,N_4588);
nand U4702 (N_4702,N_4584,N_4482);
and U4703 (N_4703,N_4531,N_4496);
or U4704 (N_4704,N_4427,N_4485);
or U4705 (N_4705,N_4545,N_4422);
nand U4706 (N_4706,N_4456,N_4529);
and U4707 (N_4707,N_4454,N_4491);
nand U4708 (N_4708,N_4424,N_4525);
nand U4709 (N_4709,N_4527,N_4419);
xnor U4710 (N_4710,N_4419,N_4596);
nand U4711 (N_4711,N_4566,N_4443);
or U4712 (N_4712,N_4580,N_4435);
or U4713 (N_4713,N_4550,N_4454);
nand U4714 (N_4714,N_4454,N_4477);
nor U4715 (N_4715,N_4454,N_4489);
or U4716 (N_4716,N_4539,N_4410);
and U4717 (N_4717,N_4509,N_4450);
nor U4718 (N_4718,N_4514,N_4511);
nand U4719 (N_4719,N_4578,N_4454);
nor U4720 (N_4720,N_4578,N_4478);
nor U4721 (N_4721,N_4557,N_4553);
nor U4722 (N_4722,N_4440,N_4562);
and U4723 (N_4723,N_4422,N_4401);
xor U4724 (N_4724,N_4432,N_4488);
nor U4725 (N_4725,N_4455,N_4471);
or U4726 (N_4726,N_4581,N_4470);
nand U4727 (N_4727,N_4414,N_4593);
nor U4728 (N_4728,N_4595,N_4444);
nand U4729 (N_4729,N_4486,N_4479);
and U4730 (N_4730,N_4434,N_4505);
or U4731 (N_4731,N_4428,N_4463);
and U4732 (N_4732,N_4482,N_4424);
nor U4733 (N_4733,N_4515,N_4574);
nor U4734 (N_4734,N_4565,N_4595);
or U4735 (N_4735,N_4501,N_4414);
or U4736 (N_4736,N_4444,N_4421);
nand U4737 (N_4737,N_4428,N_4435);
nand U4738 (N_4738,N_4507,N_4504);
or U4739 (N_4739,N_4402,N_4576);
or U4740 (N_4740,N_4509,N_4406);
and U4741 (N_4741,N_4520,N_4576);
nor U4742 (N_4742,N_4507,N_4491);
nor U4743 (N_4743,N_4471,N_4533);
nor U4744 (N_4744,N_4484,N_4540);
nor U4745 (N_4745,N_4451,N_4562);
or U4746 (N_4746,N_4483,N_4562);
nor U4747 (N_4747,N_4557,N_4596);
or U4748 (N_4748,N_4404,N_4441);
or U4749 (N_4749,N_4478,N_4443);
nor U4750 (N_4750,N_4410,N_4589);
and U4751 (N_4751,N_4451,N_4494);
or U4752 (N_4752,N_4538,N_4536);
nand U4753 (N_4753,N_4478,N_4541);
and U4754 (N_4754,N_4537,N_4443);
nor U4755 (N_4755,N_4460,N_4444);
xnor U4756 (N_4756,N_4423,N_4477);
nor U4757 (N_4757,N_4561,N_4485);
and U4758 (N_4758,N_4504,N_4533);
and U4759 (N_4759,N_4474,N_4533);
nand U4760 (N_4760,N_4519,N_4575);
and U4761 (N_4761,N_4431,N_4470);
xnor U4762 (N_4762,N_4414,N_4454);
and U4763 (N_4763,N_4548,N_4507);
nor U4764 (N_4764,N_4419,N_4522);
and U4765 (N_4765,N_4553,N_4493);
nand U4766 (N_4766,N_4422,N_4528);
and U4767 (N_4767,N_4485,N_4430);
and U4768 (N_4768,N_4496,N_4585);
xnor U4769 (N_4769,N_4543,N_4505);
and U4770 (N_4770,N_4431,N_4551);
or U4771 (N_4771,N_4420,N_4552);
or U4772 (N_4772,N_4563,N_4417);
or U4773 (N_4773,N_4442,N_4456);
nand U4774 (N_4774,N_4412,N_4569);
nor U4775 (N_4775,N_4532,N_4484);
xnor U4776 (N_4776,N_4464,N_4555);
nor U4777 (N_4777,N_4524,N_4583);
or U4778 (N_4778,N_4421,N_4591);
or U4779 (N_4779,N_4564,N_4460);
or U4780 (N_4780,N_4406,N_4541);
or U4781 (N_4781,N_4499,N_4560);
or U4782 (N_4782,N_4468,N_4458);
or U4783 (N_4783,N_4400,N_4413);
nand U4784 (N_4784,N_4411,N_4568);
and U4785 (N_4785,N_4554,N_4512);
nand U4786 (N_4786,N_4560,N_4457);
nand U4787 (N_4787,N_4468,N_4519);
and U4788 (N_4788,N_4460,N_4526);
nand U4789 (N_4789,N_4444,N_4477);
xor U4790 (N_4790,N_4408,N_4588);
or U4791 (N_4791,N_4554,N_4566);
xnor U4792 (N_4792,N_4400,N_4451);
and U4793 (N_4793,N_4481,N_4480);
or U4794 (N_4794,N_4400,N_4545);
or U4795 (N_4795,N_4543,N_4430);
and U4796 (N_4796,N_4464,N_4510);
and U4797 (N_4797,N_4551,N_4588);
or U4798 (N_4798,N_4428,N_4551);
and U4799 (N_4799,N_4463,N_4586);
and U4800 (N_4800,N_4778,N_4621);
and U4801 (N_4801,N_4761,N_4714);
xor U4802 (N_4802,N_4796,N_4786);
nor U4803 (N_4803,N_4752,N_4660);
or U4804 (N_4804,N_4722,N_4687);
and U4805 (N_4805,N_4609,N_4630);
nand U4806 (N_4806,N_4653,N_4707);
and U4807 (N_4807,N_4647,N_4725);
nor U4808 (N_4808,N_4674,N_4741);
nand U4809 (N_4809,N_4746,N_4650);
nor U4810 (N_4810,N_4709,N_4755);
and U4811 (N_4811,N_4717,N_4777);
nand U4812 (N_4812,N_4688,N_4679);
nor U4813 (N_4813,N_4624,N_4715);
or U4814 (N_4814,N_4692,N_4771);
nor U4815 (N_4815,N_4754,N_4603);
nand U4816 (N_4816,N_4618,N_4691);
nand U4817 (N_4817,N_4736,N_4774);
nand U4818 (N_4818,N_4671,N_4764);
nand U4819 (N_4819,N_4765,N_4788);
or U4820 (N_4820,N_4690,N_4610);
xnor U4821 (N_4821,N_4742,N_4727);
or U4822 (N_4822,N_4667,N_4748);
and U4823 (N_4823,N_4606,N_4661);
and U4824 (N_4824,N_4682,N_4613);
nor U4825 (N_4825,N_4625,N_4795);
or U4826 (N_4826,N_4684,N_4734);
or U4827 (N_4827,N_4602,N_4608);
or U4828 (N_4828,N_4652,N_4644);
nand U4829 (N_4829,N_4763,N_4723);
and U4830 (N_4830,N_4677,N_4782);
and U4831 (N_4831,N_4783,N_4651);
and U4832 (N_4832,N_4766,N_4750);
xnor U4833 (N_4833,N_4739,N_4798);
and U4834 (N_4834,N_4775,N_4768);
and U4835 (N_4835,N_4640,N_4749);
and U4836 (N_4836,N_4635,N_4646);
or U4837 (N_4837,N_4681,N_4601);
xnor U4838 (N_4838,N_4716,N_4797);
nand U4839 (N_4839,N_4724,N_4605);
xnor U4840 (N_4840,N_4631,N_4673);
and U4841 (N_4841,N_4637,N_4718);
and U4842 (N_4842,N_4683,N_4728);
nor U4843 (N_4843,N_4735,N_4698);
nor U4844 (N_4844,N_4669,N_4657);
and U4845 (N_4845,N_4784,N_4655);
nand U4846 (N_4846,N_4600,N_4665);
nand U4847 (N_4847,N_4738,N_4689);
and U4848 (N_4848,N_4781,N_4776);
xnor U4849 (N_4849,N_4706,N_4616);
nand U4850 (N_4850,N_4703,N_4695);
or U4851 (N_4851,N_4641,N_4792);
nor U4852 (N_4852,N_4769,N_4619);
or U4853 (N_4853,N_4634,N_4785);
and U4854 (N_4854,N_4756,N_4753);
nand U4855 (N_4855,N_4731,N_4713);
or U4856 (N_4856,N_4629,N_4611);
nand U4857 (N_4857,N_4656,N_4628);
and U4858 (N_4858,N_4666,N_4626);
xnor U4859 (N_4859,N_4614,N_4676);
xnor U4860 (N_4860,N_4649,N_4793);
nor U4861 (N_4861,N_4732,N_4789);
nor U4862 (N_4862,N_4697,N_4773);
or U4863 (N_4863,N_4708,N_4758);
nor U4864 (N_4864,N_4744,N_4699);
and U4865 (N_4865,N_4721,N_4615);
nand U4866 (N_4866,N_4643,N_4623);
nor U4867 (N_4867,N_4604,N_4730);
or U4868 (N_4868,N_4694,N_4791);
nor U4869 (N_4869,N_4638,N_4607);
and U4870 (N_4870,N_4664,N_4701);
xor U4871 (N_4871,N_4790,N_4685);
xnor U4872 (N_4872,N_4743,N_4719);
nor U4873 (N_4873,N_4747,N_4762);
nand U4874 (N_4874,N_4675,N_4711);
and U4875 (N_4875,N_4659,N_4670);
nand U4876 (N_4876,N_4693,N_4642);
nand U4877 (N_4877,N_4733,N_4726);
or U4878 (N_4878,N_4680,N_4767);
or U4879 (N_4879,N_4696,N_4612);
xor U4880 (N_4880,N_4787,N_4627);
or U4881 (N_4881,N_4794,N_4658);
xnor U4882 (N_4882,N_4751,N_4648);
and U4883 (N_4883,N_4757,N_4759);
and U4884 (N_4884,N_4705,N_4672);
and U4885 (N_4885,N_4633,N_4704);
nand U4886 (N_4886,N_4620,N_4654);
nor U4887 (N_4887,N_4645,N_4780);
and U4888 (N_4888,N_4720,N_4770);
nand U4889 (N_4889,N_4772,N_4712);
nand U4890 (N_4890,N_4729,N_4636);
or U4891 (N_4891,N_4686,N_4617);
and U4892 (N_4892,N_4745,N_4740);
nor U4893 (N_4893,N_4668,N_4700);
nand U4894 (N_4894,N_4737,N_4622);
and U4895 (N_4895,N_4678,N_4710);
or U4896 (N_4896,N_4799,N_4760);
and U4897 (N_4897,N_4702,N_4639);
nor U4898 (N_4898,N_4632,N_4663);
xor U4899 (N_4899,N_4662,N_4779);
nand U4900 (N_4900,N_4776,N_4744);
or U4901 (N_4901,N_4692,N_4661);
or U4902 (N_4902,N_4651,N_4653);
xnor U4903 (N_4903,N_4606,N_4729);
or U4904 (N_4904,N_4630,N_4771);
and U4905 (N_4905,N_4797,N_4701);
or U4906 (N_4906,N_4676,N_4769);
and U4907 (N_4907,N_4684,N_4796);
or U4908 (N_4908,N_4676,N_4776);
or U4909 (N_4909,N_4706,N_4689);
nand U4910 (N_4910,N_4701,N_4740);
or U4911 (N_4911,N_4750,N_4745);
nor U4912 (N_4912,N_4639,N_4654);
nand U4913 (N_4913,N_4648,N_4676);
nand U4914 (N_4914,N_4641,N_4661);
and U4915 (N_4915,N_4665,N_4689);
xor U4916 (N_4916,N_4785,N_4723);
nor U4917 (N_4917,N_4615,N_4636);
nor U4918 (N_4918,N_4770,N_4730);
nor U4919 (N_4919,N_4619,N_4714);
and U4920 (N_4920,N_4615,N_4611);
and U4921 (N_4921,N_4773,N_4602);
nor U4922 (N_4922,N_4681,N_4620);
xnor U4923 (N_4923,N_4609,N_4660);
or U4924 (N_4924,N_4651,N_4677);
and U4925 (N_4925,N_4682,N_4783);
nor U4926 (N_4926,N_4600,N_4795);
and U4927 (N_4927,N_4656,N_4707);
nor U4928 (N_4928,N_4704,N_4732);
nor U4929 (N_4929,N_4712,N_4672);
and U4930 (N_4930,N_4629,N_4774);
or U4931 (N_4931,N_4709,N_4756);
nor U4932 (N_4932,N_4749,N_4659);
and U4933 (N_4933,N_4746,N_4684);
and U4934 (N_4934,N_4683,N_4786);
nor U4935 (N_4935,N_4672,N_4749);
or U4936 (N_4936,N_4761,N_4619);
and U4937 (N_4937,N_4748,N_4736);
or U4938 (N_4938,N_4779,N_4641);
and U4939 (N_4939,N_4767,N_4733);
xnor U4940 (N_4940,N_4631,N_4799);
nor U4941 (N_4941,N_4753,N_4669);
or U4942 (N_4942,N_4796,N_4700);
or U4943 (N_4943,N_4786,N_4746);
and U4944 (N_4944,N_4670,N_4798);
nand U4945 (N_4945,N_4793,N_4753);
or U4946 (N_4946,N_4630,N_4705);
and U4947 (N_4947,N_4689,N_4747);
or U4948 (N_4948,N_4726,N_4727);
nor U4949 (N_4949,N_4610,N_4753);
and U4950 (N_4950,N_4685,N_4638);
xor U4951 (N_4951,N_4637,N_4600);
and U4952 (N_4952,N_4775,N_4677);
xnor U4953 (N_4953,N_4715,N_4746);
and U4954 (N_4954,N_4682,N_4645);
nand U4955 (N_4955,N_4751,N_4671);
and U4956 (N_4956,N_4763,N_4657);
or U4957 (N_4957,N_4600,N_4640);
and U4958 (N_4958,N_4796,N_4748);
nand U4959 (N_4959,N_4780,N_4754);
nor U4960 (N_4960,N_4773,N_4649);
nand U4961 (N_4961,N_4795,N_4765);
or U4962 (N_4962,N_4758,N_4754);
and U4963 (N_4963,N_4619,N_4764);
and U4964 (N_4964,N_4643,N_4685);
nor U4965 (N_4965,N_4637,N_4707);
nor U4966 (N_4966,N_4622,N_4642);
and U4967 (N_4967,N_4675,N_4688);
and U4968 (N_4968,N_4751,N_4605);
nor U4969 (N_4969,N_4636,N_4775);
nand U4970 (N_4970,N_4731,N_4774);
nor U4971 (N_4971,N_4700,N_4651);
or U4972 (N_4972,N_4619,N_4794);
or U4973 (N_4973,N_4716,N_4678);
nand U4974 (N_4974,N_4772,N_4715);
xnor U4975 (N_4975,N_4762,N_4768);
nor U4976 (N_4976,N_4614,N_4675);
and U4977 (N_4977,N_4634,N_4678);
and U4978 (N_4978,N_4641,N_4747);
nor U4979 (N_4979,N_4647,N_4785);
nand U4980 (N_4980,N_4722,N_4766);
nand U4981 (N_4981,N_4713,N_4732);
nand U4982 (N_4982,N_4727,N_4703);
nand U4983 (N_4983,N_4784,N_4694);
or U4984 (N_4984,N_4635,N_4723);
nand U4985 (N_4985,N_4710,N_4726);
or U4986 (N_4986,N_4683,N_4624);
or U4987 (N_4987,N_4618,N_4645);
and U4988 (N_4988,N_4730,N_4676);
nand U4989 (N_4989,N_4675,N_4686);
nor U4990 (N_4990,N_4638,N_4785);
or U4991 (N_4991,N_4744,N_4739);
or U4992 (N_4992,N_4721,N_4786);
or U4993 (N_4993,N_4737,N_4715);
nor U4994 (N_4994,N_4761,N_4739);
nand U4995 (N_4995,N_4709,N_4736);
nand U4996 (N_4996,N_4672,N_4711);
nor U4997 (N_4997,N_4623,N_4646);
and U4998 (N_4998,N_4762,N_4728);
nand U4999 (N_4999,N_4679,N_4663);
and U5000 (N_5000,N_4838,N_4907);
or U5001 (N_5001,N_4901,N_4833);
nand U5002 (N_5002,N_4834,N_4837);
nand U5003 (N_5003,N_4884,N_4828);
nor U5004 (N_5004,N_4869,N_4946);
nand U5005 (N_5005,N_4836,N_4807);
and U5006 (N_5006,N_4870,N_4991);
nor U5007 (N_5007,N_4862,N_4928);
or U5008 (N_5008,N_4857,N_4958);
and U5009 (N_5009,N_4831,N_4894);
or U5010 (N_5010,N_4895,N_4873);
xor U5011 (N_5011,N_4978,N_4825);
xnor U5012 (N_5012,N_4867,N_4808);
nand U5013 (N_5013,N_4802,N_4965);
nor U5014 (N_5014,N_4801,N_4902);
or U5015 (N_5015,N_4812,N_4944);
and U5016 (N_5016,N_4961,N_4875);
nand U5017 (N_5017,N_4864,N_4940);
and U5018 (N_5018,N_4856,N_4863);
nor U5019 (N_5019,N_4948,N_4954);
nand U5020 (N_5020,N_4922,N_4866);
and U5021 (N_5021,N_4981,N_4816);
nand U5022 (N_5022,N_4943,N_4906);
or U5023 (N_5023,N_4960,N_4950);
nor U5024 (N_5024,N_4971,N_4915);
or U5025 (N_5025,N_4832,N_4890);
nor U5026 (N_5026,N_4826,N_4967);
nand U5027 (N_5027,N_4865,N_4881);
nor U5028 (N_5028,N_4871,N_4973);
nand U5029 (N_5029,N_4849,N_4824);
and U5030 (N_5030,N_4880,N_4896);
nand U5031 (N_5031,N_4984,N_4927);
nor U5032 (N_5032,N_4882,N_4957);
or U5033 (N_5033,N_4912,N_4953);
and U5034 (N_5034,N_4850,N_4843);
nor U5035 (N_5035,N_4997,N_4874);
nor U5036 (N_5036,N_4989,N_4827);
or U5037 (N_5037,N_4941,N_4956);
nand U5038 (N_5038,N_4823,N_4848);
nand U5039 (N_5039,N_4962,N_4804);
and U5040 (N_5040,N_4844,N_4868);
nor U5041 (N_5041,N_4904,N_4966);
nand U5042 (N_5042,N_4969,N_4918);
nor U5043 (N_5043,N_4840,N_4921);
and U5044 (N_5044,N_4891,N_4911);
and U5045 (N_5045,N_4920,N_4820);
and U5046 (N_5046,N_4983,N_4919);
nor U5047 (N_5047,N_4932,N_4893);
xor U5048 (N_5048,N_4972,N_4990);
nand U5049 (N_5049,N_4859,N_4829);
or U5050 (N_5050,N_4817,N_4800);
or U5051 (N_5051,N_4963,N_4936);
nand U5052 (N_5052,N_4994,N_4970);
nand U5053 (N_5053,N_4839,N_4987);
and U5054 (N_5054,N_4916,N_4813);
and U5055 (N_5055,N_4803,N_4818);
nand U5056 (N_5056,N_4886,N_4988);
nor U5057 (N_5057,N_4934,N_4883);
nor U5058 (N_5058,N_4899,N_4986);
or U5059 (N_5059,N_4879,N_4974);
xnor U5060 (N_5060,N_4930,N_4842);
nand U5061 (N_5061,N_4900,N_4905);
and U5062 (N_5062,N_4992,N_4845);
and U5063 (N_5063,N_4908,N_4949);
nor U5064 (N_5064,N_4841,N_4854);
and U5065 (N_5065,N_4995,N_4830);
or U5066 (N_5066,N_4872,N_4805);
and U5067 (N_5067,N_4942,N_4924);
or U5068 (N_5068,N_4980,N_4858);
and U5069 (N_5069,N_4898,N_4996);
nand U5070 (N_5070,N_4855,N_4982);
and U5071 (N_5071,N_4917,N_4952);
nand U5072 (N_5072,N_4877,N_4810);
nor U5073 (N_5073,N_4892,N_4931);
and U5074 (N_5074,N_4819,N_4976);
nand U5075 (N_5075,N_4809,N_4897);
nand U5076 (N_5076,N_4852,N_4861);
or U5077 (N_5077,N_4853,N_4887);
nand U5078 (N_5078,N_4913,N_4888);
nand U5079 (N_5079,N_4933,N_4903);
nor U5080 (N_5080,N_4885,N_4945);
nand U5081 (N_5081,N_4977,N_4910);
and U5082 (N_5082,N_4964,N_4923);
nand U5083 (N_5083,N_4846,N_4998);
xor U5084 (N_5084,N_4993,N_4806);
or U5085 (N_5085,N_4925,N_4926);
nand U5086 (N_5086,N_4979,N_4947);
or U5087 (N_5087,N_4889,N_4959);
or U5088 (N_5088,N_4951,N_4860);
xor U5089 (N_5089,N_4835,N_4937);
nor U5090 (N_5090,N_4975,N_4878);
or U5091 (N_5091,N_4985,N_4876);
nand U5092 (N_5092,N_4822,N_4955);
nand U5093 (N_5093,N_4929,N_4815);
nand U5094 (N_5094,N_4935,N_4914);
nor U5095 (N_5095,N_4939,N_4938);
or U5096 (N_5096,N_4847,N_4814);
and U5097 (N_5097,N_4811,N_4821);
nor U5098 (N_5098,N_4999,N_4909);
nor U5099 (N_5099,N_4968,N_4851);
and U5100 (N_5100,N_4829,N_4908);
xor U5101 (N_5101,N_4894,N_4968);
nor U5102 (N_5102,N_4999,N_4816);
and U5103 (N_5103,N_4893,N_4814);
or U5104 (N_5104,N_4913,N_4993);
and U5105 (N_5105,N_4941,N_4978);
nor U5106 (N_5106,N_4855,N_4960);
nor U5107 (N_5107,N_4834,N_4895);
and U5108 (N_5108,N_4965,N_4817);
and U5109 (N_5109,N_4865,N_4836);
or U5110 (N_5110,N_4926,N_4942);
nand U5111 (N_5111,N_4899,N_4838);
and U5112 (N_5112,N_4996,N_4945);
and U5113 (N_5113,N_4880,N_4872);
nand U5114 (N_5114,N_4829,N_4850);
xnor U5115 (N_5115,N_4983,N_4985);
nand U5116 (N_5116,N_4946,N_4857);
nand U5117 (N_5117,N_4968,N_4905);
xor U5118 (N_5118,N_4946,N_4894);
nor U5119 (N_5119,N_4872,N_4946);
or U5120 (N_5120,N_4816,N_4870);
nor U5121 (N_5121,N_4982,N_4858);
or U5122 (N_5122,N_4909,N_4861);
nand U5123 (N_5123,N_4999,N_4943);
nand U5124 (N_5124,N_4881,N_4973);
and U5125 (N_5125,N_4909,N_4934);
nor U5126 (N_5126,N_4825,N_4977);
and U5127 (N_5127,N_4888,N_4959);
or U5128 (N_5128,N_4920,N_4858);
nand U5129 (N_5129,N_4885,N_4918);
nand U5130 (N_5130,N_4902,N_4939);
and U5131 (N_5131,N_4802,N_4962);
or U5132 (N_5132,N_4834,N_4826);
and U5133 (N_5133,N_4864,N_4900);
nor U5134 (N_5134,N_4963,N_4953);
or U5135 (N_5135,N_4950,N_4932);
nand U5136 (N_5136,N_4807,N_4943);
nor U5137 (N_5137,N_4967,N_4922);
nor U5138 (N_5138,N_4977,N_4959);
nand U5139 (N_5139,N_4971,N_4898);
xor U5140 (N_5140,N_4862,N_4902);
or U5141 (N_5141,N_4983,N_4927);
nor U5142 (N_5142,N_4910,N_4865);
nand U5143 (N_5143,N_4934,N_4967);
nand U5144 (N_5144,N_4931,N_4860);
or U5145 (N_5145,N_4810,N_4881);
and U5146 (N_5146,N_4846,N_4997);
nor U5147 (N_5147,N_4880,N_4902);
and U5148 (N_5148,N_4816,N_4992);
nor U5149 (N_5149,N_4960,N_4826);
nand U5150 (N_5150,N_4993,N_4896);
nor U5151 (N_5151,N_4852,N_4992);
and U5152 (N_5152,N_4896,N_4821);
and U5153 (N_5153,N_4938,N_4980);
or U5154 (N_5154,N_4934,N_4941);
and U5155 (N_5155,N_4831,N_4916);
or U5156 (N_5156,N_4838,N_4956);
nor U5157 (N_5157,N_4834,N_4829);
nor U5158 (N_5158,N_4864,N_4856);
nand U5159 (N_5159,N_4968,N_4867);
nand U5160 (N_5160,N_4926,N_4944);
or U5161 (N_5161,N_4869,N_4915);
or U5162 (N_5162,N_4892,N_4972);
nand U5163 (N_5163,N_4963,N_4912);
xor U5164 (N_5164,N_4824,N_4921);
nor U5165 (N_5165,N_4900,N_4835);
nor U5166 (N_5166,N_4941,N_4910);
nor U5167 (N_5167,N_4825,N_4994);
and U5168 (N_5168,N_4878,N_4994);
and U5169 (N_5169,N_4880,N_4851);
or U5170 (N_5170,N_4820,N_4871);
xnor U5171 (N_5171,N_4938,N_4949);
or U5172 (N_5172,N_4939,N_4952);
nor U5173 (N_5173,N_4976,N_4981);
or U5174 (N_5174,N_4893,N_4861);
nand U5175 (N_5175,N_4978,N_4880);
and U5176 (N_5176,N_4878,N_4897);
and U5177 (N_5177,N_4986,N_4979);
and U5178 (N_5178,N_4962,N_4966);
nand U5179 (N_5179,N_4954,N_4978);
nor U5180 (N_5180,N_4812,N_4931);
nand U5181 (N_5181,N_4985,N_4891);
nand U5182 (N_5182,N_4875,N_4972);
and U5183 (N_5183,N_4829,N_4819);
and U5184 (N_5184,N_4853,N_4999);
nor U5185 (N_5185,N_4901,N_4836);
nand U5186 (N_5186,N_4893,N_4941);
and U5187 (N_5187,N_4965,N_4917);
and U5188 (N_5188,N_4952,N_4897);
or U5189 (N_5189,N_4957,N_4846);
or U5190 (N_5190,N_4884,N_4945);
or U5191 (N_5191,N_4894,N_4986);
nor U5192 (N_5192,N_4873,N_4812);
nor U5193 (N_5193,N_4858,N_4933);
nor U5194 (N_5194,N_4925,N_4924);
nand U5195 (N_5195,N_4892,N_4953);
or U5196 (N_5196,N_4969,N_4806);
xor U5197 (N_5197,N_4951,N_4952);
or U5198 (N_5198,N_4857,N_4996);
nand U5199 (N_5199,N_4958,N_4810);
nor U5200 (N_5200,N_5126,N_5131);
and U5201 (N_5201,N_5146,N_5023);
nor U5202 (N_5202,N_5034,N_5123);
and U5203 (N_5203,N_5028,N_5091);
or U5204 (N_5204,N_5059,N_5120);
nand U5205 (N_5205,N_5141,N_5022);
or U5206 (N_5206,N_5187,N_5020);
or U5207 (N_5207,N_5021,N_5108);
or U5208 (N_5208,N_5064,N_5030);
nor U5209 (N_5209,N_5157,N_5144);
and U5210 (N_5210,N_5097,N_5179);
and U5211 (N_5211,N_5182,N_5162);
xor U5212 (N_5212,N_5183,N_5006);
xnor U5213 (N_5213,N_5140,N_5049);
or U5214 (N_5214,N_5009,N_5103);
and U5215 (N_5215,N_5054,N_5180);
nor U5216 (N_5216,N_5137,N_5010);
and U5217 (N_5217,N_5192,N_5112);
or U5218 (N_5218,N_5015,N_5053);
or U5219 (N_5219,N_5104,N_5124);
xnor U5220 (N_5220,N_5067,N_5148);
xor U5221 (N_5221,N_5173,N_5159);
and U5222 (N_5222,N_5114,N_5004);
or U5223 (N_5223,N_5078,N_5033);
nor U5224 (N_5224,N_5111,N_5161);
and U5225 (N_5225,N_5136,N_5106);
nor U5226 (N_5226,N_5077,N_5181);
nor U5227 (N_5227,N_5164,N_5002);
and U5228 (N_5228,N_5129,N_5011);
nand U5229 (N_5229,N_5100,N_5107);
nor U5230 (N_5230,N_5168,N_5113);
or U5231 (N_5231,N_5169,N_5166);
nor U5232 (N_5232,N_5068,N_5063);
or U5233 (N_5233,N_5007,N_5039);
nor U5234 (N_5234,N_5139,N_5081);
nand U5235 (N_5235,N_5152,N_5095);
nor U5236 (N_5236,N_5174,N_5000);
xnor U5237 (N_5237,N_5038,N_5134);
nor U5238 (N_5238,N_5153,N_5024);
or U5239 (N_5239,N_5035,N_5073);
nand U5240 (N_5240,N_5075,N_5065);
nand U5241 (N_5241,N_5090,N_5080);
and U5242 (N_5242,N_5089,N_5118);
and U5243 (N_5243,N_5191,N_5051);
nor U5244 (N_5244,N_5197,N_5199);
and U5245 (N_5245,N_5184,N_5158);
nor U5246 (N_5246,N_5071,N_5074);
nor U5247 (N_5247,N_5047,N_5060);
nand U5248 (N_5248,N_5092,N_5175);
nand U5249 (N_5249,N_5147,N_5070);
nand U5250 (N_5250,N_5149,N_5142);
or U5251 (N_5251,N_5003,N_5172);
and U5252 (N_5252,N_5177,N_5026);
nor U5253 (N_5253,N_5138,N_5195);
nor U5254 (N_5254,N_5117,N_5013);
nand U5255 (N_5255,N_5031,N_5101);
or U5256 (N_5256,N_5109,N_5072);
nand U5257 (N_5257,N_5079,N_5167);
nor U5258 (N_5258,N_5189,N_5046);
and U5259 (N_5259,N_5155,N_5151);
or U5260 (N_5260,N_5188,N_5066);
or U5261 (N_5261,N_5105,N_5084);
or U5262 (N_5262,N_5096,N_5041);
or U5263 (N_5263,N_5086,N_5121);
or U5264 (N_5264,N_5050,N_5122);
or U5265 (N_5265,N_5127,N_5132);
and U5266 (N_5266,N_5012,N_5160);
or U5267 (N_5267,N_5193,N_5008);
and U5268 (N_5268,N_5061,N_5156);
nand U5269 (N_5269,N_5019,N_5130);
nand U5270 (N_5270,N_5069,N_5027);
and U5271 (N_5271,N_5185,N_5119);
and U5272 (N_5272,N_5171,N_5163);
nand U5273 (N_5273,N_5099,N_5088);
xnor U5274 (N_5274,N_5044,N_5102);
nor U5275 (N_5275,N_5042,N_5043);
nand U5276 (N_5276,N_5085,N_5036);
nor U5277 (N_5277,N_5098,N_5116);
or U5278 (N_5278,N_5025,N_5040);
xnor U5279 (N_5279,N_5115,N_5055);
nor U5280 (N_5280,N_5186,N_5058);
nand U5281 (N_5281,N_5062,N_5093);
and U5282 (N_5282,N_5110,N_5128);
nor U5283 (N_5283,N_5029,N_5194);
and U5284 (N_5284,N_5176,N_5150);
and U5285 (N_5285,N_5190,N_5001);
or U5286 (N_5286,N_5145,N_5143);
and U5287 (N_5287,N_5052,N_5125);
xnor U5288 (N_5288,N_5170,N_5083);
nor U5289 (N_5289,N_5057,N_5017);
nor U5290 (N_5290,N_5045,N_5094);
nor U5291 (N_5291,N_5076,N_5018);
and U5292 (N_5292,N_5005,N_5014);
or U5293 (N_5293,N_5016,N_5082);
nand U5294 (N_5294,N_5178,N_5135);
nand U5295 (N_5295,N_5048,N_5056);
and U5296 (N_5296,N_5037,N_5196);
or U5297 (N_5297,N_5032,N_5133);
nor U5298 (N_5298,N_5165,N_5087);
and U5299 (N_5299,N_5198,N_5154);
nand U5300 (N_5300,N_5019,N_5015);
or U5301 (N_5301,N_5115,N_5037);
nand U5302 (N_5302,N_5004,N_5186);
nand U5303 (N_5303,N_5047,N_5027);
and U5304 (N_5304,N_5192,N_5053);
or U5305 (N_5305,N_5115,N_5174);
and U5306 (N_5306,N_5131,N_5055);
and U5307 (N_5307,N_5071,N_5185);
nand U5308 (N_5308,N_5011,N_5076);
nand U5309 (N_5309,N_5109,N_5028);
xnor U5310 (N_5310,N_5072,N_5195);
and U5311 (N_5311,N_5079,N_5120);
nor U5312 (N_5312,N_5196,N_5035);
nor U5313 (N_5313,N_5175,N_5131);
nand U5314 (N_5314,N_5086,N_5079);
nand U5315 (N_5315,N_5029,N_5073);
and U5316 (N_5316,N_5133,N_5129);
or U5317 (N_5317,N_5015,N_5118);
and U5318 (N_5318,N_5016,N_5027);
or U5319 (N_5319,N_5197,N_5181);
nor U5320 (N_5320,N_5177,N_5156);
nor U5321 (N_5321,N_5110,N_5065);
nor U5322 (N_5322,N_5116,N_5120);
nand U5323 (N_5323,N_5094,N_5136);
nand U5324 (N_5324,N_5100,N_5050);
and U5325 (N_5325,N_5039,N_5016);
and U5326 (N_5326,N_5136,N_5156);
nor U5327 (N_5327,N_5140,N_5107);
or U5328 (N_5328,N_5000,N_5194);
nor U5329 (N_5329,N_5191,N_5019);
or U5330 (N_5330,N_5065,N_5059);
and U5331 (N_5331,N_5152,N_5146);
xnor U5332 (N_5332,N_5093,N_5124);
or U5333 (N_5333,N_5066,N_5160);
nor U5334 (N_5334,N_5159,N_5068);
xnor U5335 (N_5335,N_5119,N_5090);
or U5336 (N_5336,N_5052,N_5002);
nor U5337 (N_5337,N_5024,N_5135);
and U5338 (N_5338,N_5164,N_5064);
or U5339 (N_5339,N_5175,N_5196);
and U5340 (N_5340,N_5177,N_5091);
or U5341 (N_5341,N_5198,N_5152);
and U5342 (N_5342,N_5146,N_5038);
nand U5343 (N_5343,N_5025,N_5024);
and U5344 (N_5344,N_5006,N_5114);
or U5345 (N_5345,N_5041,N_5185);
and U5346 (N_5346,N_5156,N_5128);
and U5347 (N_5347,N_5126,N_5057);
or U5348 (N_5348,N_5184,N_5005);
and U5349 (N_5349,N_5123,N_5012);
or U5350 (N_5350,N_5126,N_5017);
nand U5351 (N_5351,N_5005,N_5189);
nor U5352 (N_5352,N_5158,N_5166);
nand U5353 (N_5353,N_5099,N_5086);
or U5354 (N_5354,N_5073,N_5199);
nor U5355 (N_5355,N_5167,N_5146);
nand U5356 (N_5356,N_5028,N_5103);
nor U5357 (N_5357,N_5074,N_5028);
xor U5358 (N_5358,N_5055,N_5178);
nor U5359 (N_5359,N_5040,N_5003);
or U5360 (N_5360,N_5022,N_5050);
nor U5361 (N_5361,N_5121,N_5128);
or U5362 (N_5362,N_5065,N_5061);
xor U5363 (N_5363,N_5121,N_5129);
nand U5364 (N_5364,N_5058,N_5088);
and U5365 (N_5365,N_5023,N_5148);
and U5366 (N_5366,N_5107,N_5111);
and U5367 (N_5367,N_5188,N_5101);
xnor U5368 (N_5368,N_5072,N_5089);
or U5369 (N_5369,N_5051,N_5179);
xnor U5370 (N_5370,N_5185,N_5001);
and U5371 (N_5371,N_5144,N_5076);
nand U5372 (N_5372,N_5024,N_5119);
nand U5373 (N_5373,N_5017,N_5044);
xnor U5374 (N_5374,N_5029,N_5172);
nor U5375 (N_5375,N_5149,N_5135);
xor U5376 (N_5376,N_5026,N_5142);
nor U5377 (N_5377,N_5165,N_5012);
and U5378 (N_5378,N_5009,N_5194);
and U5379 (N_5379,N_5158,N_5182);
or U5380 (N_5380,N_5077,N_5080);
and U5381 (N_5381,N_5005,N_5115);
nand U5382 (N_5382,N_5078,N_5060);
xor U5383 (N_5383,N_5184,N_5157);
nor U5384 (N_5384,N_5149,N_5077);
nand U5385 (N_5385,N_5070,N_5166);
xnor U5386 (N_5386,N_5005,N_5045);
nand U5387 (N_5387,N_5170,N_5090);
nor U5388 (N_5388,N_5095,N_5019);
and U5389 (N_5389,N_5016,N_5122);
or U5390 (N_5390,N_5176,N_5190);
xnor U5391 (N_5391,N_5094,N_5184);
xor U5392 (N_5392,N_5038,N_5091);
xnor U5393 (N_5393,N_5007,N_5151);
or U5394 (N_5394,N_5137,N_5075);
nand U5395 (N_5395,N_5024,N_5139);
or U5396 (N_5396,N_5098,N_5052);
and U5397 (N_5397,N_5007,N_5107);
and U5398 (N_5398,N_5089,N_5027);
and U5399 (N_5399,N_5053,N_5167);
or U5400 (N_5400,N_5378,N_5310);
nor U5401 (N_5401,N_5263,N_5324);
nand U5402 (N_5402,N_5228,N_5334);
xnor U5403 (N_5403,N_5358,N_5208);
nand U5404 (N_5404,N_5346,N_5318);
and U5405 (N_5405,N_5319,N_5306);
and U5406 (N_5406,N_5385,N_5317);
nand U5407 (N_5407,N_5394,N_5256);
nor U5408 (N_5408,N_5279,N_5372);
nor U5409 (N_5409,N_5257,N_5274);
nand U5410 (N_5410,N_5227,N_5252);
nand U5411 (N_5411,N_5245,N_5261);
nor U5412 (N_5412,N_5202,N_5260);
xnor U5413 (N_5413,N_5244,N_5376);
and U5414 (N_5414,N_5299,N_5212);
nand U5415 (N_5415,N_5314,N_5297);
nor U5416 (N_5416,N_5383,N_5399);
nor U5417 (N_5417,N_5219,N_5335);
or U5418 (N_5418,N_5389,N_5226);
and U5419 (N_5419,N_5368,N_5359);
and U5420 (N_5420,N_5396,N_5238);
and U5421 (N_5421,N_5221,N_5266);
and U5422 (N_5422,N_5271,N_5330);
xor U5423 (N_5423,N_5286,N_5200);
and U5424 (N_5424,N_5269,N_5287);
and U5425 (N_5425,N_5291,N_5251);
xnor U5426 (N_5426,N_5360,N_5354);
nor U5427 (N_5427,N_5265,N_5386);
nand U5428 (N_5428,N_5384,N_5281);
or U5429 (N_5429,N_5273,N_5237);
nor U5430 (N_5430,N_5230,N_5204);
and U5431 (N_5431,N_5391,N_5272);
nand U5432 (N_5432,N_5233,N_5249);
xnor U5433 (N_5433,N_5264,N_5320);
nor U5434 (N_5434,N_5338,N_5343);
nand U5435 (N_5435,N_5213,N_5222);
nor U5436 (N_5436,N_5243,N_5203);
xnor U5437 (N_5437,N_5303,N_5387);
and U5438 (N_5438,N_5250,N_5267);
or U5439 (N_5439,N_5296,N_5283);
nor U5440 (N_5440,N_5277,N_5214);
or U5441 (N_5441,N_5300,N_5248);
nand U5442 (N_5442,N_5325,N_5367);
nor U5443 (N_5443,N_5328,N_5270);
nor U5444 (N_5444,N_5201,N_5357);
nor U5445 (N_5445,N_5290,N_5355);
nor U5446 (N_5446,N_5235,N_5315);
nor U5447 (N_5447,N_5216,N_5308);
or U5448 (N_5448,N_5371,N_5347);
nand U5449 (N_5449,N_5206,N_5345);
or U5450 (N_5450,N_5293,N_5356);
or U5451 (N_5451,N_5207,N_5285);
and U5452 (N_5452,N_5327,N_5395);
nor U5453 (N_5453,N_5381,N_5302);
nor U5454 (N_5454,N_5301,N_5333);
xnor U5455 (N_5455,N_5232,N_5284);
and U5456 (N_5456,N_5253,N_5366);
xor U5457 (N_5457,N_5331,N_5215);
or U5458 (N_5458,N_5305,N_5382);
and U5459 (N_5459,N_5350,N_5223);
xor U5460 (N_5460,N_5220,N_5362);
nand U5461 (N_5461,N_5259,N_5336);
and U5462 (N_5462,N_5210,N_5344);
nand U5463 (N_5463,N_5211,N_5316);
nor U5464 (N_5464,N_5322,N_5311);
and U5465 (N_5465,N_5294,N_5236);
nand U5466 (N_5466,N_5292,N_5280);
nand U5467 (N_5467,N_5289,N_5352);
nand U5468 (N_5468,N_5307,N_5349);
or U5469 (N_5469,N_5329,N_5370);
nand U5470 (N_5470,N_5276,N_5351);
nor U5471 (N_5471,N_5240,N_5217);
nor U5472 (N_5472,N_5390,N_5275);
or U5473 (N_5473,N_5321,N_5313);
nand U5474 (N_5474,N_5392,N_5205);
or U5475 (N_5475,N_5304,N_5298);
and U5476 (N_5476,N_5229,N_5282);
nor U5477 (N_5477,N_5241,N_5397);
nand U5478 (N_5478,N_5247,N_5231);
and U5479 (N_5479,N_5369,N_5309);
or U5480 (N_5480,N_5262,N_5239);
nor U5481 (N_5481,N_5364,N_5209);
and U5482 (N_5482,N_5348,N_5337);
nand U5483 (N_5483,N_5340,N_5288);
xor U5484 (N_5484,N_5398,N_5326);
xnor U5485 (N_5485,N_5339,N_5295);
or U5486 (N_5486,N_5246,N_5379);
nor U5487 (N_5487,N_5225,N_5374);
and U5488 (N_5488,N_5363,N_5234);
and U5489 (N_5489,N_5361,N_5254);
nor U5490 (N_5490,N_5258,N_5242);
and U5491 (N_5491,N_5268,N_5278);
and U5492 (N_5492,N_5375,N_5353);
and U5493 (N_5493,N_5323,N_5393);
nor U5494 (N_5494,N_5224,N_5341);
or U5495 (N_5495,N_5365,N_5342);
and U5496 (N_5496,N_5380,N_5377);
and U5497 (N_5497,N_5332,N_5218);
nand U5498 (N_5498,N_5255,N_5388);
and U5499 (N_5499,N_5312,N_5373);
nand U5500 (N_5500,N_5340,N_5244);
and U5501 (N_5501,N_5238,N_5291);
xor U5502 (N_5502,N_5213,N_5389);
xnor U5503 (N_5503,N_5312,N_5241);
nor U5504 (N_5504,N_5377,N_5259);
or U5505 (N_5505,N_5245,N_5383);
and U5506 (N_5506,N_5225,N_5264);
nor U5507 (N_5507,N_5213,N_5284);
nand U5508 (N_5508,N_5284,N_5311);
nor U5509 (N_5509,N_5372,N_5325);
and U5510 (N_5510,N_5242,N_5370);
or U5511 (N_5511,N_5308,N_5322);
or U5512 (N_5512,N_5211,N_5291);
nand U5513 (N_5513,N_5254,N_5384);
and U5514 (N_5514,N_5229,N_5343);
nand U5515 (N_5515,N_5342,N_5364);
xor U5516 (N_5516,N_5336,N_5377);
and U5517 (N_5517,N_5288,N_5210);
nand U5518 (N_5518,N_5315,N_5353);
or U5519 (N_5519,N_5356,N_5304);
and U5520 (N_5520,N_5242,N_5327);
nand U5521 (N_5521,N_5245,N_5235);
nand U5522 (N_5522,N_5251,N_5250);
nand U5523 (N_5523,N_5379,N_5215);
nand U5524 (N_5524,N_5324,N_5342);
or U5525 (N_5525,N_5225,N_5230);
and U5526 (N_5526,N_5235,N_5313);
nand U5527 (N_5527,N_5247,N_5348);
nor U5528 (N_5528,N_5236,N_5343);
and U5529 (N_5529,N_5316,N_5368);
nand U5530 (N_5530,N_5334,N_5263);
and U5531 (N_5531,N_5275,N_5370);
xnor U5532 (N_5532,N_5241,N_5239);
and U5533 (N_5533,N_5355,N_5229);
nor U5534 (N_5534,N_5385,N_5382);
and U5535 (N_5535,N_5237,N_5319);
and U5536 (N_5536,N_5326,N_5352);
nor U5537 (N_5537,N_5201,N_5245);
nor U5538 (N_5538,N_5324,N_5396);
or U5539 (N_5539,N_5262,N_5266);
nand U5540 (N_5540,N_5363,N_5382);
xor U5541 (N_5541,N_5393,N_5287);
nand U5542 (N_5542,N_5242,N_5332);
nand U5543 (N_5543,N_5343,N_5349);
nand U5544 (N_5544,N_5327,N_5243);
xnor U5545 (N_5545,N_5300,N_5352);
or U5546 (N_5546,N_5330,N_5237);
nor U5547 (N_5547,N_5315,N_5286);
or U5548 (N_5548,N_5346,N_5323);
or U5549 (N_5549,N_5308,N_5315);
nor U5550 (N_5550,N_5362,N_5218);
nor U5551 (N_5551,N_5381,N_5205);
nor U5552 (N_5552,N_5218,N_5246);
nor U5553 (N_5553,N_5367,N_5238);
nand U5554 (N_5554,N_5345,N_5223);
and U5555 (N_5555,N_5322,N_5223);
nor U5556 (N_5556,N_5218,N_5299);
and U5557 (N_5557,N_5336,N_5376);
nand U5558 (N_5558,N_5229,N_5208);
and U5559 (N_5559,N_5338,N_5346);
or U5560 (N_5560,N_5212,N_5358);
and U5561 (N_5561,N_5235,N_5349);
or U5562 (N_5562,N_5305,N_5346);
nand U5563 (N_5563,N_5310,N_5265);
nand U5564 (N_5564,N_5352,N_5373);
nand U5565 (N_5565,N_5288,N_5314);
nand U5566 (N_5566,N_5204,N_5258);
nand U5567 (N_5567,N_5358,N_5247);
nand U5568 (N_5568,N_5309,N_5399);
and U5569 (N_5569,N_5240,N_5366);
nor U5570 (N_5570,N_5202,N_5262);
nor U5571 (N_5571,N_5237,N_5325);
nand U5572 (N_5572,N_5201,N_5378);
and U5573 (N_5573,N_5385,N_5234);
and U5574 (N_5574,N_5268,N_5274);
nand U5575 (N_5575,N_5236,N_5314);
xor U5576 (N_5576,N_5356,N_5223);
nand U5577 (N_5577,N_5335,N_5370);
or U5578 (N_5578,N_5305,N_5249);
and U5579 (N_5579,N_5254,N_5237);
and U5580 (N_5580,N_5246,N_5224);
and U5581 (N_5581,N_5306,N_5393);
nand U5582 (N_5582,N_5230,N_5224);
and U5583 (N_5583,N_5225,N_5328);
nor U5584 (N_5584,N_5337,N_5311);
and U5585 (N_5585,N_5256,N_5311);
or U5586 (N_5586,N_5231,N_5358);
nor U5587 (N_5587,N_5255,N_5353);
or U5588 (N_5588,N_5268,N_5229);
nor U5589 (N_5589,N_5355,N_5230);
and U5590 (N_5590,N_5233,N_5220);
nor U5591 (N_5591,N_5374,N_5389);
nand U5592 (N_5592,N_5382,N_5319);
or U5593 (N_5593,N_5282,N_5226);
nand U5594 (N_5594,N_5376,N_5301);
or U5595 (N_5595,N_5205,N_5328);
nand U5596 (N_5596,N_5334,N_5397);
nand U5597 (N_5597,N_5382,N_5351);
nor U5598 (N_5598,N_5327,N_5293);
nand U5599 (N_5599,N_5246,N_5289);
or U5600 (N_5600,N_5519,N_5528);
and U5601 (N_5601,N_5540,N_5598);
xnor U5602 (N_5602,N_5555,N_5548);
or U5603 (N_5603,N_5413,N_5465);
nor U5604 (N_5604,N_5573,N_5403);
and U5605 (N_5605,N_5591,N_5406);
nor U5606 (N_5606,N_5411,N_5479);
and U5607 (N_5607,N_5524,N_5501);
or U5608 (N_5608,N_5466,N_5518);
nor U5609 (N_5609,N_5570,N_5482);
or U5610 (N_5610,N_5410,N_5564);
nor U5611 (N_5611,N_5486,N_5575);
nor U5612 (N_5612,N_5450,N_5453);
or U5613 (N_5613,N_5594,N_5496);
nor U5614 (N_5614,N_5522,N_5526);
or U5615 (N_5615,N_5455,N_5543);
nand U5616 (N_5616,N_5539,N_5529);
or U5617 (N_5617,N_5430,N_5534);
and U5618 (N_5618,N_5449,N_5472);
nand U5619 (N_5619,N_5506,N_5491);
nand U5620 (N_5620,N_5417,N_5596);
or U5621 (N_5621,N_5474,N_5437);
nand U5622 (N_5622,N_5525,N_5494);
nor U5623 (N_5623,N_5435,N_5500);
and U5624 (N_5624,N_5504,N_5419);
or U5625 (N_5625,N_5442,N_5426);
xor U5626 (N_5626,N_5432,N_5438);
and U5627 (N_5627,N_5448,N_5568);
nand U5628 (N_5628,N_5447,N_5582);
xnor U5629 (N_5629,N_5443,N_5559);
or U5630 (N_5630,N_5467,N_5561);
nand U5631 (N_5631,N_5597,N_5457);
nor U5632 (N_5632,N_5489,N_5505);
nand U5633 (N_5633,N_5495,N_5477);
or U5634 (N_5634,N_5584,N_5521);
xor U5635 (N_5635,N_5511,N_5587);
nor U5636 (N_5636,N_5512,N_5508);
and U5637 (N_5637,N_5574,N_5478);
and U5638 (N_5638,N_5420,N_5459);
and U5639 (N_5639,N_5502,N_5488);
nor U5640 (N_5640,N_5415,N_5421);
and U5641 (N_5641,N_5552,N_5473);
xnor U5642 (N_5642,N_5405,N_5412);
nor U5643 (N_5643,N_5468,N_5400);
xor U5644 (N_5644,N_5401,N_5439);
nor U5645 (N_5645,N_5445,N_5461);
nand U5646 (N_5646,N_5527,N_5414);
nand U5647 (N_5647,N_5546,N_5550);
or U5648 (N_5648,N_5560,N_5520);
or U5649 (N_5649,N_5458,N_5424);
nand U5650 (N_5650,N_5441,N_5531);
and U5651 (N_5651,N_5499,N_5446);
or U5652 (N_5652,N_5485,N_5563);
nand U5653 (N_5653,N_5576,N_5431);
xnor U5654 (N_5654,N_5422,N_5566);
and U5655 (N_5655,N_5554,N_5483);
or U5656 (N_5656,N_5593,N_5451);
nand U5657 (N_5657,N_5536,N_5452);
nor U5658 (N_5658,N_5463,N_5464);
nand U5659 (N_5659,N_5510,N_5599);
nand U5660 (N_5660,N_5416,N_5497);
nand U5661 (N_5661,N_5578,N_5462);
nand U5662 (N_5662,N_5513,N_5481);
and U5663 (N_5663,N_5558,N_5588);
or U5664 (N_5664,N_5409,N_5577);
or U5665 (N_5665,N_5565,N_5579);
nor U5666 (N_5666,N_5592,N_5538);
nand U5667 (N_5667,N_5492,N_5509);
and U5668 (N_5668,N_5476,N_5583);
xor U5669 (N_5669,N_5470,N_5586);
and U5670 (N_5670,N_5590,N_5517);
or U5671 (N_5671,N_5490,N_5557);
and U5672 (N_5672,N_5595,N_5544);
or U5673 (N_5673,N_5541,N_5454);
nand U5674 (N_5674,N_5456,N_5475);
nand U5675 (N_5675,N_5427,N_5562);
nor U5676 (N_5676,N_5533,N_5537);
and U5677 (N_5677,N_5440,N_5580);
or U5678 (N_5678,N_5581,N_5551);
nor U5679 (N_5679,N_5444,N_5542);
and U5680 (N_5680,N_5407,N_5516);
nor U5681 (N_5681,N_5535,N_5545);
nor U5682 (N_5682,N_5434,N_5436);
or U5683 (N_5683,N_5469,N_5423);
or U5684 (N_5684,N_5471,N_5589);
nand U5685 (N_5685,N_5507,N_5514);
nor U5686 (N_5686,N_5460,N_5480);
nand U5687 (N_5687,N_5532,N_5515);
nand U5688 (N_5688,N_5569,N_5553);
or U5689 (N_5689,N_5418,N_5567);
and U5690 (N_5690,N_5433,N_5493);
nor U5691 (N_5691,N_5547,N_5503);
or U5692 (N_5692,N_5572,N_5429);
nor U5693 (N_5693,N_5549,N_5425);
nand U5694 (N_5694,N_5556,N_5408);
xnor U5695 (N_5695,N_5402,N_5487);
nand U5696 (N_5696,N_5484,N_5428);
and U5697 (N_5697,N_5571,N_5498);
nor U5698 (N_5698,N_5404,N_5530);
nor U5699 (N_5699,N_5585,N_5523);
nor U5700 (N_5700,N_5531,N_5502);
or U5701 (N_5701,N_5423,N_5471);
nand U5702 (N_5702,N_5535,N_5408);
nor U5703 (N_5703,N_5469,N_5580);
nand U5704 (N_5704,N_5432,N_5405);
nor U5705 (N_5705,N_5463,N_5561);
or U5706 (N_5706,N_5411,N_5570);
xor U5707 (N_5707,N_5555,N_5402);
and U5708 (N_5708,N_5579,N_5420);
or U5709 (N_5709,N_5404,N_5525);
nand U5710 (N_5710,N_5454,N_5473);
xor U5711 (N_5711,N_5450,N_5441);
xor U5712 (N_5712,N_5510,N_5475);
xnor U5713 (N_5713,N_5453,N_5498);
nand U5714 (N_5714,N_5467,N_5422);
nand U5715 (N_5715,N_5451,N_5556);
and U5716 (N_5716,N_5431,N_5489);
nor U5717 (N_5717,N_5438,N_5404);
nand U5718 (N_5718,N_5480,N_5529);
nand U5719 (N_5719,N_5506,N_5588);
xnor U5720 (N_5720,N_5593,N_5439);
nor U5721 (N_5721,N_5409,N_5459);
xor U5722 (N_5722,N_5550,N_5412);
nor U5723 (N_5723,N_5436,N_5468);
nor U5724 (N_5724,N_5525,N_5548);
or U5725 (N_5725,N_5481,N_5436);
or U5726 (N_5726,N_5503,N_5566);
or U5727 (N_5727,N_5460,N_5520);
nor U5728 (N_5728,N_5572,N_5493);
nand U5729 (N_5729,N_5540,N_5599);
and U5730 (N_5730,N_5427,N_5431);
nand U5731 (N_5731,N_5435,N_5575);
xor U5732 (N_5732,N_5428,N_5575);
xnor U5733 (N_5733,N_5479,N_5476);
or U5734 (N_5734,N_5541,N_5506);
and U5735 (N_5735,N_5482,N_5501);
nand U5736 (N_5736,N_5591,N_5513);
and U5737 (N_5737,N_5558,N_5584);
nor U5738 (N_5738,N_5438,N_5588);
or U5739 (N_5739,N_5458,N_5580);
and U5740 (N_5740,N_5583,N_5586);
and U5741 (N_5741,N_5422,N_5521);
and U5742 (N_5742,N_5439,N_5533);
nand U5743 (N_5743,N_5502,N_5458);
and U5744 (N_5744,N_5437,N_5466);
nor U5745 (N_5745,N_5419,N_5596);
nand U5746 (N_5746,N_5556,N_5522);
nor U5747 (N_5747,N_5508,N_5513);
nor U5748 (N_5748,N_5548,N_5505);
and U5749 (N_5749,N_5411,N_5455);
and U5750 (N_5750,N_5576,N_5527);
nand U5751 (N_5751,N_5593,N_5578);
or U5752 (N_5752,N_5417,N_5535);
nand U5753 (N_5753,N_5486,N_5508);
and U5754 (N_5754,N_5552,N_5537);
nor U5755 (N_5755,N_5563,N_5575);
nand U5756 (N_5756,N_5481,N_5452);
and U5757 (N_5757,N_5413,N_5484);
nand U5758 (N_5758,N_5590,N_5532);
nor U5759 (N_5759,N_5549,N_5521);
and U5760 (N_5760,N_5493,N_5535);
nor U5761 (N_5761,N_5530,N_5571);
and U5762 (N_5762,N_5575,N_5431);
nand U5763 (N_5763,N_5449,N_5482);
and U5764 (N_5764,N_5479,N_5555);
nor U5765 (N_5765,N_5440,N_5593);
nor U5766 (N_5766,N_5559,N_5578);
nor U5767 (N_5767,N_5517,N_5549);
nor U5768 (N_5768,N_5551,N_5584);
or U5769 (N_5769,N_5433,N_5400);
or U5770 (N_5770,N_5428,N_5463);
and U5771 (N_5771,N_5425,N_5544);
or U5772 (N_5772,N_5458,N_5579);
nand U5773 (N_5773,N_5482,N_5457);
or U5774 (N_5774,N_5583,N_5491);
or U5775 (N_5775,N_5442,N_5522);
and U5776 (N_5776,N_5448,N_5454);
and U5777 (N_5777,N_5456,N_5531);
nor U5778 (N_5778,N_5435,N_5457);
xor U5779 (N_5779,N_5539,N_5495);
or U5780 (N_5780,N_5454,N_5422);
nand U5781 (N_5781,N_5554,N_5579);
nor U5782 (N_5782,N_5436,N_5510);
and U5783 (N_5783,N_5458,N_5426);
nor U5784 (N_5784,N_5491,N_5495);
nand U5785 (N_5785,N_5438,N_5528);
and U5786 (N_5786,N_5493,N_5479);
nand U5787 (N_5787,N_5401,N_5523);
nor U5788 (N_5788,N_5507,N_5460);
nand U5789 (N_5789,N_5401,N_5589);
or U5790 (N_5790,N_5523,N_5426);
or U5791 (N_5791,N_5477,N_5589);
xor U5792 (N_5792,N_5404,N_5594);
nor U5793 (N_5793,N_5469,N_5409);
nor U5794 (N_5794,N_5462,N_5591);
xor U5795 (N_5795,N_5505,N_5426);
nor U5796 (N_5796,N_5485,N_5500);
xor U5797 (N_5797,N_5585,N_5459);
and U5798 (N_5798,N_5582,N_5491);
or U5799 (N_5799,N_5582,N_5548);
or U5800 (N_5800,N_5606,N_5724);
nand U5801 (N_5801,N_5614,N_5652);
and U5802 (N_5802,N_5662,N_5741);
nand U5803 (N_5803,N_5717,N_5628);
or U5804 (N_5804,N_5657,N_5750);
nand U5805 (N_5805,N_5711,N_5648);
nor U5806 (N_5806,N_5611,N_5658);
and U5807 (N_5807,N_5646,N_5667);
and U5808 (N_5808,N_5642,N_5612);
nor U5809 (N_5809,N_5620,N_5719);
nand U5810 (N_5810,N_5782,N_5799);
or U5811 (N_5811,N_5731,N_5605);
and U5812 (N_5812,N_5604,N_5678);
or U5813 (N_5813,N_5708,N_5685);
and U5814 (N_5814,N_5749,N_5654);
nor U5815 (N_5815,N_5748,N_5755);
nand U5816 (N_5816,N_5687,N_5788);
nand U5817 (N_5817,N_5783,N_5772);
nor U5818 (N_5818,N_5745,N_5634);
nand U5819 (N_5819,N_5671,N_5784);
nand U5820 (N_5820,N_5762,N_5622);
or U5821 (N_5821,N_5680,N_5636);
and U5822 (N_5822,N_5760,N_5716);
nand U5823 (N_5823,N_5747,N_5689);
nand U5824 (N_5824,N_5608,N_5771);
and U5825 (N_5825,N_5681,N_5674);
nor U5826 (N_5826,N_5768,N_5744);
nand U5827 (N_5827,N_5617,N_5713);
or U5828 (N_5828,N_5682,N_5734);
or U5829 (N_5829,N_5781,N_5751);
nand U5830 (N_5830,N_5710,N_5673);
nor U5831 (N_5831,N_5797,N_5793);
or U5832 (N_5832,N_5633,N_5665);
nand U5833 (N_5833,N_5735,N_5676);
nor U5834 (N_5834,N_5679,N_5777);
or U5835 (N_5835,N_5677,N_5739);
or U5836 (N_5836,N_5603,N_5758);
and U5837 (N_5837,N_5703,N_5759);
xor U5838 (N_5838,N_5757,N_5718);
nand U5839 (N_5839,N_5726,N_5727);
nor U5840 (N_5840,N_5776,N_5767);
or U5841 (N_5841,N_5688,N_5638);
and U5842 (N_5842,N_5752,N_5789);
nand U5843 (N_5843,N_5743,N_5645);
and U5844 (N_5844,N_5664,N_5728);
or U5845 (N_5845,N_5641,N_5712);
and U5846 (N_5846,N_5644,N_5770);
nor U5847 (N_5847,N_5775,N_5692);
nand U5848 (N_5848,N_5729,N_5602);
nand U5849 (N_5849,N_5722,N_5730);
nor U5850 (N_5850,N_5631,N_5720);
or U5851 (N_5851,N_5696,N_5697);
nand U5852 (N_5852,N_5785,N_5740);
or U5853 (N_5853,N_5695,N_5701);
and U5854 (N_5854,N_5609,N_5610);
nor U5855 (N_5855,N_5668,N_5639);
or U5856 (N_5856,N_5663,N_5600);
or U5857 (N_5857,N_5723,N_5666);
or U5858 (N_5858,N_5669,N_5661);
or U5859 (N_5859,N_5798,N_5787);
and U5860 (N_5860,N_5700,N_5670);
or U5861 (N_5861,N_5714,N_5615);
nor U5862 (N_5862,N_5764,N_5629);
or U5863 (N_5863,N_5766,N_5626);
nand U5864 (N_5864,N_5694,N_5791);
xor U5865 (N_5865,N_5647,N_5640);
nor U5866 (N_5866,N_5721,N_5613);
and U5867 (N_5867,N_5643,N_5699);
xor U5868 (N_5868,N_5790,N_5795);
nor U5869 (N_5869,N_5754,N_5774);
nand U5870 (N_5870,N_5655,N_5773);
nand U5871 (N_5871,N_5769,N_5738);
xnor U5872 (N_5872,N_5702,N_5779);
nand U5873 (N_5873,N_5675,N_5786);
nor U5874 (N_5874,N_5630,N_5792);
nand U5875 (N_5875,N_5725,N_5650);
xor U5876 (N_5876,N_5705,N_5616);
nor U5877 (N_5877,N_5704,N_5635);
xnor U5878 (N_5878,N_5706,N_5601);
and U5879 (N_5879,N_5796,N_5627);
xnor U5880 (N_5880,N_5684,N_5794);
or U5881 (N_5881,N_5632,N_5607);
nor U5882 (N_5882,N_5707,N_5625);
and U5883 (N_5883,N_5761,N_5693);
nor U5884 (N_5884,N_5651,N_5778);
and U5885 (N_5885,N_5653,N_5746);
and U5886 (N_5886,N_5709,N_5691);
nand U5887 (N_5887,N_5756,N_5780);
or U5888 (N_5888,N_5733,N_5618);
and U5889 (N_5889,N_5736,N_5690);
nand U5890 (N_5890,N_5698,N_5649);
or U5891 (N_5891,N_5637,N_5737);
and U5892 (N_5892,N_5753,N_5683);
and U5893 (N_5893,N_5619,N_5672);
and U5894 (N_5894,N_5765,N_5660);
nand U5895 (N_5895,N_5621,N_5624);
nand U5896 (N_5896,N_5623,N_5656);
nor U5897 (N_5897,N_5732,N_5686);
nor U5898 (N_5898,N_5763,N_5659);
nand U5899 (N_5899,N_5715,N_5742);
nor U5900 (N_5900,N_5647,N_5678);
nor U5901 (N_5901,N_5629,N_5617);
xor U5902 (N_5902,N_5792,N_5717);
and U5903 (N_5903,N_5712,N_5723);
or U5904 (N_5904,N_5700,N_5711);
or U5905 (N_5905,N_5680,N_5677);
or U5906 (N_5906,N_5727,N_5671);
or U5907 (N_5907,N_5673,N_5755);
or U5908 (N_5908,N_5790,N_5725);
nand U5909 (N_5909,N_5728,N_5634);
nand U5910 (N_5910,N_5793,N_5632);
or U5911 (N_5911,N_5744,N_5714);
or U5912 (N_5912,N_5600,N_5790);
or U5913 (N_5913,N_5715,N_5727);
and U5914 (N_5914,N_5795,N_5782);
nand U5915 (N_5915,N_5779,N_5665);
nand U5916 (N_5916,N_5649,N_5720);
xnor U5917 (N_5917,N_5742,N_5633);
and U5918 (N_5918,N_5788,N_5612);
nor U5919 (N_5919,N_5731,N_5735);
nor U5920 (N_5920,N_5660,N_5732);
and U5921 (N_5921,N_5693,N_5786);
nor U5922 (N_5922,N_5702,N_5659);
nand U5923 (N_5923,N_5664,N_5628);
nor U5924 (N_5924,N_5625,N_5785);
and U5925 (N_5925,N_5778,N_5600);
and U5926 (N_5926,N_5749,N_5739);
nand U5927 (N_5927,N_5740,N_5663);
nor U5928 (N_5928,N_5784,N_5682);
or U5929 (N_5929,N_5605,N_5603);
nor U5930 (N_5930,N_5605,N_5638);
nor U5931 (N_5931,N_5620,N_5652);
nand U5932 (N_5932,N_5642,N_5623);
and U5933 (N_5933,N_5665,N_5743);
and U5934 (N_5934,N_5777,N_5632);
nand U5935 (N_5935,N_5618,N_5727);
nor U5936 (N_5936,N_5651,N_5767);
or U5937 (N_5937,N_5728,N_5708);
nand U5938 (N_5938,N_5632,N_5746);
and U5939 (N_5939,N_5624,N_5657);
nand U5940 (N_5940,N_5742,N_5744);
nand U5941 (N_5941,N_5658,N_5601);
nor U5942 (N_5942,N_5612,N_5771);
nand U5943 (N_5943,N_5653,N_5736);
nor U5944 (N_5944,N_5684,N_5790);
and U5945 (N_5945,N_5618,N_5747);
nand U5946 (N_5946,N_5701,N_5769);
and U5947 (N_5947,N_5787,N_5667);
nand U5948 (N_5948,N_5642,N_5731);
nand U5949 (N_5949,N_5767,N_5726);
nor U5950 (N_5950,N_5630,N_5752);
or U5951 (N_5951,N_5776,N_5771);
nand U5952 (N_5952,N_5794,N_5737);
nand U5953 (N_5953,N_5676,N_5793);
and U5954 (N_5954,N_5609,N_5728);
nor U5955 (N_5955,N_5760,N_5643);
xor U5956 (N_5956,N_5634,N_5707);
or U5957 (N_5957,N_5799,N_5688);
nor U5958 (N_5958,N_5729,N_5739);
and U5959 (N_5959,N_5766,N_5699);
and U5960 (N_5960,N_5694,N_5770);
nor U5961 (N_5961,N_5715,N_5627);
nand U5962 (N_5962,N_5767,N_5698);
nor U5963 (N_5963,N_5715,N_5691);
nor U5964 (N_5964,N_5646,N_5762);
nor U5965 (N_5965,N_5638,N_5668);
nor U5966 (N_5966,N_5745,N_5693);
or U5967 (N_5967,N_5606,N_5611);
nand U5968 (N_5968,N_5730,N_5633);
or U5969 (N_5969,N_5668,N_5660);
nor U5970 (N_5970,N_5734,N_5727);
nand U5971 (N_5971,N_5782,N_5656);
nor U5972 (N_5972,N_5677,N_5774);
nand U5973 (N_5973,N_5755,N_5634);
or U5974 (N_5974,N_5726,N_5630);
and U5975 (N_5975,N_5660,N_5644);
or U5976 (N_5976,N_5713,N_5772);
and U5977 (N_5977,N_5703,N_5648);
nand U5978 (N_5978,N_5662,N_5630);
nor U5979 (N_5979,N_5732,N_5718);
nor U5980 (N_5980,N_5697,N_5612);
or U5981 (N_5981,N_5731,N_5744);
nor U5982 (N_5982,N_5631,N_5775);
or U5983 (N_5983,N_5737,N_5616);
nor U5984 (N_5984,N_5727,N_5604);
xor U5985 (N_5985,N_5765,N_5740);
nand U5986 (N_5986,N_5739,N_5753);
nand U5987 (N_5987,N_5753,N_5659);
or U5988 (N_5988,N_5676,N_5754);
xnor U5989 (N_5989,N_5797,N_5738);
and U5990 (N_5990,N_5786,N_5702);
nor U5991 (N_5991,N_5673,N_5767);
or U5992 (N_5992,N_5706,N_5651);
or U5993 (N_5993,N_5605,N_5724);
nor U5994 (N_5994,N_5703,N_5666);
nand U5995 (N_5995,N_5744,N_5798);
or U5996 (N_5996,N_5657,N_5784);
xor U5997 (N_5997,N_5776,N_5662);
nor U5998 (N_5998,N_5617,N_5734);
xor U5999 (N_5999,N_5610,N_5647);
and U6000 (N_6000,N_5908,N_5803);
xor U6001 (N_6001,N_5893,N_5901);
or U6002 (N_6002,N_5991,N_5888);
or U6003 (N_6003,N_5897,N_5883);
and U6004 (N_6004,N_5932,N_5921);
xnor U6005 (N_6005,N_5909,N_5802);
or U6006 (N_6006,N_5885,N_5920);
or U6007 (N_6007,N_5984,N_5842);
xnor U6008 (N_6008,N_5959,N_5934);
xor U6009 (N_6009,N_5847,N_5986);
nand U6010 (N_6010,N_5933,N_5856);
and U6011 (N_6011,N_5840,N_5969);
nand U6012 (N_6012,N_5822,N_5823);
or U6013 (N_6013,N_5992,N_5956);
or U6014 (N_6014,N_5927,N_5819);
or U6015 (N_6015,N_5845,N_5974);
or U6016 (N_6016,N_5983,N_5943);
nor U6017 (N_6017,N_5846,N_5931);
and U6018 (N_6018,N_5994,N_5855);
or U6019 (N_6019,N_5980,N_5841);
nand U6020 (N_6020,N_5830,N_5825);
and U6021 (N_6021,N_5807,N_5961);
or U6022 (N_6022,N_5863,N_5907);
nand U6023 (N_6023,N_5915,N_5996);
nor U6024 (N_6024,N_5940,N_5820);
and U6025 (N_6025,N_5926,N_5951);
and U6026 (N_6026,N_5970,N_5862);
nor U6027 (N_6027,N_5857,N_5900);
nor U6028 (N_6028,N_5880,N_5817);
nand U6029 (N_6029,N_5896,N_5828);
xor U6030 (N_6030,N_5816,N_5844);
or U6031 (N_6031,N_5982,N_5950);
or U6032 (N_6032,N_5913,N_5884);
nor U6033 (N_6033,N_5924,N_5914);
nand U6034 (N_6034,N_5870,N_5912);
nand U6035 (N_6035,N_5916,N_5918);
nand U6036 (N_6036,N_5824,N_5800);
nor U6037 (N_6037,N_5833,N_5922);
nor U6038 (N_6038,N_5962,N_5904);
nand U6039 (N_6039,N_5902,N_5892);
nand U6040 (N_6040,N_5850,N_5910);
and U6041 (N_6041,N_5939,N_5874);
and U6042 (N_6042,N_5949,N_5942);
nor U6043 (N_6043,N_5864,N_5806);
and U6044 (N_6044,N_5854,N_5968);
xor U6045 (N_6045,N_5911,N_5865);
nand U6046 (N_6046,N_5848,N_5990);
or U6047 (N_6047,N_5919,N_5898);
nor U6048 (N_6048,N_5801,N_5960);
xnor U6049 (N_6049,N_5937,N_5946);
or U6050 (N_6050,N_5882,N_5987);
nand U6051 (N_6051,N_5938,N_5829);
nand U6052 (N_6052,N_5995,N_5835);
nand U6053 (N_6053,N_5948,N_5886);
nor U6054 (N_6054,N_5903,N_5813);
and U6055 (N_6055,N_5944,N_5941);
or U6056 (N_6056,N_5851,N_5930);
or U6057 (N_6057,N_5860,N_5836);
and U6058 (N_6058,N_5975,N_5832);
or U6059 (N_6059,N_5834,N_5977);
and U6060 (N_6060,N_5804,N_5869);
nor U6061 (N_6061,N_5853,N_5945);
and U6062 (N_6062,N_5837,N_5891);
nor U6063 (N_6063,N_5952,N_5859);
or U6064 (N_6064,N_5954,N_5867);
nor U6065 (N_6065,N_5917,N_5923);
xor U6066 (N_6066,N_5890,N_5895);
nor U6067 (N_6067,N_5811,N_5972);
nand U6068 (N_6068,N_5878,N_5973);
and U6069 (N_6069,N_5989,N_5875);
xnor U6070 (N_6070,N_5849,N_5852);
xnor U6071 (N_6071,N_5827,N_5947);
and U6072 (N_6072,N_5929,N_5861);
xnor U6073 (N_6073,N_5964,N_5858);
and U6074 (N_6074,N_5831,N_5873);
and U6075 (N_6075,N_5957,N_5818);
xor U6076 (N_6076,N_5887,N_5976);
nor U6077 (N_6077,N_5843,N_5899);
nor U6078 (N_6078,N_5905,N_5826);
and U6079 (N_6079,N_5928,N_5871);
or U6080 (N_6080,N_5971,N_5877);
nand U6081 (N_6081,N_5985,N_5935);
nor U6082 (N_6082,N_5963,N_5868);
and U6083 (N_6083,N_5815,N_5906);
and U6084 (N_6084,N_5879,N_5889);
and U6085 (N_6085,N_5988,N_5876);
and U6086 (N_6086,N_5958,N_5809);
nor U6087 (N_6087,N_5978,N_5808);
and U6088 (N_6088,N_5981,N_5965);
and U6089 (N_6089,N_5955,N_5999);
nor U6090 (N_6090,N_5821,N_5953);
and U6091 (N_6091,N_5936,N_5894);
nand U6092 (N_6092,N_5979,N_5966);
or U6093 (N_6093,N_5998,N_5997);
nor U6094 (N_6094,N_5872,N_5805);
nand U6095 (N_6095,N_5814,N_5810);
nand U6096 (N_6096,N_5881,N_5812);
nand U6097 (N_6097,N_5839,N_5925);
nand U6098 (N_6098,N_5866,N_5967);
xor U6099 (N_6099,N_5838,N_5993);
nor U6100 (N_6100,N_5924,N_5840);
nor U6101 (N_6101,N_5900,N_5829);
nor U6102 (N_6102,N_5983,N_5908);
nand U6103 (N_6103,N_5912,N_5840);
nand U6104 (N_6104,N_5899,N_5964);
xor U6105 (N_6105,N_5836,N_5930);
nor U6106 (N_6106,N_5832,N_5993);
xor U6107 (N_6107,N_5976,N_5963);
nor U6108 (N_6108,N_5844,N_5840);
nand U6109 (N_6109,N_5946,N_5831);
nor U6110 (N_6110,N_5958,N_5879);
and U6111 (N_6111,N_5903,N_5875);
nand U6112 (N_6112,N_5807,N_5958);
and U6113 (N_6113,N_5986,N_5882);
and U6114 (N_6114,N_5935,N_5995);
nor U6115 (N_6115,N_5926,N_5855);
nand U6116 (N_6116,N_5952,N_5877);
and U6117 (N_6117,N_5871,N_5938);
nand U6118 (N_6118,N_5964,N_5947);
nand U6119 (N_6119,N_5997,N_5875);
nor U6120 (N_6120,N_5879,N_5986);
and U6121 (N_6121,N_5935,N_5848);
or U6122 (N_6122,N_5997,N_5914);
nand U6123 (N_6123,N_5961,N_5863);
nand U6124 (N_6124,N_5812,N_5806);
or U6125 (N_6125,N_5995,N_5878);
nand U6126 (N_6126,N_5919,N_5872);
or U6127 (N_6127,N_5965,N_5878);
nor U6128 (N_6128,N_5995,N_5881);
or U6129 (N_6129,N_5942,N_5893);
and U6130 (N_6130,N_5913,N_5999);
xnor U6131 (N_6131,N_5955,N_5976);
and U6132 (N_6132,N_5969,N_5917);
nor U6133 (N_6133,N_5918,N_5906);
nand U6134 (N_6134,N_5821,N_5833);
nand U6135 (N_6135,N_5905,N_5801);
or U6136 (N_6136,N_5917,N_5855);
and U6137 (N_6137,N_5837,N_5841);
or U6138 (N_6138,N_5856,N_5937);
and U6139 (N_6139,N_5814,N_5956);
or U6140 (N_6140,N_5926,N_5975);
nor U6141 (N_6141,N_5982,N_5810);
or U6142 (N_6142,N_5848,N_5897);
nand U6143 (N_6143,N_5985,N_5819);
nor U6144 (N_6144,N_5885,N_5810);
nand U6145 (N_6145,N_5851,N_5966);
and U6146 (N_6146,N_5930,N_5934);
and U6147 (N_6147,N_5853,N_5854);
xor U6148 (N_6148,N_5846,N_5910);
nand U6149 (N_6149,N_5873,N_5899);
and U6150 (N_6150,N_5847,N_5859);
nor U6151 (N_6151,N_5983,N_5988);
nand U6152 (N_6152,N_5923,N_5856);
xor U6153 (N_6153,N_5875,N_5965);
and U6154 (N_6154,N_5829,N_5817);
nand U6155 (N_6155,N_5954,N_5841);
nand U6156 (N_6156,N_5956,N_5959);
nand U6157 (N_6157,N_5841,N_5828);
nor U6158 (N_6158,N_5967,N_5937);
nand U6159 (N_6159,N_5978,N_5837);
nor U6160 (N_6160,N_5847,N_5960);
nand U6161 (N_6161,N_5858,N_5894);
and U6162 (N_6162,N_5854,N_5904);
and U6163 (N_6163,N_5861,N_5847);
or U6164 (N_6164,N_5951,N_5992);
nor U6165 (N_6165,N_5800,N_5889);
and U6166 (N_6166,N_5831,N_5916);
or U6167 (N_6167,N_5921,N_5970);
and U6168 (N_6168,N_5931,N_5818);
xor U6169 (N_6169,N_5954,N_5827);
nand U6170 (N_6170,N_5813,N_5967);
and U6171 (N_6171,N_5972,N_5801);
nor U6172 (N_6172,N_5885,N_5906);
nor U6173 (N_6173,N_5960,N_5932);
nand U6174 (N_6174,N_5958,N_5802);
xnor U6175 (N_6175,N_5970,N_5927);
nor U6176 (N_6176,N_5803,N_5958);
xnor U6177 (N_6177,N_5977,N_5819);
or U6178 (N_6178,N_5850,N_5979);
xor U6179 (N_6179,N_5883,N_5806);
nor U6180 (N_6180,N_5965,N_5883);
and U6181 (N_6181,N_5963,N_5923);
and U6182 (N_6182,N_5820,N_5801);
or U6183 (N_6183,N_5864,N_5914);
and U6184 (N_6184,N_5925,N_5968);
xor U6185 (N_6185,N_5869,N_5896);
nor U6186 (N_6186,N_5934,N_5936);
nor U6187 (N_6187,N_5903,N_5802);
nand U6188 (N_6188,N_5995,N_5986);
nor U6189 (N_6189,N_5940,N_5802);
and U6190 (N_6190,N_5938,N_5977);
nor U6191 (N_6191,N_5823,N_5938);
nand U6192 (N_6192,N_5907,N_5868);
or U6193 (N_6193,N_5831,N_5867);
nor U6194 (N_6194,N_5966,N_5832);
or U6195 (N_6195,N_5929,N_5872);
nor U6196 (N_6196,N_5950,N_5921);
and U6197 (N_6197,N_5904,N_5909);
or U6198 (N_6198,N_5859,N_5875);
and U6199 (N_6199,N_5936,N_5984);
or U6200 (N_6200,N_6055,N_6049);
and U6201 (N_6201,N_6050,N_6114);
xor U6202 (N_6202,N_6152,N_6022);
nor U6203 (N_6203,N_6027,N_6193);
xor U6204 (N_6204,N_6032,N_6110);
nand U6205 (N_6205,N_6190,N_6174);
and U6206 (N_6206,N_6175,N_6011);
and U6207 (N_6207,N_6028,N_6144);
nand U6208 (N_6208,N_6093,N_6108);
nor U6209 (N_6209,N_6173,N_6184);
xor U6210 (N_6210,N_6072,N_6171);
nand U6211 (N_6211,N_6170,N_6001);
or U6212 (N_6212,N_6164,N_6165);
nand U6213 (N_6213,N_6120,N_6163);
or U6214 (N_6214,N_6155,N_6020);
or U6215 (N_6215,N_6185,N_6194);
and U6216 (N_6216,N_6141,N_6034);
or U6217 (N_6217,N_6076,N_6063);
and U6218 (N_6218,N_6062,N_6094);
nor U6219 (N_6219,N_6104,N_6147);
and U6220 (N_6220,N_6107,N_6199);
nor U6221 (N_6221,N_6159,N_6198);
nand U6222 (N_6222,N_6065,N_6189);
and U6223 (N_6223,N_6115,N_6151);
nand U6224 (N_6224,N_6187,N_6033);
nor U6225 (N_6225,N_6124,N_6186);
and U6226 (N_6226,N_6132,N_6145);
or U6227 (N_6227,N_6134,N_6161);
and U6228 (N_6228,N_6126,N_6087);
nand U6229 (N_6229,N_6018,N_6182);
nor U6230 (N_6230,N_6012,N_6168);
or U6231 (N_6231,N_6154,N_6057);
xor U6232 (N_6232,N_6118,N_6061);
and U6233 (N_6233,N_6127,N_6083);
nand U6234 (N_6234,N_6026,N_6178);
nand U6235 (N_6235,N_6024,N_6037);
xor U6236 (N_6236,N_6148,N_6162);
xnor U6237 (N_6237,N_6073,N_6074);
nand U6238 (N_6238,N_6146,N_6130);
nand U6239 (N_6239,N_6053,N_6002);
or U6240 (N_6240,N_6091,N_6166);
and U6241 (N_6241,N_6105,N_6160);
and U6242 (N_6242,N_6006,N_6112);
or U6243 (N_6243,N_6014,N_6101);
and U6244 (N_6244,N_6100,N_6111);
nand U6245 (N_6245,N_6025,N_6125);
or U6246 (N_6246,N_6128,N_6031);
and U6247 (N_6247,N_6121,N_6029);
nand U6248 (N_6248,N_6019,N_6149);
nor U6249 (N_6249,N_6113,N_6096);
nand U6250 (N_6250,N_6059,N_6188);
nand U6251 (N_6251,N_6038,N_6017);
nand U6252 (N_6252,N_6047,N_6090);
xor U6253 (N_6253,N_6004,N_6137);
xnor U6254 (N_6254,N_6139,N_6010);
nor U6255 (N_6255,N_6117,N_6181);
and U6256 (N_6256,N_6007,N_6084);
nor U6257 (N_6257,N_6157,N_6098);
or U6258 (N_6258,N_6030,N_6085);
nor U6259 (N_6259,N_6016,N_6179);
nor U6260 (N_6260,N_6092,N_6015);
nor U6261 (N_6261,N_6067,N_6080);
and U6262 (N_6262,N_6035,N_6150);
xor U6263 (N_6263,N_6099,N_6070);
xor U6264 (N_6264,N_6036,N_6068);
nand U6265 (N_6265,N_6077,N_6013);
nor U6266 (N_6266,N_6140,N_6097);
xor U6267 (N_6267,N_6088,N_6078);
and U6268 (N_6268,N_6109,N_6176);
or U6269 (N_6269,N_6039,N_6003);
or U6270 (N_6270,N_6042,N_6051);
nand U6271 (N_6271,N_6023,N_6075);
nand U6272 (N_6272,N_6046,N_6069);
nor U6273 (N_6273,N_6054,N_6143);
and U6274 (N_6274,N_6005,N_6138);
nor U6275 (N_6275,N_6066,N_6116);
nand U6276 (N_6276,N_6169,N_6060);
nor U6277 (N_6277,N_6191,N_6056);
or U6278 (N_6278,N_6177,N_6123);
nor U6279 (N_6279,N_6180,N_6009);
or U6280 (N_6280,N_6048,N_6089);
nor U6281 (N_6281,N_6196,N_6082);
and U6282 (N_6282,N_6045,N_6133);
and U6283 (N_6283,N_6122,N_6095);
nor U6284 (N_6284,N_6064,N_6041);
nor U6285 (N_6285,N_6021,N_6192);
nor U6286 (N_6286,N_6153,N_6000);
nand U6287 (N_6287,N_6142,N_6135);
or U6288 (N_6288,N_6119,N_6195);
and U6289 (N_6289,N_6129,N_6043);
nand U6290 (N_6290,N_6086,N_6197);
xnor U6291 (N_6291,N_6167,N_6071);
and U6292 (N_6292,N_6103,N_6106);
nor U6293 (N_6293,N_6079,N_6081);
nand U6294 (N_6294,N_6172,N_6136);
nor U6295 (N_6295,N_6008,N_6158);
or U6296 (N_6296,N_6058,N_6183);
nor U6297 (N_6297,N_6131,N_6102);
nor U6298 (N_6298,N_6156,N_6040);
nand U6299 (N_6299,N_6044,N_6052);
nor U6300 (N_6300,N_6030,N_6106);
and U6301 (N_6301,N_6123,N_6002);
or U6302 (N_6302,N_6036,N_6193);
nor U6303 (N_6303,N_6116,N_6165);
nand U6304 (N_6304,N_6189,N_6199);
nor U6305 (N_6305,N_6048,N_6149);
or U6306 (N_6306,N_6140,N_6134);
and U6307 (N_6307,N_6113,N_6151);
xnor U6308 (N_6308,N_6064,N_6159);
xnor U6309 (N_6309,N_6182,N_6186);
and U6310 (N_6310,N_6079,N_6067);
nor U6311 (N_6311,N_6024,N_6141);
nor U6312 (N_6312,N_6139,N_6167);
or U6313 (N_6313,N_6185,N_6159);
or U6314 (N_6314,N_6068,N_6017);
nor U6315 (N_6315,N_6028,N_6073);
or U6316 (N_6316,N_6097,N_6056);
or U6317 (N_6317,N_6117,N_6091);
nand U6318 (N_6318,N_6173,N_6059);
nand U6319 (N_6319,N_6023,N_6015);
nor U6320 (N_6320,N_6160,N_6152);
and U6321 (N_6321,N_6056,N_6078);
nand U6322 (N_6322,N_6186,N_6159);
or U6323 (N_6323,N_6131,N_6135);
nor U6324 (N_6324,N_6026,N_6053);
xor U6325 (N_6325,N_6051,N_6016);
and U6326 (N_6326,N_6092,N_6061);
nand U6327 (N_6327,N_6002,N_6129);
and U6328 (N_6328,N_6037,N_6141);
or U6329 (N_6329,N_6013,N_6190);
or U6330 (N_6330,N_6014,N_6125);
xnor U6331 (N_6331,N_6005,N_6090);
and U6332 (N_6332,N_6033,N_6100);
or U6333 (N_6333,N_6036,N_6043);
or U6334 (N_6334,N_6095,N_6030);
nand U6335 (N_6335,N_6173,N_6093);
xnor U6336 (N_6336,N_6117,N_6086);
nand U6337 (N_6337,N_6150,N_6095);
and U6338 (N_6338,N_6129,N_6101);
nand U6339 (N_6339,N_6111,N_6069);
or U6340 (N_6340,N_6181,N_6151);
xor U6341 (N_6341,N_6161,N_6063);
nand U6342 (N_6342,N_6130,N_6111);
nor U6343 (N_6343,N_6127,N_6086);
xor U6344 (N_6344,N_6125,N_6161);
and U6345 (N_6345,N_6007,N_6109);
xor U6346 (N_6346,N_6025,N_6103);
or U6347 (N_6347,N_6103,N_6141);
and U6348 (N_6348,N_6026,N_6079);
nor U6349 (N_6349,N_6146,N_6051);
or U6350 (N_6350,N_6172,N_6120);
or U6351 (N_6351,N_6106,N_6096);
and U6352 (N_6352,N_6194,N_6020);
and U6353 (N_6353,N_6032,N_6044);
and U6354 (N_6354,N_6123,N_6168);
and U6355 (N_6355,N_6163,N_6185);
or U6356 (N_6356,N_6148,N_6049);
and U6357 (N_6357,N_6168,N_6081);
or U6358 (N_6358,N_6049,N_6014);
and U6359 (N_6359,N_6128,N_6058);
nor U6360 (N_6360,N_6114,N_6007);
nor U6361 (N_6361,N_6083,N_6199);
nor U6362 (N_6362,N_6146,N_6056);
nor U6363 (N_6363,N_6194,N_6104);
or U6364 (N_6364,N_6083,N_6144);
or U6365 (N_6365,N_6086,N_6055);
xor U6366 (N_6366,N_6071,N_6096);
nand U6367 (N_6367,N_6082,N_6169);
or U6368 (N_6368,N_6089,N_6084);
or U6369 (N_6369,N_6090,N_6186);
xor U6370 (N_6370,N_6162,N_6072);
nand U6371 (N_6371,N_6024,N_6111);
and U6372 (N_6372,N_6179,N_6131);
xor U6373 (N_6373,N_6139,N_6067);
or U6374 (N_6374,N_6101,N_6065);
and U6375 (N_6375,N_6007,N_6075);
and U6376 (N_6376,N_6145,N_6118);
or U6377 (N_6377,N_6135,N_6060);
nand U6378 (N_6378,N_6176,N_6179);
and U6379 (N_6379,N_6185,N_6080);
nand U6380 (N_6380,N_6164,N_6103);
and U6381 (N_6381,N_6157,N_6155);
nor U6382 (N_6382,N_6180,N_6073);
nor U6383 (N_6383,N_6142,N_6119);
or U6384 (N_6384,N_6123,N_6062);
nand U6385 (N_6385,N_6055,N_6015);
nand U6386 (N_6386,N_6160,N_6095);
nand U6387 (N_6387,N_6105,N_6094);
nand U6388 (N_6388,N_6095,N_6076);
and U6389 (N_6389,N_6158,N_6028);
nand U6390 (N_6390,N_6185,N_6186);
or U6391 (N_6391,N_6107,N_6082);
and U6392 (N_6392,N_6150,N_6055);
and U6393 (N_6393,N_6189,N_6140);
nor U6394 (N_6394,N_6165,N_6163);
nor U6395 (N_6395,N_6129,N_6014);
nor U6396 (N_6396,N_6121,N_6060);
or U6397 (N_6397,N_6061,N_6045);
nand U6398 (N_6398,N_6156,N_6147);
nor U6399 (N_6399,N_6149,N_6136);
nand U6400 (N_6400,N_6261,N_6360);
nand U6401 (N_6401,N_6378,N_6384);
nand U6402 (N_6402,N_6367,N_6228);
or U6403 (N_6403,N_6322,N_6336);
or U6404 (N_6404,N_6220,N_6246);
or U6405 (N_6405,N_6293,N_6340);
xor U6406 (N_6406,N_6201,N_6395);
nor U6407 (N_6407,N_6390,N_6326);
nand U6408 (N_6408,N_6392,N_6234);
nor U6409 (N_6409,N_6212,N_6265);
and U6410 (N_6410,N_6352,N_6289);
nor U6411 (N_6411,N_6345,N_6240);
nor U6412 (N_6412,N_6306,N_6274);
nor U6413 (N_6413,N_6343,N_6208);
nand U6414 (N_6414,N_6210,N_6350);
nor U6415 (N_6415,N_6218,N_6215);
nand U6416 (N_6416,N_6281,N_6376);
and U6417 (N_6417,N_6248,N_6317);
and U6418 (N_6418,N_6348,N_6278);
or U6419 (N_6419,N_6233,N_6335);
nor U6420 (N_6420,N_6344,N_6205);
xnor U6421 (N_6421,N_6353,N_6391);
nor U6422 (N_6422,N_6372,N_6318);
xor U6423 (N_6423,N_6200,N_6251);
nor U6424 (N_6424,N_6374,N_6347);
and U6425 (N_6425,N_6370,N_6255);
and U6426 (N_6426,N_6332,N_6300);
or U6427 (N_6427,N_6252,N_6260);
or U6428 (N_6428,N_6341,N_6371);
xnor U6429 (N_6429,N_6280,N_6393);
nand U6430 (N_6430,N_6329,N_6387);
and U6431 (N_6431,N_6250,N_6377);
and U6432 (N_6432,N_6375,N_6364);
and U6433 (N_6433,N_6373,N_6256);
nand U6434 (N_6434,N_6295,N_6386);
nand U6435 (N_6435,N_6325,N_6357);
xnor U6436 (N_6436,N_6292,N_6365);
nor U6437 (N_6437,N_6206,N_6358);
and U6438 (N_6438,N_6238,N_6302);
nor U6439 (N_6439,N_6202,N_6346);
nor U6440 (N_6440,N_6369,N_6337);
and U6441 (N_6441,N_6224,N_6389);
and U6442 (N_6442,N_6236,N_6253);
nand U6443 (N_6443,N_6258,N_6291);
or U6444 (N_6444,N_6323,N_6383);
xor U6445 (N_6445,N_6259,N_6394);
nand U6446 (N_6446,N_6269,N_6241);
or U6447 (N_6447,N_6328,N_6270);
nand U6448 (N_6448,N_6217,N_6207);
or U6449 (N_6449,N_6320,N_6286);
nand U6450 (N_6450,N_6338,N_6361);
or U6451 (N_6451,N_6264,N_6211);
nand U6452 (N_6452,N_6223,N_6382);
or U6453 (N_6453,N_6339,N_6333);
and U6454 (N_6454,N_6214,N_6221);
or U6455 (N_6455,N_6283,N_6277);
or U6456 (N_6456,N_6307,N_6399);
or U6457 (N_6457,N_6299,N_6242);
nor U6458 (N_6458,N_6225,N_6279);
nand U6459 (N_6459,N_6355,N_6366);
xor U6460 (N_6460,N_6334,N_6310);
and U6461 (N_6461,N_6308,N_6230);
nand U6462 (N_6462,N_6349,N_6247);
nor U6463 (N_6463,N_6271,N_6237);
nand U6464 (N_6464,N_6330,N_6356);
nor U6465 (N_6465,N_6268,N_6313);
nor U6466 (N_6466,N_6213,N_6351);
or U6467 (N_6467,N_6319,N_6232);
or U6468 (N_6468,N_6362,N_6327);
nand U6469 (N_6469,N_6316,N_6231);
or U6470 (N_6470,N_6209,N_6282);
xnor U6471 (N_6471,N_6203,N_6396);
and U6472 (N_6472,N_6388,N_6312);
and U6473 (N_6473,N_6226,N_6398);
or U6474 (N_6474,N_6303,N_6311);
or U6475 (N_6475,N_6315,N_6368);
and U6476 (N_6476,N_6397,N_6273);
and U6477 (N_6477,N_6298,N_6284);
or U6478 (N_6478,N_6288,N_6229);
nand U6479 (N_6479,N_6359,N_6272);
or U6480 (N_6480,N_6235,N_6296);
or U6481 (N_6481,N_6263,N_6309);
nand U6482 (N_6482,N_6219,N_6342);
nor U6483 (N_6483,N_6324,N_6243);
or U6484 (N_6484,N_6275,N_6204);
nor U6485 (N_6485,N_6287,N_6267);
and U6486 (N_6486,N_6305,N_6257);
nor U6487 (N_6487,N_6314,N_6244);
and U6488 (N_6488,N_6354,N_6276);
and U6489 (N_6489,N_6294,N_6290);
nor U6490 (N_6490,N_6380,N_6239);
and U6491 (N_6491,N_6262,N_6254);
and U6492 (N_6492,N_6363,N_6385);
or U6493 (N_6493,N_6304,N_6249);
and U6494 (N_6494,N_6266,N_6379);
xnor U6495 (N_6495,N_6216,N_6222);
nor U6496 (N_6496,N_6285,N_6381);
nand U6497 (N_6497,N_6227,N_6321);
and U6498 (N_6498,N_6297,N_6331);
or U6499 (N_6499,N_6301,N_6245);
nand U6500 (N_6500,N_6276,N_6267);
nand U6501 (N_6501,N_6280,N_6269);
or U6502 (N_6502,N_6350,N_6373);
nand U6503 (N_6503,N_6232,N_6267);
and U6504 (N_6504,N_6250,N_6264);
and U6505 (N_6505,N_6340,N_6279);
nand U6506 (N_6506,N_6334,N_6325);
nor U6507 (N_6507,N_6280,N_6329);
and U6508 (N_6508,N_6219,N_6205);
nor U6509 (N_6509,N_6295,N_6314);
and U6510 (N_6510,N_6296,N_6239);
nor U6511 (N_6511,N_6202,N_6384);
or U6512 (N_6512,N_6200,N_6264);
or U6513 (N_6513,N_6386,N_6279);
and U6514 (N_6514,N_6220,N_6374);
nor U6515 (N_6515,N_6343,N_6366);
and U6516 (N_6516,N_6241,N_6217);
nand U6517 (N_6517,N_6237,N_6200);
nor U6518 (N_6518,N_6309,N_6287);
nor U6519 (N_6519,N_6315,N_6211);
nand U6520 (N_6520,N_6340,N_6371);
or U6521 (N_6521,N_6396,N_6278);
and U6522 (N_6522,N_6291,N_6296);
nand U6523 (N_6523,N_6272,N_6312);
nand U6524 (N_6524,N_6285,N_6307);
or U6525 (N_6525,N_6236,N_6230);
nand U6526 (N_6526,N_6220,N_6202);
and U6527 (N_6527,N_6229,N_6356);
nor U6528 (N_6528,N_6376,N_6377);
nor U6529 (N_6529,N_6338,N_6362);
nand U6530 (N_6530,N_6278,N_6219);
nor U6531 (N_6531,N_6216,N_6236);
and U6532 (N_6532,N_6318,N_6350);
nand U6533 (N_6533,N_6358,N_6366);
nor U6534 (N_6534,N_6313,N_6233);
nand U6535 (N_6535,N_6306,N_6216);
nand U6536 (N_6536,N_6224,N_6222);
nor U6537 (N_6537,N_6388,N_6334);
xnor U6538 (N_6538,N_6399,N_6260);
xor U6539 (N_6539,N_6256,N_6229);
and U6540 (N_6540,N_6329,N_6344);
or U6541 (N_6541,N_6226,N_6276);
xor U6542 (N_6542,N_6296,N_6238);
or U6543 (N_6543,N_6369,N_6280);
nand U6544 (N_6544,N_6244,N_6376);
nand U6545 (N_6545,N_6272,N_6294);
and U6546 (N_6546,N_6230,N_6262);
and U6547 (N_6547,N_6359,N_6318);
and U6548 (N_6548,N_6303,N_6316);
or U6549 (N_6549,N_6322,N_6310);
nor U6550 (N_6550,N_6373,N_6269);
nor U6551 (N_6551,N_6397,N_6308);
nand U6552 (N_6552,N_6265,N_6235);
and U6553 (N_6553,N_6296,N_6207);
and U6554 (N_6554,N_6263,N_6361);
nor U6555 (N_6555,N_6331,N_6358);
xor U6556 (N_6556,N_6233,N_6219);
and U6557 (N_6557,N_6282,N_6225);
and U6558 (N_6558,N_6201,N_6360);
and U6559 (N_6559,N_6265,N_6242);
and U6560 (N_6560,N_6250,N_6342);
nor U6561 (N_6561,N_6342,N_6308);
nor U6562 (N_6562,N_6275,N_6319);
or U6563 (N_6563,N_6232,N_6202);
nand U6564 (N_6564,N_6231,N_6349);
nor U6565 (N_6565,N_6306,N_6389);
nand U6566 (N_6566,N_6373,N_6249);
and U6567 (N_6567,N_6212,N_6323);
and U6568 (N_6568,N_6357,N_6232);
or U6569 (N_6569,N_6303,N_6375);
nand U6570 (N_6570,N_6224,N_6356);
or U6571 (N_6571,N_6392,N_6207);
or U6572 (N_6572,N_6310,N_6213);
or U6573 (N_6573,N_6346,N_6375);
or U6574 (N_6574,N_6244,N_6294);
nand U6575 (N_6575,N_6352,N_6216);
nand U6576 (N_6576,N_6350,N_6254);
and U6577 (N_6577,N_6221,N_6212);
nor U6578 (N_6578,N_6338,N_6341);
nor U6579 (N_6579,N_6284,N_6339);
nor U6580 (N_6580,N_6249,N_6379);
or U6581 (N_6581,N_6327,N_6302);
nand U6582 (N_6582,N_6223,N_6399);
and U6583 (N_6583,N_6389,N_6213);
nor U6584 (N_6584,N_6399,N_6285);
or U6585 (N_6585,N_6396,N_6241);
nor U6586 (N_6586,N_6372,N_6260);
nand U6587 (N_6587,N_6375,N_6314);
nand U6588 (N_6588,N_6367,N_6259);
or U6589 (N_6589,N_6384,N_6359);
nand U6590 (N_6590,N_6338,N_6354);
or U6591 (N_6591,N_6374,N_6354);
xnor U6592 (N_6592,N_6211,N_6283);
nand U6593 (N_6593,N_6373,N_6295);
nand U6594 (N_6594,N_6220,N_6366);
and U6595 (N_6595,N_6330,N_6235);
nor U6596 (N_6596,N_6328,N_6262);
nor U6597 (N_6597,N_6290,N_6247);
nand U6598 (N_6598,N_6326,N_6343);
and U6599 (N_6599,N_6217,N_6221);
or U6600 (N_6600,N_6426,N_6580);
or U6601 (N_6601,N_6512,N_6553);
xnor U6602 (N_6602,N_6561,N_6596);
nand U6603 (N_6603,N_6501,N_6506);
nand U6604 (N_6604,N_6481,N_6466);
nor U6605 (N_6605,N_6532,N_6443);
nor U6606 (N_6606,N_6507,N_6499);
nor U6607 (N_6607,N_6504,N_6489);
nand U6608 (N_6608,N_6471,N_6564);
xnor U6609 (N_6609,N_6413,N_6459);
and U6610 (N_6610,N_6474,N_6478);
and U6611 (N_6611,N_6505,N_6533);
and U6612 (N_6612,N_6563,N_6467);
nand U6613 (N_6613,N_6503,N_6486);
and U6614 (N_6614,N_6530,N_6531);
or U6615 (N_6615,N_6549,N_6415);
nor U6616 (N_6616,N_6482,N_6436);
nor U6617 (N_6617,N_6541,N_6452);
and U6618 (N_6618,N_6576,N_6449);
nand U6619 (N_6619,N_6516,N_6423);
xnor U6620 (N_6620,N_6416,N_6585);
and U6621 (N_6621,N_6597,N_6463);
or U6622 (N_6622,N_6528,N_6401);
and U6623 (N_6623,N_6554,N_6519);
nand U6624 (N_6624,N_6437,N_6494);
and U6625 (N_6625,N_6440,N_6404);
nand U6626 (N_6626,N_6445,N_6558);
nor U6627 (N_6627,N_6518,N_6575);
and U6628 (N_6628,N_6511,N_6570);
or U6629 (N_6629,N_6447,N_6484);
nand U6630 (N_6630,N_6525,N_6581);
and U6631 (N_6631,N_6582,N_6590);
nor U6632 (N_6632,N_6422,N_6534);
nand U6633 (N_6633,N_6565,N_6451);
nor U6634 (N_6634,N_6410,N_6599);
nand U6635 (N_6635,N_6411,N_6408);
xnor U6636 (N_6636,N_6479,N_6495);
and U6637 (N_6637,N_6450,N_6487);
or U6638 (N_6638,N_6402,N_6571);
or U6639 (N_6639,N_6557,N_6526);
or U6640 (N_6640,N_6566,N_6429);
or U6641 (N_6641,N_6417,N_6574);
nor U6642 (N_6642,N_6537,N_6591);
xor U6643 (N_6643,N_6509,N_6543);
and U6644 (N_6644,N_6588,N_6523);
or U6645 (N_6645,N_6577,N_6515);
and U6646 (N_6646,N_6435,N_6414);
nand U6647 (N_6647,N_6453,N_6510);
nand U6648 (N_6648,N_6400,N_6556);
and U6649 (N_6649,N_6475,N_6433);
and U6650 (N_6650,N_6545,N_6562);
and U6651 (N_6651,N_6444,N_6425);
nor U6652 (N_6652,N_6593,N_6418);
nand U6653 (N_6653,N_6491,N_6469);
nor U6654 (N_6654,N_6498,N_6483);
or U6655 (N_6655,N_6446,N_6420);
nand U6656 (N_6656,N_6465,N_6457);
nand U6657 (N_6657,N_6544,N_6559);
nor U6658 (N_6658,N_6522,N_6583);
nor U6659 (N_6659,N_6461,N_6555);
nand U6660 (N_6660,N_6578,N_6439);
nor U6661 (N_6661,N_6508,N_6502);
nand U6662 (N_6662,N_6527,N_6579);
nand U6663 (N_6663,N_6421,N_6595);
and U6664 (N_6664,N_6477,N_6464);
nor U6665 (N_6665,N_6455,N_6427);
nand U6666 (N_6666,N_6552,N_6535);
or U6667 (N_6667,N_6405,N_6419);
xor U6668 (N_6668,N_6517,N_6589);
nand U6669 (N_6669,N_6520,N_6598);
nor U6670 (N_6670,N_6428,N_6551);
and U6671 (N_6671,N_6536,N_6409);
and U6672 (N_6672,N_6513,N_6480);
nor U6673 (N_6673,N_6460,N_6472);
and U6674 (N_6674,N_6412,N_6406);
and U6675 (N_6675,N_6454,N_6547);
nor U6676 (N_6676,N_6485,N_6546);
or U6677 (N_6677,N_6573,N_6476);
nor U6678 (N_6678,N_6492,N_6497);
nand U6679 (N_6679,N_6458,N_6542);
and U6680 (N_6680,N_6424,N_6430);
nor U6681 (N_6681,N_6568,N_6403);
and U6682 (N_6682,N_6524,N_6540);
nand U6683 (N_6683,N_6584,N_6431);
nand U6684 (N_6684,N_6592,N_6490);
nor U6685 (N_6685,N_6468,N_6407);
or U6686 (N_6686,N_6448,N_6441);
and U6687 (N_6687,N_6496,N_6493);
nand U6688 (N_6688,N_6488,N_6500);
nor U6689 (N_6689,N_6586,N_6521);
nor U6690 (N_6690,N_6432,N_6587);
and U6691 (N_6691,N_6473,N_6550);
and U6692 (N_6692,N_6560,N_6569);
and U6693 (N_6693,N_6434,N_6548);
nand U6694 (N_6694,N_6456,N_6539);
nor U6695 (N_6695,N_6470,N_6572);
nand U6696 (N_6696,N_6438,N_6529);
nor U6697 (N_6697,N_6594,N_6567);
and U6698 (N_6698,N_6462,N_6538);
and U6699 (N_6699,N_6442,N_6514);
nor U6700 (N_6700,N_6596,N_6441);
or U6701 (N_6701,N_6588,N_6400);
or U6702 (N_6702,N_6468,N_6506);
or U6703 (N_6703,N_6456,N_6527);
nor U6704 (N_6704,N_6517,N_6451);
or U6705 (N_6705,N_6596,N_6540);
or U6706 (N_6706,N_6554,N_6470);
and U6707 (N_6707,N_6554,N_6503);
nand U6708 (N_6708,N_6522,N_6525);
xor U6709 (N_6709,N_6575,N_6567);
xor U6710 (N_6710,N_6462,N_6527);
or U6711 (N_6711,N_6429,N_6585);
xor U6712 (N_6712,N_6489,N_6442);
nand U6713 (N_6713,N_6457,N_6500);
nand U6714 (N_6714,N_6595,N_6476);
nor U6715 (N_6715,N_6495,N_6566);
and U6716 (N_6716,N_6464,N_6458);
nor U6717 (N_6717,N_6415,N_6459);
or U6718 (N_6718,N_6512,N_6561);
and U6719 (N_6719,N_6493,N_6439);
and U6720 (N_6720,N_6434,N_6554);
nor U6721 (N_6721,N_6402,N_6428);
and U6722 (N_6722,N_6596,N_6583);
and U6723 (N_6723,N_6486,N_6489);
xor U6724 (N_6724,N_6526,N_6448);
nor U6725 (N_6725,N_6536,N_6455);
nand U6726 (N_6726,N_6457,N_6452);
or U6727 (N_6727,N_6558,N_6438);
or U6728 (N_6728,N_6555,N_6519);
xor U6729 (N_6729,N_6407,N_6571);
xnor U6730 (N_6730,N_6469,N_6574);
or U6731 (N_6731,N_6479,N_6476);
nand U6732 (N_6732,N_6590,N_6545);
or U6733 (N_6733,N_6580,N_6586);
or U6734 (N_6734,N_6445,N_6420);
or U6735 (N_6735,N_6488,N_6544);
and U6736 (N_6736,N_6558,N_6471);
nor U6737 (N_6737,N_6490,N_6559);
or U6738 (N_6738,N_6584,N_6504);
and U6739 (N_6739,N_6405,N_6546);
xor U6740 (N_6740,N_6411,N_6545);
nor U6741 (N_6741,N_6540,N_6597);
nand U6742 (N_6742,N_6412,N_6445);
nand U6743 (N_6743,N_6437,N_6569);
or U6744 (N_6744,N_6542,N_6472);
xor U6745 (N_6745,N_6413,N_6480);
or U6746 (N_6746,N_6433,N_6572);
and U6747 (N_6747,N_6424,N_6508);
nor U6748 (N_6748,N_6406,N_6535);
nand U6749 (N_6749,N_6432,N_6438);
or U6750 (N_6750,N_6479,N_6459);
nor U6751 (N_6751,N_6463,N_6446);
or U6752 (N_6752,N_6562,N_6490);
or U6753 (N_6753,N_6455,N_6456);
or U6754 (N_6754,N_6499,N_6573);
or U6755 (N_6755,N_6446,N_6471);
or U6756 (N_6756,N_6443,N_6405);
and U6757 (N_6757,N_6490,N_6533);
nor U6758 (N_6758,N_6446,N_6421);
and U6759 (N_6759,N_6573,N_6570);
or U6760 (N_6760,N_6546,N_6490);
or U6761 (N_6761,N_6466,N_6505);
or U6762 (N_6762,N_6597,N_6562);
nand U6763 (N_6763,N_6557,N_6523);
nor U6764 (N_6764,N_6543,N_6435);
nand U6765 (N_6765,N_6553,N_6428);
nor U6766 (N_6766,N_6428,N_6443);
nor U6767 (N_6767,N_6555,N_6458);
or U6768 (N_6768,N_6530,N_6406);
nand U6769 (N_6769,N_6417,N_6437);
and U6770 (N_6770,N_6499,N_6581);
nand U6771 (N_6771,N_6573,N_6552);
and U6772 (N_6772,N_6593,N_6427);
nor U6773 (N_6773,N_6431,N_6497);
and U6774 (N_6774,N_6426,N_6553);
and U6775 (N_6775,N_6496,N_6582);
or U6776 (N_6776,N_6571,N_6528);
and U6777 (N_6777,N_6411,N_6420);
and U6778 (N_6778,N_6461,N_6491);
nand U6779 (N_6779,N_6464,N_6568);
or U6780 (N_6780,N_6479,N_6527);
nand U6781 (N_6781,N_6424,N_6521);
nand U6782 (N_6782,N_6518,N_6512);
nor U6783 (N_6783,N_6424,N_6421);
nand U6784 (N_6784,N_6462,N_6510);
nor U6785 (N_6785,N_6542,N_6536);
nor U6786 (N_6786,N_6571,N_6431);
and U6787 (N_6787,N_6410,N_6584);
or U6788 (N_6788,N_6543,N_6439);
or U6789 (N_6789,N_6550,N_6514);
or U6790 (N_6790,N_6506,N_6420);
nand U6791 (N_6791,N_6469,N_6417);
nand U6792 (N_6792,N_6461,N_6577);
and U6793 (N_6793,N_6438,N_6446);
nand U6794 (N_6794,N_6525,N_6560);
xnor U6795 (N_6795,N_6541,N_6521);
nand U6796 (N_6796,N_6530,N_6421);
or U6797 (N_6797,N_6583,N_6536);
and U6798 (N_6798,N_6518,N_6437);
or U6799 (N_6799,N_6415,N_6428);
nand U6800 (N_6800,N_6685,N_6705);
or U6801 (N_6801,N_6646,N_6780);
nor U6802 (N_6802,N_6601,N_6698);
nor U6803 (N_6803,N_6647,N_6747);
nor U6804 (N_6804,N_6654,N_6729);
nand U6805 (N_6805,N_6628,N_6740);
and U6806 (N_6806,N_6671,N_6795);
and U6807 (N_6807,N_6660,N_6731);
and U6808 (N_6808,N_6607,N_6641);
xnor U6809 (N_6809,N_6696,N_6781);
and U6810 (N_6810,N_6692,N_6603);
nand U6811 (N_6811,N_6694,N_6749);
or U6812 (N_6812,N_6699,N_6754);
or U6813 (N_6813,N_6663,N_6767);
nand U6814 (N_6814,N_6764,N_6703);
nand U6815 (N_6815,N_6732,N_6652);
or U6816 (N_6816,N_6612,N_6644);
or U6817 (N_6817,N_6674,N_6766);
nor U6818 (N_6818,N_6638,N_6668);
nand U6819 (N_6819,N_6773,N_6752);
and U6820 (N_6820,N_6717,N_6768);
xor U6821 (N_6821,N_6739,N_6622);
nor U6822 (N_6822,N_6742,N_6655);
nand U6823 (N_6823,N_6602,N_6770);
nand U6824 (N_6824,N_6600,N_6736);
nand U6825 (N_6825,N_6624,N_6720);
and U6826 (N_6826,N_6677,N_6621);
or U6827 (N_6827,N_6678,N_6667);
xor U6828 (N_6828,N_6799,N_6619);
nor U6829 (N_6829,N_6777,N_6785);
xor U6830 (N_6830,N_6772,N_6640);
and U6831 (N_6831,N_6711,N_6682);
nor U6832 (N_6832,N_6642,N_6750);
or U6833 (N_6833,N_6657,N_6690);
nand U6834 (N_6834,N_6760,N_6645);
and U6835 (N_6835,N_6710,N_6745);
or U6836 (N_6836,N_6616,N_6664);
and U6837 (N_6837,N_6629,N_6604);
nand U6838 (N_6838,N_6712,N_6669);
and U6839 (N_6839,N_6615,N_6700);
xnor U6840 (N_6840,N_6726,N_6709);
nand U6841 (N_6841,N_6761,N_6672);
or U6842 (N_6842,N_6613,N_6792);
or U6843 (N_6843,N_6673,N_6719);
nor U6844 (N_6844,N_6716,N_6756);
and U6845 (N_6845,N_6636,N_6730);
xnor U6846 (N_6846,N_6623,N_6786);
xor U6847 (N_6847,N_6606,N_6695);
xor U6848 (N_6848,N_6722,N_6751);
and U6849 (N_6849,N_6648,N_6693);
or U6850 (N_6850,N_6743,N_6704);
and U6851 (N_6851,N_6757,N_6630);
nand U6852 (N_6852,N_6782,N_6715);
or U6853 (N_6853,N_6775,N_6707);
or U6854 (N_6854,N_6733,N_6797);
nand U6855 (N_6855,N_6723,N_6609);
nor U6856 (N_6856,N_6608,N_6718);
nand U6857 (N_6857,N_6793,N_6683);
and U6858 (N_6858,N_6788,N_6784);
and U6859 (N_6859,N_6680,N_6681);
and U6860 (N_6860,N_6635,N_6759);
or U6861 (N_6861,N_6651,N_6627);
nand U6862 (N_6862,N_6789,N_6724);
nand U6863 (N_6863,N_6721,N_6738);
or U6864 (N_6864,N_6656,N_6611);
xor U6865 (N_6865,N_6670,N_6605);
and U6866 (N_6866,N_6637,N_6790);
and U6867 (N_6867,N_6755,N_6697);
nor U6868 (N_6868,N_6658,N_6684);
and U6869 (N_6869,N_6771,N_6686);
nor U6870 (N_6870,N_6762,N_6610);
or U6871 (N_6871,N_6714,N_6661);
xnor U6872 (N_6872,N_6735,N_6633);
nand U6873 (N_6873,N_6741,N_6713);
and U6874 (N_6874,N_6620,N_6691);
and U6875 (N_6875,N_6794,N_6769);
and U6876 (N_6876,N_6791,N_6765);
nand U6877 (N_6877,N_6702,N_6744);
xor U6878 (N_6878,N_6625,N_6676);
and U6879 (N_6879,N_6708,N_6753);
nand U6880 (N_6880,N_6779,N_6679);
nand U6881 (N_6881,N_6796,N_6798);
nor U6882 (N_6882,N_6659,N_6649);
nor U6883 (N_6883,N_6778,N_6737);
or U6884 (N_6884,N_6618,N_6643);
nand U6885 (N_6885,N_6631,N_6763);
and U6886 (N_6886,N_6758,N_6783);
and U6887 (N_6887,N_6665,N_6725);
and U6888 (N_6888,N_6776,N_6626);
xor U6889 (N_6889,N_6634,N_6688);
nor U6890 (N_6890,N_6650,N_6734);
nand U6891 (N_6891,N_6687,N_6706);
and U6892 (N_6892,N_6614,N_6728);
or U6893 (N_6893,N_6666,N_6675);
or U6894 (N_6894,N_6748,N_6662);
nand U6895 (N_6895,N_6787,N_6774);
nor U6896 (N_6896,N_6617,N_6632);
nand U6897 (N_6897,N_6639,N_6727);
nand U6898 (N_6898,N_6653,N_6746);
xor U6899 (N_6899,N_6689,N_6701);
and U6900 (N_6900,N_6795,N_6631);
nor U6901 (N_6901,N_6708,N_6700);
and U6902 (N_6902,N_6623,N_6675);
and U6903 (N_6903,N_6619,N_6641);
nor U6904 (N_6904,N_6768,N_6661);
and U6905 (N_6905,N_6733,N_6664);
or U6906 (N_6906,N_6693,N_6746);
and U6907 (N_6907,N_6750,N_6742);
nor U6908 (N_6908,N_6797,N_6650);
nand U6909 (N_6909,N_6635,N_6765);
nor U6910 (N_6910,N_6766,N_6695);
or U6911 (N_6911,N_6754,N_6783);
or U6912 (N_6912,N_6696,N_6715);
and U6913 (N_6913,N_6638,N_6738);
and U6914 (N_6914,N_6637,N_6683);
or U6915 (N_6915,N_6673,N_6726);
or U6916 (N_6916,N_6667,N_6726);
nand U6917 (N_6917,N_6795,N_6756);
xor U6918 (N_6918,N_6740,N_6694);
nand U6919 (N_6919,N_6766,N_6614);
nand U6920 (N_6920,N_6790,N_6636);
xor U6921 (N_6921,N_6766,N_6693);
and U6922 (N_6922,N_6625,N_6600);
nor U6923 (N_6923,N_6750,N_6719);
or U6924 (N_6924,N_6732,N_6741);
nand U6925 (N_6925,N_6772,N_6774);
or U6926 (N_6926,N_6620,N_6718);
nand U6927 (N_6927,N_6626,N_6623);
nor U6928 (N_6928,N_6754,N_6779);
and U6929 (N_6929,N_6643,N_6682);
nand U6930 (N_6930,N_6617,N_6746);
and U6931 (N_6931,N_6664,N_6770);
nor U6932 (N_6932,N_6667,N_6633);
nor U6933 (N_6933,N_6604,N_6761);
or U6934 (N_6934,N_6720,N_6717);
nor U6935 (N_6935,N_6785,N_6612);
nor U6936 (N_6936,N_6734,N_6614);
nand U6937 (N_6937,N_6656,N_6748);
nor U6938 (N_6938,N_6696,N_6610);
and U6939 (N_6939,N_6685,N_6677);
or U6940 (N_6940,N_6675,N_6627);
nand U6941 (N_6941,N_6628,N_6718);
nand U6942 (N_6942,N_6614,N_6778);
or U6943 (N_6943,N_6690,N_6650);
and U6944 (N_6944,N_6790,N_6799);
or U6945 (N_6945,N_6727,N_6766);
nand U6946 (N_6946,N_6769,N_6774);
xnor U6947 (N_6947,N_6651,N_6749);
and U6948 (N_6948,N_6774,N_6701);
or U6949 (N_6949,N_6781,N_6722);
nand U6950 (N_6950,N_6662,N_6654);
or U6951 (N_6951,N_6672,N_6780);
and U6952 (N_6952,N_6640,N_6777);
nor U6953 (N_6953,N_6756,N_6650);
and U6954 (N_6954,N_6716,N_6773);
nor U6955 (N_6955,N_6686,N_6765);
and U6956 (N_6956,N_6721,N_6708);
nand U6957 (N_6957,N_6727,N_6624);
nor U6958 (N_6958,N_6664,N_6737);
nand U6959 (N_6959,N_6633,N_6713);
nor U6960 (N_6960,N_6783,N_6611);
and U6961 (N_6961,N_6737,N_6622);
and U6962 (N_6962,N_6753,N_6655);
nand U6963 (N_6963,N_6682,N_6606);
and U6964 (N_6964,N_6769,N_6739);
nand U6965 (N_6965,N_6601,N_6609);
nand U6966 (N_6966,N_6759,N_6772);
nor U6967 (N_6967,N_6600,N_6639);
and U6968 (N_6968,N_6796,N_6785);
and U6969 (N_6969,N_6760,N_6749);
and U6970 (N_6970,N_6607,N_6685);
and U6971 (N_6971,N_6708,N_6733);
and U6972 (N_6972,N_6713,N_6765);
nor U6973 (N_6973,N_6736,N_6745);
nor U6974 (N_6974,N_6724,N_6619);
or U6975 (N_6975,N_6672,N_6619);
nand U6976 (N_6976,N_6659,N_6617);
or U6977 (N_6977,N_6609,N_6700);
or U6978 (N_6978,N_6698,N_6631);
nand U6979 (N_6979,N_6669,N_6746);
nand U6980 (N_6980,N_6690,N_6738);
nand U6981 (N_6981,N_6723,N_6628);
nor U6982 (N_6982,N_6671,N_6658);
and U6983 (N_6983,N_6638,N_6609);
nor U6984 (N_6984,N_6689,N_6600);
xor U6985 (N_6985,N_6603,N_6661);
nor U6986 (N_6986,N_6751,N_6750);
and U6987 (N_6987,N_6774,N_6775);
nor U6988 (N_6988,N_6789,N_6686);
or U6989 (N_6989,N_6755,N_6754);
nand U6990 (N_6990,N_6767,N_6715);
or U6991 (N_6991,N_6687,N_6673);
nand U6992 (N_6992,N_6641,N_6658);
and U6993 (N_6993,N_6734,N_6666);
nand U6994 (N_6994,N_6760,N_6717);
nand U6995 (N_6995,N_6618,N_6740);
nand U6996 (N_6996,N_6664,N_6660);
xor U6997 (N_6997,N_6730,N_6721);
and U6998 (N_6998,N_6795,N_6717);
nand U6999 (N_6999,N_6787,N_6639);
nor U7000 (N_7000,N_6820,N_6832);
nor U7001 (N_7001,N_6887,N_6828);
nor U7002 (N_7002,N_6998,N_6957);
nor U7003 (N_7003,N_6804,N_6980);
nor U7004 (N_7004,N_6912,N_6894);
xor U7005 (N_7005,N_6961,N_6837);
nor U7006 (N_7006,N_6802,N_6862);
and U7007 (N_7007,N_6928,N_6945);
and U7008 (N_7008,N_6874,N_6885);
nor U7009 (N_7009,N_6911,N_6906);
and U7010 (N_7010,N_6934,N_6960);
and U7011 (N_7011,N_6863,N_6949);
or U7012 (N_7012,N_6896,N_6989);
nand U7013 (N_7013,N_6923,N_6839);
and U7014 (N_7014,N_6956,N_6806);
and U7015 (N_7015,N_6801,N_6965);
nor U7016 (N_7016,N_6946,N_6877);
and U7017 (N_7017,N_6898,N_6937);
nor U7018 (N_7018,N_6947,N_6924);
xnor U7019 (N_7019,N_6975,N_6979);
nand U7020 (N_7020,N_6959,N_6833);
nand U7021 (N_7021,N_6994,N_6856);
and U7022 (N_7022,N_6978,N_6859);
and U7023 (N_7023,N_6963,N_6992);
nand U7024 (N_7024,N_6902,N_6890);
xor U7025 (N_7025,N_6880,N_6852);
and U7026 (N_7026,N_6920,N_6861);
nand U7027 (N_7027,N_6884,N_6931);
and U7028 (N_7028,N_6930,N_6952);
or U7029 (N_7029,N_6929,N_6846);
nand U7030 (N_7030,N_6855,N_6803);
nand U7031 (N_7031,N_6908,N_6933);
and U7032 (N_7032,N_6809,N_6962);
and U7033 (N_7033,N_6909,N_6985);
and U7034 (N_7034,N_6973,N_6891);
or U7035 (N_7035,N_6834,N_6871);
nand U7036 (N_7036,N_6948,N_6981);
nand U7037 (N_7037,N_6927,N_6984);
and U7038 (N_7038,N_6827,N_6950);
and U7039 (N_7039,N_6977,N_6889);
nor U7040 (N_7040,N_6996,N_6893);
xor U7041 (N_7041,N_6917,N_6907);
and U7042 (N_7042,N_6849,N_6899);
nor U7043 (N_7043,N_6810,N_6905);
nor U7044 (N_7044,N_6897,N_6919);
nand U7045 (N_7045,N_6858,N_6910);
nand U7046 (N_7046,N_6972,N_6967);
xor U7047 (N_7047,N_6903,N_6811);
and U7048 (N_7048,N_6879,N_6817);
nor U7049 (N_7049,N_6875,N_6938);
nor U7050 (N_7050,N_6999,N_6940);
nand U7051 (N_7051,N_6819,N_6976);
and U7052 (N_7052,N_6869,N_6857);
and U7053 (N_7053,N_6883,N_6816);
nor U7054 (N_7054,N_6860,N_6822);
nor U7055 (N_7055,N_6850,N_6926);
and U7056 (N_7056,N_6824,N_6921);
and U7057 (N_7057,N_6966,N_6969);
or U7058 (N_7058,N_6873,N_6932);
nand U7059 (N_7059,N_6821,N_6993);
or U7060 (N_7060,N_6870,N_6955);
nand U7061 (N_7061,N_6851,N_6953);
and U7062 (N_7062,N_6971,N_6968);
or U7063 (N_7063,N_6882,N_6925);
nand U7064 (N_7064,N_6941,N_6892);
xor U7065 (N_7065,N_6844,N_6922);
and U7066 (N_7066,N_6835,N_6853);
or U7067 (N_7067,N_6830,N_6991);
and U7068 (N_7068,N_6954,N_6826);
and U7069 (N_7069,N_6800,N_6836);
and U7070 (N_7070,N_6807,N_6866);
and U7071 (N_7071,N_6868,N_6838);
nand U7072 (N_7072,N_6808,N_6990);
nor U7073 (N_7073,N_6995,N_6916);
xnor U7074 (N_7074,N_6895,N_6914);
nor U7075 (N_7075,N_6878,N_6904);
nor U7076 (N_7076,N_6951,N_6841);
and U7077 (N_7077,N_6854,N_6983);
and U7078 (N_7078,N_6939,N_6936);
and U7079 (N_7079,N_6901,N_6813);
and U7080 (N_7080,N_6943,N_6815);
or U7081 (N_7081,N_6829,N_6843);
nor U7082 (N_7082,N_6900,N_6823);
or U7083 (N_7083,N_6812,N_6944);
nand U7084 (N_7084,N_6867,N_6864);
nor U7085 (N_7085,N_6986,N_6818);
nor U7086 (N_7086,N_6913,N_6970);
and U7087 (N_7087,N_6935,N_6848);
xor U7088 (N_7088,N_6840,N_6982);
nor U7089 (N_7089,N_6842,N_6845);
nor U7090 (N_7090,N_6958,N_6888);
or U7091 (N_7091,N_6988,N_6831);
nand U7092 (N_7092,N_6881,N_6915);
or U7093 (N_7093,N_6847,N_6872);
or U7094 (N_7094,N_6918,N_6865);
or U7095 (N_7095,N_6805,N_6886);
or U7096 (N_7096,N_6964,N_6997);
nor U7097 (N_7097,N_6974,N_6942);
or U7098 (N_7098,N_6814,N_6876);
or U7099 (N_7099,N_6987,N_6825);
or U7100 (N_7100,N_6815,N_6929);
and U7101 (N_7101,N_6897,N_6970);
or U7102 (N_7102,N_6966,N_6813);
or U7103 (N_7103,N_6844,N_6960);
or U7104 (N_7104,N_6958,N_6831);
and U7105 (N_7105,N_6889,N_6863);
and U7106 (N_7106,N_6850,N_6858);
and U7107 (N_7107,N_6863,N_6851);
and U7108 (N_7108,N_6805,N_6828);
and U7109 (N_7109,N_6904,N_6892);
nor U7110 (N_7110,N_6930,N_6845);
and U7111 (N_7111,N_6980,N_6928);
and U7112 (N_7112,N_6998,N_6999);
nand U7113 (N_7113,N_6871,N_6936);
xnor U7114 (N_7114,N_6891,N_6812);
nand U7115 (N_7115,N_6864,N_6909);
and U7116 (N_7116,N_6892,N_6999);
and U7117 (N_7117,N_6939,N_6863);
nand U7118 (N_7118,N_6876,N_6922);
and U7119 (N_7119,N_6846,N_6854);
nand U7120 (N_7120,N_6909,N_6937);
or U7121 (N_7121,N_6959,N_6840);
nor U7122 (N_7122,N_6811,N_6972);
nor U7123 (N_7123,N_6880,N_6803);
nor U7124 (N_7124,N_6998,N_6972);
nor U7125 (N_7125,N_6863,N_6874);
and U7126 (N_7126,N_6905,N_6840);
and U7127 (N_7127,N_6981,N_6964);
and U7128 (N_7128,N_6886,N_6957);
nor U7129 (N_7129,N_6911,N_6872);
nor U7130 (N_7130,N_6992,N_6805);
and U7131 (N_7131,N_6854,N_6973);
or U7132 (N_7132,N_6859,N_6842);
xor U7133 (N_7133,N_6997,N_6956);
or U7134 (N_7134,N_6953,N_6868);
and U7135 (N_7135,N_6916,N_6859);
or U7136 (N_7136,N_6824,N_6846);
or U7137 (N_7137,N_6847,N_6890);
or U7138 (N_7138,N_6937,N_6976);
nand U7139 (N_7139,N_6850,N_6826);
and U7140 (N_7140,N_6993,N_6851);
and U7141 (N_7141,N_6875,N_6892);
nand U7142 (N_7142,N_6802,N_6822);
and U7143 (N_7143,N_6940,N_6838);
xnor U7144 (N_7144,N_6814,N_6931);
and U7145 (N_7145,N_6906,N_6883);
or U7146 (N_7146,N_6961,N_6844);
or U7147 (N_7147,N_6943,N_6892);
xor U7148 (N_7148,N_6808,N_6944);
and U7149 (N_7149,N_6998,N_6870);
nor U7150 (N_7150,N_6918,N_6927);
nor U7151 (N_7151,N_6939,N_6814);
and U7152 (N_7152,N_6926,N_6925);
nor U7153 (N_7153,N_6972,N_6827);
nor U7154 (N_7154,N_6858,N_6958);
nor U7155 (N_7155,N_6820,N_6965);
nand U7156 (N_7156,N_6809,N_6876);
or U7157 (N_7157,N_6807,N_6926);
and U7158 (N_7158,N_6936,N_6822);
nor U7159 (N_7159,N_6918,N_6871);
or U7160 (N_7160,N_6847,N_6954);
or U7161 (N_7161,N_6969,N_6834);
or U7162 (N_7162,N_6894,N_6968);
and U7163 (N_7163,N_6937,N_6811);
and U7164 (N_7164,N_6962,N_6980);
or U7165 (N_7165,N_6819,N_6860);
nor U7166 (N_7166,N_6880,N_6941);
nor U7167 (N_7167,N_6870,N_6952);
xor U7168 (N_7168,N_6962,N_6858);
or U7169 (N_7169,N_6942,N_6957);
nand U7170 (N_7170,N_6947,N_6818);
or U7171 (N_7171,N_6997,N_6880);
nor U7172 (N_7172,N_6974,N_6937);
nor U7173 (N_7173,N_6890,N_6989);
nor U7174 (N_7174,N_6806,N_6947);
nand U7175 (N_7175,N_6857,N_6999);
nor U7176 (N_7176,N_6984,N_6866);
nand U7177 (N_7177,N_6912,N_6988);
and U7178 (N_7178,N_6885,N_6928);
or U7179 (N_7179,N_6888,N_6811);
xor U7180 (N_7180,N_6932,N_6824);
nand U7181 (N_7181,N_6940,N_6957);
and U7182 (N_7182,N_6904,N_6959);
nand U7183 (N_7183,N_6881,N_6853);
nand U7184 (N_7184,N_6874,N_6929);
nor U7185 (N_7185,N_6953,N_6882);
and U7186 (N_7186,N_6910,N_6843);
xnor U7187 (N_7187,N_6842,N_6817);
and U7188 (N_7188,N_6981,N_6889);
or U7189 (N_7189,N_6899,N_6978);
nor U7190 (N_7190,N_6992,N_6946);
and U7191 (N_7191,N_6876,N_6842);
or U7192 (N_7192,N_6983,N_6803);
or U7193 (N_7193,N_6901,N_6818);
nor U7194 (N_7194,N_6867,N_6909);
nor U7195 (N_7195,N_6902,N_6892);
and U7196 (N_7196,N_6999,N_6894);
or U7197 (N_7197,N_6924,N_6985);
xor U7198 (N_7198,N_6999,N_6943);
or U7199 (N_7199,N_6842,N_6899);
or U7200 (N_7200,N_7162,N_7096);
nand U7201 (N_7201,N_7045,N_7193);
nor U7202 (N_7202,N_7059,N_7122);
or U7203 (N_7203,N_7011,N_7126);
nand U7204 (N_7204,N_7074,N_7104);
or U7205 (N_7205,N_7119,N_7189);
nor U7206 (N_7206,N_7026,N_7056);
or U7207 (N_7207,N_7057,N_7155);
and U7208 (N_7208,N_7014,N_7060);
and U7209 (N_7209,N_7049,N_7144);
and U7210 (N_7210,N_7108,N_7164);
or U7211 (N_7211,N_7010,N_7156);
xor U7212 (N_7212,N_7152,N_7033);
or U7213 (N_7213,N_7158,N_7079);
and U7214 (N_7214,N_7041,N_7130);
and U7215 (N_7215,N_7025,N_7186);
and U7216 (N_7216,N_7006,N_7116);
or U7217 (N_7217,N_7168,N_7191);
and U7218 (N_7218,N_7050,N_7197);
or U7219 (N_7219,N_7029,N_7118);
or U7220 (N_7220,N_7019,N_7039);
and U7221 (N_7221,N_7024,N_7035);
or U7222 (N_7222,N_7027,N_7080);
or U7223 (N_7223,N_7146,N_7157);
or U7224 (N_7224,N_7196,N_7051);
nor U7225 (N_7225,N_7135,N_7117);
xnor U7226 (N_7226,N_7183,N_7061);
and U7227 (N_7227,N_7038,N_7034);
and U7228 (N_7228,N_7175,N_7100);
nor U7229 (N_7229,N_7013,N_7136);
nand U7230 (N_7230,N_7112,N_7007);
and U7231 (N_7231,N_7170,N_7048);
or U7232 (N_7232,N_7173,N_7022);
nor U7233 (N_7233,N_7052,N_7166);
nor U7234 (N_7234,N_7181,N_7005);
or U7235 (N_7235,N_7141,N_7092);
nor U7236 (N_7236,N_7192,N_7169);
and U7237 (N_7237,N_7111,N_7184);
nand U7238 (N_7238,N_7180,N_7160);
nand U7239 (N_7239,N_7083,N_7081);
nor U7240 (N_7240,N_7124,N_7161);
nand U7241 (N_7241,N_7091,N_7132);
nor U7242 (N_7242,N_7138,N_7154);
and U7243 (N_7243,N_7084,N_7077);
nor U7244 (N_7244,N_7176,N_7128);
nor U7245 (N_7245,N_7190,N_7106);
or U7246 (N_7246,N_7198,N_7020);
nor U7247 (N_7247,N_7031,N_7076);
xor U7248 (N_7248,N_7115,N_7103);
nand U7249 (N_7249,N_7093,N_7127);
nor U7250 (N_7250,N_7054,N_7167);
nand U7251 (N_7251,N_7105,N_7070);
nand U7252 (N_7252,N_7174,N_7075);
or U7253 (N_7253,N_7171,N_7037);
nor U7254 (N_7254,N_7008,N_7047);
xor U7255 (N_7255,N_7133,N_7012);
and U7256 (N_7256,N_7015,N_7134);
nand U7257 (N_7257,N_7067,N_7032);
and U7258 (N_7258,N_7131,N_7194);
or U7259 (N_7259,N_7064,N_7165);
and U7260 (N_7260,N_7109,N_7107);
nor U7261 (N_7261,N_7040,N_7142);
nor U7262 (N_7262,N_7101,N_7016);
nor U7263 (N_7263,N_7098,N_7086);
nor U7264 (N_7264,N_7095,N_7090);
nor U7265 (N_7265,N_7082,N_7018);
and U7266 (N_7266,N_7187,N_7046);
nor U7267 (N_7267,N_7143,N_7072);
or U7268 (N_7268,N_7121,N_7042);
nor U7269 (N_7269,N_7178,N_7028);
and U7270 (N_7270,N_7159,N_7129);
nand U7271 (N_7271,N_7087,N_7137);
xnor U7272 (N_7272,N_7078,N_7185);
or U7273 (N_7273,N_7088,N_7068);
nand U7274 (N_7274,N_7179,N_7120);
xnor U7275 (N_7275,N_7140,N_7055);
or U7276 (N_7276,N_7113,N_7114);
nand U7277 (N_7277,N_7110,N_7125);
or U7278 (N_7278,N_7199,N_7001);
and U7279 (N_7279,N_7188,N_7085);
and U7280 (N_7280,N_7062,N_7151);
or U7281 (N_7281,N_7145,N_7066);
and U7282 (N_7282,N_7139,N_7073);
or U7283 (N_7283,N_7147,N_7004);
nand U7284 (N_7284,N_7044,N_7094);
and U7285 (N_7285,N_7053,N_7063);
nand U7286 (N_7286,N_7009,N_7058);
nand U7287 (N_7287,N_7099,N_7002);
nor U7288 (N_7288,N_7102,N_7003);
xnor U7289 (N_7289,N_7153,N_7021);
nand U7290 (N_7290,N_7163,N_7065);
and U7291 (N_7291,N_7043,N_7150);
and U7292 (N_7292,N_7195,N_7177);
nor U7293 (N_7293,N_7089,N_7069);
or U7294 (N_7294,N_7036,N_7017);
and U7295 (N_7295,N_7148,N_7071);
and U7296 (N_7296,N_7172,N_7149);
nand U7297 (N_7297,N_7000,N_7023);
nand U7298 (N_7298,N_7030,N_7123);
or U7299 (N_7299,N_7182,N_7097);
nor U7300 (N_7300,N_7192,N_7131);
nand U7301 (N_7301,N_7062,N_7190);
or U7302 (N_7302,N_7031,N_7174);
nand U7303 (N_7303,N_7094,N_7173);
or U7304 (N_7304,N_7030,N_7059);
and U7305 (N_7305,N_7144,N_7189);
nand U7306 (N_7306,N_7188,N_7184);
xnor U7307 (N_7307,N_7000,N_7147);
and U7308 (N_7308,N_7103,N_7114);
xor U7309 (N_7309,N_7148,N_7163);
and U7310 (N_7310,N_7101,N_7193);
and U7311 (N_7311,N_7173,N_7187);
and U7312 (N_7312,N_7194,N_7144);
nand U7313 (N_7313,N_7043,N_7125);
xnor U7314 (N_7314,N_7164,N_7014);
or U7315 (N_7315,N_7075,N_7114);
and U7316 (N_7316,N_7191,N_7184);
and U7317 (N_7317,N_7060,N_7022);
nor U7318 (N_7318,N_7000,N_7112);
nand U7319 (N_7319,N_7100,N_7034);
nand U7320 (N_7320,N_7168,N_7087);
xor U7321 (N_7321,N_7094,N_7140);
or U7322 (N_7322,N_7046,N_7161);
nand U7323 (N_7323,N_7137,N_7101);
and U7324 (N_7324,N_7003,N_7103);
or U7325 (N_7325,N_7157,N_7075);
nor U7326 (N_7326,N_7014,N_7071);
nand U7327 (N_7327,N_7045,N_7188);
or U7328 (N_7328,N_7014,N_7052);
xnor U7329 (N_7329,N_7005,N_7039);
nand U7330 (N_7330,N_7194,N_7161);
or U7331 (N_7331,N_7009,N_7079);
xnor U7332 (N_7332,N_7151,N_7191);
nand U7333 (N_7333,N_7129,N_7047);
or U7334 (N_7334,N_7012,N_7005);
nand U7335 (N_7335,N_7141,N_7164);
xor U7336 (N_7336,N_7166,N_7049);
xnor U7337 (N_7337,N_7151,N_7063);
nor U7338 (N_7338,N_7159,N_7110);
xor U7339 (N_7339,N_7013,N_7027);
or U7340 (N_7340,N_7133,N_7155);
nand U7341 (N_7341,N_7063,N_7190);
or U7342 (N_7342,N_7161,N_7148);
or U7343 (N_7343,N_7062,N_7050);
and U7344 (N_7344,N_7099,N_7057);
or U7345 (N_7345,N_7125,N_7189);
nor U7346 (N_7346,N_7073,N_7002);
or U7347 (N_7347,N_7027,N_7147);
nor U7348 (N_7348,N_7191,N_7117);
or U7349 (N_7349,N_7175,N_7012);
nor U7350 (N_7350,N_7021,N_7099);
nor U7351 (N_7351,N_7094,N_7003);
xor U7352 (N_7352,N_7187,N_7010);
and U7353 (N_7353,N_7052,N_7092);
xor U7354 (N_7354,N_7108,N_7062);
nand U7355 (N_7355,N_7099,N_7190);
nand U7356 (N_7356,N_7039,N_7061);
nor U7357 (N_7357,N_7082,N_7061);
nor U7358 (N_7358,N_7056,N_7149);
and U7359 (N_7359,N_7061,N_7193);
and U7360 (N_7360,N_7032,N_7131);
or U7361 (N_7361,N_7122,N_7176);
and U7362 (N_7362,N_7150,N_7074);
nor U7363 (N_7363,N_7197,N_7110);
nor U7364 (N_7364,N_7081,N_7054);
nor U7365 (N_7365,N_7056,N_7034);
and U7366 (N_7366,N_7199,N_7180);
nor U7367 (N_7367,N_7179,N_7047);
and U7368 (N_7368,N_7004,N_7087);
and U7369 (N_7369,N_7044,N_7088);
nand U7370 (N_7370,N_7079,N_7086);
or U7371 (N_7371,N_7079,N_7168);
nand U7372 (N_7372,N_7134,N_7147);
nand U7373 (N_7373,N_7166,N_7151);
nand U7374 (N_7374,N_7142,N_7058);
and U7375 (N_7375,N_7166,N_7013);
or U7376 (N_7376,N_7086,N_7096);
or U7377 (N_7377,N_7145,N_7012);
nand U7378 (N_7378,N_7166,N_7118);
nor U7379 (N_7379,N_7188,N_7148);
nand U7380 (N_7380,N_7042,N_7159);
nand U7381 (N_7381,N_7154,N_7130);
and U7382 (N_7382,N_7177,N_7064);
and U7383 (N_7383,N_7156,N_7020);
nand U7384 (N_7384,N_7040,N_7056);
and U7385 (N_7385,N_7187,N_7124);
nand U7386 (N_7386,N_7094,N_7040);
nand U7387 (N_7387,N_7159,N_7000);
xor U7388 (N_7388,N_7094,N_7121);
or U7389 (N_7389,N_7097,N_7156);
nor U7390 (N_7390,N_7059,N_7191);
and U7391 (N_7391,N_7080,N_7099);
xor U7392 (N_7392,N_7094,N_7123);
xnor U7393 (N_7393,N_7104,N_7008);
nand U7394 (N_7394,N_7048,N_7065);
and U7395 (N_7395,N_7092,N_7169);
or U7396 (N_7396,N_7161,N_7198);
xnor U7397 (N_7397,N_7125,N_7176);
nor U7398 (N_7398,N_7099,N_7079);
nor U7399 (N_7399,N_7026,N_7067);
and U7400 (N_7400,N_7266,N_7303);
nor U7401 (N_7401,N_7362,N_7263);
nor U7402 (N_7402,N_7357,N_7331);
nor U7403 (N_7403,N_7341,N_7214);
nor U7404 (N_7404,N_7308,N_7296);
and U7405 (N_7405,N_7227,N_7345);
nand U7406 (N_7406,N_7369,N_7200);
or U7407 (N_7407,N_7238,N_7229);
nor U7408 (N_7408,N_7342,N_7203);
nor U7409 (N_7409,N_7247,N_7340);
nor U7410 (N_7410,N_7212,N_7209);
and U7411 (N_7411,N_7318,N_7388);
and U7412 (N_7412,N_7211,N_7311);
xnor U7413 (N_7413,N_7251,N_7333);
and U7414 (N_7414,N_7268,N_7233);
nand U7415 (N_7415,N_7363,N_7330);
nor U7416 (N_7416,N_7280,N_7348);
or U7417 (N_7417,N_7294,N_7383);
nand U7418 (N_7418,N_7306,N_7304);
xnor U7419 (N_7419,N_7325,N_7248);
or U7420 (N_7420,N_7213,N_7314);
and U7421 (N_7421,N_7287,N_7354);
and U7422 (N_7422,N_7335,N_7242);
xnor U7423 (N_7423,N_7290,N_7313);
nor U7424 (N_7424,N_7360,N_7270);
and U7425 (N_7425,N_7275,N_7288);
and U7426 (N_7426,N_7225,N_7201);
and U7427 (N_7427,N_7334,N_7373);
or U7428 (N_7428,N_7206,N_7385);
nor U7429 (N_7429,N_7259,N_7312);
nand U7430 (N_7430,N_7255,N_7315);
nor U7431 (N_7431,N_7283,N_7220);
or U7432 (N_7432,N_7396,N_7202);
and U7433 (N_7433,N_7232,N_7208);
and U7434 (N_7434,N_7337,N_7274);
and U7435 (N_7435,N_7349,N_7323);
and U7436 (N_7436,N_7299,N_7395);
nor U7437 (N_7437,N_7307,N_7278);
and U7438 (N_7438,N_7376,N_7366);
and U7439 (N_7439,N_7257,N_7240);
nand U7440 (N_7440,N_7228,N_7398);
and U7441 (N_7441,N_7361,N_7368);
or U7442 (N_7442,N_7320,N_7339);
nor U7443 (N_7443,N_7355,N_7205);
nand U7444 (N_7444,N_7316,N_7321);
or U7445 (N_7445,N_7298,N_7352);
nand U7446 (N_7446,N_7264,N_7353);
nor U7447 (N_7447,N_7358,N_7351);
and U7448 (N_7448,N_7281,N_7324);
nor U7449 (N_7449,N_7231,N_7262);
nand U7450 (N_7450,N_7300,N_7319);
or U7451 (N_7451,N_7365,N_7332);
nor U7452 (N_7452,N_7347,N_7356);
and U7453 (N_7453,N_7336,N_7344);
nand U7454 (N_7454,N_7261,N_7279);
xor U7455 (N_7455,N_7389,N_7387);
or U7456 (N_7456,N_7260,N_7217);
nand U7457 (N_7457,N_7381,N_7230);
nand U7458 (N_7458,N_7236,N_7284);
nor U7459 (N_7459,N_7272,N_7273);
nand U7460 (N_7460,N_7219,N_7397);
xor U7461 (N_7461,N_7377,N_7293);
nand U7462 (N_7462,N_7292,N_7329);
nor U7463 (N_7463,N_7245,N_7394);
or U7464 (N_7464,N_7223,N_7380);
xnor U7465 (N_7465,N_7301,N_7327);
and U7466 (N_7466,N_7374,N_7224);
nand U7467 (N_7467,N_7254,N_7267);
nor U7468 (N_7468,N_7309,N_7244);
or U7469 (N_7469,N_7250,N_7322);
or U7470 (N_7470,N_7221,N_7215);
and U7471 (N_7471,N_7391,N_7317);
or U7472 (N_7472,N_7285,N_7359);
nor U7473 (N_7473,N_7338,N_7234);
or U7474 (N_7474,N_7297,N_7364);
nand U7475 (N_7475,N_7269,N_7343);
nor U7476 (N_7476,N_7204,N_7286);
nand U7477 (N_7477,N_7271,N_7379);
nor U7478 (N_7478,N_7222,N_7390);
nor U7479 (N_7479,N_7258,N_7295);
and U7480 (N_7480,N_7239,N_7226);
and U7481 (N_7481,N_7382,N_7328);
or U7482 (N_7482,N_7371,N_7378);
and U7483 (N_7483,N_7277,N_7302);
xor U7484 (N_7484,N_7392,N_7249);
and U7485 (N_7485,N_7375,N_7210);
xor U7486 (N_7486,N_7289,N_7393);
nand U7487 (N_7487,N_7326,N_7256);
nor U7488 (N_7488,N_7367,N_7305);
nor U7489 (N_7489,N_7291,N_7253);
or U7490 (N_7490,N_7310,N_7399);
and U7491 (N_7491,N_7346,N_7370);
xnor U7492 (N_7492,N_7372,N_7218);
nor U7493 (N_7493,N_7276,N_7237);
nor U7494 (N_7494,N_7386,N_7282);
xor U7495 (N_7495,N_7235,N_7246);
nor U7496 (N_7496,N_7384,N_7241);
and U7497 (N_7497,N_7350,N_7207);
nand U7498 (N_7498,N_7265,N_7252);
nor U7499 (N_7499,N_7216,N_7243);
and U7500 (N_7500,N_7351,N_7219);
or U7501 (N_7501,N_7366,N_7396);
nand U7502 (N_7502,N_7307,N_7329);
nor U7503 (N_7503,N_7318,N_7251);
xor U7504 (N_7504,N_7332,N_7341);
and U7505 (N_7505,N_7353,N_7246);
nor U7506 (N_7506,N_7258,N_7280);
nand U7507 (N_7507,N_7351,N_7313);
nand U7508 (N_7508,N_7391,N_7316);
xor U7509 (N_7509,N_7386,N_7382);
or U7510 (N_7510,N_7246,N_7339);
or U7511 (N_7511,N_7234,N_7265);
and U7512 (N_7512,N_7219,N_7262);
and U7513 (N_7513,N_7272,N_7353);
or U7514 (N_7514,N_7369,N_7242);
nor U7515 (N_7515,N_7285,N_7382);
nand U7516 (N_7516,N_7353,N_7370);
nand U7517 (N_7517,N_7377,N_7216);
nand U7518 (N_7518,N_7368,N_7260);
xnor U7519 (N_7519,N_7334,N_7348);
nand U7520 (N_7520,N_7309,N_7200);
nand U7521 (N_7521,N_7225,N_7370);
and U7522 (N_7522,N_7302,N_7279);
or U7523 (N_7523,N_7256,N_7368);
nand U7524 (N_7524,N_7234,N_7376);
and U7525 (N_7525,N_7279,N_7272);
nor U7526 (N_7526,N_7277,N_7293);
and U7527 (N_7527,N_7255,N_7286);
nor U7528 (N_7528,N_7282,N_7396);
and U7529 (N_7529,N_7298,N_7335);
nand U7530 (N_7530,N_7222,N_7339);
and U7531 (N_7531,N_7203,N_7371);
and U7532 (N_7532,N_7251,N_7283);
and U7533 (N_7533,N_7217,N_7305);
or U7534 (N_7534,N_7354,N_7398);
and U7535 (N_7535,N_7327,N_7233);
nand U7536 (N_7536,N_7322,N_7371);
nand U7537 (N_7537,N_7243,N_7306);
and U7538 (N_7538,N_7226,N_7377);
nor U7539 (N_7539,N_7303,N_7261);
or U7540 (N_7540,N_7289,N_7251);
and U7541 (N_7541,N_7213,N_7396);
and U7542 (N_7542,N_7247,N_7390);
nand U7543 (N_7543,N_7279,N_7227);
nand U7544 (N_7544,N_7326,N_7272);
or U7545 (N_7545,N_7202,N_7341);
and U7546 (N_7546,N_7313,N_7267);
nor U7547 (N_7547,N_7206,N_7306);
xor U7548 (N_7548,N_7328,N_7268);
nor U7549 (N_7549,N_7270,N_7387);
or U7550 (N_7550,N_7287,N_7363);
nand U7551 (N_7551,N_7314,N_7396);
nand U7552 (N_7552,N_7282,N_7373);
nor U7553 (N_7553,N_7340,N_7252);
and U7554 (N_7554,N_7230,N_7390);
nor U7555 (N_7555,N_7258,N_7218);
and U7556 (N_7556,N_7243,N_7248);
nand U7557 (N_7557,N_7327,N_7345);
or U7558 (N_7558,N_7319,N_7331);
xor U7559 (N_7559,N_7214,N_7228);
nor U7560 (N_7560,N_7388,N_7337);
and U7561 (N_7561,N_7311,N_7206);
xor U7562 (N_7562,N_7320,N_7307);
xor U7563 (N_7563,N_7310,N_7360);
or U7564 (N_7564,N_7237,N_7225);
xor U7565 (N_7565,N_7233,N_7325);
and U7566 (N_7566,N_7380,N_7377);
and U7567 (N_7567,N_7298,N_7394);
and U7568 (N_7568,N_7325,N_7384);
and U7569 (N_7569,N_7297,N_7263);
or U7570 (N_7570,N_7245,N_7226);
nand U7571 (N_7571,N_7382,N_7215);
and U7572 (N_7572,N_7335,N_7293);
and U7573 (N_7573,N_7313,N_7367);
or U7574 (N_7574,N_7375,N_7356);
nand U7575 (N_7575,N_7318,N_7222);
or U7576 (N_7576,N_7399,N_7220);
and U7577 (N_7577,N_7359,N_7208);
or U7578 (N_7578,N_7303,N_7231);
or U7579 (N_7579,N_7387,N_7372);
xnor U7580 (N_7580,N_7235,N_7354);
nor U7581 (N_7581,N_7296,N_7399);
xor U7582 (N_7582,N_7211,N_7308);
nand U7583 (N_7583,N_7392,N_7298);
nand U7584 (N_7584,N_7262,N_7396);
nor U7585 (N_7585,N_7294,N_7395);
or U7586 (N_7586,N_7306,N_7238);
nor U7587 (N_7587,N_7329,N_7328);
or U7588 (N_7588,N_7348,N_7360);
nor U7589 (N_7589,N_7223,N_7348);
nor U7590 (N_7590,N_7283,N_7369);
nand U7591 (N_7591,N_7213,N_7370);
and U7592 (N_7592,N_7287,N_7267);
and U7593 (N_7593,N_7361,N_7231);
nor U7594 (N_7594,N_7352,N_7287);
xnor U7595 (N_7595,N_7331,N_7250);
nor U7596 (N_7596,N_7229,N_7286);
nand U7597 (N_7597,N_7236,N_7359);
or U7598 (N_7598,N_7390,N_7278);
nand U7599 (N_7599,N_7366,N_7284);
nor U7600 (N_7600,N_7441,N_7473);
and U7601 (N_7601,N_7436,N_7546);
nor U7602 (N_7602,N_7467,N_7533);
or U7603 (N_7603,N_7503,N_7404);
and U7604 (N_7604,N_7478,N_7402);
and U7605 (N_7605,N_7554,N_7418);
xor U7606 (N_7606,N_7574,N_7472);
or U7607 (N_7607,N_7568,N_7437);
nand U7608 (N_7608,N_7528,N_7460);
or U7609 (N_7609,N_7505,N_7515);
nand U7610 (N_7610,N_7576,N_7423);
and U7611 (N_7611,N_7541,N_7455);
and U7612 (N_7612,N_7484,N_7487);
nand U7613 (N_7613,N_7564,N_7491);
nor U7614 (N_7614,N_7483,N_7488);
nor U7615 (N_7615,N_7450,N_7562);
nor U7616 (N_7616,N_7531,N_7588);
and U7617 (N_7617,N_7536,N_7401);
and U7618 (N_7618,N_7407,N_7592);
or U7619 (N_7619,N_7500,N_7573);
nor U7620 (N_7620,N_7469,N_7465);
xor U7621 (N_7621,N_7525,N_7569);
nand U7622 (N_7622,N_7424,N_7405);
or U7623 (N_7623,N_7480,N_7558);
and U7624 (N_7624,N_7595,N_7501);
nor U7625 (N_7625,N_7583,N_7518);
and U7626 (N_7626,N_7477,N_7567);
nor U7627 (N_7627,N_7520,N_7449);
or U7628 (N_7628,N_7482,N_7445);
nor U7629 (N_7629,N_7556,N_7591);
nand U7630 (N_7630,N_7452,N_7542);
nor U7631 (N_7631,N_7414,N_7485);
nand U7632 (N_7632,N_7454,N_7590);
nand U7633 (N_7633,N_7585,N_7415);
nand U7634 (N_7634,N_7522,N_7470);
and U7635 (N_7635,N_7535,N_7411);
and U7636 (N_7636,N_7453,N_7462);
nor U7637 (N_7637,N_7559,N_7512);
or U7638 (N_7638,N_7519,N_7507);
xor U7639 (N_7639,N_7587,N_7502);
and U7640 (N_7640,N_7446,N_7563);
or U7641 (N_7641,N_7584,N_7527);
nand U7642 (N_7642,N_7526,N_7557);
and U7643 (N_7643,N_7457,N_7493);
or U7644 (N_7644,N_7517,N_7495);
and U7645 (N_7645,N_7551,N_7444);
or U7646 (N_7646,N_7596,N_7504);
and U7647 (N_7647,N_7476,N_7458);
or U7648 (N_7648,N_7499,N_7420);
nand U7649 (N_7649,N_7412,N_7413);
or U7650 (N_7650,N_7421,N_7432);
nand U7651 (N_7651,N_7430,N_7463);
xnor U7652 (N_7652,N_7428,N_7498);
and U7653 (N_7653,N_7425,N_7539);
nor U7654 (N_7654,N_7510,N_7534);
nor U7655 (N_7655,N_7494,N_7459);
nor U7656 (N_7656,N_7511,N_7464);
nor U7657 (N_7657,N_7581,N_7456);
nor U7658 (N_7658,N_7481,N_7417);
or U7659 (N_7659,N_7530,N_7597);
xor U7660 (N_7660,N_7489,N_7593);
and U7661 (N_7661,N_7406,N_7461);
or U7662 (N_7662,N_7426,N_7582);
or U7663 (N_7663,N_7543,N_7545);
nand U7664 (N_7664,N_7532,N_7516);
or U7665 (N_7665,N_7538,N_7442);
nor U7666 (N_7666,N_7466,N_7565);
nor U7667 (N_7667,N_7552,N_7550);
or U7668 (N_7668,N_7433,N_7408);
xnor U7669 (N_7669,N_7443,N_7553);
or U7670 (N_7670,N_7409,N_7429);
nor U7671 (N_7671,N_7447,N_7451);
nand U7672 (N_7672,N_7419,N_7410);
nor U7673 (N_7673,N_7594,N_7575);
nor U7674 (N_7674,N_7523,N_7561);
or U7675 (N_7675,N_7509,N_7589);
and U7676 (N_7676,N_7537,N_7547);
nand U7677 (N_7677,N_7403,N_7400);
nand U7678 (N_7678,N_7549,N_7416);
or U7679 (N_7679,N_7448,N_7566);
and U7680 (N_7680,N_7438,N_7580);
and U7681 (N_7681,N_7492,N_7578);
and U7682 (N_7682,N_7586,N_7471);
nand U7683 (N_7683,N_7434,N_7598);
nor U7684 (N_7684,N_7440,N_7514);
nand U7685 (N_7685,N_7435,N_7479);
nand U7686 (N_7686,N_7521,N_7529);
and U7687 (N_7687,N_7548,N_7474);
nor U7688 (N_7688,N_7599,N_7496);
and U7689 (N_7689,N_7497,N_7560);
and U7690 (N_7690,N_7513,N_7570);
or U7691 (N_7691,N_7540,N_7544);
and U7692 (N_7692,N_7486,N_7508);
nand U7693 (N_7693,N_7468,N_7439);
nand U7694 (N_7694,N_7555,N_7431);
nor U7695 (N_7695,N_7579,N_7524);
xnor U7696 (N_7696,N_7490,N_7506);
and U7697 (N_7697,N_7577,N_7427);
or U7698 (N_7698,N_7422,N_7475);
and U7699 (N_7699,N_7572,N_7571);
or U7700 (N_7700,N_7452,N_7539);
and U7701 (N_7701,N_7499,N_7440);
and U7702 (N_7702,N_7587,N_7565);
nor U7703 (N_7703,N_7518,N_7421);
or U7704 (N_7704,N_7406,N_7419);
nor U7705 (N_7705,N_7483,N_7416);
nor U7706 (N_7706,N_7427,N_7419);
nand U7707 (N_7707,N_7409,N_7593);
nand U7708 (N_7708,N_7542,N_7551);
nor U7709 (N_7709,N_7454,N_7478);
nor U7710 (N_7710,N_7410,N_7450);
nor U7711 (N_7711,N_7479,N_7513);
nor U7712 (N_7712,N_7463,N_7566);
nand U7713 (N_7713,N_7419,N_7566);
xor U7714 (N_7714,N_7587,N_7406);
and U7715 (N_7715,N_7538,N_7463);
nor U7716 (N_7716,N_7566,N_7477);
or U7717 (N_7717,N_7422,N_7531);
and U7718 (N_7718,N_7428,N_7504);
nor U7719 (N_7719,N_7547,N_7470);
or U7720 (N_7720,N_7515,N_7592);
and U7721 (N_7721,N_7429,N_7527);
and U7722 (N_7722,N_7489,N_7427);
and U7723 (N_7723,N_7492,N_7460);
xnor U7724 (N_7724,N_7443,N_7557);
and U7725 (N_7725,N_7554,N_7539);
or U7726 (N_7726,N_7450,N_7427);
nor U7727 (N_7727,N_7471,N_7561);
nor U7728 (N_7728,N_7479,N_7503);
nor U7729 (N_7729,N_7567,N_7456);
nand U7730 (N_7730,N_7574,N_7499);
nand U7731 (N_7731,N_7440,N_7565);
or U7732 (N_7732,N_7422,N_7528);
or U7733 (N_7733,N_7566,N_7451);
and U7734 (N_7734,N_7460,N_7537);
xor U7735 (N_7735,N_7504,N_7579);
and U7736 (N_7736,N_7452,N_7590);
nand U7737 (N_7737,N_7576,N_7556);
or U7738 (N_7738,N_7463,N_7516);
or U7739 (N_7739,N_7572,N_7495);
nor U7740 (N_7740,N_7488,N_7406);
nor U7741 (N_7741,N_7447,N_7519);
nor U7742 (N_7742,N_7593,N_7496);
nor U7743 (N_7743,N_7420,N_7562);
and U7744 (N_7744,N_7440,N_7534);
or U7745 (N_7745,N_7585,N_7566);
nor U7746 (N_7746,N_7478,N_7525);
and U7747 (N_7747,N_7528,N_7585);
nand U7748 (N_7748,N_7416,N_7491);
nor U7749 (N_7749,N_7485,N_7529);
and U7750 (N_7750,N_7501,N_7452);
and U7751 (N_7751,N_7588,N_7520);
nand U7752 (N_7752,N_7502,N_7518);
nor U7753 (N_7753,N_7430,N_7495);
and U7754 (N_7754,N_7557,N_7453);
nand U7755 (N_7755,N_7573,N_7436);
xor U7756 (N_7756,N_7564,N_7475);
nor U7757 (N_7757,N_7485,N_7442);
and U7758 (N_7758,N_7528,N_7586);
nor U7759 (N_7759,N_7411,N_7557);
nor U7760 (N_7760,N_7490,N_7412);
xor U7761 (N_7761,N_7426,N_7487);
and U7762 (N_7762,N_7452,N_7531);
nand U7763 (N_7763,N_7579,N_7588);
nand U7764 (N_7764,N_7572,N_7444);
nand U7765 (N_7765,N_7560,N_7574);
and U7766 (N_7766,N_7568,N_7560);
and U7767 (N_7767,N_7556,N_7474);
xnor U7768 (N_7768,N_7473,N_7458);
or U7769 (N_7769,N_7461,N_7538);
nand U7770 (N_7770,N_7416,N_7465);
nand U7771 (N_7771,N_7519,N_7546);
or U7772 (N_7772,N_7538,N_7425);
and U7773 (N_7773,N_7476,N_7435);
or U7774 (N_7774,N_7525,N_7403);
nor U7775 (N_7775,N_7518,N_7468);
xor U7776 (N_7776,N_7428,N_7588);
xnor U7777 (N_7777,N_7451,N_7457);
or U7778 (N_7778,N_7427,N_7558);
and U7779 (N_7779,N_7549,N_7446);
nand U7780 (N_7780,N_7482,N_7448);
or U7781 (N_7781,N_7572,N_7597);
xnor U7782 (N_7782,N_7447,N_7532);
and U7783 (N_7783,N_7428,N_7495);
nor U7784 (N_7784,N_7586,N_7436);
or U7785 (N_7785,N_7429,N_7541);
nor U7786 (N_7786,N_7557,N_7561);
or U7787 (N_7787,N_7441,N_7481);
nor U7788 (N_7788,N_7461,N_7517);
nand U7789 (N_7789,N_7593,N_7599);
or U7790 (N_7790,N_7481,N_7468);
or U7791 (N_7791,N_7517,N_7437);
nand U7792 (N_7792,N_7484,N_7420);
and U7793 (N_7793,N_7463,N_7520);
and U7794 (N_7794,N_7448,N_7461);
xor U7795 (N_7795,N_7507,N_7432);
nor U7796 (N_7796,N_7560,N_7488);
nand U7797 (N_7797,N_7504,N_7536);
xnor U7798 (N_7798,N_7421,N_7448);
xnor U7799 (N_7799,N_7512,N_7572);
nor U7800 (N_7800,N_7719,N_7751);
or U7801 (N_7801,N_7798,N_7718);
or U7802 (N_7802,N_7628,N_7654);
or U7803 (N_7803,N_7796,N_7780);
nand U7804 (N_7804,N_7636,N_7629);
nand U7805 (N_7805,N_7608,N_7799);
xnor U7806 (N_7806,N_7783,N_7788);
nand U7807 (N_7807,N_7601,N_7659);
nor U7808 (N_7808,N_7741,N_7637);
or U7809 (N_7809,N_7745,N_7769);
nor U7810 (N_7810,N_7770,N_7795);
nor U7811 (N_7811,N_7771,N_7641);
or U7812 (N_7812,N_7716,N_7744);
nor U7813 (N_7813,N_7701,N_7649);
or U7814 (N_7814,N_7762,N_7790);
nor U7815 (N_7815,N_7765,N_7656);
nand U7816 (N_7816,N_7616,N_7617);
nor U7817 (N_7817,N_7682,N_7779);
nand U7818 (N_7818,N_7760,N_7670);
nand U7819 (N_7819,N_7664,N_7742);
or U7820 (N_7820,N_7605,N_7688);
nand U7821 (N_7821,N_7619,N_7679);
or U7822 (N_7822,N_7603,N_7729);
nand U7823 (N_7823,N_7724,N_7615);
or U7824 (N_7824,N_7695,N_7730);
nand U7825 (N_7825,N_7657,N_7661);
or U7826 (N_7826,N_7648,N_7667);
nor U7827 (N_7827,N_7686,N_7712);
or U7828 (N_7828,N_7600,N_7792);
xnor U7829 (N_7829,N_7631,N_7728);
nor U7830 (N_7830,N_7627,N_7772);
or U7831 (N_7831,N_7713,N_7732);
or U7832 (N_7832,N_7673,N_7633);
and U7833 (N_7833,N_7700,N_7638);
or U7834 (N_7834,N_7754,N_7613);
nor U7835 (N_7835,N_7684,N_7658);
nand U7836 (N_7836,N_7773,N_7775);
nand U7837 (N_7837,N_7714,N_7642);
and U7838 (N_7838,N_7768,N_7643);
xnor U7839 (N_7839,N_7675,N_7749);
nand U7840 (N_7840,N_7696,N_7650);
nor U7841 (N_7841,N_7708,N_7694);
nor U7842 (N_7842,N_7647,N_7727);
and U7843 (N_7843,N_7738,N_7787);
nand U7844 (N_7844,N_7639,N_7709);
and U7845 (N_7845,N_7683,N_7612);
and U7846 (N_7846,N_7747,N_7609);
nand U7847 (N_7847,N_7763,N_7652);
nor U7848 (N_7848,N_7755,N_7625);
nand U7849 (N_7849,N_7689,N_7662);
or U7850 (N_7850,N_7618,N_7753);
xor U7851 (N_7851,N_7630,N_7752);
nor U7852 (N_7852,N_7774,N_7668);
nor U7853 (N_7853,N_7722,N_7703);
nor U7854 (N_7854,N_7644,N_7663);
nand U7855 (N_7855,N_7674,N_7778);
nand U7856 (N_7856,N_7785,N_7733);
nand U7857 (N_7857,N_7702,N_7794);
xnor U7858 (N_7858,N_7735,N_7746);
nand U7859 (N_7859,N_7781,N_7678);
or U7860 (N_7860,N_7666,N_7715);
nor U7861 (N_7861,N_7669,N_7604);
and U7862 (N_7862,N_7705,N_7725);
and U7863 (N_7863,N_7743,N_7672);
and U7864 (N_7864,N_7767,N_7711);
or U7865 (N_7865,N_7606,N_7634);
nor U7866 (N_7866,N_7632,N_7635);
and U7867 (N_7867,N_7782,N_7610);
xnor U7868 (N_7868,N_7739,N_7624);
nand U7869 (N_7869,N_7761,N_7766);
nor U7870 (N_7870,N_7621,N_7640);
nand U7871 (N_7871,N_7726,N_7607);
nand U7872 (N_7872,N_7687,N_7660);
nand U7873 (N_7873,N_7707,N_7758);
or U7874 (N_7874,N_7655,N_7748);
and U7875 (N_7875,N_7731,N_7697);
nor U7876 (N_7876,N_7685,N_7690);
and U7877 (N_7877,N_7721,N_7723);
nand U7878 (N_7878,N_7693,N_7665);
nor U7879 (N_7879,N_7645,N_7626);
or U7880 (N_7880,N_7691,N_7797);
and U7881 (N_7881,N_7653,N_7757);
nor U7882 (N_7882,N_7740,N_7789);
xor U7883 (N_7883,N_7681,N_7676);
nand U7884 (N_7884,N_7671,N_7756);
xor U7885 (N_7885,N_7737,N_7710);
nor U7886 (N_7886,N_7776,N_7704);
nand U7887 (N_7887,N_7602,N_7777);
nor U7888 (N_7888,N_7699,N_7651);
nand U7889 (N_7889,N_7786,N_7784);
nand U7890 (N_7890,N_7698,N_7791);
and U7891 (N_7891,N_7736,N_7750);
xnor U7892 (N_7892,N_7734,N_7646);
nor U7893 (N_7893,N_7680,N_7706);
xor U7894 (N_7894,N_7793,N_7764);
and U7895 (N_7895,N_7623,N_7692);
xor U7896 (N_7896,N_7620,N_7622);
nor U7897 (N_7897,N_7614,N_7720);
nand U7898 (N_7898,N_7677,N_7717);
or U7899 (N_7899,N_7611,N_7759);
nor U7900 (N_7900,N_7789,N_7659);
and U7901 (N_7901,N_7778,N_7655);
xnor U7902 (N_7902,N_7640,N_7742);
nand U7903 (N_7903,N_7751,N_7780);
nor U7904 (N_7904,N_7794,N_7751);
and U7905 (N_7905,N_7642,N_7729);
nand U7906 (N_7906,N_7754,N_7637);
nor U7907 (N_7907,N_7709,N_7697);
nor U7908 (N_7908,N_7730,N_7651);
nor U7909 (N_7909,N_7785,N_7767);
nand U7910 (N_7910,N_7694,N_7619);
nor U7911 (N_7911,N_7682,N_7739);
nand U7912 (N_7912,N_7709,N_7771);
nor U7913 (N_7913,N_7680,N_7628);
or U7914 (N_7914,N_7762,N_7690);
nand U7915 (N_7915,N_7615,N_7713);
nand U7916 (N_7916,N_7722,N_7781);
and U7917 (N_7917,N_7620,N_7791);
xor U7918 (N_7918,N_7657,N_7622);
nand U7919 (N_7919,N_7777,N_7692);
nor U7920 (N_7920,N_7631,N_7710);
or U7921 (N_7921,N_7767,N_7784);
and U7922 (N_7922,N_7759,N_7742);
xor U7923 (N_7923,N_7771,N_7728);
and U7924 (N_7924,N_7789,N_7667);
nand U7925 (N_7925,N_7799,N_7739);
or U7926 (N_7926,N_7790,N_7631);
and U7927 (N_7927,N_7679,N_7723);
or U7928 (N_7928,N_7674,N_7616);
nand U7929 (N_7929,N_7787,N_7749);
and U7930 (N_7930,N_7613,N_7718);
or U7931 (N_7931,N_7700,N_7798);
nand U7932 (N_7932,N_7606,N_7734);
and U7933 (N_7933,N_7646,N_7750);
and U7934 (N_7934,N_7639,N_7794);
or U7935 (N_7935,N_7684,N_7607);
or U7936 (N_7936,N_7785,N_7657);
nand U7937 (N_7937,N_7667,N_7664);
nor U7938 (N_7938,N_7685,N_7736);
or U7939 (N_7939,N_7666,N_7701);
nand U7940 (N_7940,N_7786,N_7649);
and U7941 (N_7941,N_7668,N_7659);
nand U7942 (N_7942,N_7641,N_7731);
and U7943 (N_7943,N_7705,N_7637);
nand U7944 (N_7944,N_7710,N_7661);
and U7945 (N_7945,N_7798,N_7635);
nand U7946 (N_7946,N_7698,N_7793);
nand U7947 (N_7947,N_7666,N_7631);
and U7948 (N_7948,N_7683,N_7613);
or U7949 (N_7949,N_7668,N_7651);
or U7950 (N_7950,N_7661,N_7768);
and U7951 (N_7951,N_7765,N_7711);
or U7952 (N_7952,N_7769,N_7757);
or U7953 (N_7953,N_7700,N_7659);
or U7954 (N_7954,N_7617,N_7737);
and U7955 (N_7955,N_7733,N_7674);
or U7956 (N_7956,N_7779,N_7662);
nor U7957 (N_7957,N_7662,N_7693);
and U7958 (N_7958,N_7763,N_7783);
or U7959 (N_7959,N_7721,N_7627);
or U7960 (N_7960,N_7666,N_7662);
and U7961 (N_7961,N_7749,N_7735);
and U7962 (N_7962,N_7710,N_7649);
and U7963 (N_7963,N_7787,N_7636);
xnor U7964 (N_7964,N_7717,N_7747);
and U7965 (N_7965,N_7623,N_7652);
nor U7966 (N_7966,N_7619,N_7623);
nand U7967 (N_7967,N_7772,N_7667);
xor U7968 (N_7968,N_7701,N_7727);
nor U7969 (N_7969,N_7710,N_7616);
nor U7970 (N_7970,N_7762,N_7617);
nand U7971 (N_7971,N_7604,N_7719);
or U7972 (N_7972,N_7680,N_7652);
xor U7973 (N_7973,N_7798,N_7782);
and U7974 (N_7974,N_7606,N_7639);
or U7975 (N_7975,N_7675,N_7734);
xnor U7976 (N_7976,N_7617,N_7776);
and U7977 (N_7977,N_7680,N_7740);
or U7978 (N_7978,N_7715,N_7693);
or U7979 (N_7979,N_7642,N_7785);
nor U7980 (N_7980,N_7786,N_7709);
or U7981 (N_7981,N_7745,N_7753);
nand U7982 (N_7982,N_7702,N_7669);
xor U7983 (N_7983,N_7659,N_7690);
and U7984 (N_7984,N_7744,N_7798);
xor U7985 (N_7985,N_7665,N_7651);
nor U7986 (N_7986,N_7749,N_7782);
nor U7987 (N_7987,N_7638,N_7652);
nand U7988 (N_7988,N_7775,N_7727);
nand U7989 (N_7989,N_7789,N_7653);
nor U7990 (N_7990,N_7630,N_7794);
nor U7991 (N_7991,N_7738,N_7716);
or U7992 (N_7992,N_7657,N_7610);
nor U7993 (N_7993,N_7739,N_7695);
or U7994 (N_7994,N_7724,N_7754);
nand U7995 (N_7995,N_7726,N_7654);
and U7996 (N_7996,N_7657,N_7746);
nand U7997 (N_7997,N_7694,N_7699);
nand U7998 (N_7998,N_7701,N_7751);
nor U7999 (N_7999,N_7687,N_7611);
or U8000 (N_8000,N_7946,N_7817);
and U8001 (N_8001,N_7829,N_7872);
nor U8002 (N_8002,N_7951,N_7954);
and U8003 (N_8003,N_7880,N_7800);
nand U8004 (N_8004,N_7849,N_7828);
xor U8005 (N_8005,N_7808,N_7809);
nor U8006 (N_8006,N_7933,N_7998);
nor U8007 (N_8007,N_7976,N_7968);
or U8008 (N_8008,N_7997,N_7804);
nor U8009 (N_8009,N_7993,N_7914);
nor U8010 (N_8010,N_7996,N_7881);
nor U8011 (N_8011,N_7969,N_7824);
and U8012 (N_8012,N_7831,N_7965);
and U8013 (N_8013,N_7898,N_7926);
and U8014 (N_8014,N_7897,N_7910);
nand U8015 (N_8015,N_7905,N_7967);
or U8016 (N_8016,N_7855,N_7947);
or U8017 (N_8017,N_7874,N_7932);
or U8018 (N_8018,N_7918,N_7978);
and U8019 (N_8019,N_7846,N_7981);
or U8020 (N_8020,N_7919,N_7915);
nand U8021 (N_8021,N_7823,N_7985);
or U8022 (N_8022,N_7963,N_7982);
nor U8023 (N_8023,N_7929,N_7805);
nor U8024 (N_8024,N_7973,N_7876);
and U8025 (N_8025,N_7907,N_7886);
nor U8026 (N_8026,N_7979,N_7826);
nor U8027 (N_8027,N_7801,N_7840);
nand U8028 (N_8028,N_7934,N_7901);
nor U8029 (N_8029,N_7999,N_7895);
xnor U8030 (N_8030,N_7960,N_7856);
nand U8031 (N_8031,N_7821,N_7995);
or U8032 (N_8032,N_7935,N_7812);
and U8033 (N_8033,N_7957,N_7896);
nand U8034 (N_8034,N_7852,N_7952);
xor U8035 (N_8035,N_7889,N_7866);
nand U8036 (N_8036,N_7890,N_7879);
and U8037 (N_8037,N_7888,N_7945);
xnor U8038 (N_8038,N_7814,N_7989);
or U8039 (N_8039,N_7815,N_7902);
nor U8040 (N_8040,N_7883,N_7803);
and U8041 (N_8041,N_7862,N_7830);
or U8042 (N_8042,N_7868,N_7950);
xor U8043 (N_8043,N_7865,N_7949);
nor U8044 (N_8044,N_7845,N_7974);
or U8045 (N_8045,N_7847,N_7955);
or U8046 (N_8046,N_7983,N_7953);
or U8047 (N_8047,N_7875,N_7850);
or U8048 (N_8048,N_7958,N_7835);
and U8049 (N_8049,N_7966,N_7970);
and U8050 (N_8050,N_7924,N_7972);
or U8051 (N_8051,N_7820,N_7851);
and U8052 (N_8052,N_7892,N_7956);
and U8053 (N_8053,N_7819,N_7936);
nand U8054 (N_8054,N_7882,N_7848);
nand U8055 (N_8055,N_7911,N_7900);
xnor U8056 (N_8056,N_7977,N_7806);
or U8057 (N_8057,N_7885,N_7837);
nor U8058 (N_8058,N_7807,N_7822);
and U8059 (N_8059,N_7854,N_7833);
nor U8060 (N_8060,N_7992,N_7962);
and U8061 (N_8061,N_7904,N_7884);
or U8062 (N_8062,N_7913,N_7834);
and U8063 (N_8063,N_7988,N_7873);
and U8064 (N_8064,N_7909,N_7943);
and U8065 (N_8065,N_7857,N_7991);
or U8066 (N_8066,N_7859,N_7877);
nor U8067 (N_8067,N_7938,N_7964);
or U8068 (N_8068,N_7878,N_7825);
and U8069 (N_8069,N_7813,N_7811);
and U8070 (N_8070,N_7869,N_7858);
nor U8071 (N_8071,N_7975,N_7994);
nand U8072 (N_8072,N_7987,N_7930);
nand U8073 (N_8073,N_7818,N_7853);
nor U8074 (N_8074,N_7887,N_7871);
nor U8075 (N_8075,N_7860,N_7899);
nor U8076 (N_8076,N_7894,N_7870);
and U8077 (N_8077,N_7928,N_7841);
and U8078 (N_8078,N_7912,N_7944);
or U8079 (N_8079,N_7908,N_7980);
and U8080 (N_8080,N_7802,N_7971);
and U8081 (N_8081,N_7923,N_7927);
nor U8082 (N_8082,N_7961,N_7836);
nand U8083 (N_8083,N_7843,N_7984);
xor U8084 (N_8084,N_7903,N_7959);
nand U8085 (N_8085,N_7986,N_7864);
nand U8086 (N_8086,N_7939,N_7863);
xor U8087 (N_8087,N_7942,N_7940);
or U8088 (N_8088,N_7891,N_7931);
nor U8089 (N_8089,N_7937,N_7916);
or U8090 (N_8090,N_7920,N_7906);
and U8091 (N_8091,N_7844,N_7810);
nor U8092 (N_8092,N_7838,N_7861);
nor U8093 (N_8093,N_7925,N_7922);
xor U8094 (N_8094,N_7921,N_7917);
nand U8095 (N_8095,N_7941,N_7839);
or U8096 (N_8096,N_7827,N_7948);
nand U8097 (N_8097,N_7842,N_7816);
nand U8098 (N_8098,N_7832,N_7893);
or U8099 (N_8099,N_7990,N_7867);
or U8100 (N_8100,N_7870,N_7804);
or U8101 (N_8101,N_7846,N_7823);
nand U8102 (N_8102,N_7915,N_7987);
nand U8103 (N_8103,N_7892,N_7994);
or U8104 (N_8104,N_7995,N_7983);
nand U8105 (N_8105,N_7997,N_7871);
nand U8106 (N_8106,N_7971,N_7941);
nand U8107 (N_8107,N_7935,N_7844);
nor U8108 (N_8108,N_7826,N_7823);
and U8109 (N_8109,N_7839,N_7814);
and U8110 (N_8110,N_7897,N_7860);
or U8111 (N_8111,N_7963,N_7902);
nand U8112 (N_8112,N_7906,N_7927);
nor U8113 (N_8113,N_7921,N_7880);
and U8114 (N_8114,N_7923,N_7815);
and U8115 (N_8115,N_7904,N_7920);
or U8116 (N_8116,N_7836,N_7896);
nand U8117 (N_8117,N_7870,N_7857);
or U8118 (N_8118,N_7810,N_7910);
nand U8119 (N_8119,N_7844,N_7934);
xor U8120 (N_8120,N_7800,N_7989);
xor U8121 (N_8121,N_7848,N_7966);
nand U8122 (N_8122,N_7897,N_7872);
or U8123 (N_8123,N_7957,N_7872);
nor U8124 (N_8124,N_7998,N_7976);
nor U8125 (N_8125,N_7828,N_7896);
or U8126 (N_8126,N_7997,N_7807);
and U8127 (N_8127,N_7999,N_7993);
and U8128 (N_8128,N_7932,N_7853);
and U8129 (N_8129,N_7934,N_7963);
and U8130 (N_8130,N_7957,N_7980);
nand U8131 (N_8131,N_7960,N_7902);
and U8132 (N_8132,N_7908,N_7912);
nor U8133 (N_8133,N_7900,N_7859);
and U8134 (N_8134,N_7980,N_7803);
and U8135 (N_8135,N_7805,N_7952);
nand U8136 (N_8136,N_7941,N_7876);
or U8137 (N_8137,N_7992,N_7995);
nor U8138 (N_8138,N_7845,N_7946);
nand U8139 (N_8139,N_7834,N_7823);
nor U8140 (N_8140,N_7930,N_7848);
nor U8141 (N_8141,N_7991,N_7844);
or U8142 (N_8142,N_7801,N_7874);
nor U8143 (N_8143,N_7995,N_7812);
or U8144 (N_8144,N_7938,N_7948);
or U8145 (N_8145,N_7853,N_7813);
nand U8146 (N_8146,N_7985,N_7855);
or U8147 (N_8147,N_7845,N_7932);
nor U8148 (N_8148,N_7903,N_7816);
or U8149 (N_8149,N_7898,N_7849);
xor U8150 (N_8150,N_7994,N_7999);
or U8151 (N_8151,N_7926,N_7915);
or U8152 (N_8152,N_7883,N_7811);
nor U8153 (N_8153,N_7915,N_7859);
nand U8154 (N_8154,N_7927,N_7879);
nand U8155 (N_8155,N_7846,N_7859);
nand U8156 (N_8156,N_7901,N_7886);
or U8157 (N_8157,N_7976,N_7888);
nor U8158 (N_8158,N_7894,N_7993);
or U8159 (N_8159,N_7855,N_7973);
and U8160 (N_8160,N_7990,N_7999);
or U8161 (N_8161,N_7810,N_7863);
xnor U8162 (N_8162,N_7906,N_7890);
or U8163 (N_8163,N_7969,N_7870);
xnor U8164 (N_8164,N_7957,N_7821);
or U8165 (N_8165,N_7958,N_7814);
nor U8166 (N_8166,N_7852,N_7922);
nor U8167 (N_8167,N_7808,N_7919);
and U8168 (N_8168,N_7946,N_7918);
nor U8169 (N_8169,N_7941,N_7987);
nor U8170 (N_8170,N_7905,N_7931);
nand U8171 (N_8171,N_7844,N_7820);
and U8172 (N_8172,N_7929,N_7923);
nand U8173 (N_8173,N_7968,N_7996);
or U8174 (N_8174,N_7801,N_7958);
nand U8175 (N_8175,N_7804,N_7821);
nand U8176 (N_8176,N_7965,N_7911);
xnor U8177 (N_8177,N_7909,N_7842);
xnor U8178 (N_8178,N_7879,N_7960);
nand U8179 (N_8179,N_7985,N_7839);
xnor U8180 (N_8180,N_7988,N_7911);
nor U8181 (N_8181,N_7823,N_7912);
or U8182 (N_8182,N_7999,N_7846);
and U8183 (N_8183,N_7946,N_7823);
or U8184 (N_8184,N_7975,N_7874);
nand U8185 (N_8185,N_7904,N_7963);
nor U8186 (N_8186,N_7968,N_7875);
or U8187 (N_8187,N_7889,N_7971);
nand U8188 (N_8188,N_7890,N_7824);
nand U8189 (N_8189,N_7982,N_7860);
nand U8190 (N_8190,N_7896,N_7985);
or U8191 (N_8191,N_7838,N_7878);
or U8192 (N_8192,N_7942,N_7973);
nor U8193 (N_8193,N_7978,N_7929);
and U8194 (N_8194,N_7937,N_7894);
and U8195 (N_8195,N_7979,N_7844);
or U8196 (N_8196,N_7991,N_7995);
xor U8197 (N_8197,N_7819,N_7844);
nand U8198 (N_8198,N_7942,N_7893);
or U8199 (N_8199,N_7979,N_7811);
nor U8200 (N_8200,N_8030,N_8049);
and U8201 (N_8201,N_8196,N_8040);
and U8202 (N_8202,N_8126,N_8106);
and U8203 (N_8203,N_8177,N_8138);
and U8204 (N_8204,N_8052,N_8179);
nor U8205 (N_8205,N_8152,N_8010);
and U8206 (N_8206,N_8080,N_8026);
and U8207 (N_8207,N_8147,N_8178);
nor U8208 (N_8208,N_8169,N_8087);
or U8209 (N_8209,N_8027,N_8033);
nand U8210 (N_8210,N_8176,N_8012);
xor U8211 (N_8211,N_8155,N_8174);
or U8212 (N_8212,N_8133,N_8021);
xor U8213 (N_8213,N_8113,N_8186);
nand U8214 (N_8214,N_8024,N_8017);
xnor U8215 (N_8215,N_8060,N_8139);
or U8216 (N_8216,N_8162,N_8098);
nor U8217 (N_8217,N_8154,N_8159);
xor U8218 (N_8218,N_8168,N_8130);
nor U8219 (N_8219,N_8117,N_8045);
and U8220 (N_8220,N_8032,N_8193);
and U8221 (N_8221,N_8101,N_8118);
nor U8222 (N_8222,N_8151,N_8120);
or U8223 (N_8223,N_8119,N_8056);
xor U8224 (N_8224,N_8009,N_8163);
nor U8225 (N_8225,N_8131,N_8081);
or U8226 (N_8226,N_8153,N_8016);
and U8227 (N_8227,N_8195,N_8064);
or U8228 (N_8228,N_8157,N_8020);
nor U8229 (N_8229,N_8048,N_8094);
or U8230 (N_8230,N_8028,N_8038);
nor U8231 (N_8231,N_8076,N_8002);
or U8232 (N_8232,N_8142,N_8043);
nand U8233 (N_8233,N_8011,N_8143);
and U8234 (N_8234,N_8041,N_8085);
nand U8235 (N_8235,N_8135,N_8122);
or U8236 (N_8236,N_8190,N_8145);
or U8237 (N_8237,N_8042,N_8039);
or U8238 (N_8238,N_8070,N_8127);
nand U8239 (N_8239,N_8007,N_8191);
nor U8240 (N_8240,N_8086,N_8047);
xor U8241 (N_8241,N_8099,N_8058);
and U8242 (N_8242,N_8013,N_8005);
nand U8243 (N_8243,N_8181,N_8165);
and U8244 (N_8244,N_8173,N_8171);
nor U8245 (N_8245,N_8158,N_8136);
nand U8246 (N_8246,N_8116,N_8077);
nor U8247 (N_8247,N_8180,N_8006);
nand U8248 (N_8248,N_8102,N_8062);
nand U8249 (N_8249,N_8072,N_8103);
or U8250 (N_8250,N_8059,N_8022);
or U8251 (N_8251,N_8096,N_8084);
nor U8252 (N_8252,N_8150,N_8144);
or U8253 (N_8253,N_8034,N_8053);
nor U8254 (N_8254,N_8140,N_8167);
nor U8255 (N_8255,N_8114,N_8074);
or U8256 (N_8256,N_8105,N_8075);
nor U8257 (N_8257,N_8014,N_8082);
nand U8258 (N_8258,N_8069,N_8044);
and U8259 (N_8259,N_8137,N_8199);
and U8260 (N_8260,N_8008,N_8000);
nand U8261 (N_8261,N_8115,N_8172);
or U8262 (N_8262,N_8184,N_8025);
and U8263 (N_8263,N_8164,N_8068);
nand U8264 (N_8264,N_8183,N_8067);
nor U8265 (N_8265,N_8170,N_8100);
xnor U8266 (N_8266,N_8104,N_8097);
xnor U8267 (N_8267,N_8055,N_8079);
or U8268 (N_8268,N_8166,N_8091);
nand U8269 (N_8269,N_8001,N_8054);
and U8270 (N_8270,N_8182,N_8037);
nand U8271 (N_8271,N_8095,N_8066);
or U8272 (N_8272,N_8031,N_8029);
xor U8273 (N_8273,N_8111,N_8092);
nor U8274 (N_8274,N_8057,N_8128);
nand U8275 (N_8275,N_8090,N_8071);
and U8276 (N_8276,N_8088,N_8146);
xor U8277 (N_8277,N_8073,N_8156);
and U8278 (N_8278,N_8089,N_8112);
xnor U8279 (N_8279,N_8198,N_8065);
xor U8280 (N_8280,N_8078,N_8129);
nand U8281 (N_8281,N_8093,N_8125);
or U8282 (N_8282,N_8187,N_8134);
xnor U8283 (N_8283,N_8107,N_8003);
nor U8284 (N_8284,N_8036,N_8141);
nor U8285 (N_8285,N_8015,N_8175);
nand U8286 (N_8286,N_8110,N_8197);
nor U8287 (N_8287,N_8050,N_8108);
nor U8288 (N_8288,N_8121,N_8123);
nor U8289 (N_8289,N_8148,N_8023);
or U8290 (N_8290,N_8160,N_8189);
nor U8291 (N_8291,N_8083,N_8124);
and U8292 (N_8292,N_8132,N_8046);
nor U8293 (N_8293,N_8185,N_8109);
nand U8294 (N_8294,N_8063,N_8061);
or U8295 (N_8295,N_8004,N_8019);
or U8296 (N_8296,N_8192,N_8194);
xnor U8297 (N_8297,N_8188,N_8051);
nand U8298 (N_8298,N_8035,N_8161);
xor U8299 (N_8299,N_8149,N_8018);
nor U8300 (N_8300,N_8102,N_8020);
nand U8301 (N_8301,N_8122,N_8150);
and U8302 (N_8302,N_8191,N_8199);
or U8303 (N_8303,N_8153,N_8098);
nand U8304 (N_8304,N_8090,N_8045);
nor U8305 (N_8305,N_8150,N_8125);
nor U8306 (N_8306,N_8056,N_8185);
or U8307 (N_8307,N_8015,N_8122);
xnor U8308 (N_8308,N_8011,N_8165);
xnor U8309 (N_8309,N_8109,N_8149);
xnor U8310 (N_8310,N_8149,N_8033);
nand U8311 (N_8311,N_8178,N_8018);
nor U8312 (N_8312,N_8049,N_8061);
xor U8313 (N_8313,N_8112,N_8037);
or U8314 (N_8314,N_8161,N_8129);
and U8315 (N_8315,N_8076,N_8034);
nand U8316 (N_8316,N_8075,N_8179);
and U8317 (N_8317,N_8130,N_8149);
and U8318 (N_8318,N_8034,N_8114);
or U8319 (N_8319,N_8097,N_8090);
nand U8320 (N_8320,N_8159,N_8100);
and U8321 (N_8321,N_8193,N_8062);
nand U8322 (N_8322,N_8136,N_8186);
or U8323 (N_8323,N_8045,N_8075);
nor U8324 (N_8324,N_8058,N_8005);
and U8325 (N_8325,N_8171,N_8109);
and U8326 (N_8326,N_8024,N_8023);
or U8327 (N_8327,N_8064,N_8165);
nand U8328 (N_8328,N_8049,N_8194);
nand U8329 (N_8329,N_8097,N_8186);
or U8330 (N_8330,N_8106,N_8030);
and U8331 (N_8331,N_8071,N_8066);
nand U8332 (N_8332,N_8186,N_8158);
and U8333 (N_8333,N_8109,N_8091);
or U8334 (N_8334,N_8187,N_8139);
nor U8335 (N_8335,N_8112,N_8156);
nor U8336 (N_8336,N_8185,N_8187);
or U8337 (N_8337,N_8043,N_8041);
and U8338 (N_8338,N_8030,N_8182);
xnor U8339 (N_8339,N_8003,N_8135);
and U8340 (N_8340,N_8117,N_8163);
or U8341 (N_8341,N_8114,N_8192);
and U8342 (N_8342,N_8138,N_8066);
nor U8343 (N_8343,N_8134,N_8119);
or U8344 (N_8344,N_8116,N_8069);
nor U8345 (N_8345,N_8086,N_8016);
and U8346 (N_8346,N_8015,N_8140);
nand U8347 (N_8347,N_8103,N_8009);
nand U8348 (N_8348,N_8013,N_8154);
or U8349 (N_8349,N_8128,N_8111);
nor U8350 (N_8350,N_8127,N_8146);
and U8351 (N_8351,N_8097,N_8066);
nand U8352 (N_8352,N_8056,N_8058);
or U8353 (N_8353,N_8189,N_8194);
and U8354 (N_8354,N_8080,N_8153);
or U8355 (N_8355,N_8164,N_8014);
nor U8356 (N_8356,N_8134,N_8156);
nor U8357 (N_8357,N_8005,N_8137);
and U8358 (N_8358,N_8141,N_8090);
and U8359 (N_8359,N_8151,N_8076);
xnor U8360 (N_8360,N_8040,N_8068);
or U8361 (N_8361,N_8173,N_8118);
or U8362 (N_8362,N_8164,N_8030);
nand U8363 (N_8363,N_8163,N_8005);
or U8364 (N_8364,N_8063,N_8033);
and U8365 (N_8365,N_8063,N_8182);
nor U8366 (N_8366,N_8163,N_8058);
nor U8367 (N_8367,N_8068,N_8023);
and U8368 (N_8368,N_8014,N_8116);
and U8369 (N_8369,N_8158,N_8110);
and U8370 (N_8370,N_8035,N_8137);
nor U8371 (N_8371,N_8180,N_8089);
nand U8372 (N_8372,N_8146,N_8163);
nor U8373 (N_8373,N_8159,N_8141);
or U8374 (N_8374,N_8145,N_8070);
xor U8375 (N_8375,N_8014,N_8196);
or U8376 (N_8376,N_8190,N_8159);
and U8377 (N_8377,N_8008,N_8108);
nor U8378 (N_8378,N_8001,N_8044);
nor U8379 (N_8379,N_8082,N_8035);
nor U8380 (N_8380,N_8163,N_8135);
xnor U8381 (N_8381,N_8164,N_8073);
xor U8382 (N_8382,N_8060,N_8189);
nor U8383 (N_8383,N_8012,N_8000);
nor U8384 (N_8384,N_8044,N_8119);
xor U8385 (N_8385,N_8147,N_8000);
nand U8386 (N_8386,N_8184,N_8068);
nor U8387 (N_8387,N_8110,N_8049);
nand U8388 (N_8388,N_8086,N_8124);
or U8389 (N_8389,N_8062,N_8100);
nor U8390 (N_8390,N_8163,N_8077);
nor U8391 (N_8391,N_8024,N_8057);
or U8392 (N_8392,N_8177,N_8064);
and U8393 (N_8393,N_8197,N_8036);
nand U8394 (N_8394,N_8155,N_8110);
or U8395 (N_8395,N_8124,N_8118);
or U8396 (N_8396,N_8148,N_8127);
nor U8397 (N_8397,N_8183,N_8015);
nor U8398 (N_8398,N_8000,N_8146);
nor U8399 (N_8399,N_8017,N_8049);
nor U8400 (N_8400,N_8342,N_8273);
nand U8401 (N_8401,N_8260,N_8332);
or U8402 (N_8402,N_8350,N_8339);
xor U8403 (N_8403,N_8305,N_8236);
or U8404 (N_8404,N_8203,N_8307);
nor U8405 (N_8405,N_8397,N_8221);
nand U8406 (N_8406,N_8388,N_8294);
nor U8407 (N_8407,N_8284,N_8218);
or U8408 (N_8408,N_8210,N_8275);
and U8409 (N_8409,N_8225,N_8286);
nand U8410 (N_8410,N_8291,N_8296);
or U8411 (N_8411,N_8276,N_8295);
xor U8412 (N_8412,N_8249,N_8336);
nand U8413 (N_8413,N_8292,N_8246);
and U8414 (N_8414,N_8240,N_8328);
xnor U8415 (N_8415,N_8369,N_8245);
nand U8416 (N_8416,N_8341,N_8237);
nor U8417 (N_8417,N_8337,N_8263);
or U8418 (N_8418,N_8392,N_8343);
or U8419 (N_8419,N_8206,N_8258);
or U8420 (N_8420,N_8277,N_8274);
nand U8421 (N_8421,N_8362,N_8358);
nand U8422 (N_8422,N_8361,N_8393);
nand U8423 (N_8423,N_8248,N_8242);
and U8424 (N_8424,N_8227,N_8223);
and U8425 (N_8425,N_8323,N_8304);
nand U8426 (N_8426,N_8313,N_8375);
and U8427 (N_8427,N_8387,N_8300);
or U8428 (N_8428,N_8378,N_8231);
and U8429 (N_8429,N_8257,N_8298);
or U8430 (N_8430,N_8253,N_8244);
or U8431 (N_8431,N_8303,N_8290);
and U8432 (N_8432,N_8317,N_8380);
nor U8433 (N_8433,N_8318,N_8334);
and U8434 (N_8434,N_8239,N_8368);
nand U8435 (N_8435,N_8363,N_8209);
nand U8436 (N_8436,N_8321,N_8398);
nor U8437 (N_8437,N_8391,N_8222);
nand U8438 (N_8438,N_8338,N_8234);
nor U8439 (N_8439,N_8311,N_8355);
nor U8440 (N_8440,N_8285,N_8254);
nor U8441 (N_8441,N_8312,N_8385);
nand U8442 (N_8442,N_8335,N_8308);
and U8443 (N_8443,N_8266,N_8215);
nand U8444 (N_8444,N_8394,N_8214);
and U8445 (N_8445,N_8267,N_8271);
nand U8446 (N_8446,N_8372,N_8224);
and U8447 (N_8447,N_8322,N_8264);
nor U8448 (N_8448,N_8309,N_8238);
nor U8449 (N_8449,N_8255,N_8259);
xor U8450 (N_8450,N_8326,N_8226);
and U8451 (N_8451,N_8319,N_8219);
nand U8452 (N_8452,N_8306,N_8252);
and U8453 (N_8453,N_8346,N_8359);
and U8454 (N_8454,N_8302,N_8371);
nand U8455 (N_8455,N_8384,N_8315);
and U8456 (N_8456,N_8211,N_8360);
and U8457 (N_8457,N_8233,N_8243);
nor U8458 (N_8458,N_8314,N_8316);
and U8459 (N_8459,N_8280,N_8383);
xor U8460 (N_8460,N_8289,N_8293);
xnor U8461 (N_8461,N_8217,N_8310);
nand U8462 (N_8462,N_8377,N_8349);
or U8463 (N_8463,N_8265,N_8235);
nor U8464 (N_8464,N_8212,N_8201);
nand U8465 (N_8465,N_8390,N_8353);
xnor U8466 (N_8466,N_8287,N_8325);
xor U8467 (N_8467,N_8320,N_8247);
or U8468 (N_8468,N_8354,N_8270);
nand U8469 (N_8469,N_8357,N_8268);
and U8470 (N_8470,N_8331,N_8347);
and U8471 (N_8471,N_8327,N_8205);
nand U8472 (N_8472,N_8232,N_8262);
nor U8473 (N_8473,N_8373,N_8213);
nand U8474 (N_8474,N_8324,N_8348);
nand U8475 (N_8475,N_8345,N_8365);
xor U8476 (N_8476,N_8256,N_8376);
nor U8477 (N_8477,N_8370,N_8207);
nor U8478 (N_8478,N_8208,N_8200);
xnor U8479 (N_8479,N_8356,N_8261);
nand U8480 (N_8480,N_8386,N_8204);
xor U8481 (N_8481,N_8216,N_8395);
nand U8482 (N_8482,N_8229,N_8283);
nor U8483 (N_8483,N_8381,N_8364);
or U8484 (N_8484,N_8399,N_8250);
and U8485 (N_8485,N_8367,N_8251);
and U8486 (N_8486,N_8389,N_8299);
xnor U8487 (N_8487,N_8281,N_8278);
nor U8488 (N_8488,N_8344,N_8230);
nand U8489 (N_8489,N_8301,N_8279);
or U8490 (N_8490,N_8374,N_8330);
or U8491 (N_8491,N_8351,N_8340);
and U8492 (N_8492,N_8329,N_8228);
nor U8493 (N_8493,N_8269,N_8272);
nand U8494 (N_8494,N_8282,N_8288);
and U8495 (N_8495,N_8366,N_8352);
and U8496 (N_8496,N_8220,N_8297);
and U8497 (N_8497,N_8379,N_8382);
and U8498 (N_8498,N_8333,N_8241);
nand U8499 (N_8499,N_8396,N_8202);
nand U8500 (N_8500,N_8232,N_8224);
and U8501 (N_8501,N_8252,N_8204);
nand U8502 (N_8502,N_8378,N_8201);
or U8503 (N_8503,N_8363,N_8347);
and U8504 (N_8504,N_8359,N_8276);
nand U8505 (N_8505,N_8352,N_8345);
or U8506 (N_8506,N_8295,N_8281);
xor U8507 (N_8507,N_8208,N_8202);
or U8508 (N_8508,N_8205,N_8212);
or U8509 (N_8509,N_8264,N_8380);
or U8510 (N_8510,N_8342,N_8392);
or U8511 (N_8511,N_8362,N_8396);
xor U8512 (N_8512,N_8322,N_8368);
nor U8513 (N_8513,N_8312,N_8319);
and U8514 (N_8514,N_8353,N_8372);
xnor U8515 (N_8515,N_8237,N_8365);
or U8516 (N_8516,N_8284,N_8298);
and U8517 (N_8517,N_8374,N_8264);
nor U8518 (N_8518,N_8349,N_8239);
or U8519 (N_8519,N_8230,N_8329);
nor U8520 (N_8520,N_8258,N_8307);
nor U8521 (N_8521,N_8287,N_8333);
nand U8522 (N_8522,N_8369,N_8276);
or U8523 (N_8523,N_8240,N_8351);
nor U8524 (N_8524,N_8259,N_8250);
nand U8525 (N_8525,N_8246,N_8358);
or U8526 (N_8526,N_8258,N_8239);
and U8527 (N_8527,N_8290,N_8346);
or U8528 (N_8528,N_8356,N_8333);
nor U8529 (N_8529,N_8388,N_8377);
and U8530 (N_8530,N_8257,N_8205);
and U8531 (N_8531,N_8388,N_8332);
or U8532 (N_8532,N_8299,N_8317);
and U8533 (N_8533,N_8355,N_8322);
nand U8534 (N_8534,N_8247,N_8319);
xnor U8535 (N_8535,N_8285,N_8330);
or U8536 (N_8536,N_8232,N_8382);
nor U8537 (N_8537,N_8233,N_8295);
nor U8538 (N_8538,N_8296,N_8200);
nand U8539 (N_8539,N_8341,N_8300);
or U8540 (N_8540,N_8353,N_8304);
nor U8541 (N_8541,N_8377,N_8236);
xnor U8542 (N_8542,N_8216,N_8205);
xnor U8543 (N_8543,N_8280,N_8278);
or U8544 (N_8544,N_8288,N_8269);
or U8545 (N_8545,N_8309,N_8339);
nand U8546 (N_8546,N_8321,N_8304);
nor U8547 (N_8547,N_8368,N_8236);
xnor U8548 (N_8548,N_8341,N_8388);
and U8549 (N_8549,N_8228,N_8285);
or U8550 (N_8550,N_8392,N_8242);
nand U8551 (N_8551,N_8300,N_8247);
nor U8552 (N_8552,N_8306,N_8368);
or U8553 (N_8553,N_8267,N_8278);
or U8554 (N_8554,N_8333,N_8219);
xnor U8555 (N_8555,N_8269,N_8260);
nor U8556 (N_8556,N_8339,N_8252);
or U8557 (N_8557,N_8265,N_8242);
or U8558 (N_8558,N_8278,N_8201);
or U8559 (N_8559,N_8277,N_8314);
nor U8560 (N_8560,N_8351,N_8205);
or U8561 (N_8561,N_8235,N_8216);
xnor U8562 (N_8562,N_8397,N_8288);
or U8563 (N_8563,N_8393,N_8327);
nand U8564 (N_8564,N_8244,N_8303);
nor U8565 (N_8565,N_8324,N_8279);
nand U8566 (N_8566,N_8341,N_8369);
and U8567 (N_8567,N_8355,N_8327);
nor U8568 (N_8568,N_8347,N_8359);
and U8569 (N_8569,N_8390,N_8279);
or U8570 (N_8570,N_8333,N_8229);
nand U8571 (N_8571,N_8267,N_8398);
nand U8572 (N_8572,N_8226,N_8355);
nand U8573 (N_8573,N_8329,N_8212);
and U8574 (N_8574,N_8349,N_8291);
xor U8575 (N_8575,N_8351,N_8271);
nand U8576 (N_8576,N_8297,N_8386);
nor U8577 (N_8577,N_8398,N_8290);
nor U8578 (N_8578,N_8362,N_8211);
xnor U8579 (N_8579,N_8260,N_8270);
nor U8580 (N_8580,N_8230,N_8273);
xnor U8581 (N_8581,N_8282,N_8308);
nor U8582 (N_8582,N_8394,N_8304);
and U8583 (N_8583,N_8233,N_8319);
xor U8584 (N_8584,N_8227,N_8376);
nand U8585 (N_8585,N_8316,N_8238);
or U8586 (N_8586,N_8395,N_8217);
nor U8587 (N_8587,N_8251,N_8250);
and U8588 (N_8588,N_8363,N_8361);
and U8589 (N_8589,N_8335,N_8270);
and U8590 (N_8590,N_8332,N_8365);
xor U8591 (N_8591,N_8354,N_8342);
nor U8592 (N_8592,N_8296,N_8325);
and U8593 (N_8593,N_8281,N_8340);
or U8594 (N_8594,N_8364,N_8329);
nor U8595 (N_8595,N_8202,N_8206);
or U8596 (N_8596,N_8246,N_8360);
and U8597 (N_8597,N_8240,N_8219);
and U8598 (N_8598,N_8270,N_8359);
nor U8599 (N_8599,N_8246,N_8376);
or U8600 (N_8600,N_8561,N_8416);
and U8601 (N_8601,N_8408,N_8589);
nand U8602 (N_8602,N_8420,N_8462);
nand U8603 (N_8603,N_8442,N_8432);
nand U8604 (N_8604,N_8469,N_8493);
and U8605 (N_8605,N_8487,N_8405);
or U8606 (N_8606,N_8490,N_8551);
nor U8607 (N_8607,N_8519,N_8497);
or U8608 (N_8608,N_8550,N_8477);
or U8609 (N_8609,N_8573,N_8574);
or U8610 (N_8610,N_8449,N_8591);
or U8611 (N_8611,N_8584,N_8562);
and U8612 (N_8612,N_8455,N_8407);
and U8613 (N_8613,N_8549,N_8505);
and U8614 (N_8614,N_8596,N_8412);
and U8615 (N_8615,N_8483,N_8476);
nor U8616 (N_8616,N_8475,N_8566);
and U8617 (N_8617,N_8448,N_8555);
and U8618 (N_8618,N_8576,N_8451);
and U8619 (N_8619,N_8543,N_8533);
or U8620 (N_8620,N_8521,N_8517);
nand U8621 (N_8621,N_8516,N_8542);
or U8622 (N_8622,N_8458,N_8577);
or U8623 (N_8623,N_8563,N_8464);
and U8624 (N_8624,N_8414,N_8472);
and U8625 (N_8625,N_8529,N_8447);
nor U8626 (N_8626,N_8436,N_8431);
or U8627 (N_8627,N_8488,N_8541);
and U8628 (N_8628,N_8583,N_8480);
xnor U8629 (N_8629,N_8413,N_8481);
and U8630 (N_8630,N_8444,N_8568);
and U8631 (N_8631,N_8524,N_8553);
nand U8632 (N_8632,N_8507,N_8498);
nand U8633 (N_8633,N_8482,N_8466);
xor U8634 (N_8634,N_8470,N_8578);
or U8635 (N_8635,N_8567,N_8552);
or U8636 (N_8636,N_8599,N_8425);
nor U8637 (N_8637,N_8544,N_8513);
xor U8638 (N_8638,N_8424,N_8418);
and U8639 (N_8639,N_8520,N_8426);
or U8640 (N_8640,N_8421,N_8415);
nor U8641 (N_8641,N_8588,N_8427);
nand U8642 (N_8642,N_8502,N_8459);
nor U8643 (N_8643,N_8545,N_8400);
nor U8644 (N_8644,N_8503,N_8471);
or U8645 (N_8645,N_8499,N_8523);
or U8646 (N_8646,N_8509,N_8560);
nor U8647 (N_8647,N_8546,N_8479);
xor U8648 (N_8648,N_8575,N_8539);
and U8649 (N_8649,N_8548,N_8515);
or U8650 (N_8650,N_8428,N_8440);
or U8651 (N_8651,N_8496,N_8494);
or U8652 (N_8652,N_8558,N_8463);
or U8653 (N_8653,N_8450,N_8592);
nand U8654 (N_8654,N_8441,N_8525);
nor U8655 (N_8655,N_8510,N_8406);
and U8656 (N_8656,N_8527,N_8410);
nand U8657 (N_8657,N_8586,N_8437);
xor U8658 (N_8658,N_8417,N_8535);
xor U8659 (N_8659,N_8536,N_8478);
nand U8660 (N_8660,N_8489,N_8402);
nand U8661 (N_8661,N_8508,N_8500);
nand U8662 (N_8662,N_8495,N_8429);
and U8663 (N_8663,N_8411,N_8443);
and U8664 (N_8664,N_8491,N_8595);
and U8665 (N_8665,N_8559,N_8474);
nand U8666 (N_8666,N_8556,N_8452);
and U8667 (N_8667,N_8457,N_8492);
nor U8668 (N_8668,N_8485,N_8581);
nand U8669 (N_8669,N_8531,N_8572);
and U8670 (N_8670,N_8501,N_8590);
nor U8671 (N_8671,N_8511,N_8461);
nor U8672 (N_8672,N_8473,N_8403);
nor U8673 (N_8673,N_8434,N_8404);
nand U8674 (N_8674,N_8422,N_8518);
nand U8675 (N_8675,N_8597,N_8565);
or U8676 (N_8676,N_8569,N_8438);
or U8677 (N_8677,N_8460,N_8439);
nor U8678 (N_8678,N_8594,N_8409);
and U8679 (N_8679,N_8532,N_8571);
and U8680 (N_8680,N_8504,N_8582);
nor U8681 (N_8681,N_8593,N_8423);
nor U8682 (N_8682,N_8570,N_8401);
nor U8683 (N_8683,N_8512,N_8547);
nand U8684 (N_8684,N_8468,N_8579);
nor U8685 (N_8685,N_8435,N_8419);
and U8686 (N_8686,N_8433,N_8538);
and U8687 (N_8687,N_8534,N_8554);
nand U8688 (N_8688,N_8564,N_8528);
xor U8689 (N_8689,N_8587,N_8456);
nand U8690 (N_8690,N_8506,N_8484);
nor U8691 (N_8691,N_8522,N_8530);
nand U8692 (N_8692,N_8537,N_8453);
nand U8693 (N_8693,N_8557,N_8585);
nor U8694 (N_8694,N_8467,N_8486);
nand U8695 (N_8695,N_8465,N_8514);
xor U8696 (N_8696,N_8540,N_8598);
xor U8697 (N_8697,N_8526,N_8454);
or U8698 (N_8698,N_8580,N_8446);
or U8699 (N_8699,N_8430,N_8445);
nor U8700 (N_8700,N_8464,N_8582);
or U8701 (N_8701,N_8530,N_8430);
and U8702 (N_8702,N_8492,N_8529);
nor U8703 (N_8703,N_8544,N_8468);
nor U8704 (N_8704,N_8423,N_8533);
nor U8705 (N_8705,N_8458,N_8460);
nand U8706 (N_8706,N_8509,N_8471);
or U8707 (N_8707,N_8530,N_8487);
and U8708 (N_8708,N_8560,N_8575);
nor U8709 (N_8709,N_8422,N_8588);
and U8710 (N_8710,N_8444,N_8592);
nor U8711 (N_8711,N_8486,N_8483);
or U8712 (N_8712,N_8533,N_8414);
nor U8713 (N_8713,N_8401,N_8470);
or U8714 (N_8714,N_8586,N_8599);
nand U8715 (N_8715,N_8596,N_8415);
nor U8716 (N_8716,N_8423,N_8438);
xnor U8717 (N_8717,N_8513,N_8559);
or U8718 (N_8718,N_8570,N_8592);
nor U8719 (N_8719,N_8551,N_8521);
nand U8720 (N_8720,N_8449,N_8595);
nor U8721 (N_8721,N_8466,N_8484);
or U8722 (N_8722,N_8502,N_8559);
xor U8723 (N_8723,N_8432,N_8424);
or U8724 (N_8724,N_8481,N_8599);
and U8725 (N_8725,N_8409,N_8538);
xor U8726 (N_8726,N_8507,N_8495);
or U8727 (N_8727,N_8597,N_8478);
or U8728 (N_8728,N_8430,N_8523);
and U8729 (N_8729,N_8441,N_8476);
or U8730 (N_8730,N_8545,N_8473);
nor U8731 (N_8731,N_8540,N_8510);
nor U8732 (N_8732,N_8507,N_8422);
or U8733 (N_8733,N_8454,N_8461);
nand U8734 (N_8734,N_8502,N_8519);
and U8735 (N_8735,N_8560,N_8414);
nand U8736 (N_8736,N_8409,N_8563);
nand U8737 (N_8737,N_8458,N_8555);
nand U8738 (N_8738,N_8549,N_8557);
and U8739 (N_8739,N_8428,N_8589);
and U8740 (N_8740,N_8468,N_8516);
and U8741 (N_8741,N_8482,N_8400);
nand U8742 (N_8742,N_8564,N_8591);
nand U8743 (N_8743,N_8499,N_8518);
and U8744 (N_8744,N_8443,N_8500);
and U8745 (N_8745,N_8581,N_8432);
nor U8746 (N_8746,N_8554,N_8564);
nand U8747 (N_8747,N_8408,N_8431);
nor U8748 (N_8748,N_8475,N_8543);
nand U8749 (N_8749,N_8433,N_8539);
or U8750 (N_8750,N_8567,N_8477);
or U8751 (N_8751,N_8576,N_8407);
and U8752 (N_8752,N_8433,N_8467);
or U8753 (N_8753,N_8593,N_8474);
nand U8754 (N_8754,N_8583,N_8427);
xor U8755 (N_8755,N_8534,N_8533);
or U8756 (N_8756,N_8415,N_8405);
nor U8757 (N_8757,N_8437,N_8459);
nand U8758 (N_8758,N_8405,N_8556);
xnor U8759 (N_8759,N_8534,N_8575);
or U8760 (N_8760,N_8581,N_8470);
nor U8761 (N_8761,N_8568,N_8425);
xnor U8762 (N_8762,N_8517,N_8487);
nor U8763 (N_8763,N_8417,N_8435);
nor U8764 (N_8764,N_8581,N_8563);
nand U8765 (N_8765,N_8555,N_8478);
and U8766 (N_8766,N_8465,N_8565);
nor U8767 (N_8767,N_8542,N_8410);
nor U8768 (N_8768,N_8496,N_8445);
nor U8769 (N_8769,N_8495,N_8531);
nor U8770 (N_8770,N_8576,N_8507);
or U8771 (N_8771,N_8580,N_8404);
nor U8772 (N_8772,N_8441,N_8518);
nor U8773 (N_8773,N_8593,N_8419);
and U8774 (N_8774,N_8583,N_8587);
nand U8775 (N_8775,N_8553,N_8477);
and U8776 (N_8776,N_8410,N_8487);
nor U8777 (N_8777,N_8554,N_8491);
xnor U8778 (N_8778,N_8520,N_8454);
nor U8779 (N_8779,N_8569,N_8599);
nand U8780 (N_8780,N_8514,N_8595);
xnor U8781 (N_8781,N_8411,N_8458);
nor U8782 (N_8782,N_8480,N_8424);
nand U8783 (N_8783,N_8451,N_8554);
and U8784 (N_8784,N_8523,N_8459);
nand U8785 (N_8785,N_8529,N_8473);
and U8786 (N_8786,N_8560,N_8573);
or U8787 (N_8787,N_8582,N_8491);
and U8788 (N_8788,N_8596,N_8530);
and U8789 (N_8789,N_8541,N_8528);
and U8790 (N_8790,N_8576,N_8469);
nor U8791 (N_8791,N_8540,N_8473);
nand U8792 (N_8792,N_8433,N_8552);
nand U8793 (N_8793,N_8558,N_8522);
or U8794 (N_8794,N_8498,N_8495);
nand U8795 (N_8795,N_8544,N_8588);
nand U8796 (N_8796,N_8460,N_8483);
nor U8797 (N_8797,N_8582,N_8572);
nand U8798 (N_8798,N_8403,N_8581);
nand U8799 (N_8799,N_8415,N_8449);
nor U8800 (N_8800,N_8647,N_8714);
nor U8801 (N_8801,N_8600,N_8658);
and U8802 (N_8802,N_8746,N_8664);
xor U8803 (N_8803,N_8741,N_8743);
nor U8804 (N_8804,N_8675,N_8782);
xor U8805 (N_8805,N_8739,N_8663);
nand U8806 (N_8806,N_8601,N_8642);
xor U8807 (N_8807,N_8603,N_8748);
or U8808 (N_8808,N_8711,N_8635);
and U8809 (N_8809,N_8680,N_8684);
or U8810 (N_8810,N_8662,N_8760);
and U8811 (N_8811,N_8715,N_8671);
nor U8812 (N_8812,N_8790,N_8700);
or U8813 (N_8813,N_8673,N_8606);
or U8814 (N_8814,N_8660,N_8654);
nor U8815 (N_8815,N_8645,N_8631);
or U8816 (N_8816,N_8681,N_8736);
or U8817 (N_8817,N_8689,N_8686);
nor U8818 (N_8818,N_8756,N_8722);
nor U8819 (N_8819,N_8698,N_8665);
and U8820 (N_8820,N_8707,N_8632);
and U8821 (N_8821,N_8624,N_8695);
xnor U8822 (N_8822,N_8728,N_8626);
and U8823 (N_8823,N_8786,N_8691);
nor U8824 (N_8824,N_8639,N_8781);
or U8825 (N_8825,N_8704,N_8648);
or U8826 (N_8826,N_8777,N_8633);
and U8827 (N_8827,N_8737,N_8692);
or U8828 (N_8828,N_8629,N_8751);
or U8829 (N_8829,N_8795,N_8763);
xor U8830 (N_8830,N_8716,N_8734);
nor U8831 (N_8831,N_8667,N_8609);
or U8832 (N_8832,N_8674,N_8764);
nand U8833 (N_8833,N_8646,N_8617);
xor U8834 (N_8834,N_8750,N_8668);
nand U8835 (N_8835,N_8643,N_8683);
and U8836 (N_8836,N_8669,N_8602);
and U8837 (N_8837,N_8717,N_8688);
nor U8838 (N_8838,N_8738,N_8780);
nand U8839 (N_8839,N_8725,N_8718);
xor U8840 (N_8840,N_8731,N_8727);
or U8841 (N_8841,N_8723,N_8752);
xor U8842 (N_8842,N_8693,N_8625);
nor U8843 (N_8843,N_8623,N_8670);
or U8844 (N_8844,N_8791,N_8677);
xor U8845 (N_8845,N_8701,N_8690);
or U8846 (N_8846,N_8789,N_8672);
nand U8847 (N_8847,N_8783,N_8744);
xnor U8848 (N_8848,N_8710,N_8641);
or U8849 (N_8849,N_8788,N_8769);
nor U8850 (N_8850,N_8613,N_8726);
nand U8851 (N_8851,N_8767,N_8705);
xnor U8852 (N_8852,N_8721,N_8618);
nor U8853 (N_8853,N_8720,N_8614);
or U8854 (N_8854,N_8605,N_8649);
nor U8855 (N_8855,N_8699,N_8753);
and U8856 (N_8856,N_8712,N_8657);
nand U8857 (N_8857,N_8615,N_8730);
and U8858 (N_8858,N_8676,N_8765);
nand U8859 (N_8859,N_8799,N_8794);
nand U8860 (N_8860,N_8640,N_8735);
nor U8861 (N_8861,N_8778,N_8796);
nor U8862 (N_8862,N_8733,N_8685);
and U8863 (N_8863,N_8636,N_8637);
or U8864 (N_8864,N_8679,N_8610);
and U8865 (N_8865,N_8644,N_8620);
nand U8866 (N_8866,N_8628,N_8772);
nor U8867 (N_8867,N_8619,N_8708);
nand U8868 (N_8868,N_8770,N_8621);
and U8869 (N_8869,N_8792,N_8697);
nor U8870 (N_8870,N_8754,N_8762);
nand U8871 (N_8871,N_8757,N_8634);
or U8872 (N_8872,N_8729,N_8758);
and U8873 (N_8873,N_8755,N_8775);
nand U8874 (N_8874,N_8732,N_8687);
nand U8875 (N_8875,N_8666,N_8768);
nand U8876 (N_8876,N_8793,N_8709);
or U8877 (N_8877,N_8622,N_8611);
nor U8878 (N_8878,N_8749,N_8759);
and U8879 (N_8879,N_8784,N_8798);
or U8880 (N_8880,N_8785,N_8696);
xor U8881 (N_8881,N_8612,N_8766);
and U8882 (N_8882,N_8607,N_8774);
and U8883 (N_8883,N_8682,N_8604);
nor U8884 (N_8884,N_8652,N_8747);
nand U8885 (N_8885,N_8656,N_8702);
and U8886 (N_8886,N_8661,N_8713);
and U8887 (N_8887,N_8787,N_8653);
or U8888 (N_8888,N_8742,N_8627);
nor U8889 (N_8889,N_8771,N_8630);
nand U8890 (N_8890,N_8761,N_8724);
xnor U8891 (N_8891,N_8608,N_8719);
or U8892 (N_8892,N_8779,N_8638);
nor U8893 (N_8893,N_8703,N_8776);
and U8894 (N_8894,N_8745,N_8659);
nor U8895 (N_8895,N_8773,N_8706);
nand U8896 (N_8896,N_8655,N_8797);
xor U8897 (N_8897,N_8678,N_8694);
nor U8898 (N_8898,N_8650,N_8740);
xor U8899 (N_8899,N_8616,N_8651);
or U8900 (N_8900,N_8673,N_8701);
or U8901 (N_8901,N_8709,N_8750);
and U8902 (N_8902,N_8613,N_8675);
and U8903 (N_8903,N_8671,N_8707);
nor U8904 (N_8904,N_8699,N_8745);
or U8905 (N_8905,N_8639,N_8664);
nand U8906 (N_8906,N_8757,N_8742);
and U8907 (N_8907,N_8799,N_8758);
xor U8908 (N_8908,N_8679,N_8658);
and U8909 (N_8909,N_8677,N_8657);
and U8910 (N_8910,N_8794,N_8689);
and U8911 (N_8911,N_8715,N_8777);
and U8912 (N_8912,N_8786,N_8735);
xnor U8913 (N_8913,N_8765,N_8760);
and U8914 (N_8914,N_8742,N_8792);
and U8915 (N_8915,N_8773,N_8720);
xor U8916 (N_8916,N_8670,N_8618);
or U8917 (N_8917,N_8628,N_8601);
nor U8918 (N_8918,N_8755,N_8644);
xnor U8919 (N_8919,N_8690,N_8660);
nand U8920 (N_8920,N_8688,N_8776);
xor U8921 (N_8921,N_8612,N_8722);
nand U8922 (N_8922,N_8698,N_8705);
nand U8923 (N_8923,N_8783,N_8630);
nor U8924 (N_8924,N_8726,N_8750);
xor U8925 (N_8925,N_8648,N_8778);
or U8926 (N_8926,N_8772,N_8716);
nand U8927 (N_8927,N_8655,N_8707);
xnor U8928 (N_8928,N_8719,N_8722);
nor U8929 (N_8929,N_8610,N_8774);
and U8930 (N_8930,N_8698,N_8680);
nor U8931 (N_8931,N_8772,N_8720);
nor U8932 (N_8932,N_8680,N_8601);
or U8933 (N_8933,N_8697,N_8643);
or U8934 (N_8934,N_8743,N_8721);
or U8935 (N_8935,N_8634,N_8613);
nand U8936 (N_8936,N_8762,N_8705);
xnor U8937 (N_8937,N_8753,N_8748);
xor U8938 (N_8938,N_8716,N_8731);
nand U8939 (N_8939,N_8719,N_8698);
nand U8940 (N_8940,N_8772,N_8733);
nand U8941 (N_8941,N_8645,N_8658);
or U8942 (N_8942,N_8784,N_8617);
nor U8943 (N_8943,N_8635,N_8765);
and U8944 (N_8944,N_8779,N_8672);
nor U8945 (N_8945,N_8602,N_8779);
nor U8946 (N_8946,N_8686,N_8757);
nand U8947 (N_8947,N_8621,N_8617);
nand U8948 (N_8948,N_8638,N_8798);
nand U8949 (N_8949,N_8700,N_8609);
or U8950 (N_8950,N_8737,N_8700);
nand U8951 (N_8951,N_8655,N_8648);
and U8952 (N_8952,N_8614,N_8634);
or U8953 (N_8953,N_8670,N_8774);
and U8954 (N_8954,N_8640,N_8760);
and U8955 (N_8955,N_8708,N_8677);
xor U8956 (N_8956,N_8630,N_8679);
and U8957 (N_8957,N_8745,N_8668);
or U8958 (N_8958,N_8720,N_8763);
and U8959 (N_8959,N_8685,N_8709);
nand U8960 (N_8960,N_8709,N_8707);
and U8961 (N_8961,N_8718,N_8731);
or U8962 (N_8962,N_8747,N_8798);
or U8963 (N_8963,N_8636,N_8775);
or U8964 (N_8964,N_8725,N_8759);
and U8965 (N_8965,N_8608,N_8660);
nor U8966 (N_8966,N_8644,N_8611);
and U8967 (N_8967,N_8777,N_8616);
or U8968 (N_8968,N_8741,N_8718);
xnor U8969 (N_8969,N_8623,N_8612);
or U8970 (N_8970,N_8750,N_8740);
and U8971 (N_8971,N_8647,N_8777);
or U8972 (N_8972,N_8672,N_8622);
nor U8973 (N_8973,N_8632,N_8646);
or U8974 (N_8974,N_8696,N_8711);
nor U8975 (N_8975,N_8724,N_8773);
nand U8976 (N_8976,N_8681,N_8601);
or U8977 (N_8977,N_8719,N_8792);
nor U8978 (N_8978,N_8696,N_8791);
and U8979 (N_8979,N_8784,N_8717);
or U8980 (N_8980,N_8786,N_8612);
nor U8981 (N_8981,N_8733,N_8748);
nor U8982 (N_8982,N_8678,N_8649);
nand U8983 (N_8983,N_8706,N_8673);
nor U8984 (N_8984,N_8716,N_8759);
nand U8985 (N_8985,N_8718,N_8620);
nand U8986 (N_8986,N_8630,N_8632);
nand U8987 (N_8987,N_8754,N_8683);
nand U8988 (N_8988,N_8625,N_8640);
and U8989 (N_8989,N_8641,N_8748);
or U8990 (N_8990,N_8732,N_8647);
nand U8991 (N_8991,N_8615,N_8641);
and U8992 (N_8992,N_8690,N_8773);
nand U8993 (N_8993,N_8791,N_8767);
or U8994 (N_8994,N_8798,N_8785);
and U8995 (N_8995,N_8788,N_8724);
xnor U8996 (N_8996,N_8739,N_8780);
nand U8997 (N_8997,N_8627,N_8697);
and U8998 (N_8998,N_8739,N_8775);
or U8999 (N_8999,N_8722,N_8716);
xnor U9000 (N_9000,N_8879,N_8984);
nor U9001 (N_9001,N_8847,N_8890);
xnor U9002 (N_9002,N_8924,N_8841);
nand U9003 (N_9003,N_8848,N_8878);
and U9004 (N_9004,N_8805,N_8885);
or U9005 (N_9005,N_8970,N_8854);
nor U9006 (N_9006,N_8936,N_8827);
and U9007 (N_9007,N_8903,N_8916);
and U9008 (N_9008,N_8876,N_8851);
nor U9009 (N_9009,N_8800,N_8837);
or U9010 (N_9010,N_8844,N_8815);
and U9011 (N_9011,N_8823,N_8835);
nor U9012 (N_9012,N_8930,N_8956);
nor U9013 (N_9013,N_8821,N_8958);
nor U9014 (N_9014,N_8980,N_8822);
or U9015 (N_9015,N_8873,N_8863);
nand U9016 (N_9016,N_8898,N_8866);
nand U9017 (N_9017,N_8889,N_8964);
xnor U9018 (N_9018,N_8920,N_8950);
nand U9019 (N_9019,N_8975,N_8952);
nor U9020 (N_9020,N_8824,N_8908);
nor U9021 (N_9021,N_8957,N_8902);
and U9022 (N_9022,N_8869,N_8846);
nor U9023 (N_9023,N_8899,N_8808);
and U9024 (N_9024,N_8927,N_8928);
or U9025 (N_9025,N_8926,N_8959);
xor U9026 (N_9026,N_8995,N_8922);
or U9027 (N_9027,N_8949,N_8812);
and U9028 (N_9028,N_8974,N_8921);
nor U9029 (N_9029,N_8883,N_8891);
nand U9030 (N_9030,N_8807,N_8840);
xor U9031 (N_9031,N_8831,N_8867);
and U9032 (N_9032,N_8945,N_8991);
nor U9033 (N_9033,N_8826,N_8990);
nor U9034 (N_9034,N_8986,N_8895);
nand U9035 (N_9035,N_8853,N_8966);
or U9036 (N_9036,N_8858,N_8967);
or U9037 (N_9037,N_8977,N_8850);
and U9038 (N_9038,N_8989,N_8955);
xnor U9039 (N_9039,N_8997,N_8894);
or U9040 (N_9040,N_8968,N_8913);
or U9041 (N_9041,N_8910,N_8836);
nand U9042 (N_9042,N_8811,N_8849);
nor U9043 (N_9043,N_8816,N_8804);
xnor U9044 (N_9044,N_8877,N_8829);
and U9045 (N_9045,N_8972,N_8855);
nor U9046 (N_9046,N_8982,N_8994);
and U9047 (N_9047,N_8919,N_8834);
or U9048 (N_9048,N_8999,N_8888);
nand U9049 (N_9049,N_8939,N_8833);
and U9050 (N_9050,N_8884,N_8944);
nor U9051 (N_9051,N_8985,N_8828);
nor U9052 (N_9052,N_8947,N_8933);
nand U9053 (N_9053,N_8880,N_8806);
or U9054 (N_9054,N_8983,N_8988);
nand U9055 (N_9055,N_8923,N_8912);
nand U9056 (N_9056,N_8810,N_8875);
nand U9057 (N_9057,N_8872,N_8864);
and U9058 (N_9058,N_8900,N_8857);
nand U9059 (N_9059,N_8915,N_8971);
or U9060 (N_9060,N_8932,N_8809);
nand U9061 (N_9061,N_8976,N_8992);
or U9062 (N_9062,N_8813,N_8937);
nor U9063 (N_9063,N_8830,N_8998);
or U9064 (N_9064,N_8881,N_8860);
nand U9065 (N_9065,N_8925,N_8814);
nor U9066 (N_9066,N_8819,N_8973);
nand U9067 (N_9067,N_8852,N_8948);
nor U9068 (N_9068,N_8859,N_8802);
or U9069 (N_9069,N_8901,N_8868);
nor U9070 (N_9070,N_8882,N_8963);
xnor U9071 (N_9071,N_8871,N_8865);
or U9072 (N_9072,N_8861,N_8941);
and U9073 (N_9073,N_8832,N_8942);
nand U9074 (N_9074,N_8951,N_8918);
xnor U9075 (N_9075,N_8934,N_8979);
nor U9076 (N_9076,N_8896,N_8962);
nand U9077 (N_9077,N_8820,N_8993);
nand U9078 (N_9078,N_8801,N_8935);
or U9079 (N_9079,N_8961,N_8892);
nor U9080 (N_9080,N_8917,N_8843);
and U9081 (N_9081,N_8987,N_8818);
or U9082 (N_9082,N_8996,N_8938);
nand U9083 (N_9083,N_8906,N_8943);
or U9084 (N_9084,N_8960,N_8978);
nor U9085 (N_9085,N_8825,N_8904);
nand U9086 (N_9086,N_8954,N_8897);
and U9087 (N_9087,N_8856,N_8838);
nand U9088 (N_9088,N_8874,N_8907);
or U9089 (N_9089,N_8862,N_8803);
nor U9090 (N_9090,N_8929,N_8870);
nand U9091 (N_9091,N_8931,N_8953);
and U9092 (N_9092,N_8965,N_8914);
nand U9093 (N_9093,N_8969,N_8911);
nor U9094 (N_9094,N_8893,N_8981);
nor U9095 (N_9095,N_8946,N_8886);
or U9096 (N_9096,N_8887,N_8905);
xor U9097 (N_9097,N_8940,N_8845);
nand U9098 (N_9098,N_8817,N_8839);
nand U9099 (N_9099,N_8909,N_8842);
nand U9100 (N_9100,N_8894,N_8873);
nor U9101 (N_9101,N_8968,N_8839);
or U9102 (N_9102,N_8822,N_8877);
nor U9103 (N_9103,N_8855,N_8932);
and U9104 (N_9104,N_8976,N_8952);
nor U9105 (N_9105,N_8943,N_8915);
and U9106 (N_9106,N_8818,N_8952);
xor U9107 (N_9107,N_8980,N_8886);
xor U9108 (N_9108,N_8953,N_8969);
xor U9109 (N_9109,N_8860,N_8808);
or U9110 (N_9110,N_8869,N_8848);
and U9111 (N_9111,N_8831,N_8994);
and U9112 (N_9112,N_8950,N_8944);
and U9113 (N_9113,N_8842,N_8928);
nor U9114 (N_9114,N_8829,N_8922);
nand U9115 (N_9115,N_8952,N_8963);
nand U9116 (N_9116,N_8813,N_8923);
xor U9117 (N_9117,N_8938,N_8886);
nand U9118 (N_9118,N_8865,N_8876);
or U9119 (N_9119,N_8884,N_8802);
nor U9120 (N_9120,N_8857,N_8841);
xor U9121 (N_9121,N_8935,N_8895);
and U9122 (N_9122,N_8810,N_8907);
or U9123 (N_9123,N_8835,N_8916);
xor U9124 (N_9124,N_8854,N_8922);
nor U9125 (N_9125,N_8872,N_8977);
and U9126 (N_9126,N_8827,N_8992);
or U9127 (N_9127,N_8873,N_8964);
xor U9128 (N_9128,N_8801,N_8989);
or U9129 (N_9129,N_8930,N_8989);
nand U9130 (N_9130,N_8968,N_8820);
nor U9131 (N_9131,N_8949,N_8955);
and U9132 (N_9132,N_8897,N_8832);
or U9133 (N_9133,N_8942,N_8876);
xor U9134 (N_9134,N_8854,N_8928);
or U9135 (N_9135,N_8989,N_8808);
nor U9136 (N_9136,N_8976,N_8827);
or U9137 (N_9137,N_8986,N_8841);
xor U9138 (N_9138,N_8938,N_8926);
and U9139 (N_9139,N_8992,N_8898);
nand U9140 (N_9140,N_8813,N_8855);
or U9141 (N_9141,N_8968,N_8907);
nand U9142 (N_9142,N_8903,N_8966);
nand U9143 (N_9143,N_8964,N_8896);
or U9144 (N_9144,N_8895,N_8959);
or U9145 (N_9145,N_8929,N_8907);
nand U9146 (N_9146,N_8930,N_8962);
nand U9147 (N_9147,N_8815,N_8969);
nand U9148 (N_9148,N_8972,N_8995);
and U9149 (N_9149,N_8929,N_8813);
and U9150 (N_9150,N_8954,N_8987);
nand U9151 (N_9151,N_8845,N_8805);
nor U9152 (N_9152,N_8827,N_8896);
or U9153 (N_9153,N_8806,N_8945);
nor U9154 (N_9154,N_8846,N_8897);
or U9155 (N_9155,N_8925,N_8953);
nor U9156 (N_9156,N_8939,N_8972);
or U9157 (N_9157,N_8937,N_8941);
nand U9158 (N_9158,N_8887,N_8827);
nor U9159 (N_9159,N_8952,N_8857);
xor U9160 (N_9160,N_8880,N_8827);
nor U9161 (N_9161,N_8925,N_8928);
nor U9162 (N_9162,N_8962,N_8910);
nor U9163 (N_9163,N_8885,N_8829);
nand U9164 (N_9164,N_8837,N_8953);
nor U9165 (N_9165,N_8994,N_8808);
and U9166 (N_9166,N_8867,N_8946);
nor U9167 (N_9167,N_8873,N_8817);
nor U9168 (N_9168,N_8846,N_8838);
nand U9169 (N_9169,N_8904,N_8927);
nand U9170 (N_9170,N_8961,N_8900);
nand U9171 (N_9171,N_8845,N_8921);
nand U9172 (N_9172,N_8910,N_8922);
or U9173 (N_9173,N_8811,N_8949);
or U9174 (N_9174,N_8987,N_8861);
or U9175 (N_9175,N_8938,N_8823);
nand U9176 (N_9176,N_8880,N_8808);
nor U9177 (N_9177,N_8830,N_8935);
nor U9178 (N_9178,N_8819,N_8993);
or U9179 (N_9179,N_8969,N_8864);
xnor U9180 (N_9180,N_8890,N_8807);
or U9181 (N_9181,N_8800,N_8890);
xnor U9182 (N_9182,N_8925,N_8957);
nand U9183 (N_9183,N_8860,N_8878);
nand U9184 (N_9184,N_8925,N_8913);
nor U9185 (N_9185,N_8919,N_8914);
xnor U9186 (N_9186,N_8926,N_8964);
nor U9187 (N_9187,N_8846,N_8933);
xnor U9188 (N_9188,N_8844,N_8997);
and U9189 (N_9189,N_8855,N_8887);
or U9190 (N_9190,N_8926,N_8899);
nor U9191 (N_9191,N_8897,N_8940);
xor U9192 (N_9192,N_8921,N_8872);
or U9193 (N_9193,N_8876,N_8853);
nand U9194 (N_9194,N_8932,N_8974);
nand U9195 (N_9195,N_8836,N_8878);
nand U9196 (N_9196,N_8953,N_8961);
nand U9197 (N_9197,N_8991,N_8898);
nor U9198 (N_9198,N_8997,N_8904);
nand U9199 (N_9199,N_8805,N_8855);
nor U9200 (N_9200,N_9042,N_9135);
or U9201 (N_9201,N_9075,N_9009);
and U9202 (N_9202,N_9149,N_9165);
nor U9203 (N_9203,N_9027,N_9024);
xor U9204 (N_9204,N_9010,N_9020);
or U9205 (N_9205,N_9188,N_9038);
nor U9206 (N_9206,N_9043,N_9013);
and U9207 (N_9207,N_9054,N_9172);
nor U9208 (N_9208,N_9176,N_9088);
and U9209 (N_9209,N_9130,N_9062);
nor U9210 (N_9210,N_9103,N_9067);
or U9211 (N_9211,N_9193,N_9004);
nand U9212 (N_9212,N_9059,N_9154);
xnor U9213 (N_9213,N_9179,N_9034);
and U9214 (N_9214,N_9019,N_9197);
or U9215 (N_9215,N_9146,N_9106);
or U9216 (N_9216,N_9091,N_9195);
nor U9217 (N_9217,N_9046,N_9008);
or U9218 (N_9218,N_9095,N_9039);
and U9219 (N_9219,N_9052,N_9119);
nor U9220 (N_9220,N_9035,N_9000);
and U9221 (N_9221,N_9156,N_9109);
nor U9222 (N_9222,N_9050,N_9087);
nor U9223 (N_9223,N_9073,N_9163);
and U9224 (N_9224,N_9180,N_9147);
and U9225 (N_9225,N_9061,N_9001);
and U9226 (N_9226,N_9151,N_9033);
xor U9227 (N_9227,N_9139,N_9032);
and U9228 (N_9228,N_9123,N_9170);
nor U9229 (N_9229,N_9047,N_9101);
nand U9230 (N_9230,N_9006,N_9072);
or U9231 (N_9231,N_9093,N_9028);
nand U9232 (N_9232,N_9069,N_9026);
nand U9233 (N_9233,N_9185,N_9074);
xor U9234 (N_9234,N_9107,N_9196);
nand U9235 (N_9235,N_9175,N_9153);
nor U9236 (N_9236,N_9079,N_9015);
and U9237 (N_9237,N_9104,N_9124);
or U9238 (N_9238,N_9187,N_9048);
and U9239 (N_9239,N_9071,N_9164);
or U9240 (N_9240,N_9127,N_9171);
nand U9241 (N_9241,N_9122,N_9105);
nand U9242 (N_9242,N_9118,N_9114);
nor U9243 (N_9243,N_9082,N_9057);
and U9244 (N_9244,N_9076,N_9159);
xnor U9245 (N_9245,N_9022,N_9150);
xor U9246 (N_9246,N_9060,N_9140);
nor U9247 (N_9247,N_9128,N_9141);
or U9248 (N_9248,N_9007,N_9162);
or U9249 (N_9249,N_9066,N_9189);
and U9250 (N_9250,N_9014,N_9194);
or U9251 (N_9251,N_9192,N_9112);
or U9252 (N_9252,N_9056,N_9111);
nand U9253 (N_9253,N_9025,N_9148);
nand U9254 (N_9254,N_9102,N_9068);
and U9255 (N_9255,N_9113,N_9177);
nand U9256 (N_9256,N_9011,N_9155);
xor U9257 (N_9257,N_9160,N_9115);
nand U9258 (N_9258,N_9086,N_9126);
nand U9259 (N_9259,N_9044,N_9016);
nor U9260 (N_9260,N_9186,N_9051);
or U9261 (N_9261,N_9045,N_9178);
nor U9262 (N_9262,N_9023,N_9167);
xnor U9263 (N_9263,N_9003,N_9083);
or U9264 (N_9264,N_9117,N_9081);
and U9265 (N_9265,N_9037,N_9089);
or U9266 (N_9266,N_9136,N_9173);
and U9267 (N_9267,N_9152,N_9058);
nor U9268 (N_9268,N_9096,N_9134);
or U9269 (N_9269,N_9182,N_9161);
or U9270 (N_9270,N_9005,N_9078);
nand U9271 (N_9271,N_9142,N_9132);
and U9272 (N_9272,N_9110,N_9129);
nor U9273 (N_9273,N_9121,N_9157);
or U9274 (N_9274,N_9018,N_9090);
nor U9275 (N_9275,N_9064,N_9097);
and U9276 (N_9276,N_9137,N_9131);
and U9277 (N_9277,N_9065,N_9098);
xor U9278 (N_9278,N_9031,N_9184);
xor U9279 (N_9279,N_9191,N_9092);
xnor U9280 (N_9280,N_9190,N_9125);
nor U9281 (N_9281,N_9198,N_9077);
nor U9282 (N_9282,N_9116,N_9174);
nor U9283 (N_9283,N_9012,N_9166);
xnor U9284 (N_9284,N_9080,N_9145);
nand U9285 (N_9285,N_9084,N_9183);
and U9286 (N_9286,N_9100,N_9143);
nor U9287 (N_9287,N_9199,N_9094);
nand U9288 (N_9288,N_9030,N_9169);
or U9289 (N_9289,N_9053,N_9168);
nor U9290 (N_9290,N_9138,N_9040);
and U9291 (N_9291,N_9036,N_9002);
nand U9292 (N_9292,N_9120,N_9133);
nand U9293 (N_9293,N_9158,N_9055);
or U9294 (N_9294,N_9181,N_9041);
or U9295 (N_9295,N_9029,N_9017);
and U9296 (N_9296,N_9049,N_9085);
nor U9297 (N_9297,N_9108,N_9063);
nor U9298 (N_9298,N_9144,N_9099);
or U9299 (N_9299,N_9021,N_9070);
nand U9300 (N_9300,N_9163,N_9107);
and U9301 (N_9301,N_9158,N_9007);
nand U9302 (N_9302,N_9037,N_9131);
and U9303 (N_9303,N_9199,N_9099);
or U9304 (N_9304,N_9013,N_9034);
nor U9305 (N_9305,N_9075,N_9190);
or U9306 (N_9306,N_9131,N_9004);
nand U9307 (N_9307,N_9123,N_9084);
nor U9308 (N_9308,N_9155,N_9186);
nor U9309 (N_9309,N_9075,N_9193);
nor U9310 (N_9310,N_9140,N_9135);
or U9311 (N_9311,N_9068,N_9079);
or U9312 (N_9312,N_9191,N_9073);
nor U9313 (N_9313,N_9055,N_9122);
nand U9314 (N_9314,N_9050,N_9164);
xnor U9315 (N_9315,N_9010,N_9123);
nand U9316 (N_9316,N_9145,N_9046);
nand U9317 (N_9317,N_9187,N_9190);
or U9318 (N_9318,N_9169,N_9052);
nand U9319 (N_9319,N_9043,N_9145);
nor U9320 (N_9320,N_9070,N_9077);
or U9321 (N_9321,N_9116,N_9027);
nand U9322 (N_9322,N_9191,N_9145);
nor U9323 (N_9323,N_9058,N_9062);
nand U9324 (N_9324,N_9172,N_9169);
or U9325 (N_9325,N_9186,N_9069);
nor U9326 (N_9326,N_9106,N_9171);
or U9327 (N_9327,N_9128,N_9152);
xnor U9328 (N_9328,N_9044,N_9065);
or U9329 (N_9329,N_9024,N_9016);
nor U9330 (N_9330,N_9117,N_9157);
or U9331 (N_9331,N_9054,N_9134);
and U9332 (N_9332,N_9021,N_9178);
and U9333 (N_9333,N_9089,N_9119);
nand U9334 (N_9334,N_9006,N_9109);
xnor U9335 (N_9335,N_9163,N_9092);
nor U9336 (N_9336,N_9094,N_9138);
or U9337 (N_9337,N_9157,N_9001);
and U9338 (N_9338,N_9086,N_9184);
and U9339 (N_9339,N_9189,N_9167);
and U9340 (N_9340,N_9091,N_9030);
and U9341 (N_9341,N_9076,N_9062);
xnor U9342 (N_9342,N_9131,N_9019);
nor U9343 (N_9343,N_9106,N_9013);
or U9344 (N_9344,N_9119,N_9026);
and U9345 (N_9345,N_9175,N_9091);
nand U9346 (N_9346,N_9052,N_9062);
or U9347 (N_9347,N_9066,N_9092);
and U9348 (N_9348,N_9163,N_9180);
or U9349 (N_9349,N_9047,N_9019);
nand U9350 (N_9350,N_9075,N_9058);
nor U9351 (N_9351,N_9033,N_9123);
nand U9352 (N_9352,N_9041,N_9134);
and U9353 (N_9353,N_9166,N_9057);
nor U9354 (N_9354,N_9172,N_9167);
nor U9355 (N_9355,N_9107,N_9065);
and U9356 (N_9356,N_9061,N_9085);
or U9357 (N_9357,N_9094,N_9044);
nor U9358 (N_9358,N_9127,N_9132);
or U9359 (N_9359,N_9172,N_9047);
xor U9360 (N_9360,N_9188,N_9054);
nor U9361 (N_9361,N_9140,N_9151);
and U9362 (N_9362,N_9070,N_9101);
nor U9363 (N_9363,N_9001,N_9040);
nor U9364 (N_9364,N_9124,N_9109);
nand U9365 (N_9365,N_9139,N_9128);
nor U9366 (N_9366,N_9136,N_9027);
nand U9367 (N_9367,N_9035,N_9089);
nor U9368 (N_9368,N_9137,N_9036);
nor U9369 (N_9369,N_9123,N_9103);
nand U9370 (N_9370,N_9124,N_9158);
and U9371 (N_9371,N_9117,N_9020);
and U9372 (N_9372,N_9198,N_9007);
xnor U9373 (N_9373,N_9182,N_9132);
or U9374 (N_9374,N_9188,N_9013);
and U9375 (N_9375,N_9006,N_9007);
or U9376 (N_9376,N_9086,N_9164);
nand U9377 (N_9377,N_9185,N_9132);
nor U9378 (N_9378,N_9110,N_9091);
nor U9379 (N_9379,N_9109,N_9087);
and U9380 (N_9380,N_9158,N_9156);
or U9381 (N_9381,N_9090,N_9109);
nor U9382 (N_9382,N_9141,N_9138);
and U9383 (N_9383,N_9084,N_9069);
nand U9384 (N_9384,N_9183,N_9151);
nand U9385 (N_9385,N_9024,N_9137);
nor U9386 (N_9386,N_9187,N_9198);
xor U9387 (N_9387,N_9034,N_9128);
nor U9388 (N_9388,N_9070,N_9099);
xnor U9389 (N_9389,N_9125,N_9100);
nor U9390 (N_9390,N_9020,N_9144);
or U9391 (N_9391,N_9006,N_9167);
nor U9392 (N_9392,N_9180,N_9187);
or U9393 (N_9393,N_9074,N_9194);
and U9394 (N_9394,N_9124,N_9184);
and U9395 (N_9395,N_9041,N_9006);
nand U9396 (N_9396,N_9124,N_9099);
nand U9397 (N_9397,N_9186,N_9001);
nor U9398 (N_9398,N_9059,N_9179);
and U9399 (N_9399,N_9061,N_9107);
nor U9400 (N_9400,N_9302,N_9304);
nor U9401 (N_9401,N_9316,N_9251);
xnor U9402 (N_9402,N_9318,N_9298);
or U9403 (N_9403,N_9305,N_9334);
nand U9404 (N_9404,N_9257,N_9247);
nor U9405 (N_9405,N_9208,N_9269);
and U9406 (N_9406,N_9300,N_9223);
nand U9407 (N_9407,N_9341,N_9295);
and U9408 (N_9408,N_9323,N_9356);
nor U9409 (N_9409,N_9277,N_9265);
nor U9410 (N_9410,N_9301,N_9330);
nor U9411 (N_9411,N_9350,N_9239);
xor U9412 (N_9412,N_9259,N_9238);
nor U9413 (N_9413,N_9253,N_9262);
nand U9414 (N_9414,N_9271,N_9266);
nor U9415 (N_9415,N_9307,N_9285);
and U9416 (N_9416,N_9267,N_9201);
nor U9417 (N_9417,N_9320,N_9327);
nand U9418 (N_9418,N_9210,N_9399);
or U9419 (N_9419,N_9311,N_9237);
xnor U9420 (N_9420,N_9248,N_9263);
or U9421 (N_9421,N_9335,N_9333);
nor U9422 (N_9422,N_9336,N_9383);
xnor U9423 (N_9423,N_9338,N_9264);
nand U9424 (N_9424,N_9296,N_9369);
and U9425 (N_9425,N_9309,N_9227);
nand U9426 (N_9426,N_9236,N_9331);
and U9427 (N_9427,N_9293,N_9358);
nor U9428 (N_9428,N_9287,N_9380);
or U9429 (N_9429,N_9289,N_9219);
nand U9430 (N_9430,N_9349,N_9211);
and U9431 (N_9431,N_9291,N_9243);
and U9432 (N_9432,N_9270,N_9315);
nor U9433 (N_9433,N_9368,N_9379);
and U9434 (N_9434,N_9241,N_9205);
xnor U9435 (N_9435,N_9272,N_9260);
nand U9436 (N_9436,N_9202,N_9216);
nand U9437 (N_9437,N_9206,N_9340);
nand U9438 (N_9438,N_9337,N_9360);
nand U9439 (N_9439,N_9240,N_9348);
and U9440 (N_9440,N_9388,N_9200);
or U9441 (N_9441,N_9365,N_9393);
nand U9442 (N_9442,N_9235,N_9342);
and U9443 (N_9443,N_9308,N_9203);
and U9444 (N_9444,N_9362,N_9396);
or U9445 (N_9445,N_9389,N_9347);
nor U9446 (N_9446,N_9273,N_9283);
nor U9447 (N_9447,N_9366,N_9268);
or U9448 (N_9448,N_9286,N_9261);
or U9449 (N_9449,N_9317,N_9225);
and U9450 (N_9450,N_9250,N_9370);
nand U9451 (N_9451,N_9312,N_9246);
nor U9452 (N_9452,N_9367,N_9221);
nand U9453 (N_9453,N_9339,N_9242);
xnor U9454 (N_9454,N_9215,N_9230);
nand U9455 (N_9455,N_9325,N_9288);
nand U9456 (N_9456,N_9256,N_9382);
and U9457 (N_9457,N_9294,N_9249);
xor U9458 (N_9458,N_9274,N_9281);
nor U9459 (N_9459,N_9279,N_9233);
or U9460 (N_9460,N_9390,N_9321);
nand U9461 (N_9461,N_9359,N_9232);
or U9462 (N_9462,N_9361,N_9324);
nor U9463 (N_9463,N_9231,N_9234);
nor U9464 (N_9464,N_9376,N_9299);
nand U9465 (N_9465,N_9378,N_9397);
xor U9466 (N_9466,N_9212,N_9353);
nand U9467 (N_9467,N_9275,N_9292);
or U9468 (N_9468,N_9213,N_9313);
or U9469 (N_9469,N_9254,N_9386);
nand U9470 (N_9470,N_9391,N_9229);
nand U9471 (N_9471,N_9354,N_9258);
nand U9472 (N_9472,N_9282,N_9314);
nand U9473 (N_9473,N_9375,N_9297);
nor U9474 (N_9474,N_9343,N_9384);
nor U9475 (N_9475,N_9371,N_9398);
nand U9476 (N_9476,N_9204,N_9351);
and U9477 (N_9477,N_9328,N_9310);
xnor U9478 (N_9478,N_9306,N_9374);
nor U9479 (N_9479,N_9220,N_9345);
nand U9480 (N_9480,N_9303,N_9395);
nand U9481 (N_9481,N_9226,N_9363);
or U9482 (N_9482,N_9373,N_9355);
or U9483 (N_9483,N_9290,N_9245);
and U9484 (N_9484,N_9392,N_9329);
and U9485 (N_9485,N_9332,N_9387);
or U9486 (N_9486,N_9278,N_9364);
nor U9487 (N_9487,N_9352,N_9381);
nand U9488 (N_9488,N_9385,N_9218);
nor U9489 (N_9489,N_9209,N_9222);
or U9490 (N_9490,N_9357,N_9284);
and U9491 (N_9491,N_9280,N_9344);
nand U9492 (N_9492,N_9346,N_9326);
nand U9493 (N_9493,N_9224,N_9276);
or U9494 (N_9494,N_9252,N_9228);
or U9495 (N_9495,N_9244,N_9319);
or U9496 (N_9496,N_9394,N_9217);
xnor U9497 (N_9497,N_9372,N_9255);
nand U9498 (N_9498,N_9214,N_9322);
and U9499 (N_9499,N_9377,N_9207);
or U9500 (N_9500,N_9379,N_9347);
or U9501 (N_9501,N_9203,N_9386);
nor U9502 (N_9502,N_9233,N_9253);
nor U9503 (N_9503,N_9348,N_9295);
nand U9504 (N_9504,N_9240,N_9276);
or U9505 (N_9505,N_9251,N_9314);
nor U9506 (N_9506,N_9303,N_9390);
or U9507 (N_9507,N_9226,N_9323);
and U9508 (N_9508,N_9201,N_9229);
and U9509 (N_9509,N_9216,N_9339);
nand U9510 (N_9510,N_9237,N_9293);
nand U9511 (N_9511,N_9388,N_9228);
nor U9512 (N_9512,N_9203,N_9246);
or U9513 (N_9513,N_9337,N_9323);
xor U9514 (N_9514,N_9209,N_9333);
nand U9515 (N_9515,N_9332,N_9365);
nand U9516 (N_9516,N_9320,N_9227);
or U9517 (N_9517,N_9386,N_9358);
and U9518 (N_9518,N_9216,N_9218);
nand U9519 (N_9519,N_9267,N_9369);
nor U9520 (N_9520,N_9308,N_9318);
nand U9521 (N_9521,N_9336,N_9374);
or U9522 (N_9522,N_9334,N_9294);
or U9523 (N_9523,N_9224,N_9268);
or U9524 (N_9524,N_9265,N_9320);
nor U9525 (N_9525,N_9204,N_9359);
nand U9526 (N_9526,N_9231,N_9273);
nor U9527 (N_9527,N_9229,N_9364);
nand U9528 (N_9528,N_9258,N_9358);
xor U9529 (N_9529,N_9225,N_9346);
nand U9530 (N_9530,N_9399,N_9332);
nor U9531 (N_9531,N_9211,N_9223);
or U9532 (N_9532,N_9351,N_9254);
nor U9533 (N_9533,N_9245,N_9229);
nand U9534 (N_9534,N_9316,N_9387);
nor U9535 (N_9535,N_9208,N_9291);
or U9536 (N_9536,N_9349,N_9228);
nand U9537 (N_9537,N_9302,N_9276);
nor U9538 (N_9538,N_9236,N_9387);
nand U9539 (N_9539,N_9354,N_9274);
xor U9540 (N_9540,N_9377,N_9383);
nor U9541 (N_9541,N_9239,N_9374);
nor U9542 (N_9542,N_9246,N_9279);
and U9543 (N_9543,N_9375,N_9341);
and U9544 (N_9544,N_9242,N_9356);
xor U9545 (N_9545,N_9353,N_9279);
nand U9546 (N_9546,N_9303,N_9300);
nand U9547 (N_9547,N_9313,N_9397);
nor U9548 (N_9548,N_9208,N_9310);
or U9549 (N_9549,N_9260,N_9329);
or U9550 (N_9550,N_9323,N_9210);
xnor U9551 (N_9551,N_9276,N_9292);
nor U9552 (N_9552,N_9225,N_9223);
nand U9553 (N_9553,N_9215,N_9229);
nor U9554 (N_9554,N_9204,N_9360);
or U9555 (N_9555,N_9213,N_9319);
or U9556 (N_9556,N_9271,N_9231);
nor U9557 (N_9557,N_9359,N_9283);
nand U9558 (N_9558,N_9387,N_9339);
and U9559 (N_9559,N_9328,N_9261);
nor U9560 (N_9560,N_9333,N_9229);
nand U9561 (N_9561,N_9213,N_9201);
nand U9562 (N_9562,N_9231,N_9392);
and U9563 (N_9563,N_9278,N_9244);
and U9564 (N_9564,N_9256,N_9344);
or U9565 (N_9565,N_9399,N_9386);
nor U9566 (N_9566,N_9333,N_9250);
or U9567 (N_9567,N_9355,N_9310);
nor U9568 (N_9568,N_9332,N_9389);
nor U9569 (N_9569,N_9383,N_9281);
nand U9570 (N_9570,N_9208,N_9378);
nor U9571 (N_9571,N_9378,N_9398);
and U9572 (N_9572,N_9282,N_9369);
or U9573 (N_9573,N_9372,N_9273);
and U9574 (N_9574,N_9226,N_9218);
or U9575 (N_9575,N_9204,N_9290);
nand U9576 (N_9576,N_9281,N_9327);
nor U9577 (N_9577,N_9206,N_9375);
or U9578 (N_9578,N_9332,N_9383);
nor U9579 (N_9579,N_9332,N_9360);
xnor U9580 (N_9580,N_9377,N_9238);
or U9581 (N_9581,N_9352,N_9230);
nor U9582 (N_9582,N_9395,N_9313);
nor U9583 (N_9583,N_9374,N_9388);
or U9584 (N_9584,N_9357,N_9335);
nand U9585 (N_9585,N_9342,N_9283);
xor U9586 (N_9586,N_9312,N_9275);
and U9587 (N_9587,N_9259,N_9203);
nor U9588 (N_9588,N_9371,N_9348);
and U9589 (N_9589,N_9352,N_9294);
xor U9590 (N_9590,N_9231,N_9299);
and U9591 (N_9591,N_9337,N_9234);
and U9592 (N_9592,N_9281,N_9344);
nor U9593 (N_9593,N_9366,N_9308);
nand U9594 (N_9594,N_9216,N_9352);
or U9595 (N_9595,N_9298,N_9290);
nor U9596 (N_9596,N_9396,N_9240);
and U9597 (N_9597,N_9226,N_9289);
nand U9598 (N_9598,N_9381,N_9245);
nor U9599 (N_9599,N_9280,N_9281);
or U9600 (N_9600,N_9576,N_9521);
or U9601 (N_9601,N_9544,N_9407);
or U9602 (N_9602,N_9423,N_9542);
and U9603 (N_9603,N_9522,N_9588);
or U9604 (N_9604,N_9590,N_9532);
or U9605 (N_9605,N_9543,N_9553);
xnor U9606 (N_9606,N_9546,N_9431);
or U9607 (N_9607,N_9476,N_9402);
and U9608 (N_9608,N_9595,N_9533);
and U9609 (N_9609,N_9488,N_9578);
nor U9610 (N_9610,N_9490,N_9428);
xor U9611 (N_9611,N_9409,N_9561);
and U9612 (N_9612,N_9524,N_9458);
nor U9613 (N_9613,N_9404,N_9433);
nor U9614 (N_9614,N_9517,N_9591);
nor U9615 (N_9615,N_9523,N_9474);
or U9616 (N_9616,N_9504,N_9482);
and U9617 (N_9617,N_9440,N_9573);
or U9618 (N_9618,N_9405,N_9435);
nor U9619 (N_9619,N_9575,N_9587);
nand U9620 (N_9620,N_9468,N_9406);
nand U9621 (N_9621,N_9480,N_9548);
xor U9622 (N_9622,N_9471,N_9497);
and U9623 (N_9623,N_9502,N_9594);
or U9624 (N_9624,N_9493,N_9411);
or U9625 (N_9625,N_9410,N_9572);
nand U9626 (N_9626,N_9559,N_9537);
xnor U9627 (N_9627,N_9501,N_9489);
and U9628 (N_9628,N_9424,N_9432);
and U9629 (N_9629,N_9564,N_9413);
and U9630 (N_9630,N_9492,N_9447);
or U9631 (N_9631,N_9528,N_9421);
nand U9632 (N_9632,N_9512,N_9597);
nand U9633 (N_9633,N_9557,N_9584);
or U9634 (N_9634,N_9425,N_9535);
nand U9635 (N_9635,N_9509,N_9549);
xor U9636 (N_9636,N_9451,N_9454);
and U9637 (N_9637,N_9530,N_9519);
and U9638 (N_9638,N_9547,N_9516);
and U9639 (N_9639,N_9400,N_9531);
nand U9640 (N_9640,N_9477,N_9506);
and U9641 (N_9641,N_9463,N_9574);
nand U9642 (N_9642,N_9415,N_9426);
nand U9643 (N_9643,N_9438,N_9556);
xnor U9644 (N_9644,N_9526,N_9507);
and U9645 (N_9645,N_9586,N_9496);
nand U9646 (N_9646,N_9580,N_9518);
nand U9647 (N_9647,N_9419,N_9408);
nand U9648 (N_9648,N_9403,N_9429);
nand U9649 (N_9649,N_9520,N_9487);
or U9650 (N_9650,N_9481,N_9536);
nor U9651 (N_9651,N_9508,N_9446);
and U9652 (N_9652,N_9417,N_9486);
nand U9653 (N_9653,N_9484,N_9494);
and U9654 (N_9654,N_9585,N_9583);
or U9655 (N_9655,N_9568,N_9427);
xnor U9656 (N_9656,N_9453,N_9437);
nor U9657 (N_9657,N_9554,N_9498);
or U9658 (N_9658,N_9455,N_9460);
or U9659 (N_9659,N_9418,N_9420);
nor U9660 (N_9660,N_9558,N_9444);
nor U9661 (N_9661,N_9569,N_9450);
nand U9662 (N_9662,N_9469,N_9503);
and U9663 (N_9663,N_9430,N_9582);
or U9664 (N_9664,N_9511,N_9510);
and U9665 (N_9665,N_9434,N_9422);
or U9666 (N_9666,N_9565,N_9478);
nor U9667 (N_9667,N_9529,N_9527);
or U9668 (N_9668,N_9466,N_9445);
and U9669 (N_9669,N_9473,N_9540);
or U9670 (N_9670,N_9436,N_9514);
nor U9671 (N_9671,N_9525,N_9442);
nor U9672 (N_9672,N_9416,N_9462);
nor U9673 (N_9673,N_9441,N_9539);
or U9674 (N_9674,N_9593,N_9551);
nor U9675 (N_9675,N_9461,N_9571);
nand U9676 (N_9676,N_9599,N_9500);
or U9677 (N_9677,N_9550,N_9555);
nand U9678 (N_9678,N_9464,N_9491);
nor U9679 (N_9679,N_9513,N_9439);
nand U9680 (N_9680,N_9443,N_9459);
and U9681 (N_9681,N_9567,N_9560);
nor U9682 (N_9682,N_9505,N_9515);
xor U9683 (N_9683,N_9457,N_9412);
xor U9684 (N_9684,N_9589,N_9448);
or U9685 (N_9685,N_9401,N_9592);
and U9686 (N_9686,N_9541,N_9552);
or U9687 (N_9687,N_9570,N_9475);
nand U9688 (N_9688,N_9452,N_9449);
or U9689 (N_9689,N_9545,N_9414);
or U9690 (N_9690,N_9562,N_9538);
nand U9691 (N_9691,N_9579,N_9534);
or U9692 (N_9692,N_9495,N_9563);
nor U9693 (N_9693,N_9566,N_9596);
nand U9694 (N_9694,N_9485,N_9499);
xnor U9695 (N_9695,N_9581,N_9598);
and U9696 (N_9696,N_9479,N_9467);
nand U9697 (N_9697,N_9465,N_9577);
and U9698 (N_9698,N_9470,N_9456);
xor U9699 (N_9699,N_9483,N_9472);
and U9700 (N_9700,N_9404,N_9509);
and U9701 (N_9701,N_9419,N_9516);
nand U9702 (N_9702,N_9460,N_9504);
or U9703 (N_9703,N_9478,N_9512);
nor U9704 (N_9704,N_9595,N_9548);
nor U9705 (N_9705,N_9402,N_9572);
nor U9706 (N_9706,N_9578,N_9438);
nand U9707 (N_9707,N_9421,N_9544);
or U9708 (N_9708,N_9545,N_9551);
and U9709 (N_9709,N_9437,N_9477);
xor U9710 (N_9710,N_9588,N_9410);
or U9711 (N_9711,N_9562,N_9508);
nand U9712 (N_9712,N_9440,N_9401);
and U9713 (N_9713,N_9508,N_9423);
nand U9714 (N_9714,N_9444,N_9443);
nor U9715 (N_9715,N_9450,N_9486);
or U9716 (N_9716,N_9481,N_9497);
nor U9717 (N_9717,N_9528,N_9571);
nor U9718 (N_9718,N_9518,N_9491);
nand U9719 (N_9719,N_9507,N_9499);
xnor U9720 (N_9720,N_9438,N_9530);
nand U9721 (N_9721,N_9453,N_9458);
or U9722 (N_9722,N_9465,N_9547);
and U9723 (N_9723,N_9573,N_9582);
nand U9724 (N_9724,N_9527,N_9498);
nand U9725 (N_9725,N_9426,N_9551);
and U9726 (N_9726,N_9446,N_9520);
and U9727 (N_9727,N_9417,N_9548);
nand U9728 (N_9728,N_9516,N_9596);
nand U9729 (N_9729,N_9592,N_9569);
nor U9730 (N_9730,N_9536,N_9537);
nand U9731 (N_9731,N_9549,N_9476);
and U9732 (N_9732,N_9555,N_9476);
and U9733 (N_9733,N_9512,N_9502);
or U9734 (N_9734,N_9480,N_9469);
nor U9735 (N_9735,N_9501,N_9509);
or U9736 (N_9736,N_9594,N_9498);
nand U9737 (N_9737,N_9505,N_9406);
nand U9738 (N_9738,N_9583,N_9553);
nand U9739 (N_9739,N_9522,N_9445);
nor U9740 (N_9740,N_9518,N_9463);
or U9741 (N_9741,N_9411,N_9426);
and U9742 (N_9742,N_9409,N_9404);
and U9743 (N_9743,N_9427,N_9558);
nor U9744 (N_9744,N_9589,N_9423);
and U9745 (N_9745,N_9477,N_9494);
xor U9746 (N_9746,N_9461,N_9594);
or U9747 (N_9747,N_9492,N_9415);
nand U9748 (N_9748,N_9552,N_9550);
and U9749 (N_9749,N_9549,N_9543);
or U9750 (N_9750,N_9460,N_9445);
nand U9751 (N_9751,N_9413,N_9571);
nand U9752 (N_9752,N_9461,N_9472);
nand U9753 (N_9753,N_9411,N_9408);
and U9754 (N_9754,N_9538,N_9579);
and U9755 (N_9755,N_9451,N_9409);
nor U9756 (N_9756,N_9538,N_9520);
and U9757 (N_9757,N_9565,N_9404);
xor U9758 (N_9758,N_9495,N_9476);
nand U9759 (N_9759,N_9580,N_9503);
nand U9760 (N_9760,N_9564,N_9541);
and U9761 (N_9761,N_9436,N_9493);
or U9762 (N_9762,N_9412,N_9546);
or U9763 (N_9763,N_9456,N_9474);
and U9764 (N_9764,N_9514,N_9533);
nand U9765 (N_9765,N_9481,N_9542);
xnor U9766 (N_9766,N_9409,N_9599);
xor U9767 (N_9767,N_9555,N_9401);
or U9768 (N_9768,N_9525,N_9510);
nor U9769 (N_9769,N_9568,N_9401);
or U9770 (N_9770,N_9422,N_9545);
or U9771 (N_9771,N_9573,N_9535);
nand U9772 (N_9772,N_9465,N_9406);
nand U9773 (N_9773,N_9438,N_9440);
or U9774 (N_9774,N_9418,N_9477);
nand U9775 (N_9775,N_9552,N_9494);
nor U9776 (N_9776,N_9402,N_9580);
nor U9777 (N_9777,N_9594,N_9450);
nor U9778 (N_9778,N_9423,N_9597);
xor U9779 (N_9779,N_9576,N_9529);
and U9780 (N_9780,N_9579,N_9597);
nand U9781 (N_9781,N_9424,N_9489);
xnor U9782 (N_9782,N_9593,N_9498);
xnor U9783 (N_9783,N_9521,N_9568);
or U9784 (N_9784,N_9413,N_9548);
nand U9785 (N_9785,N_9544,N_9591);
nor U9786 (N_9786,N_9531,N_9445);
nor U9787 (N_9787,N_9584,N_9469);
or U9788 (N_9788,N_9572,N_9482);
and U9789 (N_9789,N_9413,N_9505);
nand U9790 (N_9790,N_9585,N_9517);
or U9791 (N_9791,N_9556,N_9503);
nand U9792 (N_9792,N_9420,N_9447);
nand U9793 (N_9793,N_9575,N_9540);
nand U9794 (N_9794,N_9558,N_9572);
nor U9795 (N_9795,N_9555,N_9444);
or U9796 (N_9796,N_9458,N_9491);
or U9797 (N_9797,N_9564,N_9489);
or U9798 (N_9798,N_9480,N_9514);
xor U9799 (N_9799,N_9446,N_9519);
xnor U9800 (N_9800,N_9705,N_9695);
or U9801 (N_9801,N_9636,N_9655);
or U9802 (N_9802,N_9605,N_9770);
nand U9803 (N_9803,N_9703,N_9672);
nor U9804 (N_9804,N_9778,N_9744);
xnor U9805 (N_9805,N_9661,N_9781);
and U9806 (N_9806,N_9696,N_9658);
or U9807 (N_9807,N_9742,N_9666);
nand U9808 (N_9808,N_9644,N_9759);
nor U9809 (N_9809,N_9775,N_9684);
nor U9810 (N_9810,N_9794,N_9632);
or U9811 (N_9811,N_9791,N_9761);
nand U9812 (N_9812,N_9714,N_9771);
nand U9813 (N_9813,N_9722,N_9740);
nand U9814 (N_9814,N_9693,N_9782);
or U9815 (N_9815,N_9765,N_9618);
and U9816 (N_9816,N_9685,N_9649);
or U9817 (N_9817,N_9709,N_9640);
or U9818 (N_9818,N_9739,N_9774);
and U9819 (N_9819,N_9698,N_9646);
or U9820 (N_9820,N_9736,N_9601);
nand U9821 (N_9821,N_9657,N_9699);
xnor U9822 (N_9822,N_9677,N_9788);
nor U9823 (N_9823,N_9762,N_9659);
nand U9824 (N_9824,N_9748,N_9756);
or U9825 (N_9825,N_9702,N_9647);
and U9826 (N_9826,N_9630,N_9634);
or U9827 (N_9827,N_9665,N_9627);
or U9828 (N_9828,N_9745,N_9613);
or U9829 (N_9829,N_9797,N_9680);
nor U9830 (N_9830,N_9713,N_9694);
nor U9831 (N_9831,N_9689,N_9681);
nor U9832 (N_9832,N_9668,N_9784);
nand U9833 (N_9833,N_9735,N_9607);
nand U9834 (N_9834,N_9795,N_9626);
xnor U9835 (N_9835,N_9608,N_9604);
nand U9836 (N_9836,N_9747,N_9673);
nor U9837 (N_9837,N_9741,N_9675);
and U9838 (N_9838,N_9653,N_9789);
nand U9839 (N_9839,N_9642,N_9746);
and U9840 (N_9840,N_9783,N_9757);
xnor U9841 (N_9841,N_9651,N_9737);
or U9842 (N_9842,N_9718,N_9753);
xor U9843 (N_9843,N_9780,N_9793);
nand U9844 (N_9844,N_9768,N_9615);
xor U9845 (N_9845,N_9663,N_9711);
or U9846 (N_9846,N_9719,N_9776);
nand U9847 (N_9847,N_9639,N_9790);
nor U9848 (N_9848,N_9717,N_9734);
nor U9849 (N_9849,N_9792,N_9750);
nand U9850 (N_9850,N_9725,N_9625);
and U9851 (N_9851,N_9716,N_9638);
or U9852 (N_9852,N_9715,N_9721);
nand U9853 (N_9853,N_9758,N_9671);
nand U9854 (N_9854,N_9660,N_9760);
nor U9855 (N_9855,N_9664,N_9621);
or U9856 (N_9856,N_9796,N_9690);
and U9857 (N_9857,N_9691,N_9611);
and U9858 (N_9858,N_9679,N_9706);
and U9859 (N_9859,N_9730,N_9674);
nor U9860 (N_9860,N_9752,N_9704);
nor U9861 (N_9861,N_9733,N_9624);
or U9862 (N_9862,N_9751,N_9799);
nor U9863 (N_9863,N_9612,N_9610);
or U9864 (N_9864,N_9631,N_9676);
or U9865 (N_9865,N_9738,N_9682);
and U9866 (N_9866,N_9620,N_9723);
or U9867 (N_9867,N_9688,N_9669);
nor U9868 (N_9868,N_9743,N_9654);
and U9869 (N_9869,N_9623,N_9633);
nand U9870 (N_9870,N_9769,N_9600);
or U9871 (N_9871,N_9645,N_9667);
xor U9872 (N_9872,N_9766,N_9701);
or U9873 (N_9873,N_9686,N_9777);
nand U9874 (N_9874,N_9798,N_9787);
nor U9875 (N_9875,N_9700,N_9652);
nor U9876 (N_9876,N_9606,N_9754);
xnor U9877 (N_9877,N_9720,N_9724);
nand U9878 (N_9878,N_9650,N_9628);
or U9879 (N_9879,N_9617,N_9637);
and U9880 (N_9880,N_9767,N_9629);
and U9881 (N_9881,N_9779,N_9764);
or U9882 (N_9882,N_9643,N_9619);
nand U9883 (N_9883,N_9603,N_9708);
nor U9884 (N_9884,N_9707,N_9728);
or U9885 (N_9885,N_9727,N_9749);
nand U9886 (N_9886,N_9763,N_9641);
and U9887 (N_9887,N_9662,N_9712);
and U9888 (N_9888,N_9710,N_9731);
nand U9889 (N_9889,N_9772,N_9670);
nor U9890 (N_9890,N_9609,N_9697);
nor U9891 (N_9891,N_9614,N_9678);
and U9892 (N_9892,N_9729,N_9692);
and U9893 (N_9893,N_9687,N_9635);
nor U9894 (N_9894,N_9726,N_9648);
xor U9895 (N_9895,N_9616,N_9602);
or U9896 (N_9896,N_9773,N_9786);
nand U9897 (N_9897,N_9755,N_9656);
and U9898 (N_9898,N_9683,N_9622);
nor U9899 (N_9899,N_9785,N_9732);
xnor U9900 (N_9900,N_9666,N_9788);
and U9901 (N_9901,N_9645,N_9780);
nor U9902 (N_9902,N_9637,N_9728);
nand U9903 (N_9903,N_9732,N_9638);
and U9904 (N_9904,N_9705,N_9767);
nand U9905 (N_9905,N_9759,N_9709);
and U9906 (N_9906,N_9721,N_9707);
xor U9907 (N_9907,N_9631,N_9718);
nand U9908 (N_9908,N_9727,N_9786);
and U9909 (N_9909,N_9657,N_9661);
or U9910 (N_9910,N_9722,N_9737);
xnor U9911 (N_9911,N_9769,N_9750);
nand U9912 (N_9912,N_9729,N_9615);
xnor U9913 (N_9913,N_9670,N_9769);
nor U9914 (N_9914,N_9757,N_9635);
xor U9915 (N_9915,N_9624,N_9662);
nor U9916 (N_9916,N_9732,N_9662);
and U9917 (N_9917,N_9673,N_9684);
and U9918 (N_9918,N_9639,N_9698);
or U9919 (N_9919,N_9615,N_9648);
nor U9920 (N_9920,N_9793,N_9666);
nand U9921 (N_9921,N_9714,N_9641);
and U9922 (N_9922,N_9713,N_9757);
nor U9923 (N_9923,N_9659,N_9696);
and U9924 (N_9924,N_9738,N_9715);
and U9925 (N_9925,N_9622,N_9788);
nand U9926 (N_9926,N_9681,N_9620);
or U9927 (N_9927,N_9650,N_9679);
or U9928 (N_9928,N_9665,N_9700);
xor U9929 (N_9929,N_9796,N_9668);
nand U9930 (N_9930,N_9724,N_9730);
nand U9931 (N_9931,N_9627,N_9716);
nand U9932 (N_9932,N_9650,N_9735);
nand U9933 (N_9933,N_9723,N_9771);
nor U9934 (N_9934,N_9651,N_9714);
or U9935 (N_9935,N_9645,N_9712);
and U9936 (N_9936,N_9764,N_9743);
and U9937 (N_9937,N_9779,N_9661);
or U9938 (N_9938,N_9691,N_9758);
nand U9939 (N_9939,N_9788,N_9602);
or U9940 (N_9940,N_9777,N_9780);
nor U9941 (N_9941,N_9720,N_9721);
nand U9942 (N_9942,N_9694,N_9741);
nor U9943 (N_9943,N_9733,N_9632);
nor U9944 (N_9944,N_9751,N_9721);
or U9945 (N_9945,N_9715,N_9733);
or U9946 (N_9946,N_9643,N_9608);
nor U9947 (N_9947,N_9707,N_9695);
nor U9948 (N_9948,N_9676,N_9709);
and U9949 (N_9949,N_9609,N_9733);
nor U9950 (N_9950,N_9734,N_9703);
and U9951 (N_9951,N_9615,N_9751);
and U9952 (N_9952,N_9675,N_9676);
or U9953 (N_9953,N_9708,N_9630);
xnor U9954 (N_9954,N_9650,N_9710);
and U9955 (N_9955,N_9639,N_9653);
or U9956 (N_9956,N_9608,N_9611);
and U9957 (N_9957,N_9793,N_9762);
nand U9958 (N_9958,N_9653,N_9680);
or U9959 (N_9959,N_9779,N_9775);
nand U9960 (N_9960,N_9629,N_9685);
and U9961 (N_9961,N_9649,N_9728);
nand U9962 (N_9962,N_9612,N_9630);
nand U9963 (N_9963,N_9616,N_9771);
and U9964 (N_9964,N_9754,N_9644);
or U9965 (N_9965,N_9743,N_9759);
and U9966 (N_9966,N_9718,N_9796);
nand U9967 (N_9967,N_9719,N_9641);
xnor U9968 (N_9968,N_9611,N_9687);
and U9969 (N_9969,N_9642,N_9610);
and U9970 (N_9970,N_9770,N_9771);
nor U9971 (N_9971,N_9661,N_9758);
or U9972 (N_9972,N_9765,N_9748);
or U9973 (N_9973,N_9770,N_9780);
nor U9974 (N_9974,N_9765,N_9647);
nor U9975 (N_9975,N_9784,N_9781);
or U9976 (N_9976,N_9649,N_9684);
or U9977 (N_9977,N_9675,N_9610);
and U9978 (N_9978,N_9740,N_9728);
nor U9979 (N_9979,N_9777,N_9710);
nor U9980 (N_9980,N_9797,N_9611);
nand U9981 (N_9981,N_9777,N_9629);
or U9982 (N_9982,N_9718,N_9698);
nand U9983 (N_9983,N_9613,N_9771);
and U9984 (N_9984,N_9698,N_9615);
or U9985 (N_9985,N_9721,N_9760);
nor U9986 (N_9986,N_9764,N_9682);
xnor U9987 (N_9987,N_9735,N_9619);
xnor U9988 (N_9988,N_9692,N_9723);
or U9989 (N_9989,N_9763,N_9770);
nor U9990 (N_9990,N_9790,N_9757);
and U9991 (N_9991,N_9797,N_9772);
nor U9992 (N_9992,N_9684,N_9642);
nand U9993 (N_9993,N_9763,N_9760);
and U9994 (N_9994,N_9604,N_9640);
xnor U9995 (N_9995,N_9601,N_9686);
and U9996 (N_9996,N_9762,N_9676);
nand U9997 (N_9997,N_9773,N_9706);
nor U9998 (N_9998,N_9781,N_9652);
nand U9999 (N_9999,N_9607,N_9718);
nor UO_0 (O_0,N_9870,N_9873);
xor UO_1 (O_1,N_9982,N_9891);
nor UO_2 (O_2,N_9963,N_9951);
or UO_3 (O_3,N_9867,N_9970);
nor UO_4 (O_4,N_9981,N_9997);
nor UO_5 (O_5,N_9857,N_9986);
nor UO_6 (O_6,N_9843,N_9854);
and UO_7 (O_7,N_9845,N_9800);
nor UO_8 (O_8,N_9937,N_9988);
xnor UO_9 (O_9,N_9846,N_9820);
and UO_10 (O_10,N_9905,N_9996);
nand UO_11 (O_11,N_9946,N_9999);
nand UO_12 (O_12,N_9862,N_9923);
or UO_13 (O_13,N_9825,N_9987);
nand UO_14 (O_14,N_9828,N_9859);
and UO_15 (O_15,N_9885,N_9932);
and UO_16 (O_16,N_9902,N_9934);
and UO_17 (O_17,N_9831,N_9917);
or UO_18 (O_18,N_9948,N_9864);
and UO_19 (O_19,N_9971,N_9847);
nand UO_20 (O_20,N_9962,N_9920);
nand UO_21 (O_21,N_9955,N_9874);
or UO_22 (O_22,N_9903,N_9892);
or UO_23 (O_23,N_9976,N_9939);
or UO_24 (O_24,N_9929,N_9816);
nand UO_25 (O_25,N_9813,N_9959);
nand UO_26 (O_26,N_9967,N_9991);
or UO_27 (O_27,N_9899,N_9918);
nor UO_28 (O_28,N_9925,N_9850);
nor UO_29 (O_29,N_9954,N_9868);
or UO_30 (O_30,N_9830,N_9840);
and UO_31 (O_31,N_9931,N_9882);
and UO_32 (O_32,N_9802,N_9936);
nand UO_33 (O_33,N_9832,N_9947);
nand UO_34 (O_34,N_9960,N_9860);
nand UO_35 (O_35,N_9992,N_9895);
and UO_36 (O_36,N_9863,N_9869);
and UO_37 (O_37,N_9945,N_9861);
and UO_38 (O_38,N_9814,N_9811);
nor UO_39 (O_39,N_9827,N_9819);
nand UO_40 (O_40,N_9834,N_9818);
or UO_41 (O_41,N_9896,N_9808);
nor UO_42 (O_42,N_9912,N_9995);
nor UO_43 (O_43,N_9964,N_9852);
nor UO_44 (O_44,N_9890,N_9836);
nor UO_45 (O_45,N_9810,N_9848);
and UO_46 (O_46,N_9907,N_9966);
and UO_47 (O_47,N_9875,N_9953);
nand UO_48 (O_48,N_9872,N_9911);
nand UO_49 (O_49,N_9849,N_9930);
nand UO_50 (O_50,N_9804,N_9985);
nand UO_51 (O_51,N_9821,N_9824);
or UO_52 (O_52,N_9965,N_9916);
and UO_53 (O_53,N_9806,N_9933);
nand UO_54 (O_54,N_9969,N_9958);
or UO_55 (O_55,N_9952,N_9866);
and UO_56 (O_56,N_9983,N_9858);
and UO_57 (O_57,N_9968,N_9943);
nor UO_58 (O_58,N_9941,N_9979);
and UO_59 (O_59,N_9877,N_9940);
nand UO_60 (O_60,N_9871,N_9927);
or UO_61 (O_61,N_9842,N_9922);
and UO_62 (O_62,N_9898,N_9928);
nor UO_63 (O_63,N_9812,N_9926);
nor UO_64 (O_64,N_9886,N_9980);
or UO_65 (O_65,N_9949,N_9910);
nand UO_66 (O_66,N_9826,N_9990);
nor UO_67 (O_67,N_9901,N_9961);
or UO_68 (O_68,N_9888,N_9919);
nand UO_69 (O_69,N_9974,N_9900);
nand UO_70 (O_70,N_9855,N_9909);
or UO_71 (O_71,N_9876,N_9889);
nand UO_72 (O_72,N_9984,N_9822);
or UO_73 (O_73,N_9880,N_9884);
xnor UO_74 (O_74,N_9829,N_9998);
and UO_75 (O_75,N_9839,N_9883);
or UO_76 (O_76,N_9881,N_9944);
nand UO_77 (O_77,N_9989,N_9835);
xnor UO_78 (O_78,N_9805,N_9833);
or UO_79 (O_79,N_9913,N_9865);
or UO_80 (O_80,N_9893,N_9915);
nor UO_81 (O_81,N_9977,N_9956);
xnor UO_82 (O_82,N_9879,N_9817);
nand UO_83 (O_83,N_9978,N_9908);
xor UO_84 (O_84,N_9975,N_9823);
nor UO_85 (O_85,N_9994,N_9942);
or UO_86 (O_86,N_9894,N_9921);
nor UO_87 (O_87,N_9837,N_9838);
nor UO_88 (O_88,N_9938,N_9972);
or UO_89 (O_89,N_9904,N_9801);
nor UO_90 (O_90,N_9887,N_9914);
and UO_91 (O_91,N_9856,N_9924);
nand UO_92 (O_92,N_9844,N_9897);
nand UO_93 (O_93,N_9851,N_9803);
xor UO_94 (O_94,N_9815,N_9973);
nand UO_95 (O_95,N_9809,N_9878);
or UO_96 (O_96,N_9950,N_9957);
nand UO_97 (O_97,N_9935,N_9807);
nor UO_98 (O_98,N_9853,N_9841);
nor UO_99 (O_99,N_9906,N_9993);
or UO_100 (O_100,N_9850,N_9800);
and UO_101 (O_101,N_9926,N_9913);
and UO_102 (O_102,N_9934,N_9946);
and UO_103 (O_103,N_9862,N_9934);
xor UO_104 (O_104,N_9998,N_9930);
and UO_105 (O_105,N_9864,N_9909);
nand UO_106 (O_106,N_9968,N_9835);
nand UO_107 (O_107,N_9892,N_9951);
and UO_108 (O_108,N_9927,N_9977);
nor UO_109 (O_109,N_9909,N_9869);
or UO_110 (O_110,N_9955,N_9896);
nand UO_111 (O_111,N_9867,N_9841);
or UO_112 (O_112,N_9974,N_9818);
or UO_113 (O_113,N_9821,N_9911);
nor UO_114 (O_114,N_9898,N_9939);
or UO_115 (O_115,N_9982,N_9822);
or UO_116 (O_116,N_9838,N_9807);
xnor UO_117 (O_117,N_9848,N_9875);
xor UO_118 (O_118,N_9857,N_9950);
nand UO_119 (O_119,N_9897,N_9869);
nor UO_120 (O_120,N_9898,N_9885);
and UO_121 (O_121,N_9870,N_9857);
nor UO_122 (O_122,N_9946,N_9977);
or UO_123 (O_123,N_9877,N_9804);
or UO_124 (O_124,N_9804,N_9998);
and UO_125 (O_125,N_9810,N_9970);
nor UO_126 (O_126,N_9839,N_9847);
nand UO_127 (O_127,N_9820,N_9933);
nor UO_128 (O_128,N_9996,N_9875);
and UO_129 (O_129,N_9820,N_9928);
and UO_130 (O_130,N_9938,N_9836);
and UO_131 (O_131,N_9821,N_9802);
xor UO_132 (O_132,N_9866,N_9985);
and UO_133 (O_133,N_9924,N_9857);
nor UO_134 (O_134,N_9801,N_9818);
or UO_135 (O_135,N_9861,N_9919);
or UO_136 (O_136,N_9834,N_9880);
nand UO_137 (O_137,N_9936,N_9894);
nand UO_138 (O_138,N_9959,N_9933);
or UO_139 (O_139,N_9982,N_9807);
nor UO_140 (O_140,N_9907,N_9971);
xor UO_141 (O_141,N_9958,N_9911);
nand UO_142 (O_142,N_9950,N_9829);
and UO_143 (O_143,N_9917,N_9913);
nor UO_144 (O_144,N_9800,N_9945);
or UO_145 (O_145,N_9823,N_9884);
nor UO_146 (O_146,N_9933,N_9815);
nand UO_147 (O_147,N_9846,N_9971);
and UO_148 (O_148,N_9866,N_9925);
nor UO_149 (O_149,N_9922,N_9888);
nor UO_150 (O_150,N_9973,N_9824);
and UO_151 (O_151,N_9928,N_9840);
nand UO_152 (O_152,N_9806,N_9851);
and UO_153 (O_153,N_9838,N_9883);
nor UO_154 (O_154,N_9875,N_9954);
or UO_155 (O_155,N_9851,N_9819);
nor UO_156 (O_156,N_9979,N_9993);
and UO_157 (O_157,N_9906,N_9945);
or UO_158 (O_158,N_9978,N_9857);
or UO_159 (O_159,N_9935,N_9932);
xnor UO_160 (O_160,N_9982,N_9910);
nor UO_161 (O_161,N_9995,N_9953);
and UO_162 (O_162,N_9900,N_9999);
and UO_163 (O_163,N_9848,N_9890);
nor UO_164 (O_164,N_9919,N_9854);
nor UO_165 (O_165,N_9940,N_9893);
nand UO_166 (O_166,N_9952,N_9858);
or UO_167 (O_167,N_9862,N_9928);
or UO_168 (O_168,N_9891,N_9981);
and UO_169 (O_169,N_9904,N_9991);
and UO_170 (O_170,N_9932,N_9808);
or UO_171 (O_171,N_9809,N_9986);
and UO_172 (O_172,N_9810,N_9901);
nor UO_173 (O_173,N_9899,N_9963);
and UO_174 (O_174,N_9847,N_9961);
nor UO_175 (O_175,N_9933,N_9984);
nand UO_176 (O_176,N_9899,N_9800);
xnor UO_177 (O_177,N_9886,N_9820);
xnor UO_178 (O_178,N_9921,N_9979);
and UO_179 (O_179,N_9990,N_9833);
nand UO_180 (O_180,N_9841,N_9809);
nor UO_181 (O_181,N_9887,N_9981);
and UO_182 (O_182,N_9978,N_9848);
xnor UO_183 (O_183,N_9964,N_9803);
or UO_184 (O_184,N_9894,N_9822);
xor UO_185 (O_185,N_9905,N_9961);
or UO_186 (O_186,N_9857,N_9952);
and UO_187 (O_187,N_9965,N_9844);
nor UO_188 (O_188,N_9956,N_9832);
nand UO_189 (O_189,N_9888,N_9840);
nor UO_190 (O_190,N_9891,N_9972);
and UO_191 (O_191,N_9807,N_9975);
nor UO_192 (O_192,N_9879,N_9940);
or UO_193 (O_193,N_9982,N_9978);
and UO_194 (O_194,N_9801,N_9828);
nand UO_195 (O_195,N_9857,N_9958);
nor UO_196 (O_196,N_9889,N_9806);
or UO_197 (O_197,N_9811,N_9972);
and UO_198 (O_198,N_9923,N_9844);
and UO_199 (O_199,N_9857,N_9966);
nand UO_200 (O_200,N_9826,N_9844);
and UO_201 (O_201,N_9866,N_9821);
nand UO_202 (O_202,N_9832,N_9914);
nand UO_203 (O_203,N_9843,N_9847);
or UO_204 (O_204,N_9870,N_9830);
nor UO_205 (O_205,N_9972,N_9963);
and UO_206 (O_206,N_9801,N_9977);
or UO_207 (O_207,N_9927,N_9938);
or UO_208 (O_208,N_9939,N_9906);
and UO_209 (O_209,N_9939,N_9862);
nor UO_210 (O_210,N_9975,N_9833);
nor UO_211 (O_211,N_9831,N_9982);
or UO_212 (O_212,N_9875,N_9924);
nor UO_213 (O_213,N_9830,N_9993);
nand UO_214 (O_214,N_9868,N_9823);
nor UO_215 (O_215,N_9825,N_9888);
and UO_216 (O_216,N_9885,N_9802);
nor UO_217 (O_217,N_9946,N_9838);
and UO_218 (O_218,N_9852,N_9814);
and UO_219 (O_219,N_9991,N_9902);
or UO_220 (O_220,N_9849,N_9831);
nor UO_221 (O_221,N_9908,N_9867);
nor UO_222 (O_222,N_9840,N_9837);
nor UO_223 (O_223,N_9828,N_9940);
nand UO_224 (O_224,N_9859,N_9813);
and UO_225 (O_225,N_9819,N_9849);
or UO_226 (O_226,N_9857,N_9842);
nor UO_227 (O_227,N_9988,N_9902);
nand UO_228 (O_228,N_9863,N_9947);
and UO_229 (O_229,N_9801,N_9846);
nand UO_230 (O_230,N_9830,N_9984);
nor UO_231 (O_231,N_9936,N_9848);
nand UO_232 (O_232,N_9993,N_9933);
nand UO_233 (O_233,N_9968,N_9970);
nand UO_234 (O_234,N_9874,N_9918);
nor UO_235 (O_235,N_9916,N_9982);
nor UO_236 (O_236,N_9893,N_9828);
and UO_237 (O_237,N_9801,N_9946);
nand UO_238 (O_238,N_9932,N_9812);
or UO_239 (O_239,N_9829,N_9983);
or UO_240 (O_240,N_9852,N_9900);
or UO_241 (O_241,N_9871,N_9996);
nor UO_242 (O_242,N_9846,N_9828);
nor UO_243 (O_243,N_9895,N_9808);
and UO_244 (O_244,N_9825,N_9931);
nor UO_245 (O_245,N_9940,N_9862);
nand UO_246 (O_246,N_9853,N_9959);
or UO_247 (O_247,N_9997,N_9940);
or UO_248 (O_248,N_9966,N_9871);
nor UO_249 (O_249,N_9911,N_9918);
nor UO_250 (O_250,N_9987,N_9949);
or UO_251 (O_251,N_9877,N_9858);
nor UO_252 (O_252,N_9823,N_9924);
xnor UO_253 (O_253,N_9806,N_9913);
nor UO_254 (O_254,N_9829,N_9923);
or UO_255 (O_255,N_9971,N_9989);
nand UO_256 (O_256,N_9908,N_9897);
nor UO_257 (O_257,N_9970,N_9975);
nand UO_258 (O_258,N_9825,N_9848);
and UO_259 (O_259,N_9906,N_9971);
nand UO_260 (O_260,N_9825,N_9869);
and UO_261 (O_261,N_9933,N_9917);
xor UO_262 (O_262,N_9880,N_9879);
and UO_263 (O_263,N_9865,N_9862);
or UO_264 (O_264,N_9959,N_9911);
nor UO_265 (O_265,N_9950,N_9888);
and UO_266 (O_266,N_9856,N_9831);
xnor UO_267 (O_267,N_9951,N_9845);
nand UO_268 (O_268,N_9911,N_9972);
nand UO_269 (O_269,N_9831,N_9931);
or UO_270 (O_270,N_9853,N_9837);
and UO_271 (O_271,N_9882,N_9871);
or UO_272 (O_272,N_9921,N_9873);
xnor UO_273 (O_273,N_9819,N_9972);
and UO_274 (O_274,N_9985,N_9898);
xor UO_275 (O_275,N_9838,N_9869);
nor UO_276 (O_276,N_9992,N_9973);
nand UO_277 (O_277,N_9912,N_9941);
nand UO_278 (O_278,N_9979,N_9813);
or UO_279 (O_279,N_9965,N_9868);
or UO_280 (O_280,N_9975,N_9834);
or UO_281 (O_281,N_9943,N_9957);
nand UO_282 (O_282,N_9859,N_9884);
or UO_283 (O_283,N_9843,N_9882);
and UO_284 (O_284,N_9820,N_9881);
nand UO_285 (O_285,N_9965,N_9940);
and UO_286 (O_286,N_9870,N_9869);
or UO_287 (O_287,N_9843,N_9969);
nand UO_288 (O_288,N_9887,N_9879);
nand UO_289 (O_289,N_9953,N_9852);
nor UO_290 (O_290,N_9871,N_9979);
nor UO_291 (O_291,N_9884,N_9941);
and UO_292 (O_292,N_9959,N_9863);
nor UO_293 (O_293,N_9937,N_9832);
xor UO_294 (O_294,N_9845,N_9984);
xnor UO_295 (O_295,N_9852,N_9872);
and UO_296 (O_296,N_9844,N_9833);
and UO_297 (O_297,N_9816,N_9823);
and UO_298 (O_298,N_9809,N_9886);
and UO_299 (O_299,N_9898,N_9924);
or UO_300 (O_300,N_9901,N_9949);
and UO_301 (O_301,N_9890,N_9813);
nor UO_302 (O_302,N_9963,N_9924);
nand UO_303 (O_303,N_9811,N_9921);
or UO_304 (O_304,N_9892,N_9834);
and UO_305 (O_305,N_9970,N_9990);
nand UO_306 (O_306,N_9926,N_9892);
and UO_307 (O_307,N_9833,N_9999);
xnor UO_308 (O_308,N_9914,N_9859);
xor UO_309 (O_309,N_9941,N_9949);
nand UO_310 (O_310,N_9902,N_9896);
nand UO_311 (O_311,N_9987,N_9836);
nand UO_312 (O_312,N_9808,N_9930);
nor UO_313 (O_313,N_9812,N_9996);
nor UO_314 (O_314,N_9973,N_9979);
nor UO_315 (O_315,N_9965,N_9831);
nand UO_316 (O_316,N_9910,N_9879);
nand UO_317 (O_317,N_9851,N_9811);
nand UO_318 (O_318,N_9834,N_9993);
nand UO_319 (O_319,N_9945,N_9996);
and UO_320 (O_320,N_9805,N_9835);
nand UO_321 (O_321,N_9928,N_9958);
or UO_322 (O_322,N_9850,N_9930);
xnor UO_323 (O_323,N_9909,N_9868);
nor UO_324 (O_324,N_9959,N_9879);
nor UO_325 (O_325,N_9960,N_9944);
nand UO_326 (O_326,N_9986,N_9810);
and UO_327 (O_327,N_9853,N_9878);
nand UO_328 (O_328,N_9825,N_9917);
and UO_329 (O_329,N_9918,N_9851);
xnor UO_330 (O_330,N_9881,N_9863);
and UO_331 (O_331,N_9940,N_9967);
or UO_332 (O_332,N_9947,N_9906);
nand UO_333 (O_333,N_9862,N_9898);
or UO_334 (O_334,N_9909,N_9967);
nor UO_335 (O_335,N_9936,N_9974);
nor UO_336 (O_336,N_9979,N_9959);
and UO_337 (O_337,N_9950,N_9803);
xnor UO_338 (O_338,N_9817,N_9991);
and UO_339 (O_339,N_9926,N_9994);
or UO_340 (O_340,N_9965,N_9827);
or UO_341 (O_341,N_9886,N_9854);
nor UO_342 (O_342,N_9995,N_9916);
or UO_343 (O_343,N_9902,N_9875);
nand UO_344 (O_344,N_9824,N_9854);
nor UO_345 (O_345,N_9956,N_9997);
and UO_346 (O_346,N_9961,N_9924);
and UO_347 (O_347,N_9823,N_9812);
nand UO_348 (O_348,N_9892,N_9996);
nand UO_349 (O_349,N_9990,N_9815);
xnor UO_350 (O_350,N_9897,N_9927);
or UO_351 (O_351,N_9864,N_9938);
nand UO_352 (O_352,N_9944,N_9821);
and UO_353 (O_353,N_9935,N_9955);
or UO_354 (O_354,N_9825,N_9854);
nor UO_355 (O_355,N_9927,N_9933);
nor UO_356 (O_356,N_9814,N_9840);
nand UO_357 (O_357,N_9836,N_9831);
nand UO_358 (O_358,N_9804,N_9935);
nand UO_359 (O_359,N_9900,N_9953);
and UO_360 (O_360,N_9961,N_9839);
nand UO_361 (O_361,N_9947,N_9872);
nor UO_362 (O_362,N_9876,N_9958);
or UO_363 (O_363,N_9904,N_9891);
xnor UO_364 (O_364,N_9920,N_9910);
or UO_365 (O_365,N_9980,N_9887);
and UO_366 (O_366,N_9902,N_9847);
nand UO_367 (O_367,N_9801,N_9992);
nand UO_368 (O_368,N_9931,N_9905);
nand UO_369 (O_369,N_9991,N_9837);
nor UO_370 (O_370,N_9816,N_9914);
and UO_371 (O_371,N_9815,N_9922);
nor UO_372 (O_372,N_9802,N_9824);
nand UO_373 (O_373,N_9890,N_9888);
nor UO_374 (O_374,N_9867,N_9991);
nor UO_375 (O_375,N_9857,N_9932);
and UO_376 (O_376,N_9985,N_9973);
or UO_377 (O_377,N_9947,N_9877);
nor UO_378 (O_378,N_9916,N_9976);
nand UO_379 (O_379,N_9977,N_9873);
nand UO_380 (O_380,N_9936,N_9939);
or UO_381 (O_381,N_9838,N_9876);
nand UO_382 (O_382,N_9838,N_9977);
or UO_383 (O_383,N_9935,N_9948);
nand UO_384 (O_384,N_9915,N_9981);
or UO_385 (O_385,N_9975,N_9813);
and UO_386 (O_386,N_9806,N_9825);
and UO_387 (O_387,N_9915,N_9909);
or UO_388 (O_388,N_9817,N_9885);
and UO_389 (O_389,N_9993,N_9803);
nor UO_390 (O_390,N_9853,N_9834);
or UO_391 (O_391,N_9872,N_9975);
and UO_392 (O_392,N_9933,N_9822);
xor UO_393 (O_393,N_9816,N_9984);
nor UO_394 (O_394,N_9955,N_9910);
or UO_395 (O_395,N_9908,N_9928);
or UO_396 (O_396,N_9841,N_9999);
or UO_397 (O_397,N_9906,N_9864);
and UO_398 (O_398,N_9916,N_9883);
nor UO_399 (O_399,N_9908,N_9807);
nor UO_400 (O_400,N_9830,N_9962);
or UO_401 (O_401,N_9975,N_9880);
or UO_402 (O_402,N_9838,N_9998);
or UO_403 (O_403,N_9852,N_9882);
nor UO_404 (O_404,N_9949,N_9968);
or UO_405 (O_405,N_9935,N_9848);
xnor UO_406 (O_406,N_9846,N_9867);
xnor UO_407 (O_407,N_9819,N_9935);
nor UO_408 (O_408,N_9907,N_9898);
nand UO_409 (O_409,N_9983,N_9806);
nand UO_410 (O_410,N_9814,N_9944);
and UO_411 (O_411,N_9878,N_9894);
and UO_412 (O_412,N_9964,N_9924);
nand UO_413 (O_413,N_9965,N_9987);
nor UO_414 (O_414,N_9819,N_9820);
and UO_415 (O_415,N_9953,N_9917);
nand UO_416 (O_416,N_9939,N_9970);
and UO_417 (O_417,N_9937,N_9802);
and UO_418 (O_418,N_9836,N_9843);
or UO_419 (O_419,N_9897,N_9809);
or UO_420 (O_420,N_9959,N_9935);
and UO_421 (O_421,N_9911,N_9898);
nand UO_422 (O_422,N_9916,N_9892);
nand UO_423 (O_423,N_9972,N_9998);
and UO_424 (O_424,N_9949,N_9976);
or UO_425 (O_425,N_9884,N_9852);
nand UO_426 (O_426,N_9946,N_9897);
nand UO_427 (O_427,N_9924,N_9955);
and UO_428 (O_428,N_9951,N_9950);
or UO_429 (O_429,N_9974,N_9866);
nand UO_430 (O_430,N_9838,N_9979);
nand UO_431 (O_431,N_9930,N_9948);
nor UO_432 (O_432,N_9805,N_9897);
or UO_433 (O_433,N_9988,N_9987);
and UO_434 (O_434,N_9862,N_9986);
and UO_435 (O_435,N_9886,N_9966);
xor UO_436 (O_436,N_9848,N_9919);
nand UO_437 (O_437,N_9903,N_9805);
nor UO_438 (O_438,N_9908,N_9804);
or UO_439 (O_439,N_9824,N_9810);
nand UO_440 (O_440,N_9981,N_9802);
or UO_441 (O_441,N_9918,N_9809);
and UO_442 (O_442,N_9958,N_9952);
or UO_443 (O_443,N_9956,N_9931);
xnor UO_444 (O_444,N_9916,N_9829);
or UO_445 (O_445,N_9800,N_9903);
xor UO_446 (O_446,N_9901,N_9970);
and UO_447 (O_447,N_9840,N_9810);
or UO_448 (O_448,N_9965,N_9845);
nor UO_449 (O_449,N_9983,N_9937);
nor UO_450 (O_450,N_9984,N_9839);
or UO_451 (O_451,N_9920,N_9996);
and UO_452 (O_452,N_9850,N_9863);
and UO_453 (O_453,N_9838,N_9820);
or UO_454 (O_454,N_9850,N_9900);
and UO_455 (O_455,N_9911,N_9982);
or UO_456 (O_456,N_9937,N_9948);
nand UO_457 (O_457,N_9923,N_9876);
or UO_458 (O_458,N_9951,N_9972);
nor UO_459 (O_459,N_9887,N_9919);
nor UO_460 (O_460,N_9825,N_9853);
nand UO_461 (O_461,N_9950,N_9868);
or UO_462 (O_462,N_9957,N_9835);
and UO_463 (O_463,N_9855,N_9810);
and UO_464 (O_464,N_9825,N_9903);
nor UO_465 (O_465,N_9847,N_9959);
and UO_466 (O_466,N_9966,N_9888);
xnor UO_467 (O_467,N_9976,N_9814);
nor UO_468 (O_468,N_9842,N_9884);
nor UO_469 (O_469,N_9838,N_9804);
nor UO_470 (O_470,N_9826,N_9922);
nand UO_471 (O_471,N_9896,N_9855);
nand UO_472 (O_472,N_9849,N_9881);
or UO_473 (O_473,N_9811,N_9960);
or UO_474 (O_474,N_9946,N_9857);
nand UO_475 (O_475,N_9871,N_9895);
nor UO_476 (O_476,N_9895,N_9807);
and UO_477 (O_477,N_9865,N_9859);
or UO_478 (O_478,N_9952,N_9870);
and UO_479 (O_479,N_9910,N_9820);
xor UO_480 (O_480,N_9840,N_9894);
and UO_481 (O_481,N_9861,N_9804);
xor UO_482 (O_482,N_9841,N_9934);
nand UO_483 (O_483,N_9858,N_9834);
and UO_484 (O_484,N_9933,N_9910);
nand UO_485 (O_485,N_9831,N_9903);
nor UO_486 (O_486,N_9807,N_9887);
xnor UO_487 (O_487,N_9992,N_9825);
nand UO_488 (O_488,N_9900,N_9968);
nor UO_489 (O_489,N_9816,N_9869);
or UO_490 (O_490,N_9861,N_9996);
nand UO_491 (O_491,N_9843,N_9855);
and UO_492 (O_492,N_9892,N_9859);
and UO_493 (O_493,N_9835,N_9931);
or UO_494 (O_494,N_9834,N_9910);
or UO_495 (O_495,N_9992,N_9970);
nand UO_496 (O_496,N_9945,N_9986);
nand UO_497 (O_497,N_9826,N_9903);
nor UO_498 (O_498,N_9836,N_9978);
nand UO_499 (O_499,N_9944,N_9817);
nand UO_500 (O_500,N_9834,N_9898);
nand UO_501 (O_501,N_9989,N_9918);
nand UO_502 (O_502,N_9811,N_9809);
or UO_503 (O_503,N_9846,N_9966);
or UO_504 (O_504,N_9803,N_9938);
nand UO_505 (O_505,N_9815,N_9812);
and UO_506 (O_506,N_9972,N_9828);
or UO_507 (O_507,N_9855,N_9914);
nand UO_508 (O_508,N_9962,N_9879);
or UO_509 (O_509,N_9903,N_9883);
nand UO_510 (O_510,N_9846,N_9885);
or UO_511 (O_511,N_9949,N_9912);
nor UO_512 (O_512,N_9907,N_9811);
nand UO_513 (O_513,N_9927,N_9997);
nand UO_514 (O_514,N_9804,N_9966);
nand UO_515 (O_515,N_9983,N_9816);
nand UO_516 (O_516,N_9901,N_9903);
or UO_517 (O_517,N_9983,N_9935);
and UO_518 (O_518,N_9825,N_9837);
nand UO_519 (O_519,N_9944,N_9908);
and UO_520 (O_520,N_9903,N_9809);
nor UO_521 (O_521,N_9958,N_9951);
xor UO_522 (O_522,N_9930,N_9936);
or UO_523 (O_523,N_9981,N_9959);
nand UO_524 (O_524,N_9832,N_9801);
xor UO_525 (O_525,N_9908,N_9801);
nand UO_526 (O_526,N_9923,N_9835);
and UO_527 (O_527,N_9902,N_9936);
or UO_528 (O_528,N_9945,N_9894);
nand UO_529 (O_529,N_9847,N_9903);
xor UO_530 (O_530,N_9846,N_9878);
nor UO_531 (O_531,N_9965,N_9915);
nand UO_532 (O_532,N_9887,N_9830);
and UO_533 (O_533,N_9999,N_9993);
nand UO_534 (O_534,N_9904,N_9873);
nand UO_535 (O_535,N_9948,N_9838);
or UO_536 (O_536,N_9830,N_9915);
and UO_537 (O_537,N_9930,N_9912);
nand UO_538 (O_538,N_9953,N_9978);
and UO_539 (O_539,N_9841,N_9891);
nor UO_540 (O_540,N_9843,N_9941);
nand UO_541 (O_541,N_9900,N_9992);
or UO_542 (O_542,N_9936,N_9821);
nor UO_543 (O_543,N_9914,N_9892);
nand UO_544 (O_544,N_9859,N_9880);
nor UO_545 (O_545,N_9805,N_9992);
nand UO_546 (O_546,N_9910,N_9861);
nor UO_547 (O_547,N_9847,N_9888);
nand UO_548 (O_548,N_9835,N_9838);
nand UO_549 (O_549,N_9951,N_9986);
and UO_550 (O_550,N_9818,N_9874);
or UO_551 (O_551,N_9916,N_9876);
nand UO_552 (O_552,N_9878,N_9813);
nor UO_553 (O_553,N_9929,N_9907);
nand UO_554 (O_554,N_9862,N_9951);
or UO_555 (O_555,N_9888,N_9864);
xor UO_556 (O_556,N_9940,N_9873);
nand UO_557 (O_557,N_9861,N_9800);
nor UO_558 (O_558,N_9837,N_9907);
nand UO_559 (O_559,N_9850,N_9842);
nor UO_560 (O_560,N_9901,N_9867);
and UO_561 (O_561,N_9957,N_9951);
or UO_562 (O_562,N_9937,N_9843);
xnor UO_563 (O_563,N_9895,N_9867);
nand UO_564 (O_564,N_9983,N_9909);
and UO_565 (O_565,N_9979,N_9995);
nor UO_566 (O_566,N_9808,N_9852);
and UO_567 (O_567,N_9941,N_9924);
nor UO_568 (O_568,N_9926,N_9861);
and UO_569 (O_569,N_9827,N_9807);
and UO_570 (O_570,N_9903,N_9807);
nand UO_571 (O_571,N_9899,N_9922);
nand UO_572 (O_572,N_9839,N_9952);
nor UO_573 (O_573,N_9980,N_9849);
nor UO_574 (O_574,N_9960,N_9888);
and UO_575 (O_575,N_9805,N_9918);
nand UO_576 (O_576,N_9855,N_9819);
or UO_577 (O_577,N_9863,N_9901);
or UO_578 (O_578,N_9822,N_9855);
and UO_579 (O_579,N_9980,N_9870);
nor UO_580 (O_580,N_9857,N_9827);
nor UO_581 (O_581,N_9883,N_9951);
nand UO_582 (O_582,N_9910,N_9929);
xnor UO_583 (O_583,N_9922,N_9970);
xor UO_584 (O_584,N_9976,N_9802);
and UO_585 (O_585,N_9995,N_9913);
nor UO_586 (O_586,N_9899,N_9928);
nor UO_587 (O_587,N_9878,N_9953);
xor UO_588 (O_588,N_9951,N_9832);
nor UO_589 (O_589,N_9910,N_9887);
and UO_590 (O_590,N_9861,N_9859);
and UO_591 (O_591,N_9878,N_9949);
nand UO_592 (O_592,N_9919,N_9807);
or UO_593 (O_593,N_9837,N_9988);
nand UO_594 (O_594,N_9884,N_9962);
and UO_595 (O_595,N_9976,N_9963);
or UO_596 (O_596,N_9880,N_9862);
nor UO_597 (O_597,N_9831,N_9829);
or UO_598 (O_598,N_9978,N_9809);
and UO_599 (O_599,N_9900,N_9978);
nor UO_600 (O_600,N_9950,N_9958);
nor UO_601 (O_601,N_9980,N_9932);
or UO_602 (O_602,N_9989,N_9997);
or UO_603 (O_603,N_9861,N_9824);
or UO_604 (O_604,N_9862,N_9925);
nand UO_605 (O_605,N_9926,N_9987);
nor UO_606 (O_606,N_9993,N_9850);
or UO_607 (O_607,N_9825,N_9880);
nand UO_608 (O_608,N_9944,N_9898);
or UO_609 (O_609,N_9860,N_9909);
nand UO_610 (O_610,N_9938,N_9952);
nor UO_611 (O_611,N_9985,N_9937);
or UO_612 (O_612,N_9949,N_9837);
or UO_613 (O_613,N_9920,N_9808);
xor UO_614 (O_614,N_9990,N_9961);
nand UO_615 (O_615,N_9868,N_9808);
nor UO_616 (O_616,N_9905,N_9807);
xor UO_617 (O_617,N_9834,N_9925);
nor UO_618 (O_618,N_9810,N_9862);
nand UO_619 (O_619,N_9871,N_9947);
and UO_620 (O_620,N_9987,N_9964);
nand UO_621 (O_621,N_9820,N_9899);
and UO_622 (O_622,N_9814,N_9819);
nor UO_623 (O_623,N_9891,N_9900);
and UO_624 (O_624,N_9837,N_9833);
and UO_625 (O_625,N_9987,N_9982);
nand UO_626 (O_626,N_9978,N_9801);
and UO_627 (O_627,N_9879,N_9986);
nand UO_628 (O_628,N_9830,N_9847);
nor UO_629 (O_629,N_9815,N_9952);
nand UO_630 (O_630,N_9910,N_9980);
nand UO_631 (O_631,N_9984,N_9979);
nor UO_632 (O_632,N_9927,N_9958);
and UO_633 (O_633,N_9925,N_9878);
xor UO_634 (O_634,N_9892,N_9888);
nor UO_635 (O_635,N_9938,N_9868);
and UO_636 (O_636,N_9991,N_9811);
nand UO_637 (O_637,N_9926,N_9853);
nor UO_638 (O_638,N_9923,N_9974);
or UO_639 (O_639,N_9898,N_9903);
nand UO_640 (O_640,N_9848,N_9929);
nand UO_641 (O_641,N_9947,N_9858);
or UO_642 (O_642,N_9886,N_9920);
nor UO_643 (O_643,N_9863,N_9867);
nor UO_644 (O_644,N_9848,N_9996);
and UO_645 (O_645,N_9836,N_9844);
or UO_646 (O_646,N_9924,N_9984);
nand UO_647 (O_647,N_9938,N_9930);
or UO_648 (O_648,N_9960,N_9954);
nor UO_649 (O_649,N_9806,N_9839);
nand UO_650 (O_650,N_9888,N_9934);
or UO_651 (O_651,N_9846,N_9904);
nand UO_652 (O_652,N_9986,N_9821);
and UO_653 (O_653,N_9836,N_9828);
nor UO_654 (O_654,N_9980,N_9842);
nor UO_655 (O_655,N_9956,N_9815);
nor UO_656 (O_656,N_9815,N_9809);
nor UO_657 (O_657,N_9884,N_9803);
or UO_658 (O_658,N_9986,N_9929);
or UO_659 (O_659,N_9836,N_9939);
nor UO_660 (O_660,N_9989,N_9942);
and UO_661 (O_661,N_9857,N_9840);
nor UO_662 (O_662,N_9908,N_9803);
nand UO_663 (O_663,N_9851,N_9814);
xor UO_664 (O_664,N_9825,N_9863);
xnor UO_665 (O_665,N_9999,N_9921);
nand UO_666 (O_666,N_9840,N_9991);
nor UO_667 (O_667,N_9986,N_9863);
nand UO_668 (O_668,N_9964,N_9942);
nor UO_669 (O_669,N_9822,N_9942);
nor UO_670 (O_670,N_9839,N_9857);
or UO_671 (O_671,N_9802,N_9944);
nand UO_672 (O_672,N_9951,N_9997);
or UO_673 (O_673,N_9848,N_9823);
nor UO_674 (O_674,N_9838,N_9999);
and UO_675 (O_675,N_9815,N_9870);
nand UO_676 (O_676,N_9853,N_9972);
and UO_677 (O_677,N_9862,N_9845);
and UO_678 (O_678,N_9985,N_9961);
or UO_679 (O_679,N_9892,N_9864);
or UO_680 (O_680,N_9846,N_9964);
and UO_681 (O_681,N_9915,N_9976);
or UO_682 (O_682,N_9810,N_9819);
nand UO_683 (O_683,N_9986,N_9878);
nor UO_684 (O_684,N_9927,N_9976);
nand UO_685 (O_685,N_9984,N_9958);
nand UO_686 (O_686,N_9875,N_9880);
and UO_687 (O_687,N_9802,N_9960);
or UO_688 (O_688,N_9903,N_9992);
or UO_689 (O_689,N_9881,N_9932);
nor UO_690 (O_690,N_9841,N_9958);
or UO_691 (O_691,N_9916,N_9811);
nor UO_692 (O_692,N_9891,N_9896);
and UO_693 (O_693,N_9914,N_9807);
nand UO_694 (O_694,N_9866,N_9861);
nor UO_695 (O_695,N_9967,N_9861);
and UO_696 (O_696,N_9812,N_9971);
or UO_697 (O_697,N_9921,N_9944);
and UO_698 (O_698,N_9974,N_9932);
nand UO_699 (O_699,N_9902,N_9877);
or UO_700 (O_700,N_9950,N_9804);
nor UO_701 (O_701,N_9900,N_9859);
nor UO_702 (O_702,N_9823,N_9854);
xor UO_703 (O_703,N_9909,N_9947);
or UO_704 (O_704,N_9979,N_9961);
nor UO_705 (O_705,N_9936,N_9949);
nor UO_706 (O_706,N_9927,N_9811);
and UO_707 (O_707,N_9893,N_9888);
nor UO_708 (O_708,N_9856,N_9913);
and UO_709 (O_709,N_9853,N_9913);
and UO_710 (O_710,N_9800,N_9915);
nor UO_711 (O_711,N_9989,N_9808);
nor UO_712 (O_712,N_9959,N_9857);
nor UO_713 (O_713,N_9871,N_9962);
and UO_714 (O_714,N_9907,N_9965);
nor UO_715 (O_715,N_9914,N_9881);
and UO_716 (O_716,N_9857,N_9929);
nand UO_717 (O_717,N_9941,N_9940);
xor UO_718 (O_718,N_9986,N_9856);
and UO_719 (O_719,N_9888,N_9932);
and UO_720 (O_720,N_9856,N_9802);
xnor UO_721 (O_721,N_9956,N_9835);
nand UO_722 (O_722,N_9874,N_9855);
and UO_723 (O_723,N_9925,N_9845);
or UO_724 (O_724,N_9851,N_9997);
and UO_725 (O_725,N_9996,N_9894);
xor UO_726 (O_726,N_9868,N_9863);
xor UO_727 (O_727,N_9804,N_9812);
and UO_728 (O_728,N_9854,N_9800);
nor UO_729 (O_729,N_9954,N_9986);
nor UO_730 (O_730,N_9829,N_9873);
and UO_731 (O_731,N_9889,N_9955);
or UO_732 (O_732,N_9957,N_9815);
nor UO_733 (O_733,N_9900,N_9895);
and UO_734 (O_734,N_9936,N_9911);
and UO_735 (O_735,N_9873,N_9998);
nand UO_736 (O_736,N_9959,N_9997);
xor UO_737 (O_737,N_9914,N_9882);
nor UO_738 (O_738,N_9841,N_9938);
nor UO_739 (O_739,N_9909,N_9849);
xor UO_740 (O_740,N_9927,N_9982);
or UO_741 (O_741,N_9881,N_9864);
and UO_742 (O_742,N_9824,N_9939);
nand UO_743 (O_743,N_9956,N_9971);
or UO_744 (O_744,N_9938,N_9872);
or UO_745 (O_745,N_9844,N_9898);
or UO_746 (O_746,N_9855,N_9923);
and UO_747 (O_747,N_9988,N_9907);
nand UO_748 (O_748,N_9866,N_9804);
nor UO_749 (O_749,N_9917,N_9853);
xnor UO_750 (O_750,N_9894,N_9898);
and UO_751 (O_751,N_9906,N_9838);
nand UO_752 (O_752,N_9946,N_9829);
nor UO_753 (O_753,N_9947,N_9923);
nor UO_754 (O_754,N_9998,N_9929);
and UO_755 (O_755,N_9865,N_9849);
nand UO_756 (O_756,N_9851,N_9869);
nor UO_757 (O_757,N_9943,N_9936);
and UO_758 (O_758,N_9828,N_9934);
xnor UO_759 (O_759,N_9819,N_9962);
and UO_760 (O_760,N_9953,N_9948);
nor UO_761 (O_761,N_9957,N_9959);
and UO_762 (O_762,N_9839,N_9894);
nand UO_763 (O_763,N_9868,N_9934);
nor UO_764 (O_764,N_9966,N_9960);
nor UO_765 (O_765,N_9870,N_9909);
nor UO_766 (O_766,N_9920,N_9856);
or UO_767 (O_767,N_9828,N_9903);
or UO_768 (O_768,N_9995,N_9894);
and UO_769 (O_769,N_9875,N_9988);
and UO_770 (O_770,N_9886,N_9846);
nand UO_771 (O_771,N_9936,N_9982);
nor UO_772 (O_772,N_9951,N_9856);
nand UO_773 (O_773,N_9993,N_9880);
or UO_774 (O_774,N_9998,N_9808);
and UO_775 (O_775,N_9850,N_9875);
xor UO_776 (O_776,N_9978,N_9875);
nor UO_777 (O_777,N_9854,N_9994);
or UO_778 (O_778,N_9924,N_9983);
nor UO_779 (O_779,N_9841,N_9835);
or UO_780 (O_780,N_9815,N_9831);
nor UO_781 (O_781,N_9838,N_9910);
nor UO_782 (O_782,N_9976,N_9996);
xnor UO_783 (O_783,N_9873,N_9897);
or UO_784 (O_784,N_9984,N_9896);
nor UO_785 (O_785,N_9866,N_9971);
nand UO_786 (O_786,N_9897,N_9953);
nor UO_787 (O_787,N_9987,N_9829);
nand UO_788 (O_788,N_9906,N_9887);
nand UO_789 (O_789,N_9811,N_9887);
nand UO_790 (O_790,N_9929,N_9811);
or UO_791 (O_791,N_9932,N_9900);
nor UO_792 (O_792,N_9867,N_9853);
nand UO_793 (O_793,N_9839,N_9981);
and UO_794 (O_794,N_9996,N_9992);
xor UO_795 (O_795,N_9980,N_9934);
and UO_796 (O_796,N_9996,N_9828);
nor UO_797 (O_797,N_9929,N_9802);
and UO_798 (O_798,N_9861,N_9849);
or UO_799 (O_799,N_9886,N_9890);
or UO_800 (O_800,N_9814,N_9859);
nor UO_801 (O_801,N_9848,N_9854);
xnor UO_802 (O_802,N_9846,N_9880);
nand UO_803 (O_803,N_9890,N_9983);
xor UO_804 (O_804,N_9818,N_9993);
nand UO_805 (O_805,N_9972,N_9833);
and UO_806 (O_806,N_9897,N_9997);
nand UO_807 (O_807,N_9985,N_9843);
xor UO_808 (O_808,N_9952,N_9978);
nor UO_809 (O_809,N_9863,N_9968);
nor UO_810 (O_810,N_9933,N_9884);
nand UO_811 (O_811,N_9925,N_9979);
or UO_812 (O_812,N_9839,N_9867);
nand UO_813 (O_813,N_9893,N_9981);
or UO_814 (O_814,N_9870,N_9864);
or UO_815 (O_815,N_9906,N_9854);
nor UO_816 (O_816,N_9826,N_9825);
and UO_817 (O_817,N_9895,N_9868);
xor UO_818 (O_818,N_9876,N_9998);
xnor UO_819 (O_819,N_9893,N_9907);
or UO_820 (O_820,N_9878,N_9921);
and UO_821 (O_821,N_9878,N_9899);
nand UO_822 (O_822,N_9893,N_9931);
nor UO_823 (O_823,N_9926,N_9942);
or UO_824 (O_824,N_9898,N_9968);
nand UO_825 (O_825,N_9956,N_9801);
or UO_826 (O_826,N_9879,N_9979);
nor UO_827 (O_827,N_9893,N_9844);
and UO_828 (O_828,N_9826,N_9864);
nand UO_829 (O_829,N_9839,N_9936);
nand UO_830 (O_830,N_9937,N_9863);
xnor UO_831 (O_831,N_9857,N_9818);
or UO_832 (O_832,N_9818,N_9959);
xor UO_833 (O_833,N_9822,N_9971);
nand UO_834 (O_834,N_9804,N_9928);
and UO_835 (O_835,N_9867,N_9923);
and UO_836 (O_836,N_9917,N_9821);
and UO_837 (O_837,N_9837,N_9836);
nand UO_838 (O_838,N_9892,N_9967);
xnor UO_839 (O_839,N_9856,N_9849);
or UO_840 (O_840,N_9977,N_9853);
and UO_841 (O_841,N_9884,N_9892);
nor UO_842 (O_842,N_9894,N_9830);
nor UO_843 (O_843,N_9878,N_9932);
nand UO_844 (O_844,N_9922,N_9969);
nor UO_845 (O_845,N_9872,N_9817);
nand UO_846 (O_846,N_9947,N_9910);
nand UO_847 (O_847,N_9810,N_9998);
nor UO_848 (O_848,N_9914,N_9858);
nand UO_849 (O_849,N_9848,N_9956);
or UO_850 (O_850,N_9830,N_9854);
and UO_851 (O_851,N_9926,N_9842);
nor UO_852 (O_852,N_9901,N_9853);
nor UO_853 (O_853,N_9811,N_9816);
and UO_854 (O_854,N_9830,N_9855);
or UO_855 (O_855,N_9876,N_9852);
and UO_856 (O_856,N_9809,N_9860);
and UO_857 (O_857,N_9876,N_9975);
nor UO_858 (O_858,N_9958,N_9811);
and UO_859 (O_859,N_9961,N_9948);
and UO_860 (O_860,N_9955,N_9938);
nand UO_861 (O_861,N_9915,N_9952);
and UO_862 (O_862,N_9930,N_9842);
xor UO_863 (O_863,N_9913,N_9889);
nand UO_864 (O_864,N_9855,N_9827);
nor UO_865 (O_865,N_9865,N_9959);
nor UO_866 (O_866,N_9999,N_9817);
or UO_867 (O_867,N_9987,N_9938);
nor UO_868 (O_868,N_9943,N_9884);
and UO_869 (O_869,N_9973,N_9942);
or UO_870 (O_870,N_9996,N_9826);
nor UO_871 (O_871,N_9836,N_9991);
nand UO_872 (O_872,N_9816,N_9968);
nand UO_873 (O_873,N_9854,N_9968);
and UO_874 (O_874,N_9839,N_9912);
nor UO_875 (O_875,N_9819,N_9884);
xor UO_876 (O_876,N_9822,N_9873);
nand UO_877 (O_877,N_9913,N_9934);
nor UO_878 (O_878,N_9811,N_9812);
and UO_879 (O_879,N_9878,N_9826);
or UO_880 (O_880,N_9905,N_9947);
nand UO_881 (O_881,N_9937,N_9867);
nor UO_882 (O_882,N_9990,N_9820);
nor UO_883 (O_883,N_9888,N_9873);
nand UO_884 (O_884,N_9820,N_9901);
and UO_885 (O_885,N_9805,N_9868);
nor UO_886 (O_886,N_9992,N_9901);
and UO_887 (O_887,N_9935,N_9911);
nand UO_888 (O_888,N_9989,N_9864);
nor UO_889 (O_889,N_9896,N_9924);
nand UO_890 (O_890,N_9806,N_9926);
xnor UO_891 (O_891,N_9872,N_9869);
nor UO_892 (O_892,N_9976,N_9979);
nor UO_893 (O_893,N_9969,N_9837);
or UO_894 (O_894,N_9838,N_9834);
or UO_895 (O_895,N_9861,N_9840);
and UO_896 (O_896,N_9813,N_9985);
or UO_897 (O_897,N_9983,N_9999);
nand UO_898 (O_898,N_9911,N_9854);
nor UO_899 (O_899,N_9969,N_9920);
xnor UO_900 (O_900,N_9809,N_9866);
nand UO_901 (O_901,N_9923,N_9983);
or UO_902 (O_902,N_9951,N_9938);
nand UO_903 (O_903,N_9969,N_9859);
or UO_904 (O_904,N_9818,N_9878);
nand UO_905 (O_905,N_9805,N_9880);
xor UO_906 (O_906,N_9960,N_9968);
or UO_907 (O_907,N_9916,N_9928);
and UO_908 (O_908,N_9992,N_9926);
xnor UO_909 (O_909,N_9991,N_9933);
nand UO_910 (O_910,N_9867,N_9980);
and UO_911 (O_911,N_9929,N_9974);
xor UO_912 (O_912,N_9903,N_9966);
nand UO_913 (O_913,N_9806,N_9994);
nor UO_914 (O_914,N_9821,N_9847);
or UO_915 (O_915,N_9923,N_9999);
or UO_916 (O_916,N_9970,N_9915);
xor UO_917 (O_917,N_9949,N_9806);
and UO_918 (O_918,N_9928,N_9979);
nand UO_919 (O_919,N_9985,N_9816);
and UO_920 (O_920,N_9999,N_9958);
and UO_921 (O_921,N_9962,N_9811);
nor UO_922 (O_922,N_9813,N_9927);
xnor UO_923 (O_923,N_9875,N_9810);
or UO_924 (O_924,N_9914,N_9817);
nor UO_925 (O_925,N_9980,N_9834);
nor UO_926 (O_926,N_9959,N_9978);
nor UO_927 (O_927,N_9807,N_9835);
or UO_928 (O_928,N_9848,N_9923);
nand UO_929 (O_929,N_9886,N_9964);
nor UO_930 (O_930,N_9995,N_9930);
nand UO_931 (O_931,N_9974,N_9824);
nor UO_932 (O_932,N_9942,N_9838);
xor UO_933 (O_933,N_9829,N_9898);
nor UO_934 (O_934,N_9905,N_9902);
nor UO_935 (O_935,N_9938,N_9813);
nor UO_936 (O_936,N_9940,N_9846);
nand UO_937 (O_937,N_9809,N_9966);
and UO_938 (O_938,N_9914,N_9901);
or UO_939 (O_939,N_9946,N_9952);
nor UO_940 (O_940,N_9815,N_9975);
and UO_941 (O_941,N_9831,N_9946);
nor UO_942 (O_942,N_9836,N_9931);
or UO_943 (O_943,N_9907,N_9896);
and UO_944 (O_944,N_9895,N_9859);
and UO_945 (O_945,N_9869,N_9990);
or UO_946 (O_946,N_9965,N_9879);
or UO_947 (O_947,N_9990,N_9944);
or UO_948 (O_948,N_9936,N_9892);
or UO_949 (O_949,N_9808,N_9866);
and UO_950 (O_950,N_9986,N_9962);
xnor UO_951 (O_951,N_9818,N_9826);
and UO_952 (O_952,N_9912,N_9824);
or UO_953 (O_953,N_9972,N_9896);
or UO_954 (O_954,N_9901,N_9950);
xnor UO_955 (O_955,N_9813,N_9961);
and UO_956 (O_956,N_9977,N_9966);
or UO_957 (O_957,N_9873,N_9864);
nand UO_958 (O_958,N_9842,N_9835);
nor UO_959 (O_959,N_9910,N_9904);
and UO_960 (O_960,N_9921,N_9935);
nor UO_961 (O_961,N_9800,N_9807);
nor UO_962 (O_962,N_9978,N_9826);
xnor UO_963 (O_963,N_9977,N_9974);
and UO_964 (O_964,N_9834,N_9889);
or UO_965 (O_965,N_9826,N_9945);
or UO_966 (O_966,N_9844,N_9882);
and UO_967 (O_967,N_9921,N_9951);
nor UO_968 (O_968,N_9872,N_9920);
nand UO_969 (O_969,N_9948,N_9963);
xnor UO_970 (O_970,N_9824,N_9836);
nand UO_971 (O_971,N_9986,N_9941);
nand UO_972 (O_972,N_9809,N_9846);
or UO_973 (O_973,N_9818,N_9877);
xnor UO_974 (O_974,N_9892,N_9858);
xor UO_975 (O_975,N_9943,N_9985);
xor UO_976 (O_976,N_9908,N_9931);
or UO_977 (O_977,N_9851,N_9900);
nand UO_978 (O_978,N_9973,N_9935);
nand UO_979 (O_979,N_9803,N_9889);
or UO_980 (O_980,N_9808,N_9840);
or UO_981 (O_981,N_9977,N_9858);
and UO_982 (O_982,N_9880,N_9886);
nor UO_983 (O_983,N_9952,N_9954);
and UO_984 (O_984,N_9892,N_9983);
nand UO_985 (O_985,N_9835,N_9976);
or UO_986 (O_986,N_9976,N_9987);
nor UO_987 (O_987,N_9958,N_9801);
or UO_988 (O_988,N_9894,N_9834);
or UO_989 (O_989,N_9813,N_9854);
nor UO_990 (O_990,N_9836,N_9905);
nor UO_991 (O_991,N_9987,N_9930);
nand UO_992 (O_992,N_9877,N_9934);
nand UO_993 (O_993,N_9954,N_9972);
and UO_994 (O_994,N_9967,N_9881);
nor UO_995 (O_995,N_9913,N_9910);
or UO_996 (O_996,N_9979,N_9889);
and UO_997 (O_997,N_9920,N_9997);
and UO_998 (O_998,N_9842,N_9992);
nand UO_999 (O_999,N_9980,N_9962);
nand UO_1000 (O_1000,N_9835,N_9906);
and UO_1001 (O_1001,N_9932,N_9834);
xor UO_1002 (O_1002,N_9936,N_9991);
nand UO_1003 (O_1003,N_9968,N_9994);
and UO_1004 (O_1004,N_9890,N_9861);
nand UO_1005 (O_1005,N_9810,N_9927);
or UO_1006 (O_1006,N_9820,N_9874);
and UO_1007 (O_1007,N_9868,N_9995);
nor UO_1008 (O_1008,N_9976,N_9870);
xor UO_1009 (O_1009,N_9960,N_9807);
and UO_1010 (O_1010,N_9904,N_9854);
nand UO_1011 (O_1011,N_9872,N_9807);
nand UO_1012 (O_1012,N_9841,N_9969);
nand UO_1013 (O_1013,N_9906,N_9825);
or UO_1014 (O_1014,N_9913,N_9825);
nand UO_1015 (O_1015,N_9853,N_9946);
nor UO_1016 (O_1016,N_9881,N_9858);
or UO_1017 (O_1017,N_9893,N_9904);
nand UO_1018 (O_1018,N_9802,N_9888);
nand UO_1019 (O_1019,N_9841,N_9963);
xor UO_1020 (O_1020,N_9818,N_9976);
and UO_1021 (O_1021,N_9816,N_9920);
nand UO_1022 (O_1022,N_9836,N_9821);
and UO_1023 (O_1023,N_9924,N_9960);
nor UO_1024 (O_1024,N_9881,N_9884);
or UO_1025 (O_1025,N_9927,N_9847);
xnor UO_1026 (O_1026,N_9801,N_9831);
xor UO_1027 (O_1027,N_9909,N_9982);
nand UO_1028 (O_1028,N_9966,N_9900);
nor UO_1029 (O_1029,N_9987,N_9855);
and UO_1030 (O_1030,N_9991,N_9885);
nor UO_1031 (O_1031,N_9848,N_9869);
or UO_1032 (O_1032,N_9820,N_9918);
nor UO_1033 (O_1033,N_9900,N_9819);
nor UO_1034 (O_1034,N_9949,N_9981);
and UO_1035 (O_1035,N_9851,N_9886);
or UO_1036 (O_1036,N_9964,N_9979);
or UO_1037 (O_1037,N_9884,N_9869);
or UO_1038 (O_1038,N_9829,N_9891);
nand UO_1039 (O_1039,N_9877,N_9946);
or UO_1040 (O_1040,N_9826,N_9991);
nand UO_1041 (O_1041,N_9931,N_9898);
or UO_1042 (O_1042,N_9819,N_9908);
nor UO_1043 (O_1043,N_9824,N_9807);
nor UO_1044 (O_1044,N_9975,N_9830);
nand UO_1045 (O_1045,N_9933,N_9953);
nor UO_1046 (O_1046,N_9888,N_9885);
nand UO_1047 (O_1047,N_9952,N_9838);
nand UO_1048 (O_1048,N_9913,N_9918);
or UO_1049 (O_1049,N_9941,N_9841);
nor UO_1050 (O_1050,N_9842,N_9968);
and UO_1051 (O_1051,N_9971,N_9841);
nor UO_1052 (O_1052,N_9975,N_9916);
and UO_1053 (O_1053,N_9880,N_9957);
and UO_1054 (O_1054,N_9974,N_9869);
nor UO_1055 (O_1055,N_9820,N_9992);
nor UO_1056 (O_1056,N_9833,N_9989);
or UO_1057 (O_1057,N_9953,N_9960);
or UO_1058 (O_1058,N_9810,N_9919);
and UO_1059 (O_1059,N_9960,N_9926);
nor UO_1060 (O_1060,N_9879,N_9858);
xor UO_1061 (O_1061,N_9997,N_9979);
nor UO_1062 (O_1062,N_9909,N_9879);
and UO_1063 (O_1063,N_9952,N_9963);
nor UO_1064 (O_1064,N_9896,N_9957);
nand UO_1065 (O_1065,N_9985,N_9947);
or UO_1066 (O_1066,N_9810,N_9885);
and UO_1067 (O_1067,N_9818,N_9816);
and UO_1068 (O_1068,N_9994,N_9977);
nor UO_1069 (O_1069,N_9980,N_9961);
nor UO_1070 (O_1070,N_9911,N_9838);
nor UO_1071 (O_1071,N_9811,N_9970);
nand UO_1072 (O_1072,N_9920,N_9912);
nor UO_1073 (O_1073,N_9876,N_9957);
xor UO_1074 (O_1074,N_9963,N_9959);
nand UO_1075 (O_1075,N_9995,N_9908);
and UO_1076 (O_1076,N_9910,N_9845);
nor UO_1077 (O_1077,N_9820,N_9915);
nand UO_1078 (O_1078,N_9808,N_9906);
or UO_1079 (O_1079,N_9932,N_9852);
nand UO_1080 (O_1080,N_9986,N_9987);
and UO_1081 (O_1081,N_9877,N_9944);
and UO_1082 (O_1082,N_9943,N_9912);
nor UO_1083 (O_1083,N_9825,N_9881);
and UO_1084 (O_1084,N_9835,N_9967);
nand UO_1085 (O_1085,N_9930,N_9870);
nand UO_1086 (O_1086,N_9996,N_9873);
or UO_1087 (O_1087,N_9982,N_9886);
nor UO_1088 (O_1088,N_9803,N_9928);
and UO_1089 (O_1089,N_9923,N_9834);
and UO_1090 (O_1090,N_9957,N_9976);
or UO_1091 (O_1091,N_9919,N_9951);
and UO_1092 (O_1092,N_9828,N_9842);
or UO_1093 (O_1093,N_9971,N_9845);
and UO_1094 (O_1094,N_9865,N_9807);
xnor UO_1095 (O_1095,N_9929,N_9978);
nand UO_1096 (O_1096,N_9873,N_9814);
or UO_1097 (O_1097,N_9966,N_9862);
nor UO_1098 (O_1098,N_9847,N_9946);
nor UO_1099 (O_1099,N_9800,N_9970);
and UO_1100 (O_1100,N_9926,N_9928);
and UO_1101 (O_1101,N_9909,N_9862);
and UO_1102 (O_1102,N_9918,N_9876);
nor UO_1103 (O_1103,N_9986,N_9910);
nor UO_1104 (O_1104,N_9832,N_9999);
xor UO_1105 (O_1105,N_9956,N_9938);
nand UO_1106 (O_1106,N_9999,N_9814);
nor UO_1107 (O_1107,N_9988,N_9801);
nor UO_1108 (O_1108,N_9899,N_9849);
and UO_1109 (O_1109,N_9921,N_9897);
and UO_1110 (O_1110,N_9933,N_9909);
nand UO_1111 (O_1111,N_9933,N_9825);
nor UO_1112 (O_1112,N_9916,N_9929);
nand UO_1113 (O_1113,N_9925,N_9888);
nor UO_1114 (O_1114,N_9990,N_9972);
xor UO_1115 (O_1115,N_9888,N_9868);
or UO_1116 (O_1116,N_9874,N_9950);
and UO_1117 (O_1117,N_9944,N_9892);
or UO_1118 (O_1118,N_9820,N_9979);
nor UO_1119 (O_1119,N_9984,N_9902);
and UO_1120 (O_1120,N_9902,N_9974);
and UO_1121 (O_1121,N_9867,N_9883);
or UO_1122 (O_1122,N_9963,N_9973);
xor UO_1123 (O_1123,N_9856,N_9969);
nor UO_1124 (O_1124,N_9932,N_9806);
and UO_1125 (O_1125,N_9871,N_9907);
xor UO_1126 (O_1126,N_9917,N_9925);
or UO_1127 (O_1127,N_9917,N_9878);
nor UO_1128 (O_1128,N_9819,N_9913);
and UO_1129 (O_1129,N_9877,N_9922);
and UO_1130 (O_1130,N_9850,N_9912);
or UO_1131 (O_1131,N_9878,N_9919);
and UO_1132 (O_1132,N_9988,N_9892);
nand UO_1133 (O_1133,N_9946,N_9919);
nor UO_1134 (O_1134,N_9951,N_9964);
or UO_1135 (O_1135,N_9826,N_9824);
nor UO_1136 (O_1136,N_9983,N_9978);
and UO_1137 (O_1137,N_9824,N_9832);
and UO_1138 (O_1138,N_9840,N_9862);
nand UO_1139 (O_1139,N_9987,N_9805);
and UO_1140 (O_1140,N_9864,N_9872);
and UO_1141 (O_1141,N_9876,N_9854);
nand UO_1142 (O_1142,N_9931,N_9876);
nor UO_1143 (O_1143,N_9904,N_9919);
nor UO_1144 (O_1144,N_9895,N_9821);
nand UO_1145 (O_1145,N_9882,N_9997);
or UO_1146 (O_1146,N_9955,N_9833);
or UO_1147 (O_1147,N_9918,N_9907);
nand UO_1148 (O_1148,N_9992,N_9990);
nor UO_1149 (O_1149,N_9834,N_9970);
and UO_1150 (O_1150,N_9945,N_9885);
or UO_1151 (O_1151,N_9991,N_9981);
and UO_1152 (O_1152,N_9828,N_9931);
nand UO_1153 (O_1153,N_9934,N_9899);
nand UO_1154 (O_1154,N_9889,N_9982);
and UO_1155 (O_1155,N_9860,N_9859);
xnor UO_1156 (O_1156,N_9912,N_9986);
nand UO_1157 (O_1157,N_9982,N_9859);
xnor UO_1158 (O_1158,N_9886,N_9992);
and UO_1159 (O_1159,N_9860,N_9819);
nor UO_1160 (O_1160,N_9818,N_9841);
nor UO_1161 (O_1161,N_9891,N_9818);
or UO_1162 (O_1162,N_9928,N_9835);
nand UO_1163 (O_1163,N_9945,N_9967);
xor UO_1164 (O_1164,N_9920,N_9823);
nor UO_1165 (O_1165,N_9977,N_9869);
or UO_1166 (O_1166,N_9862,N_9959);
nand UO_1167 (O_1167,N_9820,N_9802);
nor UO_1168 (O_1168,N_9937,N_9881);
or UO_1169 (O_1169,N_9932,N_9827);
nor UO_1170 (O_1170,N_9963,N_9982);
xor UO_1171 (O_1171,N_9828,N_9896);
nor UO_1172 (O_1172,N_9889,N_9956);
or UO_1173 (O_1173,N_9875,N_9933);
nor UO_1174 (O_1174,N_9997,N_9875);
or UO_1175 (O_1175,N_9940,N_9913);
nor UO_1176 (O_1176,N_9925,N_9903);
and UO_1177 (O_1177,N_9977,N_9911);
and UO_1178 (O_1178,N_9894,N_9990);
and UO_1179 (O_1179,N_9855,N_9807);
nand UO_1180 (O_1180,N_9885,N_9979);
and UO_1181 (O_1181,N_9847,N_9960);
nor UO_1182 (O_1182,N_9843,N_9918);
and UO_1183 (O_1183,N_9891,N_9908);
nand UO_1184 (O_1184,N_9966,N_9974);
or UO_1185 (O_1185,N_9826,N_9934);
nor UO_1186 (O_1186,N_9833,N_9908);
nand UO_1187 (O_1187,N_9870,N_9805);
nor UO_1188 (O_1188,N_9989,N_9916);
and UO_1189 (O_1189,N_9928,N_9810);
xor UO_1190 (O_1190,N_9910,N_9968);
nand UO_1191 (O_1191,N_9930,N_9876);
xnor UO_1192 (O_1192,N_9842,N_9853);
and UO_1193 (O_1193,N_9994,N_9824);
and UO_1194 (O_1194,N_9884,N_9923);
nor UO_1195 (O_1195,N_9886,N_9979);
nand UO_1196 (O_1196,N_9905,N_9952);
or UO_1197 (O_1197,N_9856,N_9949);
nand UO_1198 (O_1198,N_9902,N_9953);
and UO_1199 (O_1199,N_9836,N_9915);
nand UO_1200 (O_1200,N_9801,N_9982);
xnor UO_1201 (O_1201,N_9994,N_9844);
nand UO_1202 (O_1202,N_9952,N_9805);
or UO_1203 (O_1203,N_9927,N_9940);
nor UO_1204 (O_1204,N_9873,N_9880);
xnor UO_1205 (O_1205,N_9958,N_9906);
nand UO_1206 (O_1206,N_9942,N_9880);
and UO_1207 (O_1207,N_9842,N_9950);
nor UO_1208 (O_1208,N_9853,N_9950);
nand UO_1209 (O_1209,N_9833,N_9985);
or UO_1210 (O_1210,N_9950,N_9830);
nor UO_1211 (O_1211,N_9953,N_9971);
nand UO_1212 (O_1212,N_9840,N_9849);
and UO_1213 (O_1213,N_9859,N_9904);
and UO_1214 (O_1214,N_9901,N_9898);
nand UO_1215 (O_1215,N_9817,N_9963);
xor UO_1216 (O_1216,N_9871,N_9976);
nand UO_1217 (O_1217,N_9916,N_9994);
and UO_1218 (O_1218,N_9969,N_9948);
nor UO_1219 (O_1219,N_9847,N_9973);
nand UO_1220 (O_1220,N_9954,N_9898);
or UO_1221 (O_1221,N_9833,N_9925);
nand UO_1222 (O_1222,N_9972,N_9877);
nand UO_1223 (O_1223,N_9958,N_9988);
nor UO_1224 (O_1224,N_9802,N_9838);
nand UO_1225 (O_1225,N_9924,N_9927);
nor UO_1226 (O_1226,N_9974,N_9839);
or UO_1227 (O_1227,N_9988,N_9946);
nor UO_1228 (O_1228,N_9953,N_9872);
nand UO_1229 (O_1229,N_9904,N_9883);
or UO_1230 (O_1230,N_9951,N_9941);
xnor UO_1231 (O_1231,N_9825,N_9894);
nor UO_1232 (O_1232,N_9938,N_9867);
and UO_1233 (O_1233,N_9908,N_9946);
xor UO_1234 (O_1234,N_9841,N_9819);
nand UO_1235 (O_1235,N_9882,N_9877);
nor UO_1236 (O_1236,N_9973,N_9946);
or UO_1237 (O_1237,N_9830,N_9926);
nand UO_1238 (O_1238,N_9986,N_9922);
nor UO_1239 (O_1239,N_9865,N_9867);
nand UO_1240 (O_1240,N_9915,N_9910);
and UO_1241 (O_1241,N_9808,N_9948);
and UO_1242 (O_1242,N_9964,N_9891);
and UO_1243 (O_1243,N_9958,N_9919);
or UO_1244 (O_1244,N_9845,N_9920);
nand UO_1245 (O_1245,N_9862,N_9858);
nor UO_1246 (O_1246,N_9903,N_9829);
nand UO_1247 (O_1247,N_9938,N_9982);
xor UO_1248 (O_1248,N_9931,N_9866);
and UO_1249 (O_1249,N_9809,N_9819);
nand UO_1250 (O_1250,N_9925,N_9829);
and UO_1251 (O_1251,N_9804,N_9829);
xor UO_1252 (O_1252,N_9975,N_9843);
nand UO_1253 (O_1253,N_9967,N_9830);
or UO_1254 (O_1254,N_9954,N_9935);
and UO_1255 (O_1255,N_9874,N_9964);
nand UO_1256 (O_1256,N_9910,N_9801);
nor UO_1257 (O_1257,N_9868,N_9944);
and UO_1258 (O_1258,N_9963,N_9927);
and UO_1259 (O_1259,N_9973,N_9819);
nor UO_1260 (O_1260,N_9945,N_9834);
nand UO_1261 (O_1261,N_9997,N_9878);
nand UO_1262 (O_1262,N_9949,N_9943);
or UO_1263 (O_1263,N_9950,N_9992);
or UO_1264 (O_1264,N_9987,N_9958);
or UO_1265 (O_1265,N_9843,N_9932);
xnor UO_1266 (O_1266,N_9822,N_9969);
or UO_1267 (O_1267,N_9864,N_9927);
and UO_1268 (O_1268,N_9888,N_9846);
or UO_1269 (O_1269,N_9885,N_9983);
nor UO_1270 (O_1270,N_9999,N_9973);
nand UO_1271 (O_1271,N_9875,N_9921);
or UO_1272 (O_1272,N_9981,N_9983);
nor UO_1273 (O_1273,N_9880,N_9995);
or UO_1274 (O_1274,N_9857,N_9933);
nor UO_1275 (O_1275,N_9920,N_9830);
or UO_1276 (O_1276,N_9809,N_9850);
and UO_1277 (O_1277,N_9827,N_9889);
or UO_1278 (O_1278,N_9947,N_9831);
or UO_1279 (O_1279,N_9995,N_9829);
nor UO_1280 (O_1280,N_9945,N_9919);
nand UO_1281 (O_1281,N_9854,N_9897);
and UO_1282 (O_1282,N_9885,N_9918);
xnor UO_1283 (O_1283,N_9839,N_9863);
nand UO_1284 (O_1284,N_9858,N_9961);
xnor UO_1285 (O_1285,N_9876,N_9894);
nor UO_1286 (O_1286,N_9866,N_9942);
nand UO_1287 (O_1287,N_9863,N_9995);
or UO_1288 (O_1288,N_9933,N_9907);
nor UO_1289 (O_1289,N_9905,N_9993);
nand UO_1290 (O_1290,N_9850,N_9955);
nor UO_1291 (O_1291,N_9967,N_9841);
nor UO_1292 (O_1292,N_9986,N_9898);
xor UO_1293 (O_1293,N_9963,N_9949);
or UO_1294 (O_1294,N_9805,N_9867);
and UO_1295 (O_1295,N_9929,N_9812);
nor UO_1296 (O_1296,N_9922,N_9858);
and UO_1297 (O_1297,N_9938,N_9960);
nand UO_1298 (O_1298,N_9860,N_9879);
and UO_1299 (O_1299,N_9924,N_9881);
nor UO_1300 (O_1300,N_9897,N_9941);
xnor UO_1301 (O_1301,N_9917,N_9857);
and UO_1302 (O_1302,N_9847,N_9944);
or UO_1303 (O_1303,N_9925,N_9943);
or UO_1304 (O_1304,N_9872,N_9937);
nor UO_1305 (O_1305,N_9955,N_9943);
xor UO_1306 (O_1306,N_9927,N_9876);
nor UO_1307 (O_1307,N_9852,N_9865);
or UO_1308 (O_1308,N_9969,N_9850);
nand UO_1309 (O_1309,N_9899,N_9931);
nor UO_1310 (O_1310,N_9984,N_9951);
or UO_1311 (O_1311,N_9808,N_9977);
or UO_1312 (O_1312,N_9907,N_9936);
nand UO_1313 (O_1313,N_9865,N_9904);
nor UO_1314 (O_1314,N_9822,N_9819);
nor UO_1315 (O_1315,N_9975,N_9961);
or UO_1316 (O_1316,N_9851,N_9937);
xor UO_1317 (O_1317,N_9989,N_9827);
nor UO_1318 (O_1318,N_9924,N_9889);
nand UO_1319 (O_1319,N_9914,N_9819);
or UO_1320 (O_1320,N_9975,N_9899);
nand UO_1321 (O_1321,N_9820,N_9810);
nor UO_1322 (O_1322,N_9847,N_9928);
and UO_1323 (O_1323,N_9915,N_9978);
xnor UO_1324 (O_1324,N_9991,N_9870);
nor UO_1325 (O_1325,N_9802,N_9908);
nor UO_1326 (O_1326,N_9822,N_9924);
nor UO_1327 (O_1327,N_9813,N_9983);
and UO_1328 (O_1328,N_9928,N_9867);
and UO_1329 (O_1329,N_9801,N_9920);
nor UO_1330 (O_1330,N_9816,N_9991);
and UO_1331 (O_1331,N_9905,N_9858);
and UO_1332 (O_1332,N_9927,N_9805);
and UO_1333 (O_1333,N_9947,N_9939);
and UO_1334 (O_1334,N_9847,N_9910);
or UO_1335 (O_1335,N_9964,N_9810);
nor UO_1336 (O_1336,N_9833,N_9950);
or UO_1337 (O_1337,N_9864,N_9960);
or UO_1338 (O_1338,N_9844,N_9922);
nand UO_1339 (O_1339,N_9961,N_9806);
nor UO_1340 (O_1340,N_9883,N_9831);
and UO_1341 (O_1341,N_9930,N_9857);
and UO_1342 (O_1342,N_9896,N_9991);
nand UO_1343 (O_1343,N_9967,N_9855);
or UO_1344 (O_1344,N_9828,N_9823);
or UO_1345 (O_1345,N_9852,N_9971);
nand UO_1346 (O_1346,N_9972,N_9969);
or UO_1347 (O_1347,N_9873,N_9867);
or UO_1348 (O_1348,N_9903,N_9938);
nor UO_1349 (O_1349,N_9950,N_9975);
and UO_1350 (O_1350,N_9870,N_9913);
nor UO_1351 (O_1351,N_9991,N_9994);
or UO_1352 (O_1352,N_9912,N_9965);
and UO_1353 (O_1353,N_9864,N_9919);
nand UO_1354 (O_1354,N_9960,N_9941);
nand UO_1355 (O_1355,N_9964,N_9833);
or UO_1356 (O_1356,N_9974,N_9958);
and UO_1357 (O_1357,N_9939,N_9830);
nor UO_1358 (O_1358,N_9952,N_9806);
nor UO_1359 (O_1359,N_9943,N_9942);
nor UO_1360 (O_1360,N_9834,N_9946);
nand UO_1361 (O_1361,N_9903,N_9907);
nor UO_1362 (O_1362,N_9901,N_9896);
nand UO_1363 (O_1363,N_9903,N_9952);
and UO_1364 (O_1364,N_9897,N_9826);
nor UO_1365 (O_1365,N_9868,N_9870);
nor UO_1366 (O_1366,N_9842,N_9863);
or UO_1367 (O_1367,N_9879,N_9847);
nand UO_1368 (O_1368,N_9911,N_9870);
nor UO_1369 (O_1369,N_9915,N_9989);
nor UO_1370 (O_1370,N_9881,N_9824);
nor UO_1371 (O_1371,N_9842,N_9846);
nor UO_1372 (O_1372,N_9859,N_9851);
or UO_1373 (O_1373,N_9893,N_9908);
or UO_1374 (O_1374,N_9890,N_9803);
nor UO_1375 (O_1375,N_9967,N_9878);
and UO_1376 (O_1376,N_9823,N_9992);
xor UO_1377 (O_1377,N_9848,N_9843);
nand UO_1378 (O_1378,N_9945,N_9853);
or UO_1379 (O_1379,N_9879,N_9856);
and UO_1380 (O_1380,N_9818,N_9973);
nor UO_1381 (O_1381,N_9927,N_9999);
nor UO_1382 (O_1382,N_9805,N_9891);
or UO_1383 (O_1383,N_9899,N_9994);
nand UO_1384 (O_1384,N_9902,N_9956);
nand UO_1385 (O_1385,N_9820,N_9885);
nor UO_1386 (O_1386,N_9958,N_9990);
xnor UO_1387 (O_1387,N_9814,N_9963);
nor UO_1388 (O_1388,N_9831,N_9999);
and UO_1389 (O_1389,N_9812,N_9866);
or UO_1390 (O_1390,N_9958,N_9966);
xor UO_1391 (O_1391,N_9950,N_9895);
and UO_1392 (O_1392,N_9850,N_9882);
and UO_1393 (O_1393,N_9894,N_9968);
or UO_1394 (O_1394,N_9844,N_9863);
nand UO_1395 (O_1395,N_9830,N_9867);
nand UO_1396 (O_1396,N_9912,N_9990);
xor UO_1397 (O_1397,N_9963,N_9974);
xor UO_1398 (O_1398,N_9918,N_9961);
or UO_1399 (O_1399,N_9925,N_9896);
and UO_1400 (O_1400,N_9979,N_9844);
or UO_1401 (O_1401,N_9847,N_9867);
nand UO_1402 (O_1402,N_9838,N_9907);
or UO_1403 (O_1403,N_9927,N_9921);
and UO_1404 (O_1404,N_9877,N_9806);
and UO_1405 (O_1405,N_9958,N_9875);
nand UO_1406 (O_1406,N_9875,N_9900);
or UO_1407 (O_1407,N_9820,N_9955);
nor UO_1408 (O_1408,N_9910,N_9944);
nand UO_1409 (O_1409,N_9995,N_9830);
xnor UO_1410 (O_1410,N_9812,N_9900);
xnor UO_1411 (O_1411,N_9933,N_9828);
nand UO_1412 (O_1412,N_9812,N_9954);
xor UO_1413 (O_1413,N_9959,N_9989);
nor UO_1414 (O_1414,N_9841,N_9889);
nor UO_1415 (O_1415,N_9837,N_9955);
or UO_1416 (O_1416,N_9982,N_9876);
and UO_1417 (O_1417,N_9955,N_9842);
nor UO_1418 (O_1418,N_9820,N_9983);
or UO_1419 (O_1419,N_9821,N_9829);
xor UO_1420 (O_1420,N_9828,N_9841);
nand UO_1421 (O_1421,N_9819,N_9832);
xor UO_1422 (O_1422,N_9813,N_9874);
xor UO_1423 (O_1423,N_9905,N_9909);
and UO_1424 (O_1424,N_9852,N_9815);
and UO_1425 (O_1425,N_9944,N_9806);
nand UO_1426 (O_1426,N_9886,N_9855);
and UO_1427 (O_1427,N_9999,N_9945);
nor UO_1428 (O_1428,N_9925,N_9991);
nand UO_1429 (O_1429,N_9888,N_9850);
nand UO_1430 (O_1430,N_9975,N_9868);
and UO_1431 (O_1431,N_9943,N_9979);
and UO_1432 (O_1432,N_9942,N_9939);
xor UO_1433 (O_1433,N_9949,N_9895);
xor UO_1434 (O_1434,N_9968,N_9961);
and UO_1435 (O_1435,N_9820,N_9837);
or UO_1436 (O_1436,N_9872,N_9912);
nor UO_1437 (O_1437,N_9813,N_9830);
or UO_1438 (O_1438,N_9972,N_9875);
or UO_1439 (O_1439,N_9982,N_9979);
nand UO_1440 (O_1440,N_9951,N_9904);
or UO_1441 (O_1441,N_9894,N_9942);
and UO_1442 (O_1442,N_9859,N_9973);
or UO_1443 (O_1443,N_9982,N_9883);
nor UO_1444 (O_1444,N_9958,N_9832);
and UO_1445 (O_1445,N_9926,N_9815);
and UO_1446 (O_1446,N_9909,N_9837);
or UO_1447 (O_1447,N_9875,N_9982);
nand UO_1448 (O_1448,N_9911,N_9817);
nand UO_1449 (O_1449,N_9811,N_9894);
or UO_1450 (O_1450,N_9973,N_9846);
and UO_1451 (O_1451,N_9913,N_9908);
nor UO_1452 (O_1452,N_9828,N_9916);
nor UO_1453 (O_1453,N_9801,N_9991);
nor UO_1454 (O_1454,N_9960,N_9857);
nor UO_1455 (O_1455,N_9806,N_9872);
nor UO_1456 (O_1456,N_9945,N_9849);
and UO_1457 (O_1457,N_9952,N_9950);
nor UO_1458 (O_1458,N_9893,N_9876);
xnor UO_1459 (O_1459,N_9833,N_9846);
and UO_1460 (O_1460,N_9870,N_9932);
nor UO_1461 (O_1461,N_9858,N_9919);
or UO_1462 (O_1462,N_9925,N_9904);
and UO_1463 (O_1463,N_9992,N_9800);
nand UO_1464 (O_1464,N_9998,N_9814);
or UO_1465 (O_1465,N_9839,N_9968);
nand UO_1466 (O_1466,N_9955,N_9821);
nand UO_1467 (O_1467,N_9950,N_9834);
xor UO_1468 (O_1468,N_9955,N_9998);
nor UO_1469 (O_1469,N_9960,N_9849);
xor UO_1470 (O_1470,N_9967,N_9834);
nand UO_1471 (O_1471,N_9830,N_9831);
nand UO_1472 (O_1472,N_9836,N_9923);
xnor UO_1473 (O_1473,N_9838,N_9816);
nor UO_1474 (O_1474,N_9995,N_9937);
xnor UO_1475 (O_1475,N_9815,N_9972);
and UO_1476 (O_1476,N_9811,N_9826);
nand UO_1477 (O_1477,N_9968,N_9933);
and UO_1478 (O_1478,N_9964,N_9894);
xor UO_1479 (O_1479,N_9847,N_9871);
nor UO_1480 (O_1480,N_9839,N_9953);
or UO_1481 (O_1481,N_9925,N_9870);
nand UO_1482 (O_1482,N_9852,N_9850);
xnor UO_1483 (O_1483,N_9859,N_9864);
or UO_1484 (O_1484,N_9994,N_9871);
and UO_1485 (O_1485,N_9868,N_9962);
and UO_1486 (O_1486,N_9973,N_9845);
and UO_1487 (O_1487,N_9918,N_9935);
nand UO_1488 (O_1488,N_9918,N_9879);
and UO_1489 (O_1489,N_9856,N_9977);
xor UO_1490 (O_1490,N_9808,N_9968);
xor UO_1491 (O_1491,N_9932,N_9895);
and UO_1492 (O_1492,N_9892,N_9879);
nand UO_1493 (O_1493,N_9836,N_9941);
nand UO_1494 (O_1494,N_9893,N_9889);
and UO_1495 (O_1495,N_9959,N_9867);
nor UO_1496 (O_1496,N_9988,N_9936);
nand UO_1497 (O_1497,N_9826,N_9801);
and UO_1498 (O_1498,N_9833,N_9829);
nor UO_1499 (O_1499,N_9935,N_9984);
endmodule