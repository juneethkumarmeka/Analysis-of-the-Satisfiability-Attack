module basic_750_5000_1000_10_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_237,In_487);
nand U1 (N_1,In_397,In_718);
nand U2 (N_2,In_591,In_406);
nor U3 (N_3,In_459,In_292);
nand U4 (N_4,In_40,In_223);
or U5 (N_5,In_144,In_364);
nor U6 (N_6,In_561,In_113);
or U7 (N_7,In_742,In_469);
nor U8 (N_8,In_383,In_568);
and U9 (N_9,In_116,In_8);
xor U10 (N_10,In_138,In_0);
xor U11 (N_11,In_282,In_450);
xor U12 (N_12,In_644,In_21);
or U13 (N_13,In_576,In_458);
nand U14 (N_14,In_334,In_102);
xor U15 (N_15,In_47,In_638);
nor U16 (N_16,In_678,In_689);
or U17 (N_17,In_225,In_79);
or U18 (N_18,In_748,In_257);
or U19 (N_19,In_457,In_170);
or U20 (N_20,In_354,In_196);
and U21 (N_21,In_268,In_195);
nand U22 (N_22,In_508,In_424);
nor U23 (N_23,In_695,In_496);
nand U24 (N_24,In_400,In_68);
and U25 (N_25,In_372,In_28);
or U26 (N_26,In_405,In_577);
nor U27 (N_27,In_410,In_722);
nand U28 (N_28,In_376,In_470);
and U29 (N_29,In_640,In_584);
and U30 (N_30,In_218,In_207);
and U31 (N_31,In_312,In_686);
or U32 (N_32,In_698,In_671);
nor U33 (N_33,In_523,In_357);
xnor U34 (N_34,In_130,In_666);
xor U35 (N_35,In_380,In_669);
and U36 (N_36,In_88,In_509);
xor U37 (N_37,In_41,In_134);
or U38 (N_38,In_707,In_513);
nand U39 (N_39,In_726,In_139);
nor U40 (N_40,In_146,In_579);
and U41 (N_41,In_180,In_403);
and U42 (N_42,In_3,In_495);
and U43 (N_43,In_586,In_433);
nand U44 (N_44,In_349,In_499);
nor U45 (N_45,In_125,In_95);
or U46 (N_46,In_725,In_562);
and U47 (N_47,In_647,In_55);
nand U48 (N_48,In_539,In_362);
or U49 (N_49,In_169,In_652);
and U50 (N_50,In_556,In_174);
nor U51 (N_51,In_699,In_384);
nand U52 (N_52,In_122,In_460);
and U53 (N_53,In_327,In_105);
or U54 (N_54,In_273,In_710);
and U55 (N_55,In_645,In_685);
or U56 (N_56,In_235,In_287);
and U57 (N_57,In_446,In_598);
nor U58 (N_58,In_542,In_330);
or U59 (N_59,In_254,In_522);
nand U60 (N_60,In_297,In_507);
nand U61 (N_61,In_503,In_515);
xnor U62 (N_62,In_226,In_590);
nand U63 (N_63,In_86,In_356);
nand U64 (N_64,In_733,In_461);
nor U65 (N_65,In_673,In_31);
xor U66 (N_66,In_670,In_94);
xnor U67 (N_67,In_259,In_262);
or U68 (N_68,In_531,In_567);
or U69 (N_69,In_6,In_176);
and U70 (N_70,In_385,In_296);
xnor U71 (N_71,In_602,In_549);
or U72 (N_72,In_680,In_119);
nand U73 (N_73,In_730,In_10);
xnor U74 (N_74,In_683,In_552);
or U75 (N_75,In_46,In_307);
and U76 (N_76,In_548,In_52);
or U77 (N_77,In_100,In_66);
or U78 (N_78,In_304,In_555);
and U79 (N_79,In_360,In_624);
or U80 (N_80,In_621,In_493);
or U81 (N_81,In_368,In_289);
nor U82 (N_82,In_172,In_107);
nor U83 (N_83,In_98,In_227);
or U84 (N_84,In_603,In_366);
nand U85 (N_85,In_242,In_738);
nand U86 (N_86,In_328,In_474);
and U87 (N_87,In_33,In_343);
nand U88 (N_88,In_715,In_371);
or U89 (N_89,In_264,In_168);
and U90 (N_90,In_581,In_422);
or U91 (N_91,In_676,In_155);
xor U92 (N_92,In_353,In_613);
nor U93 (N_93,In_202,In_420);
nand U94 (N_94,In_339,In_73);
nor U95 (N_95,In_142,In_510);
and U96 (N_96,In_261,In_608);
xor U97 (N_97,In_409,In_281);
xnor U98 (N_98,In_34,In_65);
and U99 (N_99,In_582,In_189);
nor U100 (N_100,In_49,In_306);
and U101 (N_101,In_451,In_89);
or U102 (N_102,In_150,In_244);
nand U103 (N_103,In_314,In_173);
and U104 (N_104,In_336,In_43);
or U105 (N_105,In_213,In_121);
nand U106 (N_106,In_60,In_625);
nor U107 (N_107,In_56,In_432);
xnor U108 (N_108,In_533,In_19);
or U109 (N_109,In_443,In_69);
or U110 (N_110,In_240,In_61);
nor U111 (N_111,In_452,In_723);
and U112 (N_112,In_529,In_50);
nand U113 (N_113,In_250,In_601);
nand U114 (N_114,In_160,In_425);
nand U115 (N_115,In_192,In_688);
nor U116 (N_116,In_18,In_4);
or U117 (N_117,In_232,In_208);
nand U118 (N_118,In_401,In_284);
or U119 (N_119,In_30,In_702);
and U120 (N_120,In_572,In_315);
or U121 (N_121,In_367,In_544);
nand U122 (N_122,In_481,In_378);
nand U123 (N_123,In_57,In_274);
and U124 (N_124,In_426,In_106);
nor U125 (N_125,In_323,In_236);
xnor U126 (N_126,In_298,In_662);
nor U127 (N_127,In_361,In_635);
nand U128 (N_128,In_233,In_692);
nand U129 (N_129,In_220,In_390);
nor U130 (N_130,In_436,In_74);
or U131 (N_131,In_338,In_634);
xor U132 (N_132,In_394,In_583);
and U133 (N_133,In_124,In_472);
nor U134 (N_134,In_418,In_566);
or U135 (N_135,In_82,In_157);
or U136 (N_136,In_191,In_594);
nand U137 (N_137,In_546,In_329);
nor U138 (N_138,In_745,In_27);
or U139 (N_139,In_265,In_414);
and U140 (N_140,In_99,In_325);
xor U141 (N_141,In_153,In_341);
xor U142 (N_142,In_188,In_524);
and U143 (N_143,In_628,In_267);
and U144 (N_144,In_553,In_141);
or U145 (N_145,In_616,In_462);
or U146 (N_146,In_416,In_109);
and U147 (N_147,In_363,In_381);
nor U148 (N_148,In_187,In_468);
xor U149 (N_149,In_521,In_578);
nor U150 (N_150,In_498,In_276);
nand U151 (N_151,In_517,In_681);
xnor U152 (N_152,In_76,In_547);
or U153 (N_153,In_216,In_305);
nand U154 (N_154,In_388,In_744);
nor U155 (N_155,In_739,In_610);
xnor U156 (N_156,In_271,In_534);
or U157 (N_157,In_90,In_427);
xnor U158 (N_158,In_743,In_270);
xor U159 (N_159,In_340,In_145);
nor U160 (N_160,In_588,In_351);
xor U161 (N_161,In_181,In_252);
nand U162 (N_162,In_708,In_112);
xnor U163 (N_163,In_263,In_646);
or U164 (N_164,In_516,In_171);
xor U165 (N_165,In_75,In_412);
nor U166 (N_166,In_664,In_177);
or U167 (N_167,In_637,In_313);
and U168 (N_168,In_488,In_101);
or U169 (N_169,In_727,In_489);
xor U170 (N_170,In_434,In_348);
or U171 (N_171,In_617,In_123);
xnor U172 (N_172,In_612,In_311);
xnor U173 (N_173,In_285,In_655);
nor U174 (N_174,In_614,In_622);
nor U175 (N_175,In_9,In_667);
and U176 (N_176,In_701,In_476);
nand U177 (N_177,In_370,In_447);
nor U178 (N_178,In_435,In_280);
or U179 (N_179,In_221,In_258);
or U180 (N_180,In_632,In_355);
nand U181 (N_181,In_194,In_300);
nor U182 (N_182,In_619,In_375);
and U183 (N_183,In_600,In_149);
nand U184 (N_184,In_580,In_319);
and U185 (N_185,In_127,In_716);
or U186 (N_186,In_64,In_550);
nor U187 (N_187,In_26,In_557);
nor U188 (N_188,In_411,In_293);
xnor U189 (N_189,In_231,In_663);
nand U190 (N_190,In_445,In_299);
nand U191 (N_191,In_536,In_456);
nor U192 (N_192,In_455,In_431);
or U193 (N_193,In_543,In_747);
xor U194 (N_194,In_440,In_224);
or U195 (N_195,In_165,In_120);
xor U196 (N_196,In_633,In_211);
nand U197 (N_197,In_132,In_545);
nand U198 (N_198,In_627,In_136);
xnor U199 (N_199,In_477,In_479);
nand U200 (N_200,In_604,In_260);
or U201 (N_201,In_396,In_358);
nor U202 (N_202,In_316,In_618);
xnor U203 (N_203,In_42,In_210);
and U204 (N_204,In_501,In_696);
xor U205 (N_205,In_288,In_596);
or U206 (N_206,In_156,In_185);
xor U207 (N_207,In_597,In_737);
nand U208 (N_208,In_143,In_642);
nor U209 (N_209,In_317,In_190);
nor U210 (N_210,In_255,In_514);
or U211 (N_211,In_203,In_565);
xor U212 (N_212,In_247,In_650);
xor U213 (N_213,In_643,In_337);
and U214 (N_214,In_217,In_654);
xor U215 (N_215,In_379,In_511);
xnor U216 (N_216,In_653,In_11);
xnor U217 (N_217,In_482,In_72);
nand U218 (N_218,In_326,In_2);
nor U219 (N_219,In_81,In_660);
nand U220 (N_220,In_421,In_117);
or U221 (N_221,In_148,In_661);
or U222 (N_222,In_592,In_344);
nor U223 (N_223,In_24,In_359);
nand U224 (N_224,In_465,In_694);
or U225 (N_225,In_80,In_229);
or U226 (N_226,In_182,In_20);
or U227 (N_227,In_444,In_346);
xnor U228 (N_228,In_453,In_721);
xnor U229 (N_229,In_682,In_519);
nor U230 (N_230,In_115,In_712);
xor U231 (N_231,In_184,In_746);
or U232 (N_232,In_570,In_478);
xor U233 (N_233,In_677,In_502);
nor U234 (N_234,In_96,In_729);
xor U235 (N_235,In_159,In_15);
nand U236 (N_236,In_54,In_466);
or U237 (N_237,In_560,In_67);
nor U238 (N_238,In_735,In_415);
nand U239 (N_239,In_137,In_520);
xnor U240 (N_240,In_44,In_538);
and U241 (N_241,In_286,In_162);
nor U242 (N_242,In_291,In_571);
nand U243 (N_243,In_486,In_719);
nand U244 (N_244,In_331,In_587);
xor U245 (N_245,In_382,In_183);
nand U246 (N_246,In_126,In_442);
or U247 (N_247,In_279,In_438);
and U248 (N_248,In_528,In_131);
and U249 (N_249,In_639,In_302);
xnor U250 (N_250,In_275,In_104);
or U251 (N_251,In_214,In_175);
nor U252 (N_252,In_392,In_103);
xnor U253 (N_253,In_193,In_352);
or U254 (N_254,In_732,In_483);
nand U255 (N_255,In_741,In_186);
and U256 (N_256,In_204,In_166);
and U257 (N_257,In_535,In_554);
or U258 (N_258,In_25,In_29);
xnor U259 (N_259,In_164,In_665);
nand U260 (N_260,In_1,In_249);
nand U261 (N_261,In_391,In_711);
xnor U262 (N_262,In_439,In_350);
nand U263 (N_263,In_256,In_253);
and U264 (N_264,In_705,In_114);
nor U265 (N_265,In_111,In_239);
and U266 (N_266,In_321,In_630);
and U267 (N_267,In_734,In_151);
xnor U268 (N_268,In_248,In_212);
nand U269 (N_269,In_724,In_309);
and U270 (N_270,In_527,In_691);
xor U271 (N_271,In_687,In_318);
nor U272 (N_272,In_518,In_238);
or U273 (N_273,In_564,In_492);
nand U274 (N_274,In_428,In_389);
nor U275 (N_275,In_684,In_78);
xor U276 (N_276,In_574,In_679);
xnor U277 (N_277,In_110,In_205);
xor U278 (N_278,In_266,In_589);
nand U279 (N_279,In_697,In_200);
and U280 (N_280,In_278,In_595);
xor U281 (N_281,In_463,In_310);
nor U282 (N_282,In_45,In_402);
xnor U283 (N_283,In_430,In_467);
nor U284 (N_284,In_615,In_657);
nor U285 (N_285,In_167,In_675);
nand U286 (N_286,In_373,In_648);
xnor U287 (N_287,In_419,In_7);
and U288 (N_288,In_398,In_58);
xor U289 (N_289,In_672,In_386);
and U290 (N_290,In_399,In_23);
xor U291 (N_291,In_97,In_84);
or U292 (N_292,In_599,In_651);
or U293 (N_293,In_53,In_525);
or U294 (N_294,In_706,In_484);
nand U295 (N_295,In_609,In_629);
and U296 (N_296,In_5,In_32);
and U297 (N_297,In_283,In_332);
or U298 (N_298,In_377,In_245);
xor U299 (N_299,In_728,In_393);
or U300 (N_300,In_704,In_147);
nand U301 (N_301,In_77,In_387);
or U302 (N_302,In_731,In_63);
nand U303 (N_303,In_206,In_22);
nor U304 (N_304,In_215,In_13);
nand U305 (N_305,In_623,In_636);
nor U306 (N_306,In_71,In_607);
or U307 (N_307,In_83,In_320);
and U308 (N_308,In_674,In_118);
or U309 (N_309,In_345,In_530);
xor U310 (N_310,In_85,In_605);
or U311 (N_311,In_404,In_532);
xnor U312 (N_312,In_658,In_91);
nor U313 (N_313,In_92,In_569);
xor U314 (N_314,In_690,In_133);
and U315 (N_315,In_559,In_87);
nand U316 (N_316,In_333,In_473);
or U317 (N_317,In_464,In_449);
or U318 (N_318,In_335,In_36);
nand U319 (N_319,In_693,In_407);
xnor U320 (N_320,In_611,In_230);
or U321 (N_321,In_128,In_243);
or U322 (N_322,In_140,In_199);
and U323 (N_323,In_135,In_740);
or U324 (N_324,In_369,In_16);
or U325 (N_325,In_201,In_437);
nand U326 (N_326,In_342,In_152);
and U327 (N_327,In_649,In_585);
xnor U328 (N_328,In_158,In_347);
and U329 (N_329,In_541,In_38);
nand U330 (N_330,In_504,In_197);
and U331 (N_331,In_631,In_222);
nor U332 (N_332,In_417,In_39);
xnor U333 (N_333,In_303,In_198);
nand U334 (N_334,In_626,In_620);
xnor U335 (N_335,In_37,In_540);
xnor U336 (N_336,In_365,In_272);
or U337 (N_337,In_93,In_219);
xor U338 (N_338,In_269,In_374);
nor U339 (N_339,In_277,In_228);
xnor U340 (N_340,In_59,In_471);
and U341 (N_341,In_506,In_563);
nand U342 (N_342,In_575,In_709);
or U343 (N_343,In_413,In_108);
nand U344 (N_344,In_736,In_454);
nand U345 (N_345,In_51,In_717);
nand U346 (N_346,In_324,In_512);
nand U347 (N_347,In_308,In_573);
and U348 (N_348,In_322,In_14);
nor U349 (N_349,In_70,In_161);
xnor U350 (N_350,In_749,In_251);
xnor U351 (N_351,In_593,In_526);
xnor U352 (N_352,In_163,In_35);
xor U353 (N_353,In_441,In_241);
xnor U354 (N_354,In_294,In_494);
nor U355 (N_355,In_395,In_490);
and U356 (N_356,In_659,In_17);
or U357 (N_357,In_475,In_290);
nand U358 (N_358,In_129,In_700);
and U359 (N_359,In_480,In_485);
and U360 (N_360,In_606,In_178);
nand U361 (N_361,In_154,In_500);
or U362 (N_362,In_448,In_720);
nor U363 (N_363,In_703,In_497);
and U364 (N_364,In_209,In_423);
xor U365 (N_365,In_301,In_558);
and U366 (N_366,In_62,In_246);
xor U367 (N_367,In_713,In_491);
or U368 (N_368,In_714,In_429);
nor U369 (N_369,In_295,In_12);
nand U370 (N_370,In_668,In_234);
nand U371 (N_371,In_537,In_551);
nand U372 (N_372,In_408,In_656);
xor U373 (N_373,In_48,In_641);
nand U374 (N_374,In_505,In_179);
nor U375 (N_375,In_262,In_158);
and U376 (N_376,In_129,In_532);
nor U377 (N_377,In_671,In_198);
or U378 (N_378,In_37,In_588);
and U379 (N_379,In_497,In_436);
nand U380 (N_380,In_90,In_570);
or U381 (N_381,In_671,In_56);
nand U382 (N_382,In_603,In_389);
xor U383 (N_383,In_478,In_686);
nor U384 (N_384,In_47,In_736);
and U385 (N_385,In_347,In_291);
nand U386 (N_386,In_143,In_49);
xnor U387 (N_387,In_343,In_221);
nand U388 (N_388,In_719,In_453);
nor U389 (N_389,In_565,In_653);
nand U390 (N_390,In_589,In_521);
nand U391 (N_391,In_400,In_302);
nand U392 (N_392,In_272,In_385);
nand U393 (N_393,In_188,In_544);
nand U394 (N_394,In_556,In_86);
nor U395 (N_395,In_389,In_725);
and U396 (N_396,In_677,In_16);
and U397 (N_397,In_279,In_292);
and U398 (N_398,In_92,In_383);
and U399 (N_399,In_623,In_69);
or U400 (N_400,In_399,In_552);
or U401 (N_401,In_368,In_690);
xnor U402 (N_402,In_609,In_362);
xnor U403 (N_403,In_423,In_119);
or U404 (N_404,In_543,In_305);
xnor U405 (N_405,In_311,In_235);
xnor U406 (N_406,In_33,In_350);
or U407 (N_407,In_745,In_134);
nand U408 (N_408,In_495,In_358);
and U409 (N_409,In_198,In_564);
nor U410 (N_410,In_238,In_245);
xnor U411 (N_411,In_327,In_385);
nand U412 (N_412,In_558,In_505);
nor U413 (N_413,In_387,In_68);
or U414 (N_414,In_656,In_256);
nand U415 (N_415,In_638,In_666);
nand U416 (N_416,In_109,In_511);
or U417 (N_417,In_140,In_487);
nand U418 (N_418,In_145,In_712);
xnor U419 (N_419,In_698,In_298);
or U420 (N_420,In_471,In_713);
or U421 (N_421,In_295,In_208);
or U422 (N_422,In_495,In_31);
nor U423 (N_423,In_17,In_609);
xor U424 (N_424,In_262,In_245);
nor U425 (N_425,In_529,In_127);
nor U426 (N_426,In_458,In_25);
nand U427 (N_427,In_648,In_238);
nor U428 (N_428,In_512,In_320);
xor U429 (N_429,In_697,In_38);
or U430 (N_430,In_86,In_308);
nand U431 (N_431,In_97,In_296);
and U432 (N_432,In_741,In_111);
xor U433 (N_433,In_302,In_231);
nand U434 (N_434,In_302,In_456);
nor U435 (N_435,In_298,In_608);
nor U436 (N_436,In_617,In_99);
and U437 (N_437,In_39,In_643);
nor U438 (N_438,In_493,In_14);
xnor U439 (N_439,In_78,In_515);
or U440 (N_440,In_739,In_643);
and U441 (N_441,In_556,In_571);
nand U442 (N_442,In_549,In_109);
nor U443 (N_443,In_407,In_438);
and U444 (N_444,In_286,In_38);
nand U445 (N_445,In_216,In_30);
nand U446 (N_446,In_666,In_563);
nor U447 (N_447,In_68,In_39);
nand U448 (N_448,In_278,In_244);
or U449 (N_449,In_9,In_596);
xnor U450 (N_450,In_245,In_488);
nor U451 (N_451,In_119,In_89);
nand U452 (N_452,In_137,In_77);
and U453 (N_453,In_608,In_632);
nand U454 (N_454,In_491,In_692);
nand U455 (N_455,In_176,In_227);
xor U456 (N_456,In_494,In_423);
xor U457 (N_457,In_100,In_322);
or U458 (N_458,In_526,In_82);
or U459 (N_459,In_100,In_635);
xor U460 (N_460,In_1,In_89);
or U461 (N_461,In_135,In_576);
and U462 (N_462,In_601,In_671);
or U463 (N_463,In_743,In_194);
xor U464 (N_464,In_142,In_710);
nor U465 (N_465,In_510,In_423);
nand U466 (N_466,In_247,In_674);
nand U467 (N_467,In_104,In_660);
or U468 (N_468,In_81,In_552);
or U469 (N_469,In_113,In_553);
and U470 (N_470,In_550,In_707);
or U471 (N_471,In_533,In_156);
nor U472 (N_472,In_69,In_11);
nor U473 (N_473,In_429,In_600);
xor U474 (N_474,In_30,In_232);
xnor U475 (N_475,In_482,In_425);
or U476 (N_476,In_718,In_396);
nand U477 (N_477,In_391,In_627);
or U478 (N_478,In_742,In_448);
nand U479 (N_479,In_488,In_146);
or U480 (N_480,In_495,In_450);
and U481 (N_481,In_121,In_636);
or U482 (N_482,In_108,In_161);
or U483 (N_483,In_194,In_472);
nand U484 (N_484,In_711,In_267);
nand U485 (N_485,In_518,In_313);
or U486 (N_486,In_167,In_155);
xor U487 (N_487,In_588,In_417);
or U488 (N_488,In_256,In_308);
nor U489 (N_489,In_588,In_603);
and U490 (N_490,In_197,In_355);
and U491 (N_491,In_271,In_39);
or U492 (N_492,In_440,In_676);
nor U493 (N_493,In_325,In_145);
nor U494 (N_494,In_601,In_49);
nand U495 (N_495,In_391,In_226);
nand U496 (N_496,In_664,In_20);
and U497 (N_497,In_561,In_547);
nor U498 (N_498,In_453,In_38);
and U499 (N_499,In_589,In_716);
nor U500 (N_500,N_265,N_398);
nand U501 (N_501,N_197,N_468);
xnor U502 (N_502,N_452,N_276);
and U503 (N_503,N_469,N_185);
or U504 (N_504,N_454,N_117);
or U505 (N_505,N_3,N_129);
nor U506 (N_506,N_303,N_4);
nand U507 (N_507,N_397,N_472);
nor U508 (N_508,N_278,N_118);
or U509 (N_509,N_460,N_222);
and U510 (N_510,N_194,N_270);
xor U511 (N_511,N_416,N_139);
or U512 (N_512,N_19,N_333);
and U513 (N_513,N_215,N_138);
and U514 (N_514,N_28,N_45);
and U515 (N_515,N_464,N_203);
or U516 (N_516,N_24,N_143);
and U517 (N_517,N_196,N_286);
xor U518 (N_518,N_463,N_66);
nor U519 (N_519,N_142,N_137);
and U520 (N_520,N_425,N_51);
nand U521 (N_521,N_144,N_281);
and U522 (N_522,N_422,N_1);
nor U523 (N_523,N_36,N_106);
or U524 (N_524,N_23,N_288);
nor U525 (N_525,N_348,N_52);
and U526 (N_526,N_101,N_392);
nor U527 (N_527,N_308,N_32);
or U528 (N_528,N_345,N_419);
and U529 (N_529,N_189,N_79);
and U530 (N_530,N_309,N_349);
or U531 (N_531,N_456,N_293);
xor U532 (N_532,N_104,N_376);
xnor U533 (N_533,N_103,N_93);
or U534 (N_534,N_251,N_156);
nor U535 (N_535,N_123,N_181);
xnor U536 (N_536,N_177,N_121);
xor U537 (N_537,N_290,N_410);
nand U538 (N_538,N_444,N_41);
xor U539 (N_539,N_87,N_62);
nor U540 (N_540,N_16,N_375);
xor U541 (N_541,N_343,N_307);
nor U542 (N_542,N_379,N_148);
nor U543 (N_543,N_353,N_497);
nand U544 (N_544,N_372,N_494);
nand U545 (N_545,N_172,N_279);
xor U546 (N_546,N_88,N_12);
nand U547 (N_547,N_268,N_300);
nor U548 (N_548,N_94,N_256);
nand U549 (N_549,N_183,N_433);
and U550 (N_550,N_112,N_130);
nand U551 (N_551,N_83,N_297);
xor U552 (N_552,N_26,N_445);
nor U553 (N_553,N_160,N_254);
xnor U554 (N_554,N_374,N_91);
xnor U555 (N_555,N_430,N_167);
xnor U556 (N_556,N_9,N_132);
or U557 (N_557,N_176,N_280);
nand U558 (N_558,N_33,N_367);
nand U559 (N_559,N_184,N_111);
nor U560 (N_560,N_260,N_342);
or U561 (N_561,N_25,N_340);
or U562 (N_562,N_64,N_10);
nor U563 (N_563,N_18,N_377);
nor U564 (N_564,N_238,N_237);
nor U565 (N_565,N_467,N_304);
or U566 (N_566,N_223,N_243);
nor U567 (N_567,N_490,N_318);
xor U568 (N_568,N_434,N_331);
or U569 (N_569,N_451,N_406);
or U570 (N_570,N_492,N_362);
nand U571 (N_571,N_169,N_344);
nand U572 (N_572,N_180,N_136);
nand U573 (N_573,N_283,N_306);
nor U574 (N_574,N_54,N_97);
and U575 (N_575,N_385,N_7);
xnor U576 (N_576,N_102,N_53);
nor U577 (N_577,N_248,N_43);
and U578 (N_578,N_115,N_39);
and U579 (N_579,N_21,N_239);
nor U580 (N_580,N_387,N_128);
nor U581 (N_581,N_170,N_273);
nand U582 (N_582,N_216,N_72);
and U583 (N_583,N_373,N_178);
nand U584 (N_584,N_386,N_50);
or U585 (N_585,N_393,N_69);
nor U586 (N_586,N_499,N_455);
nand U587 (N_587,N_27,N_346);
nand U588 (N_588,N_296,N_70);
or U589 (N_589,N_328,N_208);
xor U590 (N_590,N_125,N_31);
or U591 (N_591,N_165,N_120);
nor U592 (N_592,N_107,N_2);
nand U593 (N_593,N_299,N_321);
and U594 (N_594,N_229,N_60);
xor U595 (N_595,N_89,N_482);
xnor U596 (N_596,N_63,N_383);
or U597 (N_597,N_90,N_325);
nand U598 (N_598,N_449,N_480);
or U599 (N_599,N_439,N_193);
nand U600 (N_600,N_99,N_478);
xor U601 (N_601,N_302,N_242);
or U602 (N_602,N_412,N_214);
or U603 (N_603,N_166,N_359);
or U604 (N_604,N_399,N_48);
or U605 (N_605,N_76,N_105);
and U606 (N_606,N_319,N_457);
nand U607 (N_607,N_95,N_352);
or U608 (N_608,N_298,N_301);
xnor U609 (N_609,N_382,N_200);
nor U610 (N_610,N_465,N_252);
nand U611 (N_611,N_152,N_351);
and U612 (N_612,N_429,N_441);
and U613 (N_613,N_271,N_162);
nor U614 (N_614,N_59,N_255);
nor U615 (N_615,N_339,N_226);
or U616 (N_616,N_365,N_46);
or U617 (N_617,N_431,N_131);
nand U618 (N_618,N_247,N_258);
nand U619 (N_619,N_438,N_44);
nand U620 (N_620,N_71,N_440);
nand U621 (N_621,N_100,N_257);
xor U622 (N_622,N_462,N_448);
nor U623 (N_623,N_413,N_287);
and U624 (N_624,N_428,N_316);
nand U625 (N_625,N_47,N_8);
nand U626 (N_626,N_334,N_409);
nand U627 (N_627,N_487,N_175);
nand U628 (N_628,N_198,N_314);
nand U629 (N_629,N_157,N_404);
nand U630 (N_630,N_145,N_370);
nand U631 (N_631,N_199,N_380);
nand U632 (N_632,N_5,N_244);
nor U633 (N_633,N_371,N_220);
nand U634 (N_634,N_424,N_261);
nor U635 (N_635,N_496,N_42);
nand U636 (N_636,N_40,N_488);
and U637 (N_637,N_320,N_67);
and U638 (N_638,N_310,N_262);
nor U639 (N_639,N_473,N_423);
xnor U640 (N_640,N_498,N_411);
and U641 (N_641,N_161,N_394);
nor U642 (N_642,N_305,N_146);
nand U643 (N_643,N_0,N_86);
xor U644 (N_644,N_477,N_240);
nor U645 (N_645,N_135,N_447);
nor U646 (N_646,N_474,N_206);
or U647 (N_647,N_378,N_327);
xor U648 (N_648,N_360,N_329);
and U649 (N_649,N_389,N_55);
and U650 (N_650,N_401,N_159);
or U651 (N_651,N_446,N_92);
and U652 (N_652,N_154,N_493);
nor U653 (N_653,N_390,N_337);
or U654 (N_654,N_384,N_147);
nand U655 (N_655,N_292,N_210);
and U656 (N_656,N_263,N_364);
and U657 (N_657,N_275,N_6);
or U658 (N_658,N_61,N_204);
nand U659 (N_659,N_259,N_49);
xor U660 (N_660,N_332,N_173);
nand U661 (N_661,N_20,N_96);
nand U662 (N_662,N_232,N_437);
and U663 (N_663,N_124,N_479);
nor U664 (N_664,N_317,N_11);
xnor U665 (N_665,N_171,N_388);
nor U666 (N_666,N_495,N_218);
xnor U667 (N_667,N_489,N_151);
nor U668 (N_668,N_403,N_57);
nand U669 (N_669,N_35,N_289);
xnor U670 (N_670,N_164,N_187);
nand U671 (N_671,N_356,N_74);
or U672 (N_672,N_400,N_407);
xor U673 (N_673,N_98,N_75);
or U674 (N_674,N_357,N_153);
nand U675 (N_675,N_108,N_436);
xor U676 (N_676,N_217,N_420);
nor U677 (N_677,N_427,N_236);
nor U678 (N_678,N_368,N_418);
and U679 (N_679,N_81,N_491);
or U680 (N_680,N_470,N_213);
nor U681 (N_681,N_246,N_158);
and U682 (N_682,N_366,N_294);
and U683 (N_683,N_415,N_38);
xnor U684 (N_684,N_29,N_313);
and U685 (N_685,N_396,N_295);
or U686 (N_686,N_133,N_230);
and U687 (N_687,N_414,N_140);
nand U688 (N_688,N_73,N_341);
xor U689 (N_689,N_350,N_221);
nand U690 (N_690,N_234,N_127);
xnor U691 (N_691,N_188,N_483);
nor U692 (N_692,N_272,N_266);
xnor U693 (N_693,N_347,N_182);
xnor U694 (N_694,N_186,N_14);
or U695 (N_695,N_338,N_395);
or U696 (N_696,N_485,N_219);
xnor U697 (N_697,N_466,N_402);
nor U698 (N_698,N_65,N_381);
or U699 (N_699,N_282,N_227);
nand U700 (N_700,N_109,N_250);
nand U701 (N_701,N_163,N_450);
or U702 (N_702,N_458,N_225);
nor U703 (N_703,N_330,N_191);
and U704 (N_704,N_179,N_363);
nor U705 (N_705,N_476,N_56);
and U706 (N_706,N_155,N_228);
and U707 (N_707,N_274,N_355);
nand U708 (N_708,N_209,N_17);
or U709 (N_709,N_326,N_113);
nand U710 (N_710,N_249,N_82);
nand U711 (N_711,N_231,N_78);
or U712 (N_712,N_174,N_354);
nand U713 (N_713,N_212,N_122);
or U714 (N_714,N_168,N_235);
xnor U715 (N_715,N_421,N_335);
or U716 (N_716,N_211,N_37);
or U717 (N_717,N_13,N_202);
or U718 (N_718,N_34,N_481);
nand U719 (N_719,N_312,N_442);
nor U720 (N_720,N_241,N_322);
and U721 (N_721,N_150,N_417);
or U722 (N_722,N_195,N_58);
nor U723 (N_723,N_201,N_432);
and U724 (N_724,N_471,N_114);
and U725 (N_725,N_84,N_110);
nand U726 (N_726,N_284,N_192);
and U727 (N_727,N_119,N_461);
or U728 (N_728,N_369,N_267);
nor U729 (N_729,N_224,N_205);
nor U730 (N_730,N_134,N_391);
and U731 (N_731,N_324,N_116);
or U732 (N_732,N_435,N_149);
nor U733 (N_733,N_264,N_77);
nand U734 (N_734,N_22,N_285);
or U735 (N_735,N_336,N_459);
nand U736 (N_736,N_207,N_141);
nand U737 (N_737,N_291,N_15);
xnor U738 (N_738,N_405,N_85);
and U739 (N_739,N_361,N_311);
xor U740 (N_740,N_253,N_408);
nor U741 (N_741,N_233,N_453);
and U742 (N_742,N_426,N_484);
xnor U743 (N_743,N_30,N_486);
or U744 (N_744,N_68,N_277);
xnor U745 (N_745,N_269,N_475);
or U746 (N_746,N_126,N_80);
or U747 (N_747,N_315,N_358);
nor U748 (N_748,N_245,N_190);
or U749 (N_749,N_323,N_443);
xnor U750 (N_750,N_201,N_212);
xnor U751 (N_751,N_377,N_301);
nor U752 (N_752,N_346,N_347);
and U753 (N_753,N_437,N_260);
xnor U754 (N_754,N_29,N_143);
xnor U755 (N_755,N_450,N_214);
nand U756 (N_756,N_138,N_362);
nor U757 (N_757,N_64,N_12);
xor U758 (N_758,N_58,N_483);
and U759 (N_759,N_456,N_115);
or U760 (N_760,N_490,N_438);
xor U761 (N_761,N_391,N_403);
xnor U762 (N_762,N_375,N_302);
or U763 (N_763,N_279,N_248);
and U764 (N_764,N_108,N_280);
nor U765 (N_765,N_245,N_244);
and U766 (N_766,N_185,N_10);
nor U767 (N_767,N_318,N_206);
or U768 (N_768,N_58,N_427);
and U769 (N_769,N_348,N_401);
and U770 (N_770,N_196,N_362);
nor U771 (N_771,N_272,N_214);
nor U772 (N_772,N_254,N_409);
or U773 (N_773,N_486,N_394);
and U774 (N_774,N_108,N_190);
and U775 (N_775,N_277,N_409);
nor U776 (N_776,N_403,N_378);
and U777 (N_777,N_264,N_418);
nor U778 (N_778,N_359,N_177);
or U779 (N_779,N_89,N_497);
nand U780 (N_780,N_423,N_239);
or U781 (N_781,N_110,N_213);
and U782 (N_782,N_399,N_417);
xor U783 (N_783,N_116,N_132);
or U784 (N_784,N_53,N_312);
nand U785 (N_785,N_93,N_198);
and U786 (N_786,N_92,N_154);
xor U787 (N_787,N_462,N_323);
xnor U788 (N_788,N_181,N_24);
nor U789 (N_789,N_462,N_5);
xor U790 (N_790,N_415,N_167);
xor U791 (N_791,N_467,N_261);
and U792 (N_792,N_486,N_445);
or U793 (N_793,N_95,N_428);
or U794 (N_794,N_412,N_262);
nand U795 (N_795,N_52,N_459);
or U796 (N_796,N_30,N_475);
nor U797 (N_797,N_304,N_379);
or U798 (N_798,N_238,N_307);
or U799 (N_799,N_89,N_309);
xor U800 (N_800,N_364,N_351);
nor U801 (N_801,N_468,N_232);
xnor U802 (N_802,N_52,N_111);
or U803 (N_803,N_127,N_360);
or U804 (N_804,N_82,N_386);
and U805 (N_805,N_226,N_206);
nor U806 (N_806,N_73,N_381);
nor U807 (N_807,N_3,N_120);
nand U808 (N_808,N_93,N_319);
or U809 (N_809,N_449,N_335);
and U810 (N_810,N_200,N_20);
nand U811 (N_811,N_120,N_178);
nand U812 (N_812,N_10,N_343);
or U813 (N_813,N_394,N_422);
nor U814 (N_814,N_421,N_247);
or U815 (N_815,N_27,N_6);
xor U816 (N_816,N_427,N_100);
nor U817 (N_817,N_463,N_472);
and U818 (N_818,N_438,N_388);
nand U819 (N_819,N_118,N_16);
nor U820 (N_820,N_324,N_253);
xnor U821 (N_821,N_33,N_336);
xnor U822 (N_822,N_308,N_49);
xor U823 (N_823,N_434,N_416);
nand U824 (N_824,N_477,N_281);
nor U825 (N_825,N_234,N_299);
or U826 (N_826,N_148,N_425);
nand U827 (N_827,N_483,N_270);
nand U828 (N_828,N_463,N_94);
xnor U829 (N_829,N_4,N_243);
nor U830 (N_830,N_23,N_363);
nor U831 (N_831,N_267,N_496);
nand U832 (N_832,N_131,N_443);
xnor U833 (N_833,N_296,N_293);
and U834 (N_834,N_52,N_258);
nand U835 (N_835,N_100,N_487);
and U836 (N_836,N_116,N_398);
xor U837 (N_837,N_374,N_495);
or U838 (N_838,N_472,N_320);
xnor U839 (N_839,N_305,N_28);
xnor U840 (N_840,N_367,N_245);
or U841 (N_841,N_219,N_211);
and U842 (N_842,N_277,N_472);
or U843 (N_843,N_466,N_178);
xor U844 (N_844,N_301,N_463);
or U845 (N_845,N_188,N_279);
or U846 (N_846,N_10,N_108);
xor U847 (N_847,N_166,N_27);
or U848 (N_848,N_163,N_358);
or U849 (N_849,N_39,N_418);
and U850 (N_850,N_176,N_258);
and U851 (N_851,N_92,N_177);
nand U852 (N_852,N_270,N_29);
nand U853 (N_853,N_64,N_257);
or U854 (N_854,N_422,N_107);
nor U855 (N_855,N_239,N_19);
xnor U856 (N_856,N_496,N_264);
xnor U857 (N_857,N_83,N_435);
xor U858 (N_858,N_34,N_218);
nor U859 (N_859,N_198,N_125);
xnor U860 (N_860,N_118,N_372);
nand U861 (N_861,N_441,N_321);
nand U862 (N_862,N_227,N_361);
or U863 (N_863,N_238,N_58);
nand U864 (N_864,N_75,N_372);
nor U865 (N_865,N_222,N_407);
nand U866 (N_866,N_82,N_163);
nand U867 (N_867,N_235,N_110);
xnor U868 (N_868,N_322,N_268);
or U869 (N_869,N_403,N_275);
and U870 (N_870,N_120,N_33);
nor U871 (N_871,N_54,N_299);
nor U872 (N_872,N_381,N_456);
nor U873 (N_873,N_260,N_411);
nor U874 (N_874,N_424,N_351);
nor U875 (N_875,N_32,N_102);
or U876 (N_876,N_129,N_124);
or U877 (N_877,N_25,N_252);
nand U878 (N_878,N_415,N_366);
or U879 (N_879,N_467,N_125);
and U880 (N_880,N_478,N_180);
nor U881 (N_881,N_457,N_93);
nor U882 (N_882,N_389,N_134);
or U883 (N_883,N_414,N_130);
nor U884 (N_884,N_280,N_486);
and U885 (N_885,N_344,N_413);
or U886 (N_886,N_245,N_427);
or U887 (N_887,N_71,N_9);
nor U888 (N_888,N_474,N_138);
nor U889 (N_889,N_342,N_20);
or U890 (N_890,N_371,N_152);
and U891 (N_891,N_498,N_1);
nand U892 (N_892,N_483,N_277);
xnor U893 (N_893,N_262,N_445);
and U894 (N_894,N_377,N_290);
nand U895 (N_895,N_399,N_174);
and U896 (N_896,N_390,N_121);
and U897 (N_897,N_130,N_464);
xor U898 (N_898,N_284,N_342);
nor U899 (N_899,N_310,N_352);
and U900 (N_900,N_412,N_80);
or U901 (N_901,N_481,N_288);
nand U902 (N_902,N_165,N_41);
nor U903 (N_903,N_493,N_257);
xnor U904 (N_904,N_321,N_132);
xor U905 (N_905,N_194,N_366);
nand U906 (N_906,N_268,N_354);
xnor U907 (N_907,N_318,N_368);
and U908 (N_908,N_382,N_302);
nand U909 (N_909,N_100,N_324);
and U910 (N_910,N_366,N_119);
nand U911 (N_911,N_326,N_118);
and U912 (N_912,N_233,N_146);
nand U913 (N_913,N_471,N_279);
and U914 (N_914,N_351,N_444);
and U915 (N_915,N_373,N_452);
nor U916 (N_916,N_272,N_244);
xor U917 (N_917,N_331,N_431);
nor U918 (N_918,N_210,N_267);
nand U919 (N_919,N_143,N_2);
xnor U920 (N_920,N_193,N_105);
or U921 (N_921,N_174,N_377);
xor U922 (N_922,N_246,N_494);
nor U923 (N_923,N_276,N_218);
nor U924 (N_924,N_317,N_33);
nand U925 (N_925,N_383,N_488);
or U926 (N_926,N_241,N_191);
xnor U927 (N_927,N_354,N_315);
and U928 (N_928,N_437,N_321);
nor U929 (N_929,N_79,N_296);
xor U930 (N_930,N_244,N_443);
and U931 (N_931,N_397,N_284);
nor U932 (N_932,N_398,N_453);
xnor U933 (N_933,N_1,N_291);
nor U934 (N_934,N_95,N_196);
nor U935 (N_935,N_143,N_393);
or U936 (N_936,N_230,N_56);
and U937 (N_937,N_196,N_42);
xnor U938 (N_938,N_63,N_486);
xor U939 (N_939,N_357,N_229);
or U940 (N_940,N_59,N_129);
and U941 (N_941,N_348,N_32);
nand U942 (N_942,N_170,N_60);
nand U943 (N_943,N_151,N_325);
nand U944 (N_944,N_115,N_339);
xor U945 (N_945,N_174,N_473);
nor U946 (N_946,N_467,N_460);
nor U947 (N_947,N_358,N_156);
nand U948 (N_948,N_222,N_328);
nor U949 (N_949,N_143,N_162);
or U950 (N_950,N_425,N_253);
or U951 (N_951,N_410,N_221);
xor U952 (N_952,N_166,N_177);
nor U953 (N_953,N_39,N_3);
nor U954 (N_954,N_226,N_94);
nand U955 (N_955,N_392,N_301);
nand U956 (N_956,N_127,N_482);
nor U957 (N_957,N_37,N_494);
and U958 (N_958,N_422,N_363);
xor U959 (N_959,N_239,N_272);
xnor U960 (N_960,N_216,N_349);
and U961 (N_961,N_102,N_26);
or U962 (N_962,N_474,N_384);
nand U963 (N_963,N_66,N_384);
nand U964 (N_964,N_422,N_455);
nand U965 (N_965,N_9,N_415);
or U966 (N_966,N_42,N_293);
or U967 (N_967,N_299,N_172);
and U968 (N_968,N_354,N_355);
nand U969 (N_969,N_389,N_119);
and U970 (N_970,N_196,N_493);
nand U971 (N_971,N_233,N_183);
and U972 (N_972,N_220,N_496);
and U973 (N_973,N_329,N_335);
and U974 (N_974,N_320,N_25);
or U975 (N_975,N_182,N_107);
or U976 (N_976,N_247,N_182);
xnor U977 (N_977,N_102,N_264);
nor U978 (N_978,N_193,N_360);
or U979 (N_979,N_311,N_156);
xor U980 (N_980,N_353,N_319);
and U981 (N_981,N_407,N_403);
and U982 (N_982,N_120,N_1);
or U983 (N_983,N_61,N_390);
nand U984 (N_984,N_304,N_167);
xnor U985 (N_985,N_468,N_68);
nand U986 (N_986,N_24,N_275);
or U987 (N_987,N_71,N_35);
xnor U988 (N_988,N_318,N_319);
or U989 (N_989,N_305,N_338);
xor U990 (N_990,N_401,N_121);
nand U991 (N_991,N_385,N_448);
nand U992 (N_992,N_383,N_260);
xnor U993 (N_993,N_0,N_484);
xor U994 (N_994,N_395,N_92);
xnor U995 (N_995,N_78,N_5);
and U996 (N_996,N_94,N_12);
nand U997 (N_997,N_491,N_497);
xor U998 (N_998,N_295,N_190);
nor U999 (N_999,N_455,N_103);
nor U1000 (N_1000,N_992,N_942);
nand U1001 (N_1001,N_761,N_855);
or U1002 (N_1002,N_511,N_729);
nor U1003 (N_1003,N_829,N_704);
or U1004 (N_1004,N_584,N_932);
xor U1005 (N_1005,N_927,N_644);
nor U1006 (N_1006,N_772,N_899);
nor U1007 (N_1007,N_647,N_801);
xor U1008 (N_1008,N_719,N_579);
or U1009 (N_1009,N_720,N_672);
nor U1010 (N_1010,N_773,N_828);
xor U1011 (N_1011,N_895,N_521);
and U1012 (N_1012,N_503,N_770);
or U1013 (N_1013,N_702,N_824);
nand U1014 (N_1014,N_649,N_776);
nand U1015 (N_1015,N_707,N_838);
nand U1016 (N_1016,N_938,N_826);
nor U1017 (N_1017,N_953,N_916);
nand U1018 (N_1018,N_697,N_808);
and U1019 (N_1019,N_542,N_532);
and U1020 (N_1020,N_984,N_562);
xnor U1021 (N_1021,N_576,N_687);
nor U1022 (N_1022,N_849,N_548);
xnor U1023 (N_1023,N_705,N_936);
and U1024 (N_1024,N_993,N_965);
or U1025 (N_1025,N_689,N_980);
xnor U1026 (N_1026,N_646,N_901);
xor U1027 (N_1027,N_739,N_893);
or U1028 (N_1028,N_727,N_818);
or U1029 (N_1029,N_636,N_890);
and U1030 (N_1030,N_615,N_527);
and U1031 (N_1031,N_660,N_678);
xnor U1032 (N_1032,N_786,N_915);
xnor U1033 (N_1033,N_625,N_754);
nand U1034 (N_1034,N_810,N_574);
nor U1035 (N_1035,N_888,N_635);
nand U1036 (N_1036,N_785,N_633);
xor U1037 (N_1037,N_950,N_605);
and U1038 (N_1038,N_716,N_612);
xor U1039 (N_1039,N_934,N_544);
nor U1040 (N_1040,N_821,N_944);
or U1041 (N_1041,N_983,N_587);
and U1042 (N_1042,N_835,N_945);
and U1043 (N_1043,N_990,N_847);
or U1044 (N_1044,N_525,N_782);
and U1045 (N_1045,N_561,N_709);
and U1046 (N_1046,N_536,N_787);
or U1047 (N_1047,N_811,N_679);
nand U1048 (N_1048,N_820,N_753);
xor U1049 (N_1049,N_706,N_898);
and U1050 (N_1050,N_564,N_806);
xor U1051 (N_1051,N_630,N_836);
xor U1052 (N_1052,N_962,N_930);
nand U1053 (N_1053,N_712,N_710);
nor U1054 (N_1054,N_780,N_750);
nand U1055 (N_1055,N_749,N_926);
nand U1056 (N_1056,N_796,N_839);
nand U1057 (N_1057,N_831,N_653);
or U1058 (N_1058,N_571,N_853);
nand U1059 (N_1059,N_834,N_575);
and U1060 (N_1060,N_919,N_569);
and U1061 (N_1061,N_762,N_734);
xor U1062 (N_1062,N_779,N_863);
nor U1063 (N_1063,N_568,N_694);
nand U1064 (N_1064,N_682,N_833);
or U1065 (N_1065,N_939,N_940);
or U1066 (N_1066,N_583,N_790);
and U1067 (N_1067,N_658,N_931);
xnor U1068 (N_1068,N_555,N_803);
or U1069 (N_1069,N_947,N_840);
nor U1070 (N_1070,N_974,N_692);
and U1071 (N_1071,N_590,N_952);
and U1072 (N_1072,N_850,N_872);
and U1073 (N_1073,N_703,N_557);
and U1074 (N_1074,N_873,N_613);
nor U1075 (N_1075,N_763,N_908);
nor U1076 (N_1076,N_910,N_815);
nand U1077 (N_1077,N_791,N_539);
and U1078 (N_1078,N_771,N_713);
and U1079 (N_1079,N_522,N_929);
nor U1080 (N_1080,N_628,N_812);
and U1081 (N_1081,N_784,N_591);
or U1082 (N_1082,N_664,N_669);
nand U1083 (N_1083,N_900,N_600);
nor U1084 (N_1084,N_606,N_604);
xor U1085 (N_1085,N_886,N_907);
nor U1086 (N_1086,N_830,N_518);
nand U1087 (N_1087,N_912,N_502);
and U1088 (N_1088,N_645,N_816);
or U1089 (N_1089,N_756,N_875);
or U1090 (N_1090,N_923,N_500);
or U1091 (N_1091,N_730,N_566);
xnor U1092 (N_1092,N_814,N_534);
and U1093 (N_1093,N_982,N_744);
xnor U1094 (N_1094,N_686,N_832);
xnor U1095 (N_1095,N_519,N_883);
xor U1096 (N_1096,N_827,N_925);
nand U1097 (N_1097,N_954,N_531);
nor U1098 (N_1098,N_523,N_918);
xnor U1099 (N_1099,N_922,N_556);
or U1100 (N_1100,N_989,N_960);
and U1101 (N_1101,N_999,N_701);
and U1102 (N_1102,N_994,N_991);
xnor U1103 (N_1103,N_524,N_733);
xnor U1104 (N_1104,N_597,N_700);
and U1105 (N_1105,N_673,N_928);
nor U1106 (N_1106,N_963,N_608);
xor U1107 (N_1107,N_603,N_639);
nand U1108 (N_1108,N_775,N_741);
or U1109 (N_1109,N_668,N_560);
and U1110 (N_1110,N_842,N_933);
nor U1111 (N_1111,N_743,N_843);
nor U1112 (N_1112,N_817,N_854);
or U1113 (N_1113,N_959,N_663);
nor U1114 (N_1114,N_602,N_513);
or U1115 (N_1115,N_624,N_765);
nor U1116 (N_1116,N_659,N_794);
or U1117 (N_1117,N_971,N_799);
or U1118 (N_1118,N_535,N_985);
nor U1119 (N_1119,N_805,N_565);
or U1120 (N_1120,N_902,N_997);
and U1121 (N_1121,N_671,N_640);
or U1122 (N_1122,N_558,N_552);
xnor U1123 (N_1123,N_758,N_593);
nand U1124 (N_1124,N_903,N_723);
or U1125 (N_1125,N_792,N_973);
or U1126 (N_1126,N_680,N_577);
nand U1127 (N_1127,N_751,N_642);
nand U1128 (N_1128,N_882,N_964);
nand U1129 (N_1129,N_553,N_949);
or U1130 (N_1130,N_891,N_870);
nor U1131 (N_1131,N_594,N_654);
nor U1132 (N_1132,N_512,N_622);
xor U1133 (N_1133,N_978,N_547);
nand U1134 (N_1134,N_881,N_567);
xor U1135 (N_1135,N_778,N_693);
nor U1136 (N_1136,N_724,N_504);
xor U1137 (N_1137,N_586,N_867);
or U1138 (N_1138,N_698,N_788);
nor U1139 (N_1139,N_641,N_906);
and U1140 (N_1140,N_943,N_551);
nor U1141 (N_1141,N_937,N_638);
and U1142 (N_1142,N_742,N_626);
xor U1143 (N_1143,N_967,N_804);
xnor U1144 (N_1144,N_607,N_725);
nand U1145 (N_1145,N_755,N_696);
nand U1146 (N_1146,N_616,N_589);
or U1147 (N_1147,N_914,N_958);
and U1148 (N_1148,N_533,N_685);
nand U1149 (N_1149,N_987,N_889);
nand U1150 (N_1150,N_695,N_789);
nand U1151 (N_1151,N_530,N_510);
nor U1152 (N_1152,N_921,N_852);
nor U1153 (N_1153,N_924,N_878);
nor U1154 (N_1154,N_955,N_514);
or U1155 (N_1155,N_515,N_740);
and U1156 (N_1156,N_667,N_800);
or U1157 (N_1157,N_599,N_688);
and U1158 (N_1158,N_718,N_897);
and U1159 (N_1159,N_573,N_880);
and U1160 (N_1160,N_920,N_858);
and U1161 (N_1161,N_581,N_837);
and U1162 (N_1162,N_904,N_714);
xor U1163 (N_1163,N_736,N_545);
xor U1164 (N_1164,N_563,N_621);
xor U1165 (N_1165,N_506,N_728);
nand U1166 (N_1166,N_651,N_774);
xnor U1167 (N_1167,N_913,N_598);
nor U1168 (N_1168,N_911,N_711);
nand U1169 (N_1169,N_861,N_722);
nand U1170 (N_1170,N_674,N_631);
xor U1171 (N_1171,N_885,N_505);
xnor U1172 (N_1172,N_726,N_662);
nor U1173 (N_1173,N_968,N_988);
and U1174 (N_1174,N_632,N_857);
nand U1175 (N_1175,N_619,N_732);
nand U1176 (N_1176,N_528,N_699);
or U1177 (N_1177,N_580,N_737);
nand U1178 (N_1178,N_819,N_760);
or U1179 (N_1179,N_892,N_846);
xor U1180 (N_1180,N_844,N_623);
xnor U1181 (N_1181,N_657,N_559);
xnor U1182 (N_1182,N_767,N_975);
or U1183 (N_1183,N_549,N_572);
or U1184 (N_1184,N_609,N_961);
nand U1185 (N_1185,N_887,N_841);
nand U1186 (N_1186,N_865,N_884);
xor U1187 (N_1187,N_856,N_781);
xnor U1188 (N_1188,N_793,N_614);
or U1189 (N_1189,N_848,N_777);
and U1190 (N_1190,N_981,N_879);
nor U1191 (N_1191,N_909,N_894);
and U1192 (N_1192,N_748,N_617);
nor U1193 (N_1193,N_996,N_526);
or U1194 (N_1194,N_611,N_905);
nand U1195 (N_1195,N_618,N_634);
and U1196 (N_1196,N_768,N_543);
or U1197 (N_1197,N_860,N_643);
and U1198 (N_1198,N_627,N_620);
or U1199 (N_1199,N_676,N_582);
xnor U1200 (N_1200,N_979,N_665);
nand U1201 (N_1201,N_546,N_969);
nand U1202 (N_1202,N_721,N_666);
or U1203 (N_1203,N_601,N_508);
or U1204 (N_1204,N_917,N_956);
nand U1205 (N_1205,N_862,N_976);
xnor U1206 (N_1206,N_869,N_995);
or U1207 (N_1207,N_585,N_681);
and U1208 (N_1208,N_570,N_998);
and U1209 (N_1209,N_655,N_675);
xor U1210 (N_1210,N_825,N_731);
nor U1211 (N_1211,N_896,N_691);
and U1212 (N_1212,N_948,N_823);
and U1213 (N_1213,N_592,N_529);
nand U1214 (N_1214,N_690,N_684);
nor U1215 (N_1215,N_550,N_520);
and U1216 (N_1216,N_876,N_798);
and U1217 (N_1217,N_874,N_868);
xnor U1218 (N_1218,N_822,N_966);
and U1219 (N_1219,N_516,N_517);
and U1220 (N_1220,N_759,N_871);
nor U1221 (N_1221,N_629,N_807);
and U1222 (N_1222,N_851,N_745);
nor U1223 (N_1223,N_951,N_554);
nor U1224 (N_1224,N_845,N_610);
nand U1225 (N_1225,N_738,N_802);
or U1226 (N_1226,N_507,N_977);
and U1227 (N_1227,N_970,N_764);
or U1228 (N_1228,N_595,N_795);
nor U1229 (N_1229,N_708,N_783);
and U1230 (N_1230,N_661,N_957);
nand U1231 (N_1231,N_747,N_866);
or U1232 (N_1232,N_652,N_650);
or U1233 (N_1233,N_746,N_648);
or U1234 (N_1234,N_578,N_813);
nand U1235 (N_1235,N_972,N_797);
nor U1236 (N_1236,N_683,N_859);
xnor U1237 (N_1237,N_946,N_715);
and U1238 (N_1238,N_540,N_538);
xor U1239 (N_1239,N_757,N_717);
xnor U1240 (N_1240,N_509,N_752);
nor U1241 (N_1241,N_864,N_809);
and U1242 (N_1242,N_596,N_541);
nand U1243 (N_1243,N_877,N_637);
and U1244 (N_1244,N_766,N_986);
or U1245 (N_1245,N_670,N_656);
nand U1246 (N_1246,N_537,N_677);
nor U1247 (N_1247,N_501,N_588);
nand U1248 (N_1248,N_735,N_941);
or U1249 (N_1249,N_935,N_769);
and U1250 (N_1250,N_991,N_864);
nand U1251 (N_1251,N_905,N_908);
or U1252 (N_1252,N_790,N_910);
nand U1253 (N_1253,N_709,N_525);
nand U1254 (N_1254,N_947,N_885);
xor U1255 (N_1255,N_808,N_554);
nor U1256 (N_1256,N_867,N_601);
nand U1257 (N_1257,N_757,N_769);
nand U1258 (N_1258,N_571,N_524);
nand U1259 (N_1259,N_964,N_937);
nand U1260 (N_1260,N_912,N_789);
xnor U1261 (N_1261,N_719,N_661);
or U1262 (N_1262,N_730,N_661);
nor U1263 (N_1263,N_790,N_538);
or U1264 (N_1264,N_511,N_926);
nand U1265 (N_1265,N_582,N_570);
or U1266 (N_1266,N_741,N_736);
nand U1267 (N_1267,N_551,N_663);
xor U1268 (N_1268,N_572,N_995);
and U1269 (N_1269,N_908,N_805);
and U1270 (N_1270,N_747,N_676);
xnor U1271 (N_1271,N_613,N_537);
or U1272 (N_1272,N_771,N_961);
and U1273 (N_1273,N_587,N_669);
or U1274 (N_1274,N_814,N_896);
xor U1275 (N_1275,N_797,N_593);
and U1276 (N_1276,N_991,N_953);
nor U1277 (N_1277,N_770,N_706);
nand U1278 (N_1278,N_829,N_682);
xnor U1279 (N_1279,N_996,N_568);
xnor U1280 (N_1280,N_716,N_919);
nand U1281 (N_1281,N_997,N_852);
or U1282 (N_1282,N_714,N_836);
nand U1283 (N_1283,N_772,N_698);
nand U1284 (N_1284,N_980,N_766);
and U1285 (N_1285,N_886,N_667);
nor U1286 (N_1286,N_634,N_855);
or U1287 (N_1287,N_907,N_810);
xor U1288 (N_1288,N_832,N_773);
nand U1289 (N_1289,N_980,N_782);
xnor U1290 (N_1290,N_627,N_754);
nand U1291 (N_1291,N_927,N_524);
and U1292 (N_1292,N_982,N_996);
or U1293 (N_1293,N_902,N_666);
nor U1294 (N_1294,N_666,N_873);
nor U1295 (N_1295,N_718,N_992);
or U1296 (N_1296,N_975,N_937);
nor U1297 (N_1297,N_630,N_546);
or U1298 (N_1298,N_553,N_808);
or U1299 (N_1299,N_697,N_645);
and U1300 (N_1300,N_647,N_803);
or U1301 (N_1301,N_842,N_521);
xnor U1302 (N_1302,N_965,N_520);
xnor U1303 (N_1303,N_644,N_830);
and U1304 (N_1304,N_778,N_723);
nand U1305 (N_1305,N_983,N_579);
nand U1306 (N_1306,N_639,N_546);
xnor U1307 (N_1307,N_950,N_775);
and U1308 (N_1308,N_511,N_887);
and U1309 (N_1309,N_875,N_603);
nand U1310 (N_1310,N_868,N_886);
xor U1311 (N_1311,N_999,N_523);
nand U1312 (N_1312,N_610,N_735);
and U1313 (N_1313,N_984,N_675);
and U1314 (N_1314,N_576,N_742);
and U1315 (N_1315,N_679,N_629);
nor U1316 (N_1316,N_992,N_609);
nor U1317 (N_1317,N_518,N_929);
nand U1318 (N_1318,N_654,N_834);
or U1319 (N_1319,N_553,N_965);
or U1320 (N_1320,N_799,N_921);
nor U1321 (N_1321,N_514,N_960);
and U1322 (N_1322,N_869,N_729);
or U1323 (N_1323,N_866,N_629);
nand U1324 (N_1324,N_737,N_693);
or U1325 (N_1325,N_604,N_719);
or U1326 (N_1326,N_987,N_514);
xnor U1327 (N_1327,N_900,N_653);
or U1328 (N_1328,N_739,N_774);
nand U1329 (N_1329,N_927,N_680);
or U1330 (N_1330,N_818,N_630);
xor U1331 (N_1331,N_982,N_514);
and U1332 (N_1332,N_781,N_615);
nand U1333 (N_1333,N_797,N_848);
nor U1334 (N_1334,N_703,N_529);
and U1335 (N_1335,N_563,N_732);
xor U1336 (N_1336,N_938,N_929);
nor U1337 (N_1337,N_784,N_532);
and U1338 (N_1338,N_786,N_912);
nand U1339 (N_1339,N_701,N_511);
and U1340 (N_1340,N_590,N_747);
nand U1341 (N_1341,N_930,N_552);
and U1342 (N_1342,N_689,N_756);
xor U1343 (N_1343,N_595,N_696);
nand U1344 (N_1344,N_587,N_819);
xnor U1345 (N_1345,N_510,N_586);
and U1346 (N_1346,N_837,N_734);
nand U1347 (N_1347,N_652,N_959);
nor U1348 (N_1348,N_967,N_983);
nand U1349 (N_1349,N_555,N_610);
or U1350 (N_1350,N_578,N_981);
and U1351 (N_1351,N_862,N_823);
and U1352 (N_1352,N_964,N_595);
nor U1353 (N_1353,N_876,N_701);
nand U1354 (N_1354,N_636,N_620);
xnor U1355 (N_1355,N_860,N_622);
or U1356 (N_1356,N_644,N_813);
and U1357 (N_1357,N_954,N_964);
or U1358 (N_1358,N_861,N_829);
nor U1359 (N_1359,N_606,N_868);
and U1360 (N_1360,N_560,N_935);
nor U1361 (N_1361,N_887,N_686);
or U1362 (N_1362,N_790,N_811);
nor U1363 (N_1363,N_614,N_607);
xor U1364 (N_1364,N_611,N_869);
or U1365 (N_1365,N_534,N_695);
or U1366 (N_1366,N_520,N_756);
nand U1367 (N_1367,N_723,N_624);
xor U1368 (N_1368,N_646,N_576);
and U1369 (N_1369,N_687,N_820);
or U1370 (N_1370,N_749,N_527);
nand U1371 (N_1371,N_681,N_699);
xnor U1372 (N_1372,N_872,N_865);
and U1373 (N_1373,N_997,N_850);
xnor U1374 (N_1374,N_939,N_860);
nor U1375 (N_1375,N_770,N_888);
and U1376 (N_1376,N_862,N_642);
nand U1377 (N_1377,N_856,N_568);
nand U1378 (N_1378,N_972,N_905);
or U1379 (N_1379,N_888,N_984);
nand U1380 (N_1380,N_544,N_866);
nand U1381 (N_1381,N_780,N_942);
nor U1382 (N_1382,N_788,N_559);
nor U1383 (N_1383,N_703,N_588);
and U1384 (N_1384,N_782,N_671);
nor U1385 (N_1385,N_811,N_809);
and U1386 (N_1386,N_570,N_696);
nand U1387 (N_1387,N_869,N_911);
nor U1388 (N_1388,N_727,N_767);
nand U1389 (N_1389,N_757,N_745);
xnor U1390 (N_1390,N_911,N_988);
xnor U1391 (N_1391,N_555,N_556);
and U1392 (N_1392,N_874,N_879);
nand U1393 (N_1393,N_722,N_850);
xor U1394 (N_1394,N_535,N_986);
and U1395 (N_1395,N_841,N_950);
and U1396 (N_1396,N_918,N_895);
and U1397 (N_1397,N_505,N_617);
xnor U1398 (N_1398,N_759,N_893);
nand U1399 (N_1399,N_991,N_904);
nand U1400 (N_1400,N_844,N_803);
nand U1401 (N_1401,N_593,N_657);
and U1402 (N_1402,N_536,N_718);
nand U1403 (N_1403,N_837,N_550);
or U1404 (N_1404,N_635,N_881);
or U1405 (N_1405,N_611,N_901);
xor U1406 (N_1406,N_642,N_705);
xor U1407 (N_1407,N_995,N_714);
or U1408 (N_1408,N_974,N_922);
xor U1409 (N_1409,N_794,N_886);
or U1410 (N_1410,N_555,N_822);
nand U1411 (N_1411,N_954,N_536);
and U1412 (N_1412,N_624,N_856);
xor U1413 (N_1413,N_706,N_516);
xnor U1414 (N_1414,N_973,N_948);
nor U1415 (N_1415,N_502,N_889);
nand U1416 (N_1416,N_574,N_882);
xor U1417 (N_1417,N_602,N_911);
nand U1418 (N_1418,N_595,N_535);
nor U1419 (N_1419,N_835,N_778);
xnor U1420 (N_1420,N_705,N_961);
nand U1421 (N_1421,N_572,N_914);
nor U1422 (N_1422,N_933,N_911);
nor U1423 (N_1423,N_987,N_835);
or U1424 (N_1424,N_984,N_643);
nor U1425 (N_1425,N_963,N_793);
nand U1426 (N_1426,N_511,N_532);
or U1427 (N_1427,N_608,N_972);
nand U1428 (N_1428,N_989,N_957);
or U1429 (N_1429,N_505,N_534);
nand U1430 (N_1430,N_866,N_530);
xnor U1431 (N_1431,N_760,N_665);
or U1432 (N_1432,N_694,N_826);
or U1433 (N_1433,N_610,N_699);
or U1434 (N_1434,N_935,N_876);
xnor U1435 (N_1435,N_530,N_779);
xor U1436 (N_1436,N_832,N_601);
xor U1437 (N_1437,N_526,N_946);
nor U1438 (N_1438,N_927,N_529);
xor U1439 (N_1439,N_808,N_602);
nand U1440 (N_1440,N_765,N_846);
nor U1441 (N_1441,N_649,N_590);
and U1442 (N_1442,N_829,N_657);
or U1443 (N_1443,N_902,N_766);
or U1444 (N_1444,N_556,N_844);
or U1445 (N_1445,N_580,N_868);
nand U1446 (N_1446,N_611,N_785);
nand U1447 (N_1447,N_699,N_676);
and U1448 (N_1448,N_742,N_663);
nor U1449 (N_1449,N_745,N_618);
xor U1450 (N_1450,N_564,N_858);
nand U1451 (N_1451,N_658,N_568);
nor U1452 (N_1452,N_856,N_952);
xnor U1453 (N_1453,N_709,N_618);
nor U1454 (N_1454,N_618,N_925);
xnor U1455 (N_1455,N_647,N_768);
or U1456 (N_1456,N_921,N_771);
nor U1457 (N_1457,N_831,N_769);
nand U1458 (N_1458,N_706,N_809);
nand U1459 (N_1459,N_654,N_849);
nand U1460 (N_1460,N_678,N_666);
nand U1461 (N_1461,N_596,N_909);
nand U1462 (N_1462,N_539,N_509);
nor U1463 (N_1463,N_517,N_927);
or U1464 (N_1464,N_817,N_676);
xnor U1465 (N_1465,N_666,N_665);
or U1466 (N_1466,N_734,N_987);
or U1467 (N_1467,N_847,N_905);
or U1468 (N_1468,N_504,N_766);
xor U1469 (N_1469,N_865,N_537);
nand U1470 (N_1470,N_674,N_763);
xor U1471 (N_1471,N_997,N_993);
xor U1472 (N_1472,N_564,N_843);
or U1473 (N_1473,N_680,N_815);
xor U1474 (N_1474,N_553,N_845);
nor U1475 (N_1475,N_955,N_632);
or U1476 (N_1476,N_656,N_739);
xor U1477 (N_1477,N_843,N_799);
xnor U1478 (N_1478,N_558,N_917);
nor U1479 (N_1479,N_931,N_574);
xor U1480 (N_1480,N_556,N_897);
and U1481 (N_1481,N_704,N_611);
nand U1482 (N_1482,N_730,N_903);
nor U1483 (N_1483,N_549,N_736);
and U1484 (N_1484,N_997,N_531);
nor U1485 (N_1485,N_886,N_652);
and U1486 (N_1486,N_572,N_837);
and U1487 (N_1487,N_563,N_810);
xor U1488 (N_1488,N_584,N_745);
or U1489 (N_1489,N_920,N_553);
xor U1490 (N_1490,N_530,N_563);
or U1491 (N_1491,N_644,N_809);
xnor U1492 (N_1492,N_573,N_557);
nand U1493 (N_1493,N_648,N_914);
and U1494 (N_1494,N_937,N_669);
xnor U1495 (N_1495,N_510,N_757);
or U1496 (N_1496,N_718,N_519);
and U1497 (N_1497,N_822,N_789);
or U1498 (N_1498,N_603,N_757);
xor U1499 (N_1499,N_694,N_829);
and U1500 (N_1500,N_1441,N_1211);
xor U1501 (N_1501,N_1394,N_1120);
and U1502 (N_1502,N_1095,N_1022);
nor U1503 (N_1503,N_1130,N_1218);
and U1504 (N_1504,N_1264,N_1055);
xor U1505 (N_1505,N_1207,N_1242);
and U1506 (N_1506,N_1188,N_1311);
nand U1507 (N_1507,N_1252,N_1493);
or U1508 (N_1508,N_1148,N_1062);
and U1509 (N_1509,N_1116,N_1092);
xor U1510 (N_1510,N_1205,N_1097);
nand U1511 (N_1511,N_1412,N_1079);
xnor U1512 (N_1512,N_1291,N_1017);
and U1513 (N_1513,N_1359,N_1047);
or U1514 (N_1514,N_1112,N_1030);
or U1515 (N_1515,N_1370,N_1300);
xnor U1516 (N_1516,N_1201,N_1243);
xor U1517 (N_1517,N_1089,N_1115);
or U1518 (N_1518,N_1477,N_1444);
and U1519 (N_1519,N_1001,N_1103);
nor U1520 (N_1520,N_1490,N_1009);
and U1521 (N_1521,N_1471,N_1425);
and U1522 (N_1522,N_1111,N_1363);
or U1523 (N_1523,N_1183,N_1121);
nor U1524 (N_1524,N_1100,N_1373);
nor U1525 (N_1525,N_1194,N_1023);
and U1526 (N_1526,N_1048,N_1384);
xnor U1527 (N_1527,N_1074,N_1254);
and U1528 (N_1528,N_1267,N_1463);
nand U1529 (N_1529,N_1169,N_1027);
and U1530 (N_1530,N_1497,N_1261);
nand U1531 (N_1531,N_1228,N_1386);
nand U1532 (N_1532,N_1197,N_1481);
or U1533 (N_1533,N_1485,N_1449);
xnor U1534 (N_1534,N_1478,N_1126);
or U1535 (N_1535,N_1277,N_1331);
nor U1536 (N_1536,N_1230,N_1436);
or U1537 (N_1537,N_1329,N_1338);
or U1538 (N_1538,N_1305,N_1245);
and U1539 (N_1539,N_1470,N_1308);
nor U1540 (N_1540,N_1282,N_1298);
nand U1541 (N_1541,N_1202,N_1256);
xnor U1542 (N_1542,N_1145,N_1052);
xor U1543 (N_1543,N_1378,N_1339);
xor U1544 (N_1544,N_1426,N_1408);
or U1545 (N_1545,N_1283,N_1389);
and U1546 (N_1546,N_1357,N_1216);
xnor U1547 (N_1547,N_1401,N_1402);
nand U1548 (N_1548,N_1193,N_1434);
nor U1549 (N_1549,N_1281,N_1396);
xnor U1550 (N_1550,N_1446,N_1303);
nand U1551 (N_1551,N_1135,N_1072);
nor U1552 (N_1552,N_1035,N_1483);
or U1553 (N_1553,N_1102,N_1340);
nor U1554 (N_1554,N_1475,N_1117);
or U1555 (N_1555,N_1123,N_1227);
xnor U1556 (N_1556,N_1286,N_1025);
xnor U1557 (N_1557,N_1088,N_1179);
nand U1558 (N_1558,N_1270,N_1044);
xor U1559 (N_1559,N_1445,N_1204);
nor U1560 (N_1560,N_1375,N_1450);
or U1561 (N_1561,N_1390,N_1090);
nand U1562 (N_1562,N_1220,N_1301);
nor U1563 (N_1563,N_1149,N_1186);
nor U1564 (N_1564,N_1255,N_1174);
or U1565 (N_1565,N_1020,N_1209);
and U1566 (N_1566,N_1224,N_1366);
nor U1567 (N_1567,N_1101,N_1320);
nand U1568 (N_1568,N_1053,N_1353);
nand U1569 (N_1569,N_1073,N_1068);
or U1570 (N_1570,N_1365,N_1178);
xor U1571 (N_1571,N_1146,N_1181);
xnor U1572 (N_1572,N_1464,N_1295);
or U1573 (N_1573,N_1438,N_1312);
or U1574 (N_1574,N_1385,N_1292);
nor U1575 (N_1575,N_1050,N_1410);
or U1576 (N_1576,N_1031,N_1419);
nor U1577 (N_1577,N_1010,N_1461);
or U1578 (N_1578,N_1343,N_1085);
xor U1579 (N_1579,N_1422,N_1466);
nor U1580 (N_1580,N_1288,N_1119);
and U1581 (N_1581,N_1003,N_1381);
and U1582 (N_1582,N_1356,N_1240);
nand U1583 (N_1583,N_1259,N_1387);
and U1584 (N_1584,N_1223,N_1488);
or U1585 (N_1585,N_1248,N_1362);
xor U1586 (N_1586,N_1316,N_1173);
or U1587 (N_1587,N_1057,N_1236);
and U1588 (N_1588,N_1206,N_1448);
or U1589 (N_1589,N_1212,N_1491);
or U1590 (N_1590,N_1299,N_1176);
and U1591 (N_1591,N_1345,N_1285);
xnor U1592 (N_1592,N_1021,N_1302);
nor U1593 (N_1593,N_1042,N_1417);
and U1594 (N_1594,N_1274,N_1349);
nor U1595 (N_1595,N_1067,N_1170);
nand U1596 (N_1596,N_1296,N_1371);
xor U1597 (N_1597,N_1383,N_1189);
nand U1598 (N_1598,N_1162,N_1143);
nor U1599 (N_1599,N_1262,N_1087);
nand U1600 (N_1600,N_1036,N_1203);
xor U1601 (N_1601,N_1238,N_1428);
nand U1602 (N_1602,N_1225,N_1019);
xnor U1603 (N_1603,N_1219,N_1114);
or U1604 (N_1604,N_1213,N_1108);
nor U1605 (N_1605,N_1420,N_1458);
and U1606 (N_1606,N_1499,N_1451);
or U1607 (N_1607,N_1468,N_1215);
xnor U1608 (N_1608,N_1165,N_1156);
and U1609 (N_1609,N_1016,N_1004);
and U1610 (N_1610,N_1078,N_1234);
xor U1611 (N_1611,N_1495,N_1086);
and U1612 (N_1612,N_1239,N_1406);
nor U1613 (N_1613,N_1155,N_1005);
nor U1614 (N_1614,N_1226,N_1456);
or U1615 (N_1615,N_1435,N_1460);
and U1616 (N_1616,N_1352,N_1093);
nor U1617 (N_1617,N_1433,N_1138);
and U1618 (N_1618,N_1398,N_1134);
and U1619 (N_1619,N_1034,N_1026);
nor U1620 (N_1620,N_1033,N_1465);
and U1621 (N_1621,N_1071,N_1336);
xor U1622 (N_1622,N_1427,N_1000);
and U1623 (N_1623,N_1253,N_1437);
and U1624 (N_1624,N_1271,N_1018);
nand U1625 (N_1625,N_1421,N_1399);
xnor U1626 (N_1626,N_1081,N_1457);
nand U1627 (N_1627,N_1011,N_1013);
nor U1628 (N_1628,N_1147,N_1158);
nor U1629 (N_1629,N_1144,N_1309);
and U1630 (N_1630,N_1037,N_1214);
and U1631 (N_1631,N_1166,N_1258);
xor U1632 (N_1632,N_1131,N_1229);
nor U1633 (N_1633,N_1455,N_1304);
nand U1634 (N_1634,N_1342,N_1122);
xnor U1635 (N_1635,N_1452,N_1063);
or U1636 (N_1636,N_1480,N_1392);
nor U1637 (N_1637,N_1479,N_1322);
or U1638 (N_1638,N_1476,N_1064);
and U1639 (N_1639,N_1247,N_1096);
or U1640 (N_1640,N_1028,N_1473);
and U1641 (N_1641,N_1498,N_1269);
nand U1642 (N_1642,N_1196,N_1486);
or U1643 (N_1643,N_1289,N_1208);
or U1644 (N_1644,N_1182,N_1376);
nor U1645 (N_1645,N_1045,N_1418);
nand U1646 (N_1646,N_1127,N_1113);
nor U1647 (N_1647,N_1235,N_1484);
nand U1648 (N_1648,N_1335,N_1453);
nand U1649 (N_1649,N_1266,N_1374);
or U1650 (N_1650,N_1462,N_1423);
or U1651 (N_1651,N_1447,N_1040);
or U1652 (N_1652,N_1190,N_1128);
nor U1653 (N_1653,N_1327,N_1459);
nor U1654 (N_1654,N_1066,N_1132);
or U1655 (N_1655,N_1222,N_1251);
nor U1656 (N_1656,N_1391,N_1163);
nor U1657 (N_1657,N_1152,N_1429);
nor U1658 (N_1658,N_1319,N_1334);
xnor U1659 (N_1659,N_1413,N_1284);
xor U1660 (N_1660,N_1397,N_1184);
nand U1661 (N_1661,N_1325,N_1249);
xor U1662 (N_1662,N_1354,N_1210);
nor U1663 (N_1663,N_1056,N_1041);
xor U1664 (N_1664,N_1489,N_1440);
xnor U1665 (N_1665,N_1124,N_1136);
and U1666 (N_1666,N_1099,N_1257);
and U1667 (N_1667,N_1313,N_1142);
nand U1668 (N_1668,N_1054,N_1341);
and U1669 (N_1669,N_1487,N_1377);
or U1670 (N_1670,N_1180,N_1323);
nand U1671 (N_1671,N_1060,N_1175);
xor U1672 (N_1672,N_1454,N_1046);
nor U1673 (N_1673,N_1129,N_1315);
xor U1674 (N_1674,N_1008,N_1395);
xor U1675 (N_1675,N_1279,N_1109);
and U1676 (N_1676,N_1140,N_1415);
nor U1677 (N_1677,N_1405,N_1409);
nand U1678 (N_1678,N_1172,N_1012);
nor U1679 (N_1679,N_1075,N_1177);
and U1680 (N_1680,N_1107,N_1442);
xnor U1681 (N_1681,N_1159,N_1355);
nand U1682 (N_1682,N_1431,N_1082);
xnor U1683 (N_1683,N_1157,N_1091);
and U1684 (N_1684,N_1198,N_1306);
nand U1685 (N_1685,N_1039,N_1280);
nor U1686 (N_1686,N_1358,N_1348);
nor U1687 (N_1687,N_1015,N_1411);
xnor U1688 (N_1688,N_1346,N_1246);
nor U1689 (N_1689,N_1141,N_1380);
and U1690 (N_1690,N_1192,N_1344);
nor U1691 (N_1691,N_1061,N_1482);
or U1692 (N_1692,N_1199,N_1032);
nand U1693 (N_1693,N_1439,N_1098);
or U1694 (N_1694,N_1424,N_1469);
nand U1695 (N_1695,N_1195,N_1369);
xnor U1696 (N_1696,N_1058,N_1161);
xnor U1697 (N_1697,N_1231,N_1139);
nor U1698 (N_1698,N_1076,N_1432);
and U1699 (N_1699,N_1367,N_1276);
nor U1700 (N_1700,N_1250,N_1330);
xor U1701 (N_1701,N_1494,N_1029);
xnor U1702 (N_1702,N_1467,N_1038);
and U1703 (N_1703,N_1360,N_1265);
nor U1704 (N_1704,N_1492,N_1137);
nand U1705 (N_1705,N_1350,N_1400);
or U1706 (N_1706,N_1065,N_1294);
nor U1707 (N_1707,N_1070,N_1150);
nor U1708 (N_1708,N_1191,N_1154);
nand U1709 (N_1709,N_1110,N_1404);
or U1710 (N_1710,N_1043,N_1472);
nor U1711 (N_1711,N_1326,N_1407);
or U1712 (N_1712,N_1049,N_1105);
and U1713 (N_1713,N_1321,N_1151);
nor U1714 (N_1714,N_1310,N_1168);
and U1715 (N_1715,N_1187,N_1347);
or U1716 (N_1716,N_1153,N_1361);
xor U1717 (N_1717,N_1263,N_1474);
or U1718 (N_1718,N_1233,N_1443);
nand U1719 (N_1719,N_1051,N_1059);
nand U1720 (N_1720,N_1006,N_1167);
nand U1721 (N_1721,N_1317,N_1232);
nand U1722 (N_1722,N_1118,N_1297);
nor U1723 (N_1723,N_1333,N_1077);
nor U1724 (N_1724,N_1318,N_1268);
nor U1725 (N_1725,N_1379,N_1094);
nand U1726 (N_1726,N_1069,N_1244);
nand U1727 (N_1727,N_1337,N_1314);
or U1728 (N_1728,N_1241,N_1272);
xnor U1729 (N_1729,N_1382,N_1307);
and U1730 (N_1730,N_1364,N_1200);
nor U1731 (N_1731,N_1416,N_1125);
nor U1732 (N_1732,N_1278,N_1414);
and U1733 (N_1733,N_1185,N_1024);
xnor U1734 (N_1734,N_1104,N_1393);
or U1735 (N_1735,N_1293,N_1160);
nor U1736 (N_1736,N_1106,N_1084);
nand U1737 (N_1737,N_1368,N_1324);
xor U1738 (N_1738,N_1133,N_1171);
nor U1739 (N_1739,N_1328,N_1014);
nor U1740 (N_1740,N_1275,N_1080);
and U1741 (N_1741,N_1273,N_1388);
xor U1742 (N_1742,N_1002,N_1430);
or U1743 (N_1743,N_1164,N_1496);
and U1744 (N_1744,N_1221,N_1372);
nand U1745 (N_1745,N_1260,N_1332);
nor U1746 (N_1746,N_1351,N_1287);
xor U1747 (N_1747,N_1007,N_1403);
or U1748 (N_1748,N_1237,N_1217);
nand U1749 (N_1749,N_1290,N_1083);
xor U1750 (N_1750,N_1367,N_1266);
or U1751 (N_1751,N_1151,N_1007);
and U1752 (N_1752,N_1269,N_1259);
or U1753 (N_1753,N_1300,N_1434);
and U1754 (N_1754,N_1237,N_1299);
nand U1755 (N_1755,N_1151,N_1315);
nor U1756 (N_1756,N_1086,N_1354);
nand U1757 (N_1757,N_1358,N_1353);
or U1758 (N_1758,N_1124,N_1447);
nor U1759 (N_1759,N_1167,N_1370);
or U1760 (N_1760,N_1077,N_1320);
nand U1761 (N_1761,N_1162,N_1477);
nand U1762 (N_1762,N_1329,N_1297);
and U1763 (N_1763,N_1173,N_1364);
xor U1764 (N_1764,N_1203,N_1484);
xnor U1765 (N_1765,N_1397,N_1380);
nand U1766 (N_1766,N_1275,N_1372);
nand U1767 (N_1767,N_1022,N_1381);
or U1768 (N_1768,N_1438,N_1094);
or U1769 (N_1769,N_1080,N_1225);
and U1770 (N_1770,N_1329,N_1430);
and U1771 (N_1771,N_1228,N_1419);
and U1772 (N_1772,N_1297,N_1184);
xor U1773 (N_1773,N_1113,N_1061);
or U1774 (N_1774,N_1181,N_1460);
or U1775 (N_1775,N_1286,N_1180);
nor U1776 (N_1776,N_1215,N_1445);
nor U1777 (N_1777,N_1028,N_1437);
and U1778 (N_1778,N_1091,N_1325);
xnor U1779 (N_1779,N_1178,N_1033);
or U1780 (N_1780,N_1300,N_1218);
nor U1781 (N_1781,N_1284,N_1457);
xor U1782 (N_1782,N_1098,N_1218);
and U1783 (N_1783,N_1472,N_1010);
nor U1784 (N_1784,N_1148,N_1021);
and U1785 (N_1785,N_1063,N_1258);
nand U1786 (N_1786,N_1322,N_1325);
nand U1787 (N_1787,N_1205,N_1390);
or U1788 (N_1788,N_1078,N_1137);
nor U1789 (N_1789,N_1007,N_1395);
and U1790 (N_1790,N_1342,N_1051);
nor U1791 (N_1791,N_1180,N_1430);
nor U1792 (N_1792,N_1383,N_1151);
nand U1793 (N_1793,N_1484,N_1399);
or U1794 (N_1794,N_1111,N_1468);
nand U1795 (N_1795,N_1139,N_1035);
and U1796 (N_1796,N_1252,N_1241);
and U1797 (N_1797,N_1159,N_1398);
and U1798 (N_1798,N_1315,N_1093);
xnor U1799 (N_1799,N_1092,N_1406);
xnor U1800 (N_1800,N_1090,N_1384);
nand U1801 (N_1801,N_1030,N_1113);
xor U1802 (N_1802,N_1389,N_1098);
nor U1803 (N_1803,N_1071,N_1499);
nand U1804 (N_1804,N_1264,N_1389);
xnor U1805 (N_1805,N_1487,N_1224);
or U1806 (N_1806,N_1211,N_1412);
nor U1807 (N_1807,N_1381,N_1170);
nand U1808 (N_1808,N_1444,N_1177);
nand U1809 (N_1809,N_1481,N_1326);
xnor U1810 (N_1810,N_1234,N_1302);
xnor U1811 (N_1811,N_1008,N_1124);
nand U1812 (N_1812,N_1316,N_1431);
nor U1813 (N_1813,N_1127,N_1184);
nand U1814 (N_1814,N_1134,N_1086);
or U1815 (N_1815,N_1276,N_1065);
nand U1816 (N_1816,N_1257,N_1467);
xnor U1817 (N_1817,N_1400,N_1351);
nor U1818 (N_1818,N_1482,N_1210);
or U1819 (N_1819,N_1098,N_1115);
nor U1820 (N_1820,N_1334,N_1230);
nor U1821 (N_1821,N_1042,N_1457);
and U1822 (N_1822,N_1162,N_1213);
or U1823 (N_1823,N_1226,N_1074);
nor U1824 (N_1824,N_1332,N_1297);
or U1825 (N_1825,N_1253,N_1445);
and U1826 (N_1826,N_1030,N_1185);
nand U1827 (N_1827,N_1424,N_1291);
and U1828 (N_1828,N_1365,N_1094);
and U1829 (N_1829,N_1225,N_1107);
nor U1830 (N_1830,N_1134,N_1202);
and U1831 (N_1831,N_1043,N_1247);
nand U1832 (N_1832,N_1245,N_1117);
nand U1833 (N_1833,N_1451,N_1245);
and U1834 (N_1834,N_1462,N_1299);
or U1835 (N_1835,N_1368,N_1479);
nor U1836 (N_1836,N_1042,N_1102);
nor U1837 (N_1837,N_1173,N_1458);
nand U1838 (N_1838,N_1172,N_1116);
xnor U1839 (N_1839,N_1032,N_1229);
nor U1840 (N_1840,N_1345,N_1021);
nand U1841 (N_1841,N_1482,N_1193);
or U1842 (N_1842,N_1220,N_1348);
nor U1843 (N_1843,N_1267,N_1180);
xnor U1844 (N_1844,N_1346,N_1430);
and U1845 (N_1845,N_1298,N_1051);
xor U1846 (N_1846,N_1470,N_1426);
xnor U1847 (N_1847,N_1219,N_1411);
nand U1848 (N_1848,N_1406,N_1168);
nand U1849 (N_1849,N_1067,N_1182);
and U1850 (N_1850,N_1297,N_1488);
nor U1851 (N_1851,N_1249,N_1491);
xnor U1852 (N_1852,N_1329,N_1478);
nand U1853 (N_1853,N_1376,N_1387);
xnor U1854 (N_1854,N_1493,N_1365);
xnor U1855 (N_1855,N_1398,N_1392);
nand U1856 (N_1856,N_1370,N_1124);
and U1857 (N_1857,N_1459,N_1063);
or U1858 (N_1858,N_1234,N_1147);
and U1859 (N_1859,N_1411,N_1008);
nor U1860 (N_1860,N_1105,N_1397);
or U1861 (N_1861,N_1378,N_1050);
xor U1862 (N_1862,N_1157,N_1120);
nor U1863 (N_1863,N_1262,N_1489);
and U1864 (N_1864,N_1125,N_1120);
nor U1865 (N_1865,N_1349,N_1438);
or U1866 (N_1866,N_1201,N_1440);
xor U1867 (N_1867,N_1427,N_1041);
nor U1868 (N_1868,N_1486,N_1447);
xor U1869 (N_1869,N_1235,N_1343);
or U1870 (N_1870,N_1398,N_1138);
nor U1871 (N_1871,N_1370,N_1053);
nor U1872 (N_1872,N_1457,N_1304);
nand U1873 (N_1873,N_1414,N_1123);
or U1874 (N_1874,N_1249,N_1375);
nor U1875 (N_1875,N_1213,N_1188);
xor U1876 (N_1876,N_1066,N_1028);
and U1877 (N_1877,N_1166,N_1389);
xnor U1878 (N_1878,N_1246,N_1131);
nor U1879 (N_1879,N_1218,N_1305);
or U1880 (N_1880,N_1302,N_1482);
and U1881 (N_1881,N_1400,N_1146);
and U1882 (N_1882,N_1458,N_1059);
nor U1883 (N_1883,N_1329,N_1446);
nand U1884 (N_1884,N_1386,N_1137);
and U1885 (N_1885,N_1314,N_1293);
or U1886 (N_1886,N_1400,N_1409);
or U1887 (N_1887,N_1289,N_1328);
and U1888 (N_1888,N_1176,N_1200);
and U1889 (N_1889,N_1038,N_1413);
or U1890 (N_1890,N_1266,N_1394);
xor U1891 (N_1891,N_1281,N_1011);
or U1892 (N_1892,N_1253,N_1467);
xor U1893 (N_1893,N_1103,N_1382);
nor U1894 (N_1894,N_1405,N_1478);
nor U1895 (N_1895,N_1320,N_1170);
nand U1896 (N_1896,N_1457,N_1445);
and U1897 (N_1897,N_1023,N_1240);
or U1898 (N_1898,N_1162,N_1250);
nand U1899 (N_1899,N_1128,N_1424);
and U1900 (N_1900,N_1201,N_1009);
nand U1901 (N_1901,N_1339,N_1307);
and U1902 (N_1902,N_1165,N_1351);
and U1903 (N_1903,N_1459,N_1238);
and U1904 (N_1904,N_1458,N_1172);
nand U1905 (N_1905,N_1491,N_1106);
or U1906 (N_1906,N_1028,N_1347);
xor U1907 (N_1907,N_1179,N_1047);
or U1908 (N_1908,N_1420,N_1438);
nor U1909 (N_1909,N_1220,N_1365);
and U1910 (N_1910,N_1279,N_1274);
nor U1911 (N_1911,N_1491,N_1467);
nor U1912 (N_1912,N_1494,N_1205);
xnor U1913 (N_1913,N_1092,N_1101);
and U1914 (N_1914,N_1187,N_1193);
nor U1915 (N_1915,N_1383,N_1381);
nand U1916 (N_1916,N_1471,N_1262);
nand U1917 (N_1917,N_1174,N_1486);
and U1918 (N_1918,N_1075,N_1343);
nor U1919 (N_1919,N_1470,N_1211);
nor U1920 (N_1920,N_1005,N_1301);
or U1921 (N_1921,N_1145,N_1482);
nand U1922 (N_1922,N_1352,N_1243);
and U1923 (N_1923,N_1315,N_1373);
and U1924 (N_1924,N_1187,N_1108);
nor U1925 (N_1925,N_1025,N_1399);
nand U1926 (N_1926,N_1094,N_1360);
and U1927 (N_1927,N_1406,N_1124);
or U1928 (N_1928,N_1119,N_1045);
or U1929 (N_1929,N_1217,N_1134);
or U1930 (N_1930,N_1390,N_1200);
and U1931 (N_1931,N_1491,N_1446);
and U1932 (N_1932,N_1259,N_1042);
xnor U1933 (N_1933,N_1131,N_1191);
or U1934 (N_1934,N_1464,N_1074);
or U1935 (N_1935,N_1138,N_1242);
or U1936 (N_1936,N_1062,N_1491);
xnor U1937 (N_1937,N_1132,N_1292);
nor U1938 (N_1938,N_1455,N_1478);
xor U1939 (N_1939,N_1324,N_1259);
xor U1940 (N_1940,N_1022,N_1132);
nor U1941 (N_1941,N_1110,N_1421);
and U1942 (N_1942,N_1222,N_1303);
and U1943 (N_1943,N_1010,N_1290);
and U1944 (N_1944,N_1082,N_1015);
and U1945 (N_1945,N_1160,N_1056);
and U1946 (N_1946,N_1258,N_1261);
and U1947 (N_1947,N_1320,N_1471);
nor U1948 (N_1948,N_1455,N_1359);
or U1949 (N_1949,N_1379,N_1022);
nor U1950 (N_1950,N_1282,N_1172);
xor U1951 (N_1951,N_1393,N_1477);
nor U1952 (N_1952,N_1271,N_1369);
xor U1953 (N_1953,N_1217,N_1308);
nand U1954 (N_1954,N_1368,N_1373);
and U1955 (N_1955,N_1412,N_1324);
xnor U1956 (N_1956,N_1049,N_1194);
or U1957 (N_1957,N_1189,N_1154);
and U1958 (N_1958,N_1260,N_1366);
or U1959 (N_1959,N_1404,N_1378);
and U1960 (N_1960,N_1127,N_1408);
or U1961 (N_1961,N_1128,N_1488);
nand U1962 (N_1962,N_1130,N_1071);
or U1963 (N_1963,N_1255,N_1432);
and U1964 (N_1964,N_1413,N_1045);
or U1965 (N_1965,N_1116,N_1339);
and U1966 (N_1966,N_1375,N_1162);
or U1967 (N_1967,N_1001,N_1487);
nand U1968 (N_1968,N_1345,N_1449);
nand U1969 (N_1969,N_1313,N_1454);
nor U1970 (N_1970,N_1044,N_1467);
xnor U1971 (N_1971,N_1179,N_1383);
and U1972 (N_1972,N_1243,N_1033);
and U1973 (N_1973,N_1168,N_1192);
xor U1974 (N_1974,N_1274,N_1365);
nor U1975 (N_1975,N_1186,N_1238);
nand U1976 (N_1976,N_1497,N_1255);
nand U1977 (N_1977,N_1142,N_1446);
or U1978 (N_1978,N_1229,N_1435);
xnor U1979 (N_1979,N_1260,N_1450);
xnor U1980 (N_1980,N_1088,N_1337);
or U1981 (N_1981,N_1044,N_1141);
nor U1982 (N_1982,N_1120,N_1456);
and U1983 (N_1983,N_1272,N_1367);
nand U1984 (N_1984,N_1174,N_1049);
nor U1985 (N_1985,N_1382,N_1340);
nor U1986 (N_1986,N_1495,N_1381);
nand U1987 (N_1987,N_1203,N_1389);
xnor U1988 (N_1988,N_1070,N_1352);
and U1989 (N_1989,N_1209,N_1167);
xnor U1990 (N_1990,N_1370,N_1340);
xnor U1991 (N_1991,N_1266,N_1196);
xnor U1992 (N_1992,N_1371,N_1366);
nand U1993 (N_1993,N_1342,N_1007);
nand U1994 (N_1994,N_1143,N_1466);
and U1995 (N_1995,N_1186,N_1460);
or U1996 (N_1996,N_1456,N_1187);
xor U1997 (N_1997,N_1342,N_1140);
xor U1998 (N_1998,N_1322,N_1058);
xnor U1999 (N_1999,N_1233,N_1043);
nor U2000 (N_2000,N_1833,N_1748);
nand U2001 (N_2001,N_1977,N_1566);
nor U2002 (N_2002,N_1600,N_1519);
xnor U2003 (N_2003,N_1796,N_1814);
or U2004 (N_2004,N_1572,N_1969);
nor U2005 (N_2005,N_1551,N_1792);
xnor U2006 (N_2006,N_1992,N_1749);
or U2007 (N_2007,N_1608,N_1564);
and U2008 (N_2008,N_1510,N_1892);
nor U2009 (N_2009,N_1547,N_1898);
and U2010 (N_2010,N_1697,N_1918);
nand U2011 (N_2011,N_1912,N_1528);
xnor U2012 (N_2012,N_1978,N_1894);
nor U2013 (N_2013,N_1987,N_1560);
or U2014 (N_2014,N_1703,N_1944);
and U2015 (N_2015,N_1655,N_1983);
or U2016 (N_2016,N_1872,N_1934);
xnor U2017 (N_2017,N_1902,N_1895);
or U2018 (N_2018,N_1791,N_1946);
xor U2019 (N_2019,N_1900,N_1750);
and U2020 (N_2020,N_1790,N_1505);
xnor U2021 (N_2021,N_1845,N_1878);
xnor U2022 (N_2022,N_1809,N_1786);
and U2023 (N_2023,N_1881,N_1798);
xor U2024 (N_2024,N_1965,N_1532);
nand U2025 (N_2025,N_1587,N_1932);
nor U2026 (N_2026,N_1543,N_1884);
or U2027 (N_2027,N_1621,N_1803);
xor U2028 (N_2028,N_1806,N_1687);
nand U2029 (N_2029,N_1662,N_1939);
nor U2030 (N_2030,N_1901,N_1864);
or U2031 (N_2031,N_1549,N_1619);
nand U2032 (N_2032,N_1550,N_1807);
nor U2033 (N_2033,N_1695,N_1709);
nand U2034 (N_2034,N_1771,N_1778);
nor U2035 (N_2035,N_1635,N_1552);
nand U2036 (N_2036,N_1647,N_1921);
and U2037 (N_2037,N_1599,N_1653);
or U2038 (N_2038,N_1891,N_1883);
and U2039 (N_2039,N_1981,N_1512);
nor U2040 (N_2040,N_1595,N_1527);
nand U2041 (N_2041,N_1625,N_1522);
xor U2042 (N_2042,N_1772,N_1743);
nand U2043 (N_2043,N_1795,N_1908);
or U2044 (N_2044,N_1899,N_1643);
and U2045 (N_2045,N_1879,N_1514);
xor U2046 (N_2046,N_1570,N_1768);
nand U2047 (N_2047,N_1988,N_1936);
xor U2048 (N_2048,N_1553,N_1711);
xnor U2049 (N_2049,N_1859,N_1893);
or U2050 (N_2050,N_1582,N_1870);
nand U2051 (N_2051,N_1729,N_1705);
nand U2052 (N_2052,N_1913,N_1813);
xnor U2053 (N_2053,N_1802,N_1724);
xor U2054 (N_2054,N_1626,N_1673);
and U2055 (N_2055,N_1993,N_1540);
nor U2056 (N_2056,N_1741,N_1947);
and U2057 (N_2057,N_1765,N_1861);
nand U2058 (N_2058,N_1773,N_1661);
xor U2059 (N_2059,N_1829,N_1683);
nand U2060 (N_2060,N_1821,N_1825);
xnor U2061 (N_2061,N_1533,N_1628);
nor U2062 (N_2062,N_1536,N_1719);
nand U2063 (N_2063,N_1685,N_1562);
and U2064 (N_2064,N_1656,N_1822);
nor U2065 (N_2065,N_1559,N_1563);
and U2066 (N_2066,N_1660,N_1865);
nor U2067 (N_2067,N_1592,N_1907);
nor U2068 (N_2068,N_1904,N_1526);
or U2069 (N_2069,N_1797,N_1681);
nand U2070 (N_2070,N_1606,N_1590);
nand U2071 (N_2071,N_1693,N_1758);
nor U2072 (N_2072,N_1967,N_1694);
and U2073 (N_2073,N_1699,N_1708);
or U2074 (N_2074,N_1785,N_1762);
or U2075 (N_2075,N_1961,N_1945);
nand U2076 (N_2076,N_1700,N_1847);
nand U2077 (N_2077,N_1575,N_1996);
and U2078 (N_2078,N_1616,N_1634);
xor U2079 (N_2079,N_1972,N_1763);
nor U2080 (N_2080,N_1827,N_1784);
nor U2081 (N_2081,N_1620,N_1515);
xnor U2082 (N_2082,N_1554,N_1863);
xnor U2083 (N_2083,N_1816,N_1759);
nor U2084 (N_2084,N_1767,N_1935);
nand U2085 (N_2085,N_1714,N_1557);
xnor U2086 (N_2086,N_1874,N_1757);
nor U2087 (N_2087,N_1876,N_1506);
or U2088 (N_2088,N_1732,N_1530);
nor U2089 (N_2089,N_1607,N_1820);
and U2090 (N_2090,N_1648,N_1836);
xor U2091 (N_2091,N_1941,N_1818);
xnor U2092 (N_2092,N_1511,N_1531);
nor U2093 (N_2093,N_1696,N_1742);
or U2094 (N_2094,N_1672,N_1609);
nor U2095 (N_2095,N_1513,N_1556);
nand U2096 (N_2096,N_1659,N_1832);
xnor U2097 (N_2097,N_1905,N_1966);
nand U2098 (N_2098,N_1544,N_1931);
or U2099 (N_2099,N_1546,N_1594);
or U2100 (N_2100,N_1914,N_1801);
nand U2101 (N_2101,N_1523,N_1623);
or U2102 (N_2102,N_1760,N_1555);
nor U2103 (N_2103,N_1747,N_1610);
and U2104 (N_2104,N_1986,N_1886);
nor U2105 (N_2105,N_1689,N_1840);
and U2106 (N_2106,N_1985,N_1928);
xor U2107 (N_2107,N_1975,N_1999);
xnor U2108 (N_2108,N_1882,N_1835);
or U2109 (N_2109,N_1518,N_1811);
nor U2110 (N_2110,N_1869,N_1614);
xor U2111 (N_2111,N_1585,N_1989);
or U2112 (N_2112,N_1633,N_1667);
or U2113 (N_2113,N_1507,N_1657);
xor U2114 (N_2114,N_1823,N_1764);
xor U2115 (N_2115,N_1508,N_1770);
nand U2116 (N_2116,N_1670,N_1800);
xnor U2117 (N_2117,N_1520,N_1851);
nor U2118 (N_2118,N_1794,N_1777);
nand U2119 (N_2119,N_1754,N_1862);
or U2120 (N_2120,N_1578,N_1596);
nand U2121 (N_2121,N_1516,N_1871);
xnor U2122 (N_2122,N_1500,N_1730);
or U2123 (N_2123,N_1682,N_1558);
nand U2124 (N_2124,N_1929,N_1702);
xnor U2125 (N_2125,N_1644,N_1974);
nor U2126 (N_2126,N_1752,N_1678);
or U2127 (N_2127,N_1571,N_1976);
xor U2128 (N_2128,N_1715,N_1776);
xor U2129 (N_2129,N_1793,N_1873);
nand U2130 (N_2130,N_1680,N_1805);
nor U2131 (N_2131,N_1979,N_1537);
or U2132 (N_2132,N_1632,N_1538);
and U2133 (N_2133,N_1677,N_1860);
nor U2134 (N_2134,N_1915,N_1710);
nand U2135 (N_2135,N_1542,N_1775);
xor U2136 (N_2136,N_1855,N_1501);
xor U2137 (N_2137,N_1639,N_1957);
xnor U2138 (N_2138,N_1645,N_1924);
xnor U2139 (N_2139,N_1735,N_1788);
and U2140 (N_2140,N_1642,N_1938);
or U2141 (N_2141,N_1964,N_1815);
nor U2142 (N_2142,N_1545,N_1517);
nor U2143 (N_2143,N_1841,N_1927);
nand U2144 (N_2144,N_1674,N_1812);
or U2145 (N_2145,N_1712,N_1854);
and U2146 (N_2146,N_1923,N_1612);
and U2147 (N_2147,N_1630,N_1573);
and U2148 (N_2148,N_1658,N_1723);
and U2149 (N_2149,N_1991,N_1942);
or U2150 (N_2150,N_1651,N_1875);
nor U2151 (N_2151,N_1525,N_1718);
xnor U2152 (N_2152,N_1819,N_1541);
nor U2153 (N_2153,N_1997,N_1953);
or U2154 (N_2154,N_1679,N_1982);
xor U2155 (N_2155,N_1774,N_1637);
xnor U2156 (N_2156,N_1769,N_1745);
or U2157 (N_2157,N_1627,N_1713);
nor U2158 (N_2158,N_1706,N_1916);
xor U2159 (N_2159,N_1668,N_1641);
xnor U2160 (N_2160,N_1911,N_1728);
and U2161 (N_2161,N_1684,N_1605);
or U2162 (N_2162,N_1738,N_1583);
and U2163 (N_2163,N_1922,N_1624);
nor U2164 (N_2164,N_1799,N_1839);
or U2165 (N_2165,N_1910,N_1740);
nand U2166 (N_2166,N_1690,N_1720);
nand U2167 (N_2167,N_1830,N_1849);
nor U2168 (N_2168,N_1810,N_1737);
nor U2169 (N_2169,N_1579,N_1613);
nand U2170 (N_2170,N_1756,N_1604);
and U2171 (N_2171,N_1888,N_1949);
and U2172 (N_2172,N_1726,N_1828);
nand U2173 (N_2173,N_1890,N_1725);
nor U2174 (N_2174,N_1837,N_1846);
and U2175 (N_2175,N_1903,N_1733);
or U2176 (N_2176,N_1727,N_1850);
nor U2177 (N_2177,N_1868,N_1817);
nor U2178 (N_2178,N_1766,N_1780);
xor U2179 (N_2179,N_1569,N_1664);
and U2180 (N_2180,N_1686,N_1831);
xnor U2181 (N_2181,N_1521,N_1692);
xnor U2182 (N_2182,N_1652,N_1808);
xnor U2183 (N_2183,N_1958,N_1940);
xor U2184 (N_2184,N_1937,N_1843);
and U2185 (N_2185,N_1857,N_1646);
and U2186 (N_2186,N_1565,N_1885);
nor U2187 (N_2187,N_1603,N_1707);
and U2188 (N_2188,N_1926,N_1663);
nand U2189 (N_2189,N_1970,N_1804);
and U2190 (N_2190,N_1746,N_1751);
nor U2191 (N_2191,N_1834,N_1665);
or U2192 (N_2192,N_1618,N_1995);
or U2193 (N_2193,N_1971,N_1504);
nand U2194 (N_2194,N_1617,N_1950);
xor U2195 (N_2195,N_1602,N_1649);
xor U2196 (N_2196,N_1586,N_1669);
and U2197 (N_2197,N_1675,N_1755);
or U2198 (N_2198,N_1574,N_1753);
and U2199 (N_2199,N_1568,N_1920);
nand U2200 (N_2200,N_1853,N_1998);
and U2201 (N_2201,N_1848,N_1629);
nand U2202 (N_2202,N_1844,N_1704);
nand U2203 (N_2203,N_1781,N_1509);
nor U2204 (N_2204,N_1880,N_1676);
nand U2205 (N_2205,N_1638,N_1539);
nor U2206 (N_2206,N_1581,N_1734);
xnor U2207 (N_2207,N_1503,N_1994);
nand U2208 (N_2208,N_1666,N_1783);
xnor U2209 (N_2209,N_1968,N_1889);
nor U2210 (N_2210,N_1789,N_1906);
and U2211 (N_2211,N_1973,N_1593);
nor U2212 (N_2212,N_1548,N_1896);
and U2213 (N_2213,N_1866,N_1909);
xor U2214 (N_2214,N_1636,N_1650);
or U2215 (N_2215,N_1761,N_1654);
nor U2216 (N_2216,N_1561,N_1640);
and U2217 (N_2217,N_1591,N_1824);
xor U2218 (N_2218,N_1980,N_1960);
nor U2219 (N_2219,N_1739,N_1887);
xnor U2220 (N_2220,N_1826,N_1917);
and U2221 (N_2221,N_1731,N_1577);
nand U2222 (N_2222,N_1722,N_1779);
xnor U2223 (N_2223,N_1721,N_1524);
nor U2224 (N_2224,N_1535,N_1930);
and U2225 (N_2225,N_1867,N_1584);
xor U2226 (N_2226,N_1688,N_1744);
and U2227 (N_2227,N_1671,N_1601);
nor U2228 (N_2228,N_1952,N_1502);
nand U2229 (N_2229,N_1787,N_1597);
and U2230 (N_2230,N_1951,N_1838);
nand U2231 (N_2231,N_1611,N_1919);
xor U2232 (N_2232,N_1580,N_1691);
or U2233 (N_2233,N_1534,N_1856);
or U2234 (N_2234,N_1716,N_1598);
or U2235 (N_2235,N_1943,N_1588);
and U2236 (N_2236,N_1567,N_1925);
or U2237 (N_2237,N_1990,N_1576);
nor U2238 (N_2238,N_1984,N_1631);
and U2239 (N_2239,N_1736,N_1955);
and U2240 (N_2240,N_1858,N_1956);
nor U2241 (N_2241,N_1954,N_1948);
nor U2242 (N_2242,N_1959,N_1717);
or U2243 (N_2243,N_1615,N_1933);
nor U2244 (N_2244,N_1589,N_1782);
or U2245 (N_2245,N_1622,N_1897);
or U2246 (N_2246,N_1962,N_1877);
nor U2247 (N_2247,N_1698,N_1852);
xor U2248 (N_2248,N_1529,N_1701);
nand U2249 (N_2249,N_1963,N_1842);
nand U2250 (N_2250,N_1966,N_1591);
xor U2251 (N_2251,N_1932,N_1769);
nor U2252 (N_2252,N_1699,N_1711);
xnor U2253 (N_2253,N_1794,N_1830);
nor U2254 (N_2254,N_1777,N_1683);
or U2255 (N_2255,N_1813,N_1517);
nor U2256 (N_2256,N_1994,N_1820);
nand U2257 (N_2257,N_1718,N_1728);
or U2258 (N_2258,N_1770,N_1564);
or U2259 (N_2259,N_1697,N_1615);
or U2260 (N_2260,N_1983,N_1577);
xor U2261 (N_2261,N_1833,N_1766);
nand U2262 (N_2262,N_1753,N_1900);
nor U2263 (N_2263,N_1965,N_1782);
nor U2264 (N_2264,N_1567,N_1514);
xnor U2265 (N_2265,N_1556,N_1636);
or U2266 (N_2266,N_1811,N_1829);
nor U2267 (N_2267,N_1779,N_1619);
nand U2268 (N_2268,N_1680,N_1576);
nor U2269 (N_2269,N_1879,N_1778);
nor U2270 (N_2270,N_1924,N_1500);
or U2271 (N_2271,N_1645,N_1681);
xor U2272 (N_2272,N_1590,N_1768);
xor U2273 (N_2273,N_1702,N_1556);
nor U2274 (N_2274,N_1572,N_1867);
or U2275 (N_2275,N_1955,N_1613);
nand U2276 (N_2276,N_1805,N_1564);
or U2277 (N_2277,N_1815,N_1986);
nor U2278 (N_2278,N_1720,N_1765);
nand U2279 (N_2279,N_1737,N_1639);
nor U2280 (N_2280,N_1987,N_1630);
or U2281 (N_2281,N_1978,N_1827);
nor U2282 (N_2282,N_1870,N_1905);
xor U2283 (N_2283,N_1761,N_1552);
nand U2284 (N_2284,N_1821,N_1976);
nand U2285 (N_2285,N_1777,N_1764);
or U2286 (N_2286,N_1943,N_1983);
xor U2287 (N_2287,N_1588,N_1869);
and U2288 (N_2288,N_1822,N_1725);
or U2289 (N_2289,N_1685,N_1594);
xnor U2290 (N_2290,N_1709,N_1570);
or U2291 (N_2291,N_1627,N_1892);
nand U2292 (N_2292,N_1611,N_1666);
nand U2293 (N_2293,N_1918,N_1863);
or U2294 (N_2294,N_1607,N_1672);
or U2295 (N_2295,N_1895,N_1855);
nor U2296 (N_2296,N_1614,N_1767);
and U2297 (N_2297,N_1615,N_1717);
or U2298 (N_2298,N_1775,N_1862);
or U2299 (N_2299,N_1854,N_1618);
xor U2300 (N_2300,N_1779,N_1836);
nand U2301 (N_2301,N_1883,N_1607);
xor U2302 (N_2302,N_1726,N_1905);
nor U2303 (N_2303,N_1921,N_1700);
or U2304 (N_2304,N_1929,N_1899);
xor U2305 (N_2305,N_1967,N_1782);
and U2306 (N_2306,N_1656,N_1689);
nor U2307 (N_2307,N_1682,N_1688);
and U2308 (N_2308,N_1956,N_1760);
xnor U2309 (N_2309,N_1654,N_1848);
xnor U2310 (N_2310,N_1758,N_1917);
and U2311 (N_2311,N_1900,N_1963);
nand U2312 (N_2312,N_1954,N_1780);
nor U2313 (N_2313,N_1571,N_1593);
or U2314 (N_2314,N_1693,N_1517);
nor U2315 (N_2315,N_1961,N_1725);
and U2316 (N_2316,N_1533,N_1669);
xor U2317 (N_2317,N_1531,N_1526);
xor U2318 (N_2318,N_1826,N_1844);
and U2319 (N_2319,N_1610,N_1940);
or U2320 (N_2320,N_1542,N_1955);
xor U2321 (N_2321,N_1718,N_1922);
and U2322 (N_2322,N_1829,N_1660);
nand U2323 (N_2323,N_1525,N_1592);
xnor U2324 (N_2324,N_1502,N_1517);
nand U2325 (N_2325,N_1811,N_1819);
and U2326 (N_2326,N_1512,N_1721);
and U2327 (N_2327,N_1961,N_1937);
and U2328 (N_2328,N_1944,N_1686);
and U2329 (N_2329,N_1761,N_1824);
nand U2330 (N_2330,N_1664,N_1877);
nor U2331 (N_2331,N_1680,N_1523);
or U2332 (N_2332,N_1808,N_1647);
and U2333 (N_2333,N_1821,N_1583);
and U2334 (N_2334,N_1840,N_1510);
nor U2335 (N_2335,N_1597,N_1988);
nor U2336 (N_2336,N_1569,N_1882);
xor U2337 (N_2337,N_1640,N_1967);
or U2338 (N_2338,N_1945,N_1795);
xor U2339 (N_2339,N_1947,N_1720);
or U2340 (N_2340,N_1940,N_1576);
nor U2341 (N_2341,N_1879,N_1516);
xor U2342 (N_2342,N_1883,N_1525);
and U2343 (N_2343,N_1864,N_1632);
and U2344 (N_2344,N_1880,N_1793);
and U2345 (N_2345,N_1918,N_1736);
and U2346 (N_2346,N_1551,N_1989);
and U2347 (N_2347,N_1945,N_1887);
and U2348 (N_2348,N_1855,N_1955);
nand U2349 (N_2349,N_1816,N_1788);
nand U2350 (N_2350,N_1759,N_1570);
nor U2351 (N_2351,N_1554,N_1900);
xnor U2352 (N_2352,N_1857,N_1694);
and U2353 (N_2353,N_1746,N_1586);
nor U2354 (N_2354,N_1571,N_1852);
and U2355 (N_2355,N_1764,N_1960);
nor U2356 (N_2356,N_1870,N_1788);
and U2357 (N_2357,N_1673,N_1535);
xor U2358 (N_2358,N_1583,N_1790);
and U2359 (N_2359,N_1905,N_1685);
or U2360 (N_2360,N_1837,N_1987);
nand U2361 (N_2361,N_1775,N_1974);
nor U2362 (N_2362,N_1710,N_1655);
nand U2363 (N_2363,N_1788,N_1695);
or U2364 (N_2364,N_1632,N_1563);
xnor U2365 (N_2365,N_1827,N_1710);
and U2366 (N_2366,N_1536,N_1939);
or U2367 (N_2367,N_1652,N_1904);
and U2368 (N_2368,N_1875,N_1782);
nor U2369 (N_2369,N_1621,N_1652);
xor U2370 (N_2370,N_1928,N_1745);
nor U2371 (N_2371,N_1512,N_1530);
nor U2372 (N_2372,N_1540,N_1828);
or U2373 (N_2373,N_1845,N_1940);
nor U2374 (N_2374,N_1798,N_1976);
nand U2375 (N_2375,N_1816,N_1665);
nor U2376 (N_2376,N_1611,N_1624);
nor U2377 (N_2377,N_1819,N_1617);
nand U2378 (N_2378,N_1716,N_1977);
or U2379 (N_2379,N_1996,N_1877);
nand U2380 (N_2380,N_1891,N_1787);
or U2381 (N_2381,N_1869,N_1627);
nor U2382 (N_2382,N_1722,N_1534);
nor U2383 (N_2383,N_1548,N_1706);
or U2384 (N_2384,N_1621,N_1848);
nor U2385 (N_2385,N_1501,N_1789);
or U2386 (N_2386,N_1980,N_1518);
xor U2387 (N_2387,N_1536,N_1830);
nor U2388 (N_2388,N_1764,N_1732);
xnor U2389 (N_2389,N_1926,N_1543);
xor U2390 (N_2390,N_1992,N_1756);
and U2391 (N_2391,N_1564,N_1574);
nand U2392 (N_2392,N_1608,N_1553);
and U2393 (N_2393,N_1965,N_1824);
and U2394 (N_2394,N_1700,N_1761);
and U2395 (N_2395,N_1615,N_1757);
nor U2396 (N_2396,N_1573,N_1807);
or U2397 (N_2397,N_1830,N_1750);
and U2398 (N_2398,N_1514,N_1857);
nand U2399 (N_2399,N_1743,N_1886);
nand U2400 (N_2400,N_1707,N_1672);
or U2401 (N_2401,N_1888,N_1781);
nand U2402 (N_2402,N_1558,N_1724);
nand U2403 (N_2403,N_1766,N_1844);
nor U2404 (N_2404,N_1817,N_1602);
xnor U2405 (N_2405,N_1543,N_1930);
nand U2406 (N_2406,N_1572,N_1964);
and U2407 (N_2407,N_1727,N_1878);
and U2408 (N_2408,N_1786,N_1803);
and U2409 (N_2409,N_1619,N_1558);
xor U2410 (N_2410,N_1503,N_1964);
nor U2411 (N_2411,N_1647,N_1528);
nand U2412 (N_2412,N_1929,N_1761);
nand U2413 (N_2413,N_1935,N_1836);
nor U2414 (N_2414,N_1935,N_1633);
xor U2415 (N_2415,N_1748,N_1516);
nand U2416 (N_2416,N_1520,N_1701);
and U2417 (N_2417,N_1556,N_1535);
xor U2418 (N_2418,N_1803,N_1617);
or U2419 (N_2419,N_1572,N_1517);
xnor U2420 (N_2420,N_1752,N_1643);
xnor U2421 (N_2421,N_1550,N_1613);
nor U2422 (N_2422,N_1936,N_1793);
and U2423 (N_2423,N_1732,N_1659);
nor U2424 (N_2424,N_1929,N_1614);
and U2425 (N_2425,N_1909,N_1933);
and U2426 (N_2426,N_1680,N_1651);
xor U2427 (N_2427,N_1966,N_1668);
and U2428 (N_2428,N_1573,N_1658);
or U2429 (N_2429,N_1623,N_1696);
and U2430 (N_2430,N_1936,N_1905);
or U2431 (N_2431,N_1628,N_1774);
nor U2432 (N_2432,N_1928,N_1557);
xnor U2433 (N_2433,N_1934,N_1787);
and U2434 (N_2434,N_1861,N_1899);
or U2435 (N_2435,N_1814,N_1738);
or U2436 (N_2436,N_1976,N_1628);
xor U2437 (N_2437,N_1795,N_1755);
nor U2438 (N_2438,N_1777,N_1885);
nor U2439 (N_2439,N_1865,N_1763);
nor U2440 (N_2440,N_1535,N_1639);
and U2441 (N_2441,N_1985,N_1765);
nor U2442 (N_2442,N_1807,N_1938);
nor U2443 (N_2443,N_1977,N_1753);
nand U2444 (N_2444,N_1538,N_1789);
xnor U2445 (N_2445,N_1961,N_1699);
nor U2446 (N_2446,N_1719,N_1716);
xnor U2447 (N_2447,N_1595,N_1591);
xor U2448 (N_2448,N_1543,N_1527);
nand U2449 (N_2449,N_1523,N_1945);
and U2450 (N_2450,N_1987,N_1569);
and U2451 (N_2451,N_1693,N_1957);
nand U2452 (N_2452,N_1690,N_1802);
or U2453 (N_2453,N_1859,N_1670);
or U2454 (N_2454,N_1697,N_1638);
nor U2455 (N_2455,N_1773,N_1966);
or U2456 (N_2456,N_1643,N_1842);
or U2457 (N_2457,N_1541,N_1865);
nor U2458 (N_2458,N_1679,N_1657);
nor U2459 (N_2459,N_1580,N_1804);
nor U2460 (N_2460,N_1506,N_1529);
and U2461 (N_2461,N_1581,N_1851);
and U2462 (N_2462,N_1589,N_1875);
or U2463 (N_2463,N_1638,N_1503);
nand U2464 (N_2464,N_1661,N_1829);
xnor U2465 (N_2465,N_1626,N_1701);
and U2466 (N_2466,N_1738,N_1523);
xnor U2467 (N_2467,N_1660,N_1893);
and U2468 (N_2468,N_1965,N_1571);
nand U2469 (N_2469,N_1780,N_1928);
xnor U2470 (N_2470,N_1856,N_1675);
xor U2471 (N_2471,N_1644,N_1623);
and U2472 (N_2472,N_1771,N_1843);
and U2473 (N_2473,N_1986,N_1549);
or U2474 (N_2474,N_1735,N_1562);
nor U2475 (N_2475,N_1719,N_1547);
xnor U2476 (N_2476,N_1613,N_1908);
or U2477 (N_2477,N_1952,N_1504);
or U2478 (N_2478,N_1888,N_1928);
or U2479 (N_2479,N_1818,N_1656);
xor U2480 (N_2480,N_1849,N_1876);
or U2481 (N_2481,N_1741,N_1958);
nor U2482 (N_2482,N_1718,N_1565);
and U2483 (N_2483,N_1850,N_1622);
xnor U2484 (N_2484,N_1841,N_1586);
xnor U2485 (N_2485,N_1675,N_1908);
and U2486 (N_2486,N_1710,N_1935);
or U2487 (N_2487,N_1581,N_1822);
nor U2488 (N_2488,N_1751,N_1537);
and U2489 (N_2489,N_1861,N_1748);
xnor U2490 (N_2490,N_1557,N_1992);
nor U2491 (N_2491,N_1573,N_1748);
nand U2492 (N_2492,N_1516,N_1531);
and U2493 (N_2493,N_1500,N_1737);
nor U2494 (N_2494,N_1801,N_1742);
and U2495 (N_2495,N_1583,N_1632);
nor U2496 (N_2496,N_1653,N_1588);
nor U2497 (N_2497,N_1915,N_1984);
and U2498 (N_2498,N_1893,N_1908);
or U2499 (N_2499,N_1955,N_1991);
nor U2500 (N_2500,N_2361,N_2371);
nand U2501 (N_2501,N_2080,N_2155);
and U2502 (N_2502,N_2159,N_2052);
nand U2503 (N_2503,N_2026,N_2296);
xor U2504 (N_2504,N_2035,N_2477);
and U2505 (N_2505,N_2273,N_2334);
nand U2506 (N_2506,N_2187,N_2430);
or U2507 (N_2507,N_2185,N_2090);
nor U2508 (N_2508,N_2389,N_2454);
and U2509 (N_2509,N_2385,N_2332);
nor U2510 (N_2510,N_2231,N_2182);
or U2511 (N_2511,N_2481,N_2449);
or U2512 (N_2512,N_2151,N_2142);
nor U2513 (N_2513,N_2122,N_2276);
nor U2514 (N_2514,N_2176,N_2497);
nand U2515 (N_2515,N_2404,N_2260);
nor U2516 (N_2516,N_2222,N_2167);
and U2517 (N_2517,N_2432,N_2082);
and U2518 (N_2518,N_2165,N_2229);
xor U2519 (N_2519,N_2281,N_2275);
nand U2520 (N_2520,N_2403,N_2458);
nand U2521 (N_2521,N_2022,N_2425);
xnor U2522 (N_2522,N_2158,N_2189);
nand U2523 (N_2523,N_2311,N_2426);
nor U2524 (N_2524,N_2252,N_2417);
xor U2525 (N_2525,N_2150,N_2456);
and U2526 (N_2526,N_2320,N_2214);
nand U2527 (N_2527,N_2006,N_2140);
xor U2528 (N_2528,N_2435,N_2348);
nand U2529 (N_2529,N_2261,N_2094);
and U2530 (N_2530,N_2269,N_2408);
or U2531 (N_2531,N_2439,N_2009);
nor U2532 (N_2532,N_2305,N_2016);
and U2533 (N_2533,N_2444,N_2266);
or U2534 (N_2534,N_2415,N_2492);
and U2535 (N_2535,N_2490,N_2302);
xnor U2536 (N_2536,N_2085,N_2145);
xnor U2537 (N_2537,N_2431,N_2104);
nor U2538 (N_2538,N_2153,N_2205);
xnor U2539 (N_2539,N_2476,N_2154);
xor U2540 (N_2540,N_2183,N_2470);
nor U2541 (N_2541,N_2235,N_2363);
and U2542 (N_2542,N_2271,N_2148);
nor U2543 (N_2543,N_2097,N_2010);
or U2544 (N_2544,N_2460,N_2354);
nand U2545 (N_2545,N_2226,N_2466);
or U2546 (N_2546,N_2124,N_2023);
xnor U2547 (N_2547,N_2318,N_2463);
and U2548 (N_2548,N_2012,N_2491);
nor U2549 (N_2549,N_2342,N_2113);
nand U2550 (N_2550,N_2177,N_2228);
or U2551 (N_2551,N_2069,N_2230);
or U2552 (N_2552,N_2160,N_2381);
and U2553 (N_2553,N_2064,N_2411);
xor U2554 (N_2554,N_2208,N_2237);
or U2555 (N_2555,N_2060,N_2072);
xor U2556 (N_2556,N_2125,N_2393);
nand U2557 (N_2557,N_2129,N_2391);
xor U2558 (N_2558,N_2443,N_2055);
or U2559 (N_2559,N_2076,N_2001);
nand U2560 (N_2560,N_2420,N_2190);
and U2561 (N_2561,N_2327,N_2108);
nor U2562 (N_2562,N_2132,N_2002);
and U2563 (N_2563,N_2133,N_2347);
nand U2564 (N_2564,N_2288,N_2357);
and U2565 (N_2565,N_2286,N_2283);
xor U2566 (N_2566,N_2186,N_2173);
xor U2567 (N_2567,N_2204,N_2355);
and U2568 (N_2568,N_2496,N_2135);
xnor U2569 (N_2569,N_2073,N_2471);
or U2570 (N_2570,N_2114,N_2027);
nor U2571 (N_2571,N_2220,N_2370);
nand U2572 (N_2572,N_2191,N_2300);
or U2573 (N_2573,N_2171,N_2110);
and U2574 (N_2574,N_2074,N_2315);
xor U2575 (N_2575,N_2483,N_2079);
and U2576 (N_2576,N_2292,N_2268);
or U2577 (N_2577,N_2324,N_2303);
xor U2578 (N_2578,N_2170,N_2128);
nand U2579 (N_2579,N_2392,N_2067);
nand U2580 (N_2580,N_2083,N_2434);
or U2581 (N_2581,N_2338,N_2306);
nand U2582 (N_2582,N_2178,N_2089);
xnor U2583 (N_2583,N_2126,N_2298);
and U2584 (N_2584,N_2386,N_2337);
or U2585 (N_2585,N_2335,N_2467);
nor U2586 (N_2586,N_2330,N_2418);
nor U2587 (N_2587,N_2179,N_2419);
nand U2588 (N_2588,N_2345,N_2437);
nand U2589 (N_2589,N_2253,N_2096);
xnor U2590 (N_2590,N_2373,N_2499);
nand U2591 (N_2591,N_2141,N_2181);
xor U2592 (N_2592,N_2224,N_2464);
and U2593 (N_2593,N_2343,N_2336);
or U2594 (N_2594,N_2240,N_2028);
nor U2595 (N_2595,N_2485,N_2376);
and U2596 (N_2596,N_2484,N_2161);
and U2597 (N_2597,N_2003,N_2429);
nor U2598 (N_2598,N_2427,N_2211);
nor U2599 (N_2599,N_2087,N_2416);
nor U2600 (N_2600,N_2257,N_2319);
nand U2601 (N_2601,N_2441,N_2149);
nor U2602 (N_2602,N_2488,N_2207);
and U2603 (N_2603,N_2356,N_2317);
or U2604 (N_2604,N_2446,N_2007);
and U2605 (N_2605,N_2137,N_2465);
nand U2606 (N_2606,N_2424,N_2272);
and U2607 (N_2607,N_2047,N_2196);
xor U2608 (N_2608,N_2423,N_2369);
xor U2609 (N_2609,N_2455,N_2278);
nand U2610 (N_2610,N_2383,N_2015);
nor U2611 (N_2611,N_2130,N_2245);
xor U2612 (N_2612,N_2111,N_2127);
and U2613 (N_2613,N_2340,N_2041);
nand U2614 (N_2614,N_2368,N_2344);
nor U2615 (N_2615,N_2367,N_2071);
nand U2616 (N_2616,N_2310,N_2084);
and U2617 (N_2617,N_2285,N_2136);
nand U2618 (N_2618,N_2284,N_2213);
nor U2619 (N_2619,N_2495,N_2459);
nand U2620 (N_2620,N_2106,N_2445);
nand U2621 (N_2621,N_2279,N_2103);
and U2622 (N_2622,N_2414,N_2049);
and U2623 (N_2623,N_2174,N_2021);
xor U2624 (N_2624,N_2295,N_2120);
nor U2625 (N_2625,N_2221,N_2291);
xor U2626 (N_2626,N_2163,N_2390);
nand U2627 (N_2627,N_2099,N_2034);
and U2628 (N_2628,N_2293,N_2075);
and U2629 (N_2629,N_2061,N_2410);
xor U2630 (N_2630,N_2475,N_2013);
xor U2631 (N_2631,N_2197,N_2045);
or U2632 (N_2632,N_2143,N_2162);
nor U2633 (N_2633,N_2374,N_2402);
nand U2634 (N_2634,N_2290,N_2238);
xor U2635 (N_2635,N_2070,N_2109);
nand U2636 (N_2636,N_2056,N_2457);
and U2637 (N_2637,N_2025,N_2299);
nor U2638 (N_2638,N_2350,N_2452);
or U2639 (N_2639,N_2289,N_2146);
and U2640 (N_2640,N_2048,N_2428);
or U2641 (N_2641,N_2329,N_2473);
nor U2642 (N_2642,N_2262,N_2362);
nor U2643 (N_2643,N_2038,N_2387);
or U2644 (N_2644,N_2063,N_2400);
xnor U2645 (N_2645,N_2358,N_2321);
nand U2646 (N_2646,N_2379,N_2199);
nand U2647 (N_2647,N_2024,N_2494);
xnor U2648 (N_2648,N_2078,N_2037);
xor U2649 (N_2649,N_2353,N_2489);
xnor U2650 (N_2650,N_2123,N_2144);
nand U2651 (N_2651,N_2077,N_2031);
or U2652 (N_2652,N_2447,N_2019);
nor U2653 (N_2653,N_2346,N_2044);
and U2654 (N_2654,N_2264,N_2218);
nand U2655 (N_2655,N_2212,N_2407);
and U2656 (N_2656,N_2372,N_2131);
and U2657 (N_2657,N_2216,N_2206);
and U2658 (N_2658,N_2375,N_2487);
xnor U2659 (N_2659,N_2388,N_2217);
or U2660 (N_2660,N_2017,N_2088);
xor U2661 (N_2661,N_2313,N_2256);
and U2662 (N_2662,N_2394,N_2166);
nand U2663 (N_2663,N_2184,N_2051);
nand U2664 (N_2664,N_2192,N_2316);
nor U2665 (N_2665,N_2421,N_2198);
nand U2666 (N_2666,N_2223,N_2068);
xor U2667 (N_2667,N_2107,N_2210);
or U2668 (N_2668,N_2005,N_2307);
nand U2669 (N_2669,N_2092,N_2234);
nand U2670 (N_2670,N_2280,N_2247);
or U2671 (N_2671,N_2241,N_2134);
or U2672 (N_2672,N_2029,N_2039);
or U2673 (N_2673,N_2105,N_2472);
and U2674 (N_2674,N_2091,N_2117);
nor U2675 (N_2675,N_2479,N_2046);
nor U2676 (N_2676,N_2042,N_2239);
nand U2677 (N_2677,N_2004,N_2215);
or U2678 (N_2678,N_2040,N_2121);
nand U2679 (N_2679,N_2382,N_2011);
or U2680 (N_2680,N_2225,N_2246);
and U2681 (N_2681,N_2384,N_2095);
or U2682 (N_2682,N_2232,N_2498);
nand U2683 (N_2683,N_2265,N_2008);
nor U2684 (N_2684,N_2195,N_2282);
nor U2685 (N_2685,N_2274,N_2251);
or U2686 (N_2686,N_2249,N_2323);
xor U2687 (N_2687,N_2351,N_2202);
nand U2688 (N_2688,N_2364,N_2304);
xor U2689 (N_2689,N_2250,N_2469);
or U2690 (N_2690,N_2474,N_2325);
and U2691 (N_2691,N_2043,N_2312);
nand U2692 (N_2692,N_2438,N_2119);
xnor U2693 (N_2693,N_2462,N_2248);
or U2694 (N_2694,N_2209,N_2000);
nor U2695 (N_2695,N_2308,N_2433);
or U2696 (N_2696,N_2169,N_2243);
and U2697 (N_2697,N_2020,N_2062);
nor U2698 (N_2698,N_2294,N_2157);
or U2699 (N_2699,N_2254,N_2412);
xnor U2700 (N_2700,N_2339,N_2255);
and U2701 (N_2701,N_2065,N_2450);
xnor U2702 (N_2702,N_2233,N_2112);
nor U2703 (N_2703,N_2258,N_2395);
nor U2704 (N_2704,N_2328,N_2453);
nor U2705 (N_2705,N_2480,N_2396);
xor U2706 (N_2706,N_2309,N_2263);
nor U2707 (N_2707,N_2270,N_2314);
nand U2708 (N_2708,N_2359,N_2036);
nor U2709 (N_2709,N_2244,N_2018);
nand U2710 (N_2710,N_2333,N_2360);
and U2711 (N_2711,N_2448,N_2014);
and U2712 (N_2712,N_2050,N_2406);
or U2713 (N_2713,N_2482,N_2468);
or U2714 (N_2714,N_2236,N_2442);
or U2715 (N_2715,N_2352,N_2030);
nor U2716 (N_2716,N_2399,N_2301);
nor U2717 (N_2717,N_2053,N_2156);
xnor U2718 (N_2718,N_2398,N_2341);
nand U2719 (N_2719,N_2267,N_2147);
and U2720 (N_2720,N_2409,N_2377);
and U2721 (N_2721,N_2116,N_2201);
xnor U2722 (N_2722,N_2193,N_2366);
xor U2723 (N_2723,N_2413,N_2365);
xnor U2724 (N_2724,N_2138,N_2054);
xor U2725 (N_2725,N_2115,N_2378);
nand U2726 (N_2726,N_2331,N_2219);
nor U2727 (N_2727,N_2180,N_2277);
nand U2728 (N_2728,N_2405,N_2118);
nand U2729 (N_2729,N_2101,N_2172);
nor U2730 (N_2730,N_2259,N_2380);
nand U2731 (N_2731,N_2461,N_2057);
and U2732 (N_2732,N_2242,N_2436);
and U2733 (N_2733,N_2059,N_2164);
xnor U2734 (N_2734,N_2175,N_2033);
and U2735 (N_2735,N_2486,N_2287);
nand U2736 (N_2736,N_2493,N_2086);
nor U2737 (N_2737,N_2098,N_2397);
and U2738 (N_2738,N_2451,N_2168);
or U2739 (N_2739,N_2081,N_2152);
or U2740 (N_2740,N_2194,N_2401);
nor U2741 (N_2741,N_2032,N_2058);
nor U2742 (N_2742,N_2349,N_2203);
or U2743 (N_2743,N_2093,N_2200);
nand U2744 (N_2744,N_2422,N_2188);
nand U2745 (N_2745,N_2227,N_2102);
and U2746 (N_2746,N_2139,N_2066);
or U2747 (N_2747,N_2297,N_2326);
nand U2748 (N_2748,N_2440,N_2322);
and U2749 (N_2749,N_2478,N_2100);
nor U2750 (N_2750,N_2121,N_2182);
or U2751 (N_2751,N_2445,N_2368);
nor U2752 (N_2752,N_2360,N_2176);
nor U2753 (N_2753,N_2154,N_2331);
nand U2754 (N_2754,N_2373,N_2209);
xor U2755 (N_2755,N_2064,N_2243);
nor U2756 (N_2756,N_2431,N_2466);
xor U2757 (N_2757,N_2360,N_2364);
xor U2758 (N_2758,N_2187,N_2442);
nor U2759 (N_2759,N_2225,N_2025);
xor U2760 (N_2760,N_2452,N_2208);
nor U2761 (N_2761,N_2216,N_2301);
or U2762 (N_2762,N_2412,N_2351);
and U2763 (N_2763,N_2344,N_2064);
xnor U2764 (N_2764,N_2060,N_2360);
or U2765 (N_2765,N_2120,N_2156);
or U2766 (N_2766,N_2074,N_2005);
and U2767 (N_2767,N_2270,N_2148);
and U2768 (N_2768,N_2393,N_2417);
xnor U2769 (N_2769,N_2472,N_2415);
nor U2770 (N_2770,N_2045,N_2377);
nor U2771 (N_2771,N_2001,N_2269);
nor U2772 (N_2772,N_2495,N_2008);
and U2773 (N_2773,N_2263,N_2284);
xnor U2774 (N_2774,N_2212,N_2057);
or U2775 (N_2775,N_2227,N_2178);
and U2776 (N_2776,N_2490,N_2483);
nor U2777 (N_2777,N_2460,N_2494);
and U2778 (N_2778,N_2338,N_2359);
or U2779 (N_2779,N_2028,N_2253);
nor U2780 (N_2780,N_2244,N_2486);
xor U2781 (N_2781,N_2499,N_2086);
nand U2782 (N_2782,N_2263,N_2104);
and U2783 (N_2783,N_2375,N_2329);
xnor U2784 (N_2784,N_2349,N_2069);
xnor U2785 (N_2785,N_2160,N_2059);
or U2786 (N_2786,N_2302,N_2064);
and U2787 (N_2787,N_2219,N_2257);
xnor U2788 (N_2788,N_2210,N_2430);
or U2789 (N_2789,N_2410,N_2255);
nand U2790 (N_2790,N_2483,N_2192);
nor U2791 (N_2791,N_2231,N_2069);
xnor U2792 (N_2792,N_2032,N_2060);
nor U2793 (N_2793,N_2182,N_2240);
and U2794 (N_2794,N_2226,N_2147);
or U2795 (N_2795,N_2073,N_2257);
nor U2796 (N_2796,N_2000,N_2301);
xor U2797 (N_2797,N_2354,N_2377);
or U2798 (N_2798,N_2046,N_2299);
and U2799 (N_2799,N_2435,N_2382);
nand U2800 (N_2800,N_2216,N_2094);
or U2801 (N_2801,N_2063,N_2331);
nor U2802 (N_2802,N_2387,N_2273);
xnor U2803 (N_2803,N_2099,N_2025);
nand U2804 (N_2804,N_2137,N_2258);
nor U2805 (N_2805,N_2361,N_2117);
nor U2806 (N_2806,N_2362,N_2493);
and U2807 (N_2807,N_2001,N_2113);
xnor U2808 (N_2808,N_2441,N_2344);
or U2809 (N_2809,N_2410,N_2329);
xnor U2810 (N_2810,N_2244,N_2285);
and U2811 (N_2811,N_2324,N_2243);
or U2812 (N_2812,N_2473,N_2023);
or U2813 (N_2813,N_2017,N_2324);
nor U2814 (N_2814,N_2368,N_2387);
or U2815 (N_2815,N_2400,N_2288);
nor U2816 (N_2816,N_2388,N_2205);
nand U2817 (N_2817,N_2047,N_2180);
or U2818 (N_2818,N_2270,N_2176);
nand U2819 (N_2819,N_2187,N_2213);
and U2820 (N_2820,N_2280,N_2128);
xnor U2821 (N_2821,N_2281,N_2417);
nor U2822 (N_2822,N_2221,N_2154);
or U2823 (N_2823,N_2255,N_2347);
nand U2824 (N_2824,N_2474,N_2088);
nand U2825 (N_2825,N_2296,N_2098);
nor U2826 (N_2826,N_2099,N_2156);
and U2827 (N_2827,N_2088,N_2342);
and U2828 (N_2828,N_2397,N_2351);
xor U2829 (N_2829,N_2371,N_2340);
and U2830 (N_2830,N_2060,N_2316);
nor U2831 (N_2831,N_2231,N_2145);
xnor U2832 (N_2832,N_2126,N_2193);
or U2833 (N_2833,N_2363,N_2134);
or U2834 (N_2834,N_2138,N_2098);
nand U2835 (N_2835,N_2259,N_2422);
or U2836 (N_2836,N_2357,N_2290);
nand U2837 (N_2837,N_2061,N_2236);
nand U2838 (N_2838,N_2363,N_2431);
nand U2839 (N_2839,N_2196,N_2407);
nor U2840 (N_2840,N_2261,N_2097);
and U2841 (N_2841,N_2091,N_2239);
nand U2842 (N_2842,N_2289,N_2414);
or U2843 (N_2843,N_2300,N_2143);
xnor U2844 (N_2844,N_2318,N_2163);
or U2845 (N_2845,N_2485,N_2084);
nand U2846 (N_2846,N_2305,N_2445);
xor U2847 (N_2847,N_2103,N_2285);
nand U2848 (N_2848,N_2125,N_2072);
nand U2849 (N_2849,N_2010,N_2030);
nor U2850 (N_2850,N_2442,N_2408);
nor U2851 (N_2851,N_2214,N_2070);
xor U2852 (N_2852,N_2124,N_2423);
or U2853 (N_2853,N_2411,N_2059);
and U2854 (N_2854,N_2398,N_2322);
or U2855 (N_2855,N_2419,N_2259);
nand U2856 (N_2856,N_2018,N_2359);
xor U2857 (N_2857,N_2405,N_2456);
nor U2858 (N_2858,N_2304,N_2018);
and U2859 (N_2859,N_2015,N_2074);
or U2860 (N_2860,N_2485,N_2074);
nand U2861 (N_2861,N_2458,N_2211);
and U2862 (N_2862,N_2448,N_2355);
nand U2863 (N_2863,N_2285,N_2027);
and U2864 (N_2864,N_2097,N_2352);
or U2865 (N_2865,N_2295,N_2217);
and U2866 (N_2866,N_2388,N_2107);
nor U2867 (N_2867,N_2419,N_2216);
nor U2868 (N_2868,N_2213,N_2030);
nor U2869 (N_2869,N_2224,N_2310);
or U2870 (N_2870,N_2225,N_2250);
nand U2871 (N_2871,N_2053,N_2007);
and U2872 (N_2872,N_2438,N_2282);
nor U2873 (N_2873,N_2148,N_2490);
or U2874 (N_2874,N_2334,N_2200);
nand U2875 (N_2875,N_2222,N_2430);
xor U2876 (N_2876,N_2449,N_2152);
nor U2877 (N_2877,N_2057,N_2447);
and U2878 (N_2878,N_2441,N_2278);
nor U2879 (N_2879,N_2097,N_2015);
xnor U2880 (N_2880,N_2207,N_2253);
xnor U2881 (N_2881,N_2453,N_2471);
xor U2882 (N_2882,N_2267,N_2418);
nand U2883 (N_2883,N_2134,N_2027);
nand U2884 (N_2884,N_2436,N_2309);
and U2885 (N_2885,N_2272,N_2301);
and U2886 (N_2886,N_2381,N_2057);
xnor U2887 (N_2887,N_2034,N_2292);
or U2888 (N_2888,N_2139,N_2436);
xnor U2889 (N_2889,N_2102,N_2246);
or U2890 (N_2890,N_2420,N_2209);
xnor U2891 (N_2891,N_2002,N_2022);
and U2892 (N_2892,N_2411,N_2090);
nor U2893 (N_2893,N_2417,N_2073);
nor U2894 (N_2894,N_2427,N_2240);
or U2895 (N_2895,N_2117,N_2044);
nor U2896 (N_2896,N_2045,N_2273);
and U2897 (N_2897,N_2254,N_2357);
nand U2898 (N_2898,N_2061,N_2435);
and U2899 (N_2899,N_2305,N_2238);
xor U2900 (N_2900,N_2110,N_2184);
xnor U2901 (N_2901,N_2415,N_2153);
or U2902 (N_2902,N_2350,N_2205);
nand U2903 (N_2903,N_2108,N_2116);
xnor U2904 (N_2904,N_2005,N_2026);
and U2905 (N_2905,N_2042,N_2309);
nand U2906 (N_2906,N_2094,N_2204);
nand U2907 (N_2907,N_2085,N_2486);
and U2908 (N_2908,N_2240,N_2193);
and U2909 (N_2909,N_2084,N_2381);
and U2910 (N_2910,N_2207,N_2252);
nand U2911 (N_2911,N_2003,N_2233);
nor U2912 (N_2912,N_2104,N_2233);
and U2913 (N_2913,N_2091,N_2330);
xor U2914 (N_2914,N_2478,N_2302);
nor U2915 (N_2915,N_2200,N_2498);
xor U2916 (N_2916,N_2091,N_2464);
nor U2917 (N_2917,N_2386,N_2452);
and U2918 (N_2918,N_2235,N_2202);
or U2919 (N_2919,N_2344,N_2000);
nand U2920 (N_2920,N_2094,N_2434);
xnor U2921 (N_2921,N_2402,N_2495);
nand U2922 (N_2922,N_2435,N_2163);
and U2923 (N_2923,N_2146,N_2222);
and U2924 (N_2924,N_2006,N_2022);
and U2925 (N_2925,N_2165,N_2265);
nand U2926 (N_2926,N_2141,N_2136);
and U2927 (N_2927,N_2033,N_2468);
nand U2928 (N_2928,N_2251,N_2414);
nor U2929 (N_2929,N_2225,N_2309);
nor U2930 (N_2930,N_2311,N_2000);
nand U2931 (N_2931,N_2266,N_2159);
and U2932 (N_2932,N_2384,N_2190);
nor U2933 (N_2933,N_2388,N_2417);
xor U2934 (N_2934,N_2162,N_2126);
and U2935 (N_2935,N_2356,N_2411);
xnor U2936 (N_2936,N_2221,N_2432);
nor U2937 (N_2937,N_2245,N_2370);
nand U2938 (N_2938,N_2409,N_2111);
nor U2939 (N_2939,N_2279,N_2492);
or U2940 (N_2940,N_2056,N_2084);
and U2941 (N_2941,N_2163,N_2181);
xnor U2942 (N_2942,N_2200,N_2106);
or U2943 (N_2943,N_2383,N_2189);
nor U2944 (N_2944,N_2348,N_2313);
xnor U2945 (N_2945,N_2244,N_2033);
or U2946 (N_2946,N_2244,N_2301);
nand U2947 (N_2947,N_2146,N_2440);
nor U2948 (N_2948,N_2285,N_2242);
xor U2949 (N_2949,N_2272,N_2189);
nand U2950 (N_2950,N_2320,N_2139);
xnor U2951 (N_2951,N_2151,N_2408);
nor U2952 (N_2952,N_2333,N_2198);
xor U2953 (N_2953,N_2009,N_2258);
nor U2954 (N_2954,N_2388,N_2414);
and U2955 (N_2955,N_2363,N_2018);
and U2956 (N_2956,N_2373,N_2058);
and U2957 (N_2957,N_2374,N_2410);
and U2958 (N_2958,N_2399,N_2494);
nor U2959 (N_2959,N_2236,N_2403);
nor U2960 (N_2960,N_2377,N_2279);
nor U2961 (N_2961,N_2216,N_2350);
nand U2962 (N_2962,N_2412,N_2305);
xnor U2963 (N_2963,N_2078,N_2180);
xnor U2964 (N_2964,N_2218,N_2219);
nor U2965 (N_2965,N_2406,N_2158);
nor U2966 (N_2966,N_2362,N_2059);
nand U2967 (N_2967,N_2308,N_2494);
or U2968 (N_2968,N_2046,N_2473);
and U2969 (N_2969,N_2310,N_2128);
xor U2970 (N_2970,N_2290,N_2149);
xnor U2971 (N_2971,N_2023,N_2372);
nand U2972 (N_2972,N_2409,N_2394);
xor U2973 (N_2973,N_2121,N_2352);
or U2974 (N_2974,N_2255,N_2291);
and U2975 (N_2975,N_2276,N_2308);
or U2976 (N_2976,N_2079,N_2074);
nand U2977 (N_2977,N_2033,N_2473);
and U2978 (N_2978,N_2340,N_2429);
and U2979 (N_2979,N_2426,N_2254);
xor U2980 (N_2980,N_2316,N_2215);
nor U2981 (N_2981,N_2326,N_2135);
xor U2982 (N_2982,N_2498,N_2298);
and U2983 (N_2983,N_2307,N_2021);
nor U2984 (N_2984,N_2323,N_2070);
xor U2985 (N_2985,N_2139,N_2459);
xor U2986 (N_2986,N_2231,N_2213);
xor U2987 (N_2987,N_2368,N_2098);
nand U2988 (N_2988,N_2345,N_2194);
xor U2989 (N_2989,N_2400,N_2120);
xor U2990 (N_2990,N_2484,N_2233);
and U2991 (N_2991,N_2300,N_2282);
or U2992 (N_2992,N_2185,N_2056);
nor U2993 (N_2993,N_2306,N_2145);
nand U2994 (N_2994,N_2268,N_2496);
nand U2995 (N_2995,N_2482,N_2254);
nand U2996 (N_2996,N_2392,N_2411);
nor U2997 (N_2997,N_2279,N_2308);
xnor U2998 (N_2998,N_2426,N_2221);
nor U2999 (N_2999,N_2127,N_2148);
xnor U3000 (N_3000,N_2741,N_2920);
nor U3001 (N_3001,N_2719,N_2974);
xnor U3002 (N_3002,N_2911,N_2569);
nor U3003 (N_3003,N_2626,N_2971);
and U3004 (N_3004,N_2688,N_2993);
nand U3005 (N_3005,N_2597,N_2686);
nand U3006 (N_3006,N_2854,N_2750);
nand U3007 (N_3007,N_2759,N_2636);
and U3008 (N_3008,N_2559,N_2812);
or U3009 (N_3009,N_2892,N_2737);
nor U3010 (N_3010,N_2962,N_2834);
or U3011 (N_3011,N_2868,N_2501);
nor U3012 (N_3012,N_2613,N_2599);
or U3013 (N_3013,N_2745,N_2964);
xor U3014 (N_3014,N_2878,N_2988);
nand U3015 (N_3015,N_2815,N_2940);
xnor U3016 (N_3016,N_2680,N_2886);
nor U3017 (N_3017,N_2554,N_2939);
nor U3018 (N_3018,N_2508,N_2588);
and U3019 (N_3019,N_2943,N_2735);
or U3020 (N_3020,N_2604,N_2879);
nor U3021 (N_3021,N_2792,N_2596);
xnor U3022 (N_3022,N_2984,N_2823);
or U3023 (N_3023,N_2773,N_2534);
and U3024 (N_3024,N_2506,N_2934);
and U3025 (N_3025,N_2820,N_2980);
xor U3026 (N_3026,N_2789,N_2744);
xor U3027 (N_3027,N_2727,N_2708);
nor U3028 (N_3028,N_2654,N_2638);
xnor U3029 (N_3029,N_2632,N_2647);
nor U3030 (N_3030,N_2749,N_2994);
nor U3031 (N_3031,N_2998,N_2548);
nand U3032 (N_3032,N_2997,N_2866);
and U3033 (N_3033,N_2517,N_2793);
xnor U3034 (N_3034,N_2702,N_2504);
and U3035 (N_3035,N_2657,N_2844);
and U3036 (N_3036,N_2772,N_2965);
and U3037 (N_3037,N_2571,N_2500);
xnor U3038 (N_3038,N_2952,N_2583);
or U3039 (N_3039,N_2894,N_2676);
xor U3040 (N_3040,N_2992,N_2848);
xor U3041 (N_3041,N_2828,N_2889);
nor U3042 (N_3042,N_2845,N_2610);
xor U3043 (N_3043,N_2864,N_2600);
nand U3044 (N_3044,N_2849,N_2594);
and U3045 (N_3045,N_2796,N_2774);
nand U3046 (N_3046,N_2639,N_2612);
xor U3047 (N_3047,N_2584,N_2785);
or U3048 (N_3048,N_2621,N_2936);
xnor U3049 (N_3049,N_2557,N_2635);
nand U3050 (N_3050,N_2855,N_2935);
nand U3051 (N_3051,N_2549,N_2665);
nand U3052 (N_3052,N_2752,N_2701);
nor U3053 (N_3053,N_2509,N_2528);
nand U3054 (N_3054,N_2819,N_2555);
or U3055 (N_3055,N_2837,N_2558);
xor U3056 (N_3056,N_2954,N_2606);
nand U3057 (N_3057,N_2563,N_2803);
or U3058 (N_3058,N_2924,N_2995);
or U3059 (N_3059,N_2822,N_2732);
and U3060 (N_3060,N_2693,N_2791);
or U3061 (N_3061,N_2870,N_2628);
nand U3062 (N_3062,N_2533,N_2843);
and U3063 (N_3063,N_2725,N_2546);
xnor U3064 (N_3064,N_2857,N_2768);
nor U3065 (N_3065,N_2957,N_2836);
nor U3066 (N_3066,N_2991,N_2776);
nand U3067 (N_3067,N_2897,N_2784);
or U3068 (N_3068,N_2687,N_2798);
xnor U3069 (N_3069,N_2841,N_2713);
nand U3070 (N_3070,N_2721,N_2830);
or U3071 (N_3071,N_2757,N_2532);
xor U3072 (N_3072,N_2909,N_2592);
nor U3073 (N_3073,N_2705,N_2805);
and U3074 (N_3074,N_2802,N_2541);
nor U3075 (N_3075,N_2529,N_2896);
nand U3076 (N_3076,N_2675,N_2524);
or U3077 (N_3077,N_2761,N_2914);
or U3078 (N_3078,N_2955,N_2564);
xnor U3079 (N_3079,N_2967,N_2511);
nand U3080 (N_3080,N_2671,N_2673);
nor U3081 (N_3081,N_2543,N_2656);
nand U3082 (N_3082,N_2574,N_2905);
nand U3083 (N_3083,N_2523,N_2751);
nor U3084 (N_3084,N_2601,N_2666);
or U3085 (N_3085,N_2824,N_2779);
and U3086 (N_3086,N_2891,N_2888);
nand U3087 (N_3087,N_2514,N_2882);
or U3088 (N_3088,N_2781,N_2522);
or U3089 (N_3089,N_2743,N_2706);
or U3090 (N_3090,N_2865,N_2641);
and U3091 (N_3091,N_2717,N_2758);
or U3092 (N_3092,N_2832,N_2790);
or U3093 (N_3093,N_2607,N_2513);
xnor U3094 (N_3094,N_2893,N_2724);
nor U3095 (N_3095,N_2556,N_2949);
xor U3096 (N_3096,N_2672,N_2970);
nand U3097 (N_3097,N_2748,N_2609);
and U3098 (N_3098,N_2747,N_2561);
and U3099 (N_3099,N_2975,N_2567);
and U3100 (N_3100,N_2778,N_2674);
nor U3101 (N_3101,N_2867,N_2679);
or U3102 (N_3102,N_2763,N_2869);
nand U3103 (N_3103,N_2566,N_2731);
or U3104 (N_3104,N_2589,N_2503);
nor U3105 (N_3105,N_2512,N_2651);
xnor U3106 (N_3106,N_2806,N_2821);
and U3107 (N_3107,N_2616,N_2655);
and U3108 (N_3108,N_2862,N_2510);
nand U3109 (N_3109,N_2932,N_2930);
nor U3110 (N_3110,N_2907,N_2746);
xor U3111 (N_3111,N_2578,N_2950);
or U3112 (N_3112,N_2903,N_2807);
or U3113 (N_3113,N_2712,N_2643);
nand U3114 (N_3114,N_2931,N_2895);
or U3115 (N_3115,N_2987,N_2579);
nor U3116 (N_3116,N_2608,N_2670);
or U3117 (N_3117,N_2729,N_2525);
xnor U3118 (N_3118,N_2720,N_2756);
or U3119 (N_3119,N_2577,N_2826);
or U3120 (N_3120,N_2788,N_2620);
or U3121 (N_3121,N_2944,N_2669);
and U3122 (N_3122,N_2945,N_2718);
nand U3123 (N_3123,N_2703,N_2769);
nand U3124 (N_3124,N_2733,N_2538);
nor U3125 (N_3125,N_2794,N_2644);
nor U3126 (N_3126,N_2692,N_2780);
or U3127 (N_3127,N_2661,N_2921);
or U3128 (N_3128,N_2694,N_2838);
and U3129 (N_3129,N_2775,N_2540);
or U3130 (N_3130,N_2782,N_2923);
nor U3131 (N_3131,N_2753,N_2710);
and U3132 (N_3132,N_2715,N_2709);
nand U3133 (N_3133,N_2922,N_2919);
and U3134 (N_3134,N_2716,N_2736);
or U3135 (N_3135,N_2652,N_2829);
and U3136 (N_3136,N_2981,N_2633);
xor U3137 (N_3137,N_2851,N_2831);
nand U3138 (N_3138,N_2850,N_2691);
or U3139 (N_3139,N_2552,N_2799);
xor U3140 (N_3140,N_2697,N_2734);
or U3141 (N_3141,N_2625,N_2738);
xnor U3142 (N_3142,N_2978,N_2972);
nand U3143 (N_3143,N_2999,N_2797);
nand U3144 (N_3144,N_2764,N_2827);
nor U3145 (N_3145,N_2875,N_2990);
and U3146 (N_3146,N_2890,N_2518);
nand U3147 (N_3147,N_2704,N_2659);
nand U3148 (N_3148,N_2842,N_2912);
or U3149 (N_3149,N_2618,N_2969);
xnor U3150 (N_3150,N_2526,N_2904);
or U3151 (N_3151,N_2804,N_2877);
xnor U3152 (N_3152,N_2976,N_2948);
and U3153 (N_3153,N_2539,N_2739);
xor U3154 (N_3154,N_2565,N_2668);
or U3155 (N_3155,N_2861,N_2953);
nor U3156 (N_3156,N_2873,N_2622);
and U3157 (N_3157,N_2614,N_2595);
nand U3158 (N_3158,N_2960,N_2951);
nor U3159 (N_3159,N_2853,N_2572);
nor U3160 (N_3160,N_2591,N_2617);
nand U3161 (N_3161,N_2650,N_2576);
nand U3162 (N_3162,N_2928,N_2913);
nand U3163 (N_3163,N_2629,N_2726);
or U3164 (N_3164,N_2887,N_2536);
xor U3165 (N_3165,N_2663,N_2929);
nand U3166 (N_3166,N_2839,N_2570);
nand U3167 (N_3167,N_2917,N_2695);
or U3168 (N_3168,N_2956,N_2770);
nor U3169 (N_3169,N_2902,N_2553);
nor U3170 (N_3170,N_2544,N_2593);
nor U3171 (N_3171,N_2947,N_2966);
xnor U3172 (N_3172,N_2550,N_2901);
xnor U3173 (N_3173,N_2690,N_2634);
xor U3174 (N_3174,N_2925,N_2860);
nor U3175 (N_3175,N_2627,N_2927);
nor U3176 (N_3176,N_2985,N_2884);
nand U3177 (N_3177,N_2664,N_2783);
nand U3178 (N_3178,N_2502,N_2642);
nor U3179 (N_3179,N_2640,N_2810);
xor U3180 (N_3180,N_2547,N_2847);
or U3181 (N_3181,N_2730,N_2722);
xnor U3182 (N_3182,N_2937,N_2871);
xnor U3183 (N_3183,N_2602,N_2881);
or U3184 (N_3184,N_2562,N_2938);
xnor U3185 (N_3185,N_2908,N_2700);
or U3186 (N_3186,N_2840,N_2667);
and U3187 (N_3187,N_2637,N_2863);
nand U3188 (N_3188,N_2814,N_2515);
or U3189 (N_3189,N_2916,N_2977);
nor U3190 (N_3190,N_2505,N_2958);
nand U3191 (N_3191,N_2816,N_2885);
xor U3192 (N_3192,N_2520,N_2542);
or U3193 (N_3193,N_2615,N_2575);
or U3194 (N_3194,N_2959,N_2619);
xor U3195 (N_3195,N_2968,N_2982);
nand U3196 (N_3196,N_2899,N_2689);
or U3197 (N_3197,N_2811,N_2624);
or U3198 (N_3198,N_2762,N_2590);
nor U3199 (N_3199,N_2683,N_2531);
and U3200 (N_3200,N_2699,N_2755);
or U3201 (N_3201,N_2516,N_2986);
and U3202 (N_3202,N_2817,N_2519);
nor U3203 (N_3203,N_2587,N_2535);
nor U3204 (N_3204,N_2646,N_2818);
xnor U3205 (N_3205,N_2833,N_2623);
xor U3206 (N_3206,N_2537,N_2649);
or U3207 (N_3207,N_2711,N_2906);
xor U3208 (N_3208,N_2545,N_2801);
xnor U3209 (N_3209,N_2918,N_2560);
xnor U3210 (N_3210,N_2898,N_2723);
nor U3211 (N_3211,N_2777,N_2876);
xor U3212 (N_3212,N_2527,N_2800);
nor U3213 (N_3213,N_2631,N_2989);
and U3214 (N_3214,N_2787,N_2900);
nand U3215 (N_3215,N_2915,N_2581);
or U3216 (N_3216,N_2660,N_2714);
xnor U3217 (N_3217,N_2825,N_2611);
and U3218 (N_3218,N_2698,N_2973);
and U3219 (N_3219,N_2933,N_2852);
xor U3220 (N_3220,N_2813,N_2910);
xor U3221 (N_3221,N_2681,N_2585);
xor U3222 (N_3222,N_2765,N_2605);
nor U3223 (N_3223,N_2760,N_2979);
and U3224 (N_3224,N_2586,N_2961);
or U3225 (N_3225,N_2767,N_2926);
nor U3226 (N_3226,N_2880,N_2786);
or U3227 (N_3227,N_2568,N_2603);
xor U3228 (N_3228,N_2809,N_2771);
nand U3229 (N_3229,N_2846,N_2658);
nor U3230 (N_3230,N_2707,N_2872);
and U3231 (N_3231,N_2941,N_2754);
nand U3232 (N_3232,N_2728,N_2874);
or U3233 (N_3233,N_2507,N_2996);
xor U3234 (N_3234,N_2653,N_2808);
nand U3235 (N_3235,N_2580,N_2835);
nand U3236 (N_3236,N_2859,N_2983);
nor U3237 (N_3237,N_2742,N_2645);
nor U3238 (N_3238,N_2963,N_2766);
or U3239 (N_3239,N_2942,N_2521);
nand U3240 (N_3240,N_2946,N_2573);
or U3241 (N_3241,N_2648,N_2530);
nand U3242 (N_3242,N_2883,N_2630);
or U3243 (N_3243,N_2696,N_2551);
nand U3244 (N_3244,N_2682,N_2582);
or U3245 (N_3245,N_2856,N_2598);
and U3246 (N_3246,N_2662,N_2858);
nor U3247 (N_3247,N_2677,N_2685);
nor U3248 (N_3248,N_2740,N_2678);
or U3249 (N_3249,N_2795,N_2684);
nand U3250 (N_3250,N_2713,N_2749);
and U3251 (N_3251,N_2909,N_2822);
or U3252 (N_3252,N_2529,N_2805);
nand U3253 (N_3253,N_2888,N_2829);
nor U3254 (N_3254,N_2514,N_2538);
or U3255 (N_3255,N_2690,N_2843);
or U3256 (N_3256,N_2542,N_2652);
or U3257 (N_3257,N_2516,N_2982);
and U3258 (N_3258,N_2727,N_2908);
xor U3259 (N_3259,N_2973,N_2765);
nand U3260 (N_3260,N_2944,N_2919);
xor U3261 (N_3261,N_2722,N_2698);
nand U3262 (N_3262,N_2529,N_2585);
nand U3263 (N_3263,N_2728,N_2658);
nor U3264 (N_3264,N_2734,N_2714);
nor U3265 (N_3265,N_2934,N_2732);
and U3266 (N_3266,N_2614,N_2629);
nand U3267 (N_3267,N_2678,N_2852);
and U3268 (N_3268,N_2741,N_2817);
xnor U3269 (N_3269,N_2919,N_2905);
nor U3270 (N_3270,N_2591,N_2797);
xor U3271 (N_3271,N_2602,N_2890);
nor U3272 (N_3272,N_2697,N_2528);
and U3273 (N_3273,N_2864,N_2941);
nor U3274 (N_3274,N_2688,N_2787);
xor U3275 (N_3275,N_2685,N_2784);
and U3276 (N_3276,N_2699,N_2923);
nor U3277 (N_3277,N_2643,N_2544);
xor U3278 (N_3278,N_2630,N_2696);
nor U3279 (N_3279,N_2743,N_2540);
or U3280 (N_3280,N_2502,N_2510);
or U3281 (N_3281,N_2854,N_2550);
and U3282 (N_3282,N_2677,N_2782);
or U3283 (N_3283,N_2987,N_2515);
or U3284 (N_3284,N_2848,N_2602);
nor U3285 (N_3285,N_2577,N_2937);
xnor U3286 (N_3286,N_2581,N_2554);
nor U3287 (N_3287,N_2733,N_2916);
or U3288 (N_3288,N_2669,N_2941);
nand U3289 (N_3289,N_2597,N_2735);
nand U3290 (N_3290,N_2758,N_2752);
nor U3291 (N_3291,N_2726,N_2546);
and U3292 (N_3292,N_2522,N_2971);
or U3293 (N_3293,N_2710,N_2659);
and U3294 (N_3294,N_2859,N_2510);
nand U3295 (N_3295,N_2682,N_2788);
or U3296 (N_3296,N_2750,N_2994);
nand U3297 (N_3297,N_2911,N_2869);
or U3298 (N_3298,N_2718,N_2888);
nand U3299 (N_3299,N_2532,N_2533);
and U3300 (N_3300,N_2584,N_2811);
xor U3301 (N_3301,N_2848,N_2689);
and U3302 (N_3302,N_2780,N_2769);
nor U3303 (N_3303,N_2620,N_2798);
and U3304 (N_3304,N_2896,N_2944);
nand U3305 (N_3305,N_2836,N_2746);
nand U3306 (N_3306,N_2601,N_2927);
nand U3307 (N_3307,N_2805,N_2598);
xnor U3308 (N_3308,N_2950,N_2603);
nand U3309 (N_3309,N_2807,N_2853);
nor U3310 (N_3310,N_2619,N_2929);
nand U3311 (N_3311,N_2881,N_2965);
nor U3312 (N_3312,N_2734,N_2651);
nor U3313 (N_3313,N_2734,N_2758);
nor U3314 (N_3314,N_2569,N_2956);
or U3315 (N_3315,N_2951,N_2523);
and U3316 (N_3316,N_2848,N_2535);
and U3317 (N_3317,N_2815,N_2935);
xnor U3318 (N_3318,N_2746,N_2624);
nand U3319 (N_3319,N_2664,N_2998);
or U3320 (N_3320,N_2579,N_2933);
nand U3321 (N_3321,N_2946,N_2549);
nand U3322 (N_3322,N_2569,N_2929);
nand U3323 (N_3323,N_2618,N_2846);
and U3324 (N_3324,N_2557,N_2642);
nand U3325 (N_3325,N_2808,N_2530);
nand U3326 (N_3326,N_2870,N_2710);
or U3327 (N_3327,N_2779,N_2895);
nor U3328 (N_3328,N_2833,N_2651);
or U3329 (N_3329,N_2828,N_2982);
and U3330 (N_3330,N_2918,N_2551);
nor U3331 (N_3331,N_2981,N_2731);
xor U3332 (N_3332,N_2971,N_2936);
xnor U3333 (N_3333,N_2842,N_2859);
or U3334 (N_3334,N_2756,N_2767);
and U3335 (N_3335,N_2718,N_2859);
and U3336 (N_3336,N_2651,N_2971);
or U3337 (N_3337,N_2618,N_2870);
nor U3338 (N_3338,N_2992,N_2775);
xor U3339 (N_3339,N_2655,N_2920);
nand U3340 (N_3340,N_2624,N_2626);
xor U3341 (N_3341,N_2854,N_2965);
or U3342 (N_3342,N_2786,N_2682);
nor U3343 (N_3343,N_2850,N_2879);
nor U3344 (N_3344,N_2808,N_2960);
nand U3345 (N_3345,N_2502,N_2773);
and U3346 (N_3346,N_2553,N_2587);
xor U3347 (N_3347,N_2692,N_2675);
or U3348 (N_3348,N_2763,N_2772);
nand U3349 (N_3349,N_2914,N_2537);
nor U3350 (N_3350,N_2615,N_2624);
or U3351 (N_3351,N_2745,N_2618);
xor U3352 (N_3352,N_2941,N_2698);
or U3353 (N_3353,N_2958,N_2580);
and U3354 (N_3354,N_2880,N_2549);
nand U3355 (N_3355,N_2934,N_2513);
or U3356 (N_3356,N_2894,N_2911);
or U3357 (N_3357,N_2774,N_2853);
nor U3358 (N_3358,N_2528,N_2789);
nor U3359 (N_3359,N_2697,N_2973);
nand U3360 (N_3360,N_2802,N_2909);
and U3361 (N_3361,N_2761,N_2922);
nor U3362 (N_3362,N_2627,N_2560);
xor U3363 (N_3363,N_2670,N_2823);
nor U3364 (N_3364,N_2908,N_2976);
nor U3365 (N_3365,N_2801,N_2637);
or U3366 (N_3366,N_2525,N_2636);
and U3367 (N_3367,N_2637,N_2640);
nor U3368 (N_3368,N_2990,N_2806);
or U3369 (N_3369,N_2888,N_2965);
or U3370 (N_3370,N_2839,N_2539);
nor U3371 (N_3371,N_2847,N_2574);
nor U3372 (N_3372,N_2913,N_2573);
nand U3373 (N_3373,N_2972,N_2778);
and U3374 (N_3374,N_2830,N_2623);
nand U3375 (N_3375,N_2600,N_2752);
or U3376 (N_3376,N_2702,N_2979);
nor U3377 (N_3377,N_2868,N_2794);
nor U3378 (N_3378,N_2967,N_2937);
nand U3379 (N_3379,N_2520,N_2579);
and U3380 (N_3380,N_2518,N_2967);
or U3381 (N_3381,N_2656,N_2929);
or U3382 (N_3382,N_2993,N_2822);
or U3383 (N_3383,N_2700,N_2822);
nand U3384 (N_3384,N_2550,N_2513);
nand U3385 (N_3385,N_2532,N_2776);
nand U3386 (N_3386,N_2907,N_2987);
xor U3387 (N_3387,N_2973,N_2746);
nor U3388 (N_3388,N_2916,N_2778);
nor U3389 (N_3389,N_2965,N_2898);
nand U3390 (N_3390,N_2588,N_2534);
or U3391 (N_3391,N_2696,N_2979);
or U3392 (N_3392,N_2521,N_2765);
xnor U3393 (N_3393,N_2531,N_2908);
and U3394 (N_3394,N_2579,N_2596);
or U3395 (N_3395,N_2567,N_2798);
nor U3396 (N_3396,N_2602,N_2904);
nand U3397 (N_3397,N_2966,N_2860);
nand U3398 (N_3398,N_2649,N_2510);
nand U3399 (N_3399,N_2533,N_2933);
nor U3400 (N_3400,N_2997,N_2604);
nor U3401 (N_3401,N_2615,N_2838);
xnor U3402 (N_3402,N_2855,N_2693);
or U3403 (N_3403,N_2719,N_2786);
nand U3404 (N_3404,N_2674,N_2872);
and U3405 (N_3405,N_2759,N_2978);
and U3406 (N_3406,N_2629,N_2501);
or U3407 (N_3407,N_2506,N_2713);
and U3408 (N_3408,N_2755,N_2771);
nand U3409 (N_3409,N_2847,N_2661);
nor U3410 (N_3410,N_2811,N_2816);
or U3411 (N_3411,N_2781,N_2623);
nand U3412 (N_3412,N_2626,N_2693);
nand U3413 (N_3413,N_2736,N_2986);
nor U3414 (N_3414,N_2945,N_2870);
or U3415 (N_3415,N_2730,N_2529);
nand U3416 (N_3416,N_2778,N_2618);
nand U3417 (N_3417,N_2528,N_2770);
xnor U3418 (N_3418,N_2642,N_2539);
or U3419 (N_3419,N_2577,N_2688);
nor U3420 (N_3420,N_2890,N_2522);
nand U3421 (N_3421,N_2787,N_2871);
xnor U3422 (N_3422,N_2943,N_2733);
nor U3423 (N_3423,N_2634,N_2568);
nand U3424 (N_3424,N_2791,N_2893);
and U3425 (N_3425,N_2960,N_2906);
xnor U3426 (N_3426,N_2526,N_2574);
nand U3427 (N_3427,N_2921,N_2950);
nand U3428 (N_3428,N_2982,N_2881);
nand U3429 (N_3429,N_2535,N_2897);
nor U3430 (N_3430,N_2737,N_2700);
and U3431 (N_3431,N_2864,N_2984);
nor U3432 (N_3432,N_2853,N_2517);
nor U3433 (N_3433,N_2589,N_2737);
xnor U3434 (N_3434,N_2790,N_2954);
nand U3435 (N_3435,N_2985,N_2667);
xnor U3436 (N_3436,N_2711,N_2865);
nand U3437 (N_3437,N_2788,N_2689);
or U3438 (N_3438,N_2819,N_2677);
or U3439 (N_3439,N_2594,N_2542);
or U3440 (N_3440,N_2817,N_2510);
nand U3441 (N_3441,N_2824,N_2510);
xor U3442 (N_3442,N_2814,N_2805);
nand U3443 (N_3443,N_2885,N_2935);
or U3444 (N_3444,N_2563,N_2514);
nand U3445 (N_3445,N_2685,N_2737);
and U3446 (N_3446,N_2733,N_2697);
xor U3447 (N_3447,N_2643,N_2605);
or U3448 (N_3448,N_2694,N_2574);
nor U3449 (N_3449,N_2638,N_2522);
and U3450 (N_3450,N_2914,N_2987);
xnor U3451 (N_3451,N_2779,N_2892);
xnor U3452 (N_3452,N_2880,N_2662);
or U3453 (N_3453,N_2672,N_2637);
xor U3454 (N_3454,N_2841,N_2800);
nand U3455 (N_3455,N_2515,N_2871);
nor U3456 (N_3456,N_2990,N_2664);
nand U3457 (N_3457,N_2767,N_2622);
or U3458 (N_3458,N_2826,N_2862);
and U3459 (N_3459,N_2938,N_2794);
and U3460 (N_3460,N_2956,N_2883);
nand U3461 (N_3461,N_2866,N_2829);
and U3462 (N_3462,N_2602,N_2677);
and U3463 (N_3463,N_2764,N_2853);
or U3464 (N_3464,N_2733,N_2757);
and U3465 (N_3465,N_2707,N_2927);
and U3466 (N_3466,N_2708,N_2625);
and U3467 (N_3467,N_2604,N_2519);
and U3468 (N_3468,N_2562,N_2585);
nor U3469 (N_3469,N_2930,N_2724);
nand U3470 (N_3470,N_2743,N_2922);
nand U3471 (N_3471,N_2829,N_2998);
nand U3472 (N_3472,N_2682,N_2713);
nor U3473 (N_3473,N_2873,N_2620);
and U3474 (N_3474,N_2772,N_2994);
nand U3475 (N_3475,N_2549,N_2923);
nor U3476 (N_3476,N_2787,N_2848);
nor U3477 (N_3477,N_2864,N_2724);
and U3478 (N_3478,N_2935,N_2668);
xor U3479 (N_3479,N_2680,N_2757);
xnor U3480 (N_3480,N_2550,N_2823);
and U3481 (N_3481,N_2863,N_2558);
and U3482 (N_3482,N_2601,N_2853);
nor U3483 (N_3483,N_2570,N_2555);
nand U3484 (N_3484,N_2726,N_2815);
and U3485 (N_3485,N_2850,N_2709);
nand U3486 (N_3486,N_2990,N_2971);
and U3487 (N_3487,N_2988,N_2907);
xor U3488 (N_3488,N_2980,N_2735);
nor U3489 (N_3489,N_2571,N_2786);
and U3490 (N_3490,N_2645,N_2779);
or U3491 (N_3491,N_2861,N_2902);
nor U3492 (N_3492,N_2513,N_2820);
or U3493 (N_3493,N_2573,N_2574);
nor U3494 (N_3494,N_2832,N_2860);
and U3495 (N_3495,N_2818,N_2692);
nor U3496 (N_3496,N_2970,N_2569);
nor U3497 (N_3497,N_2807,N_2833);
or U3498 (N_3498,N_2521,N_2509);
nor U3499 (N_3499,N_2914,N_2950);
nand U3500 (N_3500,N_3161,N_3407);
nor U3501 (N_3501,N_3458,N_3118);
xnor U3502 (N_3502,N_3169,N_3012);
and U3503 (N_3503,N_3300,N_3324);
nor U3504 (N_3504,N_3189,N_3080);
nor U3505 (N_3505,N_3253,N_3210);
nor U3506 (N_3506,N_3475,N_3236);
xor U3507 (N_3507,N_3063,N_3402);
or U3508 (N_3508,N_3066,N_3067);
and U3509 (N_3509,N_3172,N_3282);
nor U3510 (N_3510,N_3412,N_3431);
or U3511 (N_3511,N_3427,N_3404);
and U3512 (N_3512,N_3486,N_3313);
nor U3513 (N_3513,N_3436,N_3089);
nor U3514 (N_3514,N_3054,N_3468);
xor U3515 (N_3515,N_3115,N_3037);
nand U3516 (N_3516,N_3032,N_3059);
xor U3517 (N_3517,N_3002,N_3369);
and U3518 (N_3518,N_3233,N_3117);
and U3519 (N_3519,N_3192,N_3033);
nor U3520 (N_3520,N_3040,N_3140);
nor U3521 (N_3521,N_3071,N_3353);
xor U3522 (N_3522,N_3060,N_3476);
and U3523 (N_3523,N_3223,N_3384);
xnor U3524 (N_3524,N_3241,N_3430);
xnor U3525 (N_3525,N_3309,N_3100);
and U3526 (N_3526,N_3052,N_3001);
nand U3527 (N_3527,N_3222,N_3039);
xnor U3528 (N_3528,N_3101,N_3143);
and U3529 (N_3529,N_3434,N_3102);
xnor U3530 (N_3530,N_3321,N_3417);
and U3531 (N_3531,N_3483,N_3094);
nor U3532 (N_3532,N_3280,N_3120);
or U3533 (N_3533,N_3494,N_3336);
nor U3534 (N_3534,N_3275,N_3408);
and U3535 (N_3535,N_3316,N_3165);
nor U3536 (N_3536,N_3194,N_3205);
nand U3537 (N_3537,N_3305,N_3358);
nand U3538 (N_3538,N_3278,N_3107);
nand U3539 (N_3539,N_3307,N_3145);
nor U3540 (N_3540,N_3249,N_3057);
and U3541 (N_3541,N_3003,N_3279);
nor U3542 (N_3542,N_3418,N_3461);
xor U3543 (N_3543,N_3367,N_3030);
and U3544 (N_3544,N_3329,N_3053);
and U3545 (N_3545,N_3159,N_3262);
or U3546 (N_3546,N_3320,N_3270);
and U3547 (N_3547,N_3195,N_3055);
nor U3548 (N_3548,N_3331,N_3023);
nand U3549 (N_3549,N_3413,N_3126);
nand U3550 (N_3550,N_3062,N_3184);
and U3551 (N_3551,N_3128,N_3457);
nor U3552 (N_3552,N_3371,N_3056);
and U3553 (N_3553,N_3204,N_3111);
nand U3554 (N_3554,N_3360,N_3416);
nand U3555 (N_3555,N_3050,N_3151);
nand U3556 (N_3556,N_3113,N_3209);
nand U3557 (N_3557,N_3301,N_3451);
or U3558 (N_3558,N_3293,N_3273);
and U3559 (N_3559,N_3449,N_3000);
xnor U3560 (N_3560,N_3394,N_3068);
nand U3561 (N_3561,N_3386,N_3440);
nor U3562 (N_3562,N_3011,N_3297);
or U3563 (N_3563,N_3424,N_3295);
xor U3564 (N_3564,N_3401,N_3227);
nand U3565 (N_3565,N_3382,N_3347);
nand U3566 (N_3566,N_3147,N_3229);
nor U3567 (N_3567,N_3354,N_3093);
nand U3568 (N_3568,N_3356,N_3272);
or U3569 (N_3569,N_3042,N_3377);
nor U3570 (N_3570,N_3362,N_3142);
xnor U3571 (N_3571,N_3216,N_3281);
nand U3572 (N_3572,N_3422,N_3294);
nor U3573 (N_3573,N_3467,N_3173);
or U3574 (N_3574,N_3397,N_3304);
nor U3575 (N_3575,N_3335,N_3446);
and U3576 (N_3576,N_3256,N_3420);
xnor U3577 (N_3577,N_3064,N_3363);
nand U3578 (N_3578,N_3289,N_3078);
xor U3579 (N_3579,N_3419,N_3239);
nand U3580 (N_3580,N_3084,N_3341);
or U3581 (N_3581,N_3387,N_3245);
or U3582 (N_3582,N_3099,N_3288);
and U3583 (N_3583,N_3224,N_3306);
and U3584 (N_3584,N_3477,N_3479);
nand U3585 (N_3585,N_3463,N_3423);
nor U3586 (N_3586,N_3155,N_3242);
nand U3587 (N_3587,N_3452,N_3332);
and U3588 (N_3588,N_3207,N_3315);
or U3589 (N_3589,N_3330,N_3090);
and U3590 (N_3590,N_3473,N_3237);
nand U3591 (N_3591,N_3466,N_3025);
nand U3592 (N_3592,N_3257,N_3274);
and U3593 (N_3593,N_3474,N_3203);
or U3594 (N_3594,N_3043,N_3049);
and U3595 (N_3595,N_3337,N_3160);
nand U3596 (N_3596,N_3010,N_3490);
xnor U3597 (N_3597,N_3087,N_3131);
nand U3598 (N_3598,N_3414,N_3240);
and U3599 (N_3599,N_3266,N_3497);
nor U3600 (N_3600,N_3323,N_3211);
or U3601 (N_3601,N_3103,N_3065);
xnor U3602 (N_3602,N_3044,N_3435);
and U3603 (N_3603,N_3129,N_3198);
nor U3604 (N_3604,N_3465,N_3472);
and U3605 (N_3605,N_3124,N_3439);
and U3606 (N_3606,N_3119,N_3009);
or U3607 (N_3607,N_3469,N_3459);
or U3608 (N_3608,N_3141,N_3166);
and U3609 (N_3609,N_3041,N_3244);
nor U3610 (N_3610,N_3174,N_3214);
nand U3611 (N_3611,N_3433,N_3499);
nand U3612 (N_3612,N_3136,N_3149);
or U3613 (N_3613,N_3235,N_3379);
nor U3614 (N_3614,N_3106,N_3411);
nor U3615 (N_3615,N_3208,N_3183);
and U3616 (N_3616,N_3406,N_3212);
nand U3617 (N_3617,N_3276,N_3287);
nand U3618 (N_3618,N_3082,N_3496);
or U3619 (N_3619,N_3284,N_3482);
nand U3620 (N_3620,N_3088,N_3492);
or U3621 (N_3621,N_3385,N_3154);
and U3622 (N_3622,N_3123,N_3374);
or U3623 (N_3623,N_3221,N_3074);
nand U3624 (N_3624,N_3197,N_3260);
xor U3625 (N_3625,N_3453,N_3139);
and U3626 (N_3626,N_3283,N_3188);
and U3627 (N_3627,N_3134,N_3455);
nand U3628 (N_3628,N_3248,N_3447);
or U3629 (N_3629,N_3213,N_3083);
and U3630 (N_3630,N_3020,N_3426);
or U3631 (N_3631,N_3488,N_3368);
or U3632 (N_3632,N_3398,N_3031);
or U3633 (N_3633,N_3438,N_3029);
and U3634 (N_3634,N_3125,N_3375);
nand U3635 (N_3635,N_3478,N_3327);
xnor U3636 (N_3636,N_3403,N_3421);
and U3637 (N_3637,N_3046,N_3308);
xnor U3638 (N_3638,N_3372,N_3344);
and U3639 (N_3639,N_3196,N_3092);
xor U3640 (N_3640,N_3073,N_3311);
nor U3641 (N_3641,N_3365,N_3180);
or U3642 (N_3642,N_3491,N_3013);
or U3643 (N_3643,N_3035,N_3005);
xor U3644 (N_3644,N_3376,N_3391);
nor U3645 (N_3645,N_3428,N_3069);
nor U3646 (N_3646,N_3217,N_3022);
xor U3647 (N_3647,N_3399,N_3097);
and U3648 (N_3648,N_3110,N_3314);
xor U3649 (N_3649,N_3325,N_3348);
nor U3650 (N_3650,N_3392,N_3104);
xnor U3651 (N_3651,N_3206,N_3393);
or U3652 (N_3652,N_3460,N_3004);
xor U3653 (N_3653,N_3326,N_3132);
nand U3654 (N_3654,N_3081,N_3243);
nor U3655 (N_3655,N_3410,N_3373);
xor U3656 (N_3656,N_3095,N_3077);
and U3657 (N_3657,N_3346,N_3319);
nor U3658 (N_3658,N_3310,N_3383);
or U3659 (N_3659,N_3445,N_3036);
nor U3660 (N_3660,N_3462,N_3238);
xor U3661 (N_3661,N_3230,N_3339);
and U3662 (N_3662,N_3024,N_3345);
or U3663 (N_3663,N_3163,N_3096);
nand U3664 (N_3664,N_3026,N_3286);
or U3665 (N_3665,N_3091,N_3493);
nand U3666 (N_3666,N_3109,N_3370);
or U3667 (N_3667,N_3259,N_3144);
or U3668 (N_3668,N_3138,N_3255);
and U3669 (N_3669,N_3116,N_3296);
or U3670 (N_3670,N_3034,N_3016);
and U3671 (N_3671,N_3454,N_3178);
xnor U3672 (N_3672,N_3167,N_3086);
or U3673 (N_3673,N_3015,N_3038);
nor U3674 (N_3674,N_3317,N_3157);
nand U3675 (N_3675,N_3168,N_3006);
nand U3676 (N_3676,N_3108,N_3388);
or U3677 (N_3677,N_3429,N_3498);
nand U3678 (N_3678,N_3127,N_3290);
xor U3679 (N_3679,N_3334,N_3021);
and U3680 (N_3680,N_3098,N_3400);
nand U3681 (N_3681,N_3355,N_3225);
xor U3682 (N_3682,N_3380,N_3271);
and U3683 (N_3683,N_3199,N_3340);
nand U3684 (N_3684,N_3122,N_3264);
xnor U3685 (N_3685,N_3359,N_3228);
nand U3686 (N_3686,N_3105,N_3409);
nand U3687 (N_3687,N_3170,N_3220);
nor U3688 (N_3688,N_3338,N_3051);
xor U3689 (N_3689,N_3378,N_3135);
or U3690 (N_3690,N_3470,N_3258);
or U3691 (N_3691,N_3442,N_3008);
nand U3692 (N_3692,N_3302,N_3201);
nor U3693 (N_3693,N_3246,N_3352);
or U3694 (N_3694,N_3312,N_3481);
xnor U3695 (N_3695,N_3487,N_3441);
and U3696 (N_3696,N_3017,N_3045);
xor U3697 (N_3697,N_3112,N_3121);
nand U3698 (N_3698,N_3061,N_3322);
nor U3699 (N_3699,N_3186,N_3285);
and U3700 (N_3700,N_3179,N_3269);
or U3701 (N_3701,N_3007,N_3219);
nand U3702 (N_3702,N_3218,N_3175);
nor U3703 (N_3703,N_3185,N_3234);
nand U3704 (N_3704,N_3072,N_3361);
and U3705 (N_3705,N_3158,N_3303);
or U3706 (N_3706,N_3495,N_3299);
nand U3707 (N_3707,N_3226,N_3389);
or U3708 (N_3708,N_3396,N_3190);
nand U3709 (N_3709,N_3432,N_3148);
or U3710 (N_3710,N_3471,N_3164);
and U3711 (N_3711,N_3390,N_3443);
xor U3712 (N_3712,N_3156,N_3448);
nor U3713 (N_3713,N_3079,N_3133);
nor U3714 (N_3714,N_3415,N_3152);
nand U3715 (N_3715,N_3268,N_3176);
and U3716 (N_3716,N_3027,N_3291);
or U3717 (N_3717,N_3150,N_3351);
nand U3718 (N_3718,N_3247,N_3450);
xor U3719 (N_3719,N_3267,N_3425);
nand U3720 (N_3720,N_3366,N_3485);
nor U3721 (N_3721,N_3489,N_3187);
and U3722 (N_3722,N_3328,N_3014);
xnor U3723 (N_3723,N_3200,N_3130);
or U3724 (N_3724,N_3349,N_3333);
or U3725 (N_3725,N_3181,N_3318);
and U3726 (N_3726,N_3137,N_3405);
xor U3727 (N_3727,N_3182,N_3480);
and U3728 (N_3728,N_3250,N_3381);
nand U3729 (N_3729,N_3395,N_3193);
or U3730 (N_3730,N_3456,N_3070);
xnor U3731 (N_3731,N_3177,N_3146);
nand U3732 (N_3732,N_3162,N_3085);
and U3733 (N_3733,N_3202,N_3263);
and U3734 (N_3734,N_3018,N_3254);
or U3735 (N_3735,N_3153,N_3357);
nand U3736 (N_3736,N_3075,N_3191);
or U3737 (N_3737,N_3251,N_3444);
or U3738 (N_3738,N_3484,N_3277);
nor U3739 (N_3739,N_3171,N_3231);
or U3740 (N_3740,N_3019,N_3343);
and U3741 (N_3741,N_3342,N_3350);
xnor U3742 (N_3742,N_3265,N_3261);
xnor U3743 (N_3743,N_3232,N_3114);
and U3744 (N_3744,N_3076,N_3292);
and U3745 (N_3745,N_3058,N_3464);
nor U3746 (N_3746,N_3364,N_3048);
xor U3747 (N_3747,N_3252,N_3437);
nand U3748 (N_3748,N_3298,N_3028);
xor U3749 (N_3749,N_3047,N_3215);
or U3750 (N_3750,N_3375,N_3198);
and U3751 (N_3751,N_3166,N_3022);
or U3752 (N_3752,N_3347,N_3243);
nor U3753 (N_3753,N_3006,N_3359);
or U3754 (N_3754,N_3061,N_3227);
nand U3755 (N_3755,N_3354,N_3008);
xnor U3756 (N_3756,N_3481,N_3400);
and U3757 (N_3757,N_3450,N_3106);
or U3758 (N_3758,N_3140,N_3496);
nor U3759 (N_3759,N_3254,N_3221);
nand U3760 (N_3760,N_3345,N_3007);
and U3761 (N_3761,N_3174,N_3047);
nand U3762 (N_3762,N_3260,N_3191);
or U3763 (N_3763,N_3274,N_3206);
and U3764 (N_3764,N_3124,N_3082);
nand U3765 (N_3765,N_3075,N_3478);
xnor U3766 (N_3766,N_3470,N_3117);
nand U3767 (N_3767,N_3041,N_3198);
or U3768 (N_3768,N_3027,N_3175);
nor U3769 (N_3769,N_3092,N_3498);
and U3770 (N_3770,N_3422,N_3192);
or U3771 (N_3771,N_3232,N_3486);
xnor U3772 (N_3772,N_3156,N_3185);
nand U3773 (N_3773,N_3338,N_3055);
and U3774 (N_3774,N_3343,N_3323);
nand U3775 (N_3775,N_3365,N_3159);
or U3776 (N_3776,N_3284,N_3466);
and U3777 (N_3777,N_3283,N_3038);
and U3778 (N_3778,N_3412,N_3487);
nor U3779 (N_3779,N_3303,N_3230);
or U3780 (N_3780,N_3319,N_3090);
nor U3781 (N_3781,N_3321,N_3258);
or U3782 (N_3782,N_3429,N_3127);
xor U3783 (N_3783,N_3390,N_3455);
or U3784 (N_3784,N_3060,N_3225);
nand U3785 (N_3785,N_3175,N_3239);
nor U3786 (N_3786,N_3147,N_3277);
nor U3787 (N_3787,N_3348,N_3344);
nand U3788 (N_3788,N_3354,N_3372);
xor U3789 (N_3789,N_3037,N_3282);
or U3790 (N_3790,N_3489,N_3217);
or U3791 (N_3791,N_3416,N_3173);
nand U3792 (N_3792,N_3035,N_3123);
or U3793 (N_3793,N_3004,N_3205);
nor U3794 (N_3794,N_3440,N_3109);
nand U3795 (N_3795,N_3493,N_3004);
nand U3796 (N_3796,N_3074,N_3034);
nor U3797 (N_3797,N_3075,N_3411);
nor U3798 (N_3798,N_3051,N_3278);
nand U3799 (N_3799,N_3389,N_3296);
xnor U3800 (N_3800,N_3412,N_3161);
nor U3801 (N_3801,N_3448,N_3046);
or U3802 (N_3802,N_3120,N_3182);
nor U3803 (N_3803,N_3389,N_3264);
xor U3804 (N_3804,N_3497,N_3076);
and U3805 (N_3805,N_3325,N_3385);
nor U3806 (N_3806,N_3394,N_3084);
nand U3807 (N_3807,N_3236,N_3427);
and U3808 (N_3808,N_3202,N_3155);
nor U3809 (N_3809,N_3336,N_3172);
nand U3810 (N_3810,N_3261,N_3045);
nor U3811 (N_3811,N_3424,N_3484);
nor U3812 (N_3812,N_3006,N_3120);
xor U3813 (N_3813,N_3313,N_3113);
xor U3814 (N_3814,N_3491,N_3318);
and U3815 (N_3815,N_3499,N_3495);
nor U3816 (N_3816,N_3226,N_3397);
nor U3817 (N_3817,N_3334,N_3159);
nor U3818 (N_3818,N_3298,N_3153);
or U3819 (N_3819,N_3024,N_3095);
or U3820 (N_3820,N_3025,N_3124);
xor U3821 (N_3821,N_3078,N_3126);
xor U3822 (N_3822,N_3163,N_3498);
nand U3823 (N_3823,N_3225,N_3219);
and U3824 (N_3824,N_3114,N_3024);
or U3825 (N_3825,N_3466,N_3305);
xor U3826 (N_3826,N_3117,N_3419);
nand U3827 (N_3827,N_3081,N_3263);
xnor U3828 (N_3828,N_3160,N_3016);
xor U3829 (N_3829,N_3407,N_3380);
or U3830 (N_3830,N_3473,N_3193);
nor U3831 (N_3831,N_3479,N_3128);
and U3832 (N_3832,N_3285,N_3370);
nand U3833 (N_3833,N_3109,N_3427);
nand U3834 (N_3834,N_3222,N_3317);
or U3835 (N_3835,N_3409,N_3179);
and U3836 (N_3836,N_3305,N_3092);
xor U3837 (N_3837,N_3428,N_3120);
nor U3838 (N_3838,N_3119,N_3155);
and U3839 (N_3839,N_3413,N_3168);
and U3840 (N_3840,N_3412,N_3045);
xor U3841 (N_3841,N_3021,N_3204);
or U3842 (N_3842,N_3167,N_3108);
nor U3843 (N_3843,N_3184,N_3248);
and U3844 (N_3844,N_3053,N_3404);
xnor U3845 (N_3845,N_3486,N_3330);
nand U3846 (N_3846,N_3312,N_3077);
or U3847 (N_3847,N_3096,N_3284);
and U3848 (N_3848,N_3003,N_3213);
nor U3849 (N_3849,N_3385,N_3237);
or U3850 (N_3850,N_3369,N_3340);
or U3851 (N_3851,N_3198,N_3453);
and U3852 (N_3852,N_3081,N_3120);
and U3853 (N_3853,N_3168,N_3352);
nor U3854 (N_3854,N_3336,N_3370);
nor U3855 (N_3855,N_3394,N_3143);
nand U3856 (N_3856,N_3217,N_3191);
or U3857 (N_3857,N_3496,N_3163);
or U3858 (N_3858,N_3323,N_3086);
and U3859 (N_3859,N_3418,N_3493);
xor U3860 (N_3860,N_3471,N_3304);
or U3861 (N_3861,N_3355,N_3445);
nand U3862 (N_3862,N_3084,N_3050);
or U3863 (N_3863,N_3212,N_3414);
xnor U3864 (N_3864,N_3139,N_3415);
nand U3865 (N_3865,N_3009,N_3068);
and U3866 (N_3866,N_3325,N_3193);
nor U3867 (N_3867,N_3043,N_3159);
nand U3868 (N_3868,N_3281,N_3222);
nor U3869 (N_3869,N_3242,N_3319);
nand U3870 (N_3870,N_3429,N_3120);
or U3871 (N_3871,N_3039,N_3071);
nand U3872 (N_3872,N_3032,N_3252);
nor U3873 (N_3873,N_3327,N_3158);
nand U3874 (N_3874,N_3412,N_3283);
nor U3875 (N_3875,N_3346,N_3311);
xor U3876 (N_3876,N_3390,N_3185);
nor U3877 (N_3877,N_3341,N_3220);
xnor U3878 (N_3878,N_3410,N_3339);
and U3879 (N_3879,N_3016,N_3475);
xor U3880 (N_3880,N_3293,N_3427);
nand U3881 (N_3881,N_3258,N_3187);
nor U3882 (N_3882,N_3101,N_3164);
or U3883 (N_3883,N_3222,N_3267);
or U3884 (N_3884,N_3468,N_3265);
or U3885 (N_3885,N_3009,N_3138);
nor U3886 (N_3886,N_3091,N_3419);
nand U3887 (N_3887,N_3459,N_3099);
or U3888 (N_3888,N_3216,N_3208);
nor U3889 (N_3889,N_3006,N_3285);
xor U3890 (N_3890,N_3363,N_3137);
xor U3891 (N_3891,N_3164,N_3354);
or U3892 (N_3892,N_3347,N_3289);
nand U3893 (N_3893,N_3312,N_3045);
xnor U3894 (N_3894,N_3037,N_3278);
xor U3895 (N_3895,N_3463,N_3342);
nor U3896 (N_3896,N_3403,N_3064);
xor U3897 (N_3897,N_3128,N_3148);
or U3898 (N_3898,N_3002,N_3193);
xor U3899 (N_3899,N_3107,N_3158);
xor U3900 (N_3900,N_3148,N_3072);
nand U3901 (N_3901,N_3442,N_3202);
xnor U3902 (N_3902,N_3267,N_3139);
nor U3903 (N_3903,N_3438,N_3115);
nor U3904 (N_3904,N_3256,N_3376);
nor U3905 (N_3905,N_3053,N_3077);
nand U3906 (N_3906,N_3225,N_3054);
nor U3907 (N_3907,N_3442,N_3281);
xnor U3908 (N_3908,N_3196,N_3353);
or U3909 (N_3909,N_3192,N_3497);
nand U3910 (N_3910,N_3473,N_3128);
nand U3911 (N_3911,N_3000,N_3269);
and U3912 (N_3912,N_3193,N_3352);
nand U3913 (N_3913,N_3373,N_3185);
or U3914 (N_3914,N_3215,N_3148);
and U3915 (N_3915,N_3486,N_3307);
nor U3916 (N_3916,N_3070,N_3135);
xnor U3917 (N_3917,N_3112,N_3403);
nor U3918 (N_3918,N_3025,N_3098);
and U3919 (N_3919,N_3497,N_3054);
nand U3920 (N_3920,N_3028,N_3162);
nor U3921 (N_3921,N_3123,N_3340);
xnor U3922 (N_3922,N_3061,N_3414);
and U3923 (N_3923,N_3048,N_3018);
xnor U3924 (N_3924,N_3357,N_3206);
or U3925 (N_3925,N_3034,N_3117);
or U3926 (N_3926,N_3432,N_3397);
nand U3927 (N_3927,N_3016,N_3157);
or U3928 (N_3928,N_3033,N_3267);
nand U3929 (N_3929,N_3041,N_3225);
xnor U3930 (N_3930,N_3207,N_3057);
or U3931 (N_3931,N_3214,N_3058);
nand U3932 (N_3932,N_3251,N_3409);
or U3933 (N_3933,N_3376,N_3258);
nor U3934 (N_3934,N_3148,N_3459);
nand U3935 (N_3935,N_3321,N_3282);
nand U3936 (N_3936,N_3274,N_3002);
or U3937 (N_3937,N_3014,N_3008);
nand U3938 (N_3938,N_3277,N_3016);
xnor U3939 (N_3939,N_3458,N_3256);
xnor U3940 (N_3940,N_3060,N_3152);
and U3941 (N_3941,N_3406,N_3054);
nand U3942 (N_3942,N_3084,N_3288);
or U3943 (N_3943,N_3152,N_3476);
nand U3944 (N_3944,N_3370,N_3301);
nor U3945 (N_3945,N_3022,N_3386);
or U3946 (N_3946,N_3038,N_3241);
or U3947 (N_3947,N_3423,N_3355);
and U3948 (N_3948,N_3322,N_3477);
nor U3949 (N_3949,N_3466,N_3258);
nand U3950 (N_3950,N_3311,N_3446);
nor U3951 (N_3951,N_3401,N_3201);
nor U3952 (N_3952,N_3060,N_3357);
xnor U3953 (N_3953,N_3365,N_3370);
nor U3954 (N_3954,N_3370,N_3259);
or U3955 (N_3955,N_3011,N_3299);
xor U3956 (N_3956,N_3081,N_3392);
nand U3957 (N_3957,N_3082,N_3230);
nor U3958 (N_3958,N_3399,N_3074);
nor U3959 (N_3959,N_3059,N_3403);
xor U3960 (N_3960,N_3366,N_3287);
and U3961 (N_3961,N_3379,N_3129);
or U3962 (N_3962,N_3479,N_3212);
or U3963 (N_3963,N_3183,N_3357);
or U3964 (N_3964,N_3058,N_3373);
or U3965 (N_3965,N_3311,N_3286);
xor U3966 (N_3966,N_3395,N_3062);
xor U3967 (N_3967,N_3321,N_3372);
xnor U3968 (N_3968,N_3458,N_3467);
nor U3969 (N_3969,N_3256,N_3479);
and U3970 (N_3970,N_3012,N_3192);
nor U3971 (N_3971,N_3423,N_3342);
nor U3972 (N_3972,N_3128,N_3118);
and U3973 (N_3973,N_3285,N_3478);
xor U3974 (N_3974,N_3303,N_3474);
nor U3975 (N_3975,N_3133,N_3184);
and U3976 (N_3976,N_3442,N_3457);
or U3977 (N_3977,N_3132,N_3214);
xnor U3978 (N_3978,N_3157,N_3436);
or U3979 (N_3979,N_3147,N_3138);
or U3980 (N_3980,N_3245,N_3179);
nor U3981 (N_3981,N_3428,N_3195);
nand U3982 (N_3982,N_3433,N_3289);
and U3983 (N_3983,N_3247,N_3063);
nor U3984 (N_3984,N_3123,N_3040);
or U3985 (N_3985,N_3029,N_3035);
nand U3986 (N_3986,N_3060,N_3096);
nand U3987 (N_3987,N_3018,N_3498);
nor U3988 (N_3988,N_3401,N_3473);
and U3989 (N_3989,N_3280,N_3332);
xnor U3990 (N_3990,N_3376,N_3467);
nor U3991 (N_3991,N_3114,N_3258);
nor U3992 (N_3992,N_3451,N_3130);
and U3993 (N_3993,N_3467,N_3249);
nor U3994 (N_3994,N_3490,N_3152);
xnor U3995 (N_3995,N_3111,N_3173);
nor U3996 (N_3996,N_3375,N_3474);
nor U3997 (N_3997,N_3152,N_3029);
xnor U3998 (N_3998,N_3433,N_3052);
nor U3999 (N_3999,N_3022,N_3427);
nor U4000 (N_4000,N_3807,N_3976);
nand U4001 (N_4001,N_3663,N_3787);
or U4002 (N_4002,N_3552,N_3996);
xnor U4003 (N_4003,N_3925,N_3828);
nor U4004 (N_4004,N_3887,N_3837);
xnor U4005 (N_4005,N_3739,N_3588);
xor U4006 (N_4006,N_3891,N_3578);
nand U4007 (N_4007,N_3999,N_3892);
nand U4008 (N_4008,N_3883,N_3762);
nor U4009 (N_4009,N_3812,N_3725);
nor U4010 (N_4010,N_3648,N_3558);
xor U4011 (N_4011,N_3681,N_3877);
xor U4012 (N_4012,N_3817,N_3833);
xor U4013 (N_4013,N_3577,N_3746);
nand U4014 (N_4014,N_3857,N_3628);
xnor U4015 (N_4015,N_3984,N_3820);
xor U4016 (N_4016,N_3916,N_3572);
nor U4017 (N_4017,N_3638,N_3629);
nand U4018 (N_4018,N_3599,N_3990);
nor U4019 (N_4019,N_3635,N_3709);
xnor U4020 (N_4020,N_3789,N_3566);
or U4021 (N_4021,N_3710,N_3574);
nand U4022 (N_4022,N_3611,N_3603);
xnor U4023 (N_4023,N_3604,N_3948);
and U4024 (N_4024,N_3782,N_3893);
nor U4025 (N_4025,N_3597,N_3956);
xor U4026 (N_4026,N_3672,N_3803);
and U4027 (N_4027,N_3818,N_3754);
and U4028 (N_4028,N_3840,N_3750);
and U4029 (N_4029,N_3849,N_3794);
nor U4030 (N_4030,N_3941,N_3508);
and U4031 (N_4031,N_3571,N_3796);
or U4032 (N_4032,N_3593,N_3946);
xnor U4033 (N_4033,N_3627,N_3583);
nand U4034 (N_4034,N_3717,N_3686);
or U4035 (N_4035,N_3576,N_3825);
and U4036 (N_4036,N_3591,N_3622);
xnor U4037 (N_4037,N_3748,N_3856);
and U4038 (N_4038,N_3902,N_3507);
nor U4039 (N_4039,N_3886,N_3683);
or U4040 (N_4040,N_3920,N_3871);
nor U4041 (N_4041,N_3601,N_3691);
or U4042 (N_4042,N_3685,N_3829);
xnor U4043 (N_4043,N_3696,N_3805);
xnor U4044 (N_4044,N_3503,N_3866);
nand U4045 (N_4045,N_3526,N_3510);
or U4046 (N_4046,N_3512,N_3816);
nor U4047 (N_4047,N_3934,N_3620);
and U4048 (N_4048,N_3551,N_3736);
or U4049 (N_4049,N_3617,N_3894);
or U4050 (N_4050,N_3589,N_3918);
nor U4051 (N_4051,N_3865,N_3838);
nor U4052 (N_4052,N_3878,N_3904);
or U4053 (N_4053,N_3749,N_3908);
nand U4054 (N_4054,N_3610,N_3623);
nor U4055 (N_4055,N_3722,N_3687);
or U4056 (N_4056,N_3786,N_3734);
nor U4057 (N_4057,N_3703,N_3674);
nor U4058 (N_4058,N_3826,N_3719);
and U4059 (N_4059,N_3937,N_3907);
or U4060 (N_4060,N_3567,N_3753);
xnor U4061 (N_4061,N_3783,N_3953);
nor U4062 (N_4062,N_3797,N_3940);
nor U4063 (N_4063,N_3502,N_3777);
or U4064 (N_4064,N_3835,N_3945);
and U4065 (N_4065,N_3614,N_3602);
or U4066 (N_4066,N_3778,N_3757);
nor U4067 (N_4067,N_3720,N_3671);
nand U4068 (N_4068,N_3923,N_3861);
xor U4069 (N_4069,N_3832,N_3939);
xnor U4070 (N_4070,N_3524,N_3932);
nand U4071 (N_4071,N_3693,N_3959);
nor U4072 (N_4072,N_3582,N_3520);
xor U4073 (N_4073,N_3554,N_3525);
or U4074 (N_4074,N_3884,N_3810);
or U4075 (N_4075,N_3735,N_3543);
and U4076 (N_4076,N_3718,N_3855);
nand U4077 (N_4077,N_3643,N_3901);
or U4078 (N_4078,N_3867,N_3973);
or U4079 (N_4079,N_3821,N_3788);
nor U4080 (N_4080,N_3715,N_3637);
nand U4081 (N_4081,N_3982,N_3698);
nand U4082 (N_4082,N_3542,N_3500);
nor U4083 (N_4083,N_3765,N_3701);
xor U4084 (N_4084,N_3804,N_3669);
and U4085 (N_4085,N_3966,N_3625);
xor U4086 (N_4086,N_3652,N_3596);
or U4087 (N_4087,N_3707,N_3742);
or U4088 (N_4088,N_3540,N_3708);
xor U4089 (N_4089,N_3926,N_3606);
xor U4090 (N_4090,N_3523,N_3852);
or U4091 (N_4091,N_3922,N_3899);
and U4092 (N_4092,N_3732,N_3979);
xnor U4093 (N_4093,N_3967,N_3961);
nand U4094 (N_4094,N_3724,N_3793);
and U4095 (N_4095,N_3668,N_3974);
or U4096 (N_4096,N_3522,N_3986);
or U4097 (N_4097,N_3615,N_3743);
nand U4098 (N_4098,N_3758,N_3565);
xnor U4099 (N_4099,N_3759,N_3642);
xnor U4100 (N_4100,N_3546,N_3851);
or U4101 (N_4101,N_3760,N_3532);
xor U4102 (N_4102,N_3790,N_3957);
xor U4103 (N_4103,N_3699,N_3676);
nor U4104 (N_4104,N_3859,N_3645);
nor U4105 (N_4105,N_3679,N_3933);
and U4106 (N_4106,N_3738,N_3563);
nand U4107 (N_4107,N_3983,N_3624);
nand U4108 (N_4108,N_3890,N_3590);
xnor U4109 (N_4109,N_3792,N_3665);
and U4110 (N_4110,N_3655,N_3773);
and U4111 (N_4111,N_3958,N_3533);
and U4112 (N_4112,N_3905,N_3954);
and U4113 (N_4113,N_3915,N_3801);
nand U4114 (N_4114,N_3795,N_3895);
nor U4115 (N_4115,N_3767,N_3573);
nand U4116 (N_4116,N_3869,N_3534);
or U4117 (N_4117,N_3863,N_3771);
nor U4118 (N_4118,N_3987,N_3616);
or U4119 (N_4119,N_3521,N_3694);
or U4120 (N_4120,N_3870,N_3808);
xnor U4121 (N_4121,N_3677,N_3545);
or U4122 (N_4122,N_3682,N_3666);
and U4123 (N_4123,N_3631,N_3791);
nand U4124 (N_4124,N_3650,N_3921);
xor U4125 (N_4125,N_3850,N_3761);
or U4126 (N_4126,N_3535,N_3653);
nand U4127 (N_4127,N_3721,N_3673);
or U4128 (N_4128,N_3784,N_3882);
or U4129 (N_4129,N_3539,N_3943);
or U4130 (N_4130,N_3897,N_3639);
nand U4131 (N_4131,N_3822,N_3538);
and U4132 (N_4132,N_3785,N_3704);
nand U4133 (N_4133,N_3692,N_3881);
xnor U4134 (N_4134,N_3823,N_3800);
or U4135 (N_4135,N_3579,N_3740);
or U4136 (N_4136,N_3880,N_3811);
or U4137 (N_4137,N_3872,N_3560);
nand U4138 (N_4138,N_3695,N_3705);
or U4139 (N_4139,N_3659,N_3839);
xnor U4140 (N_4140,N_3644,N_3684);
nand U4141 (N_4141,N_3667,N_3561);
or U4142 (N_4142,N_3744,N_3570);
and U4143 (N_4143,N_3930,N_3727);
xnor U4144 (N_4144,N_3978,N_3955);
nand U4145 (N_4145,N_3858,N_3547);
or U4146 (N_4146,N_3585,N_3975);
nand U4147 (N_4147,N_3711,N_3843);
or U4148 (N_4148,N_3714,N_3824);
or U4149 (N_4149,N_3947,N_3656);
xor U4150 (N_4150,N_3658,N_3556);
nand U4151 (N_4151,N_3670,N_3592);
and U4152 (N_4152,N_3609,N_3853);
nor U4153 (N_4153,N_3841,N_3848);
and U4154 (N_4154,N_3660,N_3731);
nand U4155 (N_4155,N_3917,N_3914);
or U4156 (N_4156,N_3518,N_3755);
and U4157 (N_4157,N_3944,N_3516);
and U4158 (N_4158,N_3876,N_3564);
nor U4159 (N_4159,N_3690,N_3657);
and U4160 (N_4160,N_3607,N_3621);
or U4161 (N_4161,N_3991,N_3651);
or U4162 (N_4162,N_3995,N_3557);
and U4163 (N_4163,N_3531,N_3636);
nand U4164 (N_4164,N_3594,N_3798);
nand U4165 (N_4165,N_3776,N_3548);
xor U4166 (N_4166,N_3741,N_3752);
xnor U4167 (N_4167,N_3847,N_3646);
xnor U4168 (N_4168,N_3885,N_3555);
nand U4169 (N_4169,N_3514,N_3927);
and U4170 (N_4170,N_3661,N_3649);
nand U4171 (N_4171,N_3630,N_3831);
nand U4172 (N_4172,N_3575,N_3972);
xor U4173 (N_4173,N_3536,N_3950);
nand U4174 (N_4174,N_3968,N_3780);
or U4175 (N_4175,N_3879,N_3906);
or U4176 (N_4176,N_3842,N_3772);
xnor U4177 (N_4177,N_3529,N_3504);
xor U4178 (N_4178,N_3697,N_3779);
nand U4179 (N_4179,N_3864,N_3559);
nor U4180 (N_4180,N_3900,N_3846);
nor U4181 (N_4181,N_3723,N_3912);
or U4182 (N_4182,N_3549,N_3612);
nor U4183 (N_4183,N_3550,N_3931);
and U4184 (N_4184,N_3706,N_3626);
and U4185 (N_4185,N_3598,N_3647);
nor U4186 (N_4186,N_3586,N_3938);
or U4187 (N_4187,N_3981,N_3632);
or U4188 (N_4188,N_3619,N_3888);
xor U4189 (N_4189,N_3960,N_3506);
and U4190 (N_4190,N_3909,N_3584);
and U4191 (N_4191,N_3633,N_3580);
or U4192 (N_4192,N_3913,N_3756);
or U4193 (N_4193,N_3581,N_3662);
and U4194 (N_4194,N_3595,N_3729);
xnor U4195 (N_4195,N_3997,N_3998);
or U4196 (N_4196,N_3544,N_3562);
or U4197 (N_4197,N_3541,N_3678);
nand U4198 (N_4198,N_3992,N_3827);
and U4199 (N_4199,N_3664,N_3733);
xor U4200 (N_4200,N_3952,N_3970);
nand U4201 (N_4201,N_3568,N_3688);
xor U4202 (N_4202,N_3834,N_3963);
and U4203 (N_4203,N_3889,N_3969);
nand U4204 (N_4204,N_3763,N_3587);
and U4205 (N_4205,N_3728,N_3519);
nand U4206 (N_4206,N_3702,N_3680);
nand U4207 (N_4207,N_3949,N_3769);
and U4208 (N_4208,N_3903,N_3854);
nand U4209 (N_4209,N_3962,N_3730);
xnor U4210 (N_4210,N_3689,N_3608);
nand U4211 (N_4211,N_3618,N_3745);
nand U4212 (N_4212,N_3527,N_3936);
and U4213 (N_4213,N_3814,N_3605);
nand U4214 (N_4214,N_3802,N_3509);
nand U4215 (N_4215,N_3980,N_3768);
xnor U4216 (N_4216,N_3845,N_3716);
nor U4217 (N_4217,N_3806,N_3971);
nor U4218 (N_4218,N_3553,N_3634);
nor U4219 (N_4219,N_3517,N_3712);
nand U4220 (N_4220,N_3964,N_3928);
nand U4221 (N_4221,N_3530,N_3935);
xor U4222 (N_4222,N_3988,N_3898);
nand U4223 (N_4223,N_3911,N_3860);
or U4224 (N_4224,N_3951,N_3836);
nand U4225 (N_4225,N_3813,N_3640);
nand U4226 (N_4226,N_3910,N_3700);
and U4227 (N_4227,N_3942,N_3874);
nor U4228 (N_4228,N_3799,N_3965);
and U4229 (N_4229,N_3994,N_3830);
xor U4230 (N_4230,N_3766,N_3501);
xor U4231 (N_4231,N_3809,N_3774);
and U4232 (N_4232,N_3569,N_3511);
nand U4233 (N_4233,N_3844,N_3781);
nor U4234 (N_4234,N_3815,N_3875);
or U4235 (N_4235,N_3515,N_3862);
and U4236 (N_4236,N_3989,N_3770);
nor U4237 (N_4237,N_3896,N_3924);
xor U4238 (N_4238,N_3713,N_3977);
and U4239 (N_4239,N_3513,N_3775);
nor U4240 (N_4240,N_3764,N_3613);
or U4241 (N_4241,N_3868,N_3528);
and U4242 (N_4242,N_3747,N_3737);
nand U4243 (N_4243,N_3537,N_3505);
and U4244 (N_4244,N_3919,N_3819);
and U4245 (N_4245,N_3726,N_3993);
nor U4246 (N_4246,N_3929,N_3873);
xnor U4247 (N_4247,N_3641,N_3654);
nor U4248 (N_4248,N_3675,N_3985);
nand U4249 (N_4249,N_3600,N_3751);
nand U4250 (N_4250,N_3753,N_3503);
nand U4251 (N_4251,N_3979,N_3719);
xnor U4252 (N_4252,N_3859,N_3709);
nor U4253 (N_4253,N_3584,N_3678);
nor U4254 (N_4254,N_3739,N_3512);
xnor U4255 (N_4255,N_3760,N_3998);
xnor U4256 (N_4256,N_3981,N_3656);
or U4257 (N_4257,N_3881,N_3667);
xor U4258 (N_4258,N_3623,N_3533);
nand U4259 (N_4259,N_3501,N_3739);
and U4260 (N_4260,N_3733,N_3721);
nor U4261 (N_4261,N_3781,N_3536);
nand U4262 (N_4262,N_3597,N_3941);
nor U4263 (N_4263,N_3829,N_3937);
nand U4264 (N_4264,N_3929,N_3535);
nor U4265 (N_4265,N_3790,N_3876);
nand U4266 (N_4266,N_3648,N_3603);
nand U4267 (N_4267,N_3857,N_3976);
and U4268 (N_4268,N_3635,N_3719);
nand U4269 (N_4269,N_3527,N_3686);
nor U4270 (N_4270,N_3525,N_3730);
or U4271 (N_4271,N_3629,N_3927);
xor U4272 (N_4272,N_3616,N_3998);
nor U4273 (N_4273,N_3521,N_3515);
nor U4274 (N_4274,N_3582,N_3854);
and U4275 (N_4275,N_3536,N_3517);
xor U4276 (N_4276,N_3913,N_3601);
xor U4277 (N_4277,N_3675,N_3642);
nand U4278 (N_4278,N_3951,N_3535);
nor U4279 (N_4279,N_3633,N_3689);
nor U4280 (N_4280,N_3591,N_3785);
nand U4281 (N_4281,N_3992,N_3767);
or U4282 (N_4282,N_3831,N_3922);
nor U4283 (N_4283,N_3512,N_3691);
and U4284 (N_4284,N_3950,N_3773);
and U4285 (N_4285,N_3551,N_3920);
or U4286 (N_4286,N_3653,N_3996);
or U4287 (N_4287,N_3764,N_3569);
and U4288 (N_4288,N_3614,N_3843);
or U4289 (N_4289,N_3803,N_3665);
nand U4290 (N_4290,N_3836,N_3878);
or U4291 (N_4291,N_3695,N_3657);
nor U4292 (N_4292,N_3871,N_3747);
nand U4293 (N_4293,N_3736,N_3639);
nor U4294 (N_4294,N_3601,N_3989);
xor U4295 (N_4295,N_3508,N_3518);
nand U4296 (N_4296,N_3552,N_3661);
xnor U4297 (N_4297,N_3896,N_3574);
xor U4298 (N_4298,N_3653,N_3981);
or U4299 (N_4299,N_3538,N_3834);
nor U4300 (N_4300,N_3693,N_3627);
nand U4301 (N_4301,N_3886,N_3523);
nand U4302 (N_4302,N_3752,N_3901);
xor U4303 (N_4303,N_3884,N_3962);
or U4304 (N_4304,N_3811,N_3898);
or U4305 (N_4305,N_3766,N_3511);
nor U4306 (N_4306,N_3641,N_3569);
and U4307 (N_4307,N_3821,N_3872);
nand U4308 (N_4308,N_3865,N_3642);
xnor U4309 (N_4309,N_3722,N_3716);
or U4310 (N_4310,N_3667,N_3548);
or U4311 (N_4311,N_3721,N_3624);
nor U4312 (N_4312,N_3983,N_3749);
or U4313 (N_4313,N_3806,N_3976);
and U4314 (N_4314,N_3500,N_3782);
nor U4315 (N_4315,N_3507,N_3594);
nor U4316 (N_4316,N_3806,N_3749);
nand U4317 (N_4317,N_3588,N_3676);
nand U4318 (N_4318,N_3937,N_3832);
xnor U4319 (N_4319,N_3852,N_3515);
xor U4320 (N_4320,N_3770,N_3824);
or U4321 (N_4321,N_3501,N_3540);
or U4322 (N_4322,N_3813,N_3572);
and U4323 (N_4323,N_3524,N_3713);
nor U4324 (N_4324,N_3671,N_3746);
and U4325 (N_4325,N_3782,N_3944);
or U4326 (N_4326,N_3955,N_3523);
xor U4327 (N_4327,N_3518,N_3847);
nor U4328 (N_4328,N_3559,N_3808);
nand U4329 (N_4329,N_3584,N_3906);
xnor U4330 (N_4330,N_3871,N_3973);
xor U4331 (N_4331,N_3635,N_3733);
nand U4332 (N_4332,N_3711,N_3958);
or U4333 (N_4333,N_3804,N_3848);
and U4334 (N_4334,N_3650,N_3676);
xnor U4335 (N_4335,N_3793,N_3699);
xor U4336 (N_4336,N_3744,N_3621);
xnor U4337 (N_4337,N_3774,N_3829);
and U4338 (N_4338,N_3841,N_3593);
and U4339 (N_4339,N_3960,N_3534);
nor U4340 (N_4340,N_3907,N_3881);
xor U4341 (N_4341,N_3771,N_3823);
nor U4342 (N_4342,N_3502,N_3858);
and U4343 (N_4343,N_3742,N_3538);
and U4344 (N_4344,N_3920,N_3732);
and U4345 (N_4345,N_3803,N_3849);
and U4346 (N_4346,N_3721,N_3548);
nor U4347 (N_4347,N_3662,N_3640);
xor U4348 (N_4348,N_3793,N_3727);
nand U4349 (N_4349,N_3599,N_3750);
nand U4350 (N_4350,N_3541,N_3531);
nor U4351 (N_4351,N_3928,N_3659);
and U4352 (N_4352,N_3737,N_3707);
nor U4353 (N_4353,N_3874,N_3539);
or U4354 (N_4354,N_3540,N_3926);
and U4355 (N_4355,N_3856,N_3697);
nor U4356 (N_4356,N_3727,N_3702);
and U4357 (N_4357,N_3770,N_3574);
and U4358 (N_4358,N_3673,N_3657);
nand U4359 (N_4359,N_3658,N_3996);
or U4360 (N_4360,N_3675,N_3767);
nor U4361 (N_4361,N_3935,N_3961);
xor U4362 (N_4362,N_3919,N_3623);
or U4363 (N_4363,N_3846,N_3523);
nor U4364 (N_4364,N_3899,N_3823);
or U4365 (N_4365,N_3896,N_3886);
or U4366 (N_4366,N_3741,N_3564);
and U4367 (N_4367,N_3926,N_3609);
or U4368 (N_4368,N_3966,N_3793);
xnor U4369 (N_4369,N_3859,N_3540);
nor U4370 (N_4370,N_3540,N_3751);
nand U4371 (N_4371,N_3719,N_3739);
and U4372 (N_4372,N_3529,N_3985);
and U4373 (N_4373,N_3971,N_3798);
nand U4374 (N_4374,N_3722,N_3666);
xnor U4375 (N_4375,N_3941,N_3530);
nand U4376 (N_4376,N_3532,N_3751);
or U4377 (N_4377,N_3786,N_3871);
or U4378 (N_4378,N_3890,N_3557);
and U4379 (N_4379,N_3745,N_3789);
or U4380 (N_4380,N_3573,N_3980);
xor U4381 (N_4381,N_3851,N_3612);
nor U4382 (N_4382,N_3695,N_3564);
nand U4383 (N_4383,N_3696,N_3720);
or U4384 (N_4384,N_3899,N_3526);
xnor U4385 (N_4385,N_3763,N_3955);
or U4386 (N_4386,N_3731,N_3987);
xnor U4387 (N_4387,N_3622,N_3552);
nor U4388 (N_4388,N_3646,N_3988);
and U4389 (N_4389,N_3515,N_3550);
and U4390 (N_4390,N_3547,N_3550);
nor U4391 (N_4391,N_3516,N_3725);
nand U4392 (N_4392,N_3833,N_3843);
xor U4393 (N_4393,N_3658,N_3597);
nor U4394 (N_4394,N_3779,N_3981);
and U4395 (N_4395,N_3667,N_3892);
nor U4396 (N_4396,N_3765,N_3729);
and U4397 (N_4397,N_3526,N_3512);
nand U4398 (N_4398,N_3798,N_3846);
xnor U4399 (N_4399,N_3680,N_3534);
nand U4400 (N_4400,N_3511,N_3926);
nand U4401 (N_4401,N_3615,N_3641);
nor U4402 (N_4402,N_3609,N_3604);
or U4403 (N_4403,N_3893,N_3921);
xor U4404 (N_4404,N_3518,N_3801);
nor U4405 (N_4405,N_3510,N_3720);
and U4406 (N_4406,N_3753,N_3549);
nor U4407 (N_4407,N_3679,N_3577);
xnor U4408 (N_4408,N_3970,N_3605);
or U4409 (N_4409,N_3714,N_3909);
or U4410 (N_4410,N_3732,N_3619);
or U4411 (N_4411,N_3668,N_3828);
nor U4412 (N_4412,N_3898,N_3794);
or U4413 (N_4413,N_3945,N_3809);
or U4414 (N_4414,N_3953,N_3626);
xnor U4415 (N_4415,N_3805,N_3830);
nor U4416 (N_4416,N_3507,N_3581);
and U4417 (N_4417,N_3986,N_3581);
xor U4418 (N_4418,N_3980,N_3518);
and U4419 (N_4419,N_3904,N_3744);
nand U4420 (N_4420,N_3907,N_3565);
nand U4421 (N_4421,N_3595,N_3575);
or U4422 (N_4422,N_3911,N_3849);
nand U4423 (N_4423,N_3654,N_3894);
or U4424 (N_4424,N_3827,N_3562);
xor U4425 (N_4425,N_3609,N_3747);
xor U4426 (N_4426,N_3650,N_3516);
xor U4427 (N_4427,N_3893,N_3534);
or U4428 (N_4428,N_3591,N_3786);
or U4429 (N_4429,N_3914,N_3930);
and U4430 (N_4430,N_3885,N_3646);
and U4431 (N_4431,N_3982,N_3677);
xor U4432 (N_4432,N_3962,N_3684);
or U4433 (N_4433,N_3949,N_3707);
and U4434 (N_4434,N_3783,N_3935);
xor U4435 (N_4435,N_3931,N_3529);
nand U4436 (N_4436,N_3548,N_3763);
or U4437 (N_4437,N_3578,N_3504);
xor U4438 (N_4438,N_3740,N_3591);
nor U4439 (N_4439,N_3966,N_3978);
nor U4440 (N_4440,N_3953,N_3658);
nor U4441 (N_4441,N_3537,N_3645);
and U4442 (N_4442,N_3833,N_3648);
nor U4443 (N_4443,N_3624,N_3682);
or U4444 (N_4444,N_3933,N_3650);
nand U4445 (N_4445,N_3869,N_3833);
or U4446 (N_4446,N_3839,N_3869);
xor U4447 (N_4447,N_3720,N_3952);
xor U4448 (N_4448,N_3542,N_3764);
and U4449 (N_4449,N_3900,N_3782);
and U4450 (N_4450,N_3641,N_3971);
nor U4451 (N_4451,N_3625,N_3693);
or U4452 (N_4452,N_3668,N_3774);
nand U4453 (N_4453,N_3653,N_3589);
nand U4454 (N_4454,N_3971,N_3842);
xor U4455 (N_4455,N_3878,N_3526);
nand U4456 (N_4456,N_3699,N_3701);
nor U4457 (N_4457,N_3850,N_3506);
and U4458 (N_4458,N_3830,N_3727);
nand U4459 (N_4459,N_3704,N_3510);
nor U4460 (N_4460,N_3968,N_3555);
nor U4461 (N_4461,N_3717,N_3660);
nand U4462 (N_4462,N_3679,N_3561);
and U4463 (N_4463,N_3619,N_3930);
or U4464 (N_4464,N_3921,N_3719);
xnor U4465 (N_4465,N_3904,N_3565);
or U4466 (N_4466,N_3691,N_3901);
and U4467 (N_4467,N_3866,N_3651);
nor U4468 (N_4468,N_3802,N_3929);
and U4469 (N_4469,N_3695,N_3516);
xnor U4470 (N_4470,N_3779,N_3598);
nand U4471 (N_4471,N_3667,N_3830);
nor U4472 (N_4472,N_3615,N_3856);
or U4473 (N_4473,N_3924,N_3949);
nor U4474 (N_4474,N_3802,N_3847);
nand U4475 (N_4475,N_3880,N_3691);
nand U4476 (N_4476,N_3656,N_3969);
nor U4477 (N_4477,N_3848,N_3656);
and U4478 (N_4478,N_3780,N_3779);
and U4479 (N_4479,N_3568,N_3983);
xor U4480 (N_4480,N_3971,N_3649);
nor U4481 (N_4481,N_3810,N_3863);
nor U4482 (N_4482,N_3507,N_3621);
nor U4483 (N_4483,N_3819,N_3572);
or U4484 (N_4484,N_3726,N_3870);
nand U4485 (N_4485,N_3953,N_3668);
xor U4486 (N_4486,N_3864,N_3697);
xor U4487 (N_4487,N_3547,N_3922);
or U4488 (N_4488,N_3781,N_3818);
xnor U4489 (N_4489,N_3548,N_3813);
nand U4490 (N_4490,N_3546,N_3634);
or U4491 (N_4491,N_3954,N_3741);
or U4492 (N_4492,N_3574,N_3807);
nand U4493 (N_4493,N_3599,N_3508);
and U4494 (N_4494,N_3543,N_3711);
or U4495 (N_4495,N_3527,N_3650);
nand U4496 (N_4496,N_3848,N_3789);
xnor U4497 (N_4497,N_3855,N_3733);
nand U4498 (N_4498,N_3504,N_3971);
or U4499 (N_4499,N_3937,N_3861);
nor U4500 (N_4500,N_4256,N_4214);
nand U4501 (N_4501,N_4082,N_4466);
or U4502 (N_4502,N_4370,N_4169);
or U4503 (N_4503,N_4196,N_4431);
or U4504 (N_4504,N_4405,N_4389);
or U4505 (N_4505,N_4114,N_4319);
and U4506 (N_4506,N_4206,N_4390);
and U4507 (N_4507,N_4134,N_4302);
xor U4508 (N_4508,N_4093,N_4367);
or U4509 (N_4509,N_4008,N_4351);
or U4510 (N_4510,N_4213,N_4393);
xnor U4511 (N_4511,N_4136,N_4373);
or U4512 (N_4512,N_4081,N_4440);
and U4513 (N_4513,N_4018,N_4332);
xnor U4514 (N_4514,N_4043,N_4113);
nor U4515 (N_4515,N_4178,N_4496);
xor U4516 (N_4516,N_4293,N_4062);
nand U4517 (N_4517,N_4184,N_4096);
or U4518 (N_4518,N_4479,N_4363);
and U4519 (N_4519,N_4427,N_4376);
or U4520 (N_4520,N_4139,N_4112);
xor U4521 (N_4521,N_4212,N_4333);
nor U4522 (N_4522,N_4308,N_4147);
nor U4523 (N_4523,N_4138,N_4494);
xnor U4524 (N_4524,N_4239,N_4472);
xnor U4525 (N_4525,N_4310,N_4300);
and U4526 (N_4526,N_4187,N_4452);
nor U4527 (N_4527,N_4065,N_4489);
nor U4528 (N_4528,N_4135,N_4348);
nand U4529 (N_4529,N_4451,N_4387);
nand U4530 (N_4530,N_4232,N_4357);
xnor U4531 (N_4531,N_4436,N_4072);
xor U4532 (N_4532,N_4444,N_4111);
xor U4533 (N_4533,N_4074,N_4460);
or U4534 (N_4534,N_4498,N_4437);
nor U4535 (N_4535,N_4417,N_4264);
nand U4536 (N_4536,N_4346,N_4411);
nand U4537 (N_4537,N_4281,N_4407);
nand U4538 (N_4538,N_4156,N_4443);
nor U4539 (N_4539,N_4288,N_4034);
or U4540 (N_4540,N_4092,N_4318);
and U4541 (N_4541,N_4204,N_4153);
and U4542 (N_4542,N_4192,N_4480);
nor U4543 (N_4543,N_4273,N_4224);
nor U4544 (N_4544,N_4258,N_4289);
and U4545 (N_4545,N_4492,N_4227);
xnor U4546 (N_4546,N_4179,N_4241);
or U4547 (N_4547,N_4118,N_4410);
or U4548 (N_4548,N_4108,N_4441);
nor U4549 (N_4549,N_4416,N_4091);
or U4550 (N_4550,N_4027,N_4053);
or U4551 (N_4551,N_4029,N_4025);
or U4552 (N_4552,N_4183,N_4173);
xnor U4553 (N_4553,N_4455,N_4471);
or U4554 (N_4554,N_4143,N_4328);
or U4555 (N_4555,N_4068,N_4244);
xor U4556 (N_4556,N_4197,N_4090);
nand U4557 (N_4557,N_4133,N_4282);
or U4558 (N_4558,N_4424,N_4356);
xnor U4559 (N_4559,N_4414,N_4116);
nor U4560 (N_4560,N_4304,N_4033);
and U4561 (N_4561,N_4159,N_4057);
nor U4562 (N_4562,N_4408,N_4174);
nand U4563 (N_4563,N_4209,N_4454);
and U4564 (N_4564,N_4297,N_4433);
nor U4565 (N_4565,N_4465,N_4222);
xor U4566 (N_4566,N_4352,N_4216);
xor U4567 (N_4567,N_4306,N_4166);
nor U4568 (N_4568,N_4329,N_4011);
xnor U4569 (N_4569,N_4246,N_4384);
nor U4570 (N_4570,N_4218,N_4076);
and U4571 (N_4571,N_4382,N_4228);
or U4572 (N_4572,N_4426,N_4186);
nand U4573 (N_4573,N_4117,N_4230);
or U4574 (N_4574,N_4439,N_4482);
nand U4575 (N_4575,N_4265,N_4051);
or U4576 (N_4576,N_4225,N_4128);
or U4577 (N_4577,N_4040,N_4315);
nand U4578 (N_4578,N_4045,N_4019);
xor U4579 (N_4579,N_4038,N_4481);
nor U4580 (N_4580,N_4353,N_4418);
or U4581 (N_4581,N_4080,N_4495);
nor U4582 (N_4582,N_4148,N_4267);
nor U4583 (N_4583,N_4361,N_4007);
or U4584 (N_4584,N_4342,N_4331);
or U4585 (N_4585,N_4330,N_4069);
or U4586 (N_4586,N_4110,N_4320);
or U4587 (N_4587,N_4022,N_4369);
nand U4588 (N_4588,N_4420,N_4084);
or U4589 (N_4589,N_4485,N_4185);
and U4590 (N_4590,N_4262,N_4486);
or U4591 (N_4591,N_4161,N_4151);
or U4592 (N_4592,N_4350,N_4383);
nand U4593 (N_4593,N_4359,N_4312);
nand U4594 (N_4594,N_4474,N_4176);
nor U4595 (N_4595,N_4165,N_4155);
or U4596 (N_4596,N_4044,N_4021);
and U4597 (N_4597,N_4257,N_4487);
and U4598 (N_4598,N_4002,N_4399);
and U4599 (N_4599,N_4075,N_4012);
nor U4600 (N_4600,N_4146,N_4275);
and U4601 (N_4601,N_4120,N_4326);
xnor U4602 (N_4602,N_4442,N_4321);
xnor U4603 (N_4603,N_4126,N_4154);
and U4604 (N_4604,N_4119,N_4031);
and U4605 (N_4605,N_4391,N_4396);
xor U4606 (N_4606,N_4221,N_4423);
or U4607 (N_4607,N_4255,N_4470);
nor U4608 (N_4608,N_4132,N_4272);
nand U4609 (N_4609,N_4458,N_4432);
or U4610 (N_4610,N_4398,N_4061);
and U4611 (N_4611,N_4263,N_4125);
nor U4612 (N_4612,N_4254,N_4298);
nor U4613 (N_4613,N_4368,N_4338);
nor U4614 (N_4614,N_4249,N_4371);
and U4615 (N_4615,N_4109,N_4217);
or U4616 (N_4616,N_4087,N_4234);
nor U4617 (N_4617,N_4088,N_4127);
or U4618 (N_4618,N_4296,N_4137);
xnor U4619 (N_4619,N_4462,N_4415);
xor U4620 (N_4620,N_4307,N_4064);
or U4621 (N_4621,N_4168,N_4177);
nor U4622 (N_4622,N_4236,N_4059);
xor U4623 (N_4623,N_4476,N_4469);
nand U4624 (N_4624,N_4006,N_4499);
nand U4625 (N_4625,N_4140,N_4245);
nand U4626 (N_4626,N_4419,N_4199);
nor U4627 (N_4627,N_4409,N_4028);
xor U4628 (N_4628,N_4171,N_4286);
and U4629 (N_4629,N_4467,N_4438);
nor U4630 (N_4630,N_4392,N_4477);
nand U4631 (N_4631,N_4071,N_4464);
and U4632 (N_4632,N_4106,N_4219);
nand U4633 (N_4633,N_4295,N_4400);
nand U4634 (N_4634,N_4395,N_4343);
xnor U4635 (N_4635,N_4484,N_4233);
nand U4636 (N_4636,N_4003,N_4063);
xor U4637 (N_4637,N_4172,N_4035);
nand U4638 (N_4638,N_4314,N_4129);
nand U4639 (N_4639,N_4413,N_4004);
xnor U4640 (N_4640,N_4344,N_4097);
nor U4641 (N_4641,N_4380,N_4374);
nor U4642 (N_4642,N_4149,N_4152);
or U4643 (N_4643,N_4226,N_4016);
and U4644 (N_4644,N_4340,N_4089);
and U4645 (N_4645,N_4362,N_4229);
or U4646 (N_4646,N_4290,N_4394);
or U4647 (N_4647,N_4195,N_4164);
and U4648 (N_4648,N_4381,N_4009);
nand U4649 (N_4649,N_4131,N_4180);
and U4650 (N_4650,N_4020,N_4015);
nand U4651 (N_4651,N_4223,N_4242);
or U4652 (N_4652,N_4042,N_4478);
nand U4653 (N_4653,N_4337,N_4163);
and U4654 (N_4654,N_4013,N_4378);
nand U4655 (N_4655,N_4251,N_4336);
nand U4656 (N_4656,N_4100,N_4421);
nor U4657 (N_4657,N_4294,N_4445);
nand U4658 (N_4658,N_4189,N_4317);
and U4659 (N_4659,N_4215,N_4327);
and U4660 (N_4660,N_4341,N_4130);
or U4661 (N_4661,N_4287,N_4299);
nand U4662 (N_4662,N_4123,N_4121);
nor U4663 (N_4663,N_4435,N_4162);
or U4664 (N_4664,N_4010,N_4276);
or U4665 (N_4665,N_4285,N_4124);
xor U4666 (N_4666,N_4447,N_4237);
and U4667 (N_4667,N_4201,N_4453);
nand U4668 (N_4668,N_4268,N_4490);
nor U4669 (N_4669,N_4334,N_4316);
nand U4670 (N_4670,N_4313,N_4354);
nor U4671 (N_4671,N_4190,N_4406);
or U4672 (N_4672,N_4412,N_4032);
nor U4673 (N_4673,N_4017,N_4325);
or U4674 (N_4674,N_4142,N_4349);
nand U4675 (N_4675,N_4050,N_4388);
xor U4676 (N_4676,N_4434,N_4386);
nor U4677 (N_4677,N_4150,N_4048);
or U4678 (N_4678,N_4085,N_4261);
or U4679 (N_4679,N_4014,N_4145);
xnor U4680 (N_4680,N_4203,N_4271);
nand U4681 (N_4681,N_4098,N_4055);
xor U4682 (N_4682,N_4404,N_4270);
xnor U4683 (N_4683,N_4345,N_4060);
and U4684 (N_4684,N_4083,N_4430);
xnor U4685 (N_4685,N_4323,N_4103);
xor U4686 (N_4686,N_4181,N_4364);
or U4687 (N_4687,N_4456,N_4303);
and U4688 (N_4688,N_4182,N_4001);
and U4689 (N_4689,N_4450,N_4073);
xor U4690 (N_4690,N_4122,N_4141);
nand U4691 (N_4691,N_4403,N_4066);
and U4692 (N_4692,N_4105,N_4000);
or U4693 (N_4693,N_4253,N_4079);
and U4694 (N_4694,N_4375,N_4167);
and U4695 (N_4695,N_4429,N_4335);
xor U4696 (N_4696,N_4056,N_4220);
xor U4697 (N_4697,N_4202,N_4036);
nand U4698 (N_4698,N_4301,N_4144);
or U4699 (N_4699,N_4046,N_4305);
xnor U4700 (N_4700,N_4347,N_4269);
nand U4701 (N_4701,N_4459,N_4377);
nand U4702 (N_4702,N_4366,N_4266);
or U4703 (N_4703,N_4365,N_4101);
xor U4704 (N_4704,N_4250,N_4200);
nor U4705 (N_4705,N_4231,N_4158);
xor U4706 (N_4706,N_4358,N_4026);
or U4707 (N_4707,N_4078,N_4243);
or U4708 (N_4708,N_4115,N_4292);
or U4709 (N_4709,N_4402,N_4160);
nand U4710 (N_4710,N_4457,N_4191);
xnor U4711 (N_4711,N_4274,N_4039);
xor U4712 (N_4712,N_4094,N_4425);
xor U4713 (N_4713,N_4397,N_4493);
xor U4714 (N_4714,N_4194,N_4023);
and U4715 (N_4715,N_4291,N_4461);
nor U4716 (N_4716,N_4279,N_4283);
xnor U4717 (N_4717,N_4067,N_4175);
or U4718 (N_4718,N_4193,N_4247);
nand U4719 (N_4719,N_4052,N_4448);
nand U4720 (N_4720,N_4235,N_4483);
nand U4721 (N_4721,N_4210,N_4497);
and U4722 (N_4722,N_4324,N_4449);
and U4723 (N_4723,N_4322,N_4205);
nor U4724 (N_4724,N_4104,N_4475);
xnor U4725 (N_4725,N_4339,N_4259);
xor U4726 (N_4726,N_4107,N_4280);
nor U4727 (N_4727,N_4037,N_4385);
nor U4728 (N_4728,N_4252,N_4030);
nor U4729 (N_4729,N_4372,N_4005);
nand U4730 (N_4730,N_4099,N_4355);
or U4731 (N_4731,N_4491,N_4047);
nand U4732 (N_4732,N_4207,N_4024);
nor U4733 (N_4733,N_4208,N_4054);
and U4734 (N_4734,N_4284,N_4211);
and U4735 (N_4735,N_4468,N_4238);
xor U4736 (N_4736,N_4379,N_4260);
nor U4737 (N_4737,N_4277,N_4401);
or U4738 (N_4738,N_4428,N_4041);
xor U4739 (N_4739,N_4240,N_4058);
nor U4740 (N_4740,N_4095,N_4463);
nor U4741 (N_4741,N_4248,N_4278);
xor U4742 (N_4742,N_4446,N_4473);
xor U4743 (N_4743,N_4157,N_4077);
or U4744 (N_4744,N_4311,N_4070);
and U4745 (N_4745,N_4309,N_4488);
or U4746 (N_4746,N_4198,N_4049);
xnor U4747 (N_4747,N_4188,N_4360);
xor U4748 (N_4748,N_4422,N_4086);
xor U4749 (N_4749,N_4170,N_4102);
or U4750 (N_4750,N_4156,N_4157);
and U4751 (N_4751,N_4415,N_4338);
or U4752 (N_4752,N_4040,N_4181);
nand U4753 (N_4753,N_4287,N_4290);
and U4754 (N_4754,N_4478,N_4230);
and U4755 (N_4755,N_4234,N_4217);
nor U4756 (N_4756,N_4363,N_4108);
or U4757 (N_4757,N_4499,N_4275);
or U4758 (N_4758,N_4295,N_4043);
nor U4759 (N_4759,N_4329,N_4307);
nand U4760 (N_4760,N_4428,N_4215);
and U4761 (N_4761,N_4290,N_4049);
nand U4762 (N_4762,N_4456,N_4157);
or U4763 (N_4763,N_4372,N_4270);
nand U4764 (N_4764,N_4075,N_4193);
xnor U4765 (N_4765,N_4407,N_4110);
nor U4766 (N_4766,N_4161,N_4114);
nand U4767 (N_4767,N_4397,N_4224);
or U4768 (N_4768,N_4427,N_4345);
nand U4769 (N_4769,N_4415,N_4356);
xor U4770 (N_4770,N_4478,N_4458);
and U4771 (N_4771,N_4320,N_4398);
or U4772 (N_4772,N_4192,N_4163);
nor U4773 (N_4773,N_4147,N_4199);
nand U4774 (N_4774,N_4143,N_4146);
nor U4775 (N_4775,N_4371,N_4094);
xor U4776 (N_4776,N_4018,N_4200);
or U4777 (N_4777,N_4159,N_4383);
nand U4778 (N_4778,N_4201,N_4367);
or U4779 (N_4779,N_4394,N_4383);
xor U4780 (N_4780,N_4214,N_4217);
or U4781 (N_4781,N_4318,N_4208);
or U4782 (N_4782,N_4385,N_4476);
xnor U4783 (N_4783,N_4094,N_4048);
or U4784 (N_4784,N_4429,N_4204);
and U4785 (N_4785,N_4192,N_4404);
and U4786 (N_4786,N_4116,N_4397);
or U4787 (N_4787,N_4189,N_4449);
xor U4788 (N_4788,N_4028,N_4406);
nor U4789 (N_4789,N_4159,N_4495);
or U4790 (N_4790,N_4330,N_4285);
and U4791 (N_4791,N_4457,N_4170);
nand U4792 (N_4792,N_4388,N_4255);
xor U4793 (N_4793,N_4030,N_4332);
and U4794 (N_4794,N_4390,N_4155);
nor U4795 (N_4795,N_4381,N_4329);
nor U4796 (N_4796,N_4307,N_4048);
and U4797 (N_4797,N_4239,N_4233);
or U4798 (N_4798,N_4379,N_4413);
nand U4799 (N_4799,N_4142,N_4208);
and U4800 (N_4800,N_4013,N_4107);
nand U4801 (N_4801,N_4395,N_4412);
nand U4802 (N_4802,N_4314,N_4262);
or U4803 (N_4803,N_4036,N_4082);
and U4804 (N_4804,N_4185,N_4191);
or U4805 (N_4805,N_4347,N_4239);
nor U4806 (N_4806,N_4472,N_4245);
nor U4807 (N_4807,N_4289,N_4326);
xnor U4808 (N_4808,N_4400,N_4196);
and U4809 (N_4809,N_4098,N_4154);
xnor U4810 (N_4810,N_4043,N_4403);
nor U4811 (N_4811,N_4185,N_4167);
nand U4812 (N_4812,N_4418,N_4277);
nand U4813 (N_4813,N_4105,N_4031);
nor U4814 (N_4814,N_4173,N_4402);
nand U4815 (N_4815,N_4383,N_4236);
xnor U4816 (N_4816,N_4469,N_4185);
nor U4817 (N_4817,N_4474,N_4067);
nor U4818 (N_4818,N_4197,N_4155);
and U4819 (N_4819,N_4493,N_4064);
xnor U4820 (N_4820,N_4230,N_4498);
nand U4821 (N_4821,N_4324,N_4460);
and U4822 (N_4822,N_4009,N_4331);
xnor U4823 (N_4823,N_4046,N_4090);
or U4824 (N_4824,N_4398,N_4410);
or U4825 (N_4825,N_4056,N_4343);
or U4826 (N_4826,N_4206,N_4073);
or U4827 (N_4827,N_4172,N_4021);
or U4828 (N_4828,N_4406,N_4147);
or U4829 (N_4829,N_4202,N_4013);
nand U4830 (N_4830,N_4152,N_4255);
and U4831 (N_4831,N_4259,N_4152);
and U4832 (N_4832,N_4034,N_4116);
xor U4833 (N_4833,N_4332,N_4440);
and U4834 (N_4834,N_4002,N_4042);
xor U4835 (N_4835,N_4190,N_4292);
nand U4836 (N_4836,N_4364,N_4336);
nor U4837 (N_4837,N_4466,N_4486);
and U4838 (N_4838,N_4169,N_4204);
xor U4839 (N_4839,N_4215,N_4353);
and U4840 (N_4840,N_4405,N_4325);
or U4841 (N_4841,N_4231,N_4018);
nand U4842 (N_4842,N_4036,N_4168);
xor U4843 (N_4843,N_4284,N_4047);
and U4844 (N_4844,N_4056,N_4462);
or U4845 (N_4845,N_4012,N_4063);
or U4846 (N_4846,N_4363,N_4027);
nand U4847 (N_4847,N_4163,N_4011);
nand U4848 (N_4848,N_4075,N_4155);
nor U4849 (N_4849,N_4198,N_4042);
nor U4850 (N_4850,N_4375,N_4097);
nor U4851 (N_4851,N_4250,N_4331);
xor U4852 (N_4852,N_4021,N_4278);
and U4853 (N_4853,N_4416,N_4341);
nor U4854 (N_4854,N_4059,N_4195);
nand U4855 (N_4855,N_4431,N_4231);
and U4856 (N_4856,N_4219,N_4141);
or U4857 (N_4857,N_4022,N_4089);
nor U4858 (N_4858,N_4484,N_4151);
or U4859 (N_4859,N_4094,N_4129);
or U4860 (N_4860,N_4312,N_4364);
or U4861 (N_4861,N_4306,N_4067);
xnor U4862 (N_4862,N_4009,N_4080);
or U4863 (N_4863,N_4439,N_4077);
nor U4864 (N_4864,N_4201,N_4260);
and U4865 (N_4865,N_4265,N_4429);
xnor U4866 (N_4866,N_4247,N_4331);
nor U4867 (N_4867,N_4126,N_4313);
xnor U4868 (N_4868,N_4085,N_4356);
nor U4869 (N_4869,N_4235,N_4394);
nand U4870 (N_4870,N_4114,N_4176);
xor U4871 (N_4871,N_4092,N_4062);
nor U4872 (N_4872,N_4039,N_4271);
or U4873 (N_4873,N_4212,N_4364);
and U4874 (N_4874,N_4345,N_4462);
or U4875 (N_4875,N_4305,N_4402);
nor U4876 (N_4876,N_4202,N_4187);
and U4877 (N_4877,N_4187,N_4353);
xnor U4878 (N_4878,N_4469,N_4042);
nor U4879 (N_4879,N_4072,N_4056);
nor U4880 (N_4880,N_4083,N_4211);
xnor U4881 (N_4881,N_4076,N_4279);
nor U4882 (N_4882,N_4251,N_4279);
nand U4883 (N_4883,N_4179,N_4405);
nor U4884 (N_4884,N_4484,N_4204);
xor U4885 (N_4885,N_4010,N_4351);
or U4886 (N_4886,N_4232,N_4102);
and U4887 (N_4887,N_4073,N_4275);
xor U4888 (N_4888,N_4212,N_4116);
nor U4889 (N_4889,N_4138,N_4208);
nand U4890 (N_4890,N_4114,N_4401);
xor U4891 (N_4891,N_4411,N_4133);
nor U4892 (N_4892,N_4498,N_4436);
or U4893 (N_4893,N_4384,N_4158);
and U4894 (N_4894,N_4152,N_4217);
or U4895 (N_4895,N_4364,N_4078);
or U4896 (N_4896,N_4374,N_4047);
or U4897 (N_4897,N_4121,N_4079);
and U4898 (N_4898,N_4099,N_4295);
or U4899 (N_4899,N_4125,N_4331);
and U4900 (N_4900,N_4385,N_4407);
or U4901 (N_4901,N_4108,N_4208);
or U4902 (N_4902,N_4416,N_4332);
nor U4903 (N_4903,N_4149,N_4494);
nor U4904 (N_4904,N_4404,N_4273);
nor U4905 (N_4905,N_4337,N_4342);
and U4906 (N_4906,N_4318,N_4449);
nor U4907 (N_4907,N_4075,N_4436);
and U4908 (N_4908,N_4151,N_4095);
nand U4909 (N_4909,N_4487,N_4358);
or U4910 (N_4910,N_4428,N_4116);
or U4911 (N_4911,N_4114,N_4416);
xor U4912 (N_4912,N_4270,N_4430);
xnor U4913 (N_4913,N_4370,N_4430);
and U4914 (N_4914,N_4022,N_4069);
xor U4915 (N_4915,N_4222,N_4265);
and U4916 (N_4916,N_4089,N_4001);
and U4917 (N_4917,N_4234,N_4289);
nand U4918 (N_4918,N_4109,N_4492);
and U4919 (N_4919,N_4191,N_4125);
xor U4920 (N_4920,N_4438,N_4325);
nor U4921 (N_4921,N_4271,N_4342);
or U4922 (N_4922,N_4027,N_4435);
xnor U4923 (N_4923,N_4263,N_4181);
or U4924 (N_4924,N_4395,N_4018);
xor U4925 (N_4925,N_4289,N_4284);
nor U4926 (N_4926,N_4422,N_4101);
nand U4927 (N_4927,N_4079,N_4026);
or U4928 (N_4928,N_4274,N_4007);
xnor U4929 (N_4929,N_4289,N_4195);
and U4930 (N_4930,N_4282,N_4455);
xnor U4931 (N_4931,N_4064,N_4410);
nor U4932 (N_4932,N_4211,N_4305);
nand U4933 (N_4933,N_4008,N_4337);
nand U4934 (N_4934,N_4120,N_4412);
nor U4935 (N_4935,N_4114,N_4422);
and U4936 (N_4936,N_4215,N_4037);
nand U4937 (N_4937,N_4419,N_4447);
and U4938 (N_4938,N_4029,N_4000);
xor U4939 (N_4939,N_4368,N_4119);
and U4940 (N_4940,N_4289,N_4257);
and U4941 (N_4941,N_4329,N_4171);
nand U4942 (N_4942,N_4456,N_4042);
or U4943 (N_4943,N_4367,N_4376);
or U4944 (N_4944,N_4129,N_4018);
or U4945 (N_4945,N_4301,N_4037);
and U4946 (N_4946,N_4282,N_4303);
or U4947 (N_4947,N_4415,N_4236);
nand U4948 (N_4948,N_4340,N_4044);
and U4949 (N_4949,N_4395,N_4102);
xnor U4950 (N_4950,N_4478,N_4045);
nor U4951 (N_4951,N_4155,N_4000);
or U4952 (N_4952,N_4171,N_4247);
nand U4953 (N_4953,N_4084,N_4425);
xnor U4954 (N_4954,N_4467,N_4242);
nor U4955 (N_4955,N_4117,N_4485);
nor U4956 (N_4956,N_4201,N_4097);
or U4957 (N_4957,N_4204,N_4049);
and U4958 (N_4958,N_4093,N_4375);
nor U4959 (N_4959,N_4364,N_4022);
or U4960 (N_4960,N_4435,N_4251);
xnor U4961 (N_4961,N_4334,N_4315);
nand U4962 (N_4962,N_4402,N_4207);
nand U4963 (N_4963,N_4382,N_4221);
nand U4964 (N_4964,N_4036,N_4286);
xor U4965 (N_4965,N_4228,N_4348);
or U4966 (N_4966,N_4306,N_4106);
nor U4967 (N_4967,N_4235,N_4101);
nand U4968 (N_4968,N_4079,N_4071);
or U4969 (N_4969,N_4350,N_4291);
and U4970 (N_4970,N_4292,N_4024);
or U4971 (N_4971,N_4168,N_4127);
xnor U4972 (N_4972,N_4443,N_4062);
and U4973 (N_4973,N_4288,N_4164);
nor U4974 (N_4974,N_4145,N_4419);
nand U4975 (N_4975,N_4223,N_4041);
nor U4976 (N_4976,N_4210,N_4258);
xor U4977 (N_4977,N_4407,N_4349);
nor U4978 (N_4978,N_4261,N_4162);
nand U4979 (N_4979,N_4290,N_4020);
nand U4980 (N_4980,N_4475,N_4202);
nor U4981 (N_4981,N_4023,N_4244);
xnor U4982 (N_4982,N_4269,N_4137);
and U4983 (N_4983,N_4306,N_4062);
or U4984 (N_4984,N_4229,N_4011);
or U4985 (N_4985,N_4050,N_4357);
or U4986 (N_4986,N_4077,N_4007);
nor U4987 (N_4987,N_4083,N_4168);
or U4988 (N_4988,N_4426,N_4251);
xnor U4989 (N_4989,N_4251,N_4440);
nand U4990 (N_4990,N_4003,N_4233);
xor U4991 (N_4991,N_4437,N_4446);
and U4992 (N_4992,N_4060,N_4009);
nand U4993 (N_4993,N_4224,N_4436);
and U4994 (N_4994,N_4349,N_4132);
or U4995 (N_4995,N_4334,N_4182);
nor U4996 (N_4996,N_4186,N_4215);
nor U4997 (N_4997,N_4280,N_4299);
nand U4998 (N_4998,N_4343,N_4371);
and U4999 (N_4999,N_4495,N_4141);
or UO_0 (O_0,N_4644,N_4953);
and UO_1 (O_1,N_4944,N_4979);
xnor UO_2 (O_2,N_4878,N_4701);
nor UO_3 (O_3,N_4886,N_4899);
xnor UO_4 (O_4,N_4880,N_4661);
nand UO_5 (O_5,N_4856,N_4768);
nor UO_6 (O_6,N_4746,N_4585);
or UO_7 (O_7,N_4818,N_4958);
or UO_8 (O_8,N_4674,N_4857);
and UO_9 (O_9,N_4813,N_4535);
xnor UO_10 (O_10,N_4702,N_4828);
or UO_11 (O_11,N_4714,N_4942);
nand UO_12 (O_12,N_4816,N_4810);
xnor UO_13 (O_13,N_4735,N_4935);
nand UO_14 (O_14,N_4665,N_4937);
nand UO_15 (O_15,N_4614,N_4564);
nor UO_16 (O_16,N_4704,N_4550);
nand UO_17 (O_17,N_4545,N_4985);
nand UO_18 (O_18,N_4582,N_4802);
nand UO_19 (O_19,N_4770,N_4515);
xor UO_20 (O_20,N_4962,N_4949);
nor UO_21 (O_21,N_4910,N_4596);
or UO_22 (O_22,N_4754,N_4991);
or UO_23 (O_23,N_4806,N_4881);
xor UO_24 (O_24,N_4697,N_4694);
xor UO_25 (O_25,N_4939,N_4821);
nor UO_26 (O_26,N_4926,N_4845);
or UO_27 (O_27,N_4874,N_4593);
nor UO_28 (O_28,N_4727,N_4931);
and UO_29 (O_29,N_4509,N_4505);
or UO_30 (O_30,N_4833,N_4922);
or UO_31 (O_31,N_4634,N_4521);
nand UO_32 (O_32,N_4963,N_4927);
or UO_33 (O_33,N_4720,N_4996);
nor UO_34 (O_34,N_4795,N_4978);
nand UO_35 (O_35,N_4882,N_4724);
nor UO_36 (O_36,N_4676,N_4965);
xnor UO_37 (O_37,N_4640,N_4796);
xnor UO_38 (O_38,N_4742,N_4752);
nand UO_39 (O_39,N_4906,N_4506);
xnor UO_40 (O_40,N_4737,N_4892);
xnor UO_41 (O_41,N_4688,N_4663);
nand UO_42 (O_42,N_4623,N_4872);
and UO_43 (O_43,N_4554,N_4980);
nor UO_44 (O_44,N_4556,N_4863);
or UO_45 (O_45,N_4745,N_4683);
and UO_46 (O_46,N_4586,N_4771);
or UO_47 (O_47,N_4969,N_4827);
nor UO_48 (O_48,N_4527,N_4528);
xor UO_49 (O_49,N_4900,N_4998);
xor UO_50 (O_50,N_4743,N_4782);
and UO_51 (O_51,N_4595,N_4598);
nor UO_52 (O_52,N_4657,N_4534);
or UO_53 (O_53,N_4839,N_4921);
nor UO_54 (O_54,N_4519,N_4594);
nor UO_55 (O_55,N_4639,N_4992);
or UO_56 (O_56,N_4936,N_4559);
or UO_57 (O_57,N_4600,N_4808);
nor UO_58 (O_58,N_4798,N_4797);
xor UO_59 (O_59,N_4897,N_4565);
or UO_60 (O_60,N_4829,N_4893);
xnor UO_61 (O_61,N_4999,N_4615);
or UO_62 (O_62,N_4525,N_4577);
and UO_63 (O_63,N_4987,N_4579);
and UO_64 (O_64,N_4954,N_4636);
nand UO_65 (O_65,N_4885,N_4952);
nor UO_66 (O_66,N_4513,N_4898);
nand UO_67 (O_67,N_4873,N_4604);
xnor UO_68 (O_68,N_4659,N_4756);
or UO_69 (O_69,N_4786,N_4599);
xnor UO_70 (O_70,N_4819,N_4609);
nand UO_71 (O_71,N_4847,N_4738);
nor UO_72 (O_72,N_4911,N_4864);
nand UO_73 (O_73,N_4726,N_4672);
nand UO_74 (O_74,N_4540,N_4989);
xor UO_75 (O_75,N_4976,N_4817);
or UO_76 (O_76,N_4658,N_4859);
and UO_77 (O_77,N_4971,N_4631);
nand UO_78 (O_78,N_4822,N_4815);
nand UO_79 (O_79,N_4778,N_4700);
nor UO_80 (O_80,N_4627,N_4502);
xor UO_81 (O_81,N_4500,N_4736);
and UO_82 (O_82,N_4809,N_4645);
or UO_83 (O_83,N_4924,N_4616);
nand UO_84 (O_84,N_4875,N_4548);
xnor UO_85 (O_85,N_4919,N_4673);
xor UO_86 (O_86,N_4917,N_4753);
nand UO_87 (O_87,N_4708,N_4836);
or UO_88 (O_88,N_4587,N_4693);
xor UO_89 (O_89,N_4824,N_4703);
or UO_90 (O_90,N_4914,N_4547);
nand UO_91 (O_91,N_4781,N_4890);
and UO_92 (O_92,N_4717,N_4628);
and UO_93 (O_93,N_4887,N_4855);
xor UO_94 (O_94,N_4622,N_4920);
and UO_95 (O_95,N_4718,N_4643);
or UO_96 (O_96,N_4748,N_4687);
nand UO_97 (O_97,N_4516,N_4504);
nor UO_98 (O_98,N_4961,N_4651);
nand UO_99 (O_99,N_4997,N_4633);
or UO_100 (O_100,N_4626,N_4517);
xnor UO_101 (O_101,N_4621,N_4532);
or UO_102 (O_102,N_4852,N_4563);
nor UO_103 (O_103,N_4762,N_4901);
and UO_104 (O_104,N_4758,N_4749);
nor UO_105 (O_105,N_4649,N_4733);
or UO_106 (O_106,N_4514,N_4512);
nor UO_107 (O_107,N_4576,N_4529);
nand UO_108 (O_108,N_4837,N_4705);
xnor UO_109 (O_109,N_4902,N_4788);
xnor UO_110 (O_110,N_4680,N_4841);
nand UO_111 (O_111,N_4934,N_4677);
nand UO_112 (O_112,N_4566,N_4699);
and UO_113 (O_113,N_4842,N_4889);
xnor UO_114 (O_114,N_4690,N_4904);
or UO_115 (O_115,N_4713,N_4843);
nand UO_116 (O_116,N_4691,N_4611);
nor UO_117 (O_117,N_4530,N_4570);
nand UO_118 (O_118,N_4790,N_4930);
nand UO_119 (O_119,N_4666,N_4789);
and UO_120 (O_120,N_4617,N_4950);
nor UO_121 (O_121,N_4544,N_4712);
or UO_122 (O_122,N_4832,N_4946);
nor UO_123 (O_123,N_4812,N_4807);
xnor UO_124 (O_124,N_4648,N_4723);
nand UO_125 (O_125,N_4698,N_4728);
nand UO_126 (O_126,N_4792,N_4896);
xnor UO_127 (O_127,N_4861,N_4522);
nand UO_128 (O_128,N_4603,N_4725);
nor UO_129 (O_129,N_4618,N_4681);
xnor UO_130 (O_130,N_4959,N_4684);
nor UO_131 (O_131,N_4814,N_4630);
nand UO_132 (O_132,N_4629,N_4981);
and UO_133 (O_133,N_4820,N_4755);
xnor UO_134 (O_134,N_4686,N_4669);
or UO_135 (O_135,N_4908,N_4637);
xor UO_136 (O_136,N_4647,N_4675);
nand UO_137 (O_137,N_4578,N_4909);
nand UO_138 (O_138,N_4835,N_4549);
and UO_139 (O_139,N_4562,N_4850);
nor UO_140 (O_140,N_4734,N_4923);
nor UO_141 (O_141,N_4763,N_4772);
and UO_142 (O_142,N_4776,N_4865);
nor UO_143 (O_143,N_4538,N_4613);
and UO_144 (O_144,N_4635,N_4523);
xnor UO_145 (O_145,N_4511,N_4769);
or UO_146 (O_146,N_4891,N_4866);
xnor UO_147 (O_147,N_4805,N_4883);
or UO_148 (O_148,N_4664,N_4995);
nand UO_149 (O_149,N_4912,N_4905);
nand UO_150 (O_150,N_4853,N_4597);
xnor UO_151 (O_151,N_4552,N_4916);
nor UO_152 (O_152,N_4652,N_4794);
nand UO_153 (O_153,N_4612,N_4844);
nand UO_154 (O_154,N_4678,N_4834);
or UO_155 (O_155,N_4524,N_4888);
nor UO_156 (O_156,N_4846,N_4561);
nor UO_157 (O_157,N_4574,N_4793);
or UO_158 (O_158,N_4876,N_4619);
and UO_159 (O_159,N_4695,N_4765);
and UO_160 (O_160,N_4947,N_4966);
nand UO_161 (O_161,N_4767,N_4867);
and UO_162 (O_162,N_4986,N_4655);
and UO_163 (O_163,N_4840,N_4641);
nand UO_164 (O_164,N_4968,N_4716);
and UO_165 (O_165,N_4801,N_4941);
nor UO_166 (O_166,N_4779,N_4766);
and UO_167 (O_167,N_4868,N_4625);
xnor UO_168 (O_168,N_4870,N_4775);
xor UO_169 (O_169,N_4601,N_4967);
nand UO_170 (O_170,N_4670,N_4879);
nor UO_171 (O_171,N_4903,N_4974);
or UO_172 (O_172,N_4508,N_4803);
xor UO_173 (O_173,N_4606,N_4668);
or UO_174 (O_174,N_4546,N_4571);
xnor UO_175 (O_175,N_4929,N_4589);
and UO_176 (O_176,N_4884,N_4719);
or UO_177 (O_177,N_4825,N_4679);
or UO_178 (O_178,N_4972,N_4730);
nor UO_179 (O_179,N_4860,N_4682);
xor UO_180 (O_180,N_4895,N_4588);
nor UO_181 (O_181,N_4761,N_4849);
nor UO_182 (O_182,N_4984,N_4973);
nand UO_183 (O_183,N_4709,N_4542);
and UO_184 (O_184,N_4804,N_4575);
or UO_185 (O_185,N_4988,N_4646);
xnor UO_186 (O_186,N_4791,N_4707);
or UO_187 (O_187,N_4933,N_4940);
xor UO_188 (O_188,N_4696,N_4759);
and UO_189 (O_189,N_4894,N_4826);
and UO_190 (O_190,N_4654,N_4948);
xnor UO_191 (O_191,N_4799,N_4955);
nand UO_192 (O_192,N_4581,N_4610);
nor UO_193 (O_193,N_4572,N_4518);
or UO_194 (O_194,N_4994,N_4848);
or UO_195 (O_195,N_4932,N_4671);
nor UO_196 (O_196,N_4584,N_4854);
or UO_197 (O_197,N_4590,N_4957);
or UO_198 (O_198,N_4975,N_4568);
and UO_199 (O_199,N_4773,N_4977);
or UO_200 (O_200,N_4993,N_4928);
or UO_201 (O_201,N_4722,N_4938);
nor UO_202 (O_202,N_4871,N_4862);
or UO_203 (O_203,N_4560,N_4915);
nand UO_204 (O_204,N_4787,N_4732);
xor UO_205 (O_205,N_4777,N_4638);
nor UO_206 (O_206,N_4710,N_4592);
xor UO_207 (O_207,N_4877,N_4501);
or UO_208 (O_208,N_4558,N_4608);
xor UO_209 (O_209,N_4751,N_4925);
and UO_210 (O_210,N_4520,N_4650);
and UO_211 (O_211,N_4536,N_4757);
and UO_212 (O_212,N_4685,N_4780);
and UO_213 (O_213,N_4945,N_4533);
xnor UO_214 (O_214,N_4739,N_4800);
nand UO_215 (O_215,N_4667,N_4569);
nand UO_216 (O_216,N_4731,N_4830);
or UO_217 (O_217,N_4750,N_4591);
nand UO_218 (O_218,N_4602,N_4783);
or UO_219 (O_219,N_4831,N_4531);
nor UO_220 (O_220,N_4541,N_4721);
and UO_221 (O_221,N_4960,N_4811);
and UO_222 (O_222,N_4573,N_4692);
nor UO_223 (O_223,N_4715,N_4526);
nand UO_224 (O_224,N_4706,N_4620);
and UO_225 (O_225,N_4764,N_4553);
nand UO_226 (O_226,N_4760,N_4983);
xor UO_227 (O_227,N_4607,N_4990);
or UO_228 (O_228,N_4580,N_4656);
or UO_229 (O_229,N_4583,N_4740);
or UO_230 (O_230,N_4784,N_4662);
nor UO_231 (O_231,N_4543,N_4913);
and UO_232 (O_232,N_4823,N_4907);
nor UO_233 (O_233,N_4982,N_4943);
and UO_234 (O_234,N_4642,N_4747);
xor UO_235 (O_235,N_4970,N_4539);
xor UO_236 (O_236,N_4838,N_4858);
xor UO_237 (O_237,N_4624,N_4537);
and UO_238 (O_238,N_4785,N_4503);
or UO_239 (O_239,N_4964,N_4567);
nand UO_240 (O_240,N_4510,N_4774);
xor UO_241 (O_241,N_4660,N_4632);
nand UO_242 (O_242,N_4729,N_4869);
xnor UO_243 (O_243,N_4851,N_4507);
xnor UO_244 (O_244,N_4956,N_4551);
and UO_245 (O_245,N_4741,N_4557);
or UO_246 (O_246,N_4951,N_4689);
nand UO_247 (O_247,N_4918,N_4555);
xor UO_248 (O_248,N_4653,N_4711);
and UO_249 (O_249,N_4744,N_4605);
xor UO_250 (O_250,N_4843,N_4766);
nand UO_251 (O_251,N_4589,N_4825);
nor UO_252 (O_252,N_4858,N_4881);
or UO_253 (O_253,N_4634,N_4578);
or UO_254 (O_254,N_4973,N_4719);
nor UO_255 (O_255,N_4710,N_4790);
nor UO_256 (O_256,N_4740,N_4784);
or UO_257 (O_257,N_4691,N_4944);
nor UO_258 (O_258,N_4650,N_4684);
and UO_259 (O_259,N_4957,N_4576);
nor UO_260 (O_260,N_4995,N_4908);
xor UO_261 (O_261,N_4880,N_4987);
nor UO_262 (O_262,N_4561,N_4643);
nor UO_263 (O_263,N_4741,N_4777);
nor UO_264 (O_264,N_4599,N_4549);
xnor UO_265 (O_265,N_4581,N_4541);
nand UO_266 (O_266,N_4830,N_4715);
and UO_267 (O_267,N_4628,N_4857);
nor UO_268 (O_268,N_4996,N_4820);
nand UO_269 (O_269,N_4709,N_4883);
and UO_270 (O_270,N_4921,N_4668);
nand UO_271 (O_271,N_4878,N_4752);
and UO_272 (O_272,N_4591,N_4652);
nand UO_273 (O_273,N_4671,N_4747);
nor UO_274 (O_274,N_4677,N_4693);
xnor UO_275 (O_275,N_4956,N_4838);
or UO_276 (O_276,N_4615,N_4726);
nand UO_277 (O_277,N_4832,N_4981);
or UO_278 (O_278,N_4912,N_4571);
xor UO_279 (O_279,N_4843,N_4669);
and UO_280 (O_280,N_4677,N_4973);
and UO_281 (O_281,N_4859,N_4978);
xor UO_282 (O_282,N_4712,N_4566);
nor UO_283 (O_283,N_4898,N_4906);
nor UO_284 (O_284,N_4932,N_4595);
or UO_285 (O_285,N_4632,N_4937);
xor UO_286 (O_286,N_4671,N_4781);
and UO_287 (O_287,N_4977,N_4812);
nand UO_288 (O_288,N_4758,N_4579);
nand UO_289 (O_289,N_4819,N_4728);
nand UO_290 (O_290,N_4700,N_4701);
nand UO_291 (O_291,N_4955,N_4679);
nand UO_292 (O_292,N_4888,N_4716);
xor UO_293 (O_293,N_4746,N_4511);
nor UO_294 (O_294,N_4667,N_4680);
xor UO_295 (O_295,N_4831,N_4643);
or UO_296 (O_296,N_4708,N_4724);
or UO_297 (O_297,N_4749,N_4956);
nor UO_298 (O_298,N_4954,N_4578);
or UO_299 (O_299,N_4792,N_4815);
and UO_300 (O_300,N_4638,N_4552);
nand UO_301 (O_301,N_4700,N_4510);
nor UO_302 (O_302,N_4637,N_4808);
nor UO_303 (O_303,N_4928,N_4731);
nand UO_304 (O_304,N_4830,N_4661);
or UO_305 (O_305,N_4644,N_4802);
or UO_306 (O_306,N_4592,N_4769);
or UO_307 (O_307,N_4790,N_4630);
nor UO_308 (O_308,N_4954,N_4920);
xor UO_309 (O_309,N_4575,N_4784);
or UO_310 (O_310,N_4838,N_4545);
xnor UO_311 (O_311,N_4639,N_4861);
nand UO_312 (O_312,N_4500,N_4807);
or UO_313 (O_313,N_4587,N_4988);
nor UO_314 (O_314,N_4598,N_4809);
nand UO_315 (O_315,N_4624,N_4958);
xor UO_316 (O_316,N_4612,N_4853);
xnor UO_317 (O_317,N_4875,N_4777);
nor UO_318 (O_318,N_4719,N_4601);
nor UO_319 (O_319,N_4769,N_4595);
nand UO_320 (O_320,N_4938,N_4975);
nand UO_321 (O_321,N_4573,N_4732);
nor UO_322 (O_322,N_4857,N_4503);
and UO_323 (O_323,N_4857,N_4690);
nor UO_324 (O_324,N_4893,N_4654);
nand UO_325 (O_325,N_4933,N_4880);
nor UO_326 (O_326,N_4849,N_4925);
or UO_327 (O_327,N_4514,N_4755);
and UO_328 (O_328,N_4896,N_4997);
nor UO_329 (O_329,N_4800,N_4605);
nor UO_330 (O_330,N_4938,N_4868);
and UO_331 (O_331,N_4799,N_4947);
nand UO_332 (O_332,N_4652,N_4974);
and UO_333 (O_333,N_4594,N_4588);
nor UO_334 (O_334,N_4856,N_4879);
xor UO_335 (O_335,N_4562,N_4828);
xor UO_336 (O_336,N_4996,N_4591);
nor UO_337 (O_337,N_4824,N_4608);
nor UO_338 (O_338,N_4885,N_4892);
nor UO_339 (O_339,N_4586,N_4686);
and UO_340 (O_340,N_4845,N_4703);
and UO_341 (O_341,N_4794,N_4991);
nor UO_342 (O_342,N_4817,N_4679);
nor UO_343 (O_343,N_4894,N_4699);
and UO_344 (O_344,N_4727,N_4556);
nand UO_345 (O_345,N_4943,N_4667);
and UO_346 (O_346,N_4518,N_4975);
or UO_347 (O_347,N_4744,N_4914);
xnor UO_348 (O_348,N_4523,N_4703);
and UO_349 (O_349,N_4886,N_4903);
and UO_350 (O_350,N_4772,N_4746);
nor UO_351 (O_351,N_4646,N_4578);
nand UO_352 (O_352,N_4532,N_4700);
nand UO_353 (O_353,N_4993,N_4530);
xor UO_354 (O_354,N_4574,N_4827);
nand UO_355 (O_355,N_4939,N_4953);
nor UO_356 (O_356,N_4950,N_4942);
xor UO_357 (O_357,N_4977,N_4506);
or UO_358 (O_358,N_4788,N_4598);
xnor UO_359 (O_359,N_4936,N_4733);
or UO_360 (O_360,N_4659,N_4676);
and UO_361 (O_361,N_4879,N_4570);
nand UO_362 (O_362,N_4681,N_4866);
nand UO_363 (O_363,N_4992,N_4758);
and UO_364 (O_364,N_4845,N_4586);
or UO_365 (O_365,N_4612,N_4806);
nor UO_366 (O_366,N_4922,N_4971);
xor UO_367 (O_367,N_4957,N_4572);
xor UO_368 (O_368,N_4656,N_4651);
and UO_369 (O_369,N_4920,N_4990);
nand UO_370 (O_370,N_4587,N_4934);
xnor UO_371 (O_371,N_4685,N_4691);
nand UO_372 (O_372,N_4926,N_4518);
xor UO_373 (O_373,N_4620,N_4753);
xor UO_374 (O_374,N_4840,N_4515);
nor UO_375 (O_375,N_4747,N_4854);
nor UO_376 (O_376,N_4906,N_4597);
and UO_377 (O_377,N_4686,N_4633);
nor UO_378 (O_378,N_4722,N_4986);
and UO_379 (O_379,N_4592,N_4616);
or UO_380 (O_380,N_4622,N_4771);
nand UO_381 (O_381,N_4586,N_4507);
nor UO_382 (O_382,N_4600,N_4547);
nand UO_383 (O_383,N_4982,N_4892);
or UO_384 (O_384,N_4615,N_4831);
and UO_385 (O_385,N_4888,N_4659);
and UO_386 (O_386,N_4862,N_4910);
or UO_387 (O_387,N_4535,N_4935);
nor UO_388 (O_388,N_4538,N_4773);
nand UO_389 (O_389,N_4503,N_4689);
nand UO_390 (O_390,N_4514,N_4572);
and UO_391 (O_391,N_4756,N_4590);
and UO_392 (O_392,N_4722,N_4760);
xnor UO_393 (O_393,N_4980,N_4593);
nand UO_394 (O_394,N_4697,N_4647);
xor UO_395 (O_395,N_4610,N_4628);
xnor UO_396 (O_396,N_4891,N_4584);
xor UO_397 (O_397,N_4699,N_4926);
xnor UO_398 (O_398,N_4801,N_4556);
nand UO_399 (O_399,N_4715,N_4591);
and UO_400 (O_400,N_4638,N_4779);
nand UO_401 (O_401,N_4597,N_4588);
or UO_402 (O_402,N_4661,N_4747);
xor UO_403 (O_403,N_4539,N_4689);
xor UO_404 (O_404,N_4549,N_4926);
and UO_405 (O_405,N_4867,N_4769);
or UO_406 (O_406,N_4547,N_4596);
and UO_407 (O_407,N_4863,N_4807);
xor UO_408 (O_408,N_4942,N_4740);
xor UO_409 (O_409,N_4793,N_4884);
nand UO_410 (O_410,N_4966,N_4908);
or UO_411 (O_411,N_4962,N_4521);
xnor UO_412 (O_412,N_4801,N_4799);
or UO_413 (O_413,N_4716,N_4544);
nor UO_414 (O_414,N_4755,N_4718);
xor UO_415 (O_415,N_4847,N_4902);
nor UO_416 (O_416,N_4677,N_4536);
and UO_417 (O_417,N_4733,N_4708);
and UO_418 (O_418,N_4853,N_4594);
nand UO_419 (O_419,N_4633,N_4536);
xnor UO_420 (O_420,N_4883,N_4510);
nand UO_421 (O_421,N_4763,N_4661);
or UO_422 (O_422,N_4516,N_4894);
nand UO_423 (O_423,N_4788,N_4573);
xor UO_424 (O_424,N_4882,N_4887);
nor UO_425 (O_425,N_4900,N_4838);
nor UO_426 (O_426,N_4678,N_4602);
nand UO_427 (O_427,N_4617,N_4584);
xor UO_428 (O_428,N_4500,N_4877);
or UO_429 (O_429,N_4501,N_4572);
or UO_430 (O_430,N_4765,N_4845);
or UO_431 (O_431,N_4980,N_4618);
nor UO_432 (O_432,N_4908,N_4920);
or UO_433 (O_433,N_4785,N_4702);
and UO_434 (O_434,N_4632,N_4930);
or UO_435 (O_435,N_4898,N_4612);
and UO_436 (O_436,N_4545,N_4915);
nand UO_437 (O_437,N_4681,N_4748);
xor UO_438 (O_438,N_4617,N_4943);
nand UO_439 (O_439,N_4540,N_4823);
or UO_440 (O_440,N_4761,N_4982);
nor UO_441 (O_441,N_4574,N_4603);
xnor UO_442 (O_442,N_4720,N_4505);
or UO_443 (O_443,N_4998,N_4525);
nor UO_444 (O_444,N_4548,N_4613);
nand UO_445 (O_445,N_4502,N_4894);
nor UO_446 (O_446,N_4693,N_4829);
nand UO_447 (O_447,N_4752,N_4903);
xnor UO_448 (O_448,N_4777,N_4874);
nand UO_449 (O_449,N_4736,N_4788);
and UO_450 (O_450,N_4970,N_4815);
xor UO_451 (O_451,N_4505,N_4649);
nand UO_452 (O_452,N_4589,N_4666);
and UO_453 (O_453,N_4930,N_4974);
xor UO_454 (O_454,N_4862,N_4599);
or UO_455 (O_455,N_4666,N_4821);
xor UO_456 (O_456,N_4737,N_4533);
nor UO_457 (O_457,N_4739,N_4765);
or UO_458 (O_458,N_4905,N_4991);
nor UO_459 (O_459,N_4655,N_4878);
xor UO_460 (O_460,N_4752,N_4672);
and UO_461 (O_461,N_4784,N_4626);
nor UO_462 (O_462,N_4548,N_4526);
and UO_463 (O_463,N_4767,N_4993);
nor UO_464 (O_464,N_4701,N_4595);
nand UO_465 (O_465,N_4501,N_4550);
nor UO_466 (O_466,N_4580,N_4889);
or UO_467 (O_467,N_4540,N_4831);
nand UO_468 (O_468,N_4773,N_4736);
nor UO_469 (O_469,N_4818,N_4560);
or UO_470 (O_470,N_4927,N_4577);
nand UO_471 (O_471,N_4981,N_4817);
xnor UO_472 (O_472,N_4985,N_4651);
or UO_473 (O_473,N_4767,N_4542);
nor UO_474 (O_474,N_4529,N_4947);
nor UO_475 (O_475,N_4793,N_4983);
and UO_476 (O_476,N_4635,N_4865);
and UO_477 (O_477,N_4820,N_4532);
and UO_478 (O_478,N_4960,N_4835);
or UO_479 (O_479,N_4555,N_4972);
nor UO_480 (O_480,N_4730,N_4563);
and UO_481 (O_481,N_4603,N_4660);
nor UO_482 (O_482,N_4816,N_4689);
nand UO_483 (O_483,N_4556,N_4647);
xor UO_484 (O_484,N_4712,N_4920);
nor UO_485 (O_485,N_4782,N_4702);
nand UO_486 (O_486,N_4646,N_4739);
and UO_487 (O_487,N_4552,N_4674);
nor UO_488 (O_488,N_4921,N_4995);
nand UO_489 (O_489,N_4903,N_4910);
nor UO_490 (O_490,N_4891,N_4897);
xnor UO_491 (O_491,N_4839,N_4766);
xor UO_492 (O_492,N_4706,N_4816);
and UO_493 (O_493,N_4954,N_4941);
xnor UO_494 (O_494,N_4693,N_4831);
xnor UO_495 (O_495,N_4922,N_4999);
xor UO_496 (O_496,N_4613,N_4742);
nand UO_497 (O_497,N_4721,N_4753);
nand UO_498 (O_498,N_4619,N_4937);
and UO_499 (O_499,N_4752,N_4885);
and UO_500 (O_500,N_4723,N_4507);
xor UO_501 (O_501,N_4997,N_4637);
nor UO_502 (O_502,N_4788,N_4895);
and UO_503 (O_503,N_4795,N_4684);
and UO_504 (O_504,N_4799,N_4959);
or UO_505 (O_505,N_4646,N_4610);
or UO_506 (O_506,N_4867,N_4666);
xnor UO_507 (O_507,N_4515,N_4718);
xnor UO_508 (O_508,N_4629,N_4709);
xor UO_509 (O_509,N_4784,N_4898);
nand UO_510 (O_510,N_4572,N_4823);
nand UO_511 (O_511,N_4685,N_4511);
or UO_512 (O_512,N_4657,N_4986);
nand UO_513 (O_513,N_4707,N_4852);
or UO_514 (O_514,N_4625,N_4540);
xor UO_515 (O_515,N_4765,N_4961);
nor UO_516 (O_516,N_4771,N_4854);
nand UO_517 (O_517,N_4681,N_4546);
nor UO_518 (O_518,N_4671,N_4588);
nand UO_519 (O_519,N_4955,N_4820);
xor UO_520 (O_520,N_4777,N_4786);
xnor UO_521 (O_521,N_4873,N_4627);
or UO_522 (O_522,N_4600,N_4811);
nor UO_523 (O_523,N_4834,N_4998);
xnor UO_524 (O_524,N_4812,N_4763);
or UO_525 (O_525,N_4702,N_4659);
xnor UO_526 (O_526,N_4578,N_4552);
or UO_527 (O_527,N_4911,N_4891);
and UO_528 (O_528,N_4906,N_4576);
nor UO_529 (O_529,N_4865,N_4828);
and UO_530 (O_530,N_4628,N_4543);
and UO_531 (O_531,N_4960,N_4617);
xnor UO_532 (O_532,N_4554,N_4963);
or UO_533 (O_533,N_4706,N_4659);
xor UO_534 (O_534,N_4768,N_4702);
and UO_535 (O_535,N_4764,N_4737);
xnor UO_536 (O_536,N_4786,N_4998);
and UO_537 (O_537,N_4788,N_4673);
nand UO_538 (O_538,N_4949,N_4558);
or UO_539 (O_539,N_4700,N_4653);
nand UO_540 (O_540,N_4641,N_4853);
nand UO_541 (O_541,N_4669,N_4743);
nand UO_542 (O_542,N_4788,N_4559);
or UO_543 (O_543,N_4849,N_4574);
xnor UO_544 (O_544,N_4989,N_4618);
nand UO_545 (O_545,N_4935,N_4729);
nor UO_546 (O_546,N_4570,N_4752);
nor UO_547 (O_547,N_4586,N_4802);
or UO_548 (O_548,N_4929,N_4595);
xor UO_549 (O_549,N_4628,N_4525);
and UO_550 (O_550,N_4924,N_4852);
xnor UO_551 (O_551,N_4753,N_4942);
xnor UO_552 (O_552,N_4979,N_4915);
xnor UO_553 (O_553,N_4750,N_4918);
or UO_554 (O_554,N_4891,N_4960);
and UO_555 (O_555,N_4527,N_4995);
xnor UO_556 (O_556,N_4637,N_4571);
xnor UO_557 (O_557,N_4989,N_4528);
xor UO_558 (O_558,N_4758,N_4946);
xnor UO_559 (O_559,N_4813,N_4887);
nand UO_560 (O_560,N_4558,N_4668);
nor UO_561 (O_561,N_4872,N_4911);
or UO_562 (O_562,N_4503,N_4696);
xor UO_563 (O_563,N_4998,N_4555);
xor UO_564 (O_564,N_4953,N_4536);
or UO_565 (O_565,N_4852,N_4659);
and UO_566 (O_566,N_4889,N_4535);
nor UO_567 (O_567,N_4799,N_4501);
or UO_568 (O_568,N_4505,N_4699);
and UO_569 (O_569,N_4887,N_4766);
nor UO_570 (O_570,N_4671,N_4982);
and UO_571 (O_571,N_4924,N_4590);
or UO_572 (O_572,N_4912,N_4989);
and UO_573 (O_573,N_4620,N_4847);
xnor UO_574 (O_574,N_4975,N_4881);
and UO_575 (O_575,N_4756,N_4784);
and UO_576 (O_576,N_4853,N_4722);
nor UO_577 (O_577,N_4618,N_4763);
and UO_578 (O_578,N_4698,N_4784);
nand UO_579 (O_579,N_4995,N_4894);
and UO_580 (O_580,N_4898,N_4854);
xnor UO_581 (O_581,N_4657,N_4831);
nor UO_582 (O_582,N_4837,N_4625);
nand UO_583 (O_583,N_4988,N_4591);
and UO_584 (O_584,N_4508,N_4744);
nand UO_585 (O_585,N_4825,N_4968);
nor UO_586 (O_586,N_4721,N_4810);
nand UO_587 (O_587,N_4508,N_4887);
and UO_588 (O_588,N_4892,N_4544);
xnor UO_589 (O_589,N_4557,N_4590);
nand UO_590 (O_590,N_4586,N_4600);
or UO_591 (O_591,N_4682,N_4647);
xor UO_592 (O_592,N_4535,N_4702);
nor UO_593 (O_593,N_4715,N_4908);
xor UO_594 (O_594,N_4859,N_4651);
nor UO_595 (O_595,N_4904,N_4557);
and UO_596 (O_596,N_4522,N_4716);
and UO_597 (O_597,N_4552,N_4520);
or UO_598 (O_598,N_4529,N_4558);
xnor UO_599 (O_599,N_4943,N_4995);
or UO_600 (O_600,N_4553,N_4513);
or UO_601 (O_601,N_4755,N_4702);
nor UO_602 (O_602,N_4685,N_4923);
and UO_603 (O_603,N_4828,N_4791);
xnor UO_604 (O_604,N_4737,N_4541);
xor UO_605 (O_605,N_4540,N_4773);
xor UO_606 (O_606,N_4797,N_4536);
nand UO_607 (O_607,N_4786,N_4657);
nand UO_608 (O_608,N_4844,N_4670);
or UO_609 (O_609,N_4773,N_4771);
or UO_610 (O_610,N_4942,N_4955);
nand UO_611 (O_611,N_4733,N_4697);
xnor UO_612 (O_612,N_4513,N_4545);
or UO_613 (O_613,N_4506,N_4727);
nor UO_614 (O_614,N_4829,N_4830);
or UO_615 (O_615,N_4792,N_4551);
or UO_616 (O_616,N_4621,N_4507);
and UO_617 (O_617,N_4781,N_4611);
or UO_618 (O_618,N_4975,N_4906);
nor UO_619 (O_619,N_4857,N_4899);
xnor UO_620 (O_620,N_4800,N_4755);
nand UO_621 (O_621,N_4828,N_4695);
xor UO_622 (O_622,N_4729,N_4763);
and UO_623 (O_623,N_4744,N_4865);
or UO_624 (O_624,N_4911,N_4923);
nor UO_625 (O_625,N_4515,N_4886);
and UO_626 (O_626,N_4691,N_4529);
nor UO_627 (O_627,N_4554,N_4832);
or UO_628 (O_628,N_4731,N_4773);
or UO_629 (O_629,N_4861,N_4924);
nor UO_630 (O_630,N_4630,N_4956);
or UO_631 (O_631,N_4552,N_4994);
nor UO_632 (O_632,N_4888,N_4555);
nor UO_633 (O_633,N_4913,N_4604);
and UO_634 (O_634,N_4963,N_4812);
nand UO_635 (O_635,N_4784,N_4883);
xor UO_636 (O_636,N_4926,N_4903);
nand UO_637 (O_637,N_4658,N_4764);
and UO_638 (O_638,N_4829,N_4876);
or UO_639 (O_639,N_4977,N_4594);
or UO_640 (O_640,N_4688,N_4683);
or UO_641 (O_641,N_4591,N_4816);
xor UO_642 (O_642,N_4733,N_4616);
xnor UO_643 (O_643,N_4509,N_4536);
nand UO_644 (O_644,N_4998,N_4588);
nand UO_645 (O_645,N_4864,N_4882);
nor UO_646 (O_646,N_4641,N_4632);
or UO_647 (O_647,N_4833,N_4923);
xnor UO_648 (O_648,N_4613,N_4851);
nor UO_649 (O_649,N_4835,N_4738);
nor UO_650 (O_650,N_4860,N_4651);
nand UO_651 (O_651,N_4520,N_4949);
and UO_652 (O_652,N_4849,N_4730);
or UO_653 (O_653,N_4853,N_4779);
or UO_654 (O_654,N_4545,N_4621);
and UO_655 (O_655,N_4924,N_4798);
or UO_656 (O_656,N_4500,N_4845);
or UO_657 (O_657,N_4741,N_4949);
and UO_658 (O_658,N_4820,N_4619);
nand UO_659 (O_659,N_4642,N_4679);
nor UO_660 (O_660,N_4611,N_4658);
nor UO_661 (O_661,N_4618,N_4760);
nand UO_662 (O_662,N_4820,N_4726);
xnor UO_663 (O_663,N_4743,N_4684);
or UO_664 (O_664,N_4861,N_4613);
nand UO_665 (O_665,N_4721,N_4906);
or UO_666 (O_666,N_4944,N_4943);
and UO_667 (O_667,N_4830,N_4620);
or UO_668 (O_668,N_4636,N_4546);
or UO_669 (O_669,N_4762,N_4646);
and UO_670 (O_670,N_4767,N_4656);
or UO_671 (O_671,N_4943,N_4761);
xor UO_672 (O_672,N_4787,N_4673);
nand UO_673 (O_673,N_4559,N_4900);
nor UO_674 (O_674,N_4526,N_4862);
or UO_675 (O_675,N_4620,N_4984);
nand UO_676 (O_676,N_4582,N_4654);
nor UO_677 (O_677,N_4681,N_4532);
nand UO_678 (O_678,N_4797,N_4979);
or UO_679 (O_679,N_4681,N_4939);
xor UO_680 (O_680,N_4891,N_4655);
xnor UO_681 (O_681,N_4565,N_4626);
xor UO_682 (O_682,N_4543,N_4781);
and UO_683 (O_683,N_4944,N_4977);
nand UO_684 (O_684,N_4705,N_4533);
nand UO_685 (O_685,N_4685,N_4593);
or UO_686 (O_686,N_4947,N_4931);
or UO_687 (O_687,N_4574,N_4699);
and UO_688 (O_688,N_4507,N_4527);
or UO_689 (O_689,N_4711,N_4894);
nor UO_690 (O_690,N_4663,N_4599);
or UO_691 (O_691,N_4705,N_4601);
nor UO_692 (O_692,N_4736,N_4931);
xor UO_693 (O_693,N_4755,N_4775);
xnor UO_694 (O_694,N_4815,N_4966);
and UO_695 (O_695,N_4609,N_4755);
nor UO_696 (O_696,N_4789,N_4544);
xor UO_697 (O_697,N_4965,N_4822);
nand UO_698 (O_698,N_4586,N_4989);
and UO_699 (O_699,N_4512,N_4551);
and UO_700 (O_700,N_4576,N_4920);
nand UO_701 (O_701,N_4908,N_4552);
nand UO_702 (O_702,N_4894,N_4684);
nor UO_703 (O_703,N_4759,N_4889);
nor UO_704 (O_704,N_4902,N_4988);
nor UO_705 (O_705,N_4885,N_4637);
and UO_706 (O_706,N_4679,N_4740);
nand UO_707 (O_707,N_4925,N_4649);
nand UO_708 (O_708,N_4657,N_4551);
or UO_709 (O_709,N_4941,N_4962);
xor UO_710 (O_710,N_4797,N_4772);
xor UO_711 (O_711,N_4686,N_4554);
or UO_712 (O_712,N_4790,N_4829);
and UO_713 (O_713,N_4644,N_4700);
nand UO_714 (O_714,N_4546,N_4959);
or UO_715 (O_715,N_4824,N_4511);
and UO_716 (O_716,N_4970,N_4888);
nand UO_717 (O_717,N_4989,N_4931);
and UO_718 (O_718,N_4977,N_4976);
nor UO_719 (O_719,N_4750,N_4803);
or UO_720 (O_720,N_4757,N_4731);
nand UO_721 (O_721,N_4698,N_4721);
nor UO_722 (O_722,N_4976,N_4718);
nor UO_723 (O_723,N_4716,N_4547);
or UO_724 (O_724,N_4781,N_4817);
or UO_725 (O_725,N_4736,N_4811);
xor UO_726 (O_726,N_4760,N_4679);
nand UO_727 (O_727,N_4996,N_4554);
xor UO_728 (O_728,N_4816,N_4919);
xor UO_729 (O_729,N_4814,N_4699);
xor UO_730 (O_730,N_4637,N_4632);
xnor UO_731 (O_731,N_4891,N_4689);
nand UO_732 (O_732,N_4919,N_4920);
and UO_733 (O_733,N_4952,N_4720);
and UO_734 (O_734,N_4985,N_4978);
nand UO_735 (O_735,N_4923,N_4777);
or UO_736 (O_736,N_4648,N_4722);
nor UO_737 (O_737,N_4559,N_4505);
xnor UO_738 (O_738,N_4662,N_4888);
and UO_739 (O_739,N_4538,N_4615);
and UO_740 (O_740,N_4904,N_4581);
xor UO_741 (O_741,N_4776,N_4744);
nor UO_742 (O_742,N_4969,N_4527);
nor UO_743 (O_743,N_4920,N_4854);
or UO_744 (O_744,N_4739,N_4637);
or UO_745 (O_745,N_4602,N_4736);
xor UO_746 (O_746,N_4649,N_4623);
and UO_747 (O_747,N_4685,N_4546);
or UO_748 (O_748,N_4702,N_4614);
xnor UO_749 (O_749,N_4528,N_4514);
or UO_750 (O_750,N_4954,N_4893);
xor UO_751 (O_751,N_4921,N_4501);
nor UO_752 (O_752,N_4535,N_4783);
or UO_753 (O_753,N_4859,N_4812);
and UO_754 (O_754,N_4595,N_4867);
and UO_755 (O_755,N_4539,N_4988);
xor UO_756 (O_756,N_4637,N_4775);
nand UO_757 (O_757,N_4963,N_4959);
nor UO_758 (O_758,N_4922,N_4637);
and UO_759 (O_759,N_4708,N_4820);
and UO_760 (O_760,N_4506,N_4827);
or UO_761 (O_761,N_4582,N_4501);
nor UO_762 (O_762,N_4633,N_4745);
nand UO_763 (O_763,N_4865,N_4614);
xnor UO_764 (O_764,N_4837,N_4801);
or UO_765 (O_765,N_4537,N_4910);
and UO_766 (O_766,N_4883,N_4776);
xnor UO_767 (O_767,N_4611,N_4612);
and UO_768 (O_768,N_4541,N_4612);
and UO_769 (O_769,N_4504,N_4831);
xor UO_770 (O_770,N_4638,N_4966);
xor UO_771 (O_771,N_4689,N_4980);
xor UO_772 (O_772,N_4616,N_4944);
or UO_773 (O_773,N_4936,N_4682);
xor UO_774 (O_774,N_4729,N_4705);
xnor UO_775 (O_775,N_4668,N_4785);
or UO_776 (O_776,N_4768,N_4593);
nor UO_777 (O_777,N_4971,N_4845);
xor UO_778 (O_778,N_4598,N_4802);
nor UO_779 (O_779,N_4516,N_4607);
and UO_780 (O_780,N_4986,N_4629);
nor UO_781 (O_781,N_4577,N_4851);
nor UO_782 (O_782,N_4694,N_4575);
nor UO_783 (O_783,N_4992,N_4912);
nor UO_784 (O_784,N_4505,N_4583);
xnor UO_785 (O_785,N_4807,N_4979);
nor UO_786 (O_786,N_4627,N_4703);
nor UO_787 (O_787,N_4667,N_4581);
xnor UO_788 (O_788,N_4752,N_4722);
nor UO_789 (O_789,N_4695,N_4613);
nand UO_790 (O_790,N_4996,N_4824);
or UO_791 (O_791,N_4737,N_4730);
nand UO_792 (O_792,N_4806,N_4514);
nand UO_793 (O_793,N_4654,N_4679);
and UO_794 (O_794,N_4762,N_4760);
nand UO_795 (O_795,N_4976,N_4958);
or UO_796 (O_796,N_4762,N_4990);
nand UO_797 (O_797,N_4953,N_4640);
or UO_798 (O_798,N_4715,N_4519);
nand UO_799 (O_799,N_4566,N_4767);
and UO_800 (O_800,N_4584,N_4509);
xor UO_801 (O_801,N_4891,N_4676);
nor UO_802 (O_802,N_4730,N_4562);
and UO_803 (O_803,N_4818,N_4593);
xnor UO_804 (O_804,N_4986,N_4816);
or UO_805 (O_805,N_4674,N_4539);
nand UO_806 (O_806,N_4572,N_4688);
xnor UO_807 (O_807,N_4673,N_4565);
and UO_808 (O_808,N_4533,N_4654);
and UO_809 (O_809,N_4875,N_4805);
or UO_810 (O_810,N_4697,N_4970);
or UO_811 (O_811,N_4952,N_4589);
nor UO_812 (O_812,N_4585,N_4508);
nor UO_813 (O_813,N_4629,N_4989);
or UO_814 (O_814,N_4769,N_4938);
nor UO_815 (O_815,N_4894,N_4928);
xor UO_816 (O_816,N_4930,N_4793);
nor UO_817 (O_817,N_4618,N_4854);
nor UO_818 (O_818,N_4760,N_4932);
xor UO_819 (O_819,N_4852,N_4638);
or UO_820 (O_820,N_4777,N_4747);
nand UO_821 (O_821,N_4578,N_4632);
nor UO_822 (O_822,N_4842,N_4857);
or UO_823 (O_823,N_4701,N_4575);
and UO_824 (O_824,N_4650,N_4783);
xnor UO_825 (O_825,N_4616,N_4568);
or UO_826 (O_826,N_4860,N_4901);
or UO_827 (O_827,N_4639,N_4781);
and UO_828 (O_828,N_4765,N_4975);
or UO_829 (O_829,N_4522,N_4742);
or UO_830 (O_830,N_4597,N_4644);
nor UO_831 (O_831,N_4541,N_4503);
nand UO_832 (O_832,N_4533,N_4871);
nor UO_833 (O_833,N_4994,N_4968);
nor UO_834 (O_834,N_4888,N_4735);
nor UO_835 (O_835,N_4640,N_4974);
or UO_836 (O_836,N_4510,N_4558);
or UO_837 (O_837,N_4944,N_4976);
and UO_838 (O_838,N_4595,N_4713);
xor UO_839 (O_839,N_4885,N_4573);
xor UO_840 (O_840,N_4885,N_4944);
and UO_841 (O_841,N_4791,N_4634);
or UO_842 (O_842,N_4729,N_4760);
and UO_843 (O_843,N_4573,N_4681);
or UO_844 (O_844,N_4882,N_4529);
nand UO_845 (O_845,N_4978,N_4708);
or UO_846 (O_846,N_4880,N_4734);
and UO_847 (O_847,N_4858,N_4541);
or UO_848 (O_848,N_4564,N_4854);
xor UO_849 (O_849,N_4787,N_4814);
or UO_850 (O_850,N_4947,N_4801);
xor UO_851 (O_851,N_4792,N_4718);
nor UO_852 (O_852,N_4893,N_4741);
nand UO_853 (O_853,N_4916,N_4864);
nand UO_854 (O_854,N_4724,N_4803);
and UO_855 (O_855,N_4603,N_4594);
or UO_856 (O_856,N_4901,N_4718);
xnor UO_857 (O_857,N_4539,N_4957);
nand UO_858 (O_858,N_4847,N_4779);
and UO_859 (O_859,N_4641,N_4983);
nor UO_860 (O_860,N_4957,N_4660);
or UO_861 (O_861,N_4864,N_4813);
and UO_862 (O_862,N_4591,N_4602);
nand UO_863 (O_863,N_4945,N_4661);
xor UO_864 (O_864,N_4680,N_4855);
and UO_865 (O_865,N_4554,N_4610);
and UO_866 (O_866,N_4664,N_4628);
nand UO_867 (O_867,N_4610,N_4885);
and UO_868 (O_868,N_4967,N_4969);
nor UO_869 (O_869,N_4699,N_4880);
or UO_870 (O_870,N_4730,N_4621);
nand UO_871 (O_871,N_4560,N_4866);
xor UO_872 (O_872,N_4974,N_4716);
nand UO_873 (O_873,N_4595,N_4968);
nand UO_874 (O_874,N_4792,N_4943);
or UO_875 (O_875,N_4855,N_4856);
nor UO_876 (O_876,N_4544,N_4615);
or UO_877 (O_877,N_4720,N_4913);
nand UO_878 (O_878,N_4672,N_4604);
nand UO_879 (O_879,N_4549,N_4997);
or UO_880 (O_880,N_4959,N_4531);
or UO_881 (O_881,N_4590,N_4628);
or UO_882 (O_882,N_4570,N_4678);
xnor UO_883 (O_883,N_4933,N_4791);
nor UO_884 (O_884,N_4524,N_4765);
and UO_885 (O_885,N_4512,N_4727);
xor UO_886 (O_886,N_4751,N_4728);
nor UO_887 (O_887,N_4860,N_4844);
nand UO_888 (O_888,N_4959,N_4502);
or UO_889 (O_889,N_4845,N_4659);
and UO_890 (O_890,N_4505,N_4996);
and UO_891 (O_891,N_4605,N_4505);
nor UO_892 (O_892,N_4979,N_4684);
or UO_893 (O_893,N_4763,N_4573);
nor UO_894 (O_894,N_4867,N_4936);
and UO_895 (O_895,N_4890,N_4737);
and UO_896 (O_896,N_4870,N_4743);
xor UO_897 (O_897,N_4734,N_4688);
xnor UO_898 (O_898,N_4612,N_4870);
nor UO_899 (O_899,N_4889,N_4772);
nand UO_900 (O_900,N_4705,N_4580);
nor UO_901 (O_901,N_4688,N_4863);
and UO_902 (O_902,N_4708,N_4788);
xnor UO_903 (O_903,N_4567,N_4537);
nor UO_904 (O_904,N_4680,N_4895);
nand UO_905 (O_905,N_4952,N_4555);
xor UO_906 (O_906,N_4600,N_4572);
or UO_907 (O_907,N_4784,N_4556);
and UO_908 (O_908,N_4537,N_4994);
nor UO_909 (O_909,N_4919,N_4827);
xnor UO_910 (O_910,N_4933,N_4774);
or UO_911 (O_911,N_4758,N_4904);
and UO_912 (O_912,N_4523,N_4540);
or UO_913 (O_913,N_4674,N_4568);
nor UO_914 (O_914,N_4968,N_4966);
and UO_915 (O_915,N_4731,N_4514);
nand UO_916 (O_916,N_4704,N_4647);
and UO_917 (O_917,N_4926,N_4996);
xor UO_918 (O_918,N_4564,N_4530);
and UO_919 (O_919,N_4608,N_4969);
and UO_920 (O_920,N_4634,N_4544);
and UO_921 (O_921,N_4549,N_4771);
xor UO_922 (O_922,N_4974,N_4687);
nand UO_923 (O_923,N_4581,N_4538);
nor UO_924 (O_924,N_4583,N_4924);
nor UO_925 (O_925,N_4968,N_4683);
nand UO_926 (O_926,N_4736,N_4621);
nand UO_927 (O_927,N_4673,N_4627);
and UO_928 (O_928,N_4862,N_4545);
nand UO_929 (O_929,N_4963,N_4512);
or UO_930 (O_930,N_4600,N_4849);
xor UO_931 (O_931,N_4913,N_4766);
or UO_932 (O_932,N_4877,N_4802);
and UO_933 (O_933,N_4958,N_4662);
nand UO_934 (O_934,N_4927,N_4844);
or UO_935 (O_935,N_4552,N_4627);
and UO_936 (O_936,N_4949,N_4681);
nand UO_937 (O_937,N_4569,N_4770);
or UO_938 (O_938,N_4850,N_4845);
or UO_939 (O_939,N_4759,N_4595);
xnor UO_940 (O_940,N_4507,N_4656);
nor UO_941 (O_941,N_4674,N_4604);
and UO_942 (O_942,N_4984,N_4589);
or UO_943 (O_943,N_4827,N_4520);
nor UO_944 (O_944,N_4939,N_4680);
or UO_945 (O_945,N_4773,N_4868);
nor UO_946 (O_946,N_4974,N_4924);
and UO_947 (O_947,N_4773,N_4756);
and UO_948 (O_948,N_4837,N_4636);
nand UO_949 (O_949,N_4950,N_4743);
or UO_950 (O_950,N_4919,N_4502);
xnor UO_951 (O_951,N_4959,N_4921);
nand UO_952 (O_952,N_4862,N_4993);
or UO_953 (O_953,N_4554,N_4989);
xor UO_954 (O_954,N_4525,N_4976);
xor UO_955 (O_955,N_4898,N_4590);
and UO_956 (O_956,N_4794,N_4760);
or UO_957 (O_957,N_4703,N_4612);
nor UO_958 (O_958,N_4745,N_4792);
xnor UO_959 (O_959,N_4764,N_4755);
or UO_960 (O_960,N_4502,N_4820);
or UO_961 (O_961,N_4788,N_4740);
nor UO_962 (O_962,N_4592,N_4542);
or UO_963 (O_963,N_4893,N_4982);
and UO_964 (O_964,N_4882,N_4824);
or UO_965 (O_965,N_4958,N_4767);
and UO_966 (O_966,N_4693,N_4636);
xnor UO_967 (O_967,N_4586,N_4804);
nand UO_968 (O_968,N_4946,N_4849);
xnor UO_969 (O_969,N_4669,N_4978);
nand UO_970 (O_970,N_4638,N_4863);
or UO_971 (O_971,N_4730,N_4968);
nand UO_972 (O_972,N_4560,N_4913);
nor UO_973 (O_973,N_4552,N_4860);
or UO_974 (O_974,N_4973,N_4955);
nand UO_975 (O_975,N_4898,N_4643);
nor UO_976 (O_976,N_4657,N_4845);
and UO_977 (O_977,N_4814,N_4668);
xor UO_978 (O_978,N_4520,N_4920);
xnor UO_979 (O_979,N_4813,N_4997);
or UO_980 (O_980,N_4850,N_4835);
nor UO_981 (O_981,N_4964,N_4997);
nor UO_982 (O_982,N_4671,N_4906);
xnor UO_983 (O_983,N_4579,N_4602);
and UO_984 (O_984,N_4564,N_4904);
xor UO_985 (O_985,N_4710,N_4842);
nor UO_986 (O_986,N_4803,N_4538);
nor UO_987 (O_987,N_4594,N_4886);
nor UO_988 (O_988,N_4795,N_4720);
and UO_989 (O_989,N_4644,N_4577);
nor UO_990 (O_990,N_4975,N_4685);
or UO_991 (O_991,N_4918,N_4529);
and UO_992 (O_992,N_4875,N_4641);
xor UO_993 (O_993,N_4844,N_4841);
nand UO_994 (O_994,N_4562,N_4704);
xnor UO_995 (O_995,N_4900,N_4778);
xnor UO_996 (O_996,N_4715,N_4911);
nand UO_997 (O_997,N_4800,N_4735);
and UO_998 (O_998,N_4585,N_4824);
nand UO_999 (O_999,N_4696,N_4748);
endmodule