module basic_1500_15000_2000_5_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_2,In_578);
nor U1 (N_1,In_138,In_1168);
nand U2 (N_2,In_608,In_565);
xor U3 (N_3,In_468,In_676);
nand U4 (N_4,In_948,In_639);
and U5 (N_5,In_78,In_940);
nand U6 (N_6,In_1152,In_444);
and U7 (N_7,In_835,In_1205);
nor U8 (N_8,In_386,In_654);
nor U9 (N_9,In_1295,In_1473);
or U10 (N_10,In_606,In_217);
xnor U11 (N_11,In_106,In_1171);
nor U12 (N_12,In_904,In_919);
nor U13 (N_13,In_66,In_631);
or U14 (N_14,In_636,In_1145);
and U15 (N_15,In_1148,In_462);
nand U16 (N_16,In_1355,In_1489);
and U17 (N_17,In_330,In_46);
or U18 (N_18,In_775,In_1404);
nand U19 (N_19,In_338,In_414);
or U20 (N_20,In_29,In_1276);
or U21 (N_21,In_875,In_365);
and U22 (N_22,In_1493,In_307);
xnor U23 (N_23,In_1432,In_1435);
or U24 (N_24,In_889,In_43);
xor U25 (N_25,In_558,In_1345);
nand U26 (N_26,In_1407,In_1296);
nand U27 (N_27,In_864,In_596);
or U28 (N_28,In_852,In_1056);
xnor U29 (N_29,In_980,In_734);
xnor U30 (N_30,In_1100,In_1040);
or U31 (N_31,In_149,In_272);
nor U32 (N_32,In_1313,In_1170);
xor U33 (N_33,In_866,In_94);
and U34 (N_34,In_222,In_771);
or U35 (N_35,In_197,In_661);
nand U36 (N_36,In_928,In_705);
nor U37 (N_37,In_576,In_1298);
and U38 (N_38,In_354,In_991);
nand U39 (N_39,In_477,In_1156);
and U40 (N_40,In_367,In_214);
nor U41 (N_41,In_355,In_32);
xor U42 (N_42,In_581,In_933);
or U43 (N_43,In_1034,In_746);
or U44 (N_44,In_525,In_1323);
nor U45 (N_45,In_960,In_4);
xor U46 (N_46,In_783,In_1078);
nor U47 (N_47,In_1098,In_759);
or U48 (N_48,In_303,In_333);
nor U49 (N_49,In_597,In_379);
and U50 (N_50,In_1483,In_751);
nand U51 (N_51,In_387,In_1251);
and U52 (N_52,In_1144,In_1285);
and U53 (N_53,In_473,In_259);
nor U54 (N_54,In_21,In_766);
nand U55 (N_55,In_1282,In_594);
nand U56 (N_56,In_560,In_1248);
xor U57 (N_57,In_40,In_997);
xor U58 (N_58,In_300,In_610);
and U59 (N_59,In_1362,In_84);
and U60 (N_60,In_1016,In_288);
and U61 (N_61,In_53,In_1172);
and U62 (N_62,In_906,In_1229);
and U63 (N_63,In_1390,In_1136);
xnor U64 (N_64,In_344,In_1310);
or U65 (N_65,In_1181,In_100);
or U66 (N_66,In_360,In_669);
xor U67 (N_67,In_87,In_1055);
nand U68 (N_68,In_789,In_1252);
nand U69 (N_69,In_522,In_281);
nor U70 (N_70,In_1437,In_1017);
nor U71 (N_71,In_1253,In_570);
nor U72 (N_72,In_494,In_488);
nand U73 (N_73,In_580,In_103);
nand U74 (N_74,In_125,In_1422);
nand U75 (N_75,In_611,In_1333);
xor U76 (N_76,In_811,In_953);
nand U77 (N_77,In_112,In_1399);
nand U78 (N_78,In_196,In_1480);
or U79 (N_79,In_484,In_198);
or U80 (N_80,In_859,In_151);
and U81 (N_81,In_132,In_752);
nand U82 (N_82,In_1084,In_1228);
and U83 (N_83,In_286,In_858);
nor U84 (N_84,In_1411,In_440);
and U85 (N_85,In_1268,In_265);
xnor U86 (N_86,In_25,In_184);
and U87 (N_87,In_1211,In_48);
and U88 (N_88,In_486,In_408);
nor U89 (N_89,In_709,In_1442);
and U90 (N_90,In_302,In_323);
xnor U91 (N_91,In_943,In_230);
and U92 (N_92,In_1461,In_1431);
nor U93 (N_93,In_507,In_485);
xor U94 (N_94,In_1197,In_258);
or U95 (N_95,In_1330,In_397);
and U96 (N_96,In_1352,In_917);
and U97 (N_97,In_1135,In_317);
or U98 (N_98,In_1206,In_117);
or U99 (N_99,In_218,In_795);
nor U100 (N_100,In_1004,In_1191);
and U101 (N_101,In_869,In_718);
nor U102 (N_102,In_975,In_118);
nand U103 (N_103,In_1482,In_264);
nand U104 (N_104,In_533,In_749);
nor U105 (N_105,In_1005,In_1497);
nor U106 (N_106,In_395,In_1311);
and U107 (N_107,In_1416,In_1054);
xnor U108 (N_108,In_526,In_1196);
nor U109 (N_109,In_1117,In_1121);
or U110 (N_110,In_707,In_1202);
nor U111 (N_111,In_1446,In_175);
or U112 (N_112,In_1209,In_347);
nor U113 (N_113,In_976,In_1366);
xnor U114 (N_114,In_509,In_398);
nor U115 (N_115,In_75,In_407);
xnor U116 (N_116,In_822,In_1015);
nor U117 (N_117,In_781,In_1081);
and U118 (N_118,In_529,In_260);
xnor U119 (N_119,In_320,In_511);
or U120 (N_120,In_966,In_1060);
nand U121 (N_121,In_825,In_729);
and U122 (N_122,In_814,In_492);
xnor U123 (N_123,In_1163,In_1498);
or U124 (N_124,In_1427,In_1154);
xnor U125 (N_125,In_1027,In_158);
nand U126 (N_126,In_713,In_1426);
nor U127 (N_127,In_539,In_193);
xnor U128 (N_128,In_712,In_296);
nand U129 (N_129,In_1018,In_714);
nor U130 (N_130,In_692,In_855);
and U131 (N_131,In_1468,In_1104);
and U132 (N_132,In_240,In_542);
xnor U133 (N_133,In_772,In_741);
xnor U134 (N_134,In_1457,In_1421);
nand U135 (N_135,In_737,In_8);
nor U136 (N_136,In_223,In_1300);
xnor U137 (N_137,In_845,In_1361);
xnor U138 (N_138,In_309,In_215);
or U139 (N_139,In_950,In_651);
xor U140 (N_140,In_1043,In_412);
or U141 (N_141,In_974,In_1299);
and U142 (N_142,In_1124,In_804);
and U143 (N_143,In_892,In_1091);
xnor U144 (N_144,In_527,In_37);
nand U145 (N_145,In_466,In_1237);
nor U146 (N_146,In_96,In_97);
and U147 (N_147,In_1382,In_753);
or U148 (N_148,In_1340,In_1212);
xnor U149 (N_149,In_1149,In_1302);
and U150 (N_150,In_888,In_1408);
nand U151 (N_151,In_496,In_1449);
nand U152 (N_152,In_1413,In_902);
and U153 (N_153,In_1035,In_328);
and U154 (N_154,In_1110,In_874);
nand U155 (N_155,In_1372,In_936);
or U156 (N_156,In_1021,In_767);
nor U157 (N_157,In_871,In_963);
xor U158 (N_158,In_30,In_680);
or U159 (N_159,In_798,In_124);
or U160 (N_160,In_730,In_1398);
nor U161 (N_161,In_1046,In_1453);
xor U162 (N_162,In_946,In_1256);
xor U163 (N_163,In_955,In_183);
nor U164 (N_164,In_350,In_695);
or U165 (N_165,In_1115,In_1195);
nor U166 (N_166,In_546,In_1138);
and U167 (N_167,In_479,In_1082);
nor U168 (N_168,In_778,In_489);
and U169 (N_169,In_1109,In_797);
and U170 (N_170,In_926,In_16);
and U171 (N_171,In_1491,In_1391);
nor U172 (N_172,In_615,In_277);
nor U173 (N_173,In_1113,In_1069);
xnor U174 (N_174,In_985,In_340);
xor U175 (N_175,In_1020,In_732);
or U176 (N_176,In_1047,In_817);
nand U177 (N_177,In_949,In_846);
or U178 (N_178,In_1241,In_342);
or U179 (N_179,In_847,In_979);
or U180 (N_180,In_856,In_824);
or U181 (N_181,In_982,In_881);
xnor U182 (N_182,In_135,In_474);
nand U183 (N_183,In_688,In_31);
or U184 (N_184,In_1289,In_1418);
xnor U185 (N_185,In_1327,In_22);
or U186 (N_186,In_449,In_1267);
nor U187 (N_187,In_475,In_898);
nand U188 (N_188,In_1188,In_363);
and U189 (N_189,In_878,In_1474);
or U190 (N_190,In_941,In_405);
or U191 (N_191,In_312,In_987);
nor U192 (N_192,In_1410,In_1224);
xnor U193 (N_193,In_1158,In_1093);
and U194 (N_194,In_246,In_267);
nand U195 (N_195,In_332,In_870);
or U196 (N_196,In_208,In_1266);
xor U197 (N_197,In_551,In_787);
nor U198 (N_198,In_971,In_426);
nand U199 (N_199,In_1214,In_655);
or U200 (N_200,In_957,In_1179);
xor U201 (N_201,In_69,In_704);
and U202 (N_202,In_389,In_109);
xor U203 (N_203,In_1147,In_561);
nor U204 (N_204,In_1487,In_261);
or U205 (N_205,In_463,In_1232);
xor U206 (N_206,In_1173,In_952);
xor U207 (N_207,In_429,In_577);
nor U208 (N_208,In_616,In_1233);
nor U209 (N_209,In_498,In_101);
nor U210 (N_210,In_665,In_161);
nor U211 (N_211,In_1436,In_1165);
nor U212 (N_212,In_880,In_873);
and U213 (N_213,In_262,In_506);
or U214 (N_214,In_867,In_0);
and U215 (N_215,In_1192,In_245);
and U216 (N_216,In_1119,In_588);
and U217 (N_217,In_56,In_863);
nand U218 (N_218,In_996,In_836);
and U219 (N_219,In_10,In_126);
or U220 (N_220,In_1343,In_644);
or U221 (N_221,In_165,In_838);
xnor U222 (N_222,In_186,In_357);
and U223 (N_223,In_1288,In_480);
nand U224 (N_224,In_1150,In_211);
or U225 (N_225,In_252,In_1353);
nand U226 (N_226,In_939,In_119);
nand U227 (N_227,In_791,In_1259);
and U228 (N_228,In_907,In_394);
xor U229 (N_229,In_818,In_18);
nand U230 (N_230,In_1290,In_1484);
nor U231 (N_231,In_1274,In_290);
and U232 (N_232,In_279,In_1472);
nor U233 (N_233,In_965,In_571);
nand U234 (N_234,In_1358,In_538);
nand U235 (N_235,In_1219,In_1384);
nor U236 (N_236,In_319,In_1048);
and U237 (N_237,In_83,In_219);
nand U238 (N_238,In_550,In_1280);
or U239 (N_239,In_160,In_735);
xor U240 (N_240,In_573,In_331);
nand U241 (N_241,In_912,In_1388);
nand U242 (N_242,In_1316,In_521);
nand U243 (N_243,In_1127,In_1161);
nor U244 (N_244,In_1373,In_1456);
or U245 (N_245,In_157,In_678);
nand U246 (N_246,In_154,In_456);
nor U247 (N_247,In_715,In_1466);
nor U248 (N_248,In_1080,In_883);
or U249 (N_249,In_1059,In_670);
and U250 (N_250,In_679,In_1185);
nor U251 (N_251,In_1486,In_559);
or U252 (N_252,In_796,In_553);
nor U253 (N_253,In_301,In_583);
or U254 (N_254,In_1090,In_1215);
or U255 (N_255,In_513,In_793);
or U256 (N_256,In_1007,In_537);
or U257 (N_257,In_1079,In_1178);
nor U258 (N_258,In_684,In_164);
nor U259 (N_259,In_890,In_674);
nor U260 (N_260,In_1201,In_346);
and U261 (N_261,In_809,In_1275);
and U262 (N_262,In_1063,In_435);
nand U263 (N_263,In_388,In_104);
nor U264 (N_264,In_35,In_1338);
nor U265 (N_265,In_244,In_1216);
nand U266 (N_266,In_800,In_711);
or U267 (N_267,In_1102,In_133);
nand U268 (N_268,In_231,In_931);
nor U269 (N_269,In_1208,In_652);
and U270 (N_270,In_374,In_147);
and U271 (N_271,In_587,In_39);
xnor U272 (N_272,In_994,In_853);
or U273 (N_273,In_815,In_503);
nand U274 (N_274,In_664,In_105);
or U275 (N_275,In_1106,In_122);
and U276 (N_276,In_1430,In_465);
nand U277 (N_277,In_1057,In_1469);
and U278 (N_278,In_1227,In_224);
xor U279 (N_279,In_427,In_812);
nand U280 (N_280,In_251,In_790);
nor U281 (N_281,In_321,In_885);
and U282 (N_282,In_417,In_55);
or U283 (N_283,In_436,In_1022);
nand U284 (N_284,In_114,In_1058);
xor U285 (N_285,In_326,In_68);
nand U286 (N_286,In_450,In_1061);
nor U287 (N_287,In_168,In_820);
or U288 (N_288,In_51,In_378);
nor U289 (N_289,In_210,In_134);
nand U290 (N_290,In_70,In_1346);
nor U291 (N_291,In_1264,In_834);
and U292 (N_292,In_1255,In_514);
nor U293 (N_293,In_765,In_599);
and U294 (N_294,In_603,In_842);
and U295 (N_295,In_34,In_366);
nor U296 (N_296,In_1062,In_337);
xnor U297 (N_297,In_416,In_313);
nand U298 (N_298,In_530,In_327);
xnor U299 (N_299,In_731,In_1207);
and U300 (N_300,In_769,In_140);
and U301 (N_301,In_297,In_1231);
nand U302 (N_302,In_194,In_1269);
nor U303 (N_303,In_1347,In_88);
xnor U304 (N_304,In_99,In_38);
xor U305 (N_305,In_59,In_128);
nor U306 (N_306,In_1155,In_643);
nor U307 (N_307,In_1271,In_1068);
nor U308 (N_308,In_137,In_547);
xnor U309 (N_309,In_1095,In_1126);
xor U310 (N_310,In_534,In_719);
or U311 (N_311,In_810,In_1001);
xnor U312 (N_312,In_903,In_49);
and U313 (N_313,In_255,In_1130);
xor U314 (N_314,In_9,In_1071);
or U315 (N_315,In_36,In_887);
xnor U316 (N_316,In_432,In_1332);
or U317 (N_317,In_467,In_123);
and U318 (N_318,In_1365,In_598);
or U319 (N_319,In_1439,In_799);
or U320 (N_320,In_1423,In_1257);
or U321 (N_321,In_660,In_555);
nor U322 (N_322,In_595,In_776);
and U323 (N_323,In_945,In_418);
nand U324 (N_324,In_528,In_411);
nor U325 (N_325,In_854,In_628);
xor U326 (N_326,In_287,In_794);
nor U327 (N_327,In_62,In_829);
and U328 (N_328,In_404,In_1342);
or U329 (N_329,In_633,In_1448);
nor U330 (N_330,In_1225,In_1222);
xnor U331 (N_331,In_738,In_552);
nand U332 (N_332,In_609,In_1344);
xor U333 (N_333,In_173,In_1318);
nand U334 (N_334,In_1326,In_657);
or U335 (N_335,In_1336,In_893);
nor U336 (N_336,In_413,In_1242);
or U337 (N_337,In_921,In_720);
nor U338 (N_338,In_536,In_848);
or U339 (N_339,In_461,In_1164);
or U340 (N_340,In_207,In_110);
nand U341 (N_341,In_1011,In_942);
or U342 (N_342,In_1258,In_1462);
nor U343 (N_343,In_273,In_401);
and U344 (N_344,In_1492,In_944);
nor U345 (N_345,In_382,In_620);
and U346 (N_346,In_141,In_189);
nand U347 (N_347,In_1369,In_64);
and U348 (N_348,In_677,In_770);
nor U349 (N_349,In_129,In_1169);
xor U350 (N_350,In_263,In_314);
nand U351 (N_351,In_882,In_823);
nor U352 (N_352,In_969,In_1217);
or U353 (N_353,In_433,In_425);
nor U354 (N_354,In_910,In_675);
nor U355 (N_355,In_981,In_1193);
nor U356 (N_356,In_7,In_637);
nor U357 (N_357,In_174,In_470);
nor U358 (N_358,In_243,In_142);
nor U359 (N_359,In_93,In_879);
xor U360 (N_360,In_1240,In_843);
nor U361 (N_361,In_1309,In_1329);
nor U362 (N_362,In_659,In_322);
nor U363 (N_363,In_517,In_779);
or U364 (N_364,In_499,In_185);
nor U365 (N_365,In_403,In_191);
nor U366 (N_366,In_1262,In_1401);
nand U367 (N_367,In_136,In_1180);
or U368 (N_368,In_410,In_358);
and U369 (N_369,In_1244,In_82);
nand U370 (N_370,In_6,In_85);
and U371 (N_371,In_1230,In_1103);
and U372 (N_372,In_768,In_148);
nor U373 (N_373,In_1182,In_756);
nand U374 (N_374,In_107,In_1415);
or U375 (N_375,In_562,In_1125);
or U376 (N_376,In_841,In_369);
or U377 (N_377,In_162,In_113);
xor U378 (N_378,In_819,In_1368);
nand U379 (N_379,In_1010,In_832);
and U380 (N_380,In_415,In_1286);
xnor U381 (N_381,In_1003,In_370);
nor U382 (N_382,In_1051,In_256);
and U383 (N_383,In_1375,In_755);
nand U384 (N_384,In_454,In_345);
nand U385 (N_385,In_325,In_89);
nand U386 (N_386,In_877,In_1451);
or U387 (N_387,In_977,In_697);
and U388 (N_388,In_1088,In_1350);
xnor U389 (N_389,In_428,In_763);
xnor U390 (N_390,In_341,In_523);
nor U391 (N_391,In_1014,In_472);
or U392 (N_392,In_500,In_773);
xnor U393 (N_393,In_1162,In_1499);
nor U394 (N_394,In_986,In_339);
and U395 (N_395,In_1123,In_1287);
or U396 (N_396,In_200,In_1026);
xor U397 (N_397,In_1291,In_199);
or U398 (N_398,In_723,In_970);
nand U399 (N_399,In_601,In_181);
nand U400 (N_400,In_1438,In_180);
nand U401 (N_401,In_916,In_364);
nor U402 (N_402,In_1085,In_839);
nor U403 (N_403,In_1464,In_324);
xnor U404 (N_404,In_202,In_1292);
or U405 (N_405,In_23,In_72);
nor U406 (N_406,In_187,In_1378);
or U407 (N_407,In_935,In_225);
xor U408 (N_408,In_111,In_1475);
nand U409 (N_409,In_1305,In_159);
xnor U410 (N_410,In_1194,In_1386);
and U411 (N_411,In_642,In_190);
nor U412 (N_412,In_92,In_437);
or U413 (N_413,In_351,In_516);
and U414 (N_414,In_1111,In_1297);
nand U415 (N_415,In_563,In_441);
nand U416 (N_416,In_693,In_1064);
and U417 (N_417,In_648,In_827);
or U418 (N_418,In_837,In_962);
nand U419 (N_419,In_993,In_1281);
or U420 (N_420,In_1187,In_1455);
or U421 (N_421,In_683,In_658);
or U422 (N_422,In_860,In_213);
nand U423 (N_423,In_483,In_579);
xnor U424 (N_424,In_1496,In_130);
nor U425 (N_425,In_742,In_722);
nor U426 (N_426,In_512,In_686);
nand U427 (N_427,In_98,In_895);
or U428 (N_428,In_146,In_682);
nor U429 (N_429,In_1460,In_1030);
or U430 (N_430,In_932,In_750);
xnor U431 (N_431,In_647,In_589);
nand U432 (N_432,In_491,In_1395);
nor U433 (N_433,In_192,In_285);
xnor U434 (N_434,In_681,In_393);
and U435 (N_435,In_865,In_108);
or U436 (N_436,In_14,In_761);
or U437 (N_437,In_163,In_1249);
nand U438 (N_438,In_257,In_721);
or U439 (N_439,In_634,In_1284);
xor U440 (N_440,In_925,In_1307);
nand U441 (N_441,In_619,In_1105);
nand U442 (N_442,In_1443,In_649);
xor U443 (N_443,In_937,In_45);
nand U444 (N_444,In_283,In_690);
xnor U445 (N_445,In_727,In_617);
nor U446 (N_446,In_725,In_1012);
nor U447 (N_447,In_1273,In_1153);
and U448 (N_448,In_748,In_1002);
xnor U449 (N_449,In_329,In_1320);
xnor U450 (N_450,In_816,In_65);
nand U451 (N_451,In_988,In_1128);
nand U452 (N_452,In_703,In_1471);
or U453 (N_453,In_271,In_464);
or U454 (N_454,In_1174,In_602);
xor U455 (N_455,In_574,In_335);
or U456 (N_456,In_127,In_1367);
and U457 (N_457,In_1374,In_143);
nand U458 (N_458,In_481,In_717);
nand U459 (N_459,In_1260,In_144);
nand U460 (N_460,In_782,In_1220);
or U461 (N_461,In_372,In_152);
or U462 (N_462,In_1243,In_1314);
or U463 (N_463,In_622,In_362);
nor U464 (N_464,In_908,In_11);
xnor U465 (N_465,In_24,In_73);
nand U466 (N_466,In_605,In_1247);
xor U467 (N_467,In_1076,In_457);
and U468 (N_468,In_1,In_614);
or U469 (N_469,In_316,In_278);
nand U470 (N_470,In_909,In_1210);
or U471 (N_471,In_292,In_504);
and U472 (N_472,In_972,In_294);
nand U473 (N_473,In_1234,In_204);
nand U474 (N_474,In_739,In_508);
nor U475 (N_475,In_733,In_195);
and U476 (N_476,In_918,In_638);
xor U477 (N_477,In_663,In_299);
and U478 (N_478,In_702,In_894);
xor U479 (N_479,In_188,In_627);
nor U480 (N_480,In_968,In_241);
nand U481 (N_481,In_1363,In_54);
nand U482 (N_482,In_434,In_1023);
or U483 (N_483,In_505,In_268);
and U484 (N_484,In_490,In_831);
xor U485 (N_485,In_1429,In_145);
or U486 (N_486,In_548,In_50);
and U487 (N_487,In_1476,In_1459);
nor U488 (N_488,In_736,In_1122);
nand U489 (N_489,In_802,In_830);
and U490 (N_490,In_1087,In_182);
and U491 (N_491,In_120,In_1037);
xnor U492 (N_492,In_1477,In_421);
nor U493 (N_493,In_938,In_1166);
xor U494 (N_494,In_672,In_229);
nand U495 (N_495,In_375,In_1412);
xor U496 (N_496,In_400,In_803);
nor U497 (N_497,In_1118,In_221);
nand U498 (N_498,In_169,In_376);
xor U499 (N_499,In_33,In_1131);
or U500 (N_500,In_1470,In_1381);
xor U501 (N_501,In_568,In_81);
and U502 (N_502,In_1112,In_1203);
xnor U503 (N_503,In_1074,In_584);
or U504 (N_504,In_455,In_1132);
xnor U505 (N_505,In_1417,In_612);
nand U506 (N_506,In_927,In_167);
and U507 (N_507,In_899,In_1199);
nor U508 (N_508,In_61,In_1183);
nand U509 (N_509,In_861,In_77);
and U510 (N_510,In_95,In_1392);
and U511 (N_511,In_515,In_1319);
or U512 (N_512,In_1349,In_593);
nor U513 (N_513,In_914,In_80);
nor U514 (N_514,In_390,In_150);
or U515 (N_515,In_886,In_1490);
nor U516 (N_516,In_1387,In_983);
or U517 (N_517,In_624,In_253);
or U518 (N_518,In_1032,In_478);
xor U519 (N_519,In_1325,In_1067);
xor U520 (N_520,In_998,In_250);
xor U521 (N_521,In_352,In_1385);
nor U522 (N_522,In_1006,In_274);
nor U523 (N_523,In_399,In_431);
xor U524 (N_524,In_212,In_383);
xor U525 (N_525,In_1066,In_1354);
xnor U526 (N_526,In_650,In_857);
and U527 (N_527,In_406,In_520);
or U528 (N_528,In_999,In_1039);
or U529 (N_529,In_380,In_850);
and U530 (N_530,In_60,In_1190);
or U531 (N_531,In_1175,In_178);
or U532 (N_532,In_519,In_1419);
and U533 (N_533,In_1425,In_626);
nor U534 (N_534,In_469,In_381);
nor U535 (N_535,In_1176,In_1428);
or U536 (N_536,In_269,In_724);
or U537 (N_537,In_532,In_1031);
nor U538 (N_538,In_1304,In_306);
nand U539 (N_539,In_535,In_685);
xnor U540 (N_540,In_86,In_318);
and U541 (N_541,In_786,In_623);
nor U542 (N_542,In_228,In_572);
nor U543 (N_543,In_1270,In_422);
or U544 (N_544,In_780,In_356);
nand U545 (N_545,In_1379,In_757);
or U546 (N_546,In_1420,In_291);
and U547 (N_547,In_1396,In_662);
xor U548 (N_548,In_924,In_1488);
and U549 (N_549,In_502,In_990);
nor U550 (N_550,In_216,In_420);
or U551 (N_551,In_220,In_1089);
nor U552 (N_552,In_1028,In_923);
xnor U553 (N_553,In_518,In_419);
or U554 (N_554,In_728,In_673);
and U555 (N_555,In_276,In_764);
and U556 (N_556,In_967,In_493);
and U557 (N_557,In_701,In_1479);
nor U558 (N_558,In_1221,In_1450);
or U559 (N_559,In_1177,In_964);
and U560 (N_560,In_308,In_201);
nand U561 (N_561,In_564,In_1463);
and U562 (N_562,In_613,In_1394);
or U563 (N_563,In_1389,In_52);
nor U564 (N_564,In_1445,In_876);
xnor U565 (N_565,In_635,In_833);
or U566 (N_566,In_47,In_554);
nand U567 (N_567,In_1013,In_359);
and U568 (N_568,In_1279,In_1025);
and U569 (N_569,In_760,In_1073);
nor U570 (N_570,In_233,In_1049);
or U571 (N_571,In_868,In_984);
and U572 (N_572,In_1033,In_1376);
or U573 (N_573,In_851,In_1405);
nor U574 (N_574,In_1141,In_423);
xnor U575 (N_575,In_745,In_384);
or U576 (N_576,In_1116,In_743);
or U577 (N_577,In_849,In_740);
or U578 (N_578,In_348,In_28);
nor U579 (N_579,In_600,In_762);
nand U580 (N_580,In_495,In_915);
nand U581 (N_581,In_282,In_920);
and U582 (N_582,In_961,In_1434);
or U583 (N_583,In_249,In_343);
or U584 (N_584,In_1380,In_706);
nor U585 (N_585,In_227,In_630);
nor U586 (N_586,In_947,In_973);
xor U587 (N_587,In_1322,In_153);
nor U588 (N_588,In_911,In_115);
nand U589 (N_589,In_995,In_19);
and U590 (N_590,In_353,In_1303);
and U591 (N_591,In_1397,In_1077);
and U592 (N_592,In_284,In_1009);
nand U593 (N_593,In_604,In_1424);
nand U594 (N_594,In_439,In_1334);
or U595 (N_595,In_1072,In_1465);
xor U596 (N_596,In_821,In_254);
nand U597 (N_597,In_424,In_42);
or U598 (N_598,In_646,In_691);
and U599 (N_599,In_872,In_17);
nand U600 (N_600,In_1097,In_280);
or U601 (N_601,In_929,In_569);
or U602 (N_602,In_1356,In_1050);
or U603 (N_603,In_656,In_1184);
xor U604 (N_604,In_1406,In_44);
xor U605 (N_605,In_402,In_1045);
nor U606 (N_606,In_1485,In_166);
and U607 (N_607,In_1335,In_1359);
xor U608 (N_608,In_956,In_445);
or U609 (N_609,In_726,In_807);
xor U610 (N_610,In_671,In_482);
nor U611 (N_611,In_862,In_90);
nor U612 (N_612,In_57,In_930);
nand U613 (N_613,In_540,In_170);
nor U614 (N_614,In_668,In_1277);
or U615 (N_615,In_801,In_1159);
xor U616 (N_616,In_840,In_758);
xnor U617 (N_617,In_76,In_304);
xor U618 (N_618,In_1083,In_1223);
or U619 (N_619,In_1213,In_896);
nand U620 (N_620,In_1364,In_545);
nand U621 (N_621,In_934,In_1142);
or U622 (N_622,In_270,In_203);
and U623 (N_623,In_1265,In_1370);
and U624 (N_624,In_1317,In_1283);
nor U625 (N_625,In_1478,In_1019);
or U626 (N_626,In_295,In_913);
nor U627 (N_627,In_1278,In_266);
nor U628 (N_628,In_26,In_699);
and U629 (N_629,In_1301,In_618);
xnor U630 (N_630,In_3,In_808);
nand U631 (N_631,In_1198,In_1029);
and U632 (N_632,In_1377,In_1444);
or U633 (N_633,In_1000,In_524);
or U634 (N_634,In_311,In_575);
and U635 (N_635,In_1337,In_884);
nand U636 (N_636,In_978,In_531);
nand U637 (N_637,In_777,In_442);
nand U638 (N_638,In_349,In_12);
nor U639 (N_639,In_235,In_275);
nor U640 (N_640,In_1189,In_1263);
or U641 (N_641,In_1092,In_710);
or U642 (N_642,In_901,In_1167);
or U643 (N_643,In_1331,In_1134);
or U644 (N_644,In_1261,In_1293);
xor U645 (N_645,In_237,In_900);
or U646 (N_646,In_586,In_640);
nand U647 (N_647,In_1024,In_1129);
and U648 (N_648,In_121,In_236);
nand U649 (N_649,In_792,In_1146);
nor U650 (N_650,In_497,In_1440);
or U651 (N_651,In_1139,In_716);
nand U652 (N_652,In_1052,In_334);
and U653 (N_653,In_567,In_1441);
or U654 (N_654,In_373,In_844);
or U655 (N_655,In_641,In_79);
nor U656 (N_656,In_689,In_645);
nand U657 (N_657,In_1218,In_632);
or U658 (N_658,In_1053,In_625);
nor U659 (N_659,In_543,In_566);
and U660 (N_660,In_653,In_13);
or U661 (N_661,In_1204,In_607);
or U662 (N_662,In_234,In_392);
and U663 (N_663,In_1246,In_549);
or U664 (N_664,In_451,In_1494);
nand U665 (N_665,In_409,In_242);
nor U666 (N_666,In_1403,In_1186);
nor U667 (N_667,In_1481,In_557);
nand U668 (N_668,In_590,In_1341);
xnor U669 (N_669,In_754,In_1038);
and U670 (N_670,In_1402,In_1447);
xnor U671 (N_671,In_471,In_1371);
nor U672 (N_672,In_430,In_826);
nor U673 (N_673,In_1433,In_377);
or U674 (N_674,In_700,In_396);
nand U675 (N_675,In_541,In_1454);
nand U676 (N_676,In_922,In_67);
xor U677 (N_677,In_1312,In_591);
or U678 (N_678,In_27,In_1086);
and U679 (N_679,In_1315,In_458);
nor U680 (N_680,In_667,In_368);
nand U681 (N_681,In_71,In_1409);
and U682 (N_682,In_959,In_744);
nor U683 (N_683,In_1042,In_361);
xor U684 (N_684,In_1133,In_205);
or U685 (N_685,In_116,In_1351);
xnor U686 (N_686,In_501,In_5);
nor U687 (N_687,In_1101,In_828);
nor U688 (N_688,In_177,In_747);
nor U689 (N_689,In_629,In_139);
nand U690 (N_690,In_20,In_453);
and U691 (N_691,In_905,In_315);
nor U692 (N_692,In_102,In_74);
and U693 (N_693,In_1065,In_1107);
xnor U694 (N_694,In_1348,In_209);
nand U695 (N_695,In_447,In_951);
xnor U696 (N_696,In_694,In_1400);
or U697 (N_697,In_289,In_806);
nand U698 (N_698,In_1108,In_239);
and U699 (N_699,In_460,In_891);
nand U700 (N_700,In_226,In_1360);
and U701 (N_701,In_1200,In_556);
or U702 (N_702,In_91,In_385);
nand U703 (N_703,In_1070,In_1495);
nand U704 (N_704,In_41,In_1383);
xnor U705 (N_705,In_544,In_582);
or U706 (N_706,In_63,In_989);
nor U707 (N_707,In_1137,In_1321);
xnor U708 (N_708,In_1254,In_1245);
and U709 (N_709,In_897,In_592);
and U710 (N_710,In_156,In_698);
and U711 (N_711,In_155,In_298);
or U712 (N_712,In_785,In_1226);
and U713 (N_713,In_1239,In_1044);
and U714 (N_714,In_788,In_1099);
nand U715 (N_715,In_131,In_958);
xor U716 (N_716,In_438,In_992);
or U717 (N_717,In_448,In_1160);
or U718 (N_718,In_621,In_1339);
and U719 (N_719,In_1041,In_1143);
or U720 (N_720,In_1094,In_1357);
xor U721 (N_721,In_687,In_310);
xor U722 (N_722,In_248,In_510);
and U723 (N_723,In_1308,In_1306);
nor U724 (N_724,In_487,In_171);
xor U725 (N_725,In_206,In_371);
or U726 (N_726,In_452,In_954);
nand U727 (N_727,In_1096,In_443);
nor U728 (N_728,In_247,In_1467);
and U729 (N_729,In_784,In_476);
nor U730 (N_730,In_1324,In_179);
and U731 (N_731,In_391,In_1236);
nand U732 (N_732,In_459,In_1151);
xnor U733 (N_733,In_1272,In_1114);
and U734 (N_734,In_1075,In_813);
nand U735 (N_735,In_176,In_172);
or U736 (N_736,In_232,In_696);
and U737 (N_737,In_293,In_305);
nand U738 (N_738,In_238,In_774);
nand U739 (N_739,In_708,In_1328);
or U740 (N_740,In_585,In_666);
and U741 (N_741,In_1294,In_1393);
xnor U742 (N_742,In_1458,In_1008);
nand U743 (N_743,In_1036,In_1140);
nand U744 (N_744,In_805,In_58);
or U745 (N_745,In_1157,In_1238);
xnor U746 (N_746,In_446,In_1452);
xnor U747 (N_747,In_1235,In_1120);
nand U748 (N_748,In_1414,In_336);
nand U749 (N_749,In_1250,In_15);
nor U750 (N_750,In_393,In_170);
nand U751 (N_751,In_1036,In_556);
and U752 (N_752,In_1218,In_445);
nand U753 (N_753,In_742,In_1366);
xnor U754 (N_754,In_62,In_1226);
or U755 (N_755,In_335,In_821);
xnor U756 (N_756,In_1367,In_1223);
and U757 (N_757,In_1288,In_1303);
or U758 (N_758,In_960,In_1490);
or U759 (N_759,In_232,In_327);
xor U760 (N_760,In_1180,In_383);
nor U761 (N_761,In_1431,In_601);
nand U762 (N_762,In_1369,In_84);
nand U763 (N_763,In_424,In_419);
xor U764 (N_764,In_148,In_757);
nor U765 (N_765,In_68,In_815);
and U766 (N_766,In_47,In_570);
xnor U767 (N_767,In_1247,In_728);
xor U768 (N_768,In_597,In_237);
and U769 (N_769,In_39,In_573);
xnor U770 (N_770,In_616,In_721);
nand U771 (N_771,In_305,In_599);
nor U772 (N_772,In_33,In_849);
xor U773 (N_773,In_1318,In_249);
xor U774 (N_774,In_400,In_81);
xnor U775 (N_775,In_1323,In_273);
nand U776 (N_776,In_1366,In_235);
nor U777 (N_777,In_603,In_207);
and U778 (N_778,In_452,In_309);
and U779 (N_779,In_1286,In_930);
xor U780 (N_780,In_611,In_690);
and U781 (N_781,In_364,In_353);
xnor U782 (N_782,In_626,In_396);
nand U783 (N_783,In_486,In_366);
nand U784 (N_784,In_1044,In_348);
or U785 (N_785,In_1490,In_1242);
or U786 (N_786,In_885,In_798);
nand U787 (N_787,In_296,In_105);
or U788 (N_788,In_80,In_564);
xnor U789 (N_789,In_655,In_1428);
xnor U790 (N_790,In_1233,In_145);
nand U791 (N_791,In_378,In_420);
or U792 (N_792,In_1226,In_1021);
or U793 (N_793,In_1456,In_436);
nor U794 (N_794,In_79,In_357);
nor U795 (N_795,In_71,In_1046);
xor U796 (N_796,In_606,In_682);
xnor U797 (N_797,In_1295,In_1459);
and U798 (N_798,In_913,In_527);
nand U799 (N_799,In_272,In_1481);
xnor U800 (N_800,In_982,In_1335);
nand U801 (N_801,In_1158,In_706);
xor U802 (N_802,In_863,In_332);
or U803 (N_803,In_920,In_2);
xor U804 (N_804,In_1037,In_1437);
nor U805 (N_805,In_425,In_906);
nand U806 (N_806,In_1477,In_61);
nor U807 (N_807,In_22,In_509);
xnor U808 (N_808,In_756,In_41);
or U809 (N_809,In_902,In_237);
xnor U810 (N_810,In_1427,In_648);
nor U811 (N_811,In_1235,In_1249);
and U812 (N_812,In_141,In_337);
xor U813 (N_813,In_626,In_506);
nand U814 (N_814,In_452,In_550);
xor U815 (N_815,In_196,In_1176);
or U816 (N_816,In_1025,In_1017);
or U817 (N_817,In_285,In_632);
nor U818 (N_818,In_1380,In_1344);
nor U819 (N_819,In_400,In_1004);
nand U820 (N_820,In_983,In_63);
nand U821 (N_821,In_1307,In_100);
and U822 (N_822,In_1417,In_681);
or U823 (N_823,In_1445,In_410);
nor U824 (N_824,In_547,In_1096);
nand U825 (N_825,In_1031,In_1311);
nor U826 (N_826,In_351,In_1098);
xor U827 (N_827,In_748,In_9);
nand U828 (N_828,In_478,In_1402);
nor U829 (N_829,In_1450,In_1229);
or U830 (N_830,In_1156,In_1258);
nor U831 (N_831,In_682,In_1482);
nor U832 (N_832,In_781,In_316);
xor U833 (N_833,In_682,In_942);
or U834 (N_834,In_627,In_111);
nand U835 (N_835,In_114,In_1424);
or U836 (N_836,In_198,In_208);
nand U837 (N_837,In_281,In_270);
nor U838 (N_838,In_1271,In_177);
xor U839 (N_839,In_49,In_1113);
nand U840 (N_840,In_1287,In_38);
and U841 (N_841,In_692,In_969);
or U842 (N_842,In_1142,In_1098);
xnor U843 (N_843,In_1207,In_68);
and U844 (N_844,In_988,In_242);
or U845 (N_845,In_995,In_810);
nor U846 (N_846,In_48,In_61);
xor U847 (N_847,In_907,In_511);
nand U848 (N_848,In_1395,In_1087);
and U849 (N_849,In_380,In_877);
nor U850 (N_850,In_1133,In_936);
nand U851 (N_851,In_205,In_1498);
nand U852 (N_852,In_544,In_1323);
or U853 (N_853,In_689,In_80);
nor U854 (N_854,In_1019,In_762);
and U855 (N_855,In_1173,In_526);
and U856 (N_856,In_1387,In_944);
nand U857 (N_857,In_578,In_823);
xnor U858 (N_858,In_143,In_513);
nand U859 (N_859,In_716,In_723);
or U860 (N_860,In_1455,In_1136);
nand U861 (N_861,In_1366,In_713);
xnor U862 (N_862,In_540,In_1126);
and U863 (N_863,In_186,In_436);
and U864 (N_864,In_508,In_544);
xor U865 (N_865,In_541,In_136);
or U866 (N_866,In_351,In_96);
nand U867 (N_867,In_1059,In_1261);
nor U868 (N_868,In_198,In_80);
or U869 (N_869,In_197,In_1186);
and U870 (N_870,In_21,In_436);
or U871 (N_871,In_560,In_945);
nand U872 (N_872,In_1042,In_1217);
and U873 (N_873,In_1346,In_426);
and U874 (N_874,In_1324,In_1275);
nor U875 (N_875,In_178,In_739);
nand U876 (N_876,In_758,In_732);
or U877 (N_877,In_136,In_453);
or U878 (N_878,In_1267,In_263);
and U879 (N_879,In_447,In_1359);
and U880 (N_880,In_273,In_487);
and U881 (N_881,In_1472,In_1155);
xor U882 (N_882,In_865,In_1149);
nor U883 (N_883,In_906,In_857);
or U884 (N_884,In_868,In_227);
or U885 (N_885,In_626,In_436);
and U886 (N_886,In_1314,In_644);
nand U887 (N_887,In_918,In_1490);
or U888 (N_888,In_1164,In_624);
or U889 (N_889,In_1068,In_468);
nand U890 (N_890,In_172,In_474);
xnor U891 (N_891,In_63,In_1208);
or U892 (N_892,In_410,In_202);
xnor U893 (N_893,In_282,In_807);
or U894 (N_894,In_389,In_878);
or U895 (N_895,In_1240,In_516);
or U896 (N_896,In_259,In_1043);
and U897 (N_897,In_772,In_1083);
xnor U898 (N_898,In_262,In_864);
or U899 (N_899,In_1049,In_728);
xor U900 (N_900,In_1228,In_415);
nand U901 (N_901,In_1436,In_531);
xnor U902 (N_902,In_982,In_1437);
nand U903 (N_903,In_1176,In_149);
or U904 (N_904,In_1450,In_1260);
nand U905 (N_905,In_1429,In_205);
xor U906 (N_906,In_1213,In_508);
and U907 (N_907,In_504,In_250);
and U908 (N_908,In_631,In_1358);
xnor U909 (N_909,In_1007,In_522);
and U910 (N_910,In_1378,In_206);
nand U911 (N_911,In_112,In_1006);
or U912 (N_912,In_320,In_188);
nand U913 (N_913,In_285,In_89);
and U914 (N_914,In_713,In_1264);
nand U915 (N_915,In_454,In_1050);
and U916 (N_916,In_148,In_684);
nor U917 (N_917,In_1118,In_1119);
and U918 (N_918,In_726,In_343);
nor U919 (N_919,In_1239,In_1091);
or U920 (N_920,In_589,In_985);
nor U921 (N_921,In_682,In_268);
nor U922 (N_922,In_734,In_1122);
or U923 (N_923,In_658,In_451);
nor U924 (N_924,In_1073,In_544);
and U925 (N_925,In_1275,In_612);
or U926 (N_926,In_185,In_113);
nand U927 (N_927,In_380,In_440);
nand U928 (N_928,In_223,In_1088);
and U929 (N_929,In_1373,In_68);
xnor U930 (N_930,In_475,In_435);
xor U931 (N_931,In_462,In_494);
or U932 (N_932,In_1222,In_609);
nand U933 (N_933,In_398,In_1263);
and U934 (N_934,In_841,In_507);
nor U935 (N_935,In_457,In_309);
xnor U936 (N_936,In_545,In_304);
nand U937 (N_937,In_1060,In_1479);
nand U938 (N_938,In_26,In_42);
nor U939 (N_939,In_116,In_924);
xor U940 (N_940,In_201,In_805);
nor U941 (N_941,In_83,In_1178);
and U942 (N_942,In_92,In_95);
nor U943 (N_943,In_136,In_209);
or U944 (N_944,In_939,In_747);
or U945 (N_945,In_274,In_228);
and U946 (N_946,In_57,In_503);
or U947 (N_947,In_368,In_1201);
nor U948 (N_948,In_1321,In_268);
or U949 (N_949,In_485,In_798);
or U950 (N_950,In_1106,In_832);
and U951 (N_951,In_1421,In_962);
or U952 (N_952,In_493,In_1461);
nor U953 (N_953,In_934,In_1346);
and U954 (N_954,In_487,In_351);
and U955 (N_955,In_995,In_612);
nor U956 (N_956,In_119,In_1110);
nor U957 (N_957,In_1093,In_895);
xor U958 (N_958,In_884,In_1484);
xnor U959 (N_959,In_439,In_982);
xor U960 (N_960,In_476,In_1067);
nor U961 (N_961,In_906,In_1138);
or U962 (N_962,In_1341,In_797);
or U963 (N_963,In_386,In_296);
xnor U964 (N_964,In_507,In_319);
nor U965 (N_965,In_246,In_752);
nand U966 (N_966,In_78,In_827);
or U967 (N_967,In_841,In_260);
nor U968 (N_968,In_585,In_785);
xnor U969 (N_969,In_1208,In_922);
xnor U970 (N_970,In_372,In_1387);
xnor U971 (N_971,In_571,In_1146);
or U972 (N_972,In_1130,In_1028);
nand U973 (N_973,In_103,In_804);
and U974 (N_974,In_889,In_202);
nand U975 (N_975,In_932,In_1);
nand U976 (N_976,In_872,In_1124);
nor U977 (N_977,In_830,In_1306);
nor U978 (N_978,In_600,In_954);
or U979 (N_979,In_365,In_442);
and U980 (N_980,In_1036,In_272);
nand U981 (N_981,In_183,In_82);
nand U982 (N_982,In_923,In_537);
xnor U983 (N_983,In_53,In_831);
or U984 (N_984,In_810,In_1004);
nor U985 (N_985,In_1145,In_830);
nor U986 (N_986,In_18,In_331);
and U987 (N_987,In_194,In_203);
and U988 (N_988,In_389,In_225);
or U989 (N_989,In_731,In_991);
nand U990 (N_990,In_1428,In_300);
and U991 (N_991,In_978,In_987);
or U992 (N_992,In_990,In_1111);
and U993 (N_993,In_860,In_444);
or U994 (N_994,In_1381,In_1426);
nor U995 (N_995,In_693,In_452);
xor U996 (N_996,In_1191,In_1171);
xor U997 (N_997,In_473,In_419);
or U998 (N_998,In_1255,In_1338);
nand U999 (N_999,In_583,In_1325);
or U1000 (N_1000,In_714,In_1408);
nor U1001 (N_1001,In_150,In_1366);
xor U1002 (N_1002,In_660,In_109);
nor U1003 (N_1003,In_137,In_260);
or U1004 (N_1004,In_202,In_990);
and U1005 (N_1005,In_541,In_369);
nor U1006 (N_1006,In_635,In_858);
nand U1007 (N_1007,In_875,In_895);
nand U1008 (N_1008,In_459,In_569);
nand U1009 (N_1009,In_1323,In_839);
nand U1010 (N_1010,In_382,In_1412);
nor U1011 (N_1011,In_136,In_794);
nor U1012 (N_1012,In_1134,In_436);
xnor U1013 (N_1013,In_1472,In_1020);
nor U1014 (N_1014,In_1381,In_63);
nor U1015 (N_1015,In_1174,In_906);
and U1016 (N_1016,In_358,In_927);
nor U1017 (N_1017,In_127,In_1019);
and U1018 (N_1018,In_176,In_136);
nor U1019 (N_1019,In_599,In_1361);
nor U1020 (N_1020,In_1091,In_652);
nor U1021 (N_1021,In_416,In_690);
and U1022 (N_1022,In_724,In_1359);
nor U1023 (N_1023,In_563,In_1214);
nand U1024 (N_1024,In_405,In_1012);
and U1025 (N_1025,In_859,In_615);
xor U1026 (N_1026,In_222,In_310);
or U1027 (N_1027,In_533,In_1401);
xor U1028 (N_1028,In_135,In_1094);
xor U1029 (N_1029,In_407,In_960);
xor U1030 (N_1030,In_17,In_677);
nand U1031 (N_1031,In_32,In_1311);
and U1032 (N_1032,In_722,In_980);
nor U1033 (N_1033,In_948,In_571);
and U1034 (N_1034,In_506,In_449);
or U1035 (N_1035,In_293,In_891);
xor U1036 (N_1036,In_567,In_1437);
xnor U1037 (N_1037,In_208,In_86);
nor U1038 (N_1038,In_477,In_914);
and U1039 (N_1039,In_835,In_887);
nor U1040 (N_1040,In_74,In_1391);
xnor U1041 (N_1041,In_1030,In_996);
xnor U1042 (N_1042,In_574,In_479);
xor U1043 (N_1043,In_137,In_40);
nand U1044 (N_1044,In_632,In_356);
and U1045 (N_1045,In_402,In_73);
nor U1046 (N_1046,In_987,In_1038);
nor U1047 (N_1047,In_473,In_465);
nand U1048 (N_1048,In_1467,In_428);
nor U1049 (N_1049,In_1136,In_515);
and U1050 (N_1050,In_271,In_412);
xnor U1051 (N_1051,In_85,In_475);
xor U1052 (N_1052,In_1492,In_1362);
and U1053 (N_1053,In_756,In_493);
or U1054 (N_1054,In_107,In_138);
xor U1055 (N_1055,In_150,In_746);
or U1056 (N_1056,In_595,In_62);
or U1057 (N_1057,In_608,In_917);
nor U1058 (N_1058,In_691,In_1318);
nand U1059 (N_1059,In_1206,In_217);
and U1060 (N_1060,In_1464,In_1159);
xnor U1061 (N_1061,In_988,In_450);
nor U1062 (N_1062,In_828,In_146);
and U1063 (N_1063,In_1201,In_1432);
xor U1064 (N_1064,In_478,In_1476);
nor U1065 (N_1065,In_1398,In_983);
nor U1066 (N_1066,In_759,In_1148);
nand U1067 (N_1067,In_694,In_631);
nand U1068 (N_1068,In_742,In_731);
nor U1069 (N_1069,In_681,In_525);
nand U1070 (N_1070,In_1272,In_974);
xor U1071 (N_1071,In_798,In_117);
nand U1072 (N_1072,In_218,In_1365);
or U1073 (N_1073,In_1383,In_335);
or U1074 (N_1074,In_1211,In_916);
nand U1075 (N_1075,In_611,In_1189);
nor U1076 (N_1076,In_434,In_464);
nand U1077 (N_1077,In_1104,In_357);
nor U1078 (N_1078,In_189,In_1273);
nand U1079 (N_1079,In_411,In_338);
nand U1080 (N_1080,In_1119,In_1169);
xor U1081 (N_1081,In_1070,In_167);
xnor U1082 (N_1082,In_204,In_707);
or U1083 (N_1083,In_1115,In_982);
xnor U1084 (N_1084,In_137,In_352);
and U1085 (N_1085,In_437,In_721);
nor U1086 (N_1086,In_72,In_594);
or U1087 (N_1087,In_168,In_23);
nor U1088 (N_1088,In_43,In_244);
nor U1089 (N_1089,In_1175,In_675);
and U1090 (N_1090,In_163,In_328);
and U1091 (N_1091,In_1036,In_284);
nor U1092 (N_1092,In_1055,In_1378);
or U1093 (N_1093,In_376,In_1313);
or U1094 (N_1094,In_632,In_1323);
and U1095 (N_1095,In_578,In_889);
nor U1096 (N_1096,In_1347,In_839);
or U1097 (N_1097,In_1188,In_1486);
nor U1098 (N_1098,In_816,In_1162);
nor U1099 (N_1099,In_912,In_1426);
and U1100 (N_1100,In_378,In_347);
nand U1101 (N_1101,In_213,In_1373);
xor U1102 (N_1102,In_169,In_1036);
nor U1103 (N_1103,In_1350,In_1256);
nor U1104 (N_1104,In_203,In_1005);
xnor U1105 (N_1105,In_1217,In_136);
nand U1106 (N_1106,In_780,In_722);
or U1107 (N_1107,In_310,In_1139);
nand U1108 (N_1108,In_1258,In_407);
nor U1109 (N_1109,In_601,In_1391);
and U1110 (N_1110,In_842,In_1370);
nor U1111 (N_1111,In_997,In_1048);
or U1112 (N_1112,In_982,In_1233);
or U1113 (N_1113,In_1265,In_1249);
or U1114 (N_1114,In_1140,In_493);
and U1115 (N_1115,In_1244,In_956);
or U1116 (N_1116,In_1263,In_125);
or U1117 (N_1117,In_1094,In_1117);
and U1118 (N_1118,In_913,In_502);
nand U1119 (N_1119,In_470,In_513);
nor U1120 (N_1120,In_1098,In_1360);
nand U1121 (N_1121,In_1199,In_479);
or U1122 (N_1122,In_1325,In_1130);
or U1123 (N_1123,In_777,In_1256);
and U1124 (N_1124,In_690,In_990);
xnor U1125 (N_1125,In_607,In_1279);
nand U1126 (N_1126,In_1004,In_78);
xor U1127 (N_1127,In_502,In_1473);
and U1128 (N_1128,In_965,In_134);
or U1129 (N_1129,In_886,In_1382);
xor U1130 (N_1130,In_390,In_410);
and U1131 (N_1131,In_240,In_838);
and U1132 (N_1132,In_300,In_533);
nand U1133 (N_1133,In_84,In_592);
or U1134 (N_1134,In_180,In_615);
and U1135 (N_1135,In_219,In_773);
and U1136 (N_1136,In_1224,In_1485);
and U1137 (N_1137,In_821,In_17);
nor U1138 (N_1138,In_392,In_988);
nor U1139 (N_1139,In_1102,In_1322);
nand U1140 (N_1140,In_132,In_208);
nand U1141 (N_1141,In_560,In_1052);
xor U1142 (N_1142,In_1016,In_811);
nand U1143 (N_1143,In_1004,In_777);
nor U1144 (N_1144,In_1057,In_237);
nor U1145 (N_1145,In_1259,In_1231);
and U1146 (N_1146,In_940,In_504);
xnor U1147 (N_1147,In_833,In_345);
xnor U1148 (N_1148,In_864,In_859);
and U1149 (N_1149,In_1292,In_219);
or U1150 (N_1150,In_1089,In_497);
nor U1151 (N_1151,In_995,In_730);
or U1152 (N_1152,In_379,In_1235);
nand U1153 (N_1153,In_279,In_1263);
and U1154 (N_1154,In_531,In_1319);
nand U1155 (N_1155,In_1142,In_1204);
nor U1156 (N_1156,In_1475,In_574);
xnor U1157 (N_1157,In_610,In_1103);
nand U1158 (N_1158,In_1282,In_89);
nor U1159 (N_1159,In_725,In_782);
nor U1160 (N_1160,In_114,In_1280);
nand U1161 (N_1161,In_1214,In_238);
and U1162 (N_1162,In_197,In_885);
and U1163 (N_1163,In_785,In_442);
and U1164 (N_1164,In_560,In_87);
xor U1165 (N_1165,In_786,In_1362);
nor U1166 (N_1166,In_1444,In_612);
and U1167 (N_1167,In_1027,In_438);
or U1168 (N_1168,In_1030,In_1032);
xor U1169 (N_1169,In_735,In_253);
nor U1170 (N_1170,In_1398,In_1155);
nand U1171 (N_1171,In_980,In_1117);
and U1172 (N_1172,In_842,In_878);
nand U1173 (N_1173,In_147,In_783);
xor U1174 (N_1174,In_1013,In_385);
and U1175 (N_1175,In_581,In_178);
nor U1176 (N_1176,In_749,In_1156);
and U1177 (N_1177,In_466,In_673);
xnor U1178 (N_1178,In_957,In_74);
or U1179 (N_1179,In_1294,In_436);
or U1180 (N_1180,In_880,In_897);
and U1181 (N_1181,In_88,In_1075);
or U1182 (N_1182,In_1415,In_461);
and U1183 (N_1183,In_784,In_1252);
xor U1184 (N_1184,In_1083,In_1222);
nand U1185 (N_1185,In_1381,In_675);
nand U1186 (N_1186,In_1358,In_1422);
xor U1187 (N_1187,In_95,In_827);
and U1188 (N_1188,In_1149,In_921);
and U1189 (N_1189,In_881,In_163);
nand U1190 (N_1190,In_391,In_508);
nand U1191 (N_1191,In_1473,In_1163);
nand U1192 (N_1192,In_1279,In_108);
or U1193 (N_1193,In_1223,In_994);
xor U1194 (N_1194,In_510,In_305);
or U1195 (N_1195,In_948,In_810);
nand U1196 (N_1196,In_1478,In_754);
xor U1197 (N_1197,In_1159,In_167);
nand U1198 (N_1198,In_49,In_514);
nand U1199 (N_1199,In_265,In_303);
nand U1200 (N_1200,In_228,In_1015);
nand U1201 (N_1201,In_720,In_1421);
nor U1202 (N_1202,In_1345,In_105);
xor U1203 (N_1203,In_149,In_1183);
nand U1204 (N_1204,In_1127,In_972);
or U1205 (N_1205,In_575,In_914);
xnor U1206 (N_1206,In_540,In_225);
and U1207 (N_1207,In_154,In_1127);
or U1208 (N_1208,In_1119,In_1334);
nand U1209 (N_1209,In_908,In_1094);
nor U1210 (N_1210,In_367,In_150);
or U1211 (N_1211,In_331,In_286);
xnor U1212 (N_1212,In_1098,In_328);
or U1213 (N_1213,In_172,In_411);
xor U1214 (N_1214,In_394,In_924);
nor U1215 (N_1215,In_546,In_1478);
and U1216 (N_1216,In_649,In_51);
or U1217 (N_1217,In_16,In_1172);
xor U1218 (N_1218,In_1323,In_1046);
nor U1219 (N_1219,In_854,In_1166);
or U1220 (N_1220,In_1019,In_1204);
nor U1221 (N_1221,In_1129,In_19);
and U1222 (N_1222,In_1477,In_774);
nand U1223 (N_1223,In_809,In_216);
or U1224 (N_1224,In_191,In_866);
and U1225 (N_1225,In_570,In_838);
xnor U1226 (N_1226,In_622,In_275);
xnor U1227 (N_1227,In_77,In_984);
or U1228 (N_1228,In_70,In_85);
nand U1229 (N_1229,In_953,In_1149);
nand U1230 (N_1230,In_42,In_1106);
and U1231 (N_1231,In_596,In_1209);
xor U1232 (N_1232,In_1307,In_1255);
or U1233 (N_1233,In_769,In_94);
nor U1234 (N_1234,In_1299,In_97);
nand U1235 (N_1235,In_804,In_1442);
or U1236 (N_1236,In_1447,In_1346);
or U1237 (N_1237,In_1061,In_211);
nor U1238 (N_1238,In_495,In_1307);
or U1239 (N_1239,In_292,In_665);
nand U1240 (N_1240,In_672,In_1275);
nand U1241 (N_1241,In_1281,In_692);
or U1242 (N_1242,In_260,In_621);
nor U1243 (N_1243,In_1280,In_1342);
and U1244 (N_1244,In_77,In_1397);
and U1245 (N_1245,In_1112,In_514);
and U1246 (N_1246,In_620,In_1041);
nor U1247 (N_1247,In_1377,In_1288);
nand U1248 (N_1248,In_1459,In_1426);
or U1249 (N_1249,In_451,In_1137);
xor U1250 (N_1250,In_780,In_7);
nor U1251 (N_1251,In_419,In_1108);
xnor U1252 (N_1252,In_500,In_891);
nor U1253 (N_1253,In_647,In_777);
and U1254 (N_1254,In_1318,In_169);
and U1255 (N_1255,In_351,In_798);
or U1256 (N_1256,In_234,In_553);
and U1257 (N_1257,In_699,In_1114);
nand U1258 (N_1258,In_727,In_896);
or U1259 (N_1259,In_493,In_1291);
and U1260 (N_1260,In_209,In_111);
or U1261 (N_1261,In_57,In_1068);
xor U1262 (N_1262,In_1428,In_998);
or U1263 (N_1263,In_985,In_1366);
nor U1264 (N_1264,In_205,In_611);
and U1265 (N_1265,In_518,In_544);
or U1266 (N_1266,In_58,In_1036);
nand U1267 (N_1267,In_1165,In_699);
nor U1268 (N_1268,In_965,In_937);
xor U1269 (N_1269,In_1418,In_987);
xnor U1270 (N_1270,In_470,In_517);
nor U1271 (N_1271,In_1247,In_1064);
and U1272 (N_1272,In_624,In_536);
or U1273 (N_1273,In_1301,In_569);
and U1274 (N_1274,In_405,In_713);
xnor U1275 (N_1275,In_852,In_245);
or U1276 (N_1276,In_428,In_1063);
and U1277 (N_1277,In_521,In_263);
nand U1278 (N_1278,In_840,In_990);
or U1279 (N_1279,In_260,In_20);
xnor U1280 (N_1280,In_1263,In_1338);
and U1281 (N_1281,In_154,In_959);
or U1282 (N_1282,In_1393,In_849);
nand U1283 (N_1283,In_377,In_493);
nor U1284 (N_1284,In_895,In_929);
nand U1285 (N_1285,In_847,In_912);
nand U1286 (N_1286,In_947,In_531);
xnor U1287 (N_1287,In_163,In_38);
nand U1288 (N_1288,In_1261,In_753);
or U1289 (N_1289,In_1084,In_1491);
nor U1290 (N_1290,In_414,In_616);
or U1291 (N_1291,In_687,In_1030);
nand U1292 (N_1292,In_194,In_384);
xor U1293 (N_1293,In_241,In_532);
xor U1294 (N_1294,In_155,In_597);
nor U1295 (N_1295,In_1243,In_871);
nand U1296 (N_1296,In_683,In_1062);
or U1297 (N_1297,In_489,In_1127);
and U1298 (N_1298,In_762,In_1073);
xor U1299 (N_1299,In_715,In_288);
and U1300 (N_1300,In_932,In_1458);
xor U1301 (N_1301,In_1259,In_1289);
or U1302 (N_1302,In_569,In_209);
and U1303 (N_1303,In_768,In_540);
xnor U1304 (N_1304,In_1095,In_890);
xnor U1305 (N_1305,In_517,In_126);
and U1306 (N_1306,In_1073,In_246);
nor U1307 (N_1307,In_603,In_232);
nor U1308 (N_1308,In_61,In_827);
or U1309 (N_1309,In_236,In_427);
nand U1310 (N_1310,In_64,In_700);
and U1311 (N_1311,In_605,In_425);
and U1312 (N_1312,In_169,In_367);
xor U1313 (N_1313,In_1000,In_443);
or U1314 (N_1314,In_703,In_1393);
xnor U1315 (N_1315,In_36,In_1306);
or U1316 (N_1316,In_70,In_766);
nand U1317 (N_1317,In_929,In_555);
and U1318 (N_1318,In_86,In_1417);
and U1319 (N_1319,In_1338,In_1278);
and U1320 (N_1320,In_138,In_1166);
nand U1321 (N_1321,In_283,In_1244);
nor U1322 (N_1322,In_551,In_752);
and U1323 (N_1323,In_639,In_125);
and U1324 (N_1324,In_1077,In_986);
nand U1325 (N_1325,In_251,In_1474);
and U1326 (N_1326,In_861,In_10);
nand U1327 (N_1327,In_860,In_1177);
nand U1328 (N_1328,In_505,In_1265);
xnor U1329 (N_1329,In_956,In_1374);
nand U1330 (N_1330,In_739,In_593);
nand U1331 (N_1331,In_822,In_784);
and U1332 (N_1332,In_492,In_799);
nor U1333 (N_1333,In_774,In_776);
xor U1334 (N_1334,In_303,In_335);
xor U1335 (N_1335,In_501,In_390);
nor U1336 (N_1336,In_1231,In_1473);
nand U1337 (N_1337,In_222,In_1367);
and U1338 (N_1338,In_1398,In_1374);
nand U1339 (N_1339,In_453,In_72);
nand U1340 (N_1340,In_165,In_511);
nand U1341 (N_1341,In_320,In_827);
xnor U1342 (N_1342,In_55,In_805);
and U1343 (N_1343,In_798,In_1223);
nor U1344 (N_1344,In_1189,In_143);
and U1345 (N_1345,In_775,In_170);
xnor U1346 (N_1346,In_739,In_1087);
or U1347 (N_1347,In_1087,In_683);
xnor U1348 (N_1348,In_898,In_1339);
nand U1349 (N_1349,In_1244,In_259);
and U1350 (N_1350,In_1228,In_573);
and U1351 (N_1351,In_431,In_43);
nor U1352 (N_1352,In_978,In_177);
nand U1353 (N_1353,In_1326,In_852);
nor U1354 (N_1354,In_1096,In_691);
nand U1355 (N_1355,In_232,In_29);
xor U1356 (N_1356,In_587,In_938);
nand U1357 (N_1357,In_1222,In_493);
nand U1358 (N_1358,In_555,In_145);
nand U1359 (N_1359,In_1114,In_374);
or U1360 (N_1360,In_821,In_756);
and U1361 (N_1361,In_1279,In_855);
and U1362 (N_1362,In_413,In_1102);
or U1363 (N_1363,In_797,In_923);
xnor U1364 (N_1364,In_1485,In_411);
and U1365 (N_1365,In_198,In_756);
or U1366 (N_1366,In_1197,In_457);
or U1367 (N_1367,In_1353,In_933);
and U1368 (N_1368,In_54,In_305);
xor U1369 (N_1369,In_126,In_1323);
nand U1370 (N_1370,In_1031,In_1422);
xor U1371 (N_1371,In_921,In_731);
nand U1372 (N_1372,In_458,In_680);
and U1373 (N_1373,In_1193,In_740);
nor U1374 (N_1374,In_489,In_167);
and U1375 (N_1375,In_1133,In_1132);
or U1376 (N_1376,In_785,In_1214);
nand U1377 (N_1377,In_791,In_824);
or U1378 (N_1378,In_1066,In_785);
nor U1379 (N_1379,In_35,In_1445);
xor U1380 (N_1380,In_1363,In_485);
nand U1381 (N_1381,In_474,In_696);
nand U1382 (N_1382,In_628,In_100);
nand U1383 (N_1383,In_788,In_1243);
and U1384 (N_1384,In_1420,In_510);
or U1385 (N_1385,In_1447,In_311);
nand U1386 (N_1386,In_362,In_1149);
and U1387 (N_1387,In_208,In_323);
xor U1388 (N_1388,In_936,In_518);
nand U1389 (N_1389,In_195,In_1057);
and U1390 (N_1390,In_503,In_1021);
or U1391 (N_1391,In_725,In_1353);
xor U1392 (N_1392,In_666,In_1231);
or U1393 (N_1393,In_819,In_340);
nand U1394 (N_1394,In_55,In_137);
and U1395 (N_1395,In_762,In_171);
nor U1396 (N_1396,In_927,In_519);
nor U1397 (N_1397,In_239,In_545);
and U1398 (N_1398,In_570,In_1242);
nor U1399 (N_1399,In_1141,In_946);
nand U1400 (N_1400,In_1141,In_268);
nor U1401 (N_1401,In_669,In_1274);
nand U1402 (N_1402,In_50,In_291);
or U1403 (N_1403,In_1006,In_959);
xor U1404 (N_1404,In_1303,In_1499);
nand U1405 (N_1405,In_1439,In_1137);
or U1406 (N_1406,In_1490,In_1413);
xor U1407 (N_1407,In_1084,In_166);
or U1408 (N_1408,In_1045,In_677);
and U1409 (N_1409,In_131,In_826);
and U1410 (N_1410,In_356,In_30);
nand U1411 (N_1411,In_1119,In_130);
or U1412 (N_1412,In_845,In_652);
and U1413 (N_1413,In_940,In_878);
nor U1414 (N_1414,In_1389,In_643);
nand U1415 (N_1415,In_811,In_249);
nor U1416 (N_1416,In_1398,In_234);
nor U1417 (N_1417,In_288,In_893);
and U1418 (N_1418,In_431,In_54);
xnor U1419 (N_1419,In_1067,In_609);
and U1420 (N_1420,In_636,In_391);
nand U1421 (N_1421,In_264,In_193);
and U1422 (N_1422,In_29,In_510);
nand U1423 (N_1423,In_1423,In_1487);
nor U1424 (N_1424,In_1442,In_1301);
and U1425 (N_1425,In_1195,In_137);
and U1426 (N_1426,In_645,In_1037);
xnor U1427 (N_1427,In_1447,In_1100);
and U1428 (N_1428,In_487,In_437);
nor U1429 (N_1429,In_807,In_360);
or U1430 (N_1430,In_1406,In_135);
nand U1431 (N_1431,In_1235,In_859);
nand U1432 (N_1432,In_871,In_1379);
xnor U1433 (N_1433,In_9,In_768);
nor U1434 (N_1434,In_1005,In_1297);
and U1435 (N_1435,In_829,In_665);
and U1436 (N_1436,In_1098,In_951);
nor U1437 (N_1437,In_349,In_368);
nand U1438 (N_1438,In_265,In_849);
nand U1439 (N_1439,In_715,In_669);
and U1440 (N_1440,In_1498,In_952);
xnor U1441 (N_1441,In_270,In_293);
and U1442 (N_1442,In_293,In_520);
and U1443 (N_1443,In_58,In_341);
nor U1444 (N_1444,In_928,In_386);
nor U1445 (N_1445,In_775,In_1422);
nand U1446 (N_1446,In_411,In_687);
and U1447 (N_1447,In_1117,In_174);
or U1448 (N_1448,In_122,In_1349);
xnor U1449 (N_1449,In_1251,In_717);
nand U1450 (N_1450,In_763,In_1474);
nand U1451 (N_1451,In_502,In_281);
nor U1452 (N_1452,In_1197,In_241);
nor U1453 (N_1453,In_79,In_933);
and U1454 (N_1454,In_846,In_695);
nor U1455 (N_1455,In_596,In_617);
xor U1456 (N_1456,In_1028,In_210);
or U1457 (N_1457,In_227,In_752);
xnor U1458 (N_1458,In_864,In_243);
and U1459 (N_1459,In_295,In_869);
or U1460 (N_1460,In_725,In_439);
nand U1461 (N_1461,In_995,In_5);
xnor U1462 (N_1462,In_162,In_1121);
and U1463 (N_1463,In_376,In_1371);
or U1464 (N_1464,In_1176,In_1298);
nand U1465 (N_1465,In_1401,In_135);
xor U1466 (N_1466,In_380,In_1047);
or U1467 (N_1467,In_1394,In_1429);
nand U1468 (N_1468,In_538,In_511);
and U1469 (N_1469,In_776,In_471);
xor U1470 (N_1470,In_662,In_692);
nand U1471 (N_1471,In_901,In_300);
xnor U1472 (N_1472,In_958,In_1207);
nor U1473 (N_1473,In_875,In_283);
xor U1474 (N_1474,In_1490,In_322);
and U1475 (N_1475,In_495,In_344);
xnor U1476 (N_1476,In_300,In_630);
or U1477 (N_1477,In_399,In_367);
or U1478 (N_1478,In_1028,In_458);
nand U1479 (N_1479,In_606,In_873);
xor U1480 (N_1480,In_157,In_858);
xnor U1481 (N_1481,In_418,In_550);
and U1482 (N_1482,In_459,In_325);
nor U1483 (N_1483,In_1428,In_66);
nand U1484 (N_1484,In_360,In_1183);
or U1485 (N_1485,In_1101,In_72);
or U1486 (N_1486,In_774,In_318);
xor U1487 (N_1487,In_1456,In_830);
nor U1488 (N_1488,In_1087,In_949);
nand U1489 (N_1489,In_851,In_1196);
nand U1490 (N_1490,In_381,In_791);
nand U1491 (N_1491,In_1403,In_219);
xor U1492 (N_1492,In_287,In_931);
nand U1493 (N_1493,In_987,In_813);
nor U1494 (N_1494,In_693,In_31);
or U1495 (N_1495,In_1021,In_272);
or U1496 (N_1496,In_937,In_1253);
and U1497 (N_1497,In_1304,In_707);
nand U1498 (N_1498,In_1139,In_1471);
and U1499 (N_1499,In_462,In_1471);
or U1500 (N_1500,In_503,In_863);
or U1501 (N_1501,In_1001,In_577);
xor U1502 (N_1502,In_545,In_1000);
and U1503 (N_1503,In_521,In_1179);
nor U1504 (N_1504,In_143,In_1308);
and U1505 (N_1505,In_628,In_34);
xnor U1506 (N_1506,In_1339,In_1149);
xnor U1507 (N_1507,In_134,In_656);
and U1508 (N_1508,In_21,In_1439);
nor U1509 (N_1509,In_136,In_345);
and U1510 (N_1510,In_477,In_309);
nand U1511 (N_1511,In_126,In_778);
or U1512 (N_1512,In_1061,In_1475);
xnor U1513 (N_1513,In_855,In_1114);
nor U1514 (N_1514,In_1411,In_141);
nor U1515 (N_1515,In_828,In_388);
xnor U1516 (N_1516,In_540,In_167);
or U1517 (N_1517,In_895,In_731);
or U1518 (N_1518,In_869,In_950);
nand U1519 (N_1519,In_1462,In_993);
nor U1520 (N_1520,In_1123,In_1411);
nand U1521 (N_1521,In_59,In_384);
or U1522 (N_1522,In_24,In_805);
nand U1523 (N_1523,In_1091,In_74);
and U1524 (N_1524,In_993,In_1126);
xor U1525 (N_1525,In_1105,In_658);
xor U1526 (N_1526,In_717,In_976);
xnor U1527 (N_1527,In_1409,In_102);
nor U1528 (N_1528,In_657,In_1399);
or U1529 (N_1529,In_993,In_1020);
nor U1530 (N_1530,In_608,In_1237);
and U1531 (N_1531,In_393,In_979);
nand U1532 (N_1532,In_921,In_1392);
or U1533 (N_1533,In_198,In_1156);
or U1534 (N_1534,In_364,In_248);
and U1535 (N_1535,In_49,In_1228);
or U1536 (N_1536,In_1451,In_1156);
nand U1537 (N_1537,In_227,In_387);
nor U1538 (N_1538,In_167,In_33);
or U1539 (N_1539,In_655,In_1036);
xnor U1540 (N_1540,In_739,In_792);
and U1541 (N_1541,In_327,In_399);
nor U1542 (N_1542,In_392,In_278);
and U1543 (N_1543,In_804,In_249);
or U1544 (N_1544,In_425,In_344);
or U1545 (N_1545,In_733,In_1203);
xnor U1546 (N_1546,In_1159,In_1339);
nand U1547 (N_1547,In_1257,In_561);
or U1548 (N_1548,In_1479,In_1436);
nor U1549 (N_1549,In_34,In_675);
and U1550 (N_1550,In_5,In_1066);
or U1551 (N_1551,In_833,In_1095);
or U1552 (N_1552,In_595,In_991);
nand U1553 (N_1553,In_728,In_453);
nor U1554 (N_1554,In_83,In_1108);
nand U1555 (N_1555,In_432,In_1159);
nand U1556 (N_1556,In_516,In_1415);
xnor U1557 (N_1557,In_1321,In_812);
nand U1558 (N_1558,In_1335,In_1138);
nand U1559 (N_1559,In_586,In_354);
and U1560 (N_1560,In_1274,In_1463);
or U1561 (N_1561,In_720,In_820);
and U1562 (N_1562,In_115,In_90);
or U1563 (N_1563,In_299,In_194);
or U1564 (N_1564,In_325,In_90);
or U1565 (N_1565,In_686,In_481);
xor U1566 (N_1566,In_1351,In_129);
and U1567 (N_1567,In_1138,In_782);
nor U1568 (N_1568,In_22,In_1256);
nor U1569 (N_1569,In_386,In_995);
nand U1570 (N_1570,In_376,In_1312);
and U1571 (N_1571,In_368,In_485);
xnor U1572 (N_1572,In_1455,In_199);
nor U1573 (N_1573,In_783,In_1400);
and U1574 (N_1574,In_231,In_1013);
or U1575 (N_1575,In_372,In_1487);
nor U1576 (N_1576,In_208,In_244);
xnor U1577 (N_1577,In_232,In_719);
xnor U1578 (N_1578,In_991,In_964);
xor U1579 (N_1579,In_1363,In_678);
nor U1580 (N_1580,In_86,In_1147);
and U1581 (N_1581,In_884,In_379);
or U1582 (N_1582,In_25,In_1001);
and U1583 (N_1583,In_137,In_562);
nor U1584 (N_1584,In_703,In_1463);
xnor U1585 (N_1585,In_1271,In_1088);
or U1586 (N_1586,In_724,In_1012);
xor U1587 (N_1587,In_942,In_1383);
nor U1588 (N_1588,In_1446,In_1473);
nor U1589 (N_1589,In_272,In_994);
xor U1590 (N_1590,In_373,In_1180);
nor U1591 (N_1591,In_914,In_292);
nand U1592 (N_1592,In_642,In_606);
or U1593 (N_1593,In_1243,In_1136);
or U1594 (N_1594,In_553,In_187);
nor U1595 (N_1595,In_481,In_506);
or U1596 (N_1596,In_96,In_767);
nor U1597 (N_1597,In_1100,In_1109);
and U1598 (N_1598,In_1354,In_315);
nor U1599 (N_1599,In_80,In_603);
or U1600 (N_1600,In_1172,In_441);
or U1601 (N_1601,In_1229,In_661);
xor U1602 (N_1602,In_832,In_431);
nor U1603 (N_1603,In_881,In_766);
xnor U1604 (N_1604,In_17,In_894);
or U1605 (N_1605,In_192,In_284);
xor U1606 (N_1606,In_1309,In_236);
nor U1607 (N_1607,In_580,In_787);
nand U1608 (N_1608,In_1135,In_184);
nand U1609 (N_1609,In_545,In_1363);
nor U1610 (N_1610,In_1450,In_937);
xor U1611 (N_1611,In_392,In_299);
or U1612 (N_1612,In_361,In_344);
and U1613 (N_1613,In_1442,In_842);
nor U1614 (N_1614,In_749,In_309);
or U1615 (N_1615,In_1154,In_1275);
or U1616 (N_1616,In_351,In_401);
and U1617 (N_1617,In_1435,In_539);
nor U1618 (N_1618,In_1241,In_947);
and U1619 (N_1619,In_1065,In_426);
xnor U1620 (N_1620,In_372,In_1360);
xor U1621 (N_1621,In_74,In_90);
nand U1622 (N_1622,In_1237,In_392);
nor U1623 (N_1623,In_724,In_601);
or U1624 (N_1624,In_1134,In_1329);
or U1625 (N_1625,In_414,In_1317);
or U1626 (N_1626,In_385,In_996);
or U1627 (N_1627,In_218,In_907);
or U1628 (N_1628,In_1404,In_1492);
and U1629 (N_1629,In_742,In_1044);
or U1630 (N_1630,In_1270,In_617);
nor U1631 (N_1631,In_392,In_549);
xnor U1632 (N_1632,In_86,In_354);
or U1633 (N_1633,In_82,In_1290);
or U1634 (N_1634,In_1478,In_392);
or U1635 (N_1635,In_682,In_164);
and U1636 (N_1636,In_1013,In_770);
nor U1637 (N_1637,In_499,In_27);
and U1638 (N_1638,In_561,In_1034);
nand U1639 (N_1639,In_1422,In_496);
and U1640 (N_1640,In_571,In_342);
nor U1641 (N_1641,In_17,In_544);
nor U1642 (N_1642,In_71,In_1303);
nor U1643 (N_1643,In_915,In_1437);
and U1644 (N_1644,In_503,In_1187);
nor U1645 (N_1645,In_1040,In_655);
or U1646 (N_1646,In_402,In_99);
nand U1647 (N_1647,In_944,In_568);
xor U1648 (N_1648,In_268,In_551);
or U1649 (N_1649,In_436,In_1327);
or U1650 (N_1650,In_126,In_610);
xor U1651 (N_1651,In_1453,In_1074);
xor U1652 (N_1652,In_879,In_356);
xor U1653 (N_1653,In_1446,In_426);
or U1654 (N_1654,In_847,In_893);
and U1655 (N_1655,In_476,In_116);
xor U1656 (N_1656,In_1198,In_73);
and U1657 (N_1657,In_709,In_958);
xnor U1658 (N_1658,In_279,In_1289);
or U1659 (N_1659,In_1062,In_1446);
xnor U1660 (N_1660,In_242,In_876);
or U1661 (N_1661,In_1227,In_82);
nor U1662 (N_1662,In_924,In_753);
nor U1663 (N_1663,In_1493,In_406);
nor U1664 (N_1664,In_191,In_1290);
nand U1665 (N_1665,In_1312,In_232);
nor U1666 (N_1666,In_1027,In_642);
nor U1667 (N_1667,In_1106,In_1423);
or U1668 (N_1668,In_613,In_934);
or U1669 (N_1669,In_106,In_393);
or U1670 (N_1670,In_781,In_454);
or U1671 (N_1671,In_745,In_644);
nor U1672 (N_1672,In_896,In_309);
xor U1673 (N_1673,In_1076,In_602);
or U1674 (N_1674,In_95,In_779);
nor U1675 (N_1675,In_1036,In_761);
or U1676 (N_1676,In_721,In_445);
and U1677 (N_1677,In_99,In_627);
and U1678 (N_1678,In_251,In_1303);
nand U1679 (N_1679,In_42,In_554);
xor U1680 (N_1680,In_542,In_629);
nand U1681 (N_1681,In_1233,In_1308);
or U1682 (N_1682,In_1129,In_1341);
xnor U1683 (N_1683,In_89,In_1445);
nor U1684 (N_1684,In_259,In_339);
xnor U1685 (N_1685,In_130,In_1044);
nand U1686 (N_1686,In_293,In_993);
xnor U1687 (N_1687,In_910,In_741);
nor U1688 (N_1688,In_954,In_586);
or U1689 (N_1689,In_611,In_908);
and U1690 (N_1690,In_628,In_1204);
and U1691 (N_1691,In_828,In_375);
xor U1692 (N_1692,In_92,In_324);
xor U1693 (N_1693,In_43,In_1383);
xor U1694 (N_1694,In_1488,In_1292);
or U1695 (N_1695,In_759,In_1442);
xor U1696 (N_1696,In_732,In_770);
and U1697 (N_1697,In_197,In_1019);
nor U1698 (N_1698,In_990,In_717);
or U1699 (N_1699,In_231,In_148);
and U1700 (N_1700,In_59,In_1362);
nand U1701 (N_1701,In_36,In_385);
and U1702 (N_1702,In_337,In_1214);
or U1703 (N_1703,In_518,In_857);
xnor U1704 (N_1704,In_233,In_1126);
nand U1705 (N_1705,In_532,In_266);
nand U1706 (N_1706,In_1174,In_492);
and U1707 (N_1707,In_872,In_176);
and U1708 (N_1708,In_1087,In_648);
or U1709 (N_1709,In_705,In_706);
and U1710 (N_1710,In_1239,In_1132);
nor U1711 (N_1711,In_394,In_800);
nand U1712 (N_1712,In_1011,In_871);
or U1713 (N_1713,In_1059,In_1152);
and U1714 (N_1714,In_1379,In_1468);
nand U1715 (N_1715,In_1249,In_516);
nor U1716 (N_1716,In_296,In_175);
xnor U1717 (N_1717,In_248,In_559);
nand U1718 (N_1718,In_968,In_1201);
nor U1719 (N_1719,In_1200,In_954);
nor U1720 (N_1720,In_811,In_660);
and U1721 (N_1721,In_252,In_1196);
nand U1722 (N_1722,In_735,In_638);
and U1723 (N_1723,In_879,In_294);
nand U1724 (N_1724,In_439,In_1497);
nand U1725 (N_1725,In_1411,In_1364);
nand U1726 (N_1726,In_199,In_656);
nor U1727 (N_1727,In_1468,In_27);
xnor U1728 (N_1728,In_437,In_80);
or U1729 (N_1729,In_617,In_161);
or U1730 (N_1730,In_1234,In_1395);
or U1731 (N_1731,In_580,In_1364);
or U1732 (N_1732,In_410,In_1067);
and U1733 (N_1733,In_1453,In_704);
or U1734 (N_1734,In_1085,In_997);
or U1735 (N_1735,In_638,In_492);
and U1736 (N_1736,In_287,In_953);
and U1737 (N_1737,In_1494,In_1246);
nor U1738 (N_1738,In_208,In_822);
nand U1739 (N_1739,In_1181,In_408);
nor U1740 (N_1740,In_264,In_1369);
nand U1741 (N_1741,In_105,In_397);
nor U1742 (N_1742,In_556,In_1151);
and U1743 (N_1743,In_1247,In_810);
or U1744 (N_1744,In_1095,In_0);
and U1745 (N_1745,In_310,In_209);
nor U1746 (N_1746,In_80,In_509);
nand U1747 (N_1747,In_705,In_770);
nand U1748 (N_1748,In_404,In_1295);
and U1749 (N_1749,In_1398,In_133);
and U1750 (N_1750,In_1320,In_852);
nor U1751 (N_1751,In_715,In_710);
nand U1752 (N_1752,In_1491,In_1161);
nand U1753 (N_1753,In_313,In_1194);
and U1754 (N_1754,In_453,In_568);
and U1755 (N_1755,In_1162,In_1205);
or U1756 (N_1756,In_1248,In_79);
nand U1757 (N_1757,In_353,In_735);
and U1758 (N_1758,In_931,In_67);
nor U1759 (N_1759,In_764,In_735);
and U1760 (N_1760,In_459,In_1429);
xor U1761 (N_1761,In_1031,In_222);
or U1762 (N_1762,In_224,In_1457);
xnor U1763 (N_1763,In_195,In_471);
or U1764 (N_1764,In_1382,In_950);
or U1765 (N_1765,In_761,In_1309);
nor U1766 (N_1766,In_902,In_1249);
nand U1767 (N_1767,In_1288,In_271);
xor U1768 (N_1768,In_531,In_831);
or U1769 (N_1769,In_478,In_1310);
and U1770 (N_1770,In_5,In_1310);
nand U1771 (N_1771,In_765,In_911);
nand U1772 (N_1772,In_981,In_925);
and U1773 (N_1773,In_439,In_1000);
or U1774 (N_1774,In_1260,In_1078);
xnor U1775 (N_1775,In_587,In_113);
nor U1776 (N_1776,In_1330,In_747);
or U1777 (N_1777,In_484,In_27);
or U1778 (N_1778,In_992,In_364);
and U1779 (N_1779,In_723,In_1128);
nand U1780 (N_1780,In_940,In_1230);
nand U1781 (N_1781,In_1119,In_163);
and U1782 (N_1782,In_1467,In_1222);
and U1783 (N_1783,In_608,In_1461);
xor U1784 (N_1784,In_1043,In_450);
nand U1785 (N_1785,In_454,In_1493);
xnor U1786 (N_1786,In_1138,In_823);
and U1787 (N_1787,In_1405,In_55);
xnor U1788 (N_1788,In_328,In_408);
nand U1789 (N_1789,In_535,In_1137);
nand U1790 (N_1790,In_6,In_755);
nand U1791 (N_1791,In_962,In_549);
xnor U1792 (N_1792,In_1141,In_715);
xor U1793 (N_1793,In_1398,In_1151);
xor U1794 (N_1794,In_673,In_761);
nand U1795 (N_1795,In_1421,In_650);
nor U1796 (N_1796,In_121,In_810);
nand U1797 (N_1797,In_373,In_918);
nand U1798 (N_1798,In_1171,In_685);
nand U1799 (N_1799,In_475,In_748);
nand U1800 (N_1800,In_365,In_382);
nand U1801 (N_1801,In_444,In_1185);
or U1802 (N_1802,In_442,In_1280);
or U1803 (N_1803,In_248,In_1289);
and U1804 (N_1804,In_1374,In_291);
nand U1805 (N_1805,In_808,In_1252);
and U1806 (N_1806,In_1454,In_421);
and U1807 (N_1807,In_151,In_425);
nor U1808 (N_1808,In_366,In_170);
and U1809 (N_1809,In_1463,In_1057);
or U1810 (N_1810,In_624,In_758);
nand U1811 (N_1811,In_529,In_1006);
nand U1812 (N_1812,In_1164,In_1379);
or U1813 (N_1813,In_409,In_77);
xnor U1814 (N_1814,In_45,In_540);
xnor U1815 (N_1815,In_792,In_89);
or U1816 (N_1816,In_1031,In_1270);
nor U1817 (N_1817,In_1127,In_506);
xor U1818 (N_1818,In_595,In_269);
nor U1819 (N_1819,In_997,In_749);
nor U1820 (N_1820,In_114,In_1288);
and U1821 (N_1821,In_878,In_1439);
nand U1822 (N_1822,In_693,In_1261);
xnor U1823 (N_1823,In_1015,In_1145);
or U1824 (N_1824,In_1283,In_1219);
or U1825 (N_1825,In_1413,In_1459);
xor U1826 (N_1826,In_1073,In_646);
or U1827 (N_1827,In_595,In_1420);
and U1828 (N_1828,In_1401,In_760);
nor U1829 (N_1829,In_822,In_1202);
xor U1830 (N_1830,In_1030,In_860);
nor U1831 (N_1831,In_455,In_206);
xnor U1832 (N_1832,In_637,In_719);
and U1833 (N_1833,In_287,In_1381);
nor U1834 (N_1834,In_623,In_1);
or U1835 (N_1835,In_285,In_979);
nand U1836 (N_1836,In_1267,In_1011);
or U1837 (N_1837,In_609,In_1175);
or U1838 (N_1838,In_1426,In_973);
or U1839 (N_1839,In_1409,In_1323);
xnor U1840 (N_1840,In_992,In_681);
nand U1841 (N_1841,In_634,In_267);
xnor U1842 (N_1842,In_1186,In_1059);
or U1843 (N_1843,In_970,In_122);
nand U1844 (N_1844,In_582,In_357);
or U1845 (N_1845,In_980,In_1253);
nor U1846 (N_1846,In_1137,In_1462);
and U1847 (N_1847,In_1360,In_1282);
nor U1848 (N_1848,In_757,In_1472);
nor U1849 (N_1849,In_1426,In_510);
nand U1850 (N_1850,In_912,In_1034);
or U1851 (N_1851,In_715,In_1009);
or U1852 (N_1852,In_388,In_954);
nor U1853 (N_1853,In_1298,In_775);
nand U1854 (N_1854,In_1128,In_1091);
or U1855 (N_1855,In_303,In_1160);
nor U1856 (N_1856,In_566,In_590);
nand U1857 (N_1857,In_181,In_1202);
xnor U1858 (N_1858,In_1073,In_1243);
nor U1859 (N_1859,In_697,In_1039);
nor U1860 (N_1860,In_698,In_438);
and U1861 (N_1861,In_350,In_798);
nand U1862 (N_1862,In_826,In_127);
or U1863 (N_1863,In_546,In_789);
and U1864 (N_1864,In_1491,In_1406);
nand U1865 (N_1865,In_543,In_793);
nand U1866 (N_1866,In_1044,In_174);
nand U1867 (N_1867,In_843,In_17);
and U1868 (N_1868,In_1265,In_225);
nor U1869 (N_1869,In_881,In_409);
and U1870 (N_1870,In_1276,In_140);
or U1871 (N_1871,In_311,In_921);
nand U1872 (N_1872,In_994,In_1407);
and U1873 (N_1873,In_750,In_353);
and U1874 (N_1874,In_120,In_1295);
nor U1875 (N_1875,In_29,In_1288);
xor U1876 (N_1876,In_558,In_572);
or U1877 (N_1877,In_647,In_1353);
xor U1878 (N_1878,In_536,In_1429);
and U1879 (N_1879,In_550,In_506);
xnor U1880 (N_1880,In_584,In_960);
nor U1881 (N_1881,In_1185,In_499);
nor U1882 (N_1882,In_1495,In_85);
and U1883 (N_1883,In_8,In_205);
nand U1884 (N_1884,In_101,In_1284);
and U1885 (N_1885,In_1433,In_972);
nor U1886 (N_1886,In_882,In_1220);
and U1887 (N_1887,In_564,In_331);
and U1888 (N_1888,In_1277,In_778);
xnor U1889 (N_1889,In_584,In_781);
nand U1890 (N_1890,In_41,In_1186);
or U1891 (N_1891,In_232,In_1271);
nand U1892 (N_1892,In_1453,In_829);
nand U1893 (N_1893,In_621,In_1035);
and U1894 (N_1894,In_406,In_1202);
and U1895 (N_1895,In_146,In_35);
nand U1896 (N_1896,In_939,In_212);
or U1897 (N_1897,In_370,In_237);
nor U1898 (N_1898,In_1439,In_1131);
and U1899 (N_1899,In_574,In_894);
or U1900 (N_1900,In_1447,In_1439);
nor U1901 (N_1901,In_1387,In_953);
nor U1902 (N_1902,In_1312,In_567);
or U1903 (N_1903,In_82,In_625);
nand U1904 (N_1904,In_1432,In_1153);
and U1905 (N_1905,In_697,In_1093);
nor U1906 (N_1906,In_599,In_762);
xnor U1907 (N_1907,In_1318,In_94);
nor U1908 (N_1908,In_1346,In_82);
nor U1909 (N_1909,In_737,In_861);
nor U1910 (N_1910,In_1260,In_297);
nand U1911 (N_1911,In_406,In_595);
or U1912 (N_1912,In_353,In_82);
and U1913 (N_1913,In_1172,In_902);
nand U1914 (N_1914,In_569,In_820);
nor U1915 (N_1915,In_1243,In_123);
and U1916 (N_1916,In_123,In_66);
or U1917 (N_1917,In_429,In_1489);
xnor U1918 (N_1918,In_681,In_1222);
or U1919 (N_1919,In_93,In_701);
and U1920 (N_1920,In_246,In_1405);
nor U1921 (N_1921,In_546,In_541);
or U1922 (N_1922,In_997,In_1425);
nor U1923 (N_1923,In_1372,In_720);
or U1924 (N_1924,In_181,In_1065);
and U1925 (N_1925,In_1047,In_60);
nand U1926 (N_1926,In_350,In_790);
nor U1927 (N_1927,In_217,In_1237);
nand U1928 (N_1928,In_530,In_1227);
xor U1929 (N_1929,In_1060,In_545);
or U1930 (N_1930,In_196,In_1281);
and U1931 (N_1931,In_1288,In_226);
nand U1932 (N_1932,In_554,In_296);
xnor U1933 (N_1933,In_124,In_1149);
and U1934 (N_1934,In_1130,In_1171);
or U1935 (N_1935,In_961,In_795);
or U1936 (N_1936,In_852,In_215);
or U1937 (N_1937,In_1456,In_1266);
nand U1938 (N_1938,In_1043,In_93);
nor U1939 (N_1939,In_45,In_1392);
nor U1940 (N_1940,In_914,In_1414);
nand U1941 (N_1941,In_1203,In_472);
xnor U1942 (N_1942,In_1231,In_318);
nand U1943 (N_1943,In_947,In_443);
or U1944 (N_1944,In_49,In_411);
and U1945 (N_1945,In_903,In_316);
and U1946 (N_1946,In_900,In_1399);
or U1947 (N_1947,In_110,In_1271);
or U1948 (N_1948,In_1195,In_210);
nor U1949 (N_1949,In_833,In_422);
or U1950 (N_1950,In_207,In_1185);
or U1951 (N_1951,In_135,In_1185);
xnor U1952 (N_1952,In_3,In_538);
and U1953 (N_1953,In_1152,In_313);
nand U1954 (N_1954,In_375,In_517);
nand U1955 (N_1955,In_750,In_173);
xnor U1956 (N_1956,In_1326,In_970);
or U1957 (N_1957,In_1006,In_844);
and U1958 (N_1958,In_637,In_973);
nand U1959 (N_1959,In_971,In_1061);
xnor U1960 (N_1960,In_641,In_1153);
and U1961 (N_1961,In_1361,In_592);
or U1962 (N_1962,In_657,In_185);
nor U1963 (N_1963,In_354,In_564);
and U1964 (N_1964,In_316,In_0);
or U1965 (N_1965,In_806,In_1057);
nand U1966 (N_1966,In_1261,In_34);
and U1967 (N_1967,In_459,In_594);
nor U1968 (N_1968,In_1099,In_1434);
or U1969 (N_1969,In_1057,In_74);
nor U1970 (N_1970,In_1003,In_43);
nand U1971 (N_1971,In_619,In_202);
and U1972 (N_1972,In_1105,In_1403);
nor U1973 (N_1973,In_605,In_1349);
nor U1974 (N_1974,In_1020,In_1391);
nand U1975 (N_1975,In_820,In_119);
and U1976 (N_1976,In_846,In_963);
nand U1977 (N_1977,In_814,In_762);
nor U1978 (N_1978,In_1077,In_1434);
nor U1979 (N_1979,In_1276,In_1245);
or U1980 (N_1980,In_235,In_1268);
xnor U1981 (N_1981,In_1356,In_1204);
or U1982 (N_1982,In_358,In_736);
and U1983 (N_1983,In_870,In_279);
nand U1984 (N_1984,In_1123,In_180);
nor U1985 (N_1985,In_741,In_662);
nand U1986 (N_1986,In_216,In_932);
xor U1987 (N_1987,In_363,In_907);
nor U1988 (N_1988,In_473,In_944);
and U1989 (N_1989,In_1360,In_251);
nor U1990 (N_1990,In_1287,In_464);
nand U1991 (N_1991,In_1268,In_699);
nand U1992 (N_1992,In_1443,In_1444);
nand U1993 (N_1993,In_1404,In_566);
nand U1994 (N_1994,In_1499,In_838);
nor U1995 (N_1995,In_495,In_1262);
nand U1996 (N_1996,In_352,In_1043);
xnor U1997 (N_1997,In_301,In_501);
nand U1998 (N_1998,In_319,In_1191);
or U1999 (N_1999,In_710,In_1314);
or U2000 (N_2000,In_1386,In_957);
or U2001 (N_2001,In_296,In_131);
and U2002 (N_2002,In_444,In_1283);
nand U2003 (N_2003,In_311,In_776);
nand U2004 (N_2004,In_1489,In_332);
nand U2005 (N_2005,In_804,In_1427);
nand U2006 (N_2006,In_1397,In_505);
nand U2007 (N_2007,In_18,In_728);
and U2008 (N_2008,In_265,In_191);
or U2009 (N_2009,In_190,In_1287);
and U2010 (N_2010,In_1148,In_1296);
or U2011 (N_2011,In_918,In_189);
xnor U2012 (N_2012,In_442,In_238);
xor U2013 (N_2013,In_692,In_1256);
nor U2014 (N_2014,In_961,In_98);
nor U2015 (N_2015,In_29,In_442);
xor U2016 (N_2016,In_277,In_1495);
nand U2017 (N_2017,In_303,In_953);
or U2018 (N_2018,In_1369,In_732);
nand U2019 (N_2019,In_454,In_25);
xor U2020 (N_2020,In_865,In_1092);
or U2021 (N_2021,In_689,In_1300);
and U2022 (N_2022,In_1470,In_657);
or U2023 (N_2023,In_956,In_602);
nor U2024 (N_2024,In_1474,In_1038);
nand U2025 (N_2025,In_337,In_1417);
nor U2026 (N_2026,In_1120,In_315);
xor U2027 (N_2027,In_1384,In_762);
xor U2028 (N_2028,In_526,In_456);
nand U2029 (N_2029,In_417,In_1158);
xnor U2030 (N_2030,In_1378,In_350);
nand U2031 (N_2031,In_1469,In_553);
and U2032 (N_2032,In_691,In_1439);
or U2033 (N_2033,In_196,In_249);
nor U2034 (N_2034,In_254,In_245);
nor U2035 (N_2035,In_108,In_340);
nor U2036 (N_2036,In_580,In_1267);
xnor U2037 (N_2037,In_406,In_704);
or U2038 (N_2038,In_229,In_270);
or U2039 (N_2039,In_749,In_831);
nor U2040 (N_2040,In_270,In_555);
nand U2041 (N_2041,In_665,In_1272);
and U2042 (N_2042,In_679,In_1485);
and U2043 (N_2043,In_1466,In_1023);
or U2044 (N_2044,In_832,In_46);
nand U2045 (N_2045,In_528,In_318);
or U2046 (N_2046,In_1363,In_1230);
nor U2047 (N_2047,In_1068,In_1178);
and U2048 (N_2048,In_894,In_303);
nor U2049 (N_2049,In_1326,In_664);
and U2050 (N_2050,In_1186,In_275);
xor U2051 (N_2051,In_650,In_326);
nor U2052 (N_2052,In_1240,In_748);
xor U2053 (N_2053,In_277,In_779);
xnor U2054 (N_2054,In_1070,In_406);
nor U2055 (N_2055,In_75,In_275);
nor U2056 (N_2056,In_11,In_531);
or U2057 (N_2057,In_497,In_1222);
nand U2058 (N_2058,In_1444,In_954);
and U2059 (N_2059,In_536,In_1036);
and U2060 (N_2060,In_531,In_496);
or U2061 (N_2061,In_804,In_816);
nor U2062 (N_2062,In_866,In_993);
or U2063 (N_2063,In_1236,In_1143);
nand U2064 (N_2064,In_563,In_1295);
xor U2065 (N_2065,In_769,In_1353);
nor U2066 (N_2066,In_1307,In_381);
xnor U2067 (N_2067,In_1063,In_1403);
xor U2068 (N_2068,In_1056,In_1093);
nor U2069 (N_2069,In_417,In_451);
xor U2070 (N_2070,In_57,In_217);
and U2071 (N_2071,In_1223,In_938);
xnor U2072 (N_2072,In_133,In_586);
nand U2073 (N_2073,In_207,In_619);
nor U2074 (N_2074,In_1371,In_1287);
nand U2075 (N_2075,In_945,In_972);
and U2076 (N_2076,In_96,In_1419);
xor U2077 (N_2077,In_417,In_454);
and U2078 (N_2078,In_891,In_250);
nand U2079 (N_2079,In_593,In_213);
or U2080 (N_2080,In_294,In_1348);
or U2081 (N_2081,In_319,In_1466);
xnor U2082 (N_2082,In_885,In_235);
xor U2083 (N_2083,In_604,In_1217);
or U2084 (N_2084,In_446,In_195);
xnor U2085 (N_2085,In_935,In_1001);
or U2086 (N_2086,In_1029,In_825);
xnor U2087 (N_2087,In_567,In_821);
xor U2088 (N_2088,In_1116,In_32);
and U2089 (N_2089,In_1351,In_883);
nand U2090 (N_2090,In_864,In_995);
nand U2091 (N_2091,In_34,In_1222);
nand U2092 (N_2092,In_506,In_1457);
or U2093 (N_2093,In_1259,In_23);
or U2094 (N_2094,In_665,In_1228);
nand U2095 (N_2095,In_64,In_1243);
or U2096 (N_2096,In_274,In_1499);
or U2097 (N_2097,In_1091,In_276);
and U2098 (N_2098,In_1429,In_1054);
or U2099 (N_2099,In_199,In_264);
or U2100 (N_2100,In_609,In_982);
and U2101 (N_2101,In_515,In_112);
nand U2102 (N_2102,In_359,In_1169);
nor U2103 (N_2103,In_403,In_1288);
nand U2104 (N_2104,In_1038,In_1190);
xnor U2105 (N_2105,In_746,In_1136);
nand U2106 (N_2106,In_1343,In_975);
or U2107 (N_2107,In_1362,In_580);
and U2108 (N_2108,In_350,In_1159);
nor U2109 (N_2109,In_1325,In_1465);
nand U2110 (N_2110,In_530,In_1136);
xnor U2111 (N_2111,In_90,In_878);
and U2112 (N_2112,In_560,In_1385);
or U2113 (N_2113,In_1100,In_1206);
nor U2114 (N_2114,In_789,In_1476);
nand U2115 (N_2115,In_751,In_2);
nor U2116 (N_2116,In_593,In_581);
nor U2117 (N_2117,In_356,In_306);
or U2118 (N_2118,In_640,In_706);
and U2119 (N_2119,In_525,In_1083);
nand U2120 (N_2120,In_1000,In_935);
xnor U2121 (N_2121,In_1146,In_934);
or U2122 (N_2122,In_1312,In_1004);
or U2123 (N_2123,In_596,In_1308);
nor U2124 (N_2124,In_1228,In_1441);
and U2125 (N_2125,In_173,In_167);
and U2126 (N_2126,In_282,In_103);
nor U2127 (N_2127,In_1014,In_1184);
nor U2128 (N_2128,In_1131,In_75);
and U2129 (N_2129,In_916,In_465);
and U2130 (N_2130,In_439,In_317);
and U2131 (N_2131,In_1059,In_1437);
nand U2132 (N_2132,In_1001,In_947);
or U2133 (N_2133,In_363,In_61);
or U2134 (N_2134,In_736,In_213);
xnor U2135 (N_2135,In_1320,In_1090);
nor U2136 (N_2136,In_1165,In_1372);
xor U2137 (N_2137,In_472,In_720);
nor U2138 (N_2138,In_529,In_276);
xnor U2139 (N_2139,In_1122,In_175);
or U2140 (N_2140,In_470,In_1446);
and U2141 (N_2141,In_1134,In_1004);
nand U2142 (N_2142,In_1497,In_362);
xnor U2143 (N_2143,In_217,In_1453);
nand U2144 (N_2144,In_1381,In_273);
and U2145 (N_2145,In_908,In_1072);
nand U2146 (N_2146,In_979,In_335);
nand U2147 (N_2147,In_205,In_1273);
nor U2148 (N_2148,In_359,In_538);
nand U2149 (N_2149,In_167,In_9);
and U2150 (N_2150,In_1277,In_987);
and U2151 (N_2151,In_1178,In_442);
xor U2152 (N_2152,In_324,In_102);
or U2153 (N_2153,In_1287,In_208);
and U2154 (N_2154,In_1456,In_849);
nand U2155 (N_2155,In_325,In_1172);
and U2156 (N_2156,In_428,In_828);
xnor U2157 (N_2157,In_61,In_469);
xnor U2158 (N_2158,In_1192,In_832);
nand U2159 (N_2159,In_1470,In_98);
or U2160 (N_2160,In_360,In_1009);
xor U2161 (N_2161,In_583,In_1487);
nand U2162 (N_2162,In_67,In_1237);
nor U2163 (N_2163,In_956,In_1386);
nor U2164 (N_2164,In_772,In_1071);
and U2165 (N_2165,In_250,In_1309);
xnor U2166 (N_2166,In_56,In_1245);
or U2167 (N_2167,In_204,In_1149);
or U2168 (N_2168,In_1133,In_933);
and U2169 (N_2169,In_288,In_1032);
or U2170 (N_2170,In_239,In_958);
or U2171 (N_2171,In_235,In_419);
nand U2172 (N_2172,In_213,In_461);
or U2173 (N_2173,In_1024,In_249);
or U2174 (N_2174,In_1280,In_1250);
nor U2175 (N_2175,In_218,In_40);
xnor U2176 (N_2176,In_1153,In_876);
nand U2177 (N_2177,In_1115,In_891);
nor U2178 (N_2178,In_400,In_614);
nor U2179 (N_2179,In_234,In_99);
nor U2180 (N_2180,In_135,In_1477);
xor U2181 (N_2181,In_110,In_352);
nand U2182 (N_2182,In_956,In_751);
or U2183 (N_2183,In_208,In_800);
nand U2184 (N_2184,In_407,In_1079);
nor U2185 (N_2185,In_546,In_415);
nor U2186 (N_2186,In_67,In_572);
and U2187 (N_2187,In_1208,In_876);
and U2188 (N_2188,In_119,In_723);
or U2189 (N_2189,In_1211,In_837);
nand U2190 (N_2190,In_965,In_226);
xnor U2191 (N_2191,In_1032,In_1099);
nand U2192 (N_2192,In_1078,In_973);
nor U2193 (N_2193,In_904,In_370);
nand U2194 (N_2194,In_244,In_314);
nand U2195 (N_2195,In_1396,In_560);
xor U2196 (N_2196,In_144,In_1048);
or U2197 (N_2197,In_513,In_845);
xor U2198 (N_2198,In_1270,In_551);
and U2199 (N_2199,In_49,In_1298);
or U2200 (N_2200,In_1423,In_852);
nor U2201 (N_2201,In_904,In_176);
and U2202 (N_2202,In_833,In_1341);
or U2203 (N_2203,In_354,In_440);
xor U2204 (N_2204,In_643,In_1476);
and U2205 (N_2205,In_346,In_794);
or U2206 (N_2206,In_671,In_718);
xnor U2207 (N_2207,In_1285,In_743);
nor U2208 (N_2208,In_917,In_1433);
nand U2209 (N_2209,In_687,In_1476);
or U2210 (N_2210,In_839,In_612);
and U2211 (N_2211,In_1364,In_1029);
xnor U2212 (N_2212,In_84,In_548);
xnor U2213 (N_2213,In_164,In_1126);
nand U2214 (N_2214,In_567,In_79);
xnor U2215 (N_2215,In_1409,In_642);
and U2216 (N_2216,In_194,In_28);
nor U2217 (N_2217,In_971,In_464);
and U2218 (N_2218,In_1286,In_56);
xor U2219 (N_2219,In_1005,In_582);
and U2220 (N_2220,In_345,In_664);
nor U2221 (N_2221,In_580,In_129);
or U2222 (N_2222,In_1112,In_137);
or U2223 (N_2223,In_1272,In_349);
nor U2224 (N_2224,In_135,In_1454);
or U2225 (N_2225,In_1281,In_813);
or U2226 (N_2226,In_1249,In_60);
and U2227 (N_2227,In_613,In_294);
and U2228 (N_2228,In_13,In_1227);
xor U2229 (N_2229,In_1288,In_656);
or U2230 (N_2230,In_1169,In_916);
and U2231 (N_2231,In_803,In_1126);
nor U2232 (N_2232,In_120,In_497);
or U2233 (N_2233,In_1140,In_1168);
or U2234 (N_2234,In_469,In_882);
xor U2235 (N_2235,In_784,In_625);
xor U2236 (N_2236,In_399,In_369);
and U2237 (N_2237,In_181,In_512);
nand U2238 (N_2238,In_84,In_799);
and U2239 (N_2239,In_1080,In_1391);
and U2240 (N_2240,In_1473,In_1149);
or U2241 (N_2241,In_937,In_736);
nand U2242 (N_2242,In_463,In_490);
nand U2243 (N_2243,In_1035,In_660);
and U2244 (N_2244,In_340,In_1357);
xor U2245 (N_2245,In_440,In_819);
xnor U2246 (N_2246,In_414,In_1298);
and U2247 (N_2247,In_976,In_620);
and U2248 (N_2248,In_1459,In_1099);
and U2249 (N_2249,In_1242,In_1388);
or U2250 (N_2250,In_247,In_774);
nand U2251 (N_2251,In_272,In_56);
xnor U2252 (N_2252,In_870,In_117);
nor U2253 (N_2253,In_686,In_465);
and U2254 (N_2254,In_821,In_282);
xnor U2255 (N_2255,In_24,In_136);
xnor U2256 (N_2256,In_1134,In_697);
or U2257 (N_2257,In_1302,In_1339);
or U2258 (N_2258,In_250,In_735);
nor U2259 (N_2259,In_409,In_448);
and U2260 (N_2260,In_718,In_1126);
nand U2261 (N_2261,In_836,In_312);
or U2262 (N_2262,In_839,In_868);
or U2263 (N_2263,In_857,In_984);
xnor U2264 (N_2264,In_1298,In_978);
or U2265 (N_2265,In_1278,In_443);
or U2266 (N_2266,In_1281,In_162);
and U2267 (N_2267,In_919,In_1429);
and U2268 (N_2268,In_744,In_321);
and U2269 (N_2269,In_582,In_182);
or U2270 (N_2270,In_70,In_233);
nand U2271 (N_2271,In_679,In_769);
and U2272 (N_2272,In_1415,In_8);
or U2273 (N_2273,In_524,In_1187);
or U2274 (N_2274,In_1422,In_169);
nand U2275 (N_2275,In_1240,In_794);
or U2276 (N_2276,In_144,In_1164);
or U2277 (N_2277,In_1124,In_1458);
nand U2278 (N_2278,In_411,In_625);
xor U2279 (N_2279,In_1393,In_853);
xor U2280 (N_2280,In_1117,In_1421);
or U2281 (N_2281,In_1048,In_811);
or U2282 (N_2282,In_644,In_296);
xor U2283 (N_2283,In_797,In_1054);
nand U2284 (N_2284,In_769,In_822);
xnor U2285 (N_2285,In_1323,In_1133);
nor U2286 (N_2286,In_791,In_837);
nor U2287 (N_2287,In_1334,In_592);
and U2288 (N_2288,In_468,In_1045);
or U2289 (N_2289,In_719,In_559);
nor U2290 (N_2290,In_705,In_362);
nand U2291 (N_2291,In_65,In_281);
nand U2292 (N_2292,In_1003,In_1247);
and U2293 (N_2293,In_550,In_140);
or U2294 (N_2294,In_1352,In_461);
xnor U2295 (N_2295,In_839,In_1381);
and U2296 (N_2296,In_148,In_993);
xor U2297 (N_2297,In_1149,In_342);
nor U2298 (N_2298,In_935,In_1152);
nor U2299 (N_2299,In_1488,In_28);
and U2300 (N_2300,In_338,In_454);
nor U2301 (N_2301,In_549,In_31);
or U2302 (N_2302,In_841,In_178);
nand U2303 (N_2303,In_794,In_493);
or U2304 (N_2304,In_1127,In_1306);
xnor U2305 (N_2305,In_1324,In_386);
or U2306 (N_2306,In_1251,In_1003);
nor U2307 (N_2307,In_27,In_1421);
or U2308 (N_2308,In_1116,In_631);
nor U2309 (N_2309,In_1011,In_1345);
xnor U2310 (N_2310,In_1108,In_1310);
nand U2311 (N_2311,In_581,In_619);
nand U2312 (N_2312,In_1434,In_470);
and U2313 (N_2313,In_560,In_607);
or U2314 (N_2314,In_389,In_915);
and U2315 (N_2315,In_973,In_354);
nand U2316 (N_2316,In_102,In_468);
and U2317 (N_2317,In_1198,In_310);
and U2318 (N_2318,In_390,In_1210);
or U2319 (N_2319,In_144,In_1032);
nor U2320 (N_2320,In_864,In_1345);
xnor U2321 (N_2321,In_265,In_111);
or U2322 (N_2322,In_1162,In_775);
or U2323 (N_2323,In_430,In_1076);
xor U2324 (N_2324,In_1366,In_711);
or U2325 (N_2325,In_169,In_990);
and U2326 (N_2326,In_703,In_1122);
xnor U2327 (N_2327,In_721,In_1264);
and U2328 (N_2328,In_715,In_1367);
nor U2329 (N_2329,In_690,In_900);
or U2330 (N_2330,In_1158,In_444);
nand U2331 (N_2331,In_1443,In_533);
nand U2332 (N_2332,In_1020,In_1172);
nor U2333 (N_2333,In_26,In_365);
or U2334 (N_2334,In_875,In_598);
nand U2335 (N_2335,In_987,In_876);
nand U2336 (N_2336,In_391,In_1431);
xnor U2337 (N_2337,In_245,In_794);
or U2338 (N_2338,In_1344,In_1444);
xor U2339 (N_2339,In_187,In_590);
nor U2340 (N_2340,In_274,In_320);
xnor U2341 (N_2341,In_513,In_443);
xnor U2342 (N_2342,In_98,In_867);
nand U2343 (N_2343,In_883,In_601);
and U2344 (N_2344,In_252,In_808);
and U2345 (N_2345,In_1335,In_16);
nand U2346 (N_2346,In_1194,In_562);
nand U2347 (N_2347,In_436,In_223);
or U2348 (N_2348,In_1126,In_54);
xnor U2349 (N_2349,In_1274,In_1459);
xnor U2350 (N_2350,In_561,In_1382);
or U2351 (N_2351,In_958,In_1087);
or U2352 (N_2352,In_357,In_77);
nand U2353 (N_2353,In_1232,In_426);
nor U2354 (N_2354,In_717,In_739);
nand U2355 (N_2355,In_1114,In_349);
or U2356 (N_2356,In_225,In_367);
nand U2357 (N_2357,In_1053,In_436);
or U2358 (N_2358,In_974,In_1330);
and U2359 (N_2359,In_1132,In_352);
nand U2360 (N_2360,In_561,In_1256);
nand U2361 (N_2361,In_554,In_522);
xnor U2362 (N_2362,In_116,In_664);
nand U2363 (N_2363,In_573,In_365);
and U2364 (N_2364,In_1078,In_271);
or U2365 (N_2365,In_648,In_197);
nor U2366 (N_2366,In_780,In_1365);
and U2367 (N_2367,In_1092,In_829);
and U2368 (N_2368,In_1428,In_1298);
and U2369 (N_2369,In_586,In_269);
and U2370 (N_2370,In_978,In_968);
or U2371 (N_2371,In_236,In_352);
xor U2372 (N_2372,In_1441,In_832);
nand U2373 (N_2373,In_1378,In_745);
or U2374 (N_2374,In_1394,In_216);
nand U2375 (N_2375,In_1104,In_428);
nor U2376 (N_2376,In_1210,In_335);
nand U2377 (N_2377,In_30,In_789);
and U2378 (N_2378,In_648,In_928);
xnor U2379 (N_2379,In_823,In_1462);
or U2380 (N_2380,In_1208,In_260);
nor U2381 (N_2381,In_774,In_300);
nand U2382 (N_2382,In_588,In_1470);
and U2383 (N_2383,In_507,In_358);
nand U2384 (N_2384,In_775,In_1091);
and U2385 (N_2385,In_109,In_709);
nor U2386 (N_2386,In_1066,In_1085);
or U2387 (N_2387,In_388,In_436);
xnor U2388 (N_2388,In_784,In_292);
nand U2389 (N_2389,In_694,In_311);
or U2390 (N_2390,In_850,In_804);
nand U2391 (N_2391,In_21,In_1498);
nand U2392 (N_2392,In_262,In_555);
nand U2393 (N_2393,In_982,In_385);
and U2394 (N_2394,In_429,In_1263);
xnor U2395 (N_2395,In_599,In_1076);
and U2396 (N_2396,In_106,In_179);
nor U2397 (N_2397,In_1423,In_730);
and U2398 (N_2398,In_879,In_338);
or U2399 (N_2399,In_951,In_594);
or U2400 (N_2400,In_1328,In_540);
nor U2401 (N_2401,In_559,In_1116);
nand U2402 (N_2402,In_873,In_1399);
and U2403 (N_2403,In_320,In_543);
nor U2404 (N_2404,In_1384,In_1352);
nand U2405 (N_2405,In_649,In_952);
nor U2406 (N_2406,In_759,In_542);
nor U2407 (N_2407,In_1493,In_988);
or U2408 (N_2408,In_652,In_25);
xnor U2409 (N_2409,In_721,In_1378);
xnor U2410 (N_2410,In_1121,In_498);
and U2411 (N_2411,In_120,In_1165);
and U2412 (N_2412,In_481,In_310);
nor U2413 (N_2413,In_324,In_658);
nor U2414 (N_2414,In_600,In_471);
xnor U2415 (N_2415,In_272,In_772);
or U2416 (N_2416,In_1338,In_1103);
nand U2417 (N_2417,In_470,In_1326);
nor U2418 (N_2418,In_890,In_893);
xnor U2419 (N_2419,In_1004,In_205);
xor U2420 (N_2420,In_1187,In_724);
xor U2421 (N_2421,In_647,In_1257);
nor U2422 (N_2422,In_1263,In_847);
nor U2423 (N_2423,In_87,In_1171);
nand U2424 (N_2424,In_629,In_886);
xor U2425 (N_2425,In_1297,In_1332);
xnor U2426 (N_2426,In_525,In_965);
or U2427 (N_2427,In_18,In_336);
or U2428 (N_2428,In_844,In_1118);
nand U2429 (N_2429,In_392,In_1121);
or U2430 (N_2430,In_1248,In_704);
nand U2431 (N_2431,In_935,In_631);
or U2432 (N_2432,In_1228,In_623);
xor U2433 (N_2433,In_788,In_889);
nand U2434 (N_2434,In_1348,In_1013);
or U2435 (N_2435,In_658,In_578);
nor U2436 (N_2436,In_1006,In_653);
nor U2437 (N_2437,In_24,In_614);
and U2438 (N_2438,In_1349,In_340);
nand U2439 (N_2439,In_1036,In_570);
or U2440 (N_2440,In_2,In_1459);
xnor U2441 (N_2441,In_1489,In_742);
nand U2442 (N_2442,In_163,In_762);
xor U2443 (N_2443,In_301,In_681);
or U2444 (N_2444,In_1235,In_1260);
and U2445 (N_2445,In_741,In_257);
nor U2446 (N_2446,In_1190,In_1050);
nand U2447 (N_2447,In_377,In_977);
and U2448 (N_2448,In_614,In_636);
nor U2449 (N_2449,In_1227,In_1058);
or U2450 (N_2450,In_457,In_800);
nand U2451 (N_2451,In_690,In_468);
xnor U2452 (N_2452,In_1223,In_787);
nor U2453 (N_2453,In_1396,In_448);
nor U2454 (N_2454,In_166,In_1423);
and U2455 (N_2455,In_416,In_282);
xor U2456 (N_2456,In_858,In_1098);
nor U2457 (N_2457,In_371,In_62);
and U2458 (N_2458,In_94,In_177);
or U2459 (N_2459,In_715,In_908);
nand U2460 (N_2460,In_1142,In_1440);
nor U2461 (N_2461,In_171,In_638);
nor U2462 (N_2462,In_526,In_987);
nand U2463 (N_2463,In_1334,In_414);
nand U2464 (N_2464,In_293,In_243);
and U2465 (N_2465,In_1034,In_1013);
or U2466 (N_2466,In_877,In_100);
and U2467 (N_2467,In_663,In_655);
nor U2468 (N_2468,In_1105,In_1029);
nand U2469 (N_2469,In_365,In_61);
xnor U2470 (N_2470,In_139,In_1190);
or U2471 (N_2471,In_921,In_1284);
xor U2472 (N_2472,In_135,In_212);
nand U2473 (N_2473,In_1155,In_1166);
xor U2474 (N_2474,In_1181,In_619);
or U2475 (N_2475,In_1138,In_553);
and U2476 (N_2476,In_256,In_576);
and U2477 (N_2477,In_374,In_498);
nor U2478 (N_2478,In_836,In_736);
or U2479 (N_2479,In_67,In_920);
and U2480 (N_2480,In_880,In_1465);
and U2481 (N_2481,In_603,In_1428);
nor U2482 (N_2482,In_861,In_663);
or U2483 (N_2483,In_1149,In_678);
xnor U2484 (N_2484,In_9,In_1052);
xor U2485 (N_2485,In_1268,In_300);
or U2486 (N_2486,In_1006,In_260);
nor U2487 (N_2487,In_895,In_1299);
or U2488 (N_2488,In_576,In_76);
or U2489 (N_2489,In_817,In_650);
nor U2490 (N_2490,In_1395,In_150);
nor U2491 (N_2491,In_753,In_477);
nand U2492 (N_2492,In_510,In_229);
or U2493 (N_2493,In_811,In_1304);
or U2494 (N_2494,In_191,In_24);
nor U2495 (N_2495,In_547,In_905);
nor U2496 (N_2496,In_282,In_644);
nor U2497 (N_2497,In_1473,In_395);
xor U2498 (N_2498,In_286,In_55);
or U2499 (N_2499,In_1378,In_660);
and U2500 (N_2500,In_591,In_1437);
and U2501 (N_2501,In_468,In_972);
nand U2502 (N_2502,In_957,In_202);
and U2503 (N_2503,In_233,In_393);
and U2504 (N_2504,In_1328,In_1189);
nand U2505 (N_2505,In_1365,In_573);
nand U2506 (N_2506,In_1296,In_692);
nor U2507 (N_2507,In_582,In_1026);
xnor U2508 (N_2508,In_160,In_1409);
xnor U2509 (N_2509,In_930,In_636);
and U2510 (N_2510,In_298,In_1169);
or U2511 (N_2511,In_804,In_510);
and U2512 (N_2512,In_1137,In_338);
or U2513 (N_2513,In_599,In_1161);
xnor U2514 (N_2514,In_711,In_311);
nand U2515 (N_2515,In_1124,In_832);
or U2516 (N_2516,In_924,In_541);
and U2517 (N_2517,In_133,In_473);
nor U2518 (N_2518,In_197,In_329);
and U2519 (N_2519,In_1442,In_222);
nor U2520 (N_2520,In_855,In_592);
nand U2521 (N_2521,In_579,In_199);
xor U2522 (N_2522,In_461,In_991);
and U2523 (N_2523,In_881,In_854);
xor U2524 (N_2524,In_972,In_1208);
xor U2525 (N_2525,In_459,In_1141);
nand U2526 (N_2526,In_944,In_972);
nand U2527 (N_2527,In_4,In_772);
nand U2528 (N_2528,In_396,In_16);
or U2529 (N_2529,In_598,In_1158);
nand U2530 (N_2530,In_811,In_153);
nor U2531 (N_2531,In_162,In_598);
or U2532 (N_2532,In_247,In_982);
and U2533 (N_2533,In_460,In_565);
or U2534 (N_2534,In_1421,In_637);
xor U2535 (N_2535,In_885,In_1374);
xor U2536 (N_2536,In_396,In_783);
nand U2537 (N_2537,In_683,In_398);
nand U2538 (N_2538,In_994,In_232);
nand U2539 (N_2539,In_776,In_134);
nand U2540 (N_2540,In_1189,In_132);
or U2541 (N_2541,In_596,In_951);
or U2542 (N_2542,In_737,In_1154);
xor U2543 (N_2543,In_588,In_668);
nand U2544 (N_2544,In_1459,In_601);
nand U2545 (N_2545,In_152,In_1090);
nand U2546 (N_2546,In_1032,In_346);
nor U2547 (N_2547,In_650,In_1267);
nand U2548 (N_2548,In_991,In_518);
nand U2549 (N_2549,In_1165,In_268);
and U2550 (N_2550,In_255,In_133);
or U2551 (N_2551,In_1093,In_911);
xor U2552 (N_2552,In_1301,In_328);
nand U2553 (N_2553,In_624,In_634);
xnor U2554 (N_2554,In_288,In_1157);
and U2555 (N_2555,In_989,In_689);
nand U2556 (N_2556,In_980,In_1418);
nand U2557 (N_2557,In_1050,In_1055);
nand U2558 (N_2558,In_168,In_229);
or U2559 (N_2559,In_248,In_1499);
nor U2560 (N_2560,In_894,In_604);
xnor U2561 (N_2561,In_1457,In_263);
xnor U2562 (N_2562,In_1153,In_1187);
nor U2563 (N_2563,In_587,In_1022);
nand U2564 (N_2564,In_421,In_1264);
nand U2565 (N_2565,In_634,In_140);
and U2566 (N_2566,In_368,In_30);
and U2567 (N_2567,In_597,In_1493);
nand U2568 (N_2568,In_143,In_946);
nor U2569 (N_2569,In_621,In_157);
or U2570 (N_2570,In_579,In_778);
nor U2571 (N_2571,In_417,In_511);
or U2572 (N_2572,In_300,In_107);
and U2573 (N_2573,In_228,In_331);
nor U2574 (N_2574,In_6,In_488);
and U2575 (N_2575,In_1007,In_893);
xor U2576 (N_2576,In_743,In_767);
nor U2577 (N_2577,In_1250,In_183);
nor U2578 (N_2578,In_474,In_1403);
or U2579 (N_2579,In_736,In_614);
nand U2580 (N_2580,In_1272,In_704);
and U2581 (N_2581,In_813,In_352);
xnor U2582 (N_2582,In_954,In_501);
or U2583 (N_2583,In_1142,In_626);
or U2584 (N_2584,In_983,In_1370);
xnor U2585 (N_2585,In_1086,In_961);
nand U2586 (N_2586,In_1349,In_55);
nand U2587 (N_2587,In_443,In_667);
nand U2588 (N_2588,In_1270,In_362);
xor U2589 (N_2589,In_505,In_372);
xnor U2590 (N_2590,In_210,In_1221);
or U2591 (N_2591,In_1320,In_839);
xor U2592 (N_2592,In_308,In_418);
nor U2593 (N_2593,In_765,In_647);
nor U2594 (N_2594,In_249,In_1473);
nand U2595 (N_2595,In_211,In_956);
or U2596 (N_2596,In_960,In_846);
or U2597 (N_2597,In_1257,In_748);
and U2598 (N_2598,In_1171,In_85);
or U2599 (N_2599,In_241,In_703);
xor U2600 (N_2600,In_975,In_540);
or U2601 (N_2601,In_945,In_1271);
nand U2602 (N_2602,In_929,In_1084);
xnor U2603 (N_2603,In_1167,In_1446);
or U2604 (N_2604,In_559,In_1454);
and U2605 (N_2605,In_1252,In_1040);
and U2606 (N_2606,In_843,In_1201);
and U2607 (N_2607,In_1287,In_1314);
and U2608 (N_2608,In_1320,In_1472);
nor U2609 (N_2609,In_502,In_629);
nor U2610 (N_2610,In_1324,In_271);
nand U2611 (N_2611,In_1247,In_161);
nor U2612 (N_2612,In_1369,In_1038);
nor U2613 (N_2613,In_1081,In_703);
nor U2614 (N_2614,In_1347,In_640);
nand U2615 (N_2615,In_834,In_961);
nand U2616 (N_2616,In_697,In_449);
nor U2617 (N_2617,In_1372,In_757);
xnor U2618 (N_2618,In_566,In_766);
or U2619 (N_2619,In_1459,In_332);
and U2620 (N_2620,In_1393,In_14);
nor U2621 (N_2621,In_67,In_691);
nor U2622 (N_2622,In_216,In_1445);
and U2623 (N_2623,In_1410,In_709);
nand U2624 (N_2624,In_232,In_896);
and U2625 (N_2625,In_581,In_1247);
or U2626 (N_2626,In_698,In_858);
xnor U2627 (N_2627,In_1358,In_139);
and U2628 (N_2628,In_248,In_968);
nand U2629 (N_2629,In_190,In_1271);
or U2630 (N_2630,In_63,In_1475);
and U2631 (N_2631,In_505,In_1458);
xor U2632 (N_2632,In_969,In_1113);
and U2633 (N_2633,In_1110,In_142);
nor U2634 (N_2634,In_630,In_1024);
and U2635 (N_2635,In_233,In_1331);
and U2636 (N_2636,In_870,In_1266);
nor U2637 (N_2637,In_1212,In_340);
nor U2638 (N_2638,In_1378,In_48);
and U2639 (N_2639,In_832,In_1464);
nor U2640 (N_2640,In_1179,In_172);
nand U2641 (N_2641,In_1363,In_180);
xor U2642 (N_2642,In_462,In_331);
and U2643 (N_2643,In_344,In_746);
or U2644 (N_2644,In_325,In_467);
and U2645 (N_2645,In_632,In_548);
nand U2646 (N_2646,In_762,In_35);
nor U2647 (N_2647,In_245,In_422);
nand U2648 (N_2648,In_1152,In_746);
and U2649 (N_2649,In_189,In_1116);
xor U2650 (N_2650,In_1326,In_374);
nand U2651 (N_2651,In_864,In_729);
or U2652 (N_2652,In_1093,In_1343);
and U2653 (N_2653,In_598,In_954);
nand U2654 (N_2654,In_1032,In_1201);
and U2655 (N_2655,In_1004,In_472);
nand U2656 (N_2656,In_1226,In_1383);
or U2657 (N_2657,In_1152,In_547);
and U2658 (N_2658,In_550,In_608);
or U2659 (N_2659,In_1416,In_886);
or U2660 (N_2660,In_199,In_1190);
nor U2661 (N_2661,In_652,In_1434);
and U2662 (N_2662,In_1228,In_192);
nor U2663 (N_2663,In_674,In_396);
and U2664 (N_2664,In_745,In_500);
or U2665 (N_2665,In_284,In_1034);
and U2666 (N_2666,In_399,In_599);
and U2667 (N_2667,In_277,In_1349);
nor U2668 (N_2668,In_69,In_1084);
or U2669 (N_2669,In_52,In_685);
nor U2670 (N_2670,In_136,In_1351);
nor U2671 (N_2671,In_1492,In_710);
xor U2672 (N_2672,In_1143,In_230);
nor U2673 (N_2673,In_225,In_818);
xor U2674 (N_2674,In_1126,In_1046);
nor U2675 (N_2675,In_712,In_379);
and U2676 (N_2676,In_1036,In_1032);
xnor U2677 (N_2677,In_565,In_357);
and U2678 (N_2678,In_42,In_143);
nor U2679 (N_2679,In_569,In_685);
nor U2680 (N_2680,In_128,In_325);
xnor U2681 (N_2681,In_1431,In_509);
or U2682 (N_2682,In_76,In_739);
nor U2683 (N_2683,In_711,In_730);
nor U2684 (N_2684,In_590,In_66);
nor U2685 (N_2685,In_501,In_1096);
nand U2686 (N_2686,In_1147,In_782);
nand U2687 (N_2687,In_999,In_1258);
nor U2688 (N_2688,In_395,In_282);
nor U2689 (N_2689,In_1403,In_1110);
nor U2690 (N_2690,In_1294,In_1314);
and U2691 (N_2691,In_115,In_323);
and U2692 (N_2692,In_502,In_1010);
nor U2693 (N_2693,In_141,In_967);
nor U2694 (N_2694,In_618,In_7);
xor U2695 (N_2695,In_138,In_513);
xor U2696 (N_2696,In_1077,In_359);
and U2697 (N_2697,In_1236,In_447);
nand U2698 (N_2698,In_724,In_592);
nand U2699 (N_2699,In_1081,In_32);
nor U2700 (N_2700,In_401,In_96);
and U2701 (N_2701,In_528,In_1110);
nor U2702 (N_2702,In_595,In_1098);
or U2703 (N_2703,In_493,In_1135);
or U2704 (N_2704,In_955,In_1418);
nand U2705 (N_2705,In_514,In_1240);
nand U2706 (N_2706,In_576,In_1417);
nand U2707 (N_2707,In_1345,In_278);
nor U2708 (N_2708,In_879,In_1486);
nor U2709 (N_2709,In_1463,In_198);
xnor U2710 (N_2710,In_1412,In_1480);
nand U2711 (N_2711,In_41,In_485);
nor U2712 (N_2712,In_1060,In_1431);
or U2713 (N_2713,In_1257,In_217);
or U2714 (N_2714,In_498,In_652);
nand U2715 (N_2715,In_1094,In_1108);
or U2716 (N_2716,In_455,In_601);
xnor U2717 (N_2717,In_480,In_915);
nand U2718 (N_2718,In_515,In_1029);
nand U2719 (N_2719,In_335,In_634);
xnor U2720 (N_2720,In_917,In_973);
nand U2721 (N_2721,In_488,In_531);
and U2722 (N_2722,In_131,In_974);
and U2723 (N_2723,In_1047,In_1406);
nor U2724 (N_2724,In_210,In_1375);
or U2725 (N_2725,In_1347,In_1363);
or U2726 (N_2726,In_30,In_154);
nor U2727 (N_2727,In_888,In_1040);
nand U2728 (N_2728,In_995,In_1113);
or U2729 (N_2729,In_1324,In_1011);
and U2730 (N_2730,In_400,In_867);
nor U2731 (N_2731,In_128,In_1106);
nor U2732 (N_2732,In_1310,In_657);
and U2733 (N_2733,In_722,In_1414);
xor U2734 (N_2734,In_120,In_253);
or U2735 (N_2735,In_793,In_1112);
and U2736 (N_2736,In_1201,In_128);
xor U2737 (N_2737,In_664,In_106);
or U2738 (N_2738,In_1072,In_1411);
nand U2739 (N_2739,In_1308,In_672);
nand U2740 (N_2740,In_638,In_270);
or U2741 (N_2741,In_531,In_20);
nand U2742 (N_2742,In_949,In_412);
or U2743 (N_2743,In_207,In_1280);
xnor U2744 (N_2744,In_133,In_1157);
or U2745 (N_2745,In_137,In_1369);
xnor U2746 (N_2746,In_1347,In_406);
and U2747 (N_2747,In_175,In_625);
nor U2748 (N_2748,In_130,In_17);
or U2749 (N_2749,In_1341,In_1263);
or U2750 (N_2750,In_1397,In_486);
nor U2751 (N_2751,In_1006,In_644);
nand U2752 (N_2752,In_1082,In_1066);
xor U2753 (N_2753,In_1200,In_1271);
and U2754 (N_2754,In_1373,In_1217);
nand U2755 (N_2755,In_108,In_1051);
and U2756 (N_2756,In_1275,In_1178);
or U2757 (N_2757,In_837,In_1100);
nor U2758 (N_2758,In_1170,In_1182);
or U2759 (N_2759,In_973,In_395);
xor U2760 (N_2760,In_283,In_610);
xor U2761 (N_2761,In_647,In_1383);
and U2762 (N_2762,In_271,In_997);
and U2763 (N_2763,In_1395,In_151);
and U2764 (N_2764,In_716,In_47);
nor U2765 (N_2765,In_338,In_773);
or U2766 (N_2766,In_1459,In_915);
nor U2767 (N_2767,In_527,In_237);
xor U2768 (N_2768,In_181,In_712);
or U2769 (N_2769,In_1478,In_1251);
or U2770 (N_2770,In_1453,In_1130);
and U2771 (N_2771,In_318,In_707);
and U2772 (N_2772,In_1074,In_326);
nor U2773 (N_2773,In_1167,In_1479);
xnor U2774 (N_2774,In_1453,In_761);
and U2775 (N_2775,In_74,In_1279);
nor U2776 (N_2776,In_1483,In_238);
xnor U2777 (N_2777,In_144,In_595);
nand U2778 (N_2778,In_1411,In_160);
nor U2779 (N_2779,In_485,In_1358);
or U2780 (N_2780,In_1202,In_1414);
nor U2781 (N_2781,In_492,In_1437);
nor U2782 (N_2782,In_951,In_434);
and U2783 (N_2783,In_666,In_318);
nand U2784 (N_2784,In_1386,In_1106);
or U2785 (N_2785,In_941,In_1160);
xor U2786 (N_2786,In_1003,In_106);
and U2787 (N_2787,In_1084,In_1219);
and U2788 (N_2788,In_545,In_77);
nand U2789 (N_2789,In_351,In_822);
nor U2790 (N_2790,In_718,In_1131);
or U2791 (N_2791,In_811,In_1126);
nor U2792 (N_2792,In_1442,In_94);
xor U2793 (N_2793,In_462,In_503);
xor U2794 (N_2794,In_892,In_1372);
nand U2795 (N_2795,In_312,In_1211);
xnor U2796 (N_2796,In_653,In_1191);
nand U2797 (N_2797,In_608,In_592);
or U2798 (N_2798,In_330,In_226);
nor U2799 (N_2799,In_1175,In_363);
and U2800 (N_2800,In_868,In_939);
xnor U2801 (N_2801,In_1134,In_1290);
nor U2802 (N_2802,In_346,In_1330);
xnor U2803 (N_2803,In_928,In_1410);
or U2804 (N_2804,In_1467,In_98);
nor U2805 (N_2805,In_392,In_943);
nand U2806 (N_2806,In_1062,In_1058);
nand U2807 (N_2807,In_800,In_398);
or U2808 (N_2808,In_278,In_1211);
nand U2809 (N_2809,In_345,In_692);
and U2810 (N_2810,In_1374,In_110);
or U2811 (N_2811,In_1356,In_1208);
or U2812 (N_2812,In_450,In_765);
nor U2813 (N_2813,In_1333,In_945);
nor U2814 (N_2814,In_872,In_1116);
nand U2815 (N_2815,In_1375,In_1097);
or U2816 (N_2816,In_469,In_889);
nor U2817 (N_2817,In_1237,In_1446);
and U2818 (N_2818,In_755,In_819);
or U2819 (N_2819,In_44,In_69);
or U2820 (N_2820,In_59,In_257);
xnor U2821 (N_2821,In_1197,In_894);
nor U2822 (N_2822,In_1409,In_613);
or U2823 (N_2823,In_1281,In_35);
or U2824 (N_2824,In_767,In_585);
nor U2825 (N_2825,In_80,In_1320);
or U2826 (N_2826,In_393,In_1124);
nor U2827 (N_2827,In_321,In_279);
nand U2828 (N_2828,In_1298,In_684);
nand U2829 (N_2829,In_747,In_859);
or U2830 (N_2830,In_1022,In_820);
and U2831 (N_2831,In_716,In_1020);
nor U2832 (N_2832,In_127,In_883);
nand U2833 (N_2833,In_341,In_884);
or U2834 (N_2834,In_835,In_1226);
and U2835 (N_2835,In_727,In_815);
nand U2836 (N_2836,In_951,In_431);
or U2837 (N_2837,In_736,In_361);
or U2838 (N_2838,In_606,In_227);
or U2839 (N_2839,In_60,In_1021);
nor U2840 (N_2840,In_786,In_1410);
and U2841 (N_2841,In_261,In_1266);
xor U2842 (N_2842,In_1151,In_1437);
xnor U2843 (N_2843,In_1350,In_1230);
xnor U2844 (N_2844,In_1472,In_410);
nand U2845 (N_2845,In_1131,In_1358);
nand U2846 (N_2846,In_474,In_761);
xnor U2847 (N_2847,In_332,In_1476);
and U2848 (N_2848,In_1042,In_303);
nor U2849 (N_2849,In_1403,In_1072);
and U2850 (N_2850,In_859,In_409);
xor U2851 (N_2851,In_119,In_1246);
or U2852 (N_2852,In_1421,In_215);
xnor U2853 (N_2853,In_292,In_1377);
nor U2854 (N_2854,In_1012,In_1215);
and U2855 (N_2855,In_559,In_943);
xor U2856 (N_2856,In_1493,In_47);
nand U2857 (N_2857,In_1255,In_131);
xnor U2858 (N_2858,In_18,In_1152);
nand U2859 (N_2859,In_1473,In_1443);
nor U2860 (N_2860,In_21,In_1371);
nand U2861 (N_2861,In_71,In_842);
or U2862 (N_2862,In_1495,In_1031);
nor U2863 (N_2863,In_1067,In_1073);
nor U2864 (N_2864,In_867,In_1386);
or U2865 (N_2865,In_1492,In_1282);
nor U2866 (N_2866,In_776,In_663);
and U2867 (N_2867,In_276,In_1343);
and U2868 (N_2868,In_497,In_1069);
nor U2869 (N_2869,In_1224,In_767);
and U2870 (N_2870,In_1070,In_793);
and U2871 (N_2871,In_872,In_315);
or U2872 (N_2872,In_809,In_1379);
nor U2873 (N_2873,In_484,In_883);
and U2874 (N_2874,In_231,In_210);
nand U2875 (N_2875,In_1462,In_342);
nor U2876 (N_2876,In_19,In_1292);
xnor U2877 (N_2877,In_983,In_1192);
or U2878 (N_2878,In_602,In_1024);
xor U2879 (N_2879,In_890,In_636);
or U2880 (N_2880,In_310,In_531);
nand U2881 (N_2881,In_1302,In_457);
nand U2882 (N_2882,In_590,In_1298);
nor U2883 (N_2883,In_470,In_1107);
nand U2884 (N_2884,In_778,In_1139);
nand U2885 (N_2885,In_914,In_1470);
xor U2886 (N_2886,In_329,In_68);
and U2887 (N_2887,In_224,In_1093);
or U2888 (N_2888,In_168,In_1360);
xor U2889 (N_2889,In_1373,In_404);
xor U2890 (N_2890,In_151,In_585);
nand U2891 (N_2891,In_200,In_1426);
and U2892 (N_2892,In_380,In_906);
xnor U2893 (N_2893,In_96,In_987);
and U2894 (N_2894,In_594,In_1261);
xnor U2895 (N_2895,In_244,In_477);
and U2896 (N_2896,In_856,In_236);
and U2897 (N_2897,In_99,In_762);
nor U2898 (N_2898,In_764,In_234);
and U2899 (N_2899,In_1462,In_746);
and U2900 (N_2900,In_31,In_467);
or U2901 (N_2901,In_349,In_1139);
xnor U2902 (N_2902,In_1162,In_1170);
nor U2903 (N_2903,In_78,In_1211);
nand U2904 (N_2904,In_992,In_399);
nor U2905 (N_2905,In_615,In_968);
nor U2906 (N_2906,In_67,In_741);
nand U2907 (N_2907,In_1369,In_1078);
nor U2908 (N_2908,In_246,In_670);
nand U2909 (N_2909,In_454,In_612);
or U2910 (N_2910,In_227,In_1354);
and U2911 (N_2911,In_365,In_206);
nor U2912 (N_2912,In_103,In_1082);
nor U2913 (N_2913,In_1002,In_1198);
or U2914 (N_2914,In_869,In_740);
nor U2915 (N_2915,In_781,In_516);
nor U2916 (N_2916,In_1265,In_1226);
nand U2917 (N_2917,In_892,In_926);
nor U2918 (N_2918,In_17,In_990);
or U2919 (N_2919,In_890,In_15);
xor U2920 (N_2920,In_90,In_378);
xor U2921 (N_2921,In_925,In_830);
xnor U2922 (N_2922,In_773,In_7);
and U2923 (N_2923,In_791,In_403);
or U2924 (N_2924,In_686,In_201);
nand U2925 (N_2925,In_856,In_1407);
xor U2926 (N_2926,In_469,In_548);
or U2927 (N_2927,In_375,In_185);
nor U2928 (N_2928,In_349,In_137);
and U2929 (N_2929,In_1290,In_642);
xnor U2930 (N_2930,In_1068,In_274);
nand U2931 (N_2931,In_1473,In_299);
xnor U2932 (N_2932,In_1416,In_658);
and U2933 (N_2933,In_1155,In_714);
nor U2934 (N_2934,In_1432,In_1181);
nor U2935 (N_2935,In_165,In_1030);
xor U2936 (N_2936,In_1086,In_323);
nand U2937 (N_2937,In_328,In_1258);
xor U2938 (N_2938,In_605,In_478);
or U2939 (N_2939,In_45,In_673);
nor U2940 (N_2940,In_343,In_306);
and U2941 (N_2941,In_954,In_1312);
xnor U2942 (N_2942,In_1301,In_1314);
xnor U2943 (N_2943,In_1373,In_753);
and U2944 (N_2944,In_979,In_621);
nor U2945 (N_2945,In_519,In_731);
nand U2946 (N_2946,In_217,In_985);
nor U2947 (N_2947,In_1353,In_1451);
and U2948 (N_2948,In_525,In_1269);
or U2949 (N_2949,In_171,In_52);
nor U2950 (N_2950,In_959,In_648);
and U2951 (N_2951,In_940,In_1485);
or U2952 (N_2952,In_1027,In_544);
xor U2953 (N_2953,In_350,In_479);
nor U2954 (N_2954,In_451,In_940);
nand U2955 (N_2955,In_294,In_379);
xnor U2956 (N_2956,In_862,In_1163);
nand U2957 (N_2957,In_206,In_776);
nand U2958 (N_2958,In_1272,In_1264);
and U2959 (N_2959,In_1284,In_723);
and U2960 (N_2960,In_546,In_1366);
xnor U2961 (N_2961,In_1311,In_1449);
nor U2962 (N_2962,In_1286,In_321);
and U2963 (N_2963,In_1208,In_991);
nor U2964 (N_2964,In_1360,In_317);
or U2965 (N_2965,In_959,In_1108);
nand U2966 (N_2966,In_203,In_1479);
and U2967 (N_2967,In_1396,In_377);
nor U2968 (N_2968,In_849,In_581);
nor U2969 (N_2969,In_80,In_887);
nor U2970 (N_2970,In_368,In_118);
nor U2971 (N_2971,In_676,In_18);
nand U2972 (N_2972,In_871,In_730);
nor U2973 (N_2973,In_188,In_290);
nor U2974 (N_2974,In_583,In_219);
nand U2975 (N_2975,In_789,In_954);
or U2976 (N_2976,In_677,In_1033);
or U2977 (N_2977,In_1448,In_1206);
nor U2978 (N_2978,In_898,In_1061);
nand U2979 (N_2979,In_50,In_133);
nor U2980 (N_2980,In_647,In_699);
or U2981 (N_2981,In_798,In_1350);
nor U2982 (N_2982,In_725,In_939);
and U2983 (N_2983,In_466,In_834);
or U2984 (N_2984,In_634,In_286);
nor U2985 (N_2985,In_674,In_1437);
or U2986 (N_2986,In_147,In_198);
xor U2987 (N_2987,In_616,In_1318);
nand U2988 (N_2988,In_873,In_568);
or U2989 (N_2989,In_466,In_579);
nor U2990 (N_2990,In_174,In_306);
and U2991 (N_2991,In_184,In_975);
xnor U2992 (N_2992,In_229,In_298);
and U2993 (N_2993,In_317,In_394);
xnor U2994 (N_2994,In_859,In_581);
nor U2995 (N_2995,In_1185,In_535);
nand U2996 (N_2996,In_382,In_597);
nand U2997 (N_2997,In_871,In_905);
nor U2998 (N_2998,In_1202,In_372);
and U2999 (N_2999,In_1360,In_467);
xor U3000 (N_3000,N_2045,N_2691);
nand U3001 (N_3001,N_861,N_1900);
xnor U3002 (N_3002,N_1007,N_1962);
nand U3003 (N_3003,N_1755,N_1510);
and U3004 (N_3004,N_2072,N_2767);
nor U3005 (N_3005,N_1552,N_2448);
or U3006 (N_3006,N_2737,N_1282);
and U3007 (N_3007,N_520,N_1766);
nand U3008 (N_3008,N_119,N_2046);
or U3009 (N_3009,N_1997,N_2517);
xor U3010 (N_3010,N_1194,N_2090);
nor U3011 (N_3011,N_1783,N_1916);
and U3012 (N_3012,N_2607,N_2304);
nor U3013 (N_3013,N_1173,N_2003);
and U3014 (N_3014,N_2702,N_2101);
nor U3015 (N_3015,N_329,N_1636);
and U3016 (N_3016,N_2378,N_1550);
xor U3017 (N_3017,N_2112,N_2688);
nand U3018 (N_3018,N_489,N_1349);
nand U3019 (N_3019,N_1751,N_2420);
or U3020 (N_3020,N_2703,N_1684);
nand U3021 (N_3021,N_1729,N_318);
or U3022 (N_3022,N_1655,N_1419);
xor U3023 (N_3023,N_1503,N_2163);
xor U3024 (N_3024,N_2357,N_49);
xor U3025 (N_3025,N_2575,N_105);
and U3026 (N_3026,N_2270,N_1673);
or U3027 (N_3027,N_1281,N_768);
or U3028 (N_3028,N_1789,N_2478);
nor U3029 (N_3029,N_2139,N_2274);
or U3030 (N_3030,N_441,N_1865);
xnor U3031 (N_3031,N_2418,N_1993);
nand U3032 (N_3032,N_1605,N_2155);
and U3033 (N_3033,N_1537,N_1357);
or U3034 (N_3034,N_2960,N_927);
nor U3035 (N_3035,N_2177,N_2993);
or U3036 (N_3036,N_2069,N_770);
or U3037 (N_3037,N_2059,N_482);
nand U3038 (N_3038,N_2701,N_101);
xnor U3039 (N_3039,N_1516,N_122);
nand U3040 (N_3040,N_1315,N_2999);
nor U3041 (N_3041,N_2561,N_1134);
and U3042 (N_3042,N_925,N_1512);
nor U3043 (N_3043,N_860,N_2757);
or U3044 (N_3044,N_2032,N_928);
nor U3045 (N_3045,N_2634,N_1781);
xnor U3046 (N_3046,N_236,N_2637);
or U3047 (N_3047,N_1892,N_2615);
and U3048 (N_3048,N_503,N_2589);
and U3049 (N_3049,N_64,N_2071);
nand U3050 (N_3050,N_1728,N_417);
xor U3051 (N_3051,N_2107,N_208);
and U3052 (N_3052,N_264,N_462);
xnor U3053 (N_3053,N_603,N_593);
nor U3054 (N_3054,N_1340,N_1198);
and U3055 (N_3055,N_1958,N_1578);
nor U3056 (N_3056,N_2769,N_1608);
xor U3057 (N_3057,N_2858,N_2138);
nor U3058 (N_3058,N_974,N_109);
nor U3059 (N_3059,N_2712,N_711);
xnor U3060 (N_3060,N_2754,N_1953);
and U3061 (N_3061,N_1041,N_335);
and U3062 (N_3062,N_280,N_2508);
nand U3063 (N_3063,N_2964,N_130);
xor U3064 (N_3064,N_2188,N_2797);
xnor U3065 (N_3065,N_912,N_99);
and U3066 (N_3066,N_1970,N_346);
nand U3067 (N_3067,N_2849,N_2813);
xor U3068 (N_3068,N_2472,N_2942);
and U3069 (N_3069,N_170,N_1443);
or U3070 (N_3070,N_2883,N_2037);
nor U3071 (N_3071,N_2599,N_437);
or U3072 (N_3072,N_2465,N_743);
nor U3073 (N_3073,N_2792,N_277);
xnor U3074 (N_3074,N_290,N_1476);
nor U3075 (N_3075,N_1133,N_788);
or U3076 (N_3076,N_2263,N_129);
nand U3077 (N_3077,N_2543,N_1581);
and U3078 (N_3078,N_1713,N_906);
xnor U3079 (N_3079,N_125,N_162);
nand U3080 (N_3080,N_2404,N_2531);
nand U3081 (N_3081,N_2036,N_1356);
nand U3082 (N_3082,N_314,N_874);
nor U3083 (N_3083,N_1393,N_2313);
nor U3084 (N_3084,N_1235,N_2388);
or U3085 (N_3085,N_2935,N_528);
nor U3086 (N_3086,N_1980,N_1754);
xor U3087 (N_3087,N_287,N_156);
or U3088 (N_3088,N_2565,N_1220);
xnor U3089 (N_3089,N_1272,N_1410);
and U3090 (N_3090,N_832,N_557);
and U3091 (N_3091,N_2996,N_1255);
nor U3092 (N_3092,N_1506,N_588);
or U3093 (N_3093,N_1325,N_710);
and U3094 (N_3094,N_863,N_2887);
nand U3095 (N_3095,N_1792,N_2015);
nor U3096 (N_3096,N_1870,N_2400);
or U3097 (N_3097,N_2320,N_2669);
xnor U3098 (N_3098,N_1613,N_1971);
and U3099 (N_3099,N_1278,N_1448);
xnor U3100 (N_3100,N_17,N_2641);
and U3101 (N_3101,N_2269,N_915);
xor U3102 (N_3102,N_2295,N_1224);
and U3103 (N_3103,N_2438,N_228);
or U3104 (N_3104,N_2879,N_2252);
nand U3105 (N_3105,N_1752,N_2096);
nand U3106 (N_3106,N_1029,N_2692);
or U3107 (N_3107,N_2650,N_2476);
or U3108 (N_3108,N_1875,N_2937);
or U3109 (N_3109,N_2201,N_507);
and U3110 (N_3110,N_1464,N_680);
and U3111 (N_3111,N_1565,N_418);
nor U3112 (N_3112,N_2550,N_1238);
and U3113 (N_3113,N_146,N_2548);
or U3114 (N_3114,N_1983,N_1351);
nand U3115 (N_3115,N_1364,N_334);
and U3116 (N_3116,N_357,N_944);
and U3117 (N_3117,N_853,N_972);
nand U3118 (N_3118,N_1905,N_486);
nor U3119 (N_3119,N_2770,N_732);
and U3120 (N_3120,N_2546,N_2848);
or U3121 (N_3121,N_2679,N_1482);
xor U3122 (N_3122,N_1168,N_2542);
and U3123 (N_3123,N_1172,N_1353);
or U3124 (N_3124,N_1504,N_2718);
and U3125 (N_3125,N_2804,N_1409);
xnor U3126 (N_3126,N_2827,N_851);
xnor U3127 (N_3127,N_2741,N_2065);
or U3128 (N_3128,N_960,N_103);
nand U3129 (N_3129,N_2678,N_2277);
xnor U3130 (N_3130,N_1700,N_690);
nand U3131 (N_3131,N_2834,N_426);
xnor U3132 (N_3132,N_244,N_1822);
nor U3133 (N_3133,N_717,N_1651);
nor U3134 (N_3134,N_1859,N_2549);
nor U3135 (N_3135,N_401,N_1215);
nand U3136 (N_3136,N_1470,N_2898);
and U3137 (N_3137,N_666,N_1549);
nand U3138 (N_3138,N_2401,N_794);
xnor U3139 (N_3139,N_1727,N_848);
nand U3140 (N_3140,N_903,N_2326);
or U3141 (N_3141,N_2972,N_2346);
nand U3142 (N_3142,N_2613,N_2226);
nand U3143 (N_3143,N_1279,N_2132);
and U3144 (N_3144,N_2785,N_2761);
xor U3145 (N_3145,N_982,N_1153);
nand U3146 (N_3146,N_783,N_1925);
xor U3147 (N_3147,N_31,N_2630);
nand U3148 (N_3148,N_834,N_2776);
nor U3149 (N_3149,N_530,N_923);
or U3150 (N_3150,N_1772,N_1573);
and U3151 (N_3151,N_57,N_265);
and U3152 (N_3152,N_899,N_551);
or U3153 (N_3153,N_2812,N_525);
nor U3154 (N_3154,N_694,N_2408);
nand U3155 (N_3155,N_706,N_2029);
xnor U3156 (N_3156,N_1342,N_2324);
or U3157 (N_3157,N_611,N_1844);
and U3158 (N_3158,N_1954,N_271);
or U3159 (N_3159,N_987,N_2588);
or U3160 (N_3160,N_2058,N_2953);
and U3161 (N_3161,N_2075,N_1917);
xor U3162 (N_3162,N_1780,N_2077);
and U3163 (N_3163,N_1074,N_494);
nor U3164 (N_3164,N_1525,N_2645);
nor U3165 (N_3165,N_2717,N_2413);
nand U3166 (N_3166,N_1522,N_1551);
or U3167 (N_3167,N_1439,N_2820);
and U3168 (N_3168,N_760,N_1484);
or U3169 (N_3169,N_247,N_2088);
xor U3170 (N_3170,N_2142,N_2176);
nor U3171 (N_3171,N_2219,N_839);
and U3172 (N_3172,N_402,N_273);
nand U3173 (N_3173,N_1141,N_674);
and U3174 (N_3174,N_2654,N_2869);
or U3175 (N_3175,N_1836,N_2578);
or U3176 (N_3176,N_2419,N_1231);
xnor U3177 (N_3177,N_804,N_1460);
nand U3178 (N_3178,N_1890,N_212);
and U3179 (N_3179,N_608,N_343);
nor U3180 (N_3180,N_877,N_1798);
xor U3181 (N_3181,N_1457,N_2782);
nor U3182 (N_3182,N_1668,N_498);
nor U3183 (N_3183,N_2127,N_1877);
nor U3184 (N_3184,N_1297,N_1438);
and U3185 (N_3185,N_1048,N_2405);
xnor U3186 (N_3186,N_2296,N_1248);
and U3187 (N_3187,N_1368,N_39);
nand U3188 (N_3188,N_533,N_2768);
nor U3189 (N_3189,N_2695,N_1082);
and U3190 (N_3190,N_2961,N_20);
or U3191 (N_3191,N_2113,N_1652);
xor U3192 (N_3192,N_1611,N_181);
nand U3193 (N_3193,N_1061,N_108);
or U3194 (N_3194,N_1465,N_967);
nor U3195 (N_3195,N_990,N_282);
xor U3196 (N_3196,N_1211,N_2221);
xor U3197 (N_3197,N_485,N_2467);
and U3198 (N_3198,N_398,N_270);
xnor U3199 (N_3199,N_2683,N_434);
nand U3200 (N_3200,N_427,N_1559);
nor U3201 (N_3201,N_2026,N_1534);
nand U3202 (N_3202,N_778,N_2522);
or U3203 (N_3203,N_1064,N_2507);
nor U3204 (N_3204,N_358,N_985);
nor U3205 (N_3205,N_2238,N_397);
and U3206 (N_3206,N_1968,N_283);
nor U3207 (N_3207,N_1547,N_2261);
xnor U3208 (N_3208,N_1992,N_1140);
nor U3209 (N_3209,N_759,N_667);
or U3210 (N_3210,N_2547,N_1214);
or U3211 (N_3211,N_729,N_307);
nand U3212 (N_3212,N_1285,N_591);
and U3213 (N_3213,N_1863,N_2351);
nor U3214 (N_3214,N_1112,N_2764);
xnor U3215 (N_3215,N_857,N_1533);
xor U3216 (N_3216,N_2114,N_1688);
xor U3217 (N_3217,N_2356,N_1891);
or U3218 (N_3218,N_1746,N_2699);
nand U3219 (N_3219,N_2586,N_1177);
nand U3220 (N_3220,N_1804,N_2627);
or U3221 (N_3221,N_2838,N_1286);
nor U3222 (N_3222,N_924,N_1005);
xnor U3223 (N_3223,N_1264,N_683);
or U3224 (N_3224,N_82,N_837);
xor U3225 (N_3225,N_2315,N_2681);
and U3226 (N_3226,N_1296,N_475);
nor U3227 (N_3227,N_2504,N_2605);
or U3228 (N_3228,N_1948,N_1414);
nor U3229 (N_3229,N_1878,N_275);
or U3230 (N_3230,N_471,N_1336);
nand U3231 (N_3231,N_1776,N_2134);
and U3232 (N_3232,N_1841,N_2506);
and U3233 (N_3233,N_1365,N_609);
nand U3234 (N_3234,N_180,N_563);
nand U3235 (N_3235,N_2752,N_2102);
xor U3236 (N_3236,N_703,N_1945);
and U3237 (N_3237,N_658,N_415);
or U3238 (N_3238,N_2213,N_2672);
or U3239 (N_3239,N_1190,N_2904);
or U3240 (N_3240,N_953,N_392);
and U3241 (N_3241,N_810,N_1678);
nand U3242 (N_3242,N_1429,N_2621);
xnor U3243 (N_3243,N_2924,N_1441);
nor U3244 (N_3244,N_1543,N_1692);
nor U3245 (N_3245,N_2215,N_2350);
nor U3246 (N_3246,N_2066,N_1824);
nand U3247 (N_3247,N_1160,N_2158);
nand U3248 (N_3248,N_2710,N_1389);
nand U3249 (N_3249,N_2974,N_311);
xor U3250 (N_3250,N_2122,N_1740);
nand U3251 (N_3251,N_1260,N_2020);
nor U3252 (N_3252,N_480,N_1679);
or U3253 (N_3253,N_339,N_948);
xnor U3254 (N_3254,N_2895,N_195);
nor U3255 (N_3255,N_2194,N_716);
and U3256 (N_3256,N_292,N_1136);
nand U3257 (N_3257,N_2409,N_1591);
xor U3258 (N_3258,N_223,N_204);
nor U3259 (N_3259,N_2461,N_336);
and U3260 (N_3260,N_1879,N_446);
and U3261 (N_3261,N_1720,N_2690);
xor U3262 (N_3262,N_295,N_356);
or U3263 (N_3263,N_636,N_2667);
nand U3264 (N_3264,N_980,N_2402);
and U3265 (N_3265,N_281,N_1363);
xnor U3266 (N_3266,N_1869,N_754);
nor U3267 (N_3267,N_2168,N_955);
xor U3268 (N_3268,N_1846,N_429);
or U3269 (N_3269,N_1219,N_1615);
and U3270 (N_3270,N_931,N_1629);
and U3271 (N_3271,N_2230,N_118);
xor U3272 (N_3272,N_886,N_1417);
nor U3273 (N_3273,N_341,N_2529);
xnor U3274 (N_3274,N_2369,N_2940);
nor U3275 (N_3275,N_2713,N_421);
xnor U3276 (N_3276,N_2570,N_887);
nor U3277 (N_3277,N_1753,N_1893);
nor U3278 (N_3278,N_2900,N_1873);
nand U3279 (N_3279,N_519,N_2070);
or U3280 (N_3280,N_1912,N_1817);
and U3281 (N_3281,N_308,N_896);
or U3282 (N_3282,N_1531,N_2815);
xor U3283 (N_3283,N_1000,N_278);
nor U3284 (N_3284,N_1135,N_428);
and U3285 (N_3285,N_231,N_2422);
or U3286 (N_3286,N_1070,N_2524);
and U3287 (N_3287,N_2619,N_200);
nor U3288 (N_3288,N_1797,N_882);
or U3289 (N_3289,N_2302,N_2023);
and U3290 (N_3290,N_299,N_2628);
or U3291 (N_3291,N_84,N_995);
or U3292 (N_3292,N_1094,N_2027);
or U3293 (N_3293,N_1179,N_586);
and U3294 (N_3294,N_1940,N_1697);
nor U3295 (N_3295,N_1178,N_888);
and U3296 (N_3296,N_1300,N_670);
or U3297 (N_3297,N_220,N_2911);
xnor U3298 (N_3298,N_230,N_126);
xnor U3299 (N_3299,N_2343,N_1258);
or U3300 (N_3300,N_2919,N_865);
nor U3301 (N_3301,N_2720,N_479);
and U3302 (N_3302,N_1690,N_1935);
or U3303 (N_3303,N_2731,N_1075);
nor U3304 (N_3304,N_1864,N_1583);
xnor U3305 (N_3305,N_1202,N_1084);
nor U3306 (N_3306,N_1257,N_583);
nand U3307 (N_3307,N_2079,N_306);
nor U3308 (N_3308,N_2334,N_340);
or U3309 (N_3309,N_2606,N_2923);
or U3310 (N_3310,N_2225,N_1180);
and U3311 (N_3311,N_1961,N_1164);
and U3312 (N_3312,N_545,N_1657);
and U3313 (N_3313,N_2884,N_933);
and U3314 (N_3314,N_1274,N_2178);
and U3315 (N_3315,N_391,N_2914);
and U3316 (N_3316,N_425,N_2264);
xnor U3317 (N_3317,N_1210,N_250);
and U3318 (N_3318,N_1671,N_905);
xor U3319 (N_3319,N_1100,N_2284);
nand U3320 (N_3320,N_2666,N_1721);
and U3321 (N_3321,N_2509,N_577);
or U3322 (N_3322,N_1883,N_2951);
and U3323 (N_3323,N_1350,N_1155);
nand U3324 (N_3324,N_2938,N_2514);
nor U3325 (N_3325,N_2283,N_2930);
or U3326 (N_3326,N_1062,N_504);
or U3327 (N_3327,N_1127,N_1735);
or U3328 (N_3328,N_1787,N_815);
and U3329 (N_3329,N_1032,N_2209);
or U3330 (N_3330,N_734,N_199);
nor U3331 (N_3331,N_2988,N_1696);
xor U3332 (N_3332,N_2321,N_469);
xor U3333 (N_3333,N_422,N_2187);
and U3334 (N_3334,N_590,N_1837);
xnor U3335 (N_3335,N_94,N_1520);
nor U3336 (N_3336,N_2686,N_2931);
or U3337 (N_3337,N_87,N_227);
nand U3338 (N_3338,N_2067,N_139);
or U3339 (N_3339,N_1023,N_1145);
xor U3340 (N_3340,N_1254,N_1796);
nor U3341 (N_3341,N_144,N_1313);
and U3342 (N_3342,N_1101,N_812);
xor U3343 (N_3343,N_2966,N_150);
or U3344 (N_3344,N_2427,N_387);
nand U3345 (N_3345,N_612,N_1575);
nand U3346 (N_3346,N_1239,N_613);
nand U3347 (N_3347,N_587,N_1646);
nor U3348 (N_3348,N_2245,N_2843);
and U3349 (N_3349,N_2571,N_1607);
and U3350 (N_3350,N_803,N_396);
nand U3351 (N_3351,N_645,N_1113);
nand U3352 (N_3352,N_248,N_2906);
or U3353 (N_3353,N_534,N_89);
or U3354 (N_3354,N_1816,N_1374);
xor U3355 (N_3355,N_350,N_1097);
nand U3356 (N_3356,N_112,N_739);
nor U3357 (N_3357,N_556,N_2169);
nor U3358 (N_3358,N_2104,N_1040);
xor U3359 (N_3359,N_289,N_2863);
nor U3360 (N_3360,N_1904,N_2841);
and U3361 (N_3361,N_1208,N_817);
or U3362 (N_3362,N_2493,N_328);
nor U3363 (N_3363,N_805,N_1475);
or U3364 (N_3364,N_332,N_1649);
or U3365 (N_3365,N_2925,N_268);
and U3366 (N_3366,N_2166,N_1267);
or U3367 (N_3367,N_2161,N_750);
or U3368 (N_3368,N_205,N_1977);
or U3369 (N_3369,N_1345,N_1959);
nor U3370 (N_3370,N_2994,N_2729);
nor U3371 (N_3371,N_384,N_1165);
or U3372 (N_3372,N_1014,N_1509);
nand U3373 (N_3373,N_901,N_673);
nand U3374 (N_3374,N_2028,N_2464);
nor U3375 (N_3375,N_1310,N_77);
nor U3376 (N_3376,N_2331,N_301);
nand U3377 (N_3377,N_1078,N_2362);
and U3378 (N_3378,N_259,N_1452);
and U3379 (N_3379,N_830,N_1535);
or U3380 (N_3380,N_191,N_349);
nand U3381 (N_3381,N_26,N_1631);
nor U3382 (N_3382,N_751,N_2905);
nand U3383 (N_3383,N_1137,N_9);
and U3384 (N_3384,N_1909,N_476);
nand U3385 (N_3385,N_2243,N_1944);
or U3386 (N_3386,N_2241,N_158);
xnor U3387 (N_3387,N_1502,N_23);
and U3388 (N_3388,N_309,N_194);
xnor U3389 (N_3389,N_481,N_2394);
nand U3390 (N_3390,N_876,N_1268);
and U3391 (N_3391,N_1705,N_2410);
or U3392 (N_3392,N_2762,N_366);
and U3393 (N_3393,N_727,N_1811);
xnor U3394 (N_3394,N_1790,N_1446);
or U3395 (N_3395,N_2693,N_911);
nor U3396 (N_3396,N_1401,N_2902);
xor U3397 (N_3397,N_2763,N_85);
or U3398 (N_3398,N_664,N_1329);
or U3399 (N_3399,N_1628,N_651);
or U3400 (N_3400,N_2487,N_501);
nor U3401 (N_3401,N_2826,N_1990);
nand U3402 (N_3402,N_543,N_214);
nor U3403 (N_3403,N_2748,N_1109);
nand U3404 (N_3404,N_628,N_149);
nand U3405 (N_3405,N_926,N_1191);
xor U3406 (N_3406,N_2477,N_1989);
and U3407 (N_3407,N_73,N_1610);
nor U3408 (N_3408,N_1963,N_958);
or U3409 (N_3409,N_2095,N_1926);
nand U3410 (N_3410,N_81,N_1110);
or U3411 (N_3411,N_1347,N_1730);
xnor U3412 (N_3412,N_2856,N_688);
nor U3413 (N_3413,N_1,N_74);
nand U3414 (N_3414,N_1725,N_1530);
nor U3415 (N_3415,N_1249,N_649);
nor U3416 (N_3416,N_707,N_2556);
nor U3417 (N_3417,N_2564,N_1450);
nand U3418 (N_3418,N_1913,N_477);
or U3419 (N_3419,N_1570,N_458);
and U3420 (N_3420,N_363,N_1150);
or U3421 (N_3421,N_1633,N_1229);
and U3422 (N_3422,N_1335,N_2643);
nand U3423 (N_3423,N_226,N_2483);
or U3424 (N_3424,N_1616,N_1466);
nor U3425 (N_3425,N_4,N_2894);
or U3426 (N_3426,N_2516,N_975);
xor U3427 (N_3427,N_1769,N_2352);
and U3428 (N_3428,N_1677,N_1785);
or U3429 (N_3429,N_1333,N_1732);
nand U3430 (N_3430,N_964,N_276);
xnor U3431 (N_3431,N_767,N_881);
nor U3432 (N_3432,N_2715,N_1923);
and U3433 (N_3433,N_1016,N_93);
or U3434 (N_3434,N_2668,N_1672);
xor U3435 (N_3435,N_2242,N_1698);
and U3436 (N_3436,N_2392,N_998);
nor U3437 (N_3437,N_584,N_916);
nor U3438 (N_3438,N_1719,N_672);
nor U3439 (N_3439,N_186,N_858);
nand U3440 (N_3440,N_2457,N_1632);
and U3441 (N_3441,N_2063,N_2661);
xnor U3442 (N_3442,N_1802,N_646);
or U3443 (N_3443,N_992,N_2236);
nor U3444 (N_3444,N_2677,N_2083);
or U3445 (N_3445,N_973,N_956);
or U3446 (N_3446,N_1212,N_1251);
and U3447 (N_3447,N_2256,N_597);
and U3448 (N_3448,N_1943,N_354);
or U3449 (N_3449,N_1589,N_1493);
nand U3450 (N_3450,N_2623,N_1650);
and U3451 (N_3451,N_1316,N_60);
and U3452 (N_3452,N_634,N_1232);
nand U3453 (N_3453,N_2100,N_639);
nand U3454 (N_3454,N_2287,N_2825);
and U3455 (N_3455,N_8,N_1861);
nor U3456 (N_3456,N_878,N_2437);
nand U3457 (N_3457,N_2480,N_2927);
and U3458 (N_3458,N_745,N_1588);
nor U3459 (N_3459,N_1620,N_1488);
and U3460 (N_3460,N_1277,N_2498);
nand U3461 (N_3461,N_324,N_1577);
or U3462 (N_3462,N_1236,N_852);
and U3463 (N_3463,N_2515,N_2532);
and U3464 (N_3464,N_465,N_2557);
or U3465 (N_3465,N_1002,N_2631);
nor U3466 (N_3466,N_1964,N_669);
xnor U3467 (N_3467,N_1284,N_381);
and U3468 (N_3468,N_1326,N_1116);
or U3469 (N_3469,N_1523,N_1188);
and U3470 (N_3470,N_722,N_131);
and U3471 (N_3471,N_1664,N_1920);
nor U3472 (N_3472,N_172,N_1667);
xor U3473 (N_3473,N_872,N_2053);
nor U3474 (N_3474,N_2439,N_2976);
and U3475 (N_3475,N_1969,N_2584);
and U3476 (N_3476,N_2881,N_2309);
and U3477 (N_3477,N_2329,N_2742);
or U3478 (N_3478,N_650,N_2361);
nor U3479 (N_3479,N_1169,N_576);
nand U3480 (N_3480,N_2587,N_2126);
nor U3481 (N_3481,N_1808,N_554);
or U3482 (N_3482,N_97,N_2746);
xor U3483 (N_3483,N_2195,N_827);
and U3484 (N_3484,N_1405,N_900);
xor U3485 (N_3485,N_1592,N_811);
xnor U3486 (N_3486,N_2193,N_943);
or U3487 (N_3487,N_589,N_1418);
and U3488 (N_3488,N_2829,N_2091);
nor U3489 (N_3489,N_976,N_898);
and U3490 (N_3490,N_748,N_2165);
nand U3491 (N_3491,N_1854,N_1899);
xnor U3492 (N_3492,N_1791,N_1280);
nor U3493 (N_3493,N_1461,N_1930);
and U3494 (N_3494,N_2980,N_2948);
and U3495 (N_3495,N_491,N_2198);
or U3496 (N_3496,N_1321,N_1385);
xor U3497 (N_3497,N_166,N_2794);
xnor U3498 (N_3498,N_1911,N_1095);
nand U3499 (N_3499,N_1289,N_1323);
xnor U3500 (N_3500,N_174,N_2376);
xnor U3501 (N_3501,N_1712,N_2878);
nand U3502 (N_3502,N_633,N_2445);
xnor U3503 (N_3503,N_2921,N_2779);
and U3504 (N_3504,N_2234,N_1521);
nor U3505 (N_3505,N_1931,N_1230);
nor U3506 (N_3506,N_2087,N_183);
nand U3507 (N_3507,N_936,N_2865);
nand U3508 (N_3508,N_2040,N_1747);
xor U3509 (N_3509,N_1480,N_2603);
and U3510 (N_3510,N_1731,N_431);
nor U3511 (N_3511,N_117,N_2338);
and U3512 (N_3512,N_1885,N_1225);
nor U3513 (N_3513,N_1777,N_2051);
or U3514 (N_3514,N_2470,N_136);
or U3515 (N_3515,N_1237,N_2981);
or U3516 (N_3516,N_1749,N_2482);
xor U3517 (N_3517,N_2390,N_1848);
xor U3518 (N_3518,N_2330,N_2610);
nor U3519 (N_3519,N_2220,N_258);
xnor U3520 (N_3520,N_2175,N_1782);
and U3521 (N_3521,N_1472,N_1815);
and U3522 (N_3522,N_986,N_606);
or U3523 (N_3523,N_435,N_2082);
xnor U3524 (N_3524,N_140,N_474);
nor U3525 (N_3525,N_1845,N_719);
nor U3526 (N_3526,N_430,N_2639);
nor U3527 (N_3527,N_1666,N_951);
nand U3528 (N_3528,N_2955,N_866);
nand U3529 (N_3529,N_2728,N_1361);
and U3530 (N_3530,N_1539,N_35);
nand U3531 (N_3531,N_913,N_2004);
and U3532 (N_3532,N_687,N_1233);
and U3533 (N_3533,N_2618,N_121);
or U3534 (N_3534,N_2818,N_2491);
xor U3535 (N_3535,N_55,N_371);
and U3536 (N_3536,N_1115,N_1077);
or U3537 (N_3537,N_2282,N_106);
and U3538 (N_3538,N_1079,N_1028);
or U3539 (N_3539,N_789,N_1463);
nor U3540 (N_3540,N_2760,N_2775);
nand U3541 (N_3541,N_1821,N_2459);
and U3542 (N_3542,N_1850,N_2857);
nand U3543 (N_3543,N_2105,N_133);
nor U3544 (N_3544,N_1324,N_2218);
nor U3545 (N_3545,N_27,N_2602);
nand U3546 (N_3546,N_1723,N_495);
and U3547 (N_3547,N_2796,N_1998);
nand U3548 (N_3548,N_2039,N_1043);
xor U3549 (N_3549,N_18,N_2867);
xor U3550 (N_3550,N_302,N_601);
xnor U3551 (N_3551,N_92,N_497);
and U3552 (N_3552,N_2202,N_1038);
or U3553 (N_3553,N_1431,N_1950);
and U3554 (N_3554,N_2874,N_2662);
nand U3555 (N_3555,N_1880,N_1524);
nor U3556 (N_3556,N_124,N_1445);
and U3557 (N_3557,N_1328,N_1868);
nand U3558 (N_3558,N_1057,N_66);
nor U3559 (N_3559,N_257,N_656);
xor U3560 (N_3560,N_632,N_1553);
and U3561 (N_3561,N_2093,N_61);
xnor U3562 (N_3562,N_2907,N_1283);
nand U3563 (N_3563,N_1928,N_2990);
or U3564 (N_3564,N_1974,N_2038);
or U3565 (N_3565,N_1051,N_1999);
xnor U3566 (N_3566,N_1167,N_2174);
xnor U3567 (N_3567,N_578,N_2788);
and U3568 (N_3568,N_2123,N_2012);
nor U3569 (N_3569,N_880,N_2016);
nand U3570 (N_3570,N_1176,N_2417);
xnor U3571 (N_3571,N_1453,N_2545);
nor U3572 (N_3572,N_2853,N_2021);
and U3573 (N_3573,N_1055,N_1250);
nor U3574 (N_3574,N_2222,N_405);
xor U3575 (N_3575,N_1170,N_294);
and U3576 (N_3576,N_348,N_605);
or U3577 (N_3577,N_1812,N_801);
or U3578 (N_3578,N_490,N_2789);
or U3579 (N_3579,N_2840,N_1762);
nand U3580 (N_3580,N_1091,N_2922);
and U3581 (N_3581,N_941,N_1955);
or U3582 (N_3582,N_460,N_241);
nor U3583 (N_3583,N_1704,N_1857);
nor U3584 (N_3584,N_2989,N_1492);
nand U3585 (N_3585,N_873,N_2383);
nor U3586 (N_3586,N_2018,N_390);
xnor U3587 (N_3587,N_2963,N_1189);
xor U3588 (N_3588,N_2325,N_1532);
nor U3589 (N_3589,N_2696,N_1426);
nand U3590 (N_3590,N_1120,N_2705);
and U3591 (N_3591,N_2453,N_2821);
and U3592 (N_3592,N_2246,N_2381);
or U3593 (N_3593,N_448,N_993);
xnor U3594 (N_3594,N_2181,N_631);
nand U3595 (N_3595,N_1146,N_1757);
xor U3596 (N_3596,N_2591,N_648);
or U3597 (N_3597,N_1653,N_1408);
nor U3598 (N_3598,N_274,N_2425);
xor U3599 (N_3599,N_2449,N_1087);
nand U3600 (N_3600,N_243,N_342);
nand U3601 (N_3601,N_1624,N_2952);
nand U3602 (N_3602,N_2537,N_2424);
nand U3603 (N_3603,N_2186,N_167);
nor U3604 (N_3604,N_747,N_2162);
nor U3605 (N_3605,N_455,N_2434);
nor U3606 (N_3606,N_260,N_240);
nand U3607 (N_3607,N_2511,N_2959);
or U3608 (N_3608,N_2559,N_1670);
and U3609 (N_3609,N_2382,N_671);
nor U3610 (N_3610,N_54,N_1370);
and U3611 (N_3611,N_2958,N_46);
xor U3612 (N_3612,N_2061,N_718);
or U3613 (N_3613,N_2444,N_604);
or U3614 (N_3614,N_952,N_1795);
xnor U3615 (N_3615,N_347,N_724);
nor U3616 (N_3616,N_2224,N_320);
nand U3617 (N_3617,N_1625,N_731);
xor U3618 (N_3618,N_2977,N_113);
or U3619 (N_3619,N_1148,N_285);
xor U3620 (N_3620,N_2851,N_814);
nor U3621 (N_3621,N_1501,N_1026);
xor U3622 (N_3622,N_1371,N_1567);
xnor U3623 (N_3623,N_1111,N_2010);
and U3624 (N_3624,N_2510,N_561);
nand U3625 (N_3625,N_213,N_676);
or U3626 (N_3626,N_1558,N_2626);
nor U3627 (N_3627,N_2495,N_1346);
and U3628 (N_3628,N_22,N_2913);
nand U3629 (N_3629,N_408,N_2880);
nor U3630 (N_3630,N_1378,N_654);
and U3631 (N_3631,N_893,N_1626);
and U3632 (N_3632,N_1984,N_2756);
or U3633 (N_3633,N_2594,N_2275);
nand U3634 (N_3634,N_360,N_2755);
or U3635 (N_3635,N_1487,N_524);
or U3636 (N_3636,N_592,N_351);
and U3637 (N_3637,N_1554,N_1639);
nand U3638 (N_3638,N_1621,N_1396);
and U3639 (N_3639,N_2978,N_2525);
and U3640 (N_3640,N_2502,N_681);
or U3641 (N_3641,N_678,N_2852);
and U3642 (N_3642,N_2652,N_2136);
nor U3643 (N_3643,N_412,N_1922);
xnor U3644 (N_3644,N_1433,N_785);
xnor U3645 (N_3645,N_305,N_2711);
nor U3646 (N_3646,N_1246,N_2698);
and U3647 (N_3647,N_2030,N_1689);
and U3648 (N_3648,N_1745,N_2497);
xor U3649 (N_3649,N_1528,N_574);
or U3650 (N_3650,N_553,N_2991);
and U3651 (N_3651,N_2971,N_2997);
nor U3652 (N_3652,N_1341,N_2680);
and U3653 (N_3653,N_1847,N_771);
nand U3654 (N_3654,N_2704,N_1544);
or U3655 (N_3655,N_1741,N_157);
nand U3656 (N_3656,N_2893,N_135);
or U3657 (N_3657,N_192,N_1312);
nand U3658 (N_3658,N_2787,N_777);
nand U3659 (N_3659,N_843,N_2073);
xnor U3660 (N_3660,N_1226,N_1092);
xor U3661 (N_3661,N_978,N_368);
xor U3662 (N_3662,N_1699,N_977);
xnor U3663 (N_3663,N_786,N_2771);
xor U3664 (N_3664,N_1206,N_1404);
and U3665 (N_3665,N_2656,N_2009);
and U3666 (N_3666,N_721,N_1395);
and U3667 (N_3667,N_1726,N_189);
nor U3668 (N_3668,N_145,N_1597);
or U3669 (N_3669,N_2541,N_1663);
nor U3670 (N_3670,N_1600,N_2998);
xnor U3671 (N_3671,N_1369,N_891);
and U3672 (N_3672,N_2150,N_198);
xnor U3673 (N_3673,N_2043,N_2431);
and U3674 (N_3674,N_2896,N_2866);
xnor U3675 (N_3675,N_1951,N_1978);
or U3676 (N_3676,N_2360,N_330);
and U3677 (N_3677,N_2447,N_2385);
or U3678 (N_3678,N_128,N_147);
nor U3679 (N_3679,N_464,N_1256);
xnor U3680 (N_3680,N_2665,N_1569);
and U3681 (N_3681,N_1020,N_1193);
nand U3682 (N_3682,N_1813,N_2620);
and U3683 (N_3683,N_304,N_2744);
nor U3684 (N_3684,N_1459,N_262);
and U3685 (N_3685,N_539,N_2970);
or U3686 (N_3686,N_487,N_1398);
xnor U3687 (N_3687,N_1602,N_2805);
nand U3688 (N_3688,N_746,N_1744);
nand U3689 (N_3689,N_2580,N_2740);
xor U3690 (N_3690,N_773,N_1058);
nor U3691 (N_3691,N_2778,N_2947);
and U3692 (N_3692,N_1306,N_2798);
nand U3693 (N_3693,N_516,N_2430);
and U3694 (N_3694,N_1407,N_2816);
or U3695 (N_3695,N_352,N_310);
or U3696 (N_3696,N_2137,N_457);
nand U3697 (N_3697,N_1827,N_871);
nand U3698 (N_3698,N_369,N_362);
xnor U3699 (N_3699,N_2533,N_1004);
or U3700 (N_3700,N_2854,N_1081);
and U3701 (N_3701,N_325,N_1025);
nor U3702 (N_3702,N_1656,N_1209);
nand U3703 (N_3703,N_1496,N_2086);
nor U3704 (N_3704,N_1582,N_615);
nand U3705 (N_3705,N_1008,N_715);
or U3706 (N_3706,N_1681,N_1985);
nor U3707 (N_3707,N_263,N_338);
xnor U3708 (N_3708,N_1929,N_968);
nand U3709 (N_3709,N_2373,N_1918);
nor U3710 (N_3710,N_447,N_2673);
nand U3711 (N_3711,N_1003,N_921);
and U3712 (N_3712,N_766,N_1637);
and U3713 (N_3713,N_2658,N_365);
nand U3714 (N_3714,N_2941,N_298);
nand U3715 (N_3715,N_2322,N_154);
or U3716 (N_3716,N_764,N_1083);
xnor U3717 (N_3717,N_48,N_316);
nor U3718 (N_3718,N_386,N_994);
xor U3719 (N_3719,N_2708,N_326);
nand U3720 (N_3720,N_966,N_2540);
and U3721 (N_3721,N_2379,N_2609);
nand U3722 (N_3722,N_41,N_2859);
and U3723 (N_3723,N_2055,N_2831);
or U3724 (N_3724,N_761,N_2719);
nor U3725 (N_3725,N_571,N_1163);
xnor U3726 (N_3726,N_700,N_1490);
and U3727 (N_3727,N_2278,N_1860);
and U3728 (N_3728,N_2232,N_2519);
nor U3729 (N_3729,N_1903,N_1661);
and U3730 (N_3730,N_2633,N_1413);
xor U3731 (N_3731,N_1645,N_25);
or U3732 (N_3732,N_2899,N_1151);
or U3733 (N_3733,N_2986,N_1497);
xor U3734 (N_3734,N_2266,N_296);
or U3735 (N_3735,N_470,N_1829);
xnor U3736 (N_3736,N_1818,N_744);
nand U3737 (N_3737,N_1031,N_1852);
nor U3738 (N_3738,N_2151,N_63);
and U3739 (N_3739,N_288,N_1183);
xor U3740 (N_3740,N_234,N_291);
xor U3741 (N_3741,N_1768,N_772);
xor U3742 (N_3742,N_2629,N_451);
nand U3743 (N_3743,N_337,N_846);
nor U3744 (N_3744,N_1701,N_2576);
and U3745 (N_3745,N_2239,N_2254);
and U3746 (N_3746,N_1245,N_1442);
nor U3747 (N_3747,N_2945,N_2651);
nand U3748 (N_3748,N_1665,N_232);
and U3749 (N_3749,N_902,N_2253);
nand U3750 (N_3750,N_937,N_393);
xnor U3751 (N_3751,N_1706,N_705);
and U3752 (N_3752,N_2732,N_2106);
nand U3753 (N_3753,N_29,N_463);
nand U3754 (N_3754,N_630,N_594);
and U3755 (N_3755,N_1458,N_2653);
nor U3756 (N_3756,N_2109,N_2211);
xnor U3757 (N_3757,N_2468,N_1934);
or U3758 (N_3758,N_2554,N_2423);
nand U3759 (N_3759,N_1784,N_303);
xnor U3760 (N_3760,N_741,N_1750);
nor U3761 (N_3761,N_382,N_2227);
nand U3762 (N_3762,N_1156,N_2552);
xnor U3763 (N_3763,N_2518,N_626);
or U3764 (N_3764,N_456,N_2271);
xor U3765 (N_3765,N_1674,N_970);
and U3766 (N_3766,N_188,N_211);
nor U3767 (N_3767,N_2845,N_1102);
xnor U3768 (N_3768,N_2216,N_442);
or U3769 (N_3769,N_2706,N_2359);
xnor U3770 (N_3770,N_1319,N_799);
nand U3771 (N_3771,N_1623,N_2180);
or U3772 (N_3772,N_1896,N_168);
nand U3773 (N_3773,N_930,N_2709);
nand U3774 (N_3774,N_2108,N_1449);
nor U3775 (N_3775,N_1894,N_317);
or U3776 (N_3776,N_1853,N_738);
nor U3777 (N_3777,N_752,N_2396);
nor U3778 (N_3778,N_2262,N_1643);
and U3779 (N_3779,N_685,N_897);
xor U3780 (N_3780,N_2157,N_2806);
nor U3781 (N_3781,N_2097,N_1354);
and U3782 (N_3782,N_686,N_1786);
nand U3783 (N_3783,N_708,N_1563);
or U3784 (N_3784,N_2967,N_1468);
or U3785 (N_3785,N_957,N_2929);
nand U3786 (N_3786,N_934,N_850);
xnor U3787 (N_3787,N_1018,N_2830);
and U3788 (N_3788,N_569,N_2579);
xor U3789 (N_3789,N_894,N_2707);
xnor U3790 (N_3790,N_1331,N_2407);
nor U3791 (N_3791,N_1499,N_1849);
nor U3792 (N_3792,N_468,N_2056);
or U3793 (N_3793,N_1380,N_1541);
nor U3794 (N_3794,N_2416,N_493);
nor U3795 (N_3795,N_1096,N_540);
xor U3796 (N_3796,N_2822,N_70);
xnor U3797 (N_3797,N_202,N_102);
and U3798 (N_3798,N_647,N_2110);
or U3799 (N_3799,N_515,N_689);
nand U3800 (N_3800,N_2339,N_2915);
nand U3801 (N_3801,N_1367,N_2926);
nor U3802 (N_3802,N_2057,N_2984);
and U3803 (N_3803,N_1030,N_1831);
nor U3804 (N_3804,N_266,N_2987);
nor U3805 (N_3805,N_2733,N_562);
nand U3806 (N_3806,N_2614,N_508);
or U3807 (N_3807,N_2145,N_855);
nand U3808 (N_3808,N_652,N_1301);
or U3809 (N_3809,N_907,N_2022);
nor U3810 (N_3810,N_2267,N_321);
and U3811 (N_3811,N_2888,N_2299);
xnor U3812 (N_3812,N_730,N_1640);
nor U3813 (N_3813,N_1546,N_160);
nand U3814 (N_3814,N_1069,N_665);
xnor U3815 (N_3815,N_2314,N_1838);
nor U3816 (N_3816,N_2456,N_1834);
nand U3817 (N_3817,N_2428,N_797);
or U3818 (N_3818,N_246,N_499);
and U3819 (N_3819,N_2985,N_2814);
and U3820 (N_3820,N_2837,N_1320);
nand U3821 (N_3821,N_2442,N_807);
nand U3822 (N_3822,N_34,N_617);
and U3823 (N_3823,N_2484,N_1159);
nand U3824 (N_3824,N_2292,N_2534);
nand U3825 (N_3825,N_2738,N_72);
nand U3826 (N_3826,N_2205,N_502);
xor U3827 (N_3827,N_2544,N_445);
xor U3828 (N_3828,N_2312,N_2170);
nand U3829 (N_3829,N_1222,N_229);
or U3830 (N_3830,N_1595,N_2928);
nor U3831 (N_3831,N_2625,N_1975);
nand U3832 (N_3832,N_120,N_697);
nand U3833 (N_3833,N_2835,N_781);
and U3834 (N_3834,N_641,N_2054);
xnor U3835 (N_3835,N_1538,N_159);
xor U3836 (N_3836,N_1157,N_610);
nand U3837 (N_3837,N_1855,N_353);
nor U3838 (N_3838,N_1144,N_62);
nor U3839 (N_3839,N_1252,N_2872);
or U3840 (N_3840,N_663,N_161);
and U3841 (N_3841,N_1024,N_1108);
and U3842 (N_3842,N_935,N_1764);
and U3843 (N_3843,N_2817,N_2801);
nor U3844 (N_3844,N_735,N_2574);
nand U3845 (N_3845,N_1106,N_2481);
or U3846 (N_3846,N_2739,N_1478);
nor U3847 (N_3847,N_1269,N_1474);
or U3848 (N_3848,N_922,N_2441);
nor U3849 (N_3849,N_2595,N_756);
or U3850 (N_3850,N_1598,N_818);
nor U3851 (N_3851,N_1644,N_2129);
or U3852 (N_3852,N_638,N_765);
nor U3853 (N_3853,N_2772,N_2671);
nand U3854 (N_3854,N_2365,N_454);
nor U3855 (N_3855,N_1939,N_2311);
or U3856 (N_3856,N_1760,N_884);
nor U3857 (N_3857,N_1049,N_2501);
nand U3858 (N_3858,N_370,N_2355);
or U3859 (N_3859,N_1288,N_1709);
and U3860 (N_3860,N_40,N_802);
or U3861 (N_3861,N_30,N_1139);
nor U3862 (N_3862,N_940,N_2950);
nor U3863 (N_3863,N_2882,N_2901);
nand U3864 (N_3864,N_2047,N_2463);
xnor U3865 (N_3865,N_885,N_21);
and U3866 (N_3866,N_2979,N_1383);
xnor U3867 (N_3867,N_2862,N_821);
nand U3868 (N_3868,N_1828,N_1253);
or U3869 (N_3869,N_1742,N_165);
and U3870 (N_3870,N_47,N_1748);
nor U3871 (N_3871,N_98,N_1669);
xnor U3872 (N_3872,N_2475,N_2539);
nand U3873 (N_3873,N_2196,N_1366);
xnor U3874 (N_3874,N_2406,N_2572);
nand U3875 (N_3875,N_1564,N_1710);
and U3876 (N_3876,N_971,N_2130);
nor U3877 (N_3877,N_840,N_1942);
nor U3878 (N_3878,N_868,N_380);
xor U3879 (N_3879,N_757,N_677);
and U3880 (N_3880,N_1184,N_28);
nand U3881 (N_3881,N_531,N_1519);
or U3882 (N_3882,N_914,N_1001);
nand U3883 (N_3883,N_1622,N_1199);
nand U3884 (N_3884,N_2153,N_2632);
or U3885 (N_3885,N_2192,N_12);
or U3886 (N_3886,N_1810,N_1540);
nand U3887 (N_3887,N_1914,N_2569);
xnor U3888 (N_3888,N_532,N_153);
nand U3889 (N_3889,N_787,N_2647);
nor U3890 (N_3890,N_249,N_1660);
xnor U3891 (N_3891,N_2172,N_95);
nor U3892 (N_3892,N_763,N_478);
nand U3893 (N_3893,N_2611,N_997);
nor U3894 (N_3894,N_345,N_643);
xnor U3895 (N_3895,N_1809,N_835);
nand U3896 (N_3896,N_820,N_2799);
or U3897 (N_3897,N_1105,N_2398);
and U3898 (N_3898,N_2255,N_424);
xnor U3899 (N_3899,N_225,N_107);
nor U3900 (N_3900,N_2395,N_1560);
nand U3901 (N_3901,N_1076,N_2551);
xnor U3902 (N_3902,N_2523,N_704);
nor U3903 (N_3903,N_720,N_2414);
or U3904 (N_3904,N_1047,N_2751);
nor U3905 (N_3905,N_207,N_1052);
xor U3906 (N_3906,N_2297,N_723);
or U3907 (N_3907,N_2001,N_2310);
xnor U3908 (N_3908,N_5,N_965);
nand U3909 (N_3909,N_1491,N_2513);
or U3910 (N_3910,N_1117,N_2936);
nor U3911 (N_3911,N_879,N_141);
nor U3912 (N_3912,N_2167,N_2839);
nand U3913 (N_3913,N_2660,N_1814);
nor U3914 (N_3914,N_1936,N_1218);
nor U3915 (N_3915,N_65,N_1590);
or U3916 (N_3916,N_1053,N_702);
nand U3917 (N_3917,N_596,N_1066);
xor U3918 (N_3918,N_2290,N_2116);
nor U3919 (N_3919,N_197,N_784);
xnor U3920 (N_3920,N_2520,N_2191);
nor U3921 (N_3921,N_627,N_2573);
xnor U3922 (N_3922,N_521,N_1933);
nand U3923 (N_3923,N_184,N_86);
xor U3924 (N_3924,N_550,N_2118);
nor U3925 (N_3925,N_1555,N_1067);
nor U3926 (N_3926,N_331,N_2675);
and U3927 (N_3927,N_1500,N_2212);
nand U3928 (N_3928,N_1006,N_775);
and U3929 (N_3929,N_71,N_1767);
nor U3930 (N_3930,N_2847,N_2897);
or U3931 (N_3931,N_1932,N_2766);
or U3932 (N_3932,N_1763,N_749);
or U3933 (N_3933,N_2811,N_2281);
nor U3934 (N_3934,N_2567,N_2081);
nor U3935 (N_3935,N_2140,N_2479);
or U3936 (N_3936,N_2208,N_1511);
nand U3937 (N_3937,N_2289,N_1411);
nand U3938 (N_3938,N_2159,N_1065);
and U3939 (N_3939,N_467,N_1332);
xor U3940 (N_3940,N_164,N_2060);
nor U3941 (N_3941,N_2305,N_2824);
nor U3942 (N_3942,N_185,N_75);
nor U3943 (N_3943,N_1695,N_564);
nor U3944 (N_3944,N_2340,N_2133);
xnor U3945 (N_3945,N_111,N_2934);
and U3946 (N_3946,N_1275,N_2646);
xnor U3947 (N_3947,N_2260,N_1056);
and U3948 (N_3948,N_1462,N_2214);
or U3949 (N_3949,N_2886,N_892);
nor U3950 (N_3950,N_284,N_637);
and U3951 (N_3951,N_123,N_2597);
nand U3952 (N_3952,N_148,N_1071);
or U3953 (N_3953,N_1377,N_659);
nand U3954 (N_3954,N_698,N_657);
and U3955 (N_3955,N_2349,N_1451);
or U3956 (N_3956,N_558,N_452);
nand U3957 (N_3957,N_143,N_2367);
and U3958 (N_3958,N_1734,N_1012);
nor U3959 (N_3959,N_1400,N_1303);
nor U3960 (N_3960,N_1469,N_1825);
nand U3961 (N_3961,N_2803,N_2759);
or U3962 (N_3962,N_1432,N_459);
nor U3963 (N_3963,N_2622,N_675);
or U3964 (N_3964,N_235,N_1820);
nor U3965 (N_3965,N_1976,N_2429);
nand U3966 (N_3966,N_2115,N_736);
xor U3967 (N_3967,N_1093,N_699);
nor U3968 (N_3968,N_423,N_96);
or U3969 (N_3969,N_2538,N_1343);
nor U3970 (N_3970,N_2049,N_2301);
or U3971 (N_3971,N_1242,N_379);
nand U3972 (N_3972,N_2017,N_823);
or U3973 (N_3973,N_2724,N_132);
or U3974 (N_3974,N_1390,N_419);
or U3975 (N_3975,N_1738,N_2248);
and U3976 (N_3976,N_917,N_69);
nor U3977 (N_3977,N_2784,N_2204);
or U3978 (N_3978,N_2391,N_2415);
or U3979 (N_3979,N_2199,N_1557);
nand U3980 (N_3980,N_179,N_2185);
xor U3981 (N_3981,N_2025,N_1872);
nand U3982 (N_3982,N_653,N_1680);
nor U3983 (N_3983,N_1099,N_2530);
or U3984 (N_3984,N_1648,N_315);
nand U3985 (N_3985,N_842,N_1617);
nor U3986 (N_3986,N_2426,N_2503);
or U3987 (N_3987,N_1430,N_2786);
and U3988 (N_3988,N_909,N_2307);
and U3989 (N_3989,N_361,N_1247);
and U3990 (N_3990,N_1384,N_660);
and U3991 (N_3991,N_864,N_1473);
nor U3992 (N_3992,N_1562,N_1118);
xnor U3993 (N_3993,N_709,N_961);
nand U3994 (N_3994,N_1322,N_1819);
nand U3995 (N_3995,N_1715,N_1195);
nand U3996 (N_3996,N_2111,N_1594);
nand U3997 (N_3997,N_1085,N_1103);
or U3998 (N_3998,N_555,N_2861);
xnor U3999 (N_3999,N_2317,N_2957);
nand U4000 (N_4000,N_251,N_2700);
nor U4001 (N_4001,N_1486,N_2179);
xor U4002 (N_4002,N_2585,N_2577);
nand U4003 (N_4003,N_1415,N_908);
nand U4004 (N_4004,N_1662,N_537);
nor U4005 (N_4005,N_163,N_1036);
and U4006 (N_4006,N_620,N_2014);
or U4007 (N_4007,N_261,N_216);
xor U4008 (N_4008,N_1702,N_1599);
or U4009 (N_4009,N_461,N_2050);
nand U4010 (N_4010,N_1895,N_2103);
nor U4011 (N_4011,N_695,N_1033);
or U4012 (N_4012,N_959,N_560);
and U4013 (N_4013,N_411,N_2636);
or U4014 (N_4014,N_312,N_2068);
and U4015 (N_4015,N_2203,N_2568);
or U4016 (N_4016,N_1707,N_742);
or U4017 (N_4017,N_2387,N_1886);
xor U4018 (N_4018,N_2288,N_1882);
and U4019 (N_4019,N_1759,N_1638);
or U4020 (N_4020,N_1566,N_1187);
and U4021 (N_4021,N_209,N_1758);
and U4022 (N_4022,N_15,N_1420);
nor U4023 (N_4023,N_1221,N_2436);
or U4024 (N_4024,N_1495,N_2024);
and U4025 (N_4025,N_152,N_1536);
nor U4026 (N_4026,N_2807,N_2535);
nand U4027 (N_4027,N_1119,N_573);
or U4028 (N_4028,N_822,N_1682);
and U4029 (N_4029,N_1045,N_829);
nor U4030 (N_4030,N_819,N_2146);
and U4031 (N_4031,N_753,N_1114);
nor U4032 (N_4032,N_449,N_2868);
and U4033 (N_4033,N_1424,N_378);
and U4034 (N_4034,N_693,N_1901);
or U4035 (N_4035,N_869,N_1587);
nand U4036 (N_4036,N_2160,N_190);
nand U4037 (N_4037,N_1125,N_696);
nand U4038 (N_4038,N_1060,N_2780);
nor U4039 (N_4039,N_2685,N_1527);
nor U4040 (N_4040,N_2249,N_1579);
nor U4041 (N_4041,N_2358,N_1454);
xor U4042 (N_4042,N_11,N_2917);
or U4043 (N_4043,N_725,N_1355);
nor U4044 (N_4044,N_2593,N_267);
nand U4045 (N_4045,N_1803,N_2348);
nand U4046 (N_4046,N_1130,N_2276);
and U4047 (N_4047,N_2364,N_1265);
or U4048 (N_4048,N_2286,N_518);
nor U4049 (N_4049,N_1171,N_2144);
or U4050 (N_4050,N_2013,N_3);
nor U4051 (N_4051,N_1576,N_2008);
xor U4052 (N_4052,N_1217,N_1960);
or U4053 (N_4053,N_1691,N_1881);
xnor U4054 (N_4054,N_1635,N_1308);
nand U4055 (N_4055,N_1291,N_215);
xor U4056 (N_4056,N_1456,N_2908);
nor U4057 (N_4057,N_2973,N_2600);
and U4058 (N_4058,N_500,N_1192);
xnor U4059 (N_4059,N_661,N_254);
nor U4060 (N_4060,N_989,N_2663);
nand U4061 (N_4061,N_406,N_809);
nor U4062 (N_4062,N_572,N_1915);
nand U4063 (N_4063,N_2592,N_1982);
nand U4064 (N_4064,N_1039,N_2268);
nor U4065 (N_4065,N_1035,N_2962);
nor U4066 (N_4066,N_79,N_1434);
nand U4067 (N_4067,N_2583,N_1158);
nor U4068 (N_4068,N_344,N_2616);
nor U4069 (N_4069,N_2119,N_1627);
and U4070 (N_4070,N_2257,N_1614);
xnor U4071 (N_4071,N_1344,N_1338);
nand U4072 (N_4072,N_825,N_2377);
xor U4073 (N_4073,N_580,N_1388);
nor U4074 (N_4074,N_1197,N_1489);
nand U4075 (N_4075,N_2975,N_1348);
nand U4076 (N_4076,N_2730,N_1223);
xnor U4077 (N_4077,N_1908,N_1737);
nand U4078 (N_4078,N_414,N_862);
and U4079 (N_4079,N_2892,N_910);
or U4080 (N_4080,N_2135,N_2064);
and U4081 (N_4081,N_950,N_404);
or U4082 (N_4082,N_2285,N_364);
or U4083 (N_4083,N_2259,N_1483);
nor U4084 (N_4084,N_2143,N_1924);
nand U4085 (N_4085,N_2716,N_2499);
nor U4086 (N_4086,N_782,N_10);
and U4087 (N_4087,N_962,N_1515);
xnor U4088 (N_4088,N_1572,N_2052);
nand U4089 (N_4089,N_2624,N_1833);
xnor U4090 (N_4090,N_2098,N_14);
or U4091 (N_4091,N_826,N_2697);
nor U4092 (N_4092,N_1362,N_2094);
or U4093 (N_4093,N_359,N_1887);
nor U4094 (N_4094,N_2435,N_2366);
or U4095 (N_4095,N_1471,N_932);
or U4096 (N_4096,N_2642,N_2910);
and U4097 (N_4097,N_1050,N_2223);
or U4098 (N_4098,N_1376,N_2335);
or U4099 (N_4099,N_210,N_1017);
nor U4100 (N_4100,N_473,N_1293);
and U4101 (N_4101,N_1382,N_1545);
nor U4102 (N_4102,N_513,N_1387);
xor U4103 (N_4103,N_668,N_552);
nor U4104 (N_4104,N_238,N_1862);
or U4105 (N_4105,N_2120,N_1874);
nand U4106 (N_4106,N_1427,N_2148);
or U4107 (N_4107,N_1843,N_535);
or U4108 (N_4108,N_1477,N_2684);
nand U4109 (N_4109,N_1162,N_614);
xor U4110 (N_4110,N_904,N_2612);
xnor U4111 (N_4111,N_854,N_849);
xnor U4112 (N_4112,N_2562,N_1181);
xnor U4113 (N_4113,N_1104,N_1676);
or U4114 (N_4114,N_256,N_450);
nor U4115 (N_4115,N_949,N_313);
xor U4116 (N_4116,N_76,N_222);
and U4117 (N_4117,N_2795,N_2291);
or U4118 (N_4118,N_1447,N_1981);
nand U4119 (N_4119,N_1941,N_1203);
or U4120 (N_4120,N_1603,N_1805);
or U4121 (N_4121,N_1263,N_1708);
or U4122 (N_4122,N_575,N_389);
or U4123 (N_4123,N_483,N_327);
nand U4124 (N_4124,N_2555,N_1204);
xor U4125 (N_4125,N_2891,N_2389);
or U4126 (N_4126,N_377,N_1585);
xor U4127 (N_4127,N_2933,N_2454);
xnor U4128 (N_4128,N_151,N_2034);
nand U4129 (N_4129,N_623,N_115);
nor U4130 (N_4130,N_1402,N_2657);
nand U4131 (N_4131,N_409,N_867);
nand U4132 (N_4132,N_2333,N_138);
or U4133 (N_4133,N_171,N_224);
nor U4134 (N_4134,N_1714,N_51);
and U4135 (N_4135,N_1132,N_1907);
nand U4136 (N_4136,N_217,N_2664);
or U4137 (N_4137,N_1311,N_779);
nor U4138 (N_4138,N_137,N_1807);
or U4139 (N_4139,N_2995,N_1889);
nand U4140 (N_4140,N_1073,N_253);
or U4141 (N_4141,N_1304,N_1123);
or U4142 (N_4142,N_2251,N_1683);
xnor U4143 (N_4143,N_538,N_2582);
or U4144 (N_4144,N_1010,N_1518);
and U4145 (N_4145,N_510,N_1175);
xnor U4146 (N_4146,N_1440,N_536);
and U4147 (N_4147,N_237,N_1927);
nand U4148 (N_4148,N_2125,N_774);
or U4149 (N_4149,N_1871,N_1561);
xor U4150 (N_4150,N_1919,N_2035);
or U4151 (N_4151,N_1756,N_219);
or U4152 (N_4152,N_438,N_1201);
nand U4153 (N_4153,N_2946,N_2372);
nand U4154 (N_4154,N_1778,N_644);
xnor U4155 (N_4155,N_2655,N_2800);
or U4156 (N_4156,N_1835,N_1422);
and U4157 (N_4157,N_1059,N_1302);
xor U4158 (N_4158,N_1658,N_1724);
nor U4159 (N_4159,N_2190,N_1979);
nor U4160 (N_4160,N_2873,N_1021);
or U4161 (N_4161,N_2943,N_595);
or U4162 (N_4162,N_2810,N_796);
xor U4163 (N_4163,N_1508,N_1126);
nor U4164 (N_4164,N_2128,N_2466);
xor U4165 (N_4165,N_38,N_319);
nand U4166 (N_4166,N_1779,N_1718);
or U4167 (N_4167,N_1897,N_1015);
xnor U4168 (N_4168,N_1200,N_2920);
xnor U4169 (N_4169,N_388,N_1241);
nand U4170 (N_4170,N_2397,N_1596);
nor U4171 (N_4171,N_870,N_619);
and U4172 (N_4172,N_2210,N_795);
or U4173 (N_4173,N_1381,N_1399);
xor U4174 (N_4174,N_1262,N_1358);
xnor U4175 (N_4175,N_155,N_2062);
nand U4176 (N_4176,N_1166,N_2280);
and U4177 (N_4177,N_239,N_2601);
or U4178 (N_4178,N_529,N_1722);
nor U4179 (N_4179,N_1967,N_2949);
nor U4180 (N_4180,N_2486,N_662);
and U4181 (N_4181,N_2471,N_173);
or U4182 (N_4182,N_2581,N_127);
nor U4183 (N_4183,N_1659,N_2455);
nor U4184 (N_4184,N_2117,N_440);
nor U4185 (N_4185,N_484,N_1556);
nand U4186 (N_4186,N_2124,N_988);
nor U4187 (N_4187,N_2725,N_1318);
nor U4188 (N_4188,N_56,N_831);
nor U4189 (N_4189,N_622,N_444);
or U4190 (N_4190,N_1856,N_2041);
xnor U4191 (N_4191,N_1858,N_2048);
nand U4192 (N_4192,N_1287,N_792);
nand U4193 (N_4193,N_385,N_37);
nand U4194 (N_4194,N_1360,N_374);
nand U4195 (N_4195,N_2183,N_1152);
nor U4196 (N_4196,N_293,N_2635);
nor U4197 (N_4197,N_376,N_1403);
nand U4198 (N_4198,N_2154,N_43);
nor U4199 (N_4199,N_2490,N_1921);
or U4200 (N_4200,N_517,N_355);
and U4201 (N_4201,N_1068,N_91);
nand U4202 (N_4202,N_1840,N_2909);
nand U4203 (N_4203,N_2505,N_2903);
or U4204 (N_4204,N_182,N_1124);
nor U4205 (N_4205,N_2598,N_2687);
and U4206 (N_4206,N_2864,N_1494);
and U4207 (N_4207,N_2197,N_1009);
nor U4208 (N_4208,N_1601,N_1711);
or U4209 (N_4209,N_2694,N_187);
or U4210 (N_4210,N_1266,N_889);
nand U4211 (N_4211,N_272,N_1481);
and U4212 (N_4212,N_1013,N_1485);
xnor U4213 (N_4213,N_981,N_547);
and U4214 (N_4214,N_1054,N_2446);
nand U4215 (N_4215,N_1739,N_1703);
or U4216 (N_4216,N_828,N_1088);
and U4217 (N_4217,N_2674,N_0);
nand U4218 (N_4218,N_1571,N_938);
nor U4219 (N_4219,N_2745,N_2336);
xor U4220 (N_4220,N_2458,N_2659);
nand U4221 (N_4221,N_2279,N_1654);
xnor U4222 (N_4222,N_999,N_2019);
or U4223 (N_4223,N_2939,N_1423);
and U4224 (N_4224,N_110,N_2536);
and U4225 (N_4225,N_758,N_1299);
and U4226 (N_4226,N_242,N_1080);
or U4227 (N_4227,N_544,N_1851);
nand U4228 (N_4228,N_2932,N_2173);
nor U4229 (N_4229,N_506,N_1295);
and U4230 (N_4230,N_2332,N_740);
xor U4231 (N_4231,N_824,N_413);
nand U4232 (N_4232,N_2916,N_624);
or U4233 (N_4233,N_2844,N_104);
nand U4234 (N_4234,N_568,N_1213);
nor U4235 (N_4235,N_841,N_2521);
and U4236 (N_4236,N_2485,N_52);
and U4237 (N_4237,N_2152,N_2450);
and U4238 (N_4238,N_2074,N_2494);
nand U4239 (N_4239,N_1298,N_1513);
nand U4240 (N_4240,N_375,N_1686);
and U4241 (N_4241,N_655,N_1244);
or U4242 (N_4242,N_1996,N_2386);
xnor U4243 (N_4243,N_2982,N_59);
nor U4244 (N_4244,N_2750,N_2273);
nor U4245 (N_4245,N_549,N_2247);
nand U4246 (N_4246,N_2156,N_1694);
xnor U4247 (N_4247,N_806,N_542);
xor U4248 (N_4248,N_1437,N_598);
or U4249 (N_4249,N_2604,N_1906);
nand U4250 (N_4250,N_2033,N_512);
or U4251 (N_4251,N_1305,N_1046);
xor U4252 (N_4252,N_1479,N_1339);
xor U4253 (N_4253,N_567,N_983);
nor U4254 (N_4254,N_1593,N_2876);
xor U4255 (N_4255,N_2384,N_1273);
xor U4256 (N_4256,N_2085,N_2080);
and U4257 (N_4257,N_2500,N_2560);
xor U4258 (N_4258,N_2099,N_600);
xnor U4259 (N_4259,N_1234,N_963);
nor U4260 (N_4260,N_2722,N_1687);
or U4261 (N_4261,N_2734,N_2727);
nand U4262 (N_4262,N_2006,N_1832);
or U4263 (N_4263,N_1761,N_44);
and U4264 (N_4264,N_1207,N_496);
or U4265 (N_4265,N_1196,N_2131);
and U4266 (N_4266,N_394,N_2889);
nand U4267 (N_4267,N_2676,N_2265);
nor U4268 (N_4268,N_2089,N_1444);
nand U4269 (N_4269,N_836,N_2258);
xnor U4270 (N_4270,N_2149,N_1072);
or U4271 (N_4271,N_701,N_1957);
or U4272 (N_4272,N_2306,N_890);
nand U4273 (N_4273,N_2649,N_1205);
and U4274 (N_4274,N_439,N_33);
xnor U4275 (N_4275,N_2808,N_2337);
xor U4276 (N_4276,N_991,N_2735);
nand U4277 (N_4277,N_2860,N_640);
xor U4278 (N_4278,N_206,N_2250);
nand U4279 (N_4279,N_1375,N_2875);
nor U4280 (N_4280,N_505,N_522);
nand U4281 (N_4281,N_1397,N_2836);
and U4282 (N_4282,N_1647,N_2000);
nand U4283 (N_4283,N_2380,N_1794);
or U4284 (N_4284,N_527,N_1412);
or U4285 (N_4285,N_1991,N_1276);
nor U4286 (N_4286,N_1995,N_1261);
nand U4287 (N_4287,N_1507,N_1946);
xor U4288 (N_4288,N_2670,N_2452);
or U4289 (N_4289,N_682,N_1986);
nor U4290 (N_4290,N_2492,N_2563);
xnor U4291 (N_4291,N_1034,N_1334);
nor U4292 (N_4292,N_1949,N_1406);
nand U4293 (N_4293,N_1063,N_726);
nor U4294 (N_4294,N_2007,N_2345);
and U4295 (N_4295,N_2200,N_1826);
nand U4296 (N_4296,N_1612,N_88);
nand U4297 (N_4297,N_2850,N_443);
and U4298 (N_4298,N_1089,N_2777);
nor U4299 (N_4299,N_920,N_16);
nand U4300 (N_4300,N_2871,N_969);
nand U4301 (N_4301,N_2473,N_2648);
xnor U4302 (N_4302,N_859,N_2412);
and U4303 (N_4303,N_1154,N_1128);
nor U4304 (N_4304,N_175,N_201);
nand U4305 (N_4305,N_1733,N_453);
xnor U4306 (N_4306,N_1044,N_844);
xnor U4307 (N_4307,N_416,N_714);
nor U4308 (N_4308,N_1042,N_1337);
nor U4309 (N_4309,N_1771,N_692);
xor U4310 (N_4310,N_2743,N_684);
or U4311 (N_4311,N_2,N_2229);
or U4312 (N_4312,N_1161,N_1988);
and U4313 (N_4313,N_581,N_286);
xor U4314 (N_4314,N_2308,N_1314);
or U4315 (N_4315,N_1373,N_2969);
nand U4316 (N_4316,N_2819,N_395);
and U4317 (N_4317,N_1174,N_1216);
or U4318 (N_4318,N_1788,N_116);
nand U4319 (N_4319,N_838,N_2638);
nand U4320 (N_4320,N_546,N_2965);
xnor U4321 (N_4321,N_793,N_1542);
or U4322 (N_4322,N_2078,N_2328);
nor U4323 (N_4323,N_472,N_2526);
and U4324 (N_4324,N_2189,N_2954);
nor U4325 (N_4325,N_939,N_1138);
and U4326 (N_4326,N_1290,N_2790);
nor U4327 (N_4327,N_2002,N_1574);
nand U4328 (N_4328,N_90,N_333);
and U4329 (N_4329,N_400,N_399);
or U4330 (N_4330,N_616,N_1604);
nor U4331 (N_4331,N_2512,N_1548);
and U4332 (N_4332,N_178,N_383);
nand U4333 (N_4333,N_2753,N_1586);
xnor U4334 (N_4334,N_68,N_2462);
or U4335 (N_4335,N_733,N_36);
xnor U4336 (N_4336,N_2832,N_780);
or U4337 (N_4337,N_2474,N_712);
and U4338 (N_4338,N_1526,N_1228);
or U4339 (N_4339,N_2723,N_559);
nor U4340 (N_4340,N_176,N_2147);
and U4341 (N_4341,N_13,N_1416);
nand U4342 (N_4342,N_2370,N_2528);
xnor U4343 (N_4343,N_2721,N_1641);
xor U4344 (N_4344,N_2363,N_1774);
and U4345 (N_4345,N_196,N_432);
and U4346 (N_4346,N_1956,N_67);
xnor U4347 (N_4347,N_2433,N_2855);
xnor U4348 (N_4348,N_2793,N_621);
or U4349 (N_4349,N_1421,N_776);
xor U4350 (N_4350,N_177,N_618);
nor U4351 (N_4351,N_420,N_833);
nand U4352 (N_4352,N_221,N_1011);
nor U4353 (N_4353,N_1240,N_1937);
and U4354 (N_4354,N_1830,N_1630);
nor U4355 (N_4355,N_728,N_2944);
nand U4356 (N_4356,N_625,N_1182);
or U4357 (N_4357,N_1359,N_984);
nand U4358 (N_4358,N_19,N_2005);
xnor U4359 (N_4359,N_2421,N_755);
nand U4360 (N_4360,N_2774,N_737);
xor U4361 (N_4361,N_1243,N_2327);
or U4362 (N_4362,N_1801,N_433);
nor U4363 (N_4363,N_2758,N_2488);
nand U4364 (N_4364,N_1938,N_1372);
or U4365 (N_4365,N_566,N_2164);
nor U4366 (N_4366,N_2076,N_373);
xor U4367 (N_4367,N_2749,N_2141);
or U4368 (N_4368,N_2726,N_1436);
nand U4369 (N_4369,N_2781,N_1965);
nor U4370 (N_4370,N_1122,N_1019);
and U4371 (N_4371,N_942,N_1773);
xnor U4372 (N_4372,N_83,N_1270);
xnor U4373 (N_4373,N_883,N_2374);
and U4374 (N_4374,N_322,N_50);
xor U4375 (N_4375,N_1634,N_808);
or U4376 (N_4376,N_790,N_1271);
and U4377 (N_4377,N_1947,N_2042);
nand U4378 (N_4378,N_1121,N_255);
or U4379 (N_4379,N_2347,N_1743);
nor U4380 (N_4380,N_1902,N_323);
nor U4381 (N_4381,N_492,N_2432);
or U4382 (N_4382,N_466,N_2323);
or U4383 (N_4383,N_403,N_2809);
nand U4384 (N_4384,N_2870,N_585);
xnor U4385 (N_4385,N_2469,N_1143);
or U4386 (N_4386,N_1131,N_2294);
and U4387 (N_4387,N_800,N_2527);
nor U4388 (N_4388,N_2736,N_78);
nor U4389 (N_4389,N_816,N_2316);
xnor U4390 (N_4390,N_2992,N_2773);
and U4391 (N_4391,N_2235,N_979);
and U4392 (N_4392,N_579,N_1425);
nand U4393 (N_4393,N_2171,N_1529);
xor U4394 (N_4394,N_582,N_218);
or U4395 (N_4395,N_2272,N_1799);
nand U4396 (N_4396,N_1685,N_2375);
and U4397 (N_4397,N_996,N_523);
xor U4398 (N_4398,N_1842,N_203);
xor U4399 (N_4399,N_1147,N_279);
nand U4400 (N_4400,N_1618,N_233);
xor U4401 (N_4401,N_2553,N_1876);
and U4402 (N_4402,N_1716,N_1609);
xor U4403 (N_4403,N_1107,N_1386);
nor U4404 (N_4404,N_798,N_509);
or U4405 (N_4405,N_2823,N_1806);
or U4406 (N_4406,N_2451,N_1619);
nand U4407 (N_4407,N_565,N_2918);
nand U4408 (N_4408,N_607,N_1580);
nand U4409 (N_4409,N_2912,N_1675);
and U4410 (N_4410,N_2233,N_372);
or U4411 (N_4411,N_2747,N_2403);
and U4412 (N_4412,N_918,N_2293);
xor U4413 (N_4413,N_2890,N_2217);
xnor U4414 (N_4414,N_2783,N_2341);
nand U4415 (N_4415,N_32,N_1292);
xnor U4416 (N_4416,N_1823,N_1717);
nand U4417 (N_4417,N_2590,N_2206);
nand U4418 (N_4418,N_1307,N_2596);
or U4419 (N_4419,N_1693,N_2244);
nor U4420 (N_4420,N_599,N_2640);
and U4421 (N_4421,N_845,N_1352);
nand U4422 (N_4422,N_2842,N_2121);
nor U4423 (N_4423,N_80,N_2342);
or U4424 (N_4424,N_410,N_2983);
nor U4425 (N_4425,N_1149,N_2303);
xor U4426 (N_4426,N_2689,N_929);
xnor U4427 (N_4427,N_1952,N_2608);
or U4428 (N_4428,N_2566,N_1584);
nor U4429 (N_4429,N_1090,N_875);
nor U4430 (N_4430,N_762,N_2489);
nor U4431 (N_4431,N_1765,N_2182);
or U4432 (N_4432,N_2368,N_1428);
or U4433 (N_4433,N_1505,N_2791);
or U4434 (N_4434,N_2956,N_1839);
nand U4435 (N_4435,N_1142,N_2443);
and U4436 (N_4436,N_142,N_2084);
and U4437 (N_4437,N_45,N_1392);
xnor U4438 (N_4438,N_58,N_895);
xor U4439 (N_4439,N_813,N_2877);
and U4440 (N_4440,N_1327,N_1098);
and U4441 (N_4441,N_954,N_2399);
nor U4442 (N_4442,N_1455,N_2393);
and U4443 (N_4443,N_1259,N_1770);
or U4444 (N_4444,N_1317,N_679);
nor U4445 (N_4445,N_713,N_2300);
xor U4446 (N_4446,N_1394,N_2371);
nor U4447 (N_4447,N_193,N_1884);
and U4448 (N_4448,N_2354,N_945);
nand U4449 (N_4449,N_856,N_2319);
and U4450 (N_4450,N_1866,N_245);
xor U4451 (N_4451,N_1037,N_2460);
or U4452 (N_4452,N_1391,N_2092);
nor U4453 (N_4453,N_2228,N_847);
nor U4454 (N_4454,N_269,N_2617);
xor U4455 (N_4455,N_1972,N_1309);
nor U4456 (N_4456,N_2318,N_1086);
nor U4457 (N_4457,N_1793,N_367);
xnor U4458 (N_4458,N_1910,N_602);
and U4459 (N_4459,N_2833,N_541);
nor U4460 (N_4460,N_488,N_691);
xnor U4461 (N_4461,N_548,N_2044);
or U4462 (N_4462,N_1185,N_1379);
nor U4463 (N_4463,N_1568,N_511);
xor U4464 (N_4464,N_1294,N_1514);
xnor U4465 (N_4465,N_1027,N_24);
and U4466 (N_4466,N_947,N_1330);
and U4467 (N_4467,N_2231,N_1973);
nor U4468 (N_4468,N_2558,N_2885);
nor U4469 (N_4469,N_526,N_919);
or U4470 (N_4470,N_2353,N_1498);
and U4471 (N_4471,N_1022,N_2237);
nand U4472 (N_4472,N_2828,N_1186);
nand U4473 (N_4473,N_407,N_642);
or U4474 (N_4474,N_1994,N_1517);
nand U4475 (N_4475,N_2184,N_1800);
nor U4476 (N_4476,N_2644,N_1966);
xnor U4477 (N_4477,N_297,N_114);
or U4478 (N_4478,N_1888,N_946);
or U4479 (N_4479,N_2846,N_2011);
and U4480 (N_4480,N_2298,N_1987);
and U4481 (N_4481,N_1606,N_514);
nand U4482 (N_4482,N_1129,N_169);
xor U4483 (N_4483,N_1227,N_1736);
nor U4484 (N_4484,N_1775,N_2344);
nor U4485 (N_4485,N_252,N_2765);
and U4486 (N_4486,N_635,N_2682);
or U4487 (N_4487,N_6,N_2968);
nor U4488 (N_4488,N_1467,N_100);
or U4489 (N_4489,N_2207,N_1642);
or U4490 (N_4490,N_42,N_2411);
nand U4491 (N_4491,N_2031,N_791);
and U4492 (N_4492,N_769,N_629);
nand U4493 (N_4493,N_300,N_2440);
or U4494 (N_4494,N_1867,N_7);
and U4495 (N_4495,N_53,N_2714);
nand U4496 (N_4496,N_2802,N_570);
nand U4497 (N_4497,N_134,N_1898);
or U4498 (N_4498,N_2496,N_1435);
and U4499 (N_4499,N_436,N_2240);
nor U4500 (N_4500,N_2484,N_1080);
xor U4501 (N_4501,N_104,N_2277);
or U4502 (N_4502,N_628,N_526);
xor U4503 (N_4503,N_1370,N_1387);
nor U4504 (N_4504,N_1904,N_1567);
nor U4505 (N_4505,N_1647,N_502);
nor U4506 (N_4506,N_2571,N_499);
xor U4507 (N_4507,N_2914,N_747);
nor U4508 (N_4508,N_810,N_59);
nand U4509 (N_4509,N_2200,N_298);
xor U4510 (N_4510,N_1040,N_705);
nand U4511 (N_4511,N_2746,N_711);
or U4512 (N_4512,N_3,N_1714);
xor U4513 (N_4513,N_14,N_933);
xor U4514 (N_4514,N_2224,N_2628);
or U4515 (N_4515,N_2866,N_2218);
nand U4516 (N_4516,N_1079,N_2311);
nand U4517 (N_4517,N_1464,N_880);
and U4518 (N_4518,N_539,N_2120);
xor U4519 (N_4519,N_1493,N_2295);
and U4520 (N_4520,N_1100,N_1847);
or U4521 (N_4521,N_1303,N_333);
or U4522 (N_4522,N_2314,N_251);
nand U4523 (N_4523,N_2614,N_2480);
nor U4524 (N_4524,N_1593,N_1112);
xor U4525 (N_4525,N_274,N_1815);
and U4526 (N_4526,N_2860,N_2050);
or U4527 (N_4527,N_509,N_918);
xnor U4528 (N_4528,N_1079,N_2207);
or U4529 (N_4529,N_504,N_1125);
xor U4530 (N_4530,N_2977,N_990);
or U4531 (N_4531,N_2905,N_1470);
or U4532 (N_4532,N_625,N_1747);
nand U4533 (N_4533,N_834,N_2399);
and U4534 (N_4534,N_1440,N_180);
xnor U4535 (N_4535,N_2854,N_2070);
nor U4536 (N_4536,N_2159,N_977);
and U4537 (N_4537,N_2429,N_640);
and U4538 (N_4538,N_969,N_2205);
or U4539 (N_4539,N_538,N_2654);
xnor U4540 (N_4540,N_2798,N_1783);
and U4541 (N_4541,N_1368,N_924);
and U4542 (N_4542,N_1902,N_2750);
or U4543 (N_4543,N_227,N_1834);
or U4544 (N_4544,N_2895,N_367);
nor U4545 (N_4545,N_857,N_43);
or U4546 (N_4546,N_1672,N_1773);
or U4547 (N_4547,N_511,N_1817);
xnor U4548 (N_4548,N_2948,N_902);
nand U4549 (N_4549,N_1570,N_1977);
and U4550 (N_4550,N_2462,N_2388);
nand U4551 (N_4551,N_1929,N_1304);
xor U4552 (N_4552,N_1393,N_2388);
nand U4553 (N_4553,N_2763,N_1177);
nand U4554 (N_4554,N_2100,N_2158);
and U4555 (N_4555,N_1484,N_2291);
nor U4556 (N_4556,N_2636,N_2477);
and U4557 (N_4557,N_1479,N_1372);
or U4558 (N_4558,N_595,N_1362);
xor U4559 (N_4559,N_1061,N_2014);
nor U4560 (N_4560,N_2965,N_2308);
or U4561 (N_4561,N_2937,N_2323);
xor U4562 (N_4562,N_2337,N_1335);
or U4563 (N_4563,N_776,N_2181);
and U4564 (N_4564,N_2115,N_1587);
nor U4565 (N_4565,N_982,N_2566);
or U4566 (N_4566,N_1466,N_493);
nand U4567 (N_4567,N_147,N_24);
xor U4568 (N_4568,N_1278,N_1616);
xnor U4569 (N_4569,N_627,N_2787);
and U4570 (N_4570,N_655,N_1746);
nor U4571 (N_4571,N_2126,N_2857);
and U4572 (N_4572,N_2147,N_1470);
nor U4573 (N_4573,N_839,N_2049);
xnor U4574 (N_4574,N_420,N_2507);
xor U4575 (N_4575,N_579,N_2483);
nand U4576 (N_4576,N_55,N_2377);
or U4577 (N_4577,N_777,N_195);
xnor U4578 (N_4578,N_2508,N_354);
xnor U4579 (N_4579,N_8,N_2450);
or U4580 (N_4580,N_475,N_2114);
and U4581 (N_4581,N_296,N_2318);
nand U4582 (N_4582,N_1559,N_508);
xnor U4583 (N_4583,N_685,N_765);
nand U4584 (N_4584,N_278,N_272);
nor U4585 (N_4585,N_876,N_1572);
and U4586 (N_4586,N_1835,N_521);
nor U4587 (N_4587,N_280,N_2608);
nand U4588 (N_4588,N_2647,N_683);
nor U4589 (N_4589,N_485,N_2677);
or U4590 (N_4590,N_1523,N_2338);
xnor U4591 (N_4591,N_2809,N_1811);
nor U4592 (N_4592,N_1302,N_2759);
or U4593 (N_4593,N_731,N_2589);
nand U4594 (N_4594,N_2417,N_2915);
or U4595 (N_4595,N_2367,N_1922);
nor U4596 (N_4596,N_2369,N_1050);
nand U4597 (N_4597,N_2820,N_1794);
and U4598 (N_4598,N_1674,N_2436);
or U4599 (N_4599,N_1980,N_847);
or U4600 (N_4600,N_2787,N_2061);
and U4601 (N_4601,N_115,N_1007);
or U4602 (N_4602,N_1775,N_62);
and U4603 (N_4603,N_871,N_1421);
and U4604 (N_4604,N_1134,N_598);
and U4605 (N_4605,N_2663,N_2589);
xnor U4606 (N_4606,N_1286,N_1817);
or U4607 (N_4607,N_658,N_2228);
nand U4608 (N_4608,N_1160,N_441);
nor U4609 (N_4609,N_2228,N_2544);
or U4610 (N_4610,N_2134,N_1066);
and U4611 (N_4611,N_2866,N_2079);
nor U4612 (N_4612,N_633,N_2077);
nand U4613 (N_4613,N_2730,N_1840);
nor U4614 (N_4614,N_2446,N_1760);
and U4615 (N_4615,N_1440,N_325);
nor U4616 (N_4616,N_2835,N_389);
xnor U4617 (N_4617,N_485,N_591);
or U4618 (N_4618,N_598,N_888);
or U4619 (N_4619,N_1786,N_2300);
nand U4620 (N_4620,N_1861,N_607);
or U4621 (N_4621,N_2485,N_1126);
and U4622 (N_4622,N_2387,N_461);
or U4623 (N_4623,N_2252,N_1720);
or U4624 (N_4624,N_518,N_2622);
xor U4625 (N_4625,N_2710,N_980);
and U4626 (N_4626,N_1854,N_451);
xnor U4627 (N_4627,N_1646,N_1332);
or U4628 (N_4628,N_1866,N_2538);
and U4629 (N_4629,N_1835,N_1875);
nor U4630 (N_4630,N_2755,N_1479);
xnor U4631 (N_4631,N_2993,N_1407);
nor U4632 (N_4632,N_248,N_1533);
or U4633 (N_4633,N_2082,N_1147);
nor U4634 (N_4634,N_1873,N_1083);
xnor U4635 (N_4635,N_2502,N_2724);
nor U4636 (N_4636,N_75,N_1482);
nand U4637 (N_4637,N_2759,N_1887);
nand U4638 (N_4638,N_1640,N_2147);
xnor U4639 (N_4639,N_977,N_1810);
and U4640 (N_4640,N_1899,N_2828);
xnor U4641 (N_4641,N_2723,N_2602);
and U4642 (N_4642,N_828,N_1341);
xnor U4643 (N_4643,N_2041,N_994);
or U4644 (N_4644,N_1085,N_629);
or U4645 (N_4645,N_2073,N_2562);
nor U4646 (N_4646,N_675,N_2251);
xor U4647 (N_4647,N_1215,N_120);
xnor U4648 (N_4648,N_1923,N_1894);
nor U4649 (N_4649,N_261,N_697);
and U4650 (N_4650,N_820,N_2378);
xor U4651 (N_4651,N_2844,N_621);
nor U4652 (N_4652,N_2921,N_973);
and U4653 (N_4653,N_2436,N_299);
and U4654 (N_4654,N_2083,N_2023);
or U4655 (N_4655,N_1371,N_2856);
nand U4656 (N_4656,N_108,N_1201);
or U4657 (N_4657,N_428,N_2664);
and U4658 (N_4658,N_2474,N_960);
and U4659 (N_4659,N_1691,N_2740);
and U4660 (N_4660,N_1325,N_1844);
nand U4661 (N_4661,N_2351,N_1050);
nand U4662 (N_4662,N_2602,N_862);
xnor U4663 (N_4663,N_1596,N_251);
xnor U4664 (N_4664,N_1052,N_978);
or U4665 (N_4665,N_50,N_1867);
nand U4666 (N_4666,N_2582,N_2476);
and U4667 (N_4667,N_2038,N_2553);
and U4668 (N_4668,N_622,N_2613);
or U4669 (N_4669,N_2633,N_29);
xnor U4670 (N_4670,N_1851,N_2297);
and U4671 (N_4671,N_1975,N_2869);
xor U4672 (N_4672,N_1739,N_1760);
nand U4673 (N_4673,N_2413,N_533);
nor U4674 (N_4674,N_812,N_2946);
nor U4675 (N_4675,N_240,N_2139);
or U4676 (N_4676,N_1703,N_2486);
and U4677 (N_4677,N_1601,N_78);
nor U4678 (N_4678,N_228,N_1923);
nand U4679 (N_4679,N_1826,N_888);
nor U4680 (N_4680,N_1421,N_2801);
and U4681 (N_4681,N_2099,N_706);
nand U4682 (N_4682,N_2246,N_1189);
nand U4683 (N_4683,N_1244,N_1919);
nor U4684 (N_4684,N_1008,N_2348);
or U4685 (N_4685,N_586,N_323);
xor U4686 (N_4686,N_1820,N_2961);
xnor U4687 (N_4687,N_1324,N_1786);
nand U4688 (N_4688,N_1321,N_2998);
nand U4689 (N_4689,N_1914,N_268);
and U4690 (N_4690,N_105,N_519);
xnor U4691 (N_4691,N_1382,N_1971);
xnor U4692 (N_4692,N_2808,N_700);
or U4693 (N_4693,N_2415,N_2108);
nor U4694 (N_4694,N_664,N_266);
xor U4695 (N_4695,N_1582,N_1706);
or U4696 (N_4696,N_2315,N_1692);
or U4697 (N_4697,N_1278,N_762);
and U4698 (N_4698,N_399,N_319);
nand U4699 (N_4699,N_2486,N_526);
and U4700 (N_4700,N_2039,N_1316);
and U4701 (N_4701,N_2553,N_696);
nand U4702 (N_4702,N_2954,N_1281);
or U4703 (N_4703,N_803,N_2452);
nor U4704 (N_4704,N_2688,N_2511);
nor U4705 (N_4705,N_705,N_680);
nor U4706 (N_4706,N_1843,N_425);
xnor U4707 (N_4707,N_2049,N_1414);
nand U4708 (N_4708,N_2493,N_1177);
nor U4709 (N_4709,N_689,N_336);
nor U4710 (N_4710,N_687,N_1641);
and U4711 (N_4711,N_236,N_1745);
and U4712 (N_4712,N_464,N_684);
xor U4713 (N_4713,N_1732,N_730);
nor U4714 (N_4714,N_1745,N_1233);
nor U4715 (N_4715,N_933,N_1855);
xnor U4716 (N_4716,N_292,N_41);
nor U4717 (N_4717,N_950,N_1937);
nor U4718 (N_4718,N_2960,N_863);
or U4719 (N_4719,N_1857,N_601);
or U4720 (N_4720,N_2821,N_2605);
or U4721 (N_4721,N_1546,N_176);
and U4722 (N_4722,N_2539,N_219);
or U4723 (N_4723,N_12,N_1545);
nand U4724 (N_4724,N_2310,N_263);
nor U4725 (N_4725,N_609,N_1497);
nor U4726 (N_4726,N_529,N_1803);
nand U4727 (N_4727,N_353,N_2027);
and U4728 (N_4728,N_243,N_220);
xor U4729 (N_4729,N_1584,N_1052);
nor U4730 (N_4730,N_378,N_2379);
nand U4731 (N_4731,N_1710,N_2521);
or U4732 (N_4732,N_1264,N_2666);
and U4733 (N_4733,N_2121,N_2377);
nand U4734 (N_4734,N_1814,N_1894);
nor U4735 (N_4735,N_1754,N_1360);
xnor U4736 (N_4736,N_2149,N_1829);
xor U4737 (N_4737,N_1882,N_2262);
or U4738 (N_4738,N_271,N_7);
xor U4739 (N_4739,N_280,N_1419);
nor U4740 (N_4740,N_1251,N_828);
and U4741 (N_4741,N_894,N_264);
nor U4742 (N_4742,N_2958,N_446);
or U4743 (N_4743,N_1218,N_1652);
or U4744 (N_4744,N_749,N_2019);
xnor U4745 (N_4745,N_1752,N_1696);
xor U4746 (N_4746,N_1757,N_387);
and U4747 (N_4747,N_967,N_788);
nor U4748 (N_4748,N_755,N_2256);
nand U4749 (N_4749,N_2490,N_2225);
nand U4750 (N_4750,N_1846,N_2238);
or U4751 (N_4751,N_1559,N_379);
or U4752 (N_4752,N_2322,N_2894);
xnor U4753 (N_4753,N_678,N_2378);
or U4754 (N_4754,N_2043,N_327);
nor U4755 (N_4755,N_2159,N_2316);
nand U4756 (N_4756,N_1964,N_665);
or U4757 (N_4757,N_1211,N_1625);
or U4758 (N_4758,N_2888,N_1593);
xnor U4759 (N_4759,N_893,N_115);
or U4760 (N_4760,N_1368,N_2420);
nor U4761 (N_4761,N_75,N_291);
xnor U4762 (N_4762,N_791,N_1959);
or U4763 (N_4763,N_2574,N_1788);
and U4764 (N_4764,N_2046,N_1015);
nor U4765 (N_4765,N_2118,N_2714);
nor U4766 (N_4766,N_2593,N_2223);
nand U4767 (N_4767,N_1567,N_1934);
or U4768 (N_4768,N_2760,N_2933);
nand U4769 (N_4769,N_1225,N_1377);
nor U4770 (N_4770,N_1731,N_384);
xnor U4771 (N_4771,N_902,N_618);
and U4772 (N_4772,N_328,N_2834);
xnor U4773 (N_4773,N_2286,N_589);
nor U4774 (N_4774,N_1338,N_1097);
xnor U4775 (N_4775,N_1839,N_966);
nor U4776 (N_4776,N_2312,N_2180);
xor U4777 (N_4777,N_1901,N_1518);
and U4778 (N_4778,N_890,N_508);
or U4779 (N_4779,N_404,N_2137);
nand U4780 (N_4780,N_2212,N_1806);
and U4781 (N_4781,N_518,N_1771);
or U4782 (N_4782,N_1390,N_2856);
nor U4783 (N_4783,N_679,N_63);
nand U4784 (N_4784,N_1611,N_2634);
or U4785 (N_4785,N_940,N_2121);
or U4786 (N_4786,N_278,N_2693);
nor U4787 (N_4787,N_527,N_1009);
or U4788 (N_4788,N_1773,N_2177);
and U4789 (N_4789,N_2585,N_285);
nand U4790 (N_4790,N_2588,N_2716);
and U4791 (N_4791,N_1170,N_1607);
xor U4792 (N_4792,N_2765,N_1095);
and U4793 (N_4793,N_571,N_2581);
xnor U4794 (N_4794,N_2656,N_1299);
and U4795 (N_4795,N_2791,N_1027);
and U4796 (N_4796,N_468,N_1796);
or U4797 (N_4797,N_647,N_774);
xor U4798 (N_4798,N_899,N_7);
and U4799 (N_4799,N_2591,N_1395);
xnor U4800 (N_4800,N_1114,N_2086);
and U4801 (N_4801,N_1023,N_409);
and U4802 (N_4802,N_2101,N_840);
xnor U4803 (N_4803,N_1577,N_1512);
nor U4804 (N_4804,N_2436,N_1270);
xnor U4805 (N_4805,N_2319,N_1831);
or U4806 (N_4806,N_2131,N_2694);
xnor U4807 (N_4807,N_1662,N_2834);
nand U4808 (N_4808,N_2187,N_1437);
nand U4809 (N_4809,N_33,N_596);
xnor U4810 (N_4810,N_17,N_2539);
xor U4811 (N_4811,N_494,N_1182);
or U4812 (N_4812,N_1363,N_44);
or U4813 (N_4813,N_856,N_420);
nor U4814 (N_4814,N_309,N_2553);
nand U4815 (N_4815,N_1945,N_1396);
or U4816 (N_4816,N_1288,N_2279);
and U4817 (N_4817,N_1119,N_2674);
xnor U4818 (N_4818,N_2822,N_1280);
nor U4819 (N_4819,N_2306,N_1960);
nor U4820 (N_4820,N_2252,N_2647);
nor U4821 (N_4821,N_2092,N_196);
or U4822 (N_4822,N_2390,N_737);
nor U4823 (N_4823,N_856,N_2594);
or U4824 (N_4824,N_19,N_1038);
or U4825 (N_4825,N_1204,N_435);
or U4826 (N_4826,N_2983,N_2297);
nor U4827 (N_4827,N_461,N_204);
or U4828 (N_4828,N_2823,N_734);
nor U4829 (N_4829,N_1102,N_429);
xnor U4830 (N_4830,N_2220,N_159);
nor U4831 (N_4831,N_1667,N_1983);
nor U4832 (N_4832,N_2785,N_368);
or U4833 (N_4833,N_2661,N_2513);
or U4834 (N_4834,N_1982,N_1176);
or U4835 (N_4835,N_979,N_1874);
or U4836 (N_4836,N_117,N_2189);
or U4837 (N_4837,N_58,N_473);
nand U4838 (N_4838,N_1160,N_1139);
xor U4839 (N_4839,N_519,N_1708);
nand U4840 (N_4840,N_2500,N_532);
nor U4841 (N_4841,N_588,N_644);
xor U4842 (N_4842,N_1374,N_71);
nor U4843 (N_4843,N_2720,N_1674);
and U4844 (N_4844,N_280,N_177);
or U4845 (N_4845,N_1058,N_2624);
nor U4846 (N_4846,N_933,N_2510);
xnor U4847 (N_4847,N_2535,N_1136);
nor U4848 (N_4848,N_1936,N_794);
and U4849 (N_4849,N_836,N_2584);
or U4850 (N_4850,N_1077,N_1226);
nor U4851 (N_4851,N_1653,N_1712);
and U4852 (N_4852,N_1179,N_1208);
nor U4853 (N_4853,N_2325,N_1077);
nand U4854 (N_4854,N_1895,N_2756);
xnor U4855 (N_4855,N_1870,N_2009);
nor U4856 (N_4856,N_505,N_455);
nand U4857 (N_4857,N_1254,N_2863);
xnor U4858 (N_4858,N_2983,N_2612);
or U4859 (N_4859,N_1932,N_478);
nand U4860 (N_4860,N_2284,N_1682);
or U4861 (N_4861,N_1972,N_1083);
xor U4862 (N_4862,N_159,N_750);
or U4863 (N_4863,N_2239,N_2138);
xnor U4864 (N_4864,N_2078,N_41);
and U4865 (N_4865,N_863,N_2294);
or U4866 (N_4866,N_1099,N_2962);
nand U4867 (N_4867,N_304,N_821);
and U4868 (N_4868,N_7,N_645);
xnor U4869 (N_4869,N_2931,N_2318);
xor U4870 (N_4870,N_580,N_1420);
nor U4871 (N_4871,N_1998,N_2235);
xor U4872 (N_4872,N_802,N_1548);
xnor U4873 (N_4873,N_2104,N_1968);
nor U4874 (N_4874,N_1119,N_2724);
nor U4875 (N_4875,N_744,N_239);
or U4876 (N_4876,N_21,N_750);
and U4877 (N_4877,N_2932,N_2974);
nand U4878 (N_4878,N_1612,N_1874);
nor U4879 (N_4879,N_2874,N_2043);
nand U4880 (N_4880,N_2370,N_2905);
nand U4881 (N_4881,N_650,N_1519);
xor U4882 (N_4882,N_2754,N_2766);
nand U4883 (N_4883,N_1762,N_1494);
or U4884 (N_4884,N_57,N_802);
and U4885 (N_4885,N_2843,N_2256);
xnor U4886 (N_4886,N_1905,N_2082);
xnor U4887 (N_4887,N_941,N_2447);
and U4888 (N_4888,N_2265,N_2702);
and U4889 (N_4889,N_1496,N_2445);
and U4890 (N_4890,N_2567,N_2647);
and U4891 (N_4891,N_1764,N_1370);
nor U4892 (N_4892,N_2667,N_1117);
xnor U4893 (N_4893,N_2313,N_2217);
and U4894 (N_4894,N_2244,N_2324);
or U4895 (N_4895,N_664,N_876);
and U4896 (N_4896,N_1173,N_743);
nand U4897 (N_4897,N_1843,N_1370);
xnor U4898 (N_4898,N_385,N_1703);
xnor U4899 (N_4899,N_2883,N_1457);
or U4900 (N_4900,N_2794,N_2174);
xnor U4901 (N_4901,N_2889,N_1888);
and U4902 (N_4902,N_1982,N_2257);
or U4903 (N_4903,N_2051,N_1234);
or U4904 (N_4904,N_2854,N_224);
nand U4905 (N_4905,N_475,N_1759);
nand U4906 (N_4906,N_578,N_846);
or U4907 (N_4907,N_1699,N_2910);
nand U4908 (N_4908,N_2257,N_2714);
and U4909 (N_4909,N_2926,N_1890);
xnor U4910 (N_4910,N_1041,N_2337);
nand U4911 (N_4911,N_915,N_1554);
or U4912 (N_4912,N_2378,N_2707);
xor U4913 (N_4913,N_2757,N_2825);
or U4914 (N_4914,N_2783,N_2679);
or U4915 (N_4915,N_1123,N_2188);
or U4916 (N_4916,N_1049,N_1224);
or U4917 (N_4917,N_1830,N_1637);
xor U4918 (N_4918,N_1573,N_870);
nor U4919 (N_4919,N_1755,N_24);
xnor U4920 (N_4920,N_1212,N_740);
nor U4921 (N_4921,N_466,N_629);
or U4922 (N_4922,N_633,N_2635);
and U4923 (N_4923,N_1504,N_2901);
or U4924 (N_4924,N_663,N_1890);
or U4925 (N_4925,N_2476,N_2357);
xnor U4926 (N_4926,N_2471,N_1351);
xnor U4927 (N_4927,N_557,N_2725);
nor U4928 (N_4928,N_122,N_1223);
nor U4929 (N_4929,N_245,N_2330);
nor U4930 (N_4930,N_662,N_1444);
nor U4931 (N_4931,N_2689,N_2888);
xor U4932 (N_4932,N_132,N_236);
or U4933 (N_4933,N_2232,N_2142);
or U4934 (N_4934,N_989,N_441);
nand U4935 (N_4935,N_224,N_2598);
nor U4936 (N_4936,N_801,N_1224);
and U4937 (N_4937,N_290,N_2134);
nor U4938 (N_4938,N_2591,N_777);
and U4939 (N_4939,N_414,N_1315);
and U4940 (N_4940,N_576,N_694);
nor U4941 (N_4941,N_2431,N_854);
or U4942 (N_4942,N_2285,N_2809);
and U4943 (N_4943,N_29,N_422);
and U4944 (N_4944,N_2542,N_2765);
xor U4945 (N_4945,N_1291,N_1244);
or U4946 (N_4946,N_1515,N_1486);
or U4947 (N_4947,N_1202,N_788);
nor U4948 (N_4948,N_1268,N_2945);
nor U4949 (N_4949,N_2142,N_1423);
nor U4950 (N_4950,N_1741,N_604);
nand U4951 (N_4951,N_2461,N_2869);
and U4952 (N_4952,N_1314,N_604);
xnor U4953 (N_4953,N_1166,N_2140);
nor U4954 (N_4954,N_1258,N_2769);
xor U4955 (N_4955,N_503,N_1160);
nor U4956 (N_4956,N_2333,N_2671);
nand U4957 (N_4957,N_1794,N_2292);
nor U4958 (N_4958,N_22,N_341);
nor U4959 (N_4959,N_2911,N_1699);
and U4960 (N_4960,N_2709,N_1532);
or U4961 (N_4961,N_1862,N_25);
nor U4962 (N_4962,N_510,N_310);
nor U4963 (N_4963,N_2834,N_2294);
or U4964 (N_4964,N_306,N_1720);
nand U4965 (N_4965,N_2368,N_1800);
and U4966 (N_4966,N_2646,N_804);
or U4967 (N_4967,N_52,N_47);
and U4968 (N_4968,N_204,N_794);
nor U4969 (N_4969,N_179,N_2918);
nand U4970 (N_4970,N_1512,N_760);
or U4971 (N_4971,N_607,N_633);
nor U4972 (N_4972,N_1768,N_2661);
xnor U4973 (N_4973,N_2785,N_2664);
and U4974 (N_4974,N_1791,N_2405);
or U4975 (N_4975,N_2338,N_659);
or U4976 (N_4976,N_2933,N_286);
or U4977 (N_4977,N_2887,N_84);
nor U4978 (N_4978,N_2557,N_2256);
and U4979 (N_4979,N_679,N_781);
or U4980 (N_4980,N_2192,N_2779);
xnor U4981 (N_4981,N_218,N_357);
and U4982 (N_4982,N_369,N_2928);
and U4983 (N_4983,N_2526,N_2836);
nand U4984 (N_4984,N_484,N_2874);
and U4985 (N_4985,N_2914,N_2225);
or U4986 (N_4986,N_1153,N_2786);
and U4987 (N_4987,N_2420,N_827);
xnor U4988 (N_4988,N_2509,N_652);
nand U4989 (N_4989,N_501,N_386);
nor U4990 (N_4990,N_2676,N_634);
xnor U4991 (N_4991,N_1945,N_1440);
xnor U4992 (N_4992,N_2374,N_2478);
or U4993 (N_4993,N_2502,N_1393);
and U4994 (N_4994,N_821,N_84);
nor U4995 (N_4995,N_2323,N_2154);
nor U4996 (N_4996,N_1035,N_8);
and U4997 (N_4997,N_1640,N_2209);
nand U4998 (N_4998,N_121,N_1153);
nor U4999 (N_4999,N_2551,N_642);
xor U5000 (N_5000,N_2744,N_596);
or U5001 (N_5001,N_2243,N_211);
nor U5002 (N_5002,N_2412,N_2258);
and U5003 (N_5003,N_2260,N_2930);
nand U5004 (N_5004,N_615,N_1305);
and U5005 (N_5005,N_421,N_911);
and U5006 (N_5006,N_2144,N_314);
and U5007 (N_5007,N_1608,N_776);
and U5008 (N_5008,N_2012,N_75);
nand U5009 (N_5009,N_426,N_1248);
nand U5010 (N_5010,N_1500,N_2070);
nor U5011 (N_5011,N_227,N_1890);
nor U5012 (N_5012,N_2556,N_1079);
xor U5013 (N_5013,N_2287,N_1144);
nand U5014 (N_5014,N_2972,N_1960);
and U5015 (N_5015,N_692,N_2070);
or U5016 (N_5016,N_585,N_2089);
and U5017 (N_5017,N_231,N_203);
xnor U5018 (N_5018,N_2256,N_777);
or U5019 (N_5019,N_2121,N_1670);
or U5020 (N_5020,N_1781,N_2899);
nor U5021 (N_5021,N_2378,N_1449);
nand U5022 (N_5022,N_2373,N_2375);
and U5023 (N_5023,N_2227,N_355);
xnor U5024 (N_5024,N_273,N_374);
or U5025 (N_5025,N_776,N_971);
and U5026 (N_5026,N_1823,N_799);
xor U5027 (N_5027,N_2127,N_1683);
xnor U5028 (N_5028,N_2768,N_171);
or U5029 (N_5029,N_2703,N_2042);
or U5030 (N_5030,N_1073,N_1481);
nor U5031 (N_5031,N_963,N_2587);
nand U5032 (N_5032,N_1376,N_2706);
and U5033 (N_5033,N_1985,N_1746);
and U5034 (N_5034,N_2316,N_2307);
xor U5035 (N_5035,N_363,N_1319);
or U5036 (N_5036,N_2250,N_1652);
xnor U5037 (N_5037,N_2980,N_278);
and U5038 (N_5038,N_2648,N_1786);
nand U5039 (N_5039,N_686,N_2673);
and U5040 (N_5040,N_411,N_2902);
and U5041 (N_5041,N_1883,N_1001);
nor U5042 (N_5042,N_2263,N_931);
nor U5043 (N_5043,N_232,N_1997);
and U5044 (N_5044,N_1846,N_2540);
xnor U5045 (N_5045,N_1146,N_114);
nor U5046 (N_5046,N_212,N_2781);
and U5047 (N_5047,N_1550,N_2143);
xnor U5048 (N_5048,N_2863,N_1004);
xnor U5049 (N_5049,N_1366,N_1635);
nand U5050 (N_5050,N_875,N_772);
xnor U5051 (N_5051,N_593,N_651);
xnor U5052 (N_5052,N_2995,N_85);
or U5053 (N_5053,N_1147,N_968);
nand U5054 (N_5054,N_2847,N_2551);
and U5055 (N_5055,N_2241,N_1492);
and U5056 (N_5056,N_2717,N_2755);
or U5057 (N_5057,N_233,N_82);
xor U5058 (N_5058,N_2811,N_2149);
nand U5059 (N_5059,N_1469,N_1496);
nand U5060 (N_5060,N_1890,N_1358);
nand U5061 (N_5061,N_2052,N_2513);
and U5062 (N_5062,N_2187,N_2258);
xor U5063 (N_5063,N_2654,N_110);
and U5064 (N_5064,N_757,N_1129);
xor U5065 (N_5065,N_1102,N_1241);
and U5066 (N_5066,N_2968,N_1953);
or U5067 (N_5067,N_2378,N_739);
xor U5068 (N_5068,N_1254,N_304);
nand U5069 (N_5069,N_2216,N_1140);
nor U5070 (N_5070,N_2619,N_1447);
nand U5071 (N_5071,N_2293,N_1362);
nand U5072 (N_5072,N_2216,N_1399);
nor U5073 (N_5073,N_2141,N_1125);
and U5074 (N_5074,N_2912,N_1120);
or U5075 (N_5075,N_1604,N_2287);
xor U5076 (N_5076,N_2569,N_1077);
xor U5077 (N_5077,N_2083,N_1587);
or U5078 (N_5078,N_2715,N_2083);
xor U5079 (N_5079,N_2271,N_2047);
nor U5080 (N_5080,N_1971,N_2017);
xor U5081 (N_5081,N_2447,N_2295);
nand U5082 (N_5082,N_581,N_2417);
and U5083 (N_5083,N_2525,N_688);
or U5084 (N_5084,N_392,N_2921);
xnor U5085 (N_5085,N_838,N_1090);
xnor U5086 (N_5086,N_485,N_376);
nor U5087 (N_5087,N_759,N_2837);
xnor U5088 (N_5088,N_797,N_1617);
xnor U5089 (N_5089,N_151,N_679);
xnor U5090 (N_5090,N_2588,N_2814);
nor U5091 (N_5091,N_1231,N_2261);
or U5092 (N_5092,N_2453,N_2216);
nand U5093 (N_5093,N_2287,N_1594);
nand U5094 (N_5094,N_2460,N_1035);
or U5095 (N_5095,N_2406,N_613);
xor U5096 (N_5096,N_1872,N_1377);
nand U5097 (N_5097,N_962,N_2801);
or U5098 (N_5098,N_906,N_519);
xnor U5099 (N_5099,N_1595,N_812);
nand U5100 (N_5100,N_464,N_2254);
nor U5101 (N_5101,N_567,N_1717);
xnor U5102 (N_5102,N_2939,N_2397);
xor U5103 (N_5103,N_2083,N_174);
or U5104 (N_5104,N_2413,N_1141);
xor U5105 (N_5105,N_510,N_613);
and U5106 (N_5106,N_644,N_1324);
xnor U5107 (N_5107,N_996,N_539);
xnor U5108 (N_5108,N_1680,N_729);
and U5109 (N_5109,N_1066,N_1470);
and U5110 (N_5110,N_1034,N_652);
nor U5111 (N_5111,N_2293,N_876);
or U5112 (N_5112,N_1571,N_1951);
nor U5113 (N_5113,N_148,N_2026);
nor U5114 (N_5114,N_2587,N_1943);
xnor U5115 (N_5115,N_882,N_1240);
or U5116 (N_5116,N_342,N_1115);
or U5117 (N_5117,N_2972,N_2390);
xor U5118 (N_5118,N_781,N_218);
nor U5119 (N_5119,N_2234,N_2154);
xnor U5120 (N_5120,N_102,N_295);
and U5121 (N_5121,N_2284,N_1680);
or U5122 (N_5122,N_36,N_920);
nor U5123 (N_5123,N_2570,N_2033);
or U5124 (N_5124,N_2044,N_419);
and U5125 (N_5125,N_1691,N_943);
or U5126 (N_5126,N_2585,N_1576);
or U5127 (N_5127,N_1061,N_1241);
or U5128 (N_5128,N_967,N_67);
nand U5129 (N_5129,N_650,N_2562);
nand U5130 (N_5130,N_2979,N_1957);
xnor U5131 (N_5131,N_2843,N_2065);
and U5132 (N_5132,N_846,N_2292);
or U5133 (N_5133,N_2708,N_969);
and U5134 (N_5134,N_1748,N_508);
nor U5135 (N_5135,N_28,N_2899);
and U5136 (N_5136,N_2113,N_2227);
nor U5137 (N_5137,N_2627,N_843);
nand U5138 (N_5138,N_69,N_1027);
nor U5139 (N_5139,N_425,N_19);
or U5140 (N_5140,N_1778,N_163);
nand U5141 (N_5141,N_2447,N_1979);
xor U5142 (N_5142,N_2883,N_2067);
xor U5143 (N_5143,N_1675,N_2407);
nor U5144 (N_5144,N_1395,N_1480);
nand U5145 (N_5145,N_99,N_2837);
and U5146 (N_5146,N_1690,N_534);
xor U5147 (N_5147,N_1207,N_2329);
nand U5148 (N_5148,N_2461,N_2799);
xnor U5149 (N_5149,N_301,N_1425);
and U5150 (N_5150,N_1144,N_1855);
and U5151 (N_5151,N_1771,N_1327);
nand U5152 (N_5152,N_2231,N_2706);
and U5153 (N_5153,N_136,N_1008);
nand U5154 (N_5154,N_775,N_2004);
nand U5155 (N_5155,N_356,N_441);
nand U5156 (N_5156,N_839,N_2873);
nor U5157 (N_5157,N_1452,N_875);
nor U5158 (N_5158,N_2683,N_313);
and U5159 (N_5159,N_2485,N_2924);
nand U5160 (N_5160,N_726,N_46);
xor U5161 (N_5161,N_1678,N_741);
xor U5162 (N_5162,N_1554,N_1440);
and U5163 (N_5163,N_891,N_1940);
and U5164 (N_5164,N_1907,N_1788);
or U5165 (N_5165,N_2018,N_2272);
and U5166 (N_5166,N_2820,N_842);
or U5167 (N_5167,N_1364,N_2194);
and U5168 (N_5168,N_37,N_1447);
and U5169 (N_5169,N_1531,N_108);
or U5170 (N_5170,N_769,N_788);
and U5171 (N_5171,N_1372,N_2654);
and U5172 (N_5172,N_420,N_351);
nor U5173 (N_5173,N_818,N_1365);
xor U5174 (N_5174,N_1024,N_1252);
and U5175 (N_5175,N_1327,N_2586);
and U5176 (N_5176,N_177,N_1893);
xor U5177 (N_5177,N_2718,N_1559);
xor U5178 (N_5178,N_2720,N_1844);
or U5179 (N_5179,N_2639,N_2460);
or U5180 (N_5180,N_547,N_1341);
and U5181 (N_5181,N_1427,N_2623);
and U5182 (N_5182,N_2211,N_2196);
nor U5183 (N_5183,N_1158,N_309);
nand U5184 (N_5184,N_2440,N_2185);
xor U5185 (N_5185,N_1280,N_2147);
or U5186 (N_5186,N_440,N_1079);
and U5187 (N_5187,N_1539,N_1034);
or U5188 (N_5188,N_1552,N_272);
xnor U5189 (N_5189,N_1891,N_517);
or U5190 (N_5190,N_777,N_1540);
nand U5191 (N_5191,N_1159,N_444);
and U5192 (N_5192,N_1732,N_372);
or U5193 (N_5193,N_690,N_553);
nor U5194 (N_5194,N_488,N_930);
or U5195 (N_5195,N_2874,N_1482);
nor U5196 (N_5196,N_774,N_2163);
or U5197 (N_5197,N_519,N_735);
nand U5198 (N_5198,N_2852,N_1074);
xor U5199 (N_5199,N_1372,N_1467);
nand U5200 (N_5200,N_2510,N_2364);
and U5201 (N_5201,N_383,N_1314);
or U5202 (N_5202,N_1741,N_699);
and U5203 (N_5203,N_2155,N_1912);
nand U5204 (N_5204,N_43,N_1894);
nor U5205 (N_5205,N_1878,N_335);
nor U5206 (N_5206,N_505,N_1327);
and U5207 (N_5207,N_959,N_1164);
nand U5208 (N_5208,N_2697,N_156);
nor U5209 (N_5209,N_190,N_2485);
nor U5210 (N_5210,N_1832,N_1581);
xor U5211 (N_5211,N_1523,N_159);
or U5212 (N_5212,N_353,N_1746);
xnor U5213 (N_5213,N_925,N_1071);
or U5214 (N_5214,N_2170,N_2755);
xor U5215 (N_5215,N_109,N_2470);
nor U5216 (N_5216,N_1717,N_2621);
and U5217 (N_5217,N_461,N_2844);
or U5218 (N_5218,N_995,N_563);
or U5219 (N_5219,N_1944,N_967);
xnor U5220 (N_5220,N_717,N_1022);
nand U5221 (N_5221,N_1129,N_1603);
xnor U5222 (N_5222,N_2622,N_1819);
nor U5223 (N_5223,N_2606,N_26);
xnor U5224 (N_5224,N_2364,N_2571);
or U5225 (N_5225,N_623,N_112);
xnor U5226 (N_5226,N_1534,N_552);
xnor U5227 (N_5227,N_1514,N_2581);
xnor U5228 (N_5228,N_2922,N_973);
xnor U5229 (N_5229,N_1472,N_748);
nor U5230 (N_5230,N_596,N_129);
nand U5231 (N_5231,N_477,N_1267);
nor U5232 (N_5232,N_463,N_864);
nor U5233 (N_5233,N_1831,N_2534);
and U5234 (N_5234,N_1780,N_830);
nand U5235 (N_5235,N_1024,N_2875);
nor U5236 (N_5236,N_1135,N_2319);
or U5237 (N_5237,N_1454,N_1716);
nor U5238 (N_5238,N_790,N_2594);
or U5239 (N_5239,N_1830,N_2025);
and U5240 (N_5240,N_675,N_2065);
xor U5241 (N_5241,N_1764,N_1911);
nand U5242 (N_5242,N_2029,N_255);
and U5243 (N_5243,N_589,N_1060);
or U5244 (N_5244,N_2146,N_913);
nor U5245 (N_5245,N_2085,N_128);
nor U5246 (N_5246,N_97,N_84);
xor U5247 (N_5247,N_1899,N_741);
nor U5248 (N_5248,N_2305,N_2230);
xor U5249 (N_5249,N_847,N_2695);
nand U5250 (N_5250,N_234,N_191);
nand U5251 (N_5251,N_9,N_2722);
nor U5252 (N_5252,N_2147,N_2071);
or U5253 (N_5253,N_2257,N_533);
and U5254 (N_5254,N_1,N_2298);
nand U5255 (N_5255,N_1519,N_2040);
and U5256 (N_5256,N_1117,N_1828);
and U5257 (N_5257,N_104,N_1882);
or U5258 (N_5258,N_1341,N_2891);
nand U5259 (N_5259,N_2864,N_2107);
xnor U5260 (N_5260,N_1192,N_2445);
and U5261 (N_5261,N_322,N_2362);
nand U5262 (N_5262,N_753,N_2650);
and U5263 (N_5263,N_1716,N_1554);
xnor U5264 (N_5264,N_2666,N_2147);
nor U5265 (N_5265,N_587,N_758);
nand U5266 (N_5266,N_346,N_2925);
or U5267 (N_5267,N_1089,N_2215);
nor U5268 (N_5268,N_834,N_2092);
or U5269 (N_5269,N_575,N_424);
nand U5270 (N_5270,N_164,N_1425);
xor U5271 (N_5271,N_2701,N_888);
and U5272 (N_5272,N_2717,N_2999);
xor U5273 (N_5273,N_3,N_1337);
nand U5274 (N_5274,N_2422,N_2103);
and U5275 (N_5275,N_1909,N_1306);
nand U5276 (N_5276,N_1870,N_1320);
nor U5277 (N_5277,N_1853,N_2545);
nor U5278 (N_5278,N_1432,N_494);
nor U5279 (N_5279,N_2253,N_815);
and U5280 (N_5280,N_469,N_195);
xnor U5281 (N_5281,N_2350,N_1688);
nand U5282 (N_5282,N_2158,N_1910);
and U5283 (N_5283,N_1701,N_1051);
and U5284 (N_5284,N_157,N_1373);
xnor U5285 (N_5285,N_390,N_1060);
nor U5286 (N_5286,N_621,N_1501);
nand U5287 (N_5287,N_2380,N_2221);
xnor U5288 (N_5288,N_2290,N_1865);
nor U5289 (N_5289,N_491,N_580);
and U5290 (N_5290,N_2460,N_1578);
or U5291 (N_5291,N_1460,N_2667);
and U5292 (N_5292,N_1153,N_1424);
and U5293 (N_5293,N_2593,N_1746);
nand U5294 (N_5294,N_1067,N_2951);
and U5295 (N_5295,N_2508,N_1779);
xor U5296 (N_5296,N_807,N_636);
nand U5297 (N_5297,N_2924,N_612);
xor U5298 (N_5298,N_974,N_976);
and U5299 (N_5299,N_2086,N_2883);
or U5300 (N_5300,N_2578,N_687);
xor U5301 (N_5301,N_1066,N_2629);
and U5302 (N_5302,N_1467,N_1090);
nor U5303 (N_5303,N_2800,N_795);
or U5304 (N_5304,N_685,N_849);
and U5305 (N_5305,N_2724,N_1263);
nor U5306 (N_5306,N_796,N_2465);
xor U5307 (N_5307,N_2528,N_923);
nand U5308 (N_5308,N_1693,N_180);
or U5309 (N_5309,N_2947,N_1335);
and U5310 (N_5310,N_1721,N_2002);
nor U5311 (N_5311,N_1025,N_308);
nor U5312 (N_5312,N_2306,N_1165);
and U5313 (N_5313,N_595,N_368);
nor U5314 (N_5314,N_339,N_1482);
or U5315 (N_5315,N_1793,N_1154);
nand U5316 (N_5316,N_232,N_2335);
xnor U5317 (N_5317,N_881,N_1373);
xnor U5318 (N_5318,N_1883,N_2660);
nor U5319 (N_5319,N_2879,N_1051);
nor U5320 (N_5320,N_2751,N_2714);
xnor U5321 (N_5321,N_144,N_993);
xor U5322 (N_5322,N_2408,N_863);
nand U5323 (N_5323,N_1776,N_2850);
nand U5324 (N_5324,N_1323,N_2061);
nor U5325 (N_5325,N_1871,N_227);
and U5326 (N_5326,N_2719,N_1127);
or U5327 (N_5327,N_2247,N_1846);
and U5328 (N_5328,N_1498,N_2701);
nor U5329 (N_5329,N_2420,N_2402);
and U5330 (N_5330,N_1025,N_2382);
xor U5331 (N_5331,N_2066,N_2094);
nand U5332 (N_5332,N_2224,N_2180);
nor U5333 (N_5333,N_984,N_2955);
xor U5334 (N_5334,N_137,N_488);
xor U5335 (N_5335,N_1137,N_884);
nand U5336 (N_5336,N_1092,N_2294);
or U5337 (N_5337,N_2273,N_663);
and U5338 (N_5338,N_1977,N_669);
or U5339 (N_5339,N_1144,N_1928);
and U5340 (N_5340,N_2030,N_693);
nand U5341 (N_5341,N_51,N_1563);
xnor U5342 (N_5342,N_1923,N_66);
nand U5343 (N_5343,N_2665,N_2082);
and U5344 (N_5344,N_48,N_533);
xnor U5345 (N_5345,N_2916,N_124);
nor U5346 (N_5346,N_2144,N_1207);
xnor U5347 (N_5347,N_1827,N_1313);
nor U5348 (N_5348,N_1937,N_1723);
or U5349 (N_5349,N_2424,N_929);
xnor U5350 (N_5350,N_2505,N_2161);
or U5351 (N_5351,N_2828,N_2461);
or U5352 (N_5352,N_955,N_1480);
or U5353 (N_5353,N_513,N_18);
xor U5354 (N_5354,N_804,N_2686);
xnor U5355 (N_5355,N_1294,N_1851);
or U5356 (N_5356,N_1682,N_533);
and U5357 (N_5357,N_2157,N_1127);
nand U5358 (N_5358,N_394,N_2518);
and U5359 (N_5359,N_997,N_699);
nor U5360 (N_5360,N_1472,N_255);
xor U5361 (N_5361,N_2276,N_837);
and U5362 (N_5362,N_544,N_1789);
xor U5363 (N_5363,N_990,N_2129);
or U5364 (N_5364,N_2221,N_1258);
or U5365 (N_5365,N_2673,N_2166);
and U5366 (N_5366,N_783,N_1927);
or U5367 (N_5367,N_658,N_2858);
nor U5368 (N_5368,N_1260,N_1478);
nand U5369 (N_5369,N_1392,N_2581);
xnor U5370 (N_5370,N_2964,N_780);
and U5371 (N_5371,N_278,N_1204);
xnor U5372 (N_5372,N_1380,N_2469);
xnor U5373 (N_5373,N_870,N_1312);
and U5374 (N_5374,N_2649,N_2585);
xnor U5375 (N_5375,N_671,N_2041);
xor U5376 (N_5376,N_1110,N_491);
nand U5377 (N_5377,N_1645,N_104);
or U5378 (N_5378,N_2731,N_2722);
xnor U5379 (N_5379,N_271,N_163);
and U5380 (N_5380,N_2529,N_2528);
nand U5381 (N_5381,N_1911,N_644);
xnor U5382 (N_5382,N_1734,N_241);
nor U5383 (N_5383,N_2082,N_531);
nand U5384 (N_5384,N_1783,N_1299);
xor U5385 (N_5385,N_2454,N_2101);
xor U5386 (N_5386,N_618,N_2659);
or U5387 (N_5387,N_2396,N_949);
nand U5388 (N_5388,N_2002,N_2797);
nor U5389 (N_5389,N_2543,N_332);
nand U5390 (N_5390,N_1018,N_324);
xor U5391 (N_5391,N_1898,N_1046);
and U5392 (N_5392,N_1847,N_2486);
nor U5393 (N_5393,N_2854,N_2776);
nor U5394 (N_5394,N_1147,N_92);
xnor U5395 (N_5395,N_1598,N_1101);
nor U5396 (N_5396,N_582,N_1339);
or U5397 (N_5397,N_1755,N_1005);
or U5398 (N_5398,N_1677,N_929);
xnor U5399 (N_5399,N_1084,N_1923);
nand U5400 (N_5400,N_1115,N_1907);
and U5401 (N_5401,N_364,N_2193);
and U5402 (N_5402,N_1210,N_2993);
nor U5403 (N_5403,N_155,N_1398);
and U5404 (N_5404,N_1262,N_427);
and U5405 (N_5405,N_2308,N_1516);
nor U5406 (N_5406,N_870,N_1867);
nor U5407 (N_5407,N_1142,N_1579);
nor U5408 (N_5408,N_2918,N_1980);
nor U5409 (N_5409,N_1541,N_87);
xor U5410 (N_5410,N_319,N_2235);
nand U5411 (N_5411,N_499,N_1693);
xnor U5412 (N_5412,N_1405,N_1977);
nand U5413 (N_5413,N_341,N_1309);
xor U5414 (N_5414,N_552,N_42);
or U5415 (N_5415,N_191,N_410);
nand U5416 (N_5416,N_2083,N_2493);
nor U5417 (N_5417,N_1944,N_2133);
or U5418 (N_5418,N_579,N_2388);
xor U5419 (N_5419,N_2758,N_2763);
or U5420 (N_5420,N_322,N_323);
xor U5421 (N_5421,N_2772,N_395);
xnor U5422 (N_5422,N_1035,N_531);
and U5423 (N_5423,N_2479,N_373);
nor U5424 (N_5424,N_1445,N_166);
xor U5425 (N_5425,N_1214,N_2306);
or U5426 (N_5426,N_228,N_1541);
nor U5427 (N_5427,N_407,N_1012);
xnor U5428 (N_5428,N_1837,N_1163);
and U5429 (N_5429,N_505,N_1530);
nand U5430 (N_5430,N_2707,N_1581);
nand U5431 (N_5431,N_161,N_260);
nor U5432 (N_5432,N_1235,N_812);
or U5433 (N_5433,N_2077,N_1952);
or U5434 (N_5434,N_740,N_848);
and U5435 (N_5435,N_2929,N_2979);
and U5436 (N_5436,N_2690,N_2260);
nor U5437 (N_5437,N_2634,N_981);
nand U5438 (N_5438,N_260,N_1635);
or U5439 (N_5439,N_2888,N_1558);
nor U5440 (N_5440,N_706,N_2805);
nor U5441 (N_5441,N_1397,N_2501);
nor U5442 (N_5442,N_2568,N_577);
or U5443 (N_5443,N_1437,N_407);
and U5444 (N_5444,N_2044,N_692);
or U5445 (N_5445,N_1418,N_242);
nor U5446 (N_5446,N_1157,N_706);
nand U5447 (N_5447,N_2756,N_1189);
nor U5448 (N_5448,N_2997,N_729);
nand U5449 (N_5449,N_1756,N_2591);
nand U5450 (N_5450,N_2471,N_603);
nor U5451 (N_5451,N_667,N_135);
and U5452 (N_5452,N_2720,N_2422);
or U5453 (N_5453,N_2160,N_2814);
xor U5454 (N_5454,N_2861,N_727);
or U5455 (N_5455,N_2179,N_1507);
nor U5456 (N_5456,N_460,N_2206);
xnor U5457 (N_5457,N_2583,N_2003);
or U5458 (N_5458,N_9,N_1481);
xor U5459 (N_5459,N_2841,N_1988);
nand U5460 (N_5460,N_857,N_20);
and U5461 (N_5461,N_970,N_1840);
nand U5462 (N_5462,N_2852,N_789);
xor U5463 (N_5463,N_2920,N_1);
nor U5464 (N_5464,N_251,N_185);
and U5465 (N_5465,N_644,N_2223);
nand U5466 (N_5466,N_1990,N_1052);
and U5467 (N_5467,N_1995,N_1637);
xor U5468 (N_5468,N_767,N_2429);
xnor U5469 (N_5469,N_767,N_1774);
or U5470 (N_5470,N_2041,N_987);
xnor U5471 (N_5471,N_674,N_2809);
or U5472 (N_5472,N_2691,N_2038);
nor U5473 (N_5473,N_139,N_1327);
nand U5474 (N_5474,N_2091,N_1342);
or U5475 (N_5475,N_2876,N_2073);
and U5476 (N_5476,N_2629,N_1054);
xnor U5477 (N_5477,N_2754,N_1623);
nand U5478 (N_5478,N_2491,N_2180);
nand U5479 (N_5479,N_2386,N_2508);
nor U5480 (N_5480,N_2254,N_923);
nand U5481 (N_5481,N_199,N_2770);
nand U5482 (N_5482,N_2439,N_564);
xor U5483 (N_5483,N_1681,N_1786);
nand U5484 (N_5484,N_1443,N_773);
nor U5485 (N_5485,N_255,N_182);
and U5486 (N_5486,N_361,N_2550);
and U5487 (N_5487,N_582,N_2003);
nand U5488 (N_5488,N_947,N_999);
and U5489 (N_5489,N_1287,N_1687);
or U5490 (N_5490,N_1587,N_150);
or U5491 (N_5491,N_428,N_423);
or U5492 (N_5492,N_93,N_277);
nand U5493 (N_5493,N_1792,N_2311);
nand U5494 (N_5494,N_1209,N_2373);
nand U5495 (N_5495,N_1310,N_1173);
xor U5496 (N_5496,N_323,N_1531);
xor U5497 (N_5497,N_1069,N_2405);
and U5498 (N_5498,N_467,N_2554);
xnor U5499 (N_5499,N_320,N_134);
xnor U5500 (N_5500,N_1851,N_572);
nor U5501 (N_5501,N_1215,N_1757);
nand U5502 (N_5502,N_1510,N_796);
or U5503 (N_5503,N_644,N_1682);
or U5504 (N_5504,N_453,N_132);
and U5505 (N_5505,N_2058,N_2676);
xor U5506 (N_5506,N_1072,N_2924);
nand U5507 (N_5507,N_1156,N_2124);
or U5508 (N_5508,N_1861,N_873);
nand U5509 (N_5509,N_342,N_1032);
and U5510 (N_5510,N_410,N_985);
nand U5511 (N_5511,N_2217,N_1627);
nand U5512 (N_5512,N_814,N_531);
and U5513 (N_5513,N_2296,N_216);
nor U5514 (N_5514,N_1996,N_1409);
xnor U5515 (N_5515,N_2105,N_2249);
and U5516 (N_5516,N_2413,N_817);
xor U5517 (N_5517,N_2548,N_1192);
or U5518 (N_5518,N_19,N_2055);
xnor U5519 (N_5519,N_334,N_1723);
or U5520 (N_5520,N_1184,N_442);
xor U5521 (N_5521,N_313,N_1770);
xor U5522 (N_5522,N_1223,N_1222);
and U5523 (N_5523,N_1822,N_1568);
xnor U5524 (N_5524,N_623,N_1238);
nand U5525 (N_5525,N_434,N_2265);
and U5526 (N_5526,N_245,N_1295);
and U5527 (N_5527,N_2279,N_1883);
nor U5528 (N_5528,N_310,N_364);
and U5529 (N_5529,N_2056,N_1101);
or U5530 (N_5530,N_865,N_2020);
xor U5531 (N_5531,N_2946,N_2161);
or U5532 (N_5532,N_2145,N_88);
xor U5533 (N_5533,N_2724,N_1979);
or U5534 (N_5534,N_1050,N_2852);
and U5535 (N_5535,N_1927,N_380);
or U5536 (N_5536,N_1699,N_1798);
xor U5537 (N_5537,N_1355,N_2276);
xnor U5538 (N_5538,N_694,N_408);
nand U5539 (N_5539,N_17,N_1880);
nor U5540 (N_5540,N_1405,N_253);
nand U5541 (N_5541,N_1959,N_543);
nor U5542 (N_5542,N_1712,N_2470);
nand U5543 (N_5543,N_2022,N_2712);
and U5544 (N_5544,N_408,N_2176);
nor U5545 (N_5545,N_2825,N_2330);
or U5546 (N_5546,N_2078,N_91);
nand U5547 (N_5547,N_1973,N_1919);
nor U5548 (N_5548,N_1734,N_1847);
nand U5549 (N_5549,N_1884,N_2671);
and U5550 (N_5550,N_745,N_1853);
nand U5551 (N_5551,N_1357,N_1369);
and U5552 (N_5552,N_2073,N_2685);
or U5553 (N_5553,N_2747,N_2528);
xor U5554 (N_5554,N_2934,N_474);
xnor U5555 (N_5555,N_1534,N_1559);
xor U5556 (N_5556,N_512,N_1232);
and U5557 (N_5557,N_568,N_2075);
nor U5558 (N_5558,N_634,N_85);
and U5559 (N_5559,N_188,N_902);
xnor U5560 (N_5560,N_1331,N_1503);
nand U5561 (N_5561,N_1776,N_2302);
and U5562 (N_5562,N_717,N_2935);
or U5563 (N_5563,N_1773,N_564);
nor U5564 (N_5564,N_2044,N_1042);
and U5565 (N_5565,N_1004,N_533);
xnor U5566 (N_5566,N_1477,N_2306);
xnor U5567 (N_5567,N_43,N_1023);
and U5568 (N_5568,N_2403,N_2788);
nand U5569 (N_5569,N_2222,N_1415);
or U5570 (N_5570,N_411,N_2794);
and U5571 (N_5571,N_2389,N_969);
and U5572 (N_5572,N_2076,N_2482);
nand U5573 (N_5573,N_715,N_1381);
nor U5574 (N_5574,N_2820,N_2189);
nor U5575 (N_5575,N_866,N_1662);
or U5576 (N_5576,N_1996,N_485);
and U5577 (N_5577,N_207,N_1744);
xor U5578 (N_5578,N_2735,N_2706);
nand U5579 (N_5579,N_1016,N_192);
or U5580 (N_5580,N_2974,N_2943);
and U5581 (N_5581,N_1191,N_2630);
or U5582 (N_5582,N_1642,N_2559);
and U5583 (N_5583,N_1983,N_853);
or U5584 (N_5584,N_610,N_1891);
nand U5585 (N_5585,N_1451,N_983);
and U5586 (N_5586,N_2986,N_2756);
xnor U5587 (N_5587,N_1899,N_2733);
nand U5588 (N_5588,N_2945,N_1768);
and U5589 (N_5589,N_524,N_1457);
nor U5590 (N_5590,N_1988,N_2354);
and U5591 (N_5591,N_2044,N_2521);
or U5592 (N_5592,N_1387,N_235);
nand U5593 (N_5593,N_2780,N_484);
and U5594 (N_5594,N_329,N_490);
or U5595 (N_5595,N_1626,N_1011);
nor U5596 (N_5596,N_940,N_2396);
xor U5597 (N_5597,N_1096,N_122);
and U5598 (N_5598,N_342,N_16);
nor U5599 (N_5599,N_1208,N_1619);
nor U5600 (N_5600,N_2452,N_1447);
and U5601 (N_5601,N_275,N_2633);
and U5602 (N_5602,N_1907,N_2135);
or U5603 (N_5603,N_1566,N_2797);
or U5604 (N_5604,N_2780,N_2465);
or U5605 (N_5605,N_1320,N_2486);
xor U5606 (N_5606,N_720,N_1611);
or U5607 (N_5607,N_11,N_1954);
xor U5608 (N_5608,N_1616,N_252);
nand U5609 (N_5609,N_2784,N_1875);
nand U5610 (N_5610,N_2323,N_1805);
and U5611 (N_5611,N_1520,N_1418);
nor U5612 (N_5612,N_1961,N_222);
nor U5613 (N_5613,N_2491,N_1126);
nor U5614 (N_5614,N_1244,N_310);
xnor U5615 (N_5615,N_1077,N_290);
nor U5616 (N_5616,N_1541,N_997);
nand U5617 (N_5617,N_1956,N_843);
xor U5618 (N_5618,N_5,N_2196);
nor U5619 (N_5619,N_2584,N_842);
nand U5620 (N_5620,N_2147,N_838);
nand U5621 (N_5621,N_2284,N_2387);
xnor U5622 (N_5622,N_1987,N_1221);
or U5623 (N_5623,N_879,N_1387);
nor U5624 (N_5624,N_739,N_1872);
xor U5625 (N_5625,N_1980,N_2298);
or U5626 (N_5626,N_1177,N_2829);
or U5627 (N_5627,N_804,N_901);
and U5628 (N_5628,N_2307,N_2839);
or U5629 (N_5629,N_2771,N_747);
or U5630 (N_5630,N_1257,N_379);
or U5631 (N_5631,N_1176,N_614);
nor U5632 (N_5632,N_2696,N_188);
or U5633 (N_5633,N_1789,N_101);
or U5634 (N_5634,N_1514,N_2713);
and U5635 (N_5635,N_1336,N_2064);
nor U5636 (N_5636,N_2691,N_1661);
xnor U5637 (N_5637,N_2019,N_1831);
and U5638 (N_5638,N_157,N_1537);
nand U5639 (N_5639,N_85,N_577);
or U5640 (N_5640,N_537,N_2084);
nor U5641 (N_5641,N_633,N_2457);
nand U5642 (N_5642,N_1835,N_2680);
nand U5643 (N_5643,N_247,N_930);
and U5644 (N_5644,N_1432,N_633);
or U5645 (N_5645,N_542,N_2671);
and U5646 (N_5646,N_1454,N_1900);
nor U5647 (N_5647,N_2060,N_2339);
and U5648 (N_5648,N_541,N_2165);
nor U5649 (N_5649,N_1254,N_2257);
xor U5650 (N_5650,N_2030,N_129);
and U5651 (N_5651,N_2227,N_1750);
or U5652 (N_5652,N_2897,N_905);
nor U5653 (N_5653,N_390,N_1848);
nor U5654 (N_5654,N_638,N_1111);
nor U5655 (N_5655,N_761,N_1683);
or U5656 (N_5656,N_2666,N_2671);
nor U5657 (N_5657,N_1255,N_150);
nand U5658 (N_5658,N_1614,N_1987);
or U5659 (N_5659,N_264,N_463);
nor U5660 (N_5660,N_657,N_1721);
and U5661 (N_5661,N_857,N_1677);
nor U5662 (N_5662,N_2346,N_95);
or U5663 (N_5663,N_1104,N_711);
or U5664 (N_5664,N_2762,N_241);
nor U5665 (N_5665,N_2855,N_2060);
nand U5666 (N_5666,N_2953,N_881);
nor U5667 (N_5667,N_704,N_599);
or U5668 (N_5668,N_1496,N_971);
nand U5669 (N_5669,N_789,N_450);
xnor U5670 (N_5670,N_1891,N_2237);
or U5671 (N_5671,N_684,N_1002);
and U5672 (N_5672,N_1811,N_1938);
or U5673 (N_5673,N_1058,N_2886);
or U5674 (N_5674,N_563,N_123);
nand U5675 (N_5675,N_1810,N_102);
nand U5676 (N_5676,N_2469,N_1585);
or U5677 (N_5677,N_1480,N_105);
nand U5678 (N_5678,N_667,N_1267);
nand U5679 (N_5679,N_1676,N_1612);
and U5680 (N_5680,N_1448,N_2777);
xor U5681 (N_5681,N_2986,N_2698);
nand U5682 (N_5682,N_244,N_408);
nand U5683 (N_5683,N_1881,N_339);
nand U5684 (N_5684,N_298,N_1919);
or U5685 (N_5685,N_1177,N_1818);
nand U5686 (N_5686,N_2758,N_1573);
xor U5687 (N_5687,N_1663,N_2800);
nand U5688 (N_5688,N_412,N_2488);
nor U5689 (N_5689,N_1875,N_219);
or U5690 (N_5690,N_778,N_1633);
xor U5691 (N_5691,N_1528,N_1710);
or U5692 (N_5692,N_4,N_607);
xnor U5693 (N_5693,N_1532,N_2476);
nor U5694 (N_5694,N_1036,N_2143);
or U5695 (N_5695,N_2217,N_705);
nor U5696 (N_5696,N_254,N_1992);
xor U5697 (N_5697,N_2588,N_622);
and U5698 (N_5698,N_1360,N_1403);
nor U5699 (N_5699,N_1921,N_1456);
xnor U5700 (N_5700,N_2534,N_1118);
or U5701 (N_5701,N_1431,N_359);
or U5702 (N_5702,N_2310,N_2078);
nor U5703 (N_5703,N_1983,N_2563);
nand U5704 (N_5704,N_1012,N_2915);
nor U5705 (N_5705,N_2944,N_1037);
and U5706 (N_5706,N_1487,N_1331);
or U5707 (N_5707,N_2263,N_1428);
nor U5708 (N_5708,N_1565,N_1149);
and U5709 (N_5709,N_1749,N_303);
nor U5710 (N_5710,N_1050,N_1134);
xnor U5711 (N_5711,N_992,N_165);
or U5712 (N_5712,N_640,N_2086);
nand U5713 (N_5713,N_402,N_468);
xor U5714 (N_5714,N_2911,N_2516);
and U5715 (N_5715,N_4,N_412);
nor U5716 (N_5716,N_2160,N_1366);
xnor U5717 (N_5717,N_469,N_696);
xnor U5718 (N_5718,N_1395,N_1203);
xor U5719 (N_5719,N_1776,N_1553);
or U5720 (N_5720,N_1346,N_609);
xor U5721 (N_5721,N_2276,N_1165);
or U5722 (N_5722,N_2464,N_2421);
or U5723 (N_5723,N_1290,N_539);
xnor U5724 (N_5724,N_1773,N_1954);
and U5725 (N_5725,N_2552,N_2052);
nor U5726 (N_5726,N_1194,N_2591);
xor U5727 (N_5727,N_2715,N_1025);
nor U5728 (N_5728,N_1021,N_1778);
or U5729 (N_5729,N_910,N_2389);
nand U5730 (N_5730,N_1582,N_2980);
nand U5731 (N_5731,N_2698,N_761);
nor U5732 (N_5732,N_1152,N_1289);
or U5733 (N_5733,N_2234,N_1829);
nor U5734 (N_5734,N_2014,N_2473);
or U5735 (N_5735,N_584,N_425);
xor U5736 (N_5736,N_2893,N_434);
or U5737 (N_5737,N_388,N_1878);
nor U5738 (N_5738,N_1501,N_2035);
nand U5739 (N_5739,N_1994,N_709);
nor U5740 (N_5740,N_2823,N_834);
xnor U5741 (N_5741,N_1976,N_2723);
nor U5742 (N_5742,N_1472,N_2011);
or U5743 (N_5743,N_1818,N_910);
xnor U5744 (N_5744,N_2493,N_2037);
xor U5745 (N_5745,N_2879,N_574);
or U5746 (N_5746,N_843,N_1606);
and U5747 (N_5747,N_1404,N_993);
and U5748 (N_5748,N_1102,N_86);
and U5749 (N_5749,N_2679,N_1719);
nand U5750 (N_5750,N_1068,N_881);
or U5751 (N_5751,N_1342,N_2634);
and U5752 (N_5752,N_2551,N_2132);
and U5753 (N_5753,N_1356,N_141);
xor U5754 (N_5754,N_1140,N_1641);
or U5755 (N_5755,N_1265,N_1345);
or U5756 (N_5756,N_2811,N_2871);
xnor U5757 (N_5757,N_93,N_1574);
xnor U5758 (N_5758,N_2892,N_1510);
nor U5759 (N_5759,N_2641,N_2675);
nor U5760 (N_5760,N_1050,N_1127);
or U5761 (N_5761,N_305,N_2185);
xnor U5762 (N_5762,N_2981,N_2610);
or U5763 (N_5763,N_499,N_1641);
and U5764 (N_5764,N_2190,N_493);
nor U5765 (N_5765,N_319,N_19);
xor U5766 (N_5766,N_2127,N_2021);
and U5767 (N_5767,N_667,N_2503);
nor U5768 (N_5768,N_2723,N_2851);
or U5769 (N_5769,N_1754,N_2679);
or U5770 (N_5770,N_525,N_1871);
nor U5771 (N_5771,N_1766,N_2468);
nand U5772 (N_5772,N_1608,N_1678);
nor U5773 (N_5773,N_2092,N_2003);
nand U5774 (N_5774,N_1492,N_1791);
and U5775 (N_5775,N_2513,N_1498);
xor U5776 (N_5776,N_1491,N_1285);
xor U5777 (N_5777,N_2155,N_687);
nand U5778 (N_5778,N_159,N_554);
nor U5779 (N_5779,N_2170,N_1629);
xor U5780 (N_5780,N_2151,N_324);
or U5781 (N_5781,N_2516,N_1638);
nand U5782 (N_5782,N_150,N_2510);
nor U5783 (N_5783,N_2542,N_8);
or U5784 (N_5784,N_1955,N_1341);
and U5785 (N_5785,N_1589,N_2305);
nand U5786 (N_5786,N_186,N_1965);
and U5787 (N_5787,N_2752,N_2943);
and U5788 (N_5788,N_2855,N_2944);
or U5789 (N_5789,N_277,N_114);
or U5790 (N_5790,N_156,N_496);
or U5791 (N_5791,N_2030,N_2231);
xnor U5792 (N_5792,N_2552,N_976);
and U5793 (N_5793,N_2816,N_2435);
nor U5794 (N_5794,N_1109,N_2736);
and U5795 (N_5795,N_1921,N_1293);
and U5796 (N_5796,N_2633,N_549);
xnor U5797 (N_5797,N_941,N_857);
nor U5798 (N_5798,N_2383,N_1277);
nand U5799 (N_5799,N_1178,N_805);
or U5800 (N_5800,N_1460,N_1575);
nor U5801 (N_5801,N_2695,N_870);
and U5802 (N_5802,N_714,N_1922);
and U5803 (N_5803,N_2316,N_653);
nand U5804 (N_5804,N_2751,N_1041);
and U5805 (N_5805,N_2784,N_2876);
nor U5806 (N_5806,N_90,N_1957);
nand U5807 (N_5807,N_1074,N_651);
or U5808 (N_5808,N_2685,N_551);
xor U5809 (N_5809,N_2440,N_221);
xnor U5810 (N_5810,N_494,N_2088);
or U5811 (N_5811,N_2124,N_761);
xor U5812 (N_5812,N_313,N_1392);
and U5813 (N_5813,N_248,N_2960);
and U5814 (N_5814,N_2299,N_320);
or U5815 (N_5815,N_1328,N_111);
or U5816 (N_5816,N_72,N_2942);
nor U5817 (N_5817,N_1297,N_2794);
and U5818 (N_5818,N_964,N_2942);
and U5819 (N_5819,N_720,N_505);
xor U5820 (N_5820,N_2841,N_1518);
nand U5821 (N_5821,N_1412,N_2430);
xor U5822 (N_5822,N_1737,N_1196);
or U5823 (N_5823,N_2113,N_1189);
nand U5824 (N_5824,N_1298,N_1685);
and U5825 (N_5825,N_574,N_724);
xor U5826 (N_5826,N_2697,N_1218);
nand U5827 (N_5827,N_901,N_2249);
xnor U5828 (N_5828,N_1941,N_1038);
xor U5829 (N_5829,N_1664,N_2107);
and U5830 (N_5830,N_1867,N_500);
and U5831 (N_5831,N_270,N_690);
nor U5832 (N_5832,N_339,N_2510);
and U5833 (N_5833,N_1937,N_80);
xnor U5834 (N_5834,N_596,N_1467);
or U5835 (N_5835,N_1812,N_1529);
and U5836 (N_5836,N_406,N_732);
xor U5837 (N_5837,N_1076,N_2495);
and U5838 (N_5838,N_2267,N_2338);
and U5839 (N_5839,N_913,N_368);
xor U5840 (N_5840,N_995,N_1237);
or U5841 (N_5841,N_2303,N_1335);
xor U5842 (N_5842,N_2606,N_626);
and U5843 (N_5843,N_2340,N_390);
nand U5844 (N_5844,N_1025,N_2576);
xnor U5845 (N_5845,N_2618,N_424);
or U5846 (N_5846,N_2584,N_2133);
and U5847 (N_5847,N_90,N_1935);
and U5848 (N_5848,N_2664,N_496);
or U5849 (N_5849,N_2510,N_1574);
nor U5850 (N_5850,N_2372,N_875);
nand U5851 (N_5851,N_1957,N_113);
nand U5852 (N_5852,N_1477,N_1983);
or U5853 (N_5853,N_1368,N_2054);
nand U5854 (N_5854,N_1724,N_1644);
nor U5855 (N_5855,N_1728,N_180);
nand U5856 (N_5856,N_835,N_1721);
and U5857 (N_5857,N_1293,N_1974);
and U5858 (N_5858,N_2232,N_1373);
xor U5859 (N_5859,N_1360,N_901);
nand U5860 (N_5860,N_1021,N_391);
and U5861 (N_5861,N_2380,N_2108);
nand U5862 (N_5862,N_1151,N_724);
xnor U5863 (N_5863,N_726,N_1581);
nor U5864 (N_5864,N_2167,N_453);
xor U5865 (N_5865,N_1108,N_1992);
nand U5866 (N_5866,N_637,N_2056);
or U5867 (N_5867,N_1690,N_173);
xor U5868 (N_5868,N_2539,N_2351);
xor U5869 (N_5869,N_1709,N_2064);
and U5870 (N_5870,N_85,N_1620);
and U5871 (N_5871,N_2431,N_1488);
and U5872 (N_5872,N_1071,N_475);
or U5873 (N_5873,N_1278,N_2541);
xnor U5874 (N_5874,N_2847,N_2348);
or U5875 (N_5875,N_74,N_406);
or U5876 (N_5876,N_184,N_2759);
or U5877 (N_5877,N_1208,N_701);
nand U5878 (N_5878,N_1452,N_941);
nor U5879 (N_5879,N_1480,N_7);
nand U5880 (N_5880,N_2531,N_2026);
or U5881 (N_5881,N_877,N_2311);
and U5882 (N_5882,N_776,N_513);
nand U5883 (N_5883,N_1868,N_1434);
nand U5884 (N_5884,N_2615,N_1138);
xnor U5885 (N_5885,N_2234,N_1500);
or U5886 (N_5886,N_43,N_688);
xnor U5887 (N_5887,N_2768,N_2205);
and U5888 (N_5888,N_1611,N_1898);
xnor U5889 (N_5889,N_1597,N_2602);
xor U5890 (N_5890,N_2280,N_2348);
and U5891 (N_5891,N_337,N_810);
and U5892 (N_5892,N_2167,N_699);
nor U5893 (N_5893,N_317,N_2381);
xnor U5894 (N_5894,N_875,N_2778);
and U5895 (N_5895,N_908,N_2194);
nand U5896 (N_5896,N_2109,N_765);
nand U5897 (N_5897,N_940,N_159);
xor U5898 (N_5898,N_2548,N_2643);
nor U5899 (N_5899,N_115,N_424);
nand U5900 (N_5900,N_1717,N_1349);
nand U5901 (N_5901,N_1047,N_67);
and U5902 (N_5902,N_833,N_1281);
xor U5903 (N_5903,N_1969,N_1508);
or U5904 (N_5904,N_362,N_1003);
nor U5905 (N_5905,N_1858,N_1875);
xor U5906 (N_5906,N_2479,N_1950);
nand U5907 (N_5907,N_26,N_2397);
nand U5908 (N_5908,N_2355,N_880);
nand U5909 (N_5909,N_1419,N_1464);
xnor U5910 (N_5910,N_727,N_2116);
nand U5911 (N_5911,N_2540,N_1045);
and U5912 (N_5912,N_20,N_2612);
nand U5913 (N_5913,N_2570,N_2244);
nor U5914 (N_5914,N_2300,N_2552);
or U5915 (N_5915,N_2629,N_1814);
nor U5916 (N_5916,N_482,N_1725);
and U5917 (N_5917,N_1803,N_1084);
or U5918 (N_5918,N_2540,N_2910);
and U5919 (N_5919,N_427,N_885);
xor U5920 (N_5920,N_1105,N_211);
nand U5921 (N_5921,N_1003,N_813);
or U5922 (N_5922,N_1874,N_34);
or U5923 (N_5923,N_2546,N_2878);
xnor U5924 (N_5924,N_463,N_1200);
xor U5925 (N_5925,N_1273,N_2534);
xor U5926 (N_5926,N_1933,N_1769);
nor U5927 (N_5927,N_1087,N_2787);
xor U5928 (N_5928,N_1711,N_873);
nand U5929 (N_5929,N_1715,N_99);
nand U5930 (N_5930,N_1411,N_2694);
nor U5931 (N_5931,N_1532,N_1446);
and U5932 (N_5932,N_2007,N_1807);
or U5933 (N_5933,N_2945,N_745);
nor U5934 (N_5934,N_1716,N_923);
nor U5935 (N_5935,N_1763,N_139);
xnor U5936 (N_5936,N_2323,N_2289);
xor U5937 (N_5937,N_1116,N_2373);
xnor U5938 (N_5938,N_1064,N_2757);
nand U5939 (N_5939,N_1268,N_2354);
xnor U5940 (N_5940,N_1463,N_2255);
nand U5941 (N_5941,N_99,N_663);
nand U5942 (N_5942,N_19,N_1341);
nand U5943 (N_5943,N_1656,N_36);
nand U5944 (N_5944,N_230,N_1844);
and U5945 (N_5945,N_847,N_2862);
or U5946 (N_5946,N_2140,N_1282);
or U5947 (N_5947,N_1264,N_2462);
and U5948 (N_5948,N_28,N_399);
nor U5949 (N_5949,N_2947,N_984);
and U5950 (N_5950,N_1003,N_195);
xor U5951 (N_5951,N_83,N_1804);
and U5952 (N_5952,N_358,N_380);
nand U5953 (N_5953,N_472,N_1815);
or U5954 (N_5954,N_1264,N_1327);
xnor U5955 (N_5955,N_60,N_1804);
and U5956 (N_5956,N_2051,N_334);
or U5957 (N_5957,N_1045,N_329);
or U5958 (N_5958,N_2710,N_1149);
nor U5959 (N_5959,N_2912,N_1013);
xor U5960 (N_5960,N_2603,N_1323);
xor U5961 (N_5961,N_2270,N_2401);
and U5962 (N_5962,N_246,N_1275);
xnor U5963 (N_5963,N_2251,N_2829);
or U5964 (N_5964,N_306,N_28);
or U5965 (N_5965,N_1584,N_2943);
nor U5966 (N_5966,N_1835,N_92);
nor U5967 (N_5967,N_2168,N_275);
or U5968 (N_5968,N_1500,N_1213);
xnor U5969 (N_5969,N_2123,N_1671);
xnor U5970 (N_5970,N_2861,N_467);
or U5971 (N_5971,N_2563,N_51);
and U5972 (N_5972,N_725,N_2559);
or U5973 (N_5973,N_293,N_2722);
and U5974 (N_5974,N_1391,N_2541);
or U5975 (N_5975,N_1147,N_339);
xnor U5976 (N_5976,N_8,N_1973);
nand U5977 (N_5977,N_2302,N_477);
nand U5978 (N_5978,N_2692,N_2861);
and U5979 (N_5979,N_1713,N_1844);
nor U5980 (N_5980,N_1478,N_570);
nor U5981 (N_5981,N_2603,N_2758);
and U5982 (N_5982,N_1449,N_2867);
xor U5983 (N_5983,N_1374,N_1986);
and U5984 (N_5984,N_2317,N_2823);
nand U5985 (N_5985,N_177,N_2312);
nor U5986 (N_5986,N_938,N_1018);
nand U5987 (N_5987,N_509,N_2401);
nor U5988 (N_5988,N_2617,N_1051);
nor U5989 (N_5989,N_881,N_2381);
nor U5990 (N_5990,N_215,N_222);
nor U5991 (N_5991,N_1044,N_417);
nand U5992 (N_5992,N_1291,N_1781);
nor U5993 (N_5993,N_495,N_221);
nor U5994 (N_5994,N_1291,N_1300);
or U5995 (N_5995,N_361,N_2846);
nand U5996 (N_5996,N_2052,N_1308);
nor U5997 (N_5997,N_1112,N_1068);
xnor U5998 (N_5998,N_2845,N_1077);
and U5999 (N_5999,N_2730,N_2802);
and U6000 (N_6000,N_4160,N_3151);
and U6001 (N_6001,N_4199,N_4746);
xnor U6002 (N_6002,N_5316,N_3342);
or U6003 (N_6003,N_3457,N_4586);
xor U6004 (N_6004,N_4078,N_3716);
and U6005 (N_6005,N_5386,N_4304);
nor U6006 (N_6006,N_5222,N_5132);
and U6007 (N_6007,N_3557,N_5375);
or U6008 (N_6008,N_3464,N_3926);
nor U6009 (N_6009,N_3864,N_4056);
and U6010 (N_6010,N_3204,N_5557);
nand U6011 (N_6011,N_5506,N_5959);
nor U6012 (N_6012,N_5075,N_5427);
and U6013 (N_6013,N_4456,N_4856);
nor U6014 (N_6014,N_4901,N_4531);
nand U6015 (N_6015,N_5465,N_4335);
nand U6016 (N_6016,N_4127,N_5763);
nor U6017 (N_6017,N_3205,N_5786);
or U6018 (N_6018,N_3799,N_3721);
xor U6019 (N_6019,N_4870,N_4450);
xnor U6020 (N_6020,N_5511,N_4756);
or U6021 (N_6021,N_5153,N_4336);
or U6022 (N_6022,N_5587,N_4767);
and U6023 (N_6023,N_5559,N_5814);
and U6024 (N_6024,N_4973,N_3529);
nand U6025 (N_6025,N_5522,N_4863);
and U6026 (N_6026,N_3411,N_5521);
nand U6027 (N_6027,N_3167,N_4267);
xnor U6028 (N_6028,N_4244,N_5501);
or U6029 (N_6029,N_4597,N_3299);
and U6030 (N_6030,N_4491,N_3059);
xnor U6031 (N_6031,N_5196,N_3880);
or U6032 (N_6032,N_4059,N_4754);
nand U6033 (N_6033,N_3622,N_3448);
and U6034 (N_6034,N_3596,N_5246);
or U6035 (N_6035,N_5027,N_3476);
and U6036 (N_6036,N_3128,N_5237);
xnor U6037 (N_6037,N_3691,N_5136);
and U6038 (N_6038,N_4383,N_4393);
nand U6039 (N_6039,N_5586,N_4238);
and U6040 (N_6040,N_5727,N_4681);
or U6041 (N_6041,N_5601,N_4382);
nor U6042 (N_6042,N_3994,N_4793);
and U6043 (N_6043,N_3311,N_3748);
xor U6044 (N_6044,N_3582,N_5849);
nor U6045 (N_6045,N_4709,N_3187);
or U6046 (N_6046,N_4636,N_3254);
nand U6047 (N_6047,N_5733,N_5093);
xor U6048 (N_6048,N_5900,N_5764);
nand U6049 (N_6049,N_4418,N_5867);
and U6050 (N_6050,N_4295,N_3564);
nor U6051 (N_6051,N_5998,N_3365);
or U6052 (N_6052,N_5991,N_4224);
xnor U6053 (N_6053,N_4432,N_3279);
nor U6054 (N_6054,N_5212,N_5072);
xor U6055 (N_6055,N_3608,N_3953);
nand U6056 (N_6056,N_5512,N_3911);
and U6057 (N_6057,N_4074,N_3803);
or U6058 (N_6058,N_3303,N_3966);
nand U6059 (N_6059,N_3870,N_4262);
or U6060 (N_6060,N_3895,N_4265);
nand U6061 (N_6061,N_3730,N_4807);
or U6062 (N_6062,N_3935,N_5154);
nor U6063 (N_6063,N_4520,N_4953);
or U6064 (N_6064,N_5113,N_3406);
and U6065 (N_6065,N_5757,N_5810);
or U6066 (N_6066,N_4891,N_5207);
nor U6067 (N_6067,N_5467,N_3087);
and U6068 (N_6068,N_4518,N_3758);
or U6069 (N_6069,N_3404,N_5343);
or U6070 (N_6070,N_3467,N_4678);
or U6071 (N_6071,N_5564,N_5739);
xor U6072 (N_6072,N_3751,N_5595);
or U6073 (N_6073,N_4225,N_3216);
nor U6074 (N_6074,N_4300,N_4899);
and U6075 (N_6075,N_4037,N_5852);
nor U6076 (N_6076,N_5104,N_5088);
nor U6077 (N_6077,N_4747,N_5340);
and U6078 (N_6078,N_3675,N_5156);
and U6079 (N_6079,N_5933,N_4970);
or U6080 (N_6080,N_5517,N_3732);
xnor U6081 (N_6081,N_3802,N_3416);
and U6082 (N_6082,N_4112,N_4796);
or U6083 (N_6083,N_5844,N_3274);
or U6084 (N_6084,N_3649,N_3912);
nor U6085 (N_6085,N_3019,N_4342);
xor U6086 (N_6086,N_5803,N_4632);
xor U6087 (N_6087,N_5653,N_3625);
or U6088 (N_6088,N_5001,N_4400);
and U6089 (N_6089,N_3360,N_5502);
and U6090 (N_6090,N_4490,N_4315);
nor U6091 (N_6091,N_3916,N_5215);
and U6092 (N_6092,N_4191,N_3369);
nor U6093 (N_6093,N_4405,N_5235);
and U6094 (N_6094,N_4853,N_4227);
or U6095 (N_6095,N_3735,N_3357);
nor U6096 (N_6096,N_3887,N_4539);
xnor U6097 (N_6097,N_3615,N_5974);
xnor U6098 (N_6098,N_4297,N_4394);
and U6099 (N_6099,N_3617,N_5192);
or U6100 (N_6100,N_5719,N_5090);
nor U6101 (N_6101,N_3709,N_4766);
xnor U6102 (N_6102,N_3325,N_4298);
nand U6103 (N_6103,N_3093,N_3149);
nor U6104 (N_6104,N_4617,N_4880);
nor U6105 (N_6105,N_5330,N_4446);
xnor U6106 (N_6106,N_3872,N_5297);
xnor U6107 (N_6107,N_3648,N_4163);
or U6108 (N_6108,N_3845,N_5703);
or U6109 (N_6109,N_5445,N_3373);
xor U6110 (N_6110,N_4554,N_5817);
nand U6111 (N_6111,N_3057,N_5244);
or U6112 (N_6112,N_3367,N_4139);
nor U6113 (N_6113,N_3929,N_5050);
and U6114 (N_6114,N_3745,N_4634);
or U6115 (N_6115,N_3560,N_4320);
and U6116 (N_6116,N_5681,N_4473);
nor U6117 (N_6117,N_5581,N_4562);
nor U6118 (N_6118,N_3694,N_3144);
and U6119 (N_6119,N_3066,N_4967);
or U6120 (N_6120,N_5223,N_4311);
nor U6121 (N_6121,N_5385,N_4811);
and U6122 (N_6122,N_4706,N_5528);
and U6123 (N_6123,N_5495,N_4555);
xnor U6124 (N_6124,N_3381,N_4118);
or U6125 (N_6125,N_5774,N_5463);
nand U6126 (N_6126,N_4607,N_3987);
xor U6127 (N_6127,N_5646,N_5723);
or U6128 (N_6128,N_3460,N_5578);
nand U6129 (N_6129,N_4072,N_5789);
and U6130 (N_6130,N_5802,N_4826);
and U6131 (N_6131,N_5197,N_5060);
xnor U6132 (N_6132,N_4553,N_3168);
nand U6133 (N_6133,N_3993,N_3920);
nand U6134 (N_6134,N_5069,N_3978);
and U6135 (N_6135,N_3762,N_3343);
and U6136 (N_6136,N_3296,N_4363);
nand U6137 (N_6137,N_4358,N_4557);
and U6138 (N_6138,N_3702,N_4344);
nor U6139 (N_6139,N_5538,N_4660);
or U6140 (N_6140,N_3830,N_5740);
xnor U6141 (N_6141,N_4639,N_4855);
xor U6142 (N_6142,N_5450,N_3714);
nand U6143 (N_6143,N_4338,N_3263);
nor U6144 (N_6144,N_3364,N_3842);
nor U6145 (N_6145,N_5234,N_5128);
nand U6146 (N_6146,N_3973,N_3494);
xor U6147 (N_6147,N_3697,N_3105);
xor U6148 (N_6148,N_5308,N_3772);
xnor U6149 (N_6149,N_4701,N_5031);
and U6150 (N_6150,N_3933,N_5454);
nor U6151 (N_6151,N_5364,N_5049);
nor U6152 (N_6152,N_3629,N_3248);
xor U6153 (N_6153,N_3162,N_3421);
xor U6154 (N_6154,N_3152,N_3073);
nor U6155 (N_6155,N_3155,N_4390);
and U6156 (N_6156,N_3452,N_4695);
or U6157 (N_6157,N_4522,N_5989);
or U6158 (N_6158,N_4100,N_3956);
and U6159 (N_6159,N_3388,N_3007);
and U6160 (N_6160,N_5905,N_4534);
nor U6161 (N_6161,N_4837,N_4563);
nand U6162 (N_6162,N_3042,N_4328);
or U6163 (N_6163,N_3150,N_3812);
or U6164 (N_6164,N_5206,N_5519);
xnor U6165 (N_6165,N_5143,N_5417);
and U6166 (N_6166,N_5063,N_5391);
nand U6167 (N_6167,N_5129,N_4472);
or U6168 (N_6168,N_3233,N_4571);
nor U6169 (N_6169,N_4388,N_3511);
nor U6170 (N_6170,N_4879,N_5580);
nand U6171 (N_6171,N_3711,N_5608);
or U6172 (N_6172,N_3638,N_5634);
and U6173 (N_6173,N_4349,N_5510);
or U6174 (N_6174,N_3489,N_4261);
nor U6175 (N_6175,N_3260,N_3881);
and U6176 (N_6176,N_4201,N_5529);
nor U6177 (N_6177,N_4384,N_3137);
xnor U6178 (N_6178,N_3027,N_5710);
xor U6179 (N_6179,N_5273,N_5876);
nor U6180 (N_6180,N_4887,N_5397);
nor U6181 (N_6181,N_3715,N_4969);
or U6182 (N_6182,N_3478,N_3195);
nor U6183 (N_6183,N_5535,N_4339);
or U6184 (N_6184,N_4233,N_3555);
nand U6185 (N_6185,N_5198,N_4192);
or U6186 (N_6186,N_3796,N_4448);
or U6187 (N_6187,N_4618,N_4054);
or U6188 (N_6188,N_4540,N_4172);
nand U6189 (N_6189,N_4944,N_5277);
nand U6190 (N_6190,N_4535,N_3766);
xor U6191 (N_6191,N_4376,N_3996);
and U6192 (N_6192,N_4980,N_4457);
or U6193 (N_6193,N_3614,N_5741);
nand U6194 (N_6194,N_4791,N_4246);
nor U6195 (N_6195,N_4612,N_4854);
or U6196 (N_6196,N_3484,N_5422);
and U6197 (N_6197,N_5641,N_3346);
nor U6198 (N_6198,N_5819,N_4551);
nor U6199 (N_6199,N_4442,N_5468);
xor U6200 (N_6200,N_4275,N_5761);
nand U6201 (N_6201,N_4988,N_5614);
and U6202 (N_6202,N_4596,N_3662);
or U6203 (N_6203,N_3485,N_4759);
nor U6204 (N_6204,N_3683,N_4651);
or U6205 (N_6205,N_4164,N_5765);
and U6206 (N_6206,N_4094,N_3112);
and U6207 (N_6207,N_5058,N_3655);
nor U6208 (N_6208,N_3679,N_5592);
or U6209 (N_6209,N_3992,N_3652);
nand U6210 (N_6210,N_4242,N_3193);
and U6211 (N_6211,N_4915,N_3671);
nor U6212 (N_6212,N_5806,N_4377);
or U6213 (N_6213,N_4287,N_5863);
or U6214 (N_6214,N_3164,N_3071);
nand U6215 (N_6215,N_5253,N_3665);
or U6216 (N_6216,N_5338,N_3838);
nand U6217 (N_6217,N_4273,N_3674);
nand U6218 (N_6218,N_3503,N_4114);
and U6219 (N_6219,N_5563,N_5505);
and U6220 (N_6220,N_4486,N_4061);
nand U6221 (N_6221,N_5091,N_3836);
and U6222 (N_6222,N_3451,N_3814);
xnor U6223 (N_6223,N_4169,N_3449);
nor U6224 (N_6224,N_3053,N_3639);
nand U6225 (N_6225,N_5409,N_5301);
or U6226 (N_6226,N_5248,N_3826);
nor U6227 (N_6227,N_4380,N_4185);
nand U6228 (N_6228,N_5408,N_4797);
or U6229 (N_6229,N_3191,N_5399);
nor U6230 (N_6230,N_4578,N_3862);
or U6231 (N_6231,N_3368,N_5770);
nand U6232 (N_6232,N_4728,N_3713);
or U6233 (N_6233,N_5562,N_3521);
xnor U6234 (N_6234,N_5350,N_5100);
xor U6235 (N_6235,N_4071,N_4814);
or U6236 (N_6236,N_4802,N_3526);
xnor U6237 (N_6237,N_3454,N_3182);
nor U6238 (N_6238,N_5910,N_5187);
or U6239 (N_6239,N_5281,N_5547);
or U6240 (N_6240,N_4017,N_5607);
nand U6241 (N_6241,N_3820,N_5329);
nand U6242 (N_6242,N_3969,N_3473);
xnor U6243 (N_6243,N_4036,N_4753);
nand U6244 (N_6244,N_4402,N_4296);
and U6245 (N_6245,N_4408,N_4111);
nor U6246 (N_6246,N_4708,N_3499);
nor U6247 (N_6247,N_5327,N_4626);
xor U6248 (N_6248,N_4058,N_5381);
and U6249 (N_6249,N_4454,N_5239);
xnor U6250 (N_6250,N_3946,N_4808);
xor U6251 (N_6251,N_3528,N_3703);
or U6252 (N_6252,N_5430,N_4326);
nor U6253 (N_6253,N_3861,N_5455);
xor U6254 (N_6254,N_3746,N_4070);
or U6255 (N_6255,N_4699,N_5029);
nand U6256 (N_6256,N_3349,N_5367);
xnor U6257 (N_6257,N_3479,N_5322);
or U6258 (N_6258,N_3657,N_5688);
nand U6259 (N_6259,N_4720,N_5026);
nor U6260 (N_6260,N_5161,N_3125);
and U6261 (N_6261,N_3624,N_3623);
or U6262 (N_6262,N_3919,N_4369);
nand U6263 (N_6263,N_3284,N_5992);
or U6264 (N_6264,N_5282,N_4929);
nand U6265 (N_6265,N_4444,N_3446);
nand U6266 (N_6266,N_3375,N_5285);
nand U6267 (N_6267,N_3597,N_5159);
nor U6268 (N_6268,N_4467,N_5635);
nand U6269 (N_6269,N_3447,N_3100);
xnor U6270 (N_6270,N_5176,N_5070);
or U6271 (N_6271,N_5489,N_3773);
or U6272 (N_6272,N_3395,N_5649);
nand U6273 (N_6273,N_3921,N_4313);
nand U6274 (N_6274,N_4680,N_3654);
and U6275 (N_6275,N_5326,N_3653);
and U6276 (N_6276,N_5400,N_5828);
nand U6277 (N_6277,N_4782,N_3593);
nand U6278 (N_6278,N_4080,N_4875);
and U6279 (N_6279,N_5032,N_4182);
and U6280 (N_6280,N_4375,N_5659);
and U6281 (N_6281,N_3753,N_5021);
or U6282 (N_6282,N_4868,N_4820);
or U6283 (N_6283,N_3111,N_5780);
and U6284 (N_6284,N_3483,N_4842);
and U6285 (N_6285,N_5531,N_4477);
xor U6286 (N_6286,N_5642,N_3083);
and U6287 (N_6287,N_4079,N_5271);
and U6288 (N_6288,N_5080,N_5724);
or U6289 (N_6289,N_4744,N_5262);
nor U6290 (N_6290,N_4209,N_3287);
nand U6291 (N_6291,N_5302,N_3143);
xnor U6292 (N_6292,N_3698,N_4284);
or U6293 (N_6293,N_4015,N_5439);
and U6294 (N_6294,N_3749,N_4513);
nor U6295 (N_6295,N_5389,N_5371);
and U6296 (N_6296,N_3902,N_5351);
nand U6297 (N_6297,N_5336,N_5986);
xor U6298 (N_6298,N_4737,N_4956);
nand U6299 (N_6299,N_5163,N_4960);
xor U6300 (N_6300,N_3062,N_5792);
nor U6301 (N_6301,N_4498,N_5576);
and U6302 (N_6302,N_5861,N_4568);
and U6303 (N_6303,N_5854,N_3551);
xor U6304 (N_6304,N_3372,N_3334);
xnor U6305 (N_6305,N_4628,N_3682);
xor U6306 (N_6306,N_3958,N_3659);
nor U6307 (N_6307,N_5458,N_4593);
and U6308 (N_6308,N_3177,N_4009);
or U6309 (N_6309,N_5660,N_5219);
or U6310 (N_6310,N_3009,N_5323);
and U6311 (N_6311,N_4642,N_5288);
xnor U6312 (N_6312,N_4417,N_4232);
or U6313 (N_6313,N_3206,N_4455);
or U6314 (N_6314,N_5625,N_5085);
nand U6315 (N_6315,N_5808,N_3043);
nor U6316 (N_6316,N_4406,N_3514);
and U6317 (N_6317,N_5254,N_5315);
and U6318 (N_6318,N_4102,N_5707);
xor U6319 (N_6319,N_5084,N_5729);
xor U6320 (N_6320,N_3272,N_3428);
nand U6321 (N_6321,N_3562,N_3539);
or U6322 (N_6322,N_4926,N_4995);
or U6323 (N_6323,N_5436,N_5945);
xor U6324 (N_6324,N_5024,N_3542);
nor U6325 (N_6325,N_5928,N_3658);
nand U6326 (N_6326,N_4239,N_5872);
or U6327 (N_6327,N_4395,N_5339);
or U6328 (N_6328,N_5516,N_4906);
nor U6329 (N_6329,N_5611,N_4914);
xor U6330 (N_6330,N_5444,N_4140);
nand U6331 (N_6331,N_3957,N_5842);
xnor U6332 (N_6332,N_5476,N_4487);
xnor U6333 (N_6333,N_3418,N_3630);
xor U6334 (N_6334,N_4823,N_3985);
xnor U6335 (N_6335,N_4819,N_3856);
nand U6336 (N_6336,N_5978,N_3977);
and U6337 (N_6337,N_3554,N_5145);
and U6338 (N_6338,N_3581,N_4286);
xor U6339 (N_6339,N_5286,N_3298);
xor U6340 (N_6340,N_3245,N_3183);
or U6341 (N_6341,N_3393,N_5210);
xnor U6342 (N_6342,N_5648,N_5457);
xor U6343 (N_6343,N_4096,N_5833);
xnor U6344 (N_6344,N_3747,N_5704);
nand U6345 (N_6345,N_5260,N_5200);
and U6346 (N_6346,N_5541,N_5499);
or U6347 (N_6347,N_4881,N_3626);
nand U6348 (N_6348,N_4235,N_4266);
or U6349 (N_6349,N_4218,N_4052);
nor U6350 (N_6350,N_3770,N_5868);
nand U6351 (N_6351,N_3278,N_5862);
and U6352 (N_6352,N_3378,N_3914);
and U6353 (N_6353,N_5579,N_4175);
or U6354 (N_6354,N_3505,N_4895);
nand U6355 (N_6355,N_3074,N_5894);
and U6356 (N_6356,N_5107,N_3081);
xor U6357 (N_6357,N_3795,N_3632);
or U6358 (N_6358,N_3832,N_3220);
nand U6359 (N_6359,N_5298,N_4399);
xor U6360 (N_6360,N_5878,N_3215);
xor U6361 (N_6361,N_3048,N_4035);
xor U6362 (N_6362,N_5694,N_3883);
nand U6363 (N_6363,N_5346,N_5355);
nor U6364 (N_6364,N_4585,N_5834);
nor U6365 (N_6365,N_4134,N_3901);
or U6366 (N_6366,N_5484,N_4171);
xor U6367 (N_6367,N_5575,N_4143);
and U6368 (N_6368,N_4806,N_5380);
xnor U6369 (N_6369,N_5744,N_5337);
xor U6370 (N_6370,N_4545,N_3121);
or U6371 (N_6371,N_4829,N_5447);
nand U6372 (N_6372,N_3056,N_3376);
or U6373 (N_6373,N_3174,N_4162);
nand U6374 (N_6374,N_5602,N_4379);
or U6375 (N_6375,N_5996,N_3099);
nor U6376 (N_6376,N_4846,N_5256);
and U6377 (N_6377,N_3277,N_5065);
xnor U6378 (N_6378,N_3094,N_3179);
nand U6379 (N_6379,N_3319,N_4838);
nand U6380 (N_6380,N_4504,N_5202);
nand U6381 (N_6381,N_4962,N_4088);
or U6382 (N_6382,N_3540,N_3959);
nor U6383 (N_6383,N_4635,N_3570);
and U6384 (N_6384,N_3619,N_3385);
xnor U6385 (N_6385,N_5885,N_5583);
or U6386 (N_6386,N_3684,N_3595);
nor U6387 (N_6387,N_5094,N_3673);
nand U6388 (N_6388,N_5356,N_4871);
and U6389 (N_6389,N_3333,N_5721);
and U6390 (N_6390,N_4420,N_4445);
or U6391 (N_6391,N_5162,N_4482);
nand U6392 (N_6392,N_3685,N_5233);
nand U6393 (N_6393,N_5948,N_4057);
nor U6394 (N_6394,N_4577,N_4149);
and U6395 (N_6395,N_3923,N_4279);
and U6396 (N_6396,N_3231,N_5022);
nor U6397 (N_6397,N_5300,N_5801);
and U6398 (N_6398,N_5403,N_5728);
nor U6399 (N_6399,N_3792,N_3900);
nor U6400 (N_6400,N_4961,N_5204);
nand U6401 (N_6401,N_5018,N_3873);
xor U6402 (N_6402,N_5464,N_3317);
and U6403 (N_6403,N_5686,N_5108);
xor U6404 (N_6404,N_4260,N_4775);
nand U6405 (N_6405,N_5482,N_5068);
and U6406 (N_6406,N_3510,N_4290);
nand U6407 (N_6407,N_3816,N_5172);
nand U6408 (N_6408,N_5800,N_4018);
and U6409 (N_6409,N_3192,N_5735);
nand U6410 (N_6410,N_5263,N_5048);
or U6411 (N_6411,N_4452,N_5631);
nand U6412 (N_6412,N_4422,N_3670);
and U6413 (N_6413,N_5972,N_5904);
or U6414 (N_6414,N_3991,N_5217);
or U6415 (N_6415,N_5241,N_4007);
nor U6416 (N_6416,N_5416,N_3313);
and U6417 (N_6417,N_5916,N_3998);
xnor U6418 (N_6418,N_4318,N_5428);
nand U6419 (N_6419,N_4173,N_5616);
and U6420 (N_6420,N_4966,N_4629);
nor U6421 (N_6421,N_4546,N_5979);
xor U6422 (N_6422,N_4785,N_3061);
nand U6423 (N_6423,N_5860,N_5177);
or U6424 (N_6424,N_4957,N_5255);
and U6425 (N_6425,N_3603,N_4888);
and U6426 (N_6426,N_4653,N_4489);
xnor U6427 (N_6427,N_4606,N_4833);
xor U6428 (N_6428,N_4253,N_3525);
xor U6429 (N_6429,N_3261,N_5398);
nand U6430 (N_6430,N_4240,N_4768);
nand U6431 (N_6431,N_3780,N_3898);
and U6432 (N_6432,N_4702,N_5451);
xnor U6433 (N_6433,N_5965,N_3127);
and U6434 (N_6434,N_5194,N_4582);
or U6435 (N_6435,N_3607,N_5170);
or U6436 (N_6436,N_4067,N_3480);
xor U6437 (N_6437,N_5433,N_5208);
or U6438 (N_6438,N_5086,N_3701);
nand U6439 (N_6439,N_3450,N_4116);
nor U6440 (N_6440,N_5691,N_4503);
or U6441 (N_6441,N_4048,N_4060);
or U6442 (N_6442,N_5171,N_4986);
nand U6443 (N_6443,N_4101,N_4893);
and U6444 (N_6444,N_5937,N_3806);
xor U6445 (N_6445,N_5497,N_5361);
and U6446 (N_6446,N_5665,N_4740);
nand U6447 (N_6447,N_3255,N_3332);
and U6448 (N_6448,N_3793,N_3229);
nand U6449 (N_6449,N_3080,N_3944);
nor U6450 (N_6450,N_4921,N_3647);
and U6451 (N_6451,N_4896,N_3930);
or U6452 (N_6452,N_3790,N_5790);
and U6453 (N_6453,N_3269,N_5750);
and U6454 (N_6454,N_5618,N_4451);
or U6455 (N_6455,N_5787,N_3435);
xor U6456 (N_6456,N_4144,N_4705);
or U6457 (N_6457,N_5289,N_4027);
nand U6458 (N_6458,N_4510,N_5742);
nor U6459 (N_6459,N_3178,N_5782);
xnor U6460 (N_6460,N_4347,N_4784);
and U6461 (N_6461,N_5307,N_5836);
and U6462 (N_6462,N_4126,N_4427);
xnor U6463 (N_6463,N_3469,N_3787);
nor U6464 (N_6464,N_4924,N_4549);
xnor U6465 (N_6465,N_3184,N_5655);
and U6466 (N_6466,N_5150,N_4188);
or U6467 (N_6467,N_4974,N_4258);
nor U6468 (N_6468,N_5778,N_4935);
xnor U6469 (N_6469,N_5321,N_5847);
or U6470 (N_6470,N_5483,N_3288);
nor U6471 (N_6471,N_4952,N_4329);
nand U6472 (N_6472,N_5829,N_3153);
nor U6473 (N_6473,N_5121,N_3018);
and U6474 (N_6474,N_4624,N_3202);
nand U6475 (N_6475,N_3586,N_3217);
nor U6476 (N_6476,N_3165,N_4998);
xnor U6477 (N_6477,N_3390,N_5822);
and U6478 (N_6478,N_3548,N_3733);
nand U6479 (N_6479,N_3804,N_3013);
xnor U6480 (N_6480,N_4834,N_3142);
or U6481 (N_6481,N_3271,N_4282);
or U6482 (N_6482,N_3337,N_4142);
nor U6483 (N_6483,N_3444,N_5925);
or U6484 (N_6484,N_5053,N_4174);
or U6485 (N_6485,N_5759,N_4200);
or U6486 (N_6486,N_4497,N_3869);
and U6487 (N_6487,N_3492,N_4438);
nand U6488 (N_6488,N_3208,N_5067);
nand U6489 (N_6489,N_3847,N_5283);
and U6490 (N_6490,N_3620,N_3351);
nand U6491 (N_6491,N_5677,N_4464);
nor U6492 (N_6492,N_4291,N_5961);
or U6493 (N_6493,N_5624,N_3440);
or U6494 (N_6494,N_3641,N_5264);
nand U6495 (N_6495,N_5354,N_3481);
or U6496 (N_6496,N_3610,N_4180);
nand U6497 (N_6497,N_5919,N_4928);
xnor U6498 (N_6498,N_5966,N_5908);
xor U6499 (N_6499,N_4958,N_5769);
nor U6500 (N_6500,N_3135,N_5319);
and U6501 (N_6501,N_5629,N_4356);
nor U6502 (N_6502,N_5440,N_5692);
and U6503 (N_6503,N_4830,N_4836);
xnor U6504 (N_6504,N_3282,N_4857);
xnor U6505 (N_6505,N_4665,N_5672);
and U6506 (N_6506,N_4023,N_3108);
xnor U6507 (N_6507,N_3857,N_3173);
and U6508 (N_6508,N_5475,N_3544);
or U6509 (N_6509,N_4511,N_4062);
and U6510 (N_6510,N_3871,N_5663);
and U6511 (N_6511,N_5130,N_5472);
xor U6512 (N_6512,N_5619,N_4099);
nor U6513 (N_6513,N_5395,N_5983);
nor U6514 (N_6514,N_3576,N_3771);
and U6515 (N_6515,N_3491,N_5668);
xnor U6516 (N_6516,N_4302,N_3633);
nor U6517 (N_6517,N_5066,N_5656);
xor U6518 (N_6518,N_5938,N_3955);
nor U6519 (N_6519,N_3309,N_3338);
nand U6520 (N_6520,N_5525,N_5932);
nor U6521 (N_6521,N_4724,N_4495);
and U6522 (N_6522,N_3997,N_4777);
nor U6523 (N_6523,N_3681,N_3818);
nand U6524 (N_6524,N_3030,N_5929);
or U6525 (N_6525,N_4908,N_4779);
nor U6526 (N_6526,N_4755,N_3903);
nor U6527 (N_6527,N_3218,N_3513);
or U6528 (N_6528,N_3865,N_3600);
nor U6529 (N_6529,N_3038,N_3199);
nor U6530 (N_6530,N_3877,N_5820);
nor U6531 (N_6531,N_3237,N_4983);
and U6532 (N_6532,N_3238,N_4002);
xor U6533 (N_6533,N_4044,N_5266);
nor U6534 (N_6534,N_5775,N_5591);
and U6535 (N_6535,N_5312,N_4712);
nand U6536 (N_6536,N_5008,N_4308);
nand U6537 (N_6537,N_4198,N_3858);
nand U6538 (N_6538,N_4301,N_5508);
nor U6539 (N_6539,N_4193,N_3190);
and U6540 (N_6540,N_4008,N_4972);
or U6541 (N_6541,N_3983,N_5807);
nor U6542 (N_6542,N_5035,N_3241);
or U6543 (N_6543,N_5047,N_5737);
or U6544 (N_6544,N_4374,N_5209);
or U6545 (N_6545,N_5421,N_5382);
or U6546 (N_6546,N_5556,N_3239);
and U6547 (N_6547,N_3899,N_4508);
and U6548 (N_6548,N_4250,N_5824);
xor U6549 (N_6549,N_3196,N_4798);
nor U6550 (N_6550,N_3527,N_3981);
or U6551 (N_6551,N_5539,N_4194);
and U6552 (N_6552,N_3386,N_3226);
nor U6553 (N_6553,N_4421,N_4346);
and U6554 (N_6554,N_4788,N_5042);
nor U6555 (N_6555,N_3886,N_5141);
xnor U6556 (N_6556,N_3234,N_5762);
or U6557 (N_6557,N_4909,N_4687);
nand U6558 (N_6558,N_3875,N_4673);
nand U6559 (N_6559,N_4396,N_4466);
or U6560 (N_6560,N_5857,N_3291);
nand U6561 (N_6561,N_4413,N_3072);
nand U6562 (N_6562,N_3396,N_3706);
or U6563 (N_6563,N_3295,N_5142);
nand U6564 (N_6564,N_5924,N_3024);
xor U6565 (N_6565,N_4789,N_3391);
xor U6566 (N_6566,N_4475,N_4576);
nor U6567 (N_6567,N_4312,N_4321);
or U6568 (N_6568,N_5685,N_5605);
nor U6569 (N_6569,N_5344,N_3146);
or U6570 (N_6570,N_4424,N_3722);
nor U6571 (N_6571,N_3124,N_4595);
nand U6572 (N_6572,N_4012,N_3885);
and U6573 (N_6573,N_4736,N_5490);
nand U6574 (N_6574,N_4045,N_3827);
and U6575 (N_6575,N_4662,N_4434);
xnor U6576 (N_6576,N_3707,N_5082);
or U6577 (N_6577,N_3060,N_4353);
nor U6578 (N_6578,N_4476,N_5183);
nand U6579 (N_6579,N_5305,N_5585);
nand U6580 (N_6580,N_4431,N_3423);
and U6581 (N_6581,N_4841,N_5886);
nand U6582 (N_6582,N_5477,N_3207);
xor U6583 (N_6583,N_3429,N_4307);
xor U6584 (N_6584,N_5038,N_3696);
or U6585 (N_6585,N_5549,N_3568);
nand U6586 (N_6586,N_4521,N_5189);
nand U6587 (N_6587,N_3362,N_4604);
or U6588 (N_6588,N_5713,N_3425);
nor U6589 (N_6589,N_3910,N_3091);
nand U6590 (N_6590,N_3940,N_4001);
xnor U6591 (N_6591,N_4849,N_3407);
xor U6592 (N_6592,N_5848,N_4876);
nand U6593 (N_6593,N_5376,N_4370);
and U6594 (N_6594,N_5985,N_3082);
and U6595 (N_6595,N_5374,N_4733);
nor U6596 (N_6596,N_4594,N_4337);
xnor U6597 (N_6597,N_4423,N_3757);
nand U6598 (N_6598,N_3645,N_4095);
xnor U6599 (N_6599,N_3604,N_5274);
nor U6600 (N_6600,N_3116,N_5772);
and U6601 (N_6601,N_5181,N_3839);
and U6602 (N_6602,N_5633,N_4505);
nor U6603 (N_6603,N_5211,N_3384);
or U6604 (N_6604,N_4305,N_3312);
xor U6605 (N_6605,N_4757,N_5102);
nand U6606 (N_6606,N_3635,N_4013);
or U6607 (N_6607,N_5781,N_3175);
nand U6608 (N_6608,N_5418,N_4832);
nor U6609 (N_6609,N_4426,N_3329);
nand U6610 (N_6610,N_3644,N_3613);
nand U6611 (N_6611,N_5779,N_3320);
xnor U6612 (N_6612,N_4677,N_5799);
and U6613 (N_6613,N_4692,N_3276);
nand U6614 (N_6614,N_5702,N_4877);
or U6615 (N_6615,N_4912,N_5092);
nor U6616 (N_6616,N_5951,N_5052);
xnor U6617 (N_6617,N_4316,N_3041);
xnor U6618 (N_6618,N_4707,N_3894);
and U6619 (N_6619,N_3964,N_4416);
or U6620 (N_6620,N_3535,N_5015);
and U6621 (N_6621,N_4249,N_5752);
nor U6622 (N_6622,N_4644,N_4824);
and U6623 (N_6623,N_4325,N_5368);
or U6624 (N_6624,N_4558,N_3443);
xor U6625 (N_6625,N_5590,N_5415);
nand U6626 (N_6626,N_4010,N_3426);
and U6627 (N_6627,N_3965,N_5892);
or U6628 (N_6628,N_5561,N_3477);
nand U6629 (N_6629,N_3932,N_5939);
or U6630 (N_6630,N_5907,N_4468);
and U6631 (N_6631,N_4113,N_5813);
nand U6632 (N_6632,N_5195,N_5245);
and U6633 (N_6633,N_5146,N_3039);
and U6634 (N_6634,N_5736,N_4936);
nor U6635 (N_6635,N_3695,N_3344);
or U6636 (N_6636,N_5837,N_3764);
or U6637 (N_6637,N_5335,N_3035);
and U6638 (N_6638,N_4850,N_3988);
nor U6639 (N_6639,N_5295,N_4208);
xnor U6640 (N_6640,N_3621,N_3947);
xor U6641 (N_6641,N_4150,N_4231);
xnor U6642 (N_6642,N_3323,N_3339);
nand U6643 (N_6643,N_3798,N_4637);
xnor U6644 (N_6644,N_5272,N_4991);
nor U6645 (N_6645,N_5565,N_3292);
xor U6646 (N_6646,N_3158,N_3118);
nand U6647 (N_6647,N_4069,N_4999);
and U6648 (N_6648,N_3961,N_3676);
or U6649 (N_6649,N_3672,N_3148);
xor U6650 (N_6650,N_3169,N_4459);
nand U6651 (N_6651,N_4664,N_5448);
nand U6652 (N_6652,N_3995,N_4580);
nand U6653 (N_6653,N_5227,N_4945);
nor U6654 (N_6654,N_4878,N_4918);
xnor U6655 (N_6655,N_3170,N_4366);
or U6656 (N_6656,N_3403,N_5366);
nand U6657 (N_6657,N_4572,N_5902);
xor U6658 (N_6658,N_3383,N_3776);
nand U6659 (N_6659,N_3725,N_5879);
nor U6660 (N_6660,N_5173,N_5674);
nor U6661 (N_6661,N_4911,N_5087);
and U6662 (N_6662,N_5184,N_4710);
nand U6663 (N_6663,N_4599,N_3132);
and U6664 (N_6664,N_5152,N_4530);
or U6665 (N_6665,N_5134,N_5994);
and U6666 (N_6666,N_4745,N_3356);
xnor U6667 (N_6667,N_3565,N_5096);
or U6668 (N_6668,N_4433,N_4153);
or U6669 (N_6669,N_5784,N_5423);
nand U6670 (N_6670,N_3209,N_3663);
or U6671 (N_6671,N_5037,N_3133);
or U6672 (N_6672,N_4794,N_5345);
xor U6673 (N_6673,N_4440,N_3852);
and U6674 (N_6674,N_3008,N_5696);
xnor U6675 (N_6675,N_4643,N_5324);
xnor U6676 (N_6676,N_4443,N_5160);
and U6677 (N_6677,N_4890,N_4392);
and U6678 (N_6678,N_5637,N_3070);
xnor U6679 (N_6679,N_5971,N_5682);
nor U6680 (N_6680,N_4104,N_3129);
xor U6681 (N_6681,N_3289,N_5776);
nor U6682 (N_6682,N_3336,N_3705);
and U6683 (N_6683,N_4411,N_5023);
and U6684 (N_6684,N_4309,N_3522);
and U6685 (N_6685,N_5520,N_3867);
xor U6686 (N_6686,N_4157,N_3163);
nand U6687 (N_6687,N_4154,N_3972);
or U6688 (N_6688,N_4866,N_5404);
nor U6689 (N_6689,N_5988,N_3840);
nand U6690 (N_6690,N_3461,N_3949);
or U6691 (N_6691,N_3618,N_4965);
xor U6692 (N_6692,N_4959,N_4155);
or U6693 (N_6693,N_5548,N_3286);
or U6694 (N_6694,N_3431,N_4494);
xor U6695 (N_6695,N_3110,N_4264);
nand U6696 (N_6696,N_5112,N_3265);
xnor U6697 (N_6697,N_5940,N_4089);
xnor U6698 (N_6698,N_4519,N_3688);
and U6699 (N_6699,N_3612,N_3739);
xnor U6700 (N_6700,N_3322,N_5896);
or U6701 (N_6701,N_3851,N_3999);
nor U6702 (N_6702,N_5036,N_3962);
nor U6703 (N_6703,N_4949,N_3837);
nand U6704 (N_6704,N_3907,N_4719);
nand U6705 (N_6705,N_4348,N_5083);
xnor U6706 (N_6706,N_5046,N_4658);
xor U6707 (N_6707,N_3592,N_4195);
xor U6708 (N_6708,N_4688,N_5871);
nor U6709 (N_6709,N_3777,N_3831);
xnor U6710 (N_6710,N_4146,N_3896);
or U6711 (N_6711,N_3825,N_3906);
nand U6712 (N_6712,N_3022,N_3424);
nor U6713 (N_6713,N_5588,N_5126);
nor U6714 (N_6714,N_4341,N_5334);
or U6715 (N_6715,N_3556,N_4751);
nand U6716 (N_6716,N_5751,N_4484);
or U6717 (N_6717,N_4252,N_5934);
or U6718 (N_6718,N_4014,N_5138);
xnor U6719 (N_6719,N_5480,N_4512);
nand U6720 (N_6720,N_4407,N_3243);
nand U6721 (N_6721,N_3563,N_4769);
xor U6722 (N_6722,N_5949,N_5226);
or U6723 (N_6723,N_4689,N_5911);
and U6724 (N_6724,N_3731,N_4805);
nor U6725 (N_6725,N_4270,N_5990);
or U6726 (N_6726,N_4552,N_3863);
nand U6727 (N_6727,N_4567,N_4979);
and U6728 (N_6728,N_4922,N_5004);
nor U6729 (N_6729,N_5922,N_3767);
and U6730 (N_6730,N_5243,N_4425);
or U6731 (N_6731,N_3602,N_3462);
xor U6732 (N_6732,N_3034,N_4716);
nor U6733 (N_6733,N_5390,N_4333);
xor U6734 (N_6734,N_4117,N_5122);
or U6735 (N_6735,N_5225,N_3354);
nor U6736 (N_6736,N_3301,N_4913);
nand U6737 (N_6737,N_3893,N_5882);
and U6738 (N_6738,N_4655,N_5287);
nor U6739 (N_6739,N_4207,N_5888);
and U6740 (N_6740,N_5666,N_4685);
xnor U6741 (N_6741,N_5574,N_3086);
xnor U6742 (N_6742,N_3321,N_3879);
nand U6743 (N_6743,N_5657,N_3210);
nor U6744 (N_6744,N_4925,N_3040);
nand U6745 (N_6745,N_3139,N_3710);
nand U6746 (N_6746,N_5818,N_3756);
nor U6747 (N_6747,N_3134,N_3559);
or U6748 (N_6748,N_5353,N_3589);
xor U6749 (N_6749,N_4787,N_3347);
xor U6750 (N_6750,N_4992,N_3496);
xnor U6751 (N_6751,N_5610,N_5034);
nor U6752 (N_6752,N_3001,N_4206);
or U6753 (N_6753,N_3928,N_3752);
or U6754 (N_6754,N_4862,N_3656);
and U6755 (N_6755,N_5357,N_5402);
and U6756 (N_6756,N_4386,N_5373);
and U6757 (N_6757,N_5997,N_4587);
and U6758 (N_6758,N_4843,N_5843);
nand U6759 (N_6759,N_4900,N_5767);
and U6760 (N_6760,N_4907,N_5805);
or U6761 (N_6761,N_3181,N_5504);
xnor U6762 (N_6762,N_3006,N_5701);
nor U6763 (N_6763,N_3980,N_4884);
nand U6764 (N_6764,N_3686,N_4121);
and U6765 (N_6765,N_5071,N_4063);
or U6766 (N_6766,N_4858,N_4815);
nor U6767 (N_6767,N_4365,N_4818);
and U6768 (N_6768,N_5101,N_3089);
and U6769 (N_6769,N_4828,N_5147);
xor U6770 (N_6770,N_5745,N_3157);
nand U6771 (N_6771,N_5043,N_4034);
and U6772 (N_6772,N_5275,N_4332);
xnor U6773 (N_6773,N_3145,N_4609);
nand U6774 (N_6774,N_3363,N_4758);
nor U6775 (N_6775,N_3119,N_4064);
and U6776 (N_6776,N_3067,N_3553);
nand U6777 (N_6777,N_3534,N_3422);
xor U6778 (N_6778,N_5953,N_3785);
nand U6779 (N_6779,N_3213,N_4465);
or U6780 (N_6780,N_5987,N_4463);
and U6781 (N_6781,N_3897,N_3458);
or U6782 (N_6782,N_5644,N_5669);
xor U6783 (N_6783,N_5903,N_3800);
and U6784 (N_6784,N_3922,N_5746);
nand U6785 (N_6785,N_3954,N_4605);
or U6786 (N_6786,N_3717,N_5123);
or U6787 (N_6787,N_4499,N_3516);
and U6788 (N_6788,N_4874,N_4730);
and U6789 (N_6789,N_3307,N_3084);
xor U6790 (N_6790,N_4026,N_5013);
or U6791 (N_6791,N_4460,N_4923);
xor U6792 (N_6792,N_4030,N_3294);
nand U6793 (N_6793,N_5923,N_3273);
nor U6794 (N_6794,N_4065,N_3834);
nor U6795 (N_6795,N_4255,N_5363);
or U6796 (N_6796,N_5684,N_5568);
xnor U6797 (N_6797,N_4453,N_3010);
nand U6798 (N_6798,N_4803,N_4148);
xor U6799 (N_6799,N_3138,N_4449);
or U6800 (N_6800,N_3889,N_5705);
xor U6801 (N_6801,N_3474,N_4492);
nand U6802 (N_6802,N_3353,N_4202);
nor U6803 (N_6803,N_5500,N_3297);
and U6804 (N_6804,N_3221,N_3763);
nand U6805 (N_6805,N_3524,N_3841);
nand U6806 (N_6806,N_4845,N_4671);
xnor U6807 (N_6807,N_3578,N_5513);
xor U6808 (N_6808,N_3805,N_3455);
or U6809 (N_6809,N_5362,N_3025);
nand U6810 (N_6810,N_5796,N_5798);
or U6811 (N_6811,N_5167,N_5606);
xor U6812 (N_6812,N_4694,N_5958);
xnor U6813 (N_6813,N_3270,N_3611);
and U6814 (N_6814,N_4105,N_3011);
and U6815 (N_6815,N_5257,N_4025);
nor U6816 (N_6816,N_3377,N_4226);
or U6817 (N_6817,N_3743,N_4600);
nand U6818 (N_6818,N_5284,N_5331);
nor U6819 (N_6819,N_3690,N_5826);
and U6820 (N_6820,N_5056,N_5462);
nor U6821 (N_6821,N_5182,N_3584);
nand U6822 (N_6822,N_5708,N_5662);
nor U6823 (N_6823,N_5597,N_4051);
or U6824 (N_6824,N_5109,N_3833);
xnor U6825 (N_6825,N_3667,N_3029);
xor U6826 (N_6826,N_3801,N_3975);
xor U6827 (N_6827,N_4381,N_3026);
nor U6828 (N_6828,N_5413,N_5089);
xnor U6829 (N_6829,N_5155,N_5698);
xor U6830 (N_6830,N_5045,N_3783);
nor U6831 (N_6831,N_3172,N_5626);
xor U6832 (N_6832,N_5268,N_3640);
or U6833 (N_6833,N_5317,N_3519);
or U6834 (N_6834,N_3950,N_5470);
xnor U6835 (N_6835,N_3005,N_3982);
nand U6836 (N_6836,N_4569,N_3945);
nor U6837 (N_6837,N_4963,N_3646);
and U6838 (N_6838,N_4211,N_3000);
nor U6839 (N_6839,N_4189,N_4317);
or U6840 (N_6840,N_3642,N_3585);
nor U6841 (N_6841,N_4364,N_3890);
nand U6842 (N_6842,N_5832,N_5960);
xor U6843 (N_6843,N_5981,N_4873);
or U6844 (N_6844,N_5754,N_5553);
and U6845 (N_6845,N_4715,N_5007);
nand U6846 (N_6846,N_3327,N_3076);
nand U6847 (N_6847,N_3934,N_3884);
and U6848 (N_6848,N_4219,N_3502);
and U6849 (N_6849,N_3437,N_4435);
nor U6850 (N_6850,N_4882,N_3397);
or U6851 (N_6851,N_5360,N_4550);
nand U6852 (N_6852,N_5572,N_3520);
nor U6853 (N_6853,N_3661,N_3330);
and U6854 (N_6854,N_5906,N_5821);
and U6855 (N_6855,N_5131,N_5947);
nor U6856 (N_6856,N_5074,N_5078);
or U6857 (N_6857,N_3628,N_5768);
nand U6858 (N_6858,N_5378,N_5944);
and U6859 (N_6859,N_5950,N_3064);
and U6860 (N_6860,N_4556,N_4280);
or U6861 (N_6861,N_3166,N_4638);
and U6862 (N_6862,N_4663,N_5841);
or U6863 (N_6863,N_3493,N_3247);
xor U6864 (N_6864,N_5459,N_4256);
nand U6865 (N_6865,N_3037,N_5931);
nand U6866 (N_6866,N_3228,N_3432);
or U6867 (N_6867,N_4743,N_4003);
nand U6868 (N_6868,N_3054,N_4292);
nor U6869 (N_6869,N_5899,N_5429);
nand U6870 (N_6870,N_4151,N_4004);
or U6871 (N_6871,N_4542,N_4204);
xor U6872 (N_6872,N_5918,N_4982);
nand U6873 (N_6873,N_5228,N_5627);
nand U6874 (N_6874,N_4090,N_5999);
nand U6875 (N_6875,N_3727,N_5946);
nor U6876 (N_6876,N_5369,N_5658);
and U6877 (N_6877,N_4437,N_5794);
or U6878 (N_6878,N_3669,N_5534);
nor U6879 (N_6879,N_5617,N_5895);
nand U6880 (N_6880,N_5901,N_3358);
nor U6881 (N_6881,N_3636,N_5168);
or U6882 (N_6882,N_4790,N_5640);
or U6883 (N_6883,N_5494,N_5573);
xor U6884 (N_6884,N_4303,N_4087);
and U6885 (N_6885,N_5469,N_3823);
or U6886 (N_6886,N_4288,N_3970);
nand U6887 (N_6887,N_3533,N_5749);
or U6888 (N_6888,N_3860,N_3809);
nor U6889 (N_6889,N_4676,N_5804);
or U6890 (N_6890,N_3566,N_5970);
nor U6891 (N_6891,N_3979,N_3438);
nand U6892 (N_6892,N_5140,N_5214);
or U6893 (N_6893,N_5917,N_3251);
nand U6894 (N_6894,N_3266,N_5005);
xnor U6895 (N_6895,N_4263,N_3016);
nand U6896 (N_6896,N_5594,N_3541);
nor U6897 (N_6897,N_3355,N_3791);
and U6898 (N_6898,N_4532,N_4763);
nor U6899 (N_6899,N_3044,N_4403);
and U6900 (N_6900,N_5229,N_4994);
nand U6901 (N_6901,N_5306,N_3786);
or U6902 (N_6902,N_4608,N_3668);
or U6903 (N_6903,N_5359,N_5110);
and U6904 (N_6904,N_5543,N_3106);
and U6905 (N_6905,N_3314,N_4076);
and U6906 (N_6906,N_4620,N_5628);
nand U6907 (N_6907,N_4865,N_3692);
nor U6908 (N_6908,N_5730,N_5825);
or U6909 (N_6909,N_3302,N_3352);
nand U6910 (N_6910,N_4125,N_4821);
and U6911 (N_6911,N_3392,N_5432);
nand U6912 (N_6912,N_3417,N_5982);
xnor U6913 (N_6913,N_3765,N_4996);
nand U6914 (N_6914,N_4697,N_3126);
or U6915 (N_6915,N_5201,N_3130);
xnor U6916 (N_6916,N_3101,N_5527);
nand U6917 (N_6917,N_5897,N_4848);
xnor U6918 (N_6918,N_3098,N_4137);
and U6919 (N_6919,N_5213,N_5858);
xnor U6920 (N_6920,N_3728,N_5466);
nor U6921 (N_6921,N_4931,N_4526);
xor U6922 (N_6922,N_4092,N_4667);
and U6923 (N_6923,N_5671,N_4274);
and U6924 (N_6924,N_4391,N_5967);
xor U6925 (N_6925,N_3096,N_4835);
nand U6926 (N_6926,N_5533,N_5320);
xnor U6927 (N_6927,N_5011,N_3186);
xnor U6928 (N_6928,N_3264,N_4799);
or U6929 (N_6929,N_3569,N_4462);
or U6930 (N_6930,N_3180,N_4898);
nand U6931 (N_6931,N_5017,N_4696);
or U6932 (N_6932,N_3719,N_3466);
and U6933 (N_6933,N_3835,N_4575);
xnor U6934 (N_6934,N_4579,N_5734);
and U6935 (N_6935,N_5732,N_4217);
xor U6936 (N_6936,N_3430,N_3882);
and U6937 (N_6937,N_4590,N_5434);
or U6938 (N_6938,N_4334,N_3718);
and U6939 (N_6939,N_4946,N_5431);
and U6940 (N_6940,N_3017,N_4021);
nand U6941 (N_6941,N_5105,N_4940);
nor U6942 (N_6942,N_3740,N_5276);
or U6943 (N_6943,N_5766,N_3778);
nor U6944 (N_6944,N_5236,N_4654);
and U6945 (N_6945,N_4725,N_4700);
xor U6946 (N_6946,N_4178,N_3156);
and U6947 (N_6947,N_4401,N_5057);
nor U6948 (N_6948,N_4352,N_5377);
and U6949 (N_6949,N_3200,N_5600);
nand U6950 (N_6950,N_3844,N_3281);
or U6951 (N_6951,N_3445,N_3244);
nand U6952 (N_6952,N_3572,N_4816);
and U6953 (N_6953,N_5748,N_5081);
or U6954 (N_6954,N_3486,N_4917);
xor U6955 (N_6955,N_4011,N_3189);
or U6956 (N_6956,N_3049,N_4527);
nand U6957 (N_6957,N_3759,N_5865);
xnor U6958 (N_6958,N_4968,N_4622);
or U6959 (N_6959,N_3547,N_5785);
or U6960 (N_6960,N_5252,N_4904);
or U6961 (N_6961,N_4029,N_3236);
nor U6962 (N_6962,N_5571,N_4083);
or U6963 (N_6963,N_4916,N_5148);
and U6964 (N_6964,N_3250,N_4414);
and U6965 (N_6965,N_3951,N_3811);
and U6966 (N_6966,N_4186,N_4932);
xor U6967 (N_6967,N_5424,N_4324);
and U6968 (N_6968,N_4619,N_4362);
or U6969 (N_6969,N_4955,N_4515);
or U6970 (N_6970,N_5125,N_4019);
or U6971 (N_6971,N_5124,N_4248);
and U6972 (N_6972,N_4981,N_4933);
or U6973 (N_6973,N_4130,N_3976);
and U6974 (N_6974,N_4872,N_5311);
nor U6975 (N_6975,N_3348,N_3782);
nand U6976 (N_6976,N_4005,N_5716);
nand U6977 (N_6977,N_5388,N_4770);
xor U6978 (N_6978,N_5593,N_4538);
and U6979 (N_6979,N_3819,N_4046);
nor U6980 (N_6980,N_3095,N_3577);
or U6981 (N_6981,N_3794,N_3201);
xor U6982 (N_6982,N_3442,N_3456);
and U6983 (N_6983,N_5205,N_5717);
xnor U6984 (N_6984,N_3188,N_3092);
and U6985 (N_6985,N_5435,N_5683);
and U6986 (N_6986,N_3824,N_5726);
or U6987 (N_6987,N_4184,N_4243);
or U6988 (N_6988,N_5411,N_5582);
and U6989 (N_6989,N_3036,N_5051);
or U6990 (N_6990,N_5530,N_3868);
xor U6991 (N_6991,N_3651,N_4409);
xor U6992 (N_6992,N_3316,N_3574);
or U6993 (N_6993,N_4285,N_4650);
nand U6994 (N_6994,N_4050,N_4085);
nand U6995 (N_6995,N_4223,N_4043);
or U6996 (N_6996,N_3774,N_4404);
nor U6997 (N_6997,N_5456,N_5604);
xor U6998 (N_6998,N_5584,N_3305);
nor U6999 (N_6999,N_4236,N_4611);
nand U7000 (N_7000,N_3968,N_4093);
or U7001 (N_7001,N_5251,N_5258);
or U7002 (N_7002,N_3107,N_3023);
nand U7003 (N_7003,N_5401,N_4801);
xor U7004 (N_7004,N_3490,N_4458);
xnor U7005 (N_7005,N_5639,N_5414);
and U7006 (N_7006,N_5555,N_4523);
nand U7007 (N_7007,N_5054,N_5393);
and U7008 (N_7008,N_4229,N_4447);
and U7009 (N_7009,N_5870,N_4964);
and U7010 (N_7010,N_4939,N_5887);
and U7011 (N_7011,N_3472,N_4165);
nor U7012 (N_7012,N_3203,N_4354);
nor U7013 (N_7013,N_4306,N_4749);
xor U7014 (N_7014,N_5203,N_5855);
or U7015 (N_7015,N_3306,N_4772);
or U7016 (N_7016,N_4533,N_5006);
nor U7017 (N_7017,N_4645,N_3591);
xor U7018 (N_7018,N_5392,N_5055);
xnor U7019 (N_7019,N_4997,N_3660);
or U7020 (N_7020,N_3171,N_3315);
nor U7021 (N_7021,N_5164,N_4672);
and U7022 (N_7022,N_5279,N_5968);
nor U7023 (N_7023,N_3677,N_3069);
xor U7024 (N_7024,N_3601,N_5544);
xor U7025 (N_7025,N_3813,N_5120);
or U7026 (N_7026,N_4583,N_4867);
xnor U7027 (N_7027,N_5869,N_5926);
nor U7028 (N_7028,N_4938,N_3051);
or U7029 (N_7029,N_4068,N_4589);
nand U7030 (N_7030,N_4852,N_3046);
nand U7031 (N_7031,N_3664,N_5449);
and U7032 (N_7032,N_4314,N_5545);
nand U7033 (N_7033,N_4177,N_5973);
nand U7034 (N_7034,N_4136,N_3052);
nor U7035 (N_7035,N_4038,N_4474);
or U7036 (N_7036,N_5881,N_5695);
xor U7037 (N_7037,N_4978,N_4641);
nand U7038 (N_7038,N_3769,N_4082);
nor U7039 (N_7039,N_4566,N_4742);
and U7040 (N_7040,N_3003,N_3736);
or U7041 (N_7041,N_5426,N_4221);
xor U7042 (N_7042,N_5473,N_4389);
nand U7043 (N_7043,N_4351,N_3866);
or U7044 (N_7044,N_5118,N_3065);
and U7045 (N_7045,N_3267,N_5952);
and U7046 (N_7046,N_4682,N_5720);
and U7047 (N_7047,N_5190,N_4827);
or U7048 (N_7048,N_3750,N_5039);
nand U7049 (N_7049,N_4152,N_5550);
xor U7050 (N_7050,N_5020,N_5630);
nand U7051 (N_7051,N_3909,N_3738);
or U7052 (N_7052,N_4800,N_3760);
xnor U7053 (N_7053,N_3508,N_5797);
nand U7054 (N_7054,N_3399,N_5509);
and U7055 (N_7055,N_4840,N_3185);
nor U7056 (N_7056,N_5149,N_3990);
or U7057 (N_7057,N_5823,N_5040);
nand U7058 (N_7058,N_3471,N_5370);
nand U7059 (N_7059,N_3032,N_5231);
xor U7060 (N_7060,N_5884,N_4214);
nor U7061 (N_7061,N_5012,N_4892);
and U7062 (N_7062,N_4951,N_5247);
nor U7063 (N_7063,N_3114,N_5636);
xor U7064 (N_7064,N_5303,N_4976);
nor U7065 (N_7065,N_4271,N_5777);
nand U7066 (N_7066,N_5840,N_3848);
and U7067 (N_7067,N_3382,N_4625);
nand U7068 (N_7068,N_3482,N_4216);
xnor U7069 (N_7069,N_5485,N_4373);
and U7070 (N_7070,N_5178,N_5706);
or U7071 (N_7071,N_5980,N_3412);
xor U7072 (N_7072,N_3326,N_4984);
and U7073 (N_7073,N_4804,N_3631);
and U7074 (N_7074,N_5921,N_5438);
or U7075 (N_7075,N_4183,N_5811);
nor U7076 (N_7076,N_4778,N_5310);
nand U7077 (N_7077,N_4920,N_3436);
xor U7078 (N_7078,N_5119,N_5676);
and U7079 (N_7079,N_4086,N_3974);
or U7080 (N_7080,N_4357,N_3828);
nor U7081 (N_7081,N_3504,N_5913);
or U7082 (N_7082,N_3986,N_3028);
nor U7083 (N_7083,N_5632,N_4734);
and U7084 (N_7084,N_5853,N_4905);
xnor U7085 (N_7085,N_5249,N_4343);
nand U7086 (N_7086,N_5294,N_3366);
or U7087 (N_7087,N_5412,N_4210);
nor U7088 (N_7088,N_4132,N_4739);
and U7089 (N_7089,N_3742,N_5180);
and U7090 (N_7090,N_3943,N_4345);
and U7091 (N_7091,N_5333,N_5064);
or U7092 (N_7092,N_5889,N_3573);
or U7093 (N_7093,N_5679,N_5304);
nor U7094 (N_7094,N_5941,N_5496);
nand U7095 (N_7095,N_5220,N_4764);
xor U7096 (N_7096,N_5612,N_5151);
xnor U7097 (N_7097,N_5788,N_4975);
or U7098 (N_7098,N_5224,N_5647);
or U7099 (N_7099,N_3380,N_4222);
or U7100 (N_7100,N_3088,N_3650);
or U7101 (N_7101,N_4937,N_3498);
xnor U7102 (N_7102,N_5486,N_5019);
or U7103 (N_7103,N_4190,N_5352);
nand U7104 (N_7104,N_5460,N_4591);
nand U7105 (N_7105,N_4075,N_5943);
and U7106 (N_7106,N_5514,N_4656);
and U7107 (N_7107,N_4674,N_3120);
nand U7108 (N_7108,N_5127,N_5873);
or U7109 (N_7109,N_3050,N_3937);
nor U7110 (N_7110,N_4042,N_4461);
nand U7111 (N_7111,N_5689,N_4245);
or U7112 (N_7112,N_5552,N_3020);
nor U7113 (N_7113,N_3102,N_3249);
and U7114 (N_7114,N_5567,N_3606);
nor U7115 (N_7115,N_4711,N_4559);
and U7116 (N_7116,N_3627,N_3704);
and U7117 (N_7117,N_3699,N_3908);
and U7118 (N_7118,N_4864,N_4109);
nand U7119 (N_7119,N_3859,N_5314);
nand U7120 (N_7120,N_5839,N_3497);
xor U7121 (N_7121,N_4588,N_5267);
xor U7122 (N_7122,N_5620,N_4016);
and U7123 (N_7123,N_5915,N_5809);
and U7124 (N_7124,N_5250,N_5936);
and U7125 (N_7125,N_5493,N_3888);
xor U7126 (N_7126,N_5328,N_4033);
xnor U7127 (N_7127,N_3015,N_4410);
and U7128 (N_7128,N_4780,N_3815);
and U7129 (N_7129,N_3779,N_4657);
nand U7130 (N_7130,N_4910,N_3021);
and U7131 (N_7131,N_4293,N_5098);
or U7132 (N_7132,N_4603,N_5443);
or U7133 (N_7133,N_5407,N_3509);
nand U7134 (N_7134,N_5169,N_3176);
or U7135 (N_7135,N_3634,N_3931);
and U7136 (N_7136,N_4181,N_4765);
xor U7137 (N_7137,N_5613,N_4861);
nor U7138 (N_7138,N_4006,N_5347);
and U7139 (N_7139,N_4698,N_3855);
or U7140 (N_7140,N_4581,N_5883);
nand U7141 (N_7141,N_4930,N_3427);
nor U7142 (N_7142,N_5384,N_4738);
nand U7143 (N_7143,N_3439,N_4077);
nand U7144 (N_7144,N_3744,N_5157);
xnor U7145 (N_7145,N_5654,N_4760);
xnor U7146 (N_7146,N_3543,N_5218);
or U7147 (N_7147,N_3211,N_4610);
or U7148 (N_7148,N_4031,N_3123);
xor U7149 (N_7149,N_5880,N_5700);
nor U7150 (N_7150,N_3154,N_4055);
xor U7151 (N_7151,N_4529,N_5471);
nor U7152 (N_7152,N_4517,N_4259);
and U7153 (N_7153,N_5795,N_4272);
nand U7154 (N_7154,N_4268,N_4987);
xnor U7155 (N_7155,N_3729,N_5875);
nand U7156 (N_7156,N_3567,N_5731);
and U7157 (N_7157,N_3268,N_4385);
nand U7158 (N_7158,N_4885,N_3587);
nand U7159 (N_7159,N_5615,N_5309);
nor U7160 (N_7160,N_3545,N_5405);
and U7161 (N_7161,N_4886,N_4387);
or U7162 (N_7162,N_3678,N_5673);
or U7163 (N_7163,N_4439,N_4897);
nand U7164 (N_7164,N_3219,N_5033);
nor U7165 (N_7165,N_4133,N_5690);
or U7166 (N_7166,N_4485,N_4889);
and U7167 (N_7167,N_3475,N_5387);
nor U7168 (N_7168,N_3159,N_4735);
nand U7169 (N_7169,N_4941,N_3854);
and U7170 (N_7170,N_4524,N_3918);
and U7171 (N_7171,N_4761,N_5041);
and U7172 (N_7172,N_3402,N_3530);
nor U7173 (N_7173,N_3055,N_4648);
xnor U7174 (N_7174,N_4679,N_5139);
nand U7175 (N_7175,N_4927,N_3588);
nor U7176 (N_7176,N_3488,N_4158);
or U7177 (N_7177,N_4323,N_5523);
xor U7178 (N_7178,N_5532,N_4049);
nand U7179 (N_7179,N_3258,N_5845);
xor U7180 (N_7180,N_3967,N_5687);
nor U7181 (N_7181,N_4084,N_3002);
or U7182 (N_7182,N_4138,N_4731);
or U7183 (N_7183,N_5446,N_5165);
nor U7184 (N_7184,N_5461,N_5133);
xor U7185 (N_7185,N_4573,N_4378);
or U7186 (N_7186,N_5342,N_4488);
and U7187 (N_7187,N_5420,N_4894);
nand U7188 (N_7188,N_3925,N_3117);
and U7189 (N_7189,N_3223,N_3293);
or U7190 (N_7190,N_5977,N_4330);
and U7191 (N_7191,N_4704,N_3441);
or U7192 (N_7192,N_3807,N_4156);
or U7193 (N_7193,N_3915,N_3280);
nand U7194 (N_7194,N_4501,N_5747);
xnor U7195 (N_7195,N_4714,N_4129);
or U7196 (N_7196,N_5442,N_3047);
or U7197 (N_7197,N_5487,N_5753);
xnor U7198 (N_7198,N_3571,N_4367);
or U7199 (N_7199,N_4251,N_3068);
and U7200 (N_7200,N_3468,N_3874);
xnor U7201 (N_7201,N_3605,N_3924);
and U7202 (N_7202,N_5425,N_3290);
and U7203 (N_7203,N_4668,N_4128);
nand U7204 (N_7204,N_4691,N_4934);
nand U7205 (N_7205,N_3140,N_3500);
or U7206 (N_7206,N_3963,N_3340);
xnor U7207 (N_7207,N_4839,N_5242);
xor U7208 (N_7208,N_5269,N_4598);
or U7209 (N_7209,N_5076,N_3590);
or U7210 (N_7210,N_4419,N_3723);
or U7211 (N_7211,N_4278,N_5890);
and U7212 (N_7212,N_4359,N_3817);
and U7213 (N_7213,N_4331,N_5238);
nand U7214 (N_7214,N_3952,N_3853);
or U7215 (N_7215,N_4614,N_3561);
nor U7216 (N_7216,N_3045,N_5783);
and U7217 (N_7217,N_5044,N_4666);
xor U7218 (N_7218,N_4548,N_5755);
nor U7219 (N_7219,N_5942,N_4187);
nor U7220 (N_7220,N_4990,N_5216);
and U7221 (N_7221,N_4947,N_3788);
nand U7222 (N_7222,N_5715,N_4942);
nor U7223 (N_7223,N_4592,N_3507);
or U7224 (N_7224,N_5016,N_3371);
xor U7225 (N_7225,N_4481,N_4670);
and U7226 (N_7226,N_3212,N_4289);
nand U7227 (N_7227,N_5846,N_5603);
xnor U7228 (N_7228,N_4985,N_3878);
nand U7229 (N_7229,N_3720,N_5838);
and U7230 (N_7230,N_3222,N_3666);
nand U7231 (N_7231,N_4717,N_3579);
nand U7232 (N_7232,N_4565,N_3599);
or U7233 (N_7233,N_5365,N_3784);
nand U7234 (N_7234,N_3283,N_3090);
and U7235 (N_7235,N_5498,N_5135);
and U7236 (N_7236,N_5296,N_3724);
nor U7237 (N_7237,N_4722,N_5693);
and U7238 (N_7238,N_4430,N_3768);
nor U7239 (N_7239,N_4971,N_4627);
or U7240 (N_7240,N_5293,N_3400);
or U7241 (N_7241,N_3387,N_3115);
and U7242 (N_7242,N_5379,N_5240);
xnor U7243 (N_7243,N_5166,N_4032);
nor U7244 (N_7244,N_5419,N_3741);
xnor U7245 (N_7245,N_3700,N_4350);
xnor U7246 (N_7246,N_3359,N_3580);
xnor U7247 (N_7247,N_5073,N_4234);
nand U7248 (N_7248,N_4471,N_5515);
nor U7249 (N_7249,N_3194,N_5117);
or U7250 (N_7250,N_5623,N_5554);
and U7251 (N_7251,N_3122,N_4159);
and U7252 (N_7252,N_4723,N_5569);
and U7253 (N_7253,N_5964,N_4616);
nand U7254 (N_7254,N_3708,N_4415);
xor U7255 (N_7255,N_5743,N_4684);
nand U7256 (N_7256,N_4825,N_3609);
xor U7257 (N_7257,N_4124,N_4652);
nand U7258 (N_7258,N_5174,N_4943);
and U7259 (N_7259,N_5599,N_5383);
nand U7260 (N_7260,N_4509,N_4269);
or U7261 (N_7261,N_5299,N_3246);
nor U7262 (N_7262,N_4230,N_3197);
and U7263 (N_7263,N_5158,N_3754);
xor U7264 (N_7264,N_5771,N_5114);
nand U7265 (N_7265,N_5711,N_4361);
nor U7266 (N_7266,N_3410,N_5111);
or U7267 (N_7267,N_4661,N_3575);
or U7268 (N_7268,N_4360,N_4000);
nor U7269 (N_7269,N_4750,N_5358);
or U7270 (N_7270,N_5827,N_5478);
and U7271 (N_7271,N_5831,N_5095);
nand U7272 (N_7272,N_4283,N_5137);
xor U7273 (N_7273,N_5481,N_5175);
xnor U7274 (N_7274,N_3939,N_5560);
or U7275 (N_7275,N_3643,N_3401);
or U7276 (N_7276,N_5191,N_4355);
or U7277 (N_7277,N_3103,N_3078);
nand U7278 (N_7278,N_3075,N_5898);
or U7279 (N_7279,N_4483,N_4372);
and U7280 (N_7280,N_3495,N_3389);
xnor U7281 (N_7281,N_4647,N_5638);
or U7282 (N_7282,N_4774,N_3408);
xor U7283 (N_7283,N_4669,N_3227);
nor U7284 (N_7284,N_4851,N_3259);
and U7285 (N_7285,N_4516,N_4630);
xor U7286 (N_7286,N_4781,N_4543);
nor U7287 (N_7287,N_5697,N_3550);
and U7288 (N_7288,N_3487,N_3829);
nand U7289 (N_7289,N_4537,N_3891);
nor U7290 (N_7290,N_5956,N_3583);
nor U7291 (N_7291,N_5912,N_3420);
nor U7292 (N_7292,N_4020,N_3465);
xnor U7293 (N_7293,N_4613,N_4215);
nand U7294 (N_7294,N_4493,N_4299);
xor U7295 (N_7295,N_3846,N_5261);
and U7296 (N_7296,N_5406,N_5856);
nor U7297 (N_7297,N_5864,N_3518);
xor U7298 (N_7298,N_4310,N_4228);
nor U7299 (N_7299,N_4690,N_5318);
nor U7300 (N_7300,N_3849,N_3506);
and U7301 (N_7301,N_5116,N_5546);
nor U7302 (N_7302,N_5492,N_5265);
and U7303 (N_7303,N_5348,N_4203);
xor U7304 (N_7304,N_3536,N_4039);
nor U7305 (N_7305,N_3224,N_5010);
xor U7306 (N_7306,N_5097,N_3459);
xnor U7307 (N_7307,N_4479,N_4727);
or U7308 (N_7308,N_3904,N_5622);
nand U7309 (N_7309,N_4294,N_4368);
nand U7310 (N_7310,N_3616,N_5537);
xor U7311 (N_7311,N_4831,N_4640);
and U7312 (N_7312,N_4024,N_5372);
and U7313 (N_7313,N_5199,N_5975);
or U7314 (N_7314,N_4560,N_4507);
nor U7315 (N_7315,N_5680,N_4977);
xnor U7316 (N_7316,N_3989,N_4110);
nor U7317 (N_7317,N_4170,N_4771);
or U7318 (N_7318,N_3637,N_4073);
nor U7319 (N_7319,N_4686,N_4683);
nand U7320 (N_7320,N_4584,N_4601);
xnor U7321 (N_7321,N_3058,N_3948);
xnor U7322 (N_7322,N_4135,N_4536);
and U7323 (N_7323,N_5957,N_5891);
and U7324 (N_7324,N_4844,N_3470);
and U7325 (N_7325,N_4795,N_5874);
nand U7326 (N_7326,N_5278,N_3687);
nand U7327 (N_7327,N_3253,N_5503);
or U7328 (N_7328,N_3689,N_5313);
and U7329 (N_7329,N_4081,N_3014);
xnor U7330 (N_7330,N_4621,N_5589);
nor U7331 (N_7331,N_5028,N_3214);
nand U7332 (N_7332,N_3453,N_3033);
xor U7333 (N_7333,N_4732,N_4496);
nor U7334 (N_7334,N_5773,N_5651);
or U7335 (N_7335,N_4327,N_3394);
xnor U7336 (N_7336,N_3515,N_4478);
nand U7337 (N_7337,N_3136,N_5396);
and U7338 (N_7338,N_4166,N_4721);
nor U7339 (N_7339,N_4108,N_3131);
or U7340 (N_7340,N_3240,N_4441);
and U7341 (N_7341,N_5927,N_5851);
nor U7342 (N_7342,N_3398,N_3004);
and U7343 (N_7343,N_3147,N_5756);
nand U7344 (N_7344,N_3414,N_5955);
and U7345 (N_7345,N_5621,N_4205);
and U7346 (N_7346,N_4809,N_3252);
and U7347 (N_7347,N_4119,N_3789);
or U7348 (N_7348,N_4197,N_3262);
nor U7349 (N_7349,N_5540,N_5812);
xnor U7350 (N_7350,N_5144,N_4147);
and U7351 (N_7351,N_4091,N_4659);
and U7352 (N_7352,N_5566,N_3063);
nand U7353 (N_7353,N_3079,N_5115);
and U7354 (N_7354,N_4213,N_5025);
and U7355 (N_7355,N_5280,N_5526);
nand U7356 (N_7356,N_3113,N_5232);
nor U7357 (N_7357,N_4131,N_5452);
nor U7358 (N_7358,N_4098,N_3433);
or U7359 (N_7359,N_3031,N_5725);
nand U7360 (N_7360,N_3331,N_4506);
nand U7361 (N_7361,N_4570,N_3843);
nand U7362 (N_7362,N_5760,N_5570);
xnor U7363 (N_7363,N_5030,N_5441);
or U7364 (N_7364,N_3941,N_3379);
and U7365 (N_7365,N_5002,N_3463);
xor U7366 (N_7366,N_5993,N_5059);
xor U7367 (N_7367,N_5518,N_5103);
nor U7368 (N_7368,N_4319,N_5675);
nor U7369 (N_7369,N_4810,N_5536);
nand U7370 (N_7370,N_3409,N_5577);
nand U7371 (N_7371,N_3275,N_4718);
xnor U7372 (N_7372,N_4428,N_5850);
or U7373 (N_7373,N_5963,N_4141);
nand U7374 (N_7374,N_3927,N_3104);
and U7375 (N_7375,N_4500,N_5270);
nor U7376 (N_7376,N_5014,N_4812);
or U7377 (N_7377,N_3797,N_5479);
xnor U7378 (N_7378,N_5325,N_5877);
nor U7379 (N_7379,N_4514,N_5670);
xor U7380 (N_7380,N_5106,N_4120);
nand U7381 (N_7381,N_4525,N_5714);
xor U7382 (N_7382,N_4564,N_5259);
xnor U7383 (N_7383,N_4902,N_5718);
xnor U7384 (N_7384,N_5791,N_5645);
and U7385 (N_7385,N_4123,N_5542);
and U7386 (N_7386,N_3531,N_5079);
nand U7387 (N_7387,N_3304,N_4544);
or U7388 (N_7388,N_5230,N_5609);
nand U7389 (N_7389,N_4040,N_4713);
and U7390 (N_7390,N_3734,N_3523);
xor U7391 (N_7391,N_5291,N_3256);
nand U7392 (N_7392,N_4022,N_5709);
xnor U7393 (N_7393,N_5738,N_4041);
xnor U7394 (N_7394,N_3257,N_4633);
nor U7395 (N_7395,N_3775,N_5061);
nor U7396 (N_7396,N_4277,N_3434);
nand U7397 (N_7397,N_3755,N_5650);
xor U7398 (N_7398,N_3905,N_5893);
nor U7399 (N_7399,N_4547,N_4145);
nand U7400 (N_7400,N_5712,N_5453);
and U7401 (N_7401,N_4436,N_4237);
nand U7402 (N_7402,N_4822,N_4783);
nand U7403 (N_7403,N_4602,N_4528);
nor U7404 (N_7404,N_4106,N_3726);
xor U7405 (N_7405,N_5984,N_3232);
nor U7406 (N_7406,N_3328,N_4412);
or U7407 (N_7407,N_4322,N_3984);
or U7408 (N_7408,N_4615,N_4883);
xor U7409 (N_7409,N_5643,N_3552);
or U7410 (N_7410,N_3781,N_3712);
or U7411 (N_7411,N_5598,N_3936);
or U7412 (N_7412,N_3230,N_4161);
and U7413 (N_7413,N_5962,N_3085);
nand U7414 (N_7414,N_5332,N_3517);
and U7415 (N_7415,N_3341,N_4066);
and U7416 (N_7416,N_5290,N_5185);
and U7417 (N_7417,N_3308,N_5292);
nor U7418 (N_7418,N_5859,N_4762);
nor U7419 (N_7419,N_3546,N_5930);
xor U7420 (N_7420,N_3324,N_3335);
nand U7421 (N_7421,N_5507,N_4028);
xnor U7422 (N_7422,N_4860,N_4574);
nand U7423 (N_7423,N_3012,N_5062);
or U7424 (N_7424,N_5758,N_4813);
nand U7425 (N_7425,N_3225,N_4954);
nor U7426 (N_7426,N_4741,N_4398);
nor U7427 (N_7427,N_4948,N_4752);
nand U7428 (N_7428,N_3938,N_4047);
or U7429 (N_7429,N_3160,N_4748);
xor U7430 (N_7430,N_5815,N_5099);
and U7431 (N_7431,N_3821,N_4212);
and U7432 (N_7432,N_5661,N_3594);
or U7433 (N_7433,N_5437,N_4281);
nand U7434 (N_7434,N_4107,N_5003);
nand U7435 (N_7435,N_5410,N_3532);
nor U7436 (N_7436,N_3350,N_4993);
nor U7437 (N_7437,N_5193,N_3501);
nand U7438 (N_7438,N_5909,N_4097);
xnor U7439 (N_7439,N_3097,N_3161);
and U7440 (N_7440,N_5000,N_4371);
nand U7441 (N_7441,N_5551,N_4257);
xnor U7442 (N_7442,N_4276,N_3285);
or U7443 (N_7443,N_3558,N_3345);
and U7444 (N_7444,N_3761,N_4869);
xor U7445 (N_7445,N_4167,N_5664);
and U7446 (N_7446,N_4773,N_5835);
and U7447 (N_7447,N_5954,N_4220);
nand U7448 (N_7448,N_4989,N_3419);
or U7449 (N_7449,N_4847,N_3538);
nor U7450 (N_7450,N_3300,N_4859);
or U7451 (N_7451,N_3680,N_4950);
nor U7452 (N_7452,N_4122,N_4168);
and U7453 (N_7453,N_5524,N_4703);
nor U7454 (N_7454,N_5186,N_4397);
or U7455 (N_7455,N_3109,N_4729);
nor U7456 (N_7456,N_4115,N_3822);
nand U7457 (N_7457,N_3693,N_4623);
and U7458 (N_7458,N_5995,N_5488);
xor U7459 (N_7459,N_3077,N_5667);
or U7460 (N_7460,N_4541,N_5009);
xnor U7461 (N_7461,N_5188,N_3318);
nor U7462 (N_7462,N_4254,N_4469);
xor U7463 (N_7463,N_4247,N_4480);
and U7464 (N_7464,N_5394,N_4631);
or U7465 (N_7465,N_4919,N_3537);
or U7466 (N_7466,N_5793,N_5341);
xnor U7467 (N_7467,N_5920,N_3415);
or U7468 (N_7468,N_4179,N_3876);
nand U7469 (N_7469,N_4675,N_3892);
or U7470 (N_7470,N_4561,N_4340);
and U7471 (N_7471,N_5722,N_3960);
nor U7472 (N_7472,N_5935,N_5179);
nand U7473 (N_7473,N_3374,N_3942);
nand U7474 (N_7474,N_4726,N_4786);
nor U7475 (N_7475,N_3235,N_3971);
nand U7476 (N_7476,N_5969,N_4196);
or U7477 (N_7477,N_4241,N_5558);
nor U7478 (N_7478,N_3361,N_4053);
or U7479 (N_7479,N_3512,N_4176);
nor U7480 (N_7480,N_4792,N_4470);
and U7481 (N_7481,N_4502,N_4817);
xnor U7482 (N_7482,N_4693,N_5221);
and U7483 (N_7483,N_5652,N_4103);
nand U7484 (N_7484,N_3598,N_5976);
or U7485 (N_7485,N_5866,N_5816);
nor U7486 (N_7486,N_3850,N_3913);
nor U7487 (N_7487,N_5474,N_4776);
xnor U7488 (N_7488,N_3310,N_3198);
nand U7489 (N_7489,N_3808,N_3917);
nor U7490 (N_7490,N_4903,N_3370);
nand U7491 (N_7491,N_5349,N_4429);
or U7492 (N_7492,N_3242,N_3413);
and U7493 (N_7493,N_3810,N_4646);
nand U7494 (N_7494,N_5699,N_3549);
or U7495 (N_7495,N_3141,N_5678);
nor U7496 (N_7496,N_3405,N_5914);
or U7497 (N_7497,N_4649,N_5830);
or U7498 (N_7498,N_5077,N_5491);
xnor U7499 (N_7499,N_3737,N_5596);
xor U7500 (N_7500,N_4643,N_5203);
nor U7501 (N_7501,N_5390,N_4538);
xor U7502 (N_7502,N_3817,N_4830);
nor U7503 (N_7503,N_5970,N_3233);
nor U7504 (N_7504,N_3965,N_4884);
and U7505 (N_7505,N_5037,N_3495);
nand U7506 (N_7506,N_5126,N_5619);
nor U7507 (N_7507,N_3302,N_5879);
xor U7508 (N_7508,N_4799,N_5319);
nor U7509 (N_7509,N_3263,N_3269);
nor U7510 (N_7510,N_4345,N_3798);
or U7511 (N_7511,N_3296,N_4140);
and U7512 (N_7512,N_5154,N_5389);
and U7513 (N_7513,N_3856,N_4656);
xor U7514 (N_7514,N_4605,N_3022);
nor U7515 (N_7515,N_4912,N_4631);
xor U7516 (N_7516,N_4679,N_4311);
nor U7517 (N_7517,N_5576,N_3757);
xnor U7518 (N_7518,N_3997,N_5802);
xor U7519 (N_7519,N_5793,N_3861);
nand U7520 (N_7520,N_5501,N_5007);
and U7521 (N_7521,N_5972,N_4002);
nor U7522 (N_7522,N_3339,N_5534);
nand U7523 (N_7523,N_5197,N_5250);
and U7524 (N_7524,N_3555,N_4727);
and U7525 (N_7525,N_4410,N_4871);
or U7526 (N_7526,N_3445,N_4285);
or U7527 (N_7527,N_5486,N_4536);
nor U7528 (N_7528,N_5822,N_5338);
and U7529 (N_7529,N_5153,N_5804);
nor U7530 (N_7530,N_5891,N_4714);
and U7531 (N_7531,N_3663,N_5822);
and U7532 (N_7532,N_4863,N_5741);
nand U7533 (N_7533,N_5330,N_3967);
and U7534 (N_7534,N_5369,N_5727);
or U7535 (N_7535,N_4924,N_4416);
nand U7536 (N_7536,N_5168,N_3951);
and U7537 (N_7537,N_4890,N_5465);
and U7538 (N_7538,N_5176,N_5214);
xnor U7539 (N_7539,N_3041,N_4389);
nor U7540 (N_7540,N_3094,N_4041);
nand U7541 (N_7541,N_4396,N_4787);
nor U7542 (N_7542,N_3981,N_4950);
and U7543 (N_7543,N_3009,N_3206);
nor U7544 (N_7544,N_5685,N_5487);
and U7545 (N_7545,N_5948,N_4555);
nand U7546 (N_7546,N_4951,N_4245);
nor U7547 (N_7547,N_5273,N_3975);
nor U7548 (N_7548,N_5063,N_5754);
nor U7549 (N_7549,N_3908,N_3083);
nor U7550 (N_7550,N_5770,N_3275);
or U7551 (N_7551,N_5116,N_3648);
nor U7552 (N_7552,N_5705,N_4283);
nand U7553 (N_7553,N_4670,N_4232);
nor U7554 (N_7554,N_4598,N_5045);
nor U7555 (N_7555,N_4039,N_5394);
and U7556 (N_7556,N_5842,N_5986);
nand U7557 (N_7557,N_5521,N_5522);
or U7558 (N_7558,N_4106,N_4717);
and U7559 (N_7559,N_4236,N_4554);
and U7560 (N_7560,N_4849,N_4339);
and U7561 (N_7561,N_4975,N_4665);
and U7562 (N_7562,N_3047,N_4065);
nand U7563 (N_7563,N_4430,N_4193);
xor U7564 (N_7564,N_3830,N_3416);
and U7565 (N_7565,N_3597,N_4614);
or U7566 (N_7566,N_3098,N_3233);
nand U7567 (N_7567,N_3468,N_3864);
nand U7568 (N_7568,N_3661,N_5303);
and U7569 (N_7569,N_3819,N_4092);
xnor U7570 (N_7570,N_3787,N_3698);
xnor U7571 (N_7571,N_4636,N_5366);
and U7572 (N_7572,N_3786,N_5729);
or U7573 (N_7573,N_3249,N_3697);
nand U7574 (N_7574,N_5270,N_5972);
and U7575 (N_7575,N_3879,N_3598);
or U7576 (N_7576,N_4250,N_4691);
xor U7577 (N_7577,N_3008,N_5094);
nor U7578 (N_7578,N_4626,N_4420);
xnor U7579 (N_7579,N_3457,N_4072);
or U7580 (N_7580,N_5623,N_5032);
nand U7581 (N_7581,N_4544,N_5757);
and U7582 (N_7582,N_4177,N_3048);
or U7583 (N_7583,N_5585,N_3549);
or U7584 (N_7584,N_3790,N_3160);
and U7585 (N_7585,N_3128,N_5873);
or U7586 (N_7586,N_5303,N_3051);
and U7587 (N_7587,N_3492,N_5645);
or U7588 (N_7588,N_4450,N_4177);
nor U7589 (N_7589,N_5906,N_3698);
xor U7590 (N_7590,N_4713,N_5796);
and U7591 (N_7591,N_4647,N_4578);
nand U7592 (N_7592,N_4180,N_3230);
xor U7593 (N_7593,N_5094,N_4429);
and U7594 (N_7594,N_4724,N_3972);
nand U7595 (N_7595,N_5860,N_3340);
or U7596 (N_7596,N_3363,N_3939);
or U7597 (N_7597,N_4168,N_5282);
nor U7598 (N_7598,N_3127,N_4748);
xor U7599 (N_7599,N_3283,N_5229);
and U7600 (N_7600,N_4703,N_3816);
nor U7601 (N_7601,N_3685,N_3991);
nand U7602 (N_7602,N_4276,N_3034);
nor U7603 (N_7603,N_4822,N_5674);
nand U7604 (N_7604,N_4000,N_5293);
and U7605 (N_7605,N_5787,N_4945);
and U7606 (N_7606,N_5640,N_4357);
or U7607 (N_7607,N_5627,N_5618);
nor U7608 (N_7608,N_4879,N_5379);
or U7609 (N_7609,N_5583,N_5930);
or U7610 (N_7610,N_5034,N_3416);
nand U7611 (N_7611,N_5426,N_3010);
xor U7612 (N_7612,N_5618,N_4802);
nand U7613 (N_7613,N_5199,N_3120);
and U7614 (N_7614,N_3107,N_5396);
xnor U7615 (N_7615,N_4649,N_4114);
and U7616 (N_7616,N_4416,N_3197);
xnor U7617 (N_7617,N_3792,N_3783);
nand U7618 (N_7618,N_3665,N_3112);
nor U7619 (N_7619,N_4508,N_3806);
and U7620 (N_7620,N_5870,N_3195);
or U7621 (N_7621,N_4531,N_5227);
nand U7622 (N_7622,N_5224,N_5740);
or U7623 (N_7623,N_3859,N_3131);
xor U7624 (N_7624,N_4772,N_4204);
xnor U7625 (N_7625,N_4834,N_4987);
nor U7626 (N_7626,N_4557,N_4910);
nor U7627 (N_7627,N_5336,N_4367);
xnor U7628 (N_7628,N_4783,N_3032);
and U7629 (N_7629,N_4851,N_5441);
nor U7630 (N_7630,N_4514,N_4334);
nand U7631 (N_7631,N_3902,N_3314);
and U7632 (N_7632,N_5154,N_3460);
and U7633 (N_7633,N_3304,N_5506);
and U7634 (N_7634,N_4418,N_4211);
or U7635 (N_7635,N_4376,N_4756);
nand U7636 (N_7636,N_4489,N_4940);
nand U7637 (N_7637,N_4767,N_4265);
xor U7638 (N_7638,N_4378,N_5756);
and U7639 (N_7639,N_4097,N_3858);
xnor U7640 (N_7640,N_3833,N_3275);
nand U7641 (N_7641,N_3392,N_3275);
xor U7642 (N_7642,N_4289,N_3210);
nor U7643 (N_7643,N_5702,N_4435);
nor U7644 (N_7644,N_3174,N_5981);
nand U7645 (N_7645,N_3686,N_3141);
xor U7646 (N_7646,N_3089,N_3917);
or U7647 (N_7647,N_3192,N_4617);
nor U7648 (N_7648,N_5828,N_3284);
or U7649 (N_7649,N_5474,N_5350);
nor U7650 (N_7650,N_3426,N_4530);
or U7651 (N_7651,N_5043,N_4087);
xnor U7652 (N_7652,N_3782,N_5326);
and U7653 (N_7653,N_3074,N_4892);
and U7654 (N_7654,N_4047,N_4177);
nand U7655 (N_7655,N_5222,N_4091);
or U7656 (N_7656,N_3622,N_3494);
and U7657 (N_7657,N_3505,N_4695);
or U7658 (N_7658,N_3698,N_4335);
xor U7659 (N_7659,N_5776,N_5103);
and U7660 (N_7660,N_3513,N_4894);
and U7661 (N_7661,N_4628,N_4153);
and U7662 (N_7662,N_5839,N_3197);
xnor U7663 (N_7663,N_4472,N_5164);
nor U7664 (N_7664,N_4934,N_5142);
xor U7665 (N_7665,N_5158,N_3716);
and U7666 (N_7666,N_3079,N_4917);
and U7667 (N_7667,N_3475,N_5436);
or U7668 (N_7668,N_5168,N_3642);
or U7669 (N_7669,N_3783,N_4610);
nand U7670 (N_7670,N_5938,N_5128);
nor U7671 (N_7671,N_4784,N_4991);
and U7672 (N_7672,N_3144,N_3732);
and U7673 (N_7673,N_5548,N_3396);
nand U7674 (N_7674,N_5949,N_4618);
nand U7675 (N_7675,N_5229,N_3144);
nand U7676 (N_7676,N_3950,N_4123);
and U7677 (N_7677,N_5634,N_4741);
and U7678 (N_7678,N_4655,N_3689);
nand U7679 (N_7679,N_3021,N_3486);
xnor U7680 (N_7680,N_4062,N_3233);
nor U7681 (N_7681,N_5799,N_3328);
nor U7682 (N_7682,N_3797,N_3141);
nor U7683 (N_7683,N_4886,N_3455);
nor U7684 (N_7684,N_5895,N_4387);
or U7685 (N_7685,N_5843,N_3883);
nor U7686 (N_7686,N_4372,N_4254);
and U7687 (N_7687,N_5930,N_4890);
nand U7688 (N_7688,N_3691,N_5730);
or U7689 (N_7689,N_3379,N_4225);
and U7690 (N_7690,N_3684,N_4854);
and U7691 (N_7691,N_3090,N_4491);
nor U7692 (N_7692,N_4518,N_3449);
and U7693 (N_7693,N_5747,N_4780);
xnor U7694 (N_7694,N_5268,N_4827);
xor U7695 (N_7695,N_5055,N_4780);
nor U7696 (N_7696,N_3237,N_3591);
xnor U7697 (N_7697,N_5887,N_4683);
and U7698 (N_7698,N_5054,N_5248);
or U7699 (N_7699,N_3648,N_4143);
nand U7700 (N_7700,N_3888,N_5931);
nand U7701 (N_7701,N_3732,N_5523);
nor U7702 (N_7702,N_3487,N_3112);
nand U7703 (N_7703,N_4683,N_4483);
and U7704 (N_7704,N_5978,N_5574);
nand U7705 (N_7705,N_4693,N_4105);
or U7706 (N_7706,N_3492,N_4488);
xor U7707 (N_7707,N_4970,N_5221);
nor U7708 (N_7708,N_3316,N_3597);
xor U7709 (N_7709,N_4072,N_5673);
or U7710 (N_7710,N_3067,N_5155);
and U7711 (N_7711,N_3440,N_4175);
or U7712 (N_7712,N_3847,N_3977);
nand U7713 (N_7713,N_4237,N_5257);
nor U7714 (N_7714,N_3739,N_4901);
and U7715 (N_7715,N_4128,N_5081);
nand U7716 (N_7716,N_5436,N_5259);
and U7717 (N_7717,N_4955,N_3324);
nand U7718 (N_7718,N_5881,N_3983);
and U7719 (N_7719,N_4798,N_4455);
nand U7720 (N_7720,N_3350,N_4239);
nand U7721 (N_7721,N_4416,N_4425);
or U7722 (N_7722,N_3115,N_4935);
or U7723 (N_7723,N_4290,N_4235);
nand U7724 (N_7724,N_5577,N_4130);
nand U7725 (N_7725,N_3322,N_3002);
nand U7726 (N_7726,N_5210,N_4355);
nor U7727 (N_7727,N_4422,N_3058);
nor U7728 (N_7728,N_5583,N_5924);
nand U7729 (N_7729,N_5805,N_3535);
and U7730 (N_7730,N_3960,N_3142);
xnor U7731 (N_7731,N_5250,N_3754);
xor U7732 (N_7732,N_3402,N_5351);
or U7733 (N_7733,N_4742,N_5689);
nor U7734 (N_7734,N_5058,N_4466);
xor U7735 (N_7735,N_3577,N_3040);
nand U7736 (N_7736,N_3768,N_4593);
nand U7737 (N_7737,N_3840,N_5020);
nor U7738 (N_7738,N_3403,N_4474);
or U7739 (N_7739,N_5708,N_4220);
nor U7740 (N_7740,N_3029,N_4102);
nor U7741 (N_7741,N_3087,N_4568);
or U7742 (N_7742,N_5070,N_3086);
or U7743 (N_7743,N_4698,N_3014);
nor U7744 (N_7744,N_3032,N_3851);
xnor U7745 (N_7745,N_5483,N_3095);
or U7746 (N_7746,N_3275,N_3055);
nor U7747 (N_7747,N_5438,N_4707);
nor U7748 (N_7748,N_4759,N_5660);
nand U7749 (N_7749,N_3034,N_4321);
nor U7750 (N_7750,N_5984,N_3864);
nand U7751 (N_7751,N_3674,N_3850);
xor U7752 (N_7752,N_3187,N_3084);
or U7753 (N_7753,N_3505,N_5869);
xor U7754 (N_7754,N_4402,N_3834);
and U7755 (N_7755,N_3683,N_4634);
nor U7756 (N_7756,N_3102,N_3263);
or U7757 (N_7757,N_4708,N_4076);
and U7758 (N_7758,N_3102,N_4805);
xnor U7759 (N_7759,N_5768,N_4461);
xnor U7760 (N_7760,N_5018,N_3530);
xor U7761 (N_7761,N_3359,N_3225);
or U7762 (N_7762,N_3908,N_4036);
and U7763 (N_7763,N_4155,N_3688);
nor U7764 (N_7764,N_5006,N_4084);
nor U7765 (N_7765,N_5920,N_4438);
or U7766 (N_7766,N_5743,N_5980);
nor U7767 (N_7767,N_4129,N_3283);
or U7768 (N_7768,N_4431,N_4318);
and U7769 (N_7769,N_4668,N_5774);
or U7770 (N_7770,N_4207,N_5932);
and U7771 (N_7771,N_5372,N_4088);
and U7772 (N_7772,N_4948,N_3458);
nor U7773 (N_7773,N_4031,N_5845);
or U7774 (N_7774,N_3894,N_4208);
nand U7775 (N_7775,N_3244,N_3728);
nand U7776 (N_7776,N_5713,N_5063);
nand U7777 (N_7777,N_5065,N_4725);
nand U7778 (N_7778,N_3339,N_3745);
nand U7779 (N_7779,N_5105,N_4848);
xor U7780 (N_7780,N_5465,N_5243);
and U7781 (N_7781,N_4210,N_5910);
nor U7782 (N_7782,N_4296,N_4704);
or U7783 (N_7783,N_5276,N_5712);
nand U7784 (N_7784,N_5553,N_4268);
xor U7785 (N_7785,N_3245,N_4063);
nand U7786 (N_7786,N_5808,N_4945);
nor U7787 (N_7787,N_5534,N_4133);
or U7788 (N_7788,N_3008,N_5630);
or U7789 (N_7789,N_4181,N_3455);
xnor U7790 (N_7790,N_3719,N_5564);
xor U7791 (N_7791,N_5356,N_3381);
nand U7792 (N_7792,N_5934,N_5902);
xnor U7793 (N_7793,N_5061,N_5277);
and U7794 (N_7794,N_3442,N_5886);
or U7795 (N_7795,N_3101,N_5105);
nand U7796 (N_7796,N_3362,N_3347);
xnor U7797 (N_7797,N_5933,N_3931);
and U7798 (N_7798,N_4789,N_3363);
xor U7799 (N_7799,N_3312,N_5659);
nand U7800 (N_7800,N_3870,N_4622);
xnor U7801 (N_7801,N_3612,N_3424);
or U7802 (N_7802,N_5913,N_4335);
nor U7803 (N_7803,N_4996,N_3495);
nor U7804 (N_7804,N_5468,N_5119);
and U7805 (N_7805,N_5937,N_4635);
and U7806 (N_7806,N_3548,N_4153);
and U7807 (N_7807,N_4971,N_3860);
xnor U7808 (N_7808,N_4461,N_4675);
nand U7809 (N_7809,N_4963,N_5226);
and U7810 (N_7810,N_5037,N_4388);
nand U7811 (N_7811,N_5961,N_5919);
xnor U7812 (N_7812,N_4843,N_4543);
xor U7813 (N_7813,N_4959,N_5622);
nor U7814 (N_7814,N_5180,N_3633);
xor U7815 (N_7815,N_4838,N_3616);
or U7816 (N_7816,N_5593,N_3178);
and U7817 (N_7817,N_4946,N_5996);
and U7818 (N_7818,N_5177,N_4792);
or U7819 (N_7819,N_3002,N_5989);
nor U7820 (N_7820,N_3188,N_5990);
and U7821 (N_7821,N_5753,N_3288);
and U7822 (N_7822,N_3143,N_5434);
xor U7823 (N_7823,N_4599,N_5091);
or U7824 (N_7824,N_5348,N_3161);
nand U7825 (N_7825,N_5628,N_3626);
or U7826 (N_7826,N_5450,N_4161);
nand U7827 (N_7827,N_4048,N_5869);
xor U7828 (N_7828,N_4526,N_3355);
or U7829 (N_7829,N_4147,N_5735);
xnor U7830 (N_7830,N_3674,N_5992);
nor U7831 (N_7831,N_5382,N_4569);
nand U7832 (N_7832,N_4215,N_3747);
xor U7833 (N_7833,N_3752,N_5741);
nor U7834 (N_7834,N_4476,N_4498);
nor U7835 (N_7835,N_4347,N_3697);
xnor U7836 (N_7836,N_3741,N_3773);
or U7837 (N_7837,N_3946,N_5237);
or U7838 (N_7838,N_4673,N_3903);
xor U7839 (N_7839,N_4539,N_3733);
and U7840 (N_7840,N_3461,N_5276);
and U7841 (N_7841,N_3214,N_5715);
xnor U7842 (N_7842,N_4556,N_4151);
nor U7843 (N_7843,N_5243,N_4745);
xor U7844 (N_7844,N_3026,N_4568);
and U7845 (N_7845,N_5282,N_5611);
nand U7846 (N_7846,N_3428,N_3766);
nor U7847 (N_7847,N_3359,N_4771);
and U7848 (N_7848,N_4238,N_4717);
and U7849 (N_7849,N_4788,N_4078);
nor U7850 (N_7850,N_3119,N_4992);
nand U7851 (N_7851,N_3041,N_5030);
nor U7852 (N_7852,N_3971,N_4642);
or U7853 (N_7853,N_5838,N_3969);
or U7854 (N_7854,N_5758,N_3938);
nor U7855 (N_7855,N_4952,N_4454);
nand U7856 (N_7856,N_5652,N_5301);
and U7857 (N_7857,N_4089,N_4630);
and U7858 (N_7858,N_3428,N_3389);
and U7859 (N_7859,N_5721,N_3162);
and U7860 (N_7860,N_5467,N_4031);
and U7861 (N_7861,N_5469,N_5264);
nand U7862 (N_7862,N_3254,N_4100);
and U7863 (N_7863,N_3415,N_4698);
nor U7864 (N_7864,N_5516,N_4073);
xnor U7865 (N_7865,N_5082,N_3042);
or U7866 (N_7866,N_4474,N_3971);
or U7867 (N_7867,N_5385,N_5612);
nor U7868 (N_7868,N_4753,N_4235);
nand U7869 (N_7869,N_4508,N_5942);
or U7870 (N_7870,N_3255,N_4469);
nand U7871 (N_7871,N_5554,N_4618);
or U7872 (N_7872,N_4474,N_3141);
and U7873 (N_7873,N_4094,N_5004);
nand U7874 (N_7874,N_3210,N_4484);
or U7875 (N_7875,N_4178,N_4115);
and U7876 (N_7876,N_5272,N_4472);
or U7877 (N_7877,N_5347,N_4566);
nand U7878 (N_7878,N_3478,N_4317);
and U7879 (N_7879,N_5438,N_3621);
xor U7880 (N_7880,N_3062,N_5244);
nor U7881 (N_7881,N_5770,N_5969);
and U7882 (N_7882,N_3952,N_3745);
or U7883 (N_7883,N_3011,N_5195);
xor U7884 (N_7884,N_5343,N_5633);
or U7885 (N_7885,N_5829,N_4310);
xnor U7886 (N_7886,N_5886,N_5497);
xnor U7887 (N_7887,N_4583,N_4465);
or U7888 (N_7888,N_3431,N_4227);
xnor U7889 (N_7889,N_4876,N_4760);
xnor U7890 (N_7890,N_3708,N_3840);
and U7891 (N_7891,N_3049,N_3334);
nor U7892 (N_7892,N_3531,N_4281);
xnor U7893 (N_7893,N_3902,N_4151);
nand U7894 (N_7894,N_3192,N_5673);
nor U7895 (N_7895,N_5302,N_4390);
nand U7896 (N_7896,N_5892,N_3872);
nand U7897 (N_7897,N_3163,N_4520);
or U7898 (N_7898,N_4888,N_3951);
nand U7899 (N_7899,N_3594,N_5371);
or U7900 (N_7900,N_5668,N_4202);
or U7901 (N_7901,N_3558,N_4612);
nor U7902 (N_7902,N_5968,N_3952);
nor U7903 (N_7903,N_4602,N_5353);
or U7904 (N_7904,N_4790,N_3491);
nor U7905 (N_7905,N_5892,N_4165);
or U7906 (N_7906,N_4491,N_5071);
xnor U7907 (N_7907,N_5300,N_5680);
or U7908 (N_7908,N_3587,N_3166);
or U7909 (N_7909,N_5929,N_3544);
nand U7910 (N_7910,N_5830,N_3522);
and U7911 (N_7911,N_5511,N_5931);
or U7912 (N_7912,N_5331,N_3881);
and U7913 (N_7913,N_5023,N_3368);
nor U7914 (N_7914,N_4801,N_3919);
and U7915 (N_7915,N_4755,N_5830);
and U7916 (N_7916,N_3581,N_5138);
nor U7917 (N_7917,N_5265,N_3714);
nor U7918 (N_7918,N_5914,N_3254);
and U7919 (N_7919,N_5601,N_5003);
nor U7920 (N_7920,N_3478,N_4782);
xnor U7921 (N_7921,N_4745,N_3951);
or U7922 (N_7922,N_4086,N_4879);
and U7923 (N_7923,N_4175,N_3372);
and U7924 (N_7924,N_3074,N_5263);
nor U7925 (N_7925,N_4400,N_5385);
nor U7926 (N_7926,N_5788,N_5306);
or U7927 (N_7927,N_4335,N_5300);
nand U7928 (N_7928,N_3630,N_5584);
or U7929 (N_7929,N_5241,N_4168);
or U7930 (N_7930,N_5437,N_5594);
and U7931 (N_7931,N_5240,N_3097);
nor U7932 (N_7932,N_5413,N_3513);
nor U7933 (N_7933,N_4332,N_3869);
xnor U7934 (N_7934,N_4749,N_5022);
nand U7935 (N_7935,N_4224,N_5637);
xnor U7936 (N_7936,N_5033,N_5944);
nand U7937 (N_7937,N_4634,N_5749);
nor U7938 (N_7938,N_4956,N_5843);
xnor U7939 (N_7939,N_5108,N_4417);
nor U7940 (N_7940,N_3671,N_4676);
nor U7941 (N_7941,N_3294,N_5209);
xnor U7942 (N_7942,N_4778,N_3489);
xor U7943 (N_7943,N_5363,N_3403);
or U7944 (N_7944,N_3855,N_3306);
or U7945 (N_7945,N_5085,N_3974);
and U7946 (N_7946,N_4753,N_4023);
nor U7947 (N_7947,N_5343,N_5541);
xnor U7948 (N_7948,N_5454,N_5207);
nand U7949 (N_7949,N_5886,N_4600);
nand U7950 (N_7950,N_5279,N_4775);
or U7951 (N_7951,N_3542,N_4345);
nor U7952 (N_7952,N_4738,N_4265);
or U7953 (N_7953,N_4967,N_5598);
or U7954 (N_7954,N_4066,N_3972);
nor U7955 (N_7955,N_4372,N_5701);
nor U7956 (N_7956,N_4026,N_3826);
xnor U7957 (N_7957,N_4040,N_5598);
nand U7958 (N_7958,N_5970,N_4576);
or U7959 (N_7959,N_5209,N_4956);
nor U7960 (N_7960,N_3788,N_5542);
nand U7961 (N_7961,N_5925,N_5398);
xnor U7962 (N_7962,N_4323,N_3514);
or U7963 (N_7963,N_5652,N_5727);
nand U7964 (N_7964,N_5482,N_4925);
and U7965 (N_7965,N_4997,N_5535);
nor U7966 (N_7966,N_4614,N_4097);
or U7967 (N_7967,N_5172,N_4070);
or U7968 (N_7968,N_3785,N_4053);
nor U7969 (N_7969,N_5115,N_5690);
and U7970 (N_7970,N_3612,N_5095);
nand U7971 (N_7971,N_4779,N_4227);
nor U7972 (N_7972,N_4735,N_5509);
and U7973 (N_7973,N_4914,N_5045);
xor U7974 (N_7974,N_3042,N_5546);
nand U7975 (N_7975,N_4978,N_4364);
and U7976 (N_7976,N_4004,N_4513);
nand U7977 (N_7977,N_4324,N_3671);
nor U7978 (N_7978,N_4526,N_3066);
nor U7979 (N_7979,N_4658,N_4031);
xor U7980 (N_7980,N_4422,N_5713);
nor U7981 (N_7981,N_4819,N_3616);
xnor U7982 (N_7982,N_5470,N_5300);
or U7983 (N_7983,N_3483,N_5963);
or U7984 (N_7984,N_3038,N_4728);
or U7985 (N_7985,N_5151,N_3507);
nor U7986 (N_7986,N_3169,N_5895);
nand U7987 (N_7987,N_3572,N_4432);
nand U7988 (N_7988,N_4608,N_5792);
nor U7989 (N_7989,N_4225,N_3748);
xor U7990 (N_7990,N_4155,N_3164);
and U7991 (N_7991,N_4133,N_3489);
nand U7992 (N_7992,N_4097,N_4649);
and U7993 (N_7993,N_5797,N_5212);
or U7994 (N_7994,N_5767,N_3916);
and U7995 (N_7995,N_4869,N_5201);
nor U7996 (N_7996,N_4755,N_5709);
and U7997 (N_7997,N_4900,N_5125);
xor U7998 (N_7998,N_3845,N_4703);
nor U7999 (N_7999,N_3464,N_4537);
xnor U8000 (N_8000,N_3247,N_4514);
or U8001 (N_8001,N_3166,N_5911);
or U8002 (N_8002,N_3148,N_5224);
nand U8003 (N_8003,N_3722,N_5050);
xnor U8004 (N_8004,N_4301,N_3428);
or U8005 (N_8005,N_3986,N_4798);
nand U8006 (N_8006,N_3046,N_4184);
nor U8007 (N_8007,N_3208,N_3091);
xnor U8008 (N_8008,N_5300,N_5711);
nand U8009 (N_8009,N_3314,N_5647);
and U8010 (N_8010,N_3179,N_5968);
and U8011 (N_8011,N_3084,N_5443);
and U8012 (N_8012,N_5382,N_4078);
nand U8013 (N_8013,N_5812,N_4105);
and U8014 (N_8014,N_5709,N_5427);
nand U8015 (N_8015,N_4872,N_3574);
or U8016 (N_8016,N_4130,N_5144);
xor U8017 (N_8017,N_4356,N_4999);
nand U8018 (N_8018,N_3902,N_3482);
xor U8019 (N_8019,N_5585,N_3793);
nand U8020 (N_8020,N_3317,N_4961);
xnor U8021 (N_8021,N_5654,N_4686);
nor U8022 (N_8022,N_5466,N_4922);
and U8023 (N_8023,N_4227,N_3978);
nand U8024 (N_8024,N_4629,N_3435);
xnor U8025 (N_8025,N_5494,N_3996);
nand U8026 (N_8026,N_3619,N_4473);
and U8027 (N_8027,N_5533,N_5862);
nand U8028 (N_8028,N_4457,N_5981);
nor U8029 (N_8029,N_4520,N_5224);
nand U8030 (N_8030,N_4739,N_3180);
nor U8031 (N_8031,N_4085,N_4379);
and U8032 (N_8032,N_5758,N_4180);
and U8033 (N_8033,N_5750,N_3039);
and U8034 (N_8034,N_5734,N_3137);
or U8035 (N_8035,N_5032,N_5730);
nand U8036 (N_8036,N_4664,N_3004);
nor U8037 (N_8037,N_4629,N_5336);
and U8038 (N_8038,N_3662,N_5606);
or U8039 (N_8039,N_3635,N_5780);
nor U8040 (N_8040,N_4090,N_3448);
or U8041 (N_8041,N_3377,N_4120);
and U8042 (N_8042,N_4990,N_5231);
and U8043 (N_8043,N_3145,N_4514);
nand U8044 (N_8044,N_4203,N_3703);
or U8045 (N_8045,N_3702,N_5761);
nor U8046 (N_8046,N_5794,N_4880);
xor U8047 (N_8047,N_3749,N_4613);
and U8048 (N_8048,N_5669,N_5594);
and U8049 (N_8049,N_4409,N_5120);
and U8050 (N_8050,N_3985,N_5076);
xor U8051 (N_8051,N_4497,N_4684);
xor U8052 (N_8052,N_3339,N_5348);
or U8053 (N_8053,N_3198,N_5164);
nor U8054 (N_8054,N_3765,N_4280);
nand U8055 (N_8055,N_4287,N_4119);
or U8056 (N_8056,N_4989,N_3504);
xor U8057 (N_8057,N_3487,N_4624);
xor U8058 (N_8058,N_4094,N_3583);
nor U8059 (N_8059,N_5026,N_5181);
xnor U8060 (N_8060,N_5453,N_4711);
and U8061 (N_8061,N_4694,N_3282);
nor U8062 (N_8062,N_5007,N_4968);
or U8063 (N_8063,N_5885,N_4188);
nand U8064 (N_8064,N_4227,N_4185);
and U8065 (N_8065,N_3161,N_5602);
and U8066 (N_8066,N_5152,N_3372);
or U8067 (N_8067,N_4785,N_3870);
xnor U8068 (N_8068,N_3099,N_4321);
nor U8069 (N_8069,N_3972,N_3775);
and U8070 (N_8070,N_5659,N_3902);
and U8071 (N_8071,N_4381,N_4776);
xnor U8072 (N_8072,N_3607,N_4487);
xnor U8073 (N_8073,N_4218,N_5616);
or U8074 (N_8074,N_5930,N_5966);
nor U8075 (N_8075,N_4913,N_3467);
xnor U8076 (N_8076,N_3140,N_5223);
nand U8077 (N_8077,N_4631,N_5909);
and U8078 (N_8078,N_3938,N_3449);
and U8079 (N_8079,N_4528,N_4829);
or U8080 (N_8080,N_4474,N_5360);
or U8081 (N_8081,N_5036,N_4579);
nand U8082 (N_8082,N_3133,N_4856);
and U8083 (N_8083,N_3787,N_4982);
nand U8084 (N_8084,N_5815,N_5476);
or U8085 (N_8085,N_3315,N_4957);
and U8086 (N_8086,N_3173,N_5745);
nor U8087 (N_8087,N_4300,N_4480);
and U8088 (N_8088,N_5778,N_5274);
xor U8089 (N_8089,N_3240,N_5095);
xor U8090 (N_8090,N_5467,N_5082);
nand U8091 (N_8091,N_5032,N_4523);
or U8092 (N_8092,N_4741,N_3741);
or U8093 (N_8093,N_3412,N_5805);
and U8094 (N_8094,N_3560,N_4087);
nand U8095 (N_8095,N_3455,N_5002);
nand U8096 (N_8096,N_4058,N_4411);
xnor U8097 (N_8097,N_5168,N_5970);
nor U8098 (N_8098,N_3346,N_5812);
nor U8099 (N_8099,N_5910,N_3802);
and U8100 (N_8100,N_5260,N_3310);
and U8101 (N_8101,N_5359,N_4428);
xnor U8102 (N_8102,N_5193,N_3134);
xnor U8103 (N_8103,N_5184,N_3614);
xor U8104 (N_8104,N_4207,N_5110);
and U8105 (N_8105,N_4488,N_3602);
or U8106 (N_8106,N_3369,N_4163);
and U8107 (N_8107,N_4667,N_5328);
and U8108 (N_8108,N_3861,N_3400);
and U8109 (N_8109,N_5613,N_4607);
nor U8110 (N_8110,N_5977,N_3466);
or U8111 (N_8111,N_4208,N_3343);
nand U8112 (N_8112,N_4256,N_3556);
nor U8113 (N_8113,N_4464,N_4107);
and U8114 (N_8114,N_3242,N_4700);
xnor U8115 (N_8115,N_5852,N_5918);
xnor U8116 (N_8116,N_4422,N_4272);
and U8117 (N_8117,N_3379,N_5675);
xnor U8118 (N_8118,N_4502,N_5472);
xnor U8119 (N_8119,N_4059,N_5417);
xnor U8120 (N_8120,N_3482,N_3959);
nand U8121 (N_8121,N_4847,N_3007);
nor U8122 (N_8122,N_5255,N_4270);
nor U8123 (N_8123,N_3635,N_3325);
nor U8124 (N_8124,N_4174,N_3179);
nand U8125 (N_8125,N_5117,N_4255);
nor U8126 (N_8126,N_3429,N_5134);
or U8127 (N_8127,N_5227,N_3234);
xor U8128 (N_8128,N_5942,N_3794);
nor U8129 (N_8129,N_5585,N_5162);
and U8130 (N_8130,N_3318,N_3884);
xor U8131 (N_8131,N_5083,N_4438);
xor U8132 (N_8132,N_4032,N_3947);
nor U8133 (N_8133,N_4290,N_3332);
nand U8134 (N_8134,N_5836,N_5528);
and U8135 (N_8135,N_3993,N_4948);
or U8136 (N_8136,N_5647,N_4784);
or U8137 (N_8137,N_3417,N_3138);
or U8138 (N_8138,N_5466,N_3650);
xnor U8139 (N_8139,N_4781,N_5795);
nor U8140 (N_8140,N_4452,N_3929);
nand U8141 (N_8141,N_5835,N_5895);
and U8142 (N_8142,N_3039,N_5982);
and U8143 (N_8143,N_3874,N_4381);
or U8144 (N_8144,N_4984,N_4306);
or U8145 (N_8145,N_4739,N_5522);
and U8146 (N_8146,N_4804,N_3160);
xnor U8147 (N_8147,N_4698,N_3478);
or U8148 (N_8148,N_5564,N_3029);
and U8149 (N_8149,N_4886,N_4127);
or U8150 (N_8150,N_4746,N_5370);
or U8151 (N_8151,N_4406,N_3846);
nand U8152 (N_8152,N_3795,N_3620);
or U8153 (N_8153,N_4857,N_4671);
or U8154 (N_8154,N_4758,N_3069);
or U8155 (N_8155,N_3740,N_5376);
and U8156 (N_8156,N_5668,N_4868);
nor U8157 (N_8157,N_4208,N_3851);
and U8158 (N_8158,N_4755,N_4076);
nand U8159 (N_8159,N_3507,N_4211);
xnor U8160 (N_8160,N_4903,N_5539);
nor U8161 (N_8161,N_5150,N_3783);
xnor U8162 (N_8162,N_3315,N_5803);
nand U8163 (N_8163,N_4974,N_5386);
nor U8164 (N_8164,N_4830,N_4568);
and U8165 (N_8165,N_3621,N_5627);
nand U8166 (N_8166,N_4155,N_3510);
nand U8167 (N_8167,N_3656,N_4648);
and U8168 (N_8168,N_3301,N_4837);
or U8169 (N_8169,N_5780,N_3519);
and U8170 (N_8170,N_3596,N_5019);
or U8171 (N_8171,N_3966,N_5730);
xor U8172 (N_8172,N_5633,N_4916);
and U8173 (N_8173,N_3766,N_3372);
xor U8174 (N_8174,N_4815,N_4373);
xnor U8175 (N_8175,N_4771,N_5979);
nand U8176 (N_8176,N_4000,N_5720);
or U8177 (N_8177,N_5329,N_4270);
and U8178 (N_8178,N_4810,N_5859);
nor U8179 (N_8179,N_3934,N_4659);
nand U8180 (N_8180,N_5046,N_3688);
xnor U8181 (N_8181,N_4341,N_5128);
or U8182 (N_8182,N_3085,N_3924);
nor U8183 (N_8183,N_4841,N_5916);
nand U8184 (N_8184,N_3962,N_3492);
nand U8185 (N_8185,N_4926,N_4856);
nor U8186 (N_8186,N_3074,N_5196);
xor U8187 (N_8187,N_3760,N_3355);
or U8188 (N_8188,N_5223,N_5098);
or U8189 (N_8189,N_3755,N_3469);
xor U8190 (N_8190,N_4388,N_3433);
xnor U8191 (N_8191,N_3386,N_4896);
and U8192 (N_8192,N_4799,N_4280);
nor U8193 (N_8193,N_3424,N_4774);
xnor U8194 (N_8194,N_5431,N_3056);
xnor U8195 (N_8195,N_4526,N_5352);
or U8196 (N_8196,N_4421,N_3586);
nand U8197 (N_8197,N_3280,N_5373);
or U8198 (N_8198,N_3125,N_3101);
or U8199 (N_8199,N_4052,N_3545);
xnor U8200 (N_8200,N_3543,N_3050);
nor U8201 (N_8201,N_3824,N_5325);
nand U8202 (N_8202,N_3468,N_5179);
and U8203 (N_8203,N_5761,N_3007);
nor U8204 (N_8204,N_5625,N_4221);
or U8205 (N_8205,N_5681,N_3244);
nor U8206 (N_8206,N_4204,N_4175);
nand U8207 (N_8207,N_5066,N_3716);
nand U8208 (N_8208,N_5438,N_5149);
nor U8209 (N_8209,N_3531,N_5671);
nor U8210 (N_8210,N_5282,N_4770);
nor U8211 (N_8211,N_3407,N_4472);
or U8212 (N_8212,N_5688,N_3065);
nand U8213 (N_8213,N_3634,N_3242);
and U8214 (N_8214,N_5062,N_5801);
or U8215 (N_8215,N_5908,N_5962);
nor U8216 (N_8216,N_5831,N_3441);
nor U8217 (N_8217,N_3613,N_4266);
or U8218 (N_8218,N_3822,N_4632);
nor U8219 (N_8219,N_5774,N_4929);
xor U8220 (N_8220,N_3338,N_4437);
xnor U8221 (N_8221,N_5858,N_5068);
xnor U8222 (N_8222,N_5051,N_4592);
xor U8223 (N_8223,N_5722,N_5606);
and U8224 (N_8224,N_5748,N_4083);
and U8225 (N_8225,N_3579,N_3647);
xnor U8226 (N_8226,N_5752,N_5513);
xor U8227 (N_8227,N_4205,N_5996);
or U8228 (N_8228,N_3931,N_3854);
or U8229 (N_8229,N_3283,N_3592);
or U8230 (N_8230,N_5615,N_4105);
and U8231 (N_8231,N_3590,N_5250);
or U8232 (N_8232,N_5925,N_4700);
or U8233 (N_8233,N_4912,N_4634);
xnor U8234 (N_8234,N_5693,N_4861);
nand U8235 (N_8235,N_5169,N_3114);
nor U8236 (N_8236,N_3346,N_5413);
or U8237 (N_8237,N_5736,N_5019);
or U8238 (N_8238,N_5329,N_3924);
xor U8239 (N_8239,N_5681,N_4854);
nor U8240 (N_8240,N_4114,N_4176);
nand U8241 (N_8241,N_3972,N_5082);
and U8242 (N_8242,N_4858,N_5549);
or U8243 (N_8243,N_5683,N_5879);
nand U8244 (N_8244,N_4153,N_3363);
and U8245 (N_8245,N_3126,N_3606);
nand U8246 (N_8246,N_4966,N_5746);
or U8247 (N_8247,N_3311,N_4518);
xnor U8248 (N_8248,N_3411,N_4062);
xnor U8249 (N_8249,N_5088,N_5787);
nor U8250 (N_8250,N_5189,N_5950);
and U8251 (N_8251,N_4296,N_5705);
or U8252 (N_8252,N_5093,N_4112);
nor U8253 (N_8253,N_3430,N_5848);
or U8254 (N_8254,N_3239,N_4956);
or U8255 (N_8255,N_5790,N_4004);
xnor U8256 (N_8256,N_4216,N_5885);
and U8257 (N_8257,N_4420,N_5292);
nor U8258 (N_8258,N_5044,N_3133);
nor U8259 (N_8259,N_4269,N_3962);
nor U8260 (N_8260,N_5138,N_4669);
and U8261 (N_8261,N_4516,N_3311);
or U8262 (N_8262,N_5542,N_4079);
nand U8263 (N_8263,N_3773,N_4455);
and U8264 (N_8264,N_4013,N_5219);
or U8265 (N_8265,N_3424,N_4547);
xnor U8266 (N_8266,N_3388,N_3341);
nand U8267 (N_8267,N_5504,N_3047);
and U8268 (N_8268,N_4567,N_4679);
or U8269 (N_8269,N_5918,N_5393);
or U8270 (N_8270,N_5273,N_5013);
or U8271 (N_8271,N_4537,N_4339);
or U8272 (N_8272,N_3066,N_4638);
nor U8273 (N_8273,N_5172,N_3922);
xnor U8274 (N_8274,N_5560,N_3818);
nor U8275 (N_8275,N_4704,N_3577);
nand U8276 (N_8276,N_5811,N_5158);
nand U8277 (N_8277,N_4665,N_3723);
and U8278 (N_8278,N_4492,N_5330);
xor U8279 (N_8279,N_4037,N_4645);
nor U8280 (N_8280,N_3299,N_3474);
or U8281 (N_8281,N_5600,N_3217);
nand U8282 (N_8282,N_3957,N_4654);
xor U8283 (N_8283,N_3241,N_4974);
or U8284 (N_8284,N_3837,N_4957);
nand U8285 (N_8285,N_5919,N_5901);
nand U8286 (N_8286,N_5592,N_3451);
nor U8287 (N_8287,N_5639,N_3316);
nand U8288 (N_8288,N_5832,N_5564);
and U8289 (N_8289,N_4275,N_5100);
nor U8290 (N_8290,N_5271,N_4859);
nor U8291 (N_8291,N_5286,N_4293);
and U8292 (N_8292,N_4919,N_5540);
and U8293 (N_8293,N_3892,N_4318);
and U8294 (N_8294,N_3863,N_4407);
nor U8295 (N_8295,N_5917,N_5385);
xnor U8296 (N_8296,N_4773,N_3568);
xor U8297 (N_8297,N_3510,N_3547);
xor U8298 (N_8298,N_3905,N_5711);
and U8299 (N_8299,N_4131,N_3245);
or U8300 (N_8300,N_5444,N_4434);
xor U8301 (N_8301,N_4344,N_5521);
and U8302 (N_8302,N_4359,N_4261);
xnor U8303 (N_8303,N_4023,N_5234);
or U8304 (N_8304,N_4781,N_5806);
and U8305 (N_8305,N_4278,N_3409);
nand U8306 (N_8306,N_5601,N_4166);
nor U8307 (N_8307,N_4792,N_5661);
xnor U8308 (N_8308,N_4527,N_5338);
nand U8309 (N_8309,N_4746,N_3074);
or U8310 (N_8310,N_5634,N_5073);
nor U8311 (N_8311,N_5867,N_5749);
and U8312 (N_8312,N_3371,N_3117);
or U8313 (N_8313,N_5727,N_5640);
nand U8314 (N_8314,N_5036,N_5300);
or U8315 (N_8315,N_5243,N_4006);
nor U8316 (N_8316,N_5702,N_4688);
nor U8317 (N_8317,N_4523,N_5791);
or U8318 (N_8318,N_4707,N_4513);
nor U8319 (N_8319,N_4510,N_5810);
nor U8320 (N_8320,N_5194,N_4710);
nand U8321 (N_8321,N_3278,N_3197);
xor U8322 (N_8322,N_3220,N_4520);
and U8323 (N_8323,N_3738,N_4083);
xnor U8324 (N_8324,N_5989,N_4677);
nor U8325 (N_8325,N_5116,N_5413);
or U8326 (N_8326,N_5346,N_5628);
xor U8327 (N_8327,N_3971,N_5120);
nand U8328 (N_8328,N_3966,N_3969);
or U8329 (N_8329,N_3730,N_3758);
and U8330 (N_8330,N_3600,N_3769);
xor U8331 (N_8331,N_3043,N_4535);
or U8332 (N_8332,N_3383,N_3941);
nor U8333 (N_8333,N_3480,N_3124);
nand U8334 (N_8334,N_4514,N_3267);
nor U8335 (N_8335,N_5390,N_3614);
nand U8336 (N_8336,N_3736,N_4314);
or U8337 (N_8337,N_3519,N_5540);
or U8338 (N_8338,N_3859,N_3555);
nand U8339 (N_8339,N_3989,N_3880);
nand U8340 (N_8340,N_5368,N_3760);
or U8341 (N_8341,N_4946,N_4597);
and U8342 (N_8342,N_5713,N_4741);
or U8343 (N_8343,N_5708,N_4006);
or U8344 (N_8344,N_5216,N_3880);
nand U8345 (N_8345,N_5329,N_3784);
and U8346 (N_8346,N_4027,N_5910);
nand U8347 (N_8347,N_4171,N_4857);
nor U8348 (N_8348,N_4932,N_5641);
nand U8349 (N_8349,N_3284,N_3603);
xnor U8350 (N_8350,N_4609,N_5332);
nand U8351 (N_8351,N_3960,N_4346);
or U8352 (N_8352,N_4652,N_4095);
or U8353 (N_8353,N_4177,N_4872);
and U8354 (N_8354,N_5149,N_5318);
nand U8355 (N_8355,N_3238,N_4607);
nor U8356 (N_8356,N_5460,N_3531);
or U8357 (N_8357,N_4530,N_5993);
and U8358 (N_8358,N_3439,N_3965);
nand U8359 (N_8359,N_5706,N_4487);
nand U8360 (N_8360,N_4885,N_5368);
or U8361 (N_8361,N_4297,N_4323);
or U8362 (N_8362,N_5577,N_3642);
or U8363 (N_8363,N_4754,N_5510);
and U8364 (N_8364,N_4117,N_3418);
or U8365 (N_8365,N_4231,N_3471);
and U8366 (N_8366,N_4006,N_4485);
nand U8367 (N_8367,N_5547,N_5067);
nand U8368 (N_8368,N_4448,N_5387);
nand U8369 (N_8369,N_4006,N_4182);
or U8370 (N_8370,N_5657,N_3737);
nand U8371 (N_8371,N_3940,N_4690);
nor U8372 (N_8372,N_5733,N_4749);
xnor U8373 (N_8373,N_5954,N_4748);
nand U8374 (N_8374,N_3353,N_5063);
nand U8375 (N_8375,N_5049,N_3762);
and U8376 (N_8376,N_5730,N_5120);
xnor U8377 (N_8377,N_4984,N_5121);
xnor U8378 (N_8378,N_3100,N_3391);
xor U8379 (N_8379,N_5007,N_3875);
and U8380 (N_8380,N_4358,N_5828);
nor U8381 (N_8381,N_4832,N_4666);
and U8382 (N_8382,N_4396,N_5164);
nor U8383 (N_8383,N_4462,N_3314);
nor U8384 (N_8384,N_4501,N_4777);
or U8385 (N_8385,N_4531,N_4097);
or U8386 (N_8386,N_4215,N_5138);
nand U8387 (N_8387,N_5662,N_3805);
nor U8388 (N_8388,N_5359,N_5325);
nand U8389 (N_8389,N_5274,N_3066);
nor U8390 (N_8390,N_5110,N_3957);
or U8391 (N_8391,N_4013,N_3225);
and U8392 (N_8392,N_5468,N_5344);
nand U8393 (N_8393,N_4246,N_4036);
nand U8394 (N_8394,N_5481,N_5373);
nand U8395 (N_8395,N_3057,N_4936);
or U8396 (N_8396,N_5698,N_3883);
nor U8397 (N_8397,N_3257,N_5357);
or U8398 (N_8398,N_4847,N_4247);
xor U8399 (N_8399,N_5182,N_5156);
nand U8400 (N_8400,N_3966,N_5137);
and U8401 (N_8401,N_3578,N_5779);
nand U8402 (N_8402,N_5760,N_3242);
and U8403 (N_8403,N_5073,N_4404);
and U8404 (N_8404,N_5939,N_4297);
xor U8405 (N_8405,N_4897,N_3331);
or U8406 (N_8406,N_5327,N_4054);
xnor U8407 (N_8407,N_5017,N_5945);
nand U8408 (N_8408,N_3298,N_5125);
or U8409 (N_8409,N_4385,N_4684);
and U8410 (N_8410,N_3306,N_3284);
and U8411 (N_8411,N_5550,N_5368);
and U8412 (N_8412,N_3616,N_3903);
nand U8413 (N_8413,N_3278,N_4861);
and U8414 (N_8414,N_4938,N_3116);
xor U8415 (N_8415,N_5149,N_5102);
or U8416 (N_8416,N_3749,N_3117);
xor U8417 (N_8417,N_5419,N_3032);
nor U8418 (N_8418,N_3670,N_5533);
or U8419 (N_8419,N_3492,N_4958);
xor U8420 (N_8420,N_5377,N_4650);
xor U8421 (N_8421,N_3305,N_4208);
nor U8422 (N_8422,N_4324,N_5042);
and U8423 (N_8423,N_4826,N_3269);
nor U8424 (N_8424,N_5835,N_5747);
and U8425 (N_8425,N_5680,N_5020);
or U8426 (N_8426,N_4280,N_4175);
nor U8427 (N_8427,N_4485,N_4625);
nand U8428 (N_8428,N_3418,N_5202);
nor U8429 (N_8429,N_4171,N_5488);
and U8430 (N_8430,N_5953,N_3633);
or U8431 (N_8431,N_5478,N_3435);
and U8432 (N_8432,N_5246,N_5054);
nand U8433 (N_8433,N_4334,N_4748);
nor U8434 (N_8434,N_4495,N_3940);
and U8435 (N_8435,N_3014,N_4495);
or U8436 (N_8436,N_3925,N_5120);
xnor U8437 (N_8437,N_4258,N_5643);
nor U8438 (N_8438,N_5793,N_3190);
nor U8439 (N_8439,N_3319,N_3374);
nor U8440 (N_8440,N_3012,N_4025);
nand U8441 (N_8441,N_5731,N_3906);
or U8442 (N_8442,N_3226,N_3304);
nand U8443 (N_8443,N_4534,N_4751);
or U8444 (N_8444,N_5214,N_5698);
nor U8445 (N_8445,N_4259,N_5511);
or U8446 (N_8446,N_5090,N_4088);
nor U8447 (N_8447,N_5424,N_5015);
xnor U8448 (N_8448,N_5132,N_4352);
nor U8449 (N_8449,N_3665,N_5457);
nor U8450 (N_8450,N_3105,N_4715);
and U8451 (N_8451,N_3660,N_3040);
xor U8452 (N_8452,N_3572,N_4608);
nand U8453 (N_8453,N_5571,N_3551);
or U8454 (N_8454,N_3087,N_3084);
xnor U8455 (N_8455,N_3080,N_4166);
xor U8456 (N_8456,N_4229,N_4445);
xor U8457 (N_8457,N_4604,N_5157);
nor U8458 (N_8458,N_3929,N_4803);
nand U8459 (N_8459,N_5486,N_3262);
nor U8460 (N_8460,N_4004,N_4284);
and U8461 (N_8461,N_3930,N_3434);
or U8462 (N_8462,N_3109,N_3946);
nor U8463 (N_8463,N_5110,N_3179);
and U8464 (N_8464,N_4838,N_5191);
xnor U8465 (N_8465,N_4321,N_4377);
xnor U8466 (N_8466,N_5608,N_4110);
xnor U8467 (N_8467,N_4340,N_4628);
and U8468 (N_8468,N_4594,N_5374);
nand U8469 (N_8469,N_5978,N_4693);
and U8470 (N_8470,N_5405,N_4068);
or U8471 (N_8471,N_4248,N_4347);
xnor U8472 (N_8472,N_5661,N_3100);
or U8473 (N_8473,N_3976,N_3583);
and U8474 (N_8474,N_4384,N_5997);
nor U8475 (N_8475,N_3585,N_5370);
xor U8476 (N_8476,N_4248,N_3729);
and U8477 (N_8477,N_4215,N_4746);
or U8478 (N_8478,N_3216,N_5540);
nor U8479 (N_8479,N_3828,N_3612);
nand U8480 (N_8480,N_3545,N_4607);
nand U8481 (N_8481,N_3043,N_5336);
nand U8482 (N_8482,N_5615,N_3112);
or U8483 (N_8483,N_4911,N_5825);
nor U8484 (N_8484,N_5887,N_4903);
xor U8485 (N_8485,N_3596,N_4619);
nor U8486 (N_8486,N_5696,N_3477);
nor U8487 (N_8487,N_5815,N_5555);
and U8488 (N_8488,N_4958,N_3605);
xor U8489 (N_8489,N_5197,N_5789);
nand U8490 (N_8490,N_4089,N_5337);
nor U8491 (N_8491,N_5689,N_3862);
and U8492 (N_8492,N_4845,N_3195);
nand U8493 (N_8493,N_4903,N_3052);
nor U8494 (N_8494,N_3894,N_3297);
and U8495 (N_8495,N_4346,N_5071);
or U8496 (N_8496,N_3654,N_4040);
and U8497 (N_8497,N_3583,N_3261);
and U8498 (N_8498,N_3393,N_5926);
xnor U8499 (N_8499,N_3504,N_5766);
nand U8500 (N_8500,N_4094,N_4811);
and U8501 (N_8501,N_5579,N_4450);
xor U8502 (N_8502,N_4008,N_4454);
xnor U8503 (N_8503,N_4733,N_4837);
xnor U8504 (N_8504,N_5179,N_3435);
xor U8505 (N_8505,N_4274,N_4596);
xor U8506 (N_8506,N_5514,N_5229);
xnor U8507 (N_8507,N_3040,N_4822);
nor U8508 (N_8508,N_4906,N_4456);
or U8509 (N_8509,N_5791,N_3273);
or U8510 (N_8510,N_3971,N_5255);
or U8511 (N_8511,N_4607,N_5844);
and U8512 (N_8512,N_4746,N_4094);
and U8513 (N_8513,N_4468,N_4192);
nor U8514 (N_8514,N_4508,N_3579);
xor U8515 (N_8515,N_5928,N_3635);
xor U8516 (N_8516,N_4717,N_5046);
nor U8517 (N_8517,N_4521,N_4772);
or U8518 (N_8518,N_3866,N_4937);
xor U8519 (N_8519,N_4283,N_4767);
nor U8520 (N_8520,N_5517,N_3675);
and U8521 (N_8521,N_5811,N_4674);
xor U8522 (N_8522,N_3762,N_5967);
xnor U8523 (N_8523,N_3103,N_4985);
nor U8524 (N_8524,N_3841,N_5082);
nand U8525 (N_8525,N_4703,N_5446);
or U8526 (N_8526,N_5436,N_3325);
xor U8527 (N_8527,N_4949,N_4912);
xnor U8528 (N_8528,N_4707,N_5483);
and U8529 (N_8529,N_5179,N_4868);
or U8530 (N_8530,N_5972,N_5494);
or U8531 (N_8531,N_4621,N_3406);
nand U8532 (N_8532,N_3443,N_5894);
nor U8533 (N_8533,N_5093,N_5696);
or U8534 (N_8534,N_5322,N_5912);
or U8535 (N_8535,N_4885,N_5100);
or U8536 (N_8536,N_4443,N_4277);
or U8537 (N_8537,N_3535,N_3391);
or U8538 (N_8538,N_3864,N_5270);
xor U8539 (N_8539,N_4041,N_4236);
and U8540 (N_8540,N_4510,N_5461);
nor U8541 (N_8541,N_4048,N_5260);
and U8542 (N_8542,N_4616,N_4775);
and U8543 (N_8543,N_3645,N_4687);
nand U8544 (N_8544,N_4997,N_4667);
nand U8545 (N_8545,N_4969,N_5814);
nand U8546 (N_8546,N_4953,N_5667);
or U8547 (N_8547,N_5554,N_4014);
and U8548 (N_8548,N_5442,N_3685);
nand U8549 (N_8549,N_3761,N_5214);
nand U8550 (N_8550,N_3883,N_5527);
nand U8551 (N_8551,N_4462,N_3345);
nand U8552 (N_8552,N_3853,N_4495);
nand U8553 (N_8553,N_4766,N_3484);
or U8554 (N_8554,N_3789,N_3546);
nand U8555 (N_8555,N_5437,N_3039);
nor U8556 (N_8556,N_3063,N_4572);
nor U8557 (N_8557,N_5431,N_3505);
or U8558 (N_8558,N_4283,N_5477);
xor U8559 (N_8559,N_3808,N_3294);
nand U8560 (N_8560,N_4250,N_3360);
nor U8561 (N_8561,N_4833,N_5821);
nand U8562 (N_8562,N_3537,N_3313);
or U8563 (N_8563,N_4516,N_5430);
xnor U8564 (N_8564,N_5983,N_4994);
and U8565 (N_8565,N_4566,N_4250);
or U8566 (N_8566,N_4723,N_4016);
nor U8567 (N_8567,N_4062,N_3183);
and U8568 (N_8568,N_5261,N_4914);
nand U8569 (N_8569,N_4526,N_3630);
nand U8570 (N_8570,N_4652,N_4246);
and U8571 (N_8571,N_5950,N_4954);
nand U8572 (N_8572,N_3872,N_3571);
or U8573 (N_8573,N_5066,N_4882);
or U8574 (N_8574,N_5695,N_3821);
and U8575 (N_8575,N_5519,N_4524);
nand U8576 (N_8576,N_5949,N_3520);
and U8577 (N_8577,N_4487,N_4383);
and U8578 (N_8578,N_4745,N_3493);
nor U8579 (N_8579,N_3105,N_3568);
xor U8580 (N_8580,N_4872,N_3494);
nand U8581 (N_8581,N_3670,N_5490);
nor U8582 (N_8582,N_3620,N_3265);
xor U8583 (N_8583,N_5155,N_3871);
nand U8584 (N_8584,N_5859,N_3750);
or U8585 (N_8585,N_3127,N_3519);
xnor U8586 (N_8586,N_3174,N_4710);
xor U8587 (N_8587,N_4682,N_3835);
nor U8588 (N_8588,N_4169,N_3857);
xor U8589 (N_8589,N_3923,N_4757);
or U8590 (N_8590,N_5301,N_5430);
nor U8591 (N_8591,N_3549,N_4432);
xor U8592 (N_8592,N_3348,N_4673);
nand U8593 (N_8593,N_4883,N_5938);
nand U8594 (N_8594,N_5725,N_4735);
and U8595 (N_8595,N_5662,N_3327);
nand U8596 (N_8596,N_4156,N_3736);
or U8597 (N_8597,N_4759,N_5223);
or U8598 (N_8598,N_4299,N_4476);
xnor U8599 (N_8599,N_3775,N_5961);
nor U8600 (N_8600,N_3187,N_4009);
xor U8601 (N_8601,N_5566,N_4006);
nor U8602 (N_8602,N_5568,N_5242);
xor U8603 (N_8603,N_3334,N_3609);
nand U8604 (N_8604,N_3145,N_3747);
or U8605 (N_8605,N_4355,N_3246);
or U8606 (N_8606,N_5430,N_3148);
nand U8607 (N_8607,N_3106,N_4069);
and U8608 (N_8608,N_3016,N_5470);
or U8609 (N_8609,N_5802,N_3384);
nor U8610 (N_8610,N_4657,N_5779);
or U8611 (N_8611,N_5898,N_3769);
and U8612 (N_8612,N_4109,N_5157);
nor U8613 (N_8613,N_5091,N_5246);
nand U8614 (N_8614,N_5639,N_3611);
and U8615 (N_8615,N_4151,N_3785);
xor U8616 (N_8616,N_4621,N_3492);
and U8617 (N_8617,N_3887,N_3389);
and U8618 (N_8618,N_3316,N_3610);
or U8619 (N_8619,N_4569,N_5402);
or U8620 (N_8620,N_5106,N_4498);
or U8621 (N_8621,N_3037,N_4131);
nand U8622 (N_8622,N_4344,N_5573);
or U8623 (N_8623,N_5710,N_3482);
nand U8624 (N_8624,N_5787,N_3968);
and U8625 (N_8625,N_5117,N_5741);
nor U8626 (N_8626,N_3956,N_4792);
nor U8627 (N_8627,N_4323,N_3109);
and U8628 (N_8628,N_4565,N_4322);
xnor U8629 (N_8629,N_5808,N_3215);
xnor U8630 (N_8630,N_4714,N_5751);
and U8631 (N_8631,N_4143,N_3820);
nor U8632 (N_8632,N_4483,N_3335);
and U8633 (N_8633,N_3880,N_3205);
nor U8634 (N_8634,N_3960,N_3982);
and U8635 (N_8635,N_3037,N_3743);
nand U8636 (N_8636,N_5846,N_5008);
nor U8637 (N_8637,N_3596,N_3242);
nand U8638 (N_8638,N_3042,N_5826);
xnor U8639 (N_8639,N_4590,N_3558);
xnor U8640 (N_8640,N_5750,N_4693);
nand U8641 (N_8641,N_4472,N_5220);
or U8642 (N_8642,N_3397,N_3183);
nor U8643 (N_8643,N_4738,N_4194);
nand U8644 (N_8644,N_4421,N_5145);
and U8645 (N_8645,N_5284,N_3956);
nand U8646 (N_8646,N_4213,N_4084);
or U8647 (N_8647,N_4483,N_4773);
xnor U8648 (N_8648,N_5756,N_4153);
or U8649 (N_8649,N_4748,N_3759);
and U8650 (N_8650,N_5079,N_3056);
or U8651 (N_8651,N_4431,N_4737);
nand U8652 (N_8652,N_4236,N_3394);
or U8653 (N_8653,N_4606,N_5107);
nor U8654 (N_8654,N_4010,N_4463);
xnor U8655 (N_8655,N_5371,N_4191);
and U8656 (N_8656,N_3301,N_3099);
xnor U8657 (N_8657,N_5776,N_5855);
nand U8658 (N_8658,N_4096,N_3266);
or U8659 (N_8659,N_3131,N_3735);
nor U8660 (N_8660,N_3259,N_5189);
nor U8661 (N_8661,N_5598,N_3723);
and U8662 (N_8662,N_5685,N_3393);
xor U8663 (N_8663,N_4033,N_4222);
xor U8664 (N_8664,N_3481,N_4266);
or U8665 (N_8665,N_3178,N_3590);
or U8666 (N_8666,N_3669,N_5247);
or U8667 (N_8667,N_4147,N_5646);
and U8668 (N_8668,N_4407,N_3088);
and U8669 (N_8669,N_3154,N_4516);
and U8670 (N_8670,N_4278,N_5785);
or U8671 (N_8671,N_3388,N_3842);
or U8672 (N_8672,N_4163,N_3636);
xnor U8673 (N_8673,N_4253,N_4014);
and U8674 (N_8674,N_5529,N_5323);
or U8675 (N_8675,N_3217,N_4905);
xor U8676 (N_8676,N_3523,N_5149);
nor U8677 (N_8677,N_5058,N_3888);
or U8678 (N_8678,N_3743,N_5133);
xor U8679 (N_8679,N_5429,N_5951);
and U8680 (N_8680,N_3575,N_3302);
xor U8681 (N_8681,N_5292,N_4991);
nand U8682 (N_8682,N_4964,N_5864);
or U8683 (N_8683,N_5493,N_4213);
or U8684 (N_8684,N_3391,N_5257);
nor U8685 (N_8685,N_5960,N_5310);
nand U8686 (N_8686,N_3129,N_5312);
nor U8687 (N_8687,N_4040,N_4982);
nand U8688 (N_8688,N_3196,N_4689);
or U8689 (N_8689,N_5181,N_5184);
nor U8690 (N_8690,N_4376,N_4581);
and U8691 (N_8691,N_5264,N_5431);
and U8692 (N_8692,N_4456,N_5080);
xnor U8693 (N_8693,N_5571,N_3636);
xor U8694 (N_8694,N_5542,N_3316);
or U8695 (N_8695,N_5071,N_3437);
nand U8696 (N_8696,N_4677,N_3872);
xor U8697 (N_8697,N_3252,N_5024);
or U8698 (N_8698,N_4152,N_3562);
xor U8699 (N_8699,N_4826,N_4813);
and U8700 (N_8700,N_4357,N_3099);
nand U8701 (N_8701,N_5199,N_5013);
nand U8702 (N_8702,N_4344,N_3412);
nor U8703 (N_8703,N_4954,N_3186);
nor U8704 (N_8704,N_4650,N_3723);
xor U8705 (N_8705,N_4954,N_5799);
and U8706 (N_8706,N_5606,N_4926);
nor U8707 (N_8707,N_3611,N_5281);
nand U8708 (N_8708,N_3940,N_4124);
and U8709 (N_8709,N_5478,N_3070);
nand U8710 (N_8710,N_5932,N_3751);
nand U8711 (N_8711,N_3290,N_4576);
xor U8712 (N_8712,N_4110,N_4295);
or U8713 (N_8713,N_5857,N_4412);
or U8714 (N_8714,N_5202,N_3551);
or U8715 (N_8715,N_3165,N_3833);
and U8716 (N_8716,N_4727,N_4060);
xor U8717 (N_8717,N_3122,N_5731);
or U8718 (N_8718,N_5949,N_3814);
and U8719 (N_8719,N_5642,N_5531);
nand U8720 (N_8720,N_5936,N_5795);
or U8721 (N_8721,N_3921,N_5858);
nand U8722 (N_8722,N_4954,N_4241);
and U8723 (N_8723,N_3341,N_3472);
and U8724 (N_8724,N_4611,N_5830);
nor U8725 (N_8725,N_4373,N_5081);
xnor U8726 (N_8726,N_5711,N_4037);
or U8727 (N_8727,N_4516,N_3433);
or U8728 (N_8728,N_4176,N_4448);
xor U8729 (N_8729,N_4640,N_5241);
nor U8730 (N_8730,N_3882,N_5104);
nor U8731 (N_8731,N_4352,N_3834);
xnor U8732 (N_8732,N_4508,N_4609);
xnor U8733 (N_8733,N_5040,N_5520);
xnor U8734 (N_8734,N_5291,N_5418);
nand U8735 (N_8735,N_4518,N_3346);
or U8736 (N_8736,N_4517,N_3275);
or U8737 (N_8737,N_4756,N_4503);
xor U8738 (N_8738,N_3955,N_3939);
xnor U8739 (N_8739,N_4055,N_3342);
or U8740 (N_8740,N_4432,N_5508);
nor U8741 (N_8741,N_4202,N_3217);
and U8742 (N_8742,N_5843,N_4650);
nor U8743 (N_8743,N_3515,N_4389);
nand U8744 (N_8744,N_5704,N_3019);
nand U8745 (N_8745,N_4076,N_4128);
and U8746 (N_8746,N_4706,N_4206);
xor U8747 (N_8747,N_3024,N_5564);
and U8748 (N_8748,N_3267,N_5726);
xnor U8749 (N_8749,N_4824,N_4738);
and U8750 (N_8750,N_5134,N_5605);
nand U8751 (N_8751,N_5906,N_3714);
and U8752 (N_8752,N_5618,N_5884);
nand U8753 (N_8753,N_4092,N_3642);
and U8754 (N_8754,N_4526,N_4863);
and U8755 (N_8755,N_5935,N_3598);
nand U8756 (N_8756,N_3756,N_5847);
nand U8757 (N_8757,N_4603,N_5365);
or U8758 (N_8758,N_3907,N_3338);
or U8759 (N_8759,N_4428,N_4561);
and U8760 (N_8760,N_5885,N_5069);
and U8761 (N_8761,N_4133,N_5436);
nand U8762 (N_8762,N_3321,N_4700);
xnor U8763 (N_8763,N_3028,N_5253);
xor U8764 (N_8764,N_5141,N_4695);
xor U8765 (N_8765,N_3834,N_4347);
or U8766 (N_8766,N_3854,N_5780);
or U8767 (N_8767,N_3287,N_4625);
and U8768 (N_8768,N_4885,N_3358);
and U8769 (N_8769,N_3100,N_5467);
or U8770 (N_8770,N_4226,N_3861);
nor U8771 (N_8771,N_3308,N_4185);
or U8772 (N_8772,N_4860,N_4487);
or U8773 (N_8773,N_4738,N_5871);
nand U8774 (N_8774,N_3517,N_4511);
nor U8775 (N_8775,N_5122,N_4638);
nor U8776 (N_8776,N_5865,N_4775);
nor U8777 (N_8777,N_5066,N_5791);
xnor U8778 (N_8778,N_5102,N_3280);
xor U8779 (N_8779,N_4812,N_5624);
nand U8780 (N_8780,N_3499,N_3075);
or U8781 (N_8781,N_5186,N_3100);
and U8782 (N_8782,N_5537,N_4338);
or U8783 (N_8783,N_3131,N_5818);
nand U8784 (N_8784,N_4676,N_3842);
and U8785 (N_8785,N_3638,N_5934);
xor U8786 (N_8786,N_5816,N_3572);
xor U8787 (N_8787,N_5806,N_3743);
and U8788 (N_8788,N_5603,N_4011);
nor U8789 (N_8789,N_5777,N_4962);
or U8790 (N_8790,N_4168,N_4525);
nor U8791 (N_8791,N_4215,N_4741);
or U8792 (N_8792,N_3572,N_4287);
nand U8793 (N_8793,N_5795,N_5676);
xor U8794 (N_8794,N_5105,N_3531);
xnor U8795 (N_8795,N_3085,N_3861);
nand U8796 (N_8796,N_4667,N_4404);
nand U8797 (N_8797,N_5981,N_5253);
and U8798 (N_8798,N_4053,N_3390);
nor U8799 (N_8799,N_4282,N_5115);
and U8800 (N_8800,N_5381,N_4796);
nand U8801 (N_8801,N_4198,N_4303);
and U8802 (N_8802,N_3532,N_3679);
and U8803 (N_8803,N_5660,N_5569);
nor U8804 (N_8804,N_4704,N_5456);
xor U8805 (N_8805,N_4340,N_4849);
nand U8806 (N_8806,N_5138,N_4136);
and U8807 (N_8807,N_4550,N_4941);
nand U8808 (N_8808,N_3570,N_4925);
nand U8809 (N_8809,N_5358,N_5546);
nand U8810 (N_8810,N_5389,N_5481);
or U8811 (N_8811,N_5990,N_4461);
xor U8812 (N_8812,N_3188,N_4486);
and U8813 (N_8813,N_3956,N_5257);
or U8814 (N_8814,N_3442,N_4406);
nand U8815 (N_8815,N_4159,N_5749);
or U8816 (N_8816,N_4387,N_3963);
xor U8817 (N_8817,N_4559,N_5305);
and U8818 (N_8818,N_4073,N_5250);
and U8819 (N_8819,N_3390,N_5582);
nand U8820 (N_8820,N_3083,N_5478);
nand U8821 (N_8821,N_3455,N_3699);
or U8822 (N_8822,N_4895,N_5075);
xor U8823 (N_8823,N_3400,N_5173);
nand U8824 (N_8824,N_5429,N_3751);
nand U8825 (N_8825,N_5724,N_3051);
nor U8826 (N_8826,N_5789,N_3562);
nand U8827 (N_8827,N_3711,N_4246);
nand U8828 (N_8828,N_3618,N_3151);
nand U8829 (N_8829,N_3794,N_4083);
xnor U8830 (N_8830,N_4317,N_5216);
nand U8831 (N_8831,N_3096,N_3051);
nor U8832 (N_8832,N_4500,N_3783);
xnor U8833 (N_8833,N_3694,N_4315);
or U8834 (N_8834,N_4408,N_5780);
and U8835 (N_8835,N_4201,N_5633);
and U8836 (N_8836,N_5083,N_3006);
nand U8837 (N_8837,N_4663,N_5826);
nor U8838 (N_8838,N_5181,N_4339);
nor U8839 (N_8839,N_5872,N_4762);
and U8840 (N_8840,N_3040,N_5561);
nand U8841 (N_8841,N_5519,N_5677);
nand U8842 (N_8842,N_3103,N_3849);
nor U8843 (N_8843,N_5776,N_3702);
or U8844 (N_8844,N_5650,N_5431);
nand U8845 (N_8845,N_5608,N_5892);
xor U8846 (N_8846,N_5639,N_5635);
xnor U8847 (N_8847,N_5820,N_4787);
nor U8848 (N_8848,N_3236,N_4321);
or U8849 (N_8849,N_4399,N_3452);
or U8850 (N_8850,N_5713,N_3641);
and U8851 (N_8851,N_4461,N_3705);
nor U8852 (N_8852,N_5807,N_3881);
xor U8853 (N_8853,N_5419,N_5090);
xnor U8854 (N_8854,N_3896,N_4958);
nand U8855 (N_8855,N_5544,N_5966);
nor U8856 (N_8856,N_5176,N_3920);
nor U8857 (N_8857,N_5118,N_4838);
nor U8858 (N_8858,N_3341,N_5243);
nor U8859 (N_8859,N_3989,N_5218);
and U8860 (N_8860,N_4201,N_4381);
nor U8861 (N_8861,N_3367,N_3178);
and U8862 (N_8862,N_4291,N_4835);
nor U8863 (N_8863,N_3474,N_5042);
xnor U8864 (N_8864,N_4857,N_5531);
or U8865 (N_8865,N_3576,N_3669);
nor U8866 (N_8866,N_3068,N_5523);
xor U8867 (N_8867,N_3136,N_3524);
or U8868 (N_8868,N_4485,N_5773);
and U8869 (N_8869,N_4669,N_4390);
nand U8870 (N_8870,N_5815,N_3484);
nor U8871 (N_8871,N_3035,N_4932);
nand U8872 (N_8872,N_5410,N_3116);
xor U8873 (N_8873,N_3680,N_4415);
xnor U8874 (N_8874,N_3945,N_5244);
nor U8875 (N_8875,N_4901,N_3348);
and U8876 (N_8876,N_5631,N_5306);
nand U8877 (N_8877,N_4221,N_4337);
nand U8878 (N_8878,N_4831,N_4950);
nand U8879 (N_8879,N_4102,N_5177);
or U8880 (N_8880,N_4907,N_4597);
or U8881 (N_8881,N_3979,N_5663);
and U8882 (N_8882,N_3734,N_3700);
and U8883 (N_8883,N_5895,N_5968);
and U8884 (N_8884,N_5690,N_5463);
nand U8885 (N_8885,N_4466,N_5875);
or U8886 (N_8886,N_3311,N_3881);
or U8887 (N_8887,N_5073,N_5031);
xnor U8888 (N_8888,N_5759,N_3606);
and U8889 (N_8889,N_3042,N_4324);
nor U8890 (N_8890,N_4342,N_4096);
nor U8891 (N_8891,N_5462,N_4334);
nand U8892 (N_8892,N_5651,N_5166);
nor U8893 (N_8893,N_3317,N_4768);
and U8894 (N_8894,N_3981,N_4951);
or U8895 (N_8895,N_5173,N_5207);
nor U8896 (N_8896,N_5070,N_5241);
nand U8897 (N_8897,N_5884,N_3365);
nor U8898 (N_8898,N_5706,N_4164);
or U8899 (N_8899,N_4471,N_3916);
nor U8900 (N_8900,N_4648,N_4539);
nand U8901 (N_8901,N_3598,N_4493);
and U8902 (N_8902,N_3412,N_4620);
nor U8903 (N_8903,N_5139,N_5485);
nand U8904 (N_8904,N_4082,N_3099);
or U8905 (N_8905,N_3608,N_5927);
nand U8906 (N_8906,N_3385,N_4674);
or U8907 (N_8907,N_5681,N_4740);
or U8908 (N_8908,N_5152,N_3569);
xnor U8909 (N_8909,N_5475,N_4507);
or U8910 (N_8910,N_5499,N_4248);
nor U8911 (N_8911,N_4137,N_3209);
nand U8912 (N_8912,N_3086,N_5211);
nand U8913 (N_8913,N_3584,N_3396);
and U8914 (N_8914,N_3197,N_4037);
and U8915 (N_8915,N_3604,N_4376);
or U8916 (N_8916,N_4002,N_5506);
nor U8917 (N_8917,N_4390,N_3222);
nand U8918 (N_8918,N_4633,N_5250);
xnor U8919 (N_8919,N_5894,N_4320);
or U8920 (N_8920,N_4731,N_3017);
nor U8921 (N_8921,N_3302,N_4103);
xnor U8922 (N_8922,N_4157,N_5252);
xnor U8923 (N_8923,N_4416,N_5729);
nor U8924 (N_8924,N_3950,N_3497);
nand U8925 (N_8925,N_4975,N_5591);
nor U8926 (N_8926,N_5537,N_4500);
or U8927 (N_8927,N_3337,N_3362);
nand U8928 (N_8928,N_4638,N_3200);
and U8929 (N_8929,N_3470,N_3274);
xor U8930 (N_8930,N_4408,N_4151);
or U8931 (N_8931,N_3191,N_5555);
nand U8932 (N_8932,N_5097,N_5614);
xnor U8933 (N_8933,N_4205,N_4959);
xor U8934 (N_8934,N_4608,N_3921);
and U8935 (N_8935,N_5266,N_4010);
nor U8936 (N_8936,N_3548,N_3461);
nor U8937 (N_8937,N_5853,N_4608);
nand U8938 (N_8938,N_5471,N_4775);
nor U8939 (N_8939,N_5149,N_3621);
or U8940 (N_8940,N_5789,N_3967);
and U8941 (N_8941,N_3630,N_4890);
or U8942 (N_8942,N_5139,N_3100);
xor U8943 (N_8943,N_3543,N_5895);
and U8944 (N_8944,N_4339,N_4672);
or U8945 (N_8945,N_4313,N_4972);
xor U8946 (N_8946,N_4549,N_3011);
xor U8947 (N_8947,N_3836,N_4416);
nand U8948 (N_8948,N_3529,N_4802);
nand U8949 (N_8949,N_3804,N_5276);
nand U8950 (N_8950,N_3352,N_4085);
xor U8951 (N_8951,N_4238,N_3023);
nand U8952 (N_8952,N_3314,N_5319);
xor U8953 (N_8953,N_3701,N_5465);
nor U8954 (N_8954,N_5605,N_3384);
xnor U8955 (N_8955,N_4371,N_3955);
xnor U8956 (N_8956,N_3536,N_3072);
or U8957 (N_8957,N_3026,N_4400);
and U8958 (N_8958,N_3092,N_4059);
nor U8959 (N_8959,N_5365,N_5066);
and U8960 (N_8960,N_4497,N_3571);
xnor U8961 (N_8961,N_3940,N_4093);
nor U8962 (N_8962,N_5228,N_4418);
xor U8963 (N_8963,N_5116,N_5977);
or U8964 (N_8964,N_4272,N_4360);
nor U8965 (N_8965,N_4238,N_4949);
nand U8966 (N_8966,N_3934,N_3063);
nor U8967 (N_8967,N_5378,N_4074);
xor U8968 (N_8968,N_4345,N_4660);
nand U8969 (N_8969,N_4960,N_4067);
nor U8970 (N_8970,N_4874,N_4580);
xor U8971 (N_8971,N_5048,N_3943);
or U8972 (N_8972,N_3691,N_4393);
nor U8973 (N_8973,N_4274,N_5485);
nand U8974 (N_8974,N_3510,N_3780);
nor U8975 (N_8975,N_4004,N_4313);
nor U8976 (N_8976,N_3725,N_3662);
xnor U8977 (N_8977,N_3131,N_3471);
nand U8978 (N_8978,N_5026,N_3468);
nor U8979 (N_8979,N_4943,N_5471);
or U8980 (N_8980,N_3625,N_3225);
and U8981 (N_8981,N_3667,N_4241);
xor U8982 (N_8982,N_4678,N_5492);
nor U8983 (N_8983,N_5948,N_5605);
xor U8984 (N_8984,N_4222,N_4988);
and U8985 (N_8985,N_4448,N_3619);
xnor U8986 (N_8986,N_3646,N_4993);
nand U8987 (N_8987,N_3378,N_5973);
xnor U8988 (N_8988,N_4361,N_3592);
nor U8989 (N_8989,N_4183,N_4352);
nand U8990 (N_8990,N_5354,N_4989);
nand U8991 (N_8991,N_4609,N_3220);
xnor U8992 (N_8992,N_3580,N_3660);
and U8993 (N_8993,N_5511,N_5798);
xnor U8994 (N_8994,N_4842,N_5368);
or U8995 (N_8995,N_5466,N_5760);
xnor U8996 (N_8996,N_5342,N_4951);
or U8997 (N_8997,N_5433,N_5597);
nor U8998 (N_8998,N_4369,N_3549);
or U8999 (N_8999,N_3760,N_3083);
or U9000 (N_9000,N_8053,N_7350);
xnor U9001 (N_9001,N_8649,N_8580);
or U9002 (N_9002,N_7266,N_6405);
xor U9003 (N_9003,N_7883,N_6248);
xor U9004 (N_9004,N_7074,N_8797);
or U9005 (N_9005,N_6069,N_8047);
nor U9006 (N_9006,N_6275,N_7815);
nand U9007 (N_9007,N_6931,N_6397);
nand U9008 (N_9008,N_8656,N_8727);
nor U9009 (N_9009,N_8618,N_7889);
nand U9010 (N_9010,N_7015,N_6823);
nor U9011 (N_9011,N_7417,N_7060);
nor U9012 (N_9012,N_6052,N_6856);
and U9013 (N_9013,N_7032,N_6260);
or U9014 (N_9014,N_7274,N_7606);
and U9015 (N_9015,N_6630,N_6735);
or U9016 (N_9016,N_7813,N_7081);
nand U9017 (N_9017,N_6632,N_8723);
nand U9018 (N_9018,N_8241,N_8542);
nand U9019 (N_9019,N_7721,N_6624);
nor U9020 (N_9020,N_8225,N_8718);
xnor U9021 (N_9021,N_8486,N_7628);
xor U9022 (N_9022,N_6374,N_6106);
nand U9023 (N_9023,N_7657,N_8264);
nand U9024 (N_9024,N_8413,N_8434);
xnor U9025 (N_9025,N_8508,N_7441);
and U9026 (N_9026,N_7142,N_8666);
xor U9027 (N_9027,N_8479,N_7533);
nor U9028 (N_9028,N_8040,N_8891);
nand U9029 (N_9029,N_7182,N_6977);
and U9030 (N_9030,N_8669,N_7428);
xor U9031 (N_9031,N_8537,N_6576);
and U9032 (N_9032,N_7347,N_8122);
nor U9033 (N_9033,N_6765,N_8562);
and U9034 (N_9034,N_6080,N_8771);
nand U9035 (N_9035,N_7946,N_7555);
and U9036 (N_9036,N_7808,N_6693);
nor U9037 (N_9037,N_6269,N_7311);
or U9038 (N_9038,N_8871,N_7020);
nand U9039 (N_9039,N_6398,N_8118);
and U9040 (N_9040,N_6682,N_7478);
or U9041 (N_9041,N_7245,N_8152);
and U9042 (N_9042,N_8108,N_8176);
nor U9043 (N_9043,N_6886,N_6120);
nand U9044 (N_9044,N_6998,N_6510);
nor U9045 (N_9045,N_7974,N_7470);
nand U9046 (N_9046,N_8004,N_7850);
nand U9047 (N_9047,N_6512,N_7246);
and U9048 (N_9048,N_8136,N_6980);
xor U9049 (N_9049,N_7139,N_6564);
xnor U9050 (N_9050,N_7586,N_8557);
and U9051 (N_9051,N_8138,N_8127);
nor U9052 (N_9052,N_6831,N_6007);
xor U9053 (N_9053,N_7854,N_8412);
nor U9054 (N_9054,N_6759,N_7297);
and U9055 (N_9055,N_7689,N_6708);
and U9056 (N_9056,N_6150,N_6699);
nor U9057 (N_9057,N_8731,N_6905);
xnor U9058 (N_9058,N_6943,N_8778);
nand U9059 (N_9059,N_8392,N_7123);
xor U9060 (N_9060,N_8359,N_7022);
nand U9061 (N_9061,N_6655,N_7528);
or U9062 (N_9062,N_7408,N_6770);
nor U9063 (N_9063,N_7140,N_7442);
or U9064 (N_9064,N_6393,N_8998);
nand U9065 (N_9065,N_8515,N_8023);
nand U9066 (N_9066,N_7039,N_7371);
xnor U9067 (N_9067,N_8282,N_8450);
or U9068 (N_9068,N_8583,N_6557);
and U9069 (N_9069,N_7093,N_6111);
and U9070 (N_9070,N_8112,N_6263);
nor U9071 (N_9071,N_7686,N_6809);
nor U9072 (N_9072,N_7930,N_6800);
xor U9073 (N_9073,N_6361,N_7698);
and U9074 (N_9074,N_8010,N_6928);
and U9075 (N_9075,N_8663,N_8061);
nor U9076 (N_9076,N_6306,N_7783);
and U9077 (N_9077,N_7121,N_8608);
and U9078 (N_9078,N_8978,N_7531);
or U9079 (N_9079,N_6371,N_6684);
or U9080 (N_9080,N_7912,N_8157);
and U9081 (N_9081,N_7503,N_6417);
nor U9082 (N_9082,N_8875,N_7100);
xnor U9083 (N_9083,N_7413,N_7460);
and U9084 (N_9084,N_6554,N_7435);
nand U9085 (N_9085,N_7087,N_7083);
nand U9086 (N_9086,N_6135,N_7208);
or U9087 (N_9087,N_6325,N_8383);
and U9088 (N_9088,N_8992,N_7876);
xor U9089 (N_9089,N_7482,N_8020);
and U9090 (N_9090,N_8699,N_8624);
xor U9091 (N_9091,N_7711,N_7046);
nor U9092 (N_9092,N_6020,N_8469);
or U9093 (N_9093,N_8726,N_7702);
and U9094 (N_9094,N_8953,N_6854);
xnor U9095 (N_9095,N_8928,N_6565);
nor U9096 (N_9096,N_6331,N_8623);
nor U9097 (N_9097,N_7222,N_7937);
or U9098 (N_9098,N_7444,N_7249);
and U9099 (N_9099,N_7017,N_6567);
nand U9100 (N_9100,N_6382,N_7013);
xor U9101 (N_9101,N_6047,N_7061);
xnor U9102 (N_9102,N_6024,N_6816);
and U9103 (N_9103,N_6220,N_8711);
nand U9104 (N_9104,N_6340,N_8814);
and U9105 (N_9105,N_6502,N_7469);
or U9106 (N_9106,N_7364,N_6232);
xor U9107 (N_9107,N_8568,N_7621);
or U9108 (N_9108,N_8346,N_6892);
xor U9109 (N_9109,N_7498,N_7181);
xor U9110 (N_9110,N_7668,N_6863);
nor U9111 (N_9111,N_6021,N_7662);
or U9112 (N_9112,N_7986,N_7941);
and U9113 (N_9113,N_6857,N_8237);
xor U9114 (N_9114,N_7614,N_7525);
xor U9115 (N_9115,N_8252,N_6256);
xnor U9116 (N_9116,N_7664,N_6312);
and U9117 (N_9117,N_7105,N_8251);
nor U9118 (N_9118,N_7911,N_6960);
or U9119 (N_9119,N_8552,N_8193);
and U9120 (N_9120,N_7737,N_7620);
and U9121 (N_9121,N_8043,N_6776);
or U9122 (N_9122,N_7197,N_8309);
xor U9123 (N_9123,N_6546,N_7701);
or U9124 (N_9124,N_6628,N_8038);
nor U9125 (N_9125,N_8103,N_7573);
or U9126 (N_9126,N_8235,N_6240);
or U9127 (N_9127,N_8086,N_7425);
and U9128 (N_9128,N_6391,N_8394);
and U9129 (N_9129,N_8179,N_7284);
xnor U9130 (N_9130,N_7908,N_7910);
xor U9131 (N_9131,N_7881,N_8214);
and U9132 (N_9132,N_6710,N_6721);
nand U9133 (N_9133,N_7491,N_8400);
and U9134 (N_9134,N_7127,N_7199);
nand U9135 (N_9135,N_8211,N_8755);
or U9136 (N_9136,N_8801,N_7501);
xor U9137 (N_9137,N_6638,N_6797);
nand U9138 (N_9138,N_7654,N_6430);
nor U9139 (N_9139,N_6437,N_8472);
nor U9140 (N_9140,N_7424,N_8824);
or U9141 (N_9141,N_8795,N_8279);
nand U9142 (N_9142,N_7273,N_6200);
nor U9143 (N_9143,N_6744,N_8156);
and U9144 (N_9144,N_7844,N_6485);
xnor U9145 (N_9145,N_7134,N_8027);
nand U9146 (N_9146,N_7118,N_6817);
and U9147 (N_9147,N_7892,N_6073);
nor U9148 (N_9148,N_8949,N_8126);
or U9149 (N_9149,N_8606,N_8387);
xor U9150 (N_9150,N_8367,N_7331);
or U9151 (N_9151,N_8312,N_8599);
nor U9152 (N_9152,N_8072,N_6184);
nor U9153 (N_9153,N_7079,N_6303);
xor U9154 (N_9154,N_8826,N_8658);
or U9155 (N_9155,N_6468,N_8468);
or U9156 (N_9156,N_7151,N_8742);
xnor U9157 (N_9157,N_6246,N_8338);
nand U9158 (N_9158,N_6734,N_6631);
nand U9159 (N_9159,N_8952,N_8044);
or U9160 (N_9160,N_8737,N_8407);
nor U9161 (N_9161,N_8498,N_8739);
nor U9162 (N_9162,N_7292,N_7630);
or U9163 (N_9163,N_7680,N_8673);
xnor U9164 (N_9164,N_6652,N_7097);
and U9165 (N_9165,N_6225,N_7120);
nor U9166 (N_9166,N_8900,N_6364);
and U9167 (N_9167,N_6044,N_8328);
nor U9168 (N_9168,N_6566,N_7302);
nand U9169 (N_9169,N_6757,N_7314);
nand U9170 (N_9170,N_8194,N_8465);
nor U9171 (N_9171,N_8474,N_6028);
or U9172 (N_9172,N_7597,N_8230);
nor U9173 (N_9173,N_8477,N_6660);
and U9174 (N_9174,N_6948,N_8728);
nor U9175 (N_9175,N_8389,N_6849);
and U9176 (N_9176,N_7027,N_7923);
xor U9177 (N_9177,N_6491,N_7148);
xor U9178 (N_9178,N_7255,N_7465);
xor U9179 (N_9179,N_8262,N_8811);
nand U9180 (N_9180,N_7530,N_6792);
or U9181 (N_9181,N_6054,N_7564);
and U9182 (N_9182,N_6968,N_8182);
nand U9183 (N_9183,N_7797,N_7426);
and U9184 (N_9184,N_7798,N_7637);
nand U9185 (N_9185,N_7014,N_8266);
nor U9186 (N_9186,N_7994,N_8609);
xor U9187 (N_9187,N_7320,N_6846);
nand U9188 (N_9188,N_8594,N_8117);
xnor U9189 (N_9189,N_7190,N_6100);
and U9190 (N_9190,N_8839,N_8153);
and U9191 (N_9191,N_7975,N_7366);
xnor U9192 (N_9192,N_7295,N_7078);
xnor U9193 (N_9193,N_6223,N_7861);
nand U9194 (N_9194,N_8749,N_8935);
nor U9195 (N_9195,N_7834,N_6992);
xnor U9196 (N_9196,N_6818,N_8816);
nor U9197 (N_9197,N_8294,N_7965);
xor U9198 (N_9198,N_8793,N_7751);
xnor U9199 (N_9199,N_8089,N_8854);
or U9200 (N_9200,N_6961,N_8591);
and U9201 (N_9201,N_7972,N_8827);
nand U9202 (N_9202,N_8031,N_8948);
and U9203 (N_9203,N_6089,N_6473);
xor U9204 (N_9204,N_7349,N_7041);
xnor U9205 (N_9205,N_7040,N_6455);
nor U9206 (N_9206,N_7997,N_6134);
and U9207 (N_9207,N_8535,N_7542);
nand U9208 (N_9208,N_6467,N_6066);
nor U9209 (N_9209,N_6890,N_8621);
and U9210 (N_9210,N_8203,N_8180);
nor U9211 (N_9211,N_7155,N_8614);
nand U9212 (N_9212,N_8734,N_8188);
nand U9213 (N_9213,N_7432,N_7033);
nand U9214 (N_9214,N_6379,N_6456);
nor U9215 (N_9215,N_7944,N_7954);
and U9216 (N_9216,N_7045,N_8912);
xor U9217 (N_9217,N_6577,N_7192);
and U9218 (N_9218,N_8611,N_7259);
xnor U9219 (N_9219,N_7541,N_8751);
xnor U9220 (N_9220,N_8448,N_7277);
or U9221 (N_9221,N_6880,N_8961);
xnor U9222 (N_9222,N_6019,N_8841);
nand U9223 (N_9223,N_8996,N_7981);
nand U9224 (N_9224,N_8925,N_8989);
nor U9225 (N_9225,N_6940,N_7544);
nand U9226 (N_9226,N_7452,N_8698);
xnor U9227 (N_9227,N_7323,N_6471);
xnor U9228 (N_9228,N_6585,N_6844);
or U9229 (N_9229,N_7740,N_7567);
and U9230 (N_9230,N_8725,N_7260);
nor U9231 (N_9231,N_6193,N_6032);
or U9232 (N_9232,N_7005,N_8140);
nor U9233 (N_9233,N_8784,N_7955);
nor U9234 (N_9234,N_6017,N_8246);
or U9235 (N_9235,N_8914,N_8813);
nor U9236 (N_9236,N_6582,N_7096);
xnor U9237 (N_9237,N_8414,N_7308);
and U9238 (N_9238,N_8098,N_8019);
or U9239 (N_9239,N_6202,N_8372);
nor U9240 (N_9240,N_7703,N_8765);
or U9241 (N_9241,N_6683,N_7310);
nand U9242 (N_9242,N_6380,N_6216);
nor U9243 (N_9243,N_7514,N_6443);
or U9244 (N_9244,N_7560,N_7028);
or U9245 (N_9245,N_6974,N_8085);
and U9246 (N_9246,N_6668,N_7227);
nand U9247 (N_9247,N_6899,N_7925);
and U9248 (N_9248,N_6215,N_6501);
and U9249 (N_9249,N_8348,N_7440);
or U9250 (N_9250,N_7601,N_7485);
nor U9251 (N_9251,N_6506,N_8073);
xor U9252 (N_9252,N_8482,N_6090);
or U9253 (N_9253,N_8582,N_6581);
nor U9254 (N_9254,N_7261,N_6571);
nand U9255 (N_9255,N_6056,N_7539);
and U9256 (N_9256,N_7879,N_8025);
nand U9257 (N_9257,N_8101,N_6698);
or U9258 (N_9258,N_8364,N_7901);
and U9259 (N_9259,N_7557,N_8872);
xor U9260 (N_9260,N_7769,N_7419);
nand U9261 (N_9261,N_6213,N_7860);
or U9262 (N_9262,N_7782,N_6038);
nand U9263 (N_9263,N_8286,N_7644);
nand U9264 (N_9264,N_6715,N_8870);
nand U9265 (N_9265,N_6040,N_6014);
nor U9266 (N_9266,N_7177,N_6167);
xnor U9267 (N_9267,N_8759,N_7696);
or U9268 (N_9268,N_8955,N_8302);
nor U9269 (N_9269,N_7859,N_7619);
and U9270 (N_9270,N_6690,N_6808);
nand U9271 (N_9271,N_6094,N_8080);
or U9272 (N_9272,N_6913,N_7629);
xnor U9273 (N_9273,N_6423,N_7225);
nand U9274 (N_9274,N_7642,N_8090);
nor U9275 (N_9275,N_7509,N_7653);
xor U9276 (N_9276,N_7993,N_8837);
or U9277 (N_9277,N_8183,N_7483);
nor U9278 (N_9278,N_6142,N_6489);
xor U9279 (N_9279,N_7256,N_8174);
and U9280 (N_9280,N_8172,N_8067);
and U9281 (N_9281,N_8524,N_6874);
or U9282 (N_9282,N_6869,N_7552);
or U9283 (N_9283,N_7907,N_8499);
nand U9284 (N_9284,N_6716,N_6908);
and U9285 (N_9285,N_7112,N_6815);
nand U9286 (N_9286,N_8865,N_8598);
xor U9287 (N_9287,N_8459,N_7391);
xnor U9288 (N_9288,N_6560,N_6114);
nand U9289 (N_9289,N_8306,N_7089);
nor U9290 (N_9290,N_7523,N_6933);
or U9291 (N_9291,N_8066,N_8794);
or U9292 (N_9292,N_6401,N_8075);
nor U9293 (N_9293,N_7300,N_7400);
and U9294 (N_9294,N_6426,N_7729);
nand U9295 (N_9295,N_8260,N_6626);
and U9296 (N_9296,N_6877,N_7857);
nand U9297 (N_9297,N_7195,N_6763);
and U9298 (N_9298,N_7145,N_7158);
and U9299 (N_9299,N_7149,N_7681);
nor U9300 (N_9300,N_7584,N_7734);
nor U9301 (N_9301,N_8132,N_6420);
xor U9302 (N_9302,N_8983,N_8485);
or U9303 (N_9303,N_8154,N_7571);
and U9304 (N_9304,N_8944,N_7720);
nor U9305 (N_9305,N_7431,N_6299);
and U9306 (N_9306,N_6592,N_6962);
nand U9307 (N_9307,N_8984,N_6875);
xor U9308 (N_9308,N_8631,N_7404);
nand U9309 (N_9309,N_6300,N_8950);
or U9310 (N_9310,N_8269,N_7461);
and U9311 (N_9311,N_7447,N_7753);
or U9312 (N_9312,N_7126,N_7507);
xnor U9313 (N_9313,N_7655,N_8045);
or U9314 (N_9314,N_8095,N_7385);
and U9315 (N_9315,N_8972,N_6217);
nor U9316 (N_9316,N_6733,N_8936);
or U9317 (N_9317,N_8377,N_6677);
nor U9318 (N_9318,N_7414,N_7612);
or U9319 (N_9319,N_7237,N_6870);
nand U9320 (N_9320,N_8494,N_8847);
nor U9321 (N_9321,N_6568,N_7421);
xor U9322 (N_9322,N_6357,N_7239);
and U9323 (N_9323,N_7392,N_7229);
nand U9324 (N_9324,N_6894,N_7489);
nand U9325 (N_9325,N_6450,N_6258);
nor U9326 (N_9326,N_8920,N_7026);
nand U9327 (N_9327,N_6952,N_7477);
nand U9328 (N_9328,N_7024,N_6889);
nor U9329 (N_9329,N_8300,N_6058);
and U9330 (N_9330,N_6151,N_6459);
and U9331 (N_9331,N_7914,N_6589);
nand U9332 (N_9332,N_6127,N_6881);
nand U9333 (N_9333,N_8908,N_6505);
nand U9334 (N_9334,N_7618,N_8595);
xor U9335 (N_9335,N_8283,N_6041);
and U9336 (N_9336,N_7835,N_7104);
and U9337 (N_9337,N_6686,N_8504);
nand U9338 (N_9338,N_6729,N_8069);
nand U9339 (N_9339,N_6453,N_7982);
nor U9340 (N_9340,N_8777,N_8428);
and U9341 (N_9341,N_8810,N_6376);
nor U9342 (N_9342,N_6647,N_6230);
xnor U9343 (N_9343,N_6309,N_8626);
and U9344 (N_9344,N_7138,N_7167);
and U9345 (N_9345,N_6915,N_7639);
and U9346 (N_9346,N_8643,N_8454);
or U9347 (N_9347,N_7108,N_7231);
and U9348 (N_9348,N_8048,N_6646);
or U9349 (N_9349,N_6483,N_6852);
and U9350 (N_9350,N_6117,N_7880);
nand U9351 (N_9351,N_6556,N_6113);
nand U9352 (N_9352,N_8079,N_8977);
and U9353 (N_9353,N_6137,N_6971);
and U9354 (N_9354,N_6146,N_8789);
xnor U9355 (N_9355,N_7738,N_8886);
or U9356 (N_9356,N_8703,N_6820);
and U9357 (N_9357,N_7152,N_8767);
or U9358 (N_9358,N_6641,N_7742);
and U9359 (N_9359,N_8956,N_6249);
nand U9360 (N_9360,N_8615,N_8701);
nor U9361 (N_9361,N_8327,N_8245);
or U9362 (N_9362,N_6558,N_7257);
or U9363 (N_9363,N_8016,N_6487);
nor U9364 (N_9364,N_7929,N_7464);
and U9365 (N_9365,N_7538,N_6280);
nand U9366 (N_9366,N_8408,N_6995);
or U9367 (N_9367,N_7852,N_7887);
and U9368 (N_9368,N_8976,N_8966);
nor U9369 (N_9369,N_8880,N_8253);
or U9370 (N_9370,N_6742,N_7438);
and U9371 (N_9371,N_7189,N_7793);
xnor U9372 (N_9372,N_6685,N_6779);
or U9373 (N_9373,N_7504,N_6944);
xor U9374 (N_9374,N_7580,N_7842);
and U9375 (N_9375,N_6062,N_8487);
nor U9376 (N_9376,N_6415,N_6621);
or U9377 (N_9377,N_6553,N_7900);
nor U9378 (N_9378,N_8363,N_7563);
nand U9379 (N_9379,N_8274,N_8541);
nor U9380 (N_9380,N_7018,N_6295);
xnor U9381 (N_9381,N_7577,N_7502);
and U9382 (N_9382,N_8980,N_7940);
xor U9383 (N_9383,N_7643,N_8052);
or U9384 (N_9384,N_7691,N_8005);
and U9385 (N_9385,N_6713,N_8566);
xor U9386 (N_9386,N_8417,N_8772);
xnor U9387 (N_9387,N_8858,N_6001);
xor U9388 (N_9388,N_6804,N_7473);
xor U9389 (N_9389,N_8753,N_6222);
nor U9390 (N_9390,N_8714,N_6738);
nor U9391 (N_9391,N_6344,N_7379);
or U9392 (N_9392,N_6039,N_6907);
nand U9393 (N_9393,N_6527,N_8916);
nand U9394 (N_9394,N_6946,N_7267);
nor U9395 (N_9395,N_7180,N_8890);
nand U9396 (N_9396,N_7114,N_6287);
or U9397 (N_9397,N_6709,N_7168);
xor U9398 (N_9398,N_7500,N_7232);
or U9399 (N_9399,N_7770,N_7520);
xnor U9400 (N_9400,N_7117,N_7547);
nor U9401 (N_9401,N_8201,N_8491);
nor U9402 (N_9402,N_7462,N_8330);
nor U9403 (N_9403,N_8799,N_6182);
nor U9404 (N_9404,N_8804,N_8213);
nor U9405 (N_9405,N_8342,N_6356);
nand U9406 (N_9406,N_7820,N_6659);
and U9407 (N_9407,N_7367,N_6065);
xnor U9408 (N_9408,N_7160,N_6525);
and U9409 (N_9409,N_6707,N_7561);
nor U9410 (N_9410,N_8340,N_8226);
xor U9411 (N_9411,N_8934,N_6172);
nand U9412 (N_9412,N_7848,N_6609);
and U9413 (N_9413,N_7951,N_8446);
or U9414 (N_9414,N_8848,N_8165);
nand U9415 (N_9415,N_8868,N_7186);
nand U9416 (N_9416,N_8303,N_6937);
xnor U9417 (N_9417,N_6323,N_7365);
nand U9418 (N_9418,N_6504,N_7915);
nand U9419 (N_9419,N_8273,N_8385);
nor U9420 (N_9420,N_7672,N_8313);
nand U9421 (N_9421,N_6500,N_7700);
nor U9422 (N_9422,N_8395,N_7480);
and U9423 (N_9423,N_7344,N_8320);
xor U9424 (N_9424,N_8644,N_6319);
and U9425 (N_9425,N_6425,N_7904);
xor U9426 (N_9426,N_7992,N_6392);
xor U9427 (N_9427,N_6787,N_8242);
nor U9428 (N_9428,N_7518,N_7037);
nand U9429 (N_9429,N_6231,N_8050);
nor U9430 (N_9430,N_6718,N_6802);
xor U9431 (N_9431,N_8790,N_7913);
xor U9432 (N_9432,N_8500,N_6131);
or U9433 (N_9433,N_7437,N_8105);
xor U9434 (N_9434,N_8605,N_8798);
nand U9435 (N_9435,N_8191,N_7775);
or U9436 (N_9436,N_8011,N_7157);
xor U9437 (N_9437,N_6979,N_6756);
xnor U9438 (N_9438,N_6949,N_7023);
and U9439 (N_9439,N_6214,N_7652);
xor U9440 (N_9440,N_7673,N_6692);
xnor U9441 (N_9441,N_8445,N_7002);
and U9442 (N_9442,N_8145,N_6318);
and U9443 (N_9443,N_6178,N_8693);
and U9444 (N_9444,N_6611,N_6446);
xor U9445 (N_9445,N_8365,N_6221);
or U9446 (N_9446,N_7694,N_6798);
and U9447 (N_9447,N_8985,N_6695);
or U9448 (N_9448,N_7690,N_8233);
or U9449 (N_9449,N_8710,N_8512);
and U9450 (N_9450,N_6691,N_8271);
xor U9451 (N_9451,N_6761,N_6706);
and U9452 (N_9452,N_8054,N_6334);
nand U9453 (N_9453,N_6158,N_8863);
and U9454 (N_9454,N_8604,N_6368);
or U9455 (N_9455,N_8310,N_7355);
nand U9456 (N_9456,N_8779,N_7317);
or U9457 (N_9457,N_6935,N_8785);
xor U9458 (N_9458,N_8807,N_7724);
nand U9459 (N_9459,N_7886,N_6896);
and U9460 (N_9460,N_7304,N_7136);
nand U9461 (N_9461,N_8135,N_6769);
nand U9462 (N_9462,N_8292,N_8440);
or U9463 (N_9463,N_7316,N_6128);
nor U9464 (N_9464,N_7617,N_7307);
nand U9465 (N_9465,N_8037,N_8563);
and U9466 (N_9466,N_7293,N_7803);
nor U9467 (N_9467,N_7692,N_8760);
or U9468 (N_9468,N_6369,N_6270);
xnor U9469 (N_9469,N_7263,N_8888);
nand U9470 (N_9470,N_7056,N_7905);
nor U9471 (N_9471,N_6110,N_6234);
and U9472 (N_9472,N_7334,N_7236);
nand U9473 (N_9473,N_6345,N_8256);
nand U9474 (N_9474,N_6067,N_8697);
and U9475 (N_9475,N_7247,N_8208);
nor U9476 (N_9476,N_8991,N_8918);
nand U9477 (N_9477,N_8489,N_6244);
and U9478 (N_9478,N_6042,N_7932);
nand U9479 (N_9479,N_6916,N_6520);
and U9480 (N_9480,N_7741,N_7987);
nor U9481 (N_9481,N_8325,N_7458);
nor U9482 (N_9482,N_6827,N_7807);
or U9483 (N_9483,N_8349,N_7745);
nand U9484 (N_9484,N_8046,N_6136);
or U9485 (N_9485,N_8409,N_8821);
nand U9486 (N_9486,N_8166,N_8336);
and U9487 (N_9487,N_7822,N_6834);
nand U9488 (N_9488,N_6600,N_7732);
nand U9489 (N_9489,N_6956,N_7402);
nor U9490 (N_9490,N_7383,N_7983);
and U9491 (N_9491,N_6012,N_8775);
nand U9492 (N_9492,N_6601,N_7632);
nand U9493 (N_9493,N_8993,N_6112);
and U9494 (N_9494,N_8097,N_6918);
and U9495 (N_9495,N_6604,N_8616);
nor U9496 (N_9496,N_7059,N_8899);
or U9497 (N_9497,N_7873,N_8736);
nand U9498 (N_9498,N_8796,N_6183);
and U9499 (N_9499,N_8752,N_7771);
and U9500 (N_9500,N_8932,N_8943);
or U9501 (N_9501,N_7439,N_7384);
nand U9502 (N_9502,N_6986,N_6917);
and U9503 (N_9503,N_8661,N_7960);
nor U9504 (N_9504,N_6388,N_7615);
or U9505 (N_9505,N_6281,N_8116);
nand U9506 (N_9506,N_8036,N_7279);
nand U9507 (N_9507,N_7570,N_8014);
nand U9508 (N_9508,N_6464,N_6068);
xor U9509 (N_9509,N_7159,N_8903);
and U9510 (N_9510,N_6465,N_8818);
or U9511 (N_9511,N_8741,N_8184);
xnor U9512 (N_9512,N_6236,N_7095);
and U9513 (N_9513,N_6845,N_7853);
nor U9514 (N_9514,N_7786,N_8567);
xor U9515 (N_9515,N_6700,N_6064);
and U9516 (N_9516,N_8493,N_7147);
and U9517 (N_9517,N_7877,N_7113);
and U9518 (N_9518,N_6720,N_6255);
and U9519 (N_9519,N_7812,N_6101);
nand U9520 (N_9520,N_8534,N_8913);
and U9521 (N_9521,N_8404,N_8426);
xnor U9522 (N_9522,N_6351,N_6758);
nand U9523 (N_9523,N_8039,N_6201);
xor U9524 (N_9524,N_7496,N_8322);
xor U9525 (N_9525,N_6517,N_8746);
xnor U9526 (N_9526,N_6194,N_8685);
nor U9527 (N_9527,N_8704,N_7343);
or U9528 (N_9528,N_8261,N_8945);
and U9529 (N_9529,N_7731,N_6274);
and U9530 (N_9530,N_8319,N_6088);
or U9531 (N_9531,N_8887,N_7631);
nand U9532 (N_9532,N_6651,N_8593);
nand U9533 (N_9533,N_8973,N_7235);
nor U9534 (N_9534,N_8375,N_8828);
or U9535 (N_9535,N_6662,N_7341);
xnor U9536 (N_9536,N_7084,N_6478);
nand U9537 (N_9537,N_6469,N_6022);
nor U9538 (N_9538,N_6257,N_7036);
xnor U9539 (N_9539,N_7513,N_7517);
nand U9540 (N_9540,N_7090,N_8366);
and U9541 (N_9541,N_8478,N_6503);
nand U9542 (N_9542,N_8447,N_7685);
xor U9543 (N_9543,N_8062,N_8545);
or U9544 (N_9544,N_7339,N_8231);
xnor U9545 (N_9545,N_6132,N_6555);
nand U9546 (N_9546,N_7362,N_6644);
and U9547 (N_9547,N_8690,N_8284);
or U9548 (N_9548,N_6623,N_7991);
nand U9549 (N_9549,N_6003,N_7012);
and U9550 (N_9550,N_7757,N_8502);
and U9551 (N_9551,N_7966,N_8373);
or U9552 (N_9552,N_7143,N_8293);
nor U9553 (N_9553,N_7154,N_8307);
or U9554 (N_9554,N_7602,N_6627);
nor U9555 (N_9555,N_7928,N_8059);
and U9556 (N_9556,N_8715,N_7931);
or U9557 (N_9557,N_6259,N_6121);
or U9558 (N_9558,N_6472,N_7213);
nor U9559 (N_9559,N_7758,N_8436);
and U9560 (N_9560,N_8190,N_8558);
nor U9561 (N_9561,N_7053,N_8559);
and U9562 (N_9562,N_8679,N_8382);
xor U9563 (N_9563,N_7959,N_8250);
xor U9564 (N_9564,N_7324,N_8204);
xor U9565 (N_9565,N_7169,N_8124);
nand U9566 (N_9566,N_8628,N_7851);
and U9567 (N_9567,N_8924,N_6495);
and U9568 (N_9568,N_7948,N_8345);
xnor U9569 (N_9569,N_6910,N_6206);
or U9570 (N_9570,N_6180,N_8405);
or U9571 (N_9571,N_7254,N_8911);
nand U9572 (N_9572,N_6634,N_7710);
or U9573 (N_9573,N_6123,N_7380);
nor U9574 (N_9574,N_8141,N_6059);
nand U9575 (N_9575,N_8756,N_6511);
or U9576 (N_9576,N_8461,N_6588);
nor U9577 (N_9577,N_6959,N_8682);
xnor U9578 (N_9578,N_7575,N_6777);
xnor U9579 (N_9579,N_6951,N_7683);
nor U9580 (N_9580,N_6574,N_6330);
and U9581 (N_9581,N_8331,N_7728);
or U9582 (N_9582,N_7133,N_8719);
nor U9583 (N_9583,N_8695,N_8104);
and U9584 (N_9584,N_8662,N_6622);
and U9585 (N_9585,N_8243,N_7072);
xnor U9586 (N_9586,N_6786,N_6989);
xnor U9587 (N_9587,N_8889,N_7796);
xnor U9588 (N_9588,N_7752,N_8432);
xor U9589 (N_9589,N_6023,N_6705);
or U9590 (N_9590,N_7163,N_8155);
xnor U9591 (N_9591,N_7764,N_7823);
xor U9592 (N_9592,N_7537,N_8287);
nor U9593 (N_9593,N_7636,N_7927);
and U9594 (N_9594,N_7754,N_7649);
nand U9595 (N_9595,N_7258,N_6205);
xor U9596 (N_9596,N_7170,N_8505);
or U9597 (N_9597,N_7451,N_8692);
or U9598 (N_9598,N_6605,N_7129);
or U9599 (N_9599,N_8003,N_8951);
and U9600 (N_9600,N_7203,N_8159);
or U9601 (N_9601,N_8483,N_7902);
nand U9602 (N_9602,N_7472,N_6104);
nand U9603 (N_9603,N_8276,N_8909);
nand U9604 (N_9604,N_6154,N_8119);
nand U9605 (N_9605,N_6129,N_6057);
and U9606 (N_9606,N_6790,N_6541);
nand U9607 (N_9607,N_6728,N_6235);
or U9608 (N_9608,N_6882,N_6987);
nor U9609 (N_9609,N_6840,N_6612);
or U9610 (N_9610,N_7568,N_8411);
nand U9611 (N_9611,N_8522,N_6399);
nor U9612 (N_9612,N_6806,N_6164);
and U9613 (N_9613,N_7368,N_7466);
xor U9614 (N_9614,N_6837,N_6261);
nor U9615 (N_9615,N_7800,N_8437);
and U9616 (N_9616,N_7209,N_8556);
nand U9617 (N_9617,N_6412,N_7875);
xor U9618 (N_9618,N_6814,N_7166);
and U9619 (N_9619,N_7942,N_7616);
nor U9620 (N_9620,N_8380,N_7869);
xor U9621 (N_9621,N_7356,N_6550);
and U9622 (N_9622,N_7193,N_8721);
nand U9623 (N_9623,N_7824,N_6526);
nor U9624 (N_9624,N_8637,N_6452);
and U9625 (N_9625,N_8851,N_6189);
nor U9626 (N_9626,N_7976,N_8809);
and U9627 (N_9627,N_6533,N_7953);
or U9628 (N_9628,N_7009,N_6324);
or U9629 (N_9629,N_6276,N_8532);
xor U9630 (N_9630,N_6640,N_7663);
nor U9631 (N_9631,N_7395,N_8906);
and U9632 (N_9632,N_6428,N_6925);
nand U9633 (N_9633,N_6670,N_6703);
nor U9634 (N_9634,N_7184,N_8974);
xor U9635 (N_9635,N_7545,N_8351);
and U9636 (N_9636,N_6642,N_6593);
xor U9637 (N_9637,N_7433,N_8270);
or U9638 (N_9638,N_8519,N_6615);
xor U9639 (N_9639,N_7527,N_8987);
xnor U9640 (N_9640,N_8901,N_6887);
nor U9641 (N_9641,N_8540,N_6370);
nor U9642 (N_9642,N_8647,N_7936);
or U9643 (N_9643,N_8185,N_7080);
and U9644 (N_9644,N_6492,N_8379);
xor U9645 (N_9645,N_7596,N_8940);
xor U9646 (N_9646,N_6864,N_6613);
nor U9647 (N_9647,N_6375,N_8792);
xor U9648 (N_9648,N_8764,N_8329);
nor U9649 (N_9649,N_8744,N_6580);
nand U9650 (N_9650,N_6930,N_7998);
nor U9651 (N_9651,N_6619,N_6451);
nand U9652 (N_9652,N_7581,N_6667);
nand U9653 (N_9653,N_6620,N_8257);
and U9654 (N_9654,N_8982,N_6247);
and U9655 (N_9655,N_7963,N_6942);
or U9656 (N_9656,N_7064,N_6378);
and U9657 (N_9657,N_7788,N_6181);
or U9658 (N_9658,N_6536,N_8438);
xor U9659 (N_9659,N_8403,N_7445);
nand U9660 (N_9660,N_7895,N_7727);
and U9661 (N_9661,N_6210,N_6507);
and U9662 (N_9662,N_8106,N_7042);
and U9663 (N_9663,N_8885,N_8645);
xor U9664 (N_9664,N_8947,N_7234);
xnor U9665 (N_9665,N_7950,N_8578);
nor U9666 (N_9666,N_7010,N_7540);
and U9667 (N_9667,N_8186,N_7086);
nor U9668 (N_9668,N_7382,N_7933);
xor U9669 (N_9669,N_7200,N_6532);
nor U9670 (N_9670,N_7623,N_6116);
nor U9671 (N_9671,N_8852,N_6636);
nor U9672 (N_9672,N_8018,N_6603);
nor U9673 (N_9673,N_8939,N_8747);
and U9674 (N_9674,N_7958,N_8898);
nand U9675 (N_9675,N_7947,N_7863);
or U9676 (N_9676,N_7223,N_7280);
or U9677 (N_9677,N_6932,N_8773);
nand U9678 (N_9678,N_7389,N_6271);
or U9679 (N_9679,N_6618,N_8768);
xor U9680 (N_9680,N_6519,N_6199);
and U9681 (N_9681,N_6152,N_8410);
xor U9682 (N_9682,N_7830,N_7579);
nand U9683 (N_9683,N_8750,N_7888);
nor U9684 (N_9684,N_7318,N_7457);
nor U9685 (N_9685,N_8905,N_7122);
xnor U9686 (N_9686,N_6403,N_6138);
xnor U9687 (N_9687,N_6289,N_6402);
or U9688 (N_9688,N_8575,N_7588);
nand U9689 (N_9689,N_7962,N_7092);
nand U9690 (N_9690,N_7146,N_6883);
or U9691 (N_9691,N_6460,N_7467);
or U9692 (N_9692,N_8560,N_8592);
xor U9693 (N_9693,N_6075,N_8544);
or U9694 (N_9694,N_7381,N_7106);
nor U9695 (N_9695,N_7583,N_7410);
xnor U9696 (N_9696,N_6976,N_7488);
nor U9697 (N_9697,N_6445,N_6165);
nor U9698 (N_9698,N_7187,N_7969);
or U9699 (N_9699,N_7137,N_7215);
or U9700 (N_9700,N_6811,N_6537);
nand U9701 (N_9701,N_8415,N_6964);
or U9702 (N_9702,N_6141,N_8171);
nand U9703 (N_9703,N_7825,N_8195);
xor U9704 (N_9704,N_6878,N_8210);
xnor U9705 (N_9705,N_6538,N_7406);
xnor U9706 (N_9706,N_8496,N_8218);
nand U9707 (N_9707,N_6329,N_8653);
xnor U9708 (N_9708,N_7369,N_8716);
or U9709 (N_9709,N_8860,N_8492);
nor U9710 (N_9710,N_8528,N_8634);
nor U9711 (N_9711,N_7885,N_7572);
nand U9712 (N_9712,N_7091,N_7766);
nor U9713 (N_9713,N_8882,N_6074);
nand U9714 (N_9714,N_7048,N_8758);
and U9715 (N_9715,N_7719,N_6544);
xor U9716 (N_9716,N_8234,N_8170);
nor U9717 (N_9717,N_8812,N_6290);
and U9718 (N_9718,N_8093,N_6904);
nand U9719 (N_9719,N_8012,N_6144);
nor U9720 (N_9720,N_8678,N_8421);
nand U9721 (N_9721,N_7396,N_8268);
nor U9722 (N_9722,N_7870,N_8840);
or U9723 (N_9723,N_8808,N_8833);
or U9724 (N_9724,N_8370,N_8846);
nor U9725 (N_9725,N_6307,N_7534);
xor U9726 (N_9726,N_8518,N_6025);
nand U9727 (N_9727,N_7019,N_7656);
or U9728 (N_9728,N_7282,N_8708);
nand U9729 (N_9729,N_6359,N_6785);
nand U9730 (N_9730,N_7826,N_8463);
and U9731 (N_9731,N_6678,N_6339);
and U9732 (N_9732,N_8143,N_7776);
or U9733 (N_9733,N_8503,N_8921);
xor U9734 (N_9734,N_6799,N_6161);
nand U9735 (N_9735,N_8406,N_6163);
xnor U9736 (N_9736,N_8696,N_8896);
nand U9737 (N_9737,N_6984,N_8057);
nor U9738 (N_9738,N_6867,N_8129);
nand U9739 (N_9739,N_6851,N_8391);
nand U9740 (N_9740,N_7101,N_6513);
nand U9741 (N_9741,N_6994,N_6317);
nor U9742 (N_9742,N_8633,N_8894);
xor U9743 (N_9743,N_7748,N_6458);
or U9744 (N_9744,N_6305,N_7872);
and U9745 (N_9745,N_6396,N_7667);
xor U9746 (N_9746,N_6083,N_7674);
nand U9747 (N_9747,N_7210,N_7750);
and U9748 (N_9748,N_8904,N_6578);
xnor U9749 (N_9749,N_7212,N_7474);
and U9750 (N_9750,N_7874,N_7817);
or U9751 (N_9751,N_8553,N_7495);
and U9752 (N_9752,N_7856,N_8239);
nor U9753 (N_9753,N_7336,N_7198);
and U9754 (N_9754,N_8670,N_6803);
nor U9755 (N_9755,N_6671,N_6086);
nand U9756 (N_9756,N_7806,N_7306);
and U9757 (N_9757,N_7576,N_7298);
nand U9758 (N_9758,N_6521,N_6233);
nand U9759 (N_9759,N_7454,N_6608);
xor U9760 (N_9760,N_8430,N_6103);
xnor U9761 (N_9761,N_6098,N_6291);
nor U9762 (N_9762,N_7841,N_7050);
and U9763 (N_9763,N_6035,N_8219);
and U9764 (N_9764,N_7819,N_6633);
and U9765 (N_9765,N_6963,N_8001);
and U9766 (N_9766,N_6635,N_7211);
xnor U9767 (N_9767,N_7352,N_8702);
nor U9768 (N_9768,N_7744,N_8930);
nor U9769 (N_9769,N_7607,N_6159);
xnor U9770 (N_9770,N_8393,N_8774);
xor U9771 (N_9771,N_7481,N_6482);
or U9772 (N_9772,N_6304,N_8296);
nor U9773 (N_9773,N_8381,N_8607);
nand U9774 (N_9774,N_7000,N_7319);
or U9775 (N_9775,N_8110,N_8946);
and U9776 (N_9776,N_8927,N_6360);
nand U9777 (N_9777,N_8596,N_6078);
and U9778 (N_9778,N_7175,N_7669);
nand U9779 (N_9779,N_8551,N_6767);
nand U9780 (N_9780,N_8577,N_6562);
xnor U9781 (N_9781,N_6447,N_8209);
nor U9782 (N_9782,N_7858,N_8601);
and U9783 (N_9783,N_6801,N_6938);
or U9784 (N_9784,N_7021,N_7511);
or U9785 (N_9785,N_6751,N_8278);
nor U9786 (N_9786,N_7403,N_8687);
nor U9787 (N_9787,N_8509,N_7346);
xor U9788 (N_9788,N_6410,N_8137);
xnor U9789 (N_9789,N_8081,N_8192);
or U9790 (N_9790,N_8074,N_6496);
nor U9791 (N_9791,N_7594,N_6975);
nand U9792 (N_9792,N_7599,N_6196);
nor U9793 (N_9793,N_8333,N_6696);
or U9794 (N_9794,N_7399,N_7723);
or U9795 (N_9795,N_6170,N_7939);
nand U9796 (N_9796,N_8311,N_6740);
xor U9797 (N_9797,N_6829,N_7251);
xnor U9798 (N_9798,N_8971,N_8548);
and U9799 (N_9799,N_8042,N_6160);
xor U9800 (N_9800,N_6676,N_7240);
and U9801 (N_9801,N_8009,N_8091);
nor U9802 (N_9802,N_8724,N_8902);
xnor U9803 (N_9803,N_8398,N_7499);
and U9804 (N_9804,N_6422,N_6885);
and U9805 (N_9805,N_8056,N_7898);
or U9806 (N_9806,N_8007,N_8689);
xor U9807 (N_9807,N_6755,N_6175);
and U9808 (N_9808,N_6348,N_8429);
nor U9809 (N_9809,N_7508,N_7165);
nor U9810 (N_9810,N_8574,N_8817);
and U9811 (N_9811,N_6509,N_6071);
nor U9812 (N_9812,N_6866,N_8263);
and U9813 (N_9813,N_6982,N_6865);
xor U9814 (N_9814,N_6188,N_7768);
or U9815 (N_9815,N_7739,N_7827);
nor U9816 (N_9816,N_8280,N_6148);
and U9817 (N_9817,N_6018,N_7094);
nor U9818 (N_9818,N_6063,N_8642);
nand U9819 (N_9819,N_6945,N_7566);
or U9820 (N_9820,N_8275,N_8981);
and U9821 (N_9821,N_7526,N_8248);
nand U9822 (N_9822,N_6173,N_6494);
xnor U9823 (N_9823,N_8139,N_8651);
and U9824 (N_9824,N_7110,N_6912);
nor U9825 (N_9825,N_7763,N_6203);
and U9826 (N_9826,N_8150,N_8665);
or U9827 (N_9827,N_7593,N_6288);
and U9828 (N_9828,N_8467,N_6737);
nand U9829 (N_9829,N_8488,N_6373);
nand U9830 (N_9830,N_8063,N_8441);
nand U9831 (N_9831,N_8458,N_6789);
nor U9832 (N_9832,N_6051,N_7287);
xnor U9833 (N_9833,N_8207,N_6372);
nor U9834 (N_9834,N_8738,N_6614);
nor U9835 (N_9835,N_7967,N_6484);
nand U9836 (N_9836,N_6909,N_7957);
nand U9837 (N_9837,N_6587,N_7516);
nand U9838 (N_9838,N_8371,N_8397);
xnor U9839 (N_9839,N_6990,N_8125);
and U9840 (N_9840,N_7204,N_7281);
xnor U9841 (N_9841,N_8783,N_7479);
nand U9842 (N_9842,N_8922,N_6448);
or U9843 (N_9843,N_6539,N_6224);
nand U9844 (N_9844,N_6850,N_7265);
nand U9845 (N_9845,N_6479,N_6848);
nand U9846 (N_9846,N_7647,N_7153);
nor U9847 (N_9847,N_8206,N_6186);
and U9848 (N_9848,N_6680,N_8674);
nor U9849 (N_9849,N_7638,N_7244);
nand U9850 (N_9850,N_8590,N_8748);
nor U9851 (N_9851,N_8092,N_7228);
nor U9852 (N_9852,N_7781,N_7801);
nand U9853 (N_9853,N_8017,N_6661);
and U9854 (N_9854,N_6596,N_8058);
nor U9855 (N_9855,N_8022,N_6383);
xnor U9856 (N_9856,N_8964,N_6584);
xor U9857 (N_9857,N_7756,N_8082);
xnor U9858 (N_9858,N_6868,N_6897);
or U9859 (N_9859,N_7338,N_7809);
nand U9860 (N_9860,N_7354,N_8836);
nand U9861 (N_9861,N_6830,N_6418);
nor U9862 (N_9862,N_6876,N_8962);
nand U9863 (N_9863,N_8561,N_8160);
nand U9864 (N_9864,N_8470,N_7828);
and U9865 (N_9865,N_6997,N_8162);
nand U9866 (N_9866,N_7264,N_8632);
or U9867 (N_9867,N_8533,N_8168);
and U9868 (N_9868,N_7818,N_6498);
and U9869 (N_9869,N_7272,N_7077);
or U9870 (N_9870,N_8652,N_7057);
or U9871 (N_9871,N_8041,N_8424);
nor U9872 (N_9872,N_8369,N_6993);
and U9873 (N_9873,N_8076,N_6583);
nand U9874 (N_9874,N_8295,N_7838);
or U9875 (N_9875,N_8919,N_7979);
nand U9876 (N_9876,N_8355,N_6653);
and U9877 (N_9877,N_8507,N_8315);
xor U9878 (N_9878,N_6922,N_7676);
and U9879 (N_9879,N_6286,N_8029);
or U9880 (N_9880,N_8770,N_6753);
and U9881 (N_9881,N_6549,N_8427);
or U9882 (N_9882,N_8815,N_7063);
and U9883 (N_9883,N_6669,N_7678);
nor U9884 (N_9884,N_7755,N_7589);
nor U9885 (N_9885,N_6981,N_8049);
nor U9886 (N_9886,N_7661,N_6704);
xor U9887 (N_9887,N_6791,N_6884);
xnor U9888 (N_9888,N_7604,N_7840);
and U9889 (N_9889,N_8857,N_8337);
xor U9890 (N_9890,N_7415,N_6872);
nand U9891 (N_9891,N_8099,N_7641);
or U9892 (N_9892,N_7031,N_7938);
nor U9893 (N_9893,N_8915,N_6341);
xor U9894 (N_9894,N_6543,N_8439);
and U9895 (N_9895,N_6590,N_7713);
and U9896 (N_9896,N_7493,N_7759);
nand U9897 (N_9897,N_6315,N_8431);
xor U9898 (N_9898,N_8672,N_8705);
nor U9899 (N_9899,N_6853,N_8581);
nor U9900 (N_9900,N_8869,N_6316);
xnor U9901 (N_9901,N_7390,N_6124);
nor U9902 (N_9902,N_8289,N_8763);
nand U9903 (N_9903,N_8521,N_7330);
xnor U9904 (N_9904,N_8959,N_8212);
xor U9905 (N_9905,N_8034,N_8511);
nand U9906 (N_9906,N_8362,N_8938);
xnor U9907 (N_9907,N_8660,N_8802);
nand U9908 (N_9908,N_8979,N_6043);
xor U9909 (N_9909,N_6352,N_7328);
or U9910 (N_9910,N_6272,N_7761);
xor U9911 (N_9911,N_7132,N_6727);
nor U9912 (N_9912,N_7543,N_6835);
and U9913 (N_9913,N_8510,N_8221);
or U9914 (N_9914,N_8757,N_7811);
xnor U9915 (N_9915,N_8884,N_8344);
nor U9916 (N_9916,N_6717,N_7714);
or U9917 (N_9917,N_6431,N_8671);
and U9918 (N_9918,N_7574,N_6595);
and U9919 (N_9919,N_7558,N_6725);
nand U9920 (N_9920,N_6466,N_6133);
or U9921 (N_9921,N_6195,N_6711);
and U9922 (N_9922,N_6654,N_6805);
xnor U9923 (N_9923,N_7335,N_6934);
and U9924 (N_9924,N_8199,N_8304);
nand U9925 (N_9925,N_7903,N_7608);
or U9926 (N_9926,N_7715,N_6292);
nor U9927 (N_9927,N_8088,N_6366);
or U9928 (N_9928,N_6902,N_8754);
or U9929 (N_9929,N_6586,N_7007);
or U9930 (N_9930,N_7085,N_6675);
and U9931 (N_9931,N_8228,N_8549);
or U9932 (N_9932,N_6076,N_6031);
nor U9933 (N_9933,N_8435,N_7288);
or U9934 (N_9934,N_6616,N_7144);
xnor U9935 (N_9935,N_6463,N_7423);
xnor U9936 (N_9936,N_7373,N_7357);
xnor U9937 (N_9937,N_7289,N_8730);
nand U9938 (N_9938,N_7119,N_8917);
nand U9939 (N_9939,N_7285,N_8173);
nor U9940 (N_9940,N_7535,N_8030);
or U9941 (N_9941,N_7891,N_6780);
nand U9942 (N_9942,N_7436,N_6606);
and U9943 (N_9943,N_8684,N_7099);
or U9944 (N_9944,N_6122,N_7076);
nand U9945 (N_9945,N_8803,N_8782);
nand U9946 (N_9946,N_7605,N_8215);
nand U9947 (N_9947,N_6534,N_6528);
and U9948 (N_9948,N_8820,N_6746);
nor U9949 (N_9949,N_6461,N_7471);
xnor U9950 (N_9950,N_7650,N_8051);
nor U9951 (N_9951,N_7916,N_7218);
nor U9952 (N_9952,N_7961,N_6906);
nand U9953 (N_9953,N_7329,N_7670);
nand U9954 (N_9954,N_6924,N_7345);
nor U9955 (N_9955,N_8546,N_8788);
nand U9956 (N_9956,N_6724,N_6381);
or U9957 (N_9957,N_8350,N_8495);
xor U9958 (N_9958,N_8013,N_7735);
nand U9959 (N_9959,N_7188,N_7613);
xor U9960 (N_9960,N_7360,N_6268);
xnor U9961 (N_9961,N_7468,N_7216);
xnor U9962 (N_9962,N_7103,N_7309);
or U9963 (N_9963,N_6687,N_7627);
nand U9964 (N_9964,N_8677,N_7660);
xnor U9965 (N_9965,N_7387,N_7546);
and U9966 (N_9966,N_7548,N_8994);
nor U9967 (N_9967,N_8480,N_7956);
and U9968 (N_9968,N_6354,N_7065);
and U9969 (N_9969,N_7677,N_8077);
nor U9970 (N_9970,N_8612,N_6508);
nor U9971 (N_9971,N_8655,N_7420);
xor U9972 (N_9972,N_7351,N_7183);
nor U9973 (N_9973,N_7592,N_7665);
or U9974 (N_9974,N_7332,N_7679);
or U9975 (N_9975,N_8555,N_7866);
nor U9976 (N_9976,N_8892,N_6242);
nand U9977 (N_9977,N_7376,N_6264);
nor U9978 (N_9978,N_8457,N_7202);
or U9979 (N_9979,N_8639,N_6747);
xnor U9980 (N_9980,N_8196,N_8198);
or U9981 (N_9981,N_7906,N_7224);
and U9982 (N_9982,N_8357,N_6783);
nor U9983 (N_9983,N_8862,N_6481);
xor U9984 (N_9984,N_8975,N_6954);
and U9985 (N_9985,N_6726,N_8128);
or U9986 (N_9986,N_6273,N_8187);
and U9987 (N_9987,N_7178,N_7446);
and U9988 (N_9988,N_8867,N_7964);
nor U9989 (N_9989,N_6637,N_7810);
xor U9990 (N_9990,N_6563,N_6861);
nand U9991 (N_9991,N_7393,N_6176);
nand U9992 (N_9992,N_6891,N_7109);
nand U9993 (N_9993,N_6400,N_6092);
nor U9994 (N_9994,N_6657,N_7062);
nor U9995 (N_9995,N_6523,N_6005);
and U9996 (N_9996,N_8388,N_7427);
and U9997 (N_9997,N_6731,N_6750);
and U9998 (N_9998,N_6822,N_8200);
nor U9999 (N_9999,N_8339,N_8740);
nand U10000 (N_10000,N_6545,N_7896);
nand U10001 (N_10001,N_8843,N_6284);
nand U10002 (N_10002,N_7088,N_7238);
nand U10003 (N_10003,N_6665,N_8825);
and U10004 (N_10004,N_7459,N_8464);
nand U10005 (N_10005,N_6162,N_6722);
xor U10006 (N_10006,N_8015,N_8954);
xnor U10007 (N_10007,N_7221,N_7846);
nand U10008 (N_10008,N_8178,N_7551);
nand U10009 (N_10009,N_6575,N_8094);
nand U10010 (N_10010,N_6434,N_8332);
nand U10011 (N_10011,N_8368,N_6923);
xor U10012 (N_10012,N_7780,N_6921);
nor U10013 (N_10013,N_8627,N_6424);
or U10014 (N_10014,N_6996,N_8849);
xnor U10015 (N_10015,N_7894,N_6298);
and U10016 (N_10016,N_8931,N_6743);
nor U10017 (N_10017,N_6253,N_6475);
and U10018 (N_10018,N_6037,N_6322);
or U10019 (N_10019,N_8396,N_8378);
xnor U10020 (N_10020,N_7920,N_8308);
nor U10021 (N_10021,N_8401,N_8834);
nor U10022 (N_10022,N_6547,N_8416);
xnor U10023 (N_10023,N_8842,N_7135);
nand U10024 (N_10024,N_7283,N_6824);
xnor U10025 (N_10025,N_6034,N_7730);
nor U10026 (N_10026,N_7839,N_7286);
nor U10027 (N_10027,N_7709,N_6406);
or U10028 (N_10028,N_8321,N_7675);
xnor U10029 (N_10029,N_7926,N_7098);
or U10030 (N_10030,N_7760,N_8265);
or U10031 (N_10031,N_6629,N_8576);
nor U10032 (N_10032,N_6060,N_6579);
and U10033 (N_10033,N_7043,N_6591);
nand U10034 (N_10034,N_7008,N_8822);
or U10035 (N_10035,N_8776,N_8272);
xor U10036 (N_10036,N_7582,N_8547);
or U10037 (N_10037,N_6004,N_8227);
nor U10038 (N_10038,N_7837,N_8571);
xnor U10039 (N_10039,N_8806,N_8167);
xor U10040 (N_10040,N_6283,N_8694);
xnor U10041 (N_10041,N_7659,N_8202);
or U10042 (N_10042,N_8630,N_8877);
and U10043 (N_10043,N_8028,N_8668);
nand U10044 (N_10044,N_8937,N_6859);
xor U10045 (N_10045,N_8229,N_7363);
and U10046 (N_10046,N_7943,N_7695);
or U10047 (N_10047,N_7785,N_8565);
and U10048 (N_10048,N_8829,N_8923);
and U10049 (N_10049,N_6251,N_6313);
nor U10050 (N_10050,N_6119,N_7791);
and U10051 (N_10051,N_6771,N_8720);
and U10052 (N_10052,N_6046,N_6321);
or U10053 (N_10053,N_7985,N_7506);
nand U10054 (N_10054,N_7434,N_8999);
or U10055 (N_10055,N_7591,N_6435);
nor U10056 (N_10056,N_7845,N_6625);
or U10057 (N_10057,N_8070,N_8223);
and U10058 (N_10058,N_8780,N_6561);
or U10059 (N_10059,N_8895,N_8147);
and U10060 (N_10060,N_6839,N_6841);
nand U10061 (N_10061,N_8873,N_8879);
nand U10062 (N_10062,N_6282,N_6363);
and U10063 (N_10063,N_8957,N_6697);
or U10064 (N_10064,N_8142,N_7342);
xnor U10065 (N_10065,N_8654,N_8481);
nand U10066 (N_10066,N_6347,N_7161);
xor U10067 (N_10067,N_6377,N_8791);
nand U10068 (N_10068,N_8823,N_7868);
nor U10069 (N_10069,N_6442,N_8686);
and U10070 (N_10070,N_6470,N_6768);
nand U10071 (N_10071,N_6953,N_6285);
nor U10072 (N_10072,N_8374,N_8990);
and U10073 (N_10073,N_8926,N_7191);
nand U10074 (N_10074,N_8418,N_7174);
nor U10075 (N_10075,N_7977,N_7882);
nor U10076 (N_10076,N_6096,N_6929);
and U10077 (N_10077,N_8650,N_7569);
and U10078 (N_10078,N_7816,N_7276);
nand U10079 (N_10079,N_6522,N_7172);
xor U10080 (N_10080,N_6749,N_8299);
nand U10081 (N_10081,N_7712,N_7625);
xor U10082 (N_10082,N_6741,N_7747);
nor U10083 (N_10083,N_8893,N_6821);
xor U10084 (N_10084,N_6252,N_7271);
nand U10085 (N_10085,N_8729,N_7038);
or U10086 (N_10086,N_6796,N_7054);
nor U10087 (N_10087,N_6266,N_8114);
and U10088 (N_10088,N_6107,N_6277);
nor U10089 (N_10089,N_7897,N_7847);
or U10090 (N_10090,N_6832,N_6871);
xnor U10091 (N_10091,N_7921,N_8033);
nor U10092 (N_10092,N_6988,N_7671);
nand U10093 (N_10093,N_6535,N_8855);
and U10094 (N_10094,N_6079,N_7378);
and U10095 (N_10095,N_6149,N_6927);
nand U10096 (N_10096,N_7162,N_8249);
nor U10097 (N_10097,N_7726,N_6598);
and U10098 (N_10098,N_8501,N_6985);
nor U10099 (N_10099,N_8933,N_7475);
nor U10100 (N_10100,N_6529,N_7484);
and U10101 (N_10101,N_8444,N_8620);
or U10102 (N_10102,N_6419,N_7762);
and U10103 (N_10103,N_8021,N_8352);
nor U10104 (N_10104,N_7666,N_8120);
nor U10105 (N_10105,N_7029,N_8897);
nand U10106 (N_10106,N_8539,N_6085);
or U10107 (N_10107,N_6108,N_8569);
and U10108 (N_10108,N_8883,N_8681);
xor U10109 (N_10109,N_6082,N_7624);
or U10110 (N_10110,N_6957,N_6983);
nand U10111 (N_10111,N_6179,N_6663);
nand U10112 (N_10112,N_7313,N_7422);
xor U10113 (N_10113,N_6414,N_8356);
and U10114 (N_10114,N_7952,N_8360);
nand U10115 (N_10115,N_6760,N_6006);
nor U10116 (N_10116,N_8353,N_7795);
nor U10117 (N_10117,N_8613,N_7884);
nor U10118 (N_10118,N_7401,N_6411);
xnor U10119 (N_10119,N_6237,N_6404);
nor U10120 (N_10120,N_7073,N_8527);
and U10121 (N_10121,N_6914,N_7486);
nor U10122 (N_10122,N_6858,N_8244);
nor U10123 (N_10123,N_6000,N_8060);
nand U10124 (N_10124,N_6353,N_7340);
and U10125 (N_10125,N_6072,N_6095);
or U10126 (N_10126,N_6384,N_6888);
xor U10127 (N_10127,N_6250,N_6155);
nand U10128 (N_10128,N_7587,N_8475);
and U10129 (N_10129,N_6518,N_8290);
and U10130 (N_10130,N_6838,N_8969);
nor U10131 (N_10131,N_8717,N_7219);
xor U10132 (N_10132,N_6901,N_8462);
nor U10133 (N_10133,N_7704,N_8967);
xor U10134 (N_10134,N_8423,N_8133);
and U10135 (N_10135,N_7590,N_6649);
xnor U10136 (N_10136,N_7268,N_6061);
nand U10137 (N_10137,N_8460,N_6226);
and U10138 (N_10138,N_7025,N_7075);
xnor U10139 (N_10139,N_6355,N_6828);
xor U10140 (N_10140,N_8297,N_6328);
and U10141 (N_10141,N_6314,N_8543);
nand U10142 (N_10142,N_6147,N_8845);
and U10143 (N_10143,N_8205,N_6045);
and U10144 (N_10144,N_8706,N_6723);
or U10145 (N_10145,N_6297,N_6389);
xnor U10146 (N_10146,N_7890,N_8832);
or U10147 (N_10147,N_6825,N_6926);
nand U10148 (N_10148,N_7315,N_8850);
nor U10149 (N_10149,N_6333,N_7004);
nand U10150 (N_10150,N_7131,N_7125);
or U10151 (N_10151,N_6327,N_7291);
nor U10152 (N_10152,N_6843,N_7252);
or U10153 (N_10153,N_7778,N_8420);
xor U10154 (N_10154,N_8700,N_7497);
and U10155 (N_10155,N_6552,N_7549);
and U10156 (N_10156,N_6516,N_8625);
nand U10157 (N_10157,N_6436,N_8830);
nor U10158 (N_10158,N_6462,N_8347);
or U10159 (N_10159,N_7377,N_8131);
xor U10160 (N_10160,N_7262,N_7749);
nor U10161 (N_10161,N_6736,N_7456);
or U10162 (N_10162,N_7787,N_6903);
or U10163 (N_10163,N_8376,N_7418);
xnor U10164 (N_10164,N_8055,N_7412);
and U10165 (N_10165,N_8113,N_7519);
and U10166 (N_10166,N_6813,N_6387);
and U10167 (N_10167,N_6185,N_7707);
xor U10168 (N_10168,N_8997,N_6764);
and U10169 (N_10169,N_8083,N_8761);
nor U10170 (N_10170,N_7578,N_7450);
xnor U10171 (N_10171,N_6301,N_6597);
nand U10172 (N_10172,N_8531,N_6819);
nand U10173 (N_10173,N_6860,N_8722);
or U10174 (N_10174,N_8657,N_8636);
nor U10175 (N_10175,N_8864,N_8968);
or U10176 (N_10176,N_8181,N_8134);
nor U10177 (N_10177,N_7733,N_6394);
or U10178 (N_10178,N_8006,N_8255);
and U10179 (N_10179,N_6782,N_8466);
or U10180 (N_10180,N_6190,N_7388);
nor U10181 (N_10181,N_7374,N_8301);
xor U10182 (N_10182,N_7069,N_8564);
xor U10183 (N_10183,N_7322,N_6030);
or U10184 (N_10184,N_6346,N_6440);
nor U10185 (N_10185,N_8958,N_8433);
and U10186 (N_10186,N_7550,N_8111);
nor U10187 (N_10187,N_8646,N_8087);
nor U10188 (N_10188,N_7693,N_7565);
or U10189 (N_10189,N_7522,N_6939);
nor U10190 (N_10190,N_8513,N_7358);
and U10191 (N_10191,N_6099,N_7156);
and U10192 (N_10192,N_8732,N_6570);
xnor U10193 (N_10193,N_6572,N_7230);
and U10194 (N_10194,N_8456,N_8713);
or U10195 (N_10195,N_8314,N_6218);
and U10196 (N_10196,N_7150,N_8064);
nor U10197 (N_10197,N_7633,N_6480);
nand U10198 (N_10198,N_7990,N_6573);
nor U10199 (N_10199,N_7115,N_7082);
nor U10200 (N_10200,N_8490,N_8451);
and U10201 (N_10201,N_7804,N_6308);
xor U10202 (N_10202,N_7865,N_7449);
xnor U10203 (N_10203,N_8530,N_7492);
nor U10204 (N_10204,N_7658,N_8907);
and U10205 (N_10205,N_8224,N_7487);
nand U10206 (N_10206,N_6362,N_8586);
xnor U10207 (N_10207,N_6081,N_6349);
nor U10208 (N_10208,N_8238,N_6955);
and U10209 (N_10209,N_8317,N_8878);
xor U10210 (N_10210,N_6444,N_7233);
and U10211 (N_10211,N_8988,N_6766);
xor U10212 (N_10212,N_6745,N_8189);
or U10213 (N_10213,N_7790,N_7305);
xnor U10214 (N_10214,N_7001,N_8520);
xnor U10215 (N_10215,N_6730,N_7717);
nor U10216 (N_10216,N_6617,N_8735);
nor U10217 (N_10217,N_8659,N_6239);
nor U10218 (N_10218,N_8676,N_6293);
nor U10219 (N_10219,N_7934,N_6477);
nor U10220 (N_10220,N_7532,N_8573);
nand U10221 (N_10221,N_7871,N_7794);
nand U10222 (N_10222,N_6594,N_8733);
nor U10223 (N_10223,N_7767,N_6499);
nand U10224 (N_10224,N_7051,N_8449);
nand U10225 (N_10225,N_8529,N_6664);
or U10226 (N_10226,N_7370,N_7595);
xor U10227 (N_10227,N_7185,N_8158);
nand U10228 (N_10228,N_6267,N_7554);
or U10229 (N_10229,N_8600,N_6438);
nor U10230 (N_10230,N_6812,N_7529);
xor U10231 (N_10231,N_8443,N_7301);
nand U10232 (N_10232,N_8476,N_7052);
xnor U10233 (N_10233,N_7448,N_6102);
and U10234 (N_10234,N_7194,N_8874);
nor U10235 (N_10235,N_8277,N_7648);
nand U10236 (N_10236,N_6648,N_7359);
or U10237 (N_10237,N_7862,N_8910);
and U10238 (N_10238,N_8169,N_6413);
nor U10239 (N_10239,N_7030,N_6920);
or U10240 (N_10240,N_7536,N_6973);
xnor U10241 (N_10241,N_7988,N_7337);
and U10242 (N_10242,N_8161,N_6409);
nor U10243 (N_10243,N_7070,N_8584);
xnor U10244 (N_10244,N_8597,N_8100);
or U10245 (N_10245,N_8570,N_8769);
nor U10246 (N_10246,N_6408,N_7682);
nor U10247 (N_10247,N_8589,N_7935);
and U10248 (N_10248,N_8554,N_7980);
and U10249 (N_10249,N_8622,N_8258);
nor U10250 (N_10250,N_6337,N_8354);
nor U10251 (N_10251,N_8929,N_7716);
nor U10252 (N_10252,N_8175,N_8452);
and U10253 (N_10253,N_6336,N_6936);
xnor U10254 (N_10254,N_6191,N_8745);
or U10255 (N_10255,N_7044,N_8805);
or U10256 (N_10256,N_8071,N_6702);
nor U10257 (N_10257,N_7699,N_8148);
nand U10258 (N_10258,N_6343,N_6212);
nand U10259 (N_10259,N_8667,N_7353);
or U10260 (N_10260,N_7821,N_7179);
and U10261 (N_10261,N_7833,N_7490);
nor U10262 (N_10262,N_6241,N_6542);
and U10263 (N_10263,N_7124,N_8232);
or U10264 (N_10264,N_6941,N_7327);
and U10265 (N_10265,N_8629,N_7524);
and U10266 (N_10266,N_8361,N_8866);
nor U10267 (N_10267,N_7843,N_7878);
or U10268 (N_10268,N_6967,N_6666);
and U10269 (N_10269,N_6053,N_8032);
nor U10270 (N_10270,N_7407,N_8675);
or U10271 (N_10271,N_7651,N_7919);
nand U10272 (N_10272,N_6278,N_7611);
or U10273 (N_10273,N_7626,N_8149);
or U10274 (N_10274,N_7684,N_6157);
or U10275 (N_10275,N_6009,N_8335);
nor U10276 (N_10276,N_8358,N_6156);
nand U10277 (N_10277,N_7725,N_8240);
or U10278 (N_10278,N_7107,N_6036);
xnor U10279 (N_10279,N_6778,N_8326);
and U10280 (N_10280,N_6332,N_6211);
xnor U10281 (N_10281,N_7164,N_8008);
and U10282 (N_10282,N_7805,N_7207);
xor U10283 (N_10283,N_7443,N_8217);
and U10284 (N_10284,N_6207,N_8550);
nor U10285 (N_10285,N_7968,N_6497);
nand U10286 (N_10286,N_8844,N_6972);
nor U10287 (N_10287,N_6449,N_6145);
xor U10288 (N_10288,N_6530,N_7984);
and U10289 (N_10289,N_6833,N_8123);
xor U10290 (N_10290,N_6177,N_8096);
nor U10291 (N_10291,N_6486,N_7688);
or U10292 (N_10292,N_6643,N_6245);
nand U10293 (N_10293,N_6855,N_7743);
and U10294 (N_10294,N_8281,N_8144);
nor U10295 (N_10295,N_8648,N_6775);
nand U10296 (N_10296,N_8455,N_7206);
xor U10297 (N_10297,N_6457,N_8635);
or U10298 (N_10298,N_8587,N_8163);
and U10299 (N_10299,N_6748,N_6048);
or U10300 (N_10300,N_7697,N_7945);
nor U10301 (N_10301,N_6754,N_8688);
and U10302 (N_10302,N_6143,N_6559);
and U10303 (N_10303,N_7058,N_8216);
or U10304 (N_10304,N_8115,N_7836);
nand U10305 (N_10305,N_8386,N_8881);
nand U10306 (N_10306,N_8107,N_7802);
or U10307 (N_10307,N_6395,N_7242);
nand U10308 (N_10308,N_7855,N_7867);
or U10309 (N_10309,N_7398,N_8026);
nor U10310 (N_10310,N_6794,N_7176);
and U10311 (N_10311,N_7765,N_7463);
xnor U10312 (N_10312,N_8712,N_6810);
nand U10313 (N_10313,N_6187,N_6416);
or U10314 (N_10314,N_8254,N_7899);
or U10315 (N_10315,N_6279,N_7924);
and U10316 (N_10316,N_8318,N_6911);
or U10317 (N_10317,N_7243,N_8995);
and U10318 (N_10318,N_8177,N_6488);
and U10319 (N_10319,N_7989,N_7777);
nand U10320 (N_10320,N_8291,N_6126);
xor U10321 (N_10321,N_7718,N_6978);
nor U10322 (N_10322,N_6991,N_7333);
or U10323 (N_10323,N_6476,N_7405);
nand U10324 (N_10324,N_6788,N_6772);
xor U10325 (N_10325,N_7706,N_7375);
nand U10326 (N_10326,N_6033,N_6732);
and U10327 (N_10327,N_6093,N_8453);
nand U10328 (N_10328,N_6050,N_8343);
or U10329 (N_10329,N_8471,N_8121);
nand U10330 (N_10330,N_6493,N_8536);
xor U10331 (N_10331,N_6681,N_8151);
and U10332 (N_10332,N_7722,N_7128);
nor U10333 (N_10333,N_8762,N_6432);
nand U10334 (N_10334,N_6169,N_6548);
and U10335 (N_10335,N_8419,N_6795);
or U10336 (N_10336,N_7970,N_7792);
nor U10337 (N_10337,N_6026,N_6139);
or U10338 (N_10338,N_7705,N_7562);
or U10339 (N_10339,N_8787,N_7779);
nor U10340 (N_10340,N_6514,N_6390);
nand U10341 (N_10341,N_7799,N_7687);
xor U10342 (N_10342,N_6140,N_7556);
nor U10343 (N_10343,N_7173,N_6714);
or U10344 (N_10344,N_8960,N_7515);
or U10345 (N_10345,N_6599,N_6773);
nand U10346 (N_10346,N_6125,N_8709);
and U10347 (N_10347,N_6847,N_6171);
or U10348 (N_10348,N_6429,N_6310);
nor U10349 (N_10349,N_7034,N_6294);
nand U10350 (N_10350,N_8617,N_8267);
nand U10351 (N_10351,N_6335,N_7372);
nor U10352 (N_10352,N_6842,N_6679);
nor U10353 (N_10353,N_7521,N_7598);
nand U10354 (N_10354,N_6919,N_7708);
nand U10355 (N_10355,N_7068,N_6130);
nor U10356 (N_10356,N_8579,N_7646);
and U10357 (N_10357,N_6873,N_8970);
nand U10358 (N_10358,N_7326,N_6966);
nor U10359 (N_10359,N_8390,N_7996);
nand U10360 (N_10360,N_7973,N_8861);
nand U10361 (N_10361,N_7011,N_6793);
or U10362 (N_10362,N_7922,N_8035);
xnor U10363 (N_10363,N_7111,N_6427);
or U10364 (N_10364,N_6540,N_8068);
nor U10365 (N_10365,N_6569,N_7559);
nor U10366 (N_10366,N_8523,N_7299);
nand U10367 (N_10367,N_8835,N_8109);
nand U10368 (N_10368,N_8146,N_6197);
nor U10369 (N_10369,N_8786,N_8572);
or U10370 (N_10370,N_8497,N_6311);
or U10371 (N_10371,N_7909,N_6950);
and U10372 (N_10372,N_8963,N_6689);
nor U10373 (N_10373,N_7585,N_8965);
nor U10374 (N_10374,N_8986,N_7201);
nand U10375 (N_10375,N_7294,N_6229);
and U10376 (N_10376,N_6807,N_7430);
nor U10377 (N_10377,N_7772,N_8130);
nand U10378 (N_10378,N_7949,N_7505);
nor U10379 (N_10379,N_6893,N_6265);
or U10380 (N_10380,N_6105,N_6016);
xnor U10381 (N_10381,N_7736,N_6490);
xor U10382 (N_10382,N_8102,N_7429);
and U10383 (N_10383,N_6610,N_7141);
nand U10384 (N_10384,N_6774,N_6365);
nor U10385 (N_10385,N_7494,N_8664);
xnor U10386 (N_10386,N_8065,N_7196);
xnor U10387 (N_10387,N_6204,N_8588);
nand U10388 (N_10388,N_8442,N_8585);
and U10389 (N_10389,N_6219,N_7918);
nor U10390 (N_10390,N_6198,N_7386);
nor U10391 (N_10391,N_6441,N_8197);
nand U10392 (N_10392,N_8638,N_6227);
nand U10393 (N_10393,N_8484,N_8078);
or U10394 (N_10394,N_6781,N_8941);
nor U10395 (N_10395,N_7006,N_6895);
and U10396 (N_10396,N_7999,N_7116);
nand U10397 (N_10397,N_8743,N_8084);
and U10398 (N_10398,N_7171,N_7253);
xnor U10399 (N_10399,N_8220,N_6658);
nand U10400 (N_10400,N_6013,N_7321);
and U10401 (N_10401,N_7250,N_6739);
xnor U10402 (N_10402,N_8602,N_6958);
or U10403 (N_10403,N_6243,N_8691);
and U10404 (N_10404,N_6719,N_8853);
or U10405 (N_10405,N_6118,N_8603);
nor U10406 (N_10406,N_7774,N_6077);
or U10407 (N_10407,N_6192,N_6645);
xor U10408 (N_10408,N_7290,N_8384);
and U10409 (N_10409,N_8334,N_7510);
nand U10410 (N_10410,N_6350,N_7248);
and U10411 (N_10411,N_6688,N_7789);
xor U10412 (N_10412,N_6209,N_6965);
and U10413 (N_10413,N_8526,N_6900);
and U10414 (N_10414,N_6673,N_8683);
xor U10415 (N_10415,N_6784,N_7773);
xor U10416 (N_10416,N_6879,N_8610);
xor U10417 (N_10417,N_7003,N_7829);
nor U10418 (N_10418,N_7634,N_6109);
xnor U10419 (N_10419,N_7296,N_8838);
or U10420 (N_10420,N_8859,N_6153);
and U10421 (N_10421,N_7832,N_8619);
xor U10422 (N_10422,N_8766,N_6439);
nor U10423 (N_10423,N_7455,N_7971);
or U10424 (N_10424,N_6055,N_7995);
and U10425 (N_10425,N_6656,N_7214);
nand U10426 (N_10426,N_8831,N_7831);
xor U10427 (N_10427,N_6367,N_8516);
nand U10428 (N_10428,N_8473,N_6296);
and U10429 (N_10429,N_8525,N_8324);
xnor U10430 (N_10430,N_7361,N_8305);
or U10431 (N_10431,N_7269,N_6386);
and U10432 (N_10432,N_6002,N_6898);
nor U10433 (N_10433,N_6524,N_6836);
nor U10434 (N_10434,N_7278,N_7205);
nor U10435 (N_10435,N_6531,N_6097);
or U10436 (N_10436,N_7600,N_6639);
nor U10437 (N_10437,N_6228,N_7035);
nand U10438 (N_10438,N_8514,N_7978);
nor U10439 (N_10439,N_6027,N_7055);
nor U10440 (N_10440,N_7411,N_8323);
and U10441 (N_10441,N_7610,N_6607);
xnor U10442 (N_10442,N_8002,N_6407);
or U10443 (N_10443,N_7047,N_8000);
xor U10444 (N_10444,N_6338,N_6421);
nor U10445 (N_10445,N_8680,N_7067);
nor U10446 (N_10446,N_8247,N_8288);
or U10447 (N_10447,N_7640,N_8402);
xor U10448 (N_10448,N_7102,N_8222);
nor U10449 (N_10449,N_6454,N_7049);
nand U10450 (N_10450,N_7394,N_8707);
or U10451 (N_10451,N_6320,N_7553);
nand U10452 (N_10452,N_6701,N_7512);
nand U10453 (N_10453,N_7303,N_7784);
and U10454 (N_10454,N_6551,N_7635);
and U10455 (N_10455,N_7609,N_7917);
or U10456 (N_10456,N_7603,N_6672);
nand U10457 (N_10457,N_6087,N_8259);
nor U10458 (N_10458,N_6474,N_6862);
xor U10459 (N_10459,N_7071,N_7397);
or U10460 (N_10460,N_6008,N_6010);
and U10461 (N_10461,N_6674,N_6999);
nand U10462 (N_10462,N_7226,N_8285);
and U10463 (N_10463,N_7814,N_8819);
nor U10464 (N_10464,N_6168,N_8641);
nand U10465 (N_10465,N_8341,N_7893);
and U10466 (N_10466,N_6970,N_8876);
nand U10467 (N_10467,N_7645,N_6166);
nand U10468 (N_10468,N_7270,N_6174);
xor U10469 (N_10469,N_6091,N_6762);
nand U10470 (N_10470,N_6326,N_8856);
nor U10471 (N_10471,N_7130,N_8425);
nand U10472 (N_10472,N_8781,N_7217);
xnor U10473 (N_10473,N_8399,N_6650);
nor U10474 (N_10474,N_8164,N_6752);
nor U10475 (N_10475,N_6070,N_6602);
and U10476 (N_10476,N_6358,N_6262);
xor U10477 (N_10477,N_8422,N_8942);
or U10478 (N_10478,N_7849,N_7409);
or U10479 (N_10479,N_7016,N_8800);
xor U10480 (N_10480,N_7453,N_7864);
xnor U10481 (N_10481,N_7066,N_6029);
or U10482 (N_10482,N_8517,N_8506);
nand U10483 (N_10483,N_6515,N_6015);
and U10484 (N_10484,N_7746,N_7220);
or U10485 (N_10485,N_7241,N_6712);
and U10486 (N_10486,N_6011,N_6947);
and U10487 (N_10487,N_6694,N_7348);
or U10488 (N_10488,N_6084,N_8316);
nor U10489 (N_10489,N_8024,N_7325);
nor U10490 (N_10490,N_6342,N_6302);
or U10491 (N_10491,N_6254,N_8298);
nand U10492 (N_10492,N_7622,N_6208);
xor U10493 (N_10493,N_8640,N_7416);
nor U10494 (N_10494,N_6238,N_8538);
xor U10495 (N_10495,N_7476,N_6433);
or U10496 (N_10496,N_6115,N_6049);
nand U10497 (N_10497,N_8236,N_7275);
and U10498 (N_10498,N_6385,N_6826);
nor U10499 (N_10499,N_7312,N_6969);
and U10500 (N_10500,N_8439,N_8892);
nand U10501 (N_10501,N_6939,N_8212);
and U10502 (N_10502,N_6616,N_8221);
xnor U10503 (N_10503,N_8524,N_8370);
and U10504 (N_10504,N_6525,N_7027);
and U10505 (N_10505,N_6020,N_7148);
nor U10506 (N_10506,N_8199,N_6465);
or U10507 (N_10507,N_8812,N_7753);
nor U10508 (N_10508,N_7804,N_8187);
nand U10509 (N_10509,N_8347,N_6951);
and U10510 (N_10510,N_6657,N_7182);
or U10511 (N_10511,N_8023,N_7125);
xor U10512 (N_10512,N_8316,N_8989);
nand U10513 (N_10513,N_8642,N_8286);
xor U10514 (N_10514,N_8993,N_6542);
xor U10515 (N_10515,N_8211,N_8230);
nand U10516 (N_10516,N_7976,N_7946);
xnor U10517 (N_10517,N_8820,N_7888);
nor U10518 (N_10518,N_8899,N_7016);
xor U10519 (N_10519,N_6744,N_6600);
and U10520 (N_10520,N_6516,N_6204);
nor U10521 (N_10521,N_6505,N_8012);
xnor U10522 (N_10522,N_7708,N_6390);
nor U10523 (N_10523,N_8155,N_7937);
nand U10524 (N_10524,N_7773,N_6171);
and U10525 (N_10525,N_6697,N_8712);
and U10526 (N_10526,N_8448,N_8935);
nor U10527 (N_10527,N_8099,N_8167);
nor U10528 (N_10528,N_7287,N_8597);
nand U10529 (N_10529,N_6003,N_7986);
nor U10530 (N_10530,N_8906,N_6041);
xor U10531 (N_10531,N_6201,N_6327);
or U10532 (N_10532,N_6754,N_7404);
and U10533 (N_10533,N_8640,N_7111);
xor U10534 (N_10534,N_7250,N_8880);
nor U10535 (N_10535,N_7920,N_6392);
xnor U10536 (N_10536,N_6711,N_7949);
nor U10537 (N_10537,N_8555,N_6924);
xnor U10538 (N_10538,N_7333,N_8219);
or U10539 (N_10539,N_7865,N_6188);
xor U10540 (N_10540,N_7977,N_8359);
and U10541 (N_10541,N_6374,N_6161);
xor U10542 (N_10542,N_8764,N_8725);
nand U10543 (N_10543,N_7678,N_7614);
xnor U10544 (N_10544,N_8907,N_7761);
or U10545 (N_10545,N_8722,N_7164);
nor U10546 (N_10546,N_7564,N_8319);
nor U10547 (N_10547,N_8141,N_7540);
nand U10548 (N_10548,N_8790,N_7724);
and U10549 (N_10549,N_7129,N_7401);
xnor U10550 (N_10550,N_7905,N_6054);
or U10551 (N_10551,N_8713,N_6035);
and U10552 (N_10552,N_6419,N_6888);
xnor U10553 (N_10553,N_6193,N_6327);
nand U10554 (N_10554,N_6740,N_6387);
or U10555 (N_10555,N_8287,N_8987);
or U10556 (N_10556,N_6541,N_7165);
xnor U10557 (N_10557,N_8524,N_7800);
xnor U10558 (N_10558,N_7670,N_7727);
nor U10559 (N_10559,N_6817,N_8583);
and U10560 (N_10560,N_6839,N_7501);
or U10561 (N_10561,N_7063,N_8050);
xor U10562 (N_10562,N_6623,N_7144);
nand U10563 (N_10563,N_7529,N_6030);
and U10564 (N_10564,N_6435,N_7195);
nor U10565 (N_10565,N_6710,N_8106);
or U10566 (N_10566,N_7457,N_8767);
and U10567 (N_10567,N_8831,N_7894);
and U10568 (N_10568,N_8807,N_7119);
and U10569 (N_10569,N_8349,N_8711);
nand U10570 (N_10570,N_6904,N_6681);
and U10571 (N_10571,N_6792,N_7697);
xnor U10572 (N_10572,N_6005,N_6226);
nor U10573 (N_10573,N_6010,N_8953);
xor U10574 (N_10574,N_8712,N_6345);
nand U10575 (N_10575,N_6983,N_6665);
xnor U10576 (N_10576,N_7779,N_7719);
nor U10577 (N_10577,N_7920,N_6368);
xor U10578 (N_10578,N_7255,N_8382);
and U10579 (N_10579,N_7450,N_8737);
nor U10580 (N_10580,N_8533,N_7545);
nor U10581 (N_10581,N_7374,N_8358);
or U10582 (N_10582,N_8014,N_6409);
xnor U10583 (N_10583,N_7910,N_8832);
nand U10584 (N_10584,N_8656,N_8790);
xnor U10585 (N_10585,N_8988,N_6214);
nor U10586 (N_10586,N_7690,N_8252);
or U10587 (N_10587,N_8935,N_7619);
nor U10588 (N_10588,N_6583,N_6463);
nand U10589 (N_10589,N_6691,N_8748);
or U10590 (N_10590,N_8911,N_7955);
nor U10591 (N_10591,N_6356,N_6043);
or U10592 (N_10592,N_6128,N_8642);
xor U10593 (N_10593,N_7305,N_6976);
and U10594 (N_10594,N_6369,N_7670);
or U10595 (N_10595,N_7010,N_6074);
xor U10596 (N_10596,N_7365,N_6619);
and U10597 (N_10597,N_7933,N_8856);
xnor U10598 (N_10598,N_6571,N_8210);
nand U10599 (N_10599,N_8659,N_8622);
and U10600 (N_10600,N_6139,N_6852);
nor U10601 (N_10601,N_8050,N_6202);
nand U10602 (N_10602,N_7815,N_7846);
and U10603 (N_10603,N_7296,N_7655);
nand U10604 (N_10604,N_7599,N_7232);
or U10605 (N_10605,N_7556,N_8518);
nor U10606 (N_10606,N_7710,N_6177);
nor U10607 (N_10607,N_8851,N_6733);
or U10608 (N_10608,N_7629,N_6018);
nor U10609 (N_10609,N_8863,N_8224);
or U10610 (N_10610,N_7517,N_7914);
xnor U10611 (N_10611,N_7872,N_8601);
nand U10612 (N_10612,N_7801,N_8778);
nand U10613 (N_10613,N_7478,N_7770);
nand U10614 (N_10614,N_7244,N_6240);
or U10615 (N_10615,N_8442,N_8842);
and U10616 (N_10616,N_6740,N_8994);
or U10617 (N_10617,N_8272,N_6889);
nor U10618 (N_10618,N_7449,N_6415);
nor U10619 (N_10619,N_8038,N_8141);
xnor U10620 (N_10620,N_7937,N_8687);
nand U10621 (N_10621,N_7690,N_6033);
and U10622 (N_10622,N_8028,N_8228);
or U10623 (N_10623,N_7851,N_7416);
xor U10624 (N_10624,N_8427,N_7131);
xor U10625 (N_10625,N_8767,N_7683);
or U10626 (N_10626,N_7775,N_8891);
or U10627 (N_10627,N_6048,N_8222);
xor U10628 (N_10628,N_8757,N_7588);
and U10629 (N_10629,N_6570,N_6700);
nand U10630 (N_10630,N_8910,N_7071);
or U10631 (N_10631,N_6664,N_7233);
and U10632 (N_10632,N_8057,N_8909);
nor U10633 (N_10633,N_7989,N_7215);
nand U10634 (N_10634,N_7951,N_8664);
or U10635 (N_10635,N_6995,N_7313);
and U10636 (N_10636,N_7384,N_7855);
or U10637 (N_10637,N_7141,N_6954);
and U10638 (N_10638,N_7704,N_7050);
nand U10639 (N_10639,N_6142,N_8615);
or U10640 (N_10640,N_7679,N_7293);
nand U10641 (N_10641,N_7831,N_8485);
xnor U10642 (N_10642,N_6140,N_8862);
and U10643 (N_10643,N_7491,N_7481);
nand U10644 (N_10644,N_7373,N_6308);
nor U10645 (N_10645,N_7749,N_8337);
nor U10646 (N_10646,N_8417,N_6912);
xnor U10647 (N_10647,N_6120,N_6681);
nor U10648 (N_10648,N_7574,N_7472);
xor U10649 (N_10649,N_6837,N_8961);
or U10650 (N_10650,N_6628,N_8285);
nand U10651 (N_10651,N_8631,N_6026);
or U10652 (N_10652,N_6529,N_7704);
nand U10653 (N_10653,N_6692,N_7093);
xnor U10654 (N_10654,N_8178,N_7933);
or U10655 (N_10655,N_8060,N_7937);
and U10656 (N_10656,N_6371,N_6701);
nand U10657 (N_10657,N_8924,N_8756);
or U10658 (N_10658,N_8765,N_8233);
nand U10659 (N_10659,N_7523,N_6853);
nand U10660 (N_10660,N_8424,N_8090);
or U10661 (N_10661,N_7613,N_7615);
nor U10662 (N_10662,N_8193,N_7319);
and U10663 (N_10663,N_6162,N_6373);
xnor U10664 (N_10664,N_8209,N_8651);
nor U10665 (N_10665,N_7216,N_6329);
nor U10666 (N_10666,N_8970,N_8386);
and U10667 (N_10667,N_7402,N_7619);
nor U10668 (N_10668,N_7127,N_6424);
nand U10669 (N_10669,N_7741,N_8142);
and U10670 (N_10670,N_7893,N_6856);
or U10671 (N_10671,N_6799,N_6232);
or U10672 (N_10672,N_8940,N_8703);
nand U10673 (N_10673,N_6880,N_7950);
and U10674 (N_10674,N_7273,N_7539);
xor U10675 (N_10675,N_7644,N_7970);
and U10676 (N_10676,N_8519,N_7320);
xnor U10677 (N_10677,N_6883,N_6714);
or U10678 (N_10678,N_6923,N_6493);
and U10679 (N_10679,N_6941,N_8413);
nand U10680 (N_10680,N_8138,N_8923);
and U10681 (N_10681,N_8544,N_7033);
and U10682 (N_10682,N_8249,N_8621);
and U10683 (N_10683,N_6155,N_6460);
nand U10684 (N_10684,N_7136,N_8138);
nor U10685 (N_10685,N_8020,N_6599);
or U10686 (N_10686,N_7782,N_7455);
nor U10687 (N_10687,N_7633,N_6070);
nand U10688 (N_10688,N_7138,N_7173);
xnor U10689 (N_10689,N_6649,N_8444);
and U10690 (N_10690,N_6344,N_8896);
nor U10691 (N_10691,N_6912,N_6467);
nand U10692 (N_10692,N_8275,N_6075);
nand U10693 (N_10693,N_7394,N_6029);
nand U10694 (N_10694,N_6560,N_7151);
nand U10695 (N_10695,N_7101,N_8760);
nor U10696 (N_10696,N_8538,N_8573);
and U10697 (N_10697,N_8335,N_8640);
nand U10698 (N_10698,N_6002,N_7248);
nor U10699 (N_10699,N_6135,N_7268);
and U10700 (N_10700,N_6085,N_6139);
or U10701 (N_10701,N_6757,N_7952);
nand U10702 (N_10702,N_8442,N_6867);
nor U10703 (N_10703,N_7112,N_8213);
xor U10704 (N_10704,N_8246,N_7560);
nor U10705 (N_10705,N_7872,N_6632);
nor U10706 (N_10706,N_8984,N_8746);
nand U10707 (N_10707,N_7772,N_6718);
and U10708 (N_10708,N_8069,N_6008);
and U10709 (N_10709,N_7902,N_6571);
and U10710 (N_10710,N_7730,N_8667);
and U10711 (N_10711,N_6419,N_8747);
nand U10712 (N_10712,N_7482,N_7805);
nor U10713 (N_10713,N_8442,N_8117);
xnor U10714 (N_10714,N_6776,N_7123);
or U10715 (N_10715,N_7887,N_8680);
nor U10716 (N_10716,N_6222,N_6738);
xor U10717 (N_10717,N_7918,N_7169);
nor U10718 (N_10718,N_7432,N_6188);
nor U10719 (N_10719,N_7375,N_8670);
nand U10720 (N_10720,N_6798,N_7752);
nor U10721 (N_10721,N_7369,N_8417);
and U10722 (N_10722,N_6340,N_8148);
nor U10723 (N_10723,N_6387,N_8690);
nand U10724 (N_10724,N_7358,N_7853);
nand U10725 (N_10725,N_6554,N_8532);
or U10726 (N_10726,N_8329,N_8723);
nor U10727 (N_10727,N_6629,N_6132);
or U10728 (N_10728,N_8060,N_6344);
and U10729 (N_10729,N_7561,N_7400);
xor U10730 (N_10730,N_8186,N_7870);
and U10731 (N_10731,N_6674,N_8101);
nor U10732 (N_10732,N_7239,N_6671);
and U10733 (N_10733,N_6185,N_8744);
nand U10734 (N_10734,N_6749,N_6991);
and U10735 (N_10735,N_6444,N_6578);
nand U10736 (N_10736,N_7849,N_8957);
xor U10737 (N_10737,N_6582,N_6081);
nand U10738 (N_10738,N_6256,N_6392);
nor U10739 (N_10739,N_7473,N_6466);
nor U10740 (N_10740,N_6967,N_6450);
and U10741 (N_10741,N_6009,N_6877);
nor U10742 (N_10742,N_7320,N_6123);
and U10743 (N_10743,N_6506,N_7498);
xnor U10744 (N_10744,N_8630,N_7533);
nor U10745 (N_10745,N_7434,N_7518);
nor U10746 (N_10746,N_6929,N_7196);
xor U10747 (N_10747,N_7950,N_7432);
and U10748 (N_10748,N_7272,N_7732);
nand U10749 (N_10749,N_6654,N_7035);
xnor U10750 (N_10750,N_8142,N_7264);
nand U10751 (N_10751,N_8459,N_8812);
nand U10752 (N_10752,N_6264,N_6523);
and U10753 (N_10753,N_7499,N_6982);
or U10754 (N_10754,N_8084,N_7214);
or U10755 (N_10755,N_6776,N_6154);
nand U10756 (N_10756,N_7023,N_7404);
and U10757 (N_10757,N_8444,N_6367);
nand U10758 (N_10758,N_8980,N_6749);
nand U10759 (N_10759,N_8240,N_6311);
nand U10760 (N_10760,N_6752,N_8740);
nor U10761 (N_10761,N_7114,N_6429);
and U10762 (N_10762,N_8394,N_8462);
nand U10763 (N_10763,N_6492,N_8295);
nor U10764 (N_10764,N_7434,N_7265);
xor U10765 (N_10765,N_8245,N_6445);
or U10766 (N_10766,N_6803,N_6999);
and U10767 (N_10767,N_7097,N_7720);
xnor U10768 (N_10768,N_6589,N_6705);
or U10769 (N_10769,N_8873,N_6795);
nand U10770 (N_10770,N_7877,N_8422);
and U10771 (N_10771,N_7022,N_7308);
xnor U10772 (N_10772,N_7263,N_7547);
and U10773 (N_10773,N_7201,N_7295);
nor U10774 (N_10774,N_6302,N_8069);
xnor U10775 (N_10775,N_7161,N_7524);
and U10776 (N_10776,N_8693,N_6340);
nor U10777 (N_10777,N_7153,N_6813);
xnor U10778 (N_10778,N_6276,N_7233);
nand U10779 (N_10779,N_6604,N_8521);
or U10780 (N_10780,N_7887,N_6892);
nor U10781 (N_10781,N_6056,N_8550);
and U10782 (N_10782,N_6404,N_7970);
nand U10783 (N_10783,N_6463,N_6852);
and U10784 (N_10784,N_6489,N_7871);
and U10785 (N_10785,N_8282,N_7309);
xor U10786 (N_10786,N_8917,N_6236);
or U10787 (N_10787,N_6328,N_7131);
nand U10788 (N_10788,N_7009,N_6755);
or U10789 (N_10789,N_8985,N_8215);
xnor U10790 (N_10790,N_7006,N_6783);
xor U10791 (N_10791,N_6339,N_7529);
nor U10792 (N_10792,N_8328,N_7065);
nor U10793 (N_10793,N_6415,N_7770);
nand U10794 (N_10794,N_7632,N_7657);
and U10795 (N_10795,N_8988,N_8333);
nand U10796 (N_10796,N_6381,N_8134);
nand U10797 (N_10797,N_7058,N_8011);
xnor U10798 (N_10798,N_6978,N_7586);
xor U10799 (N_10799,N_8867,N_6256);
or U10800 (N_10800,N_6548,N_6259);
nor U10801 (N_10801,N_7958,N_7331);
nor U10802 (N_10802,N_7909,N_6282);
or U10803 (N_10803,N_6369,N_8837);
and U10804 (N_10804,N_8276,N_7624);
nor U10805 (N_10805,N_7042,N_6585);
nor U10806 (N_10806,N_6924,N_8136);
or U10807 (N_10807,N_8222,N_6609);
nor U10808 (N_10808,N_8031,N_6860);
xnor U10809 (N_10809,N_8398,N_8595);
or U10810 (N_10810,N_7057,N_6679);
and U10811 (N_10811,N_7886,N_8546);
xor U10812 (N_10812,N_7754,N_7971);
xnor U10813 (N_10813,N_7755,N_6176);
nand U10814 (N_10814,N_6775,N_7903);
and U10815 (N_10815,N_8797,N_6810);
xnor U10816 (N_10816,N_8267,N_6641);
nor U10817 (N_10817,N_8637,N_8317);
nand U10818 (N_10818,N_6021,N_8943);
and U10819 (N_10819,N_6070,N_7261);
and U10820 (N_10820,N_6436,N_6221);
xnor U10821 (N_10821,N_7716,N_6571);
or U10822 (N_10822,N_6899,N_7711);
xnor U10823 (N_10823,N_8959,N_8671);
or U10824 (N_10824,N_7989,N_8174);
nor U10825 (N_10825,N_6909,N_7389);
and U10826 (N_10826,N_7964,N_7035);
or U10827 (N_10827,N_6467,N_7790);
or U10828 (N_10828,N_7403,N_7517);
xor U10829 (N_10829,N_6414,N_7209);
nor U10830 (N_10830,N_7113,N_8684);
nand U10831 (N_10831,N_6101,N_6669);
and U10832 (N_10832,N_8790,N_6277);
nor U10833 (N_10833,N_7799,N_7270);
xor U10834 (N_10834,N_8393,N_7252);
nand U10835 (N_10835,N_6552,N_7300);
xnor U10836 (N_10836,N_7212,N_6553);
nor U10837 (N_10837,N_6164,N_7406);
nand U10838 (N_10838,N_7665,N_8113);
xor U10839 (N_10839,N_7362,N_8090);
nor U10840 (N_10840,N_6770,N_7194);
nor U10841 (N_10841,N_7226,N_8460);
and U10842 (N_10842,N_7567,N_7110);
nand U10843 (N_10843,N_6054,N_7769);
xor U10844 (N_10844,N_7491,N_8792);
nand U10845 (N_10845,N_7042,N_6075);
nor U10846 (N_10846,N_6816,N_7395);
and U10847 (N_10847,N_7590,N_7413);
and U10848 (N_10848,N_6507,N_7588);
xor U10849 (N_10849,N_8252,N_8405);
xor U10850 (N_10850,N_8677,N_8891);
xnor U10851 (N_10851,N_6158,N_8579);
nor U10852 (N_10852,N_7011,N_7396);
or U10853 (N_10853,N_6420,N_6314);
and U10854 (N_10854,N_8117,N_7870);
and U10855 (N_10855,N_7603,N_7908);
nand U10856 (N_10856,N_8779,N_8888);
or U10857 (N_10857,N_7350,N_8726);
nand U10858 (N_10858,N_6401,N_8170);
nor U10859 (N_10859,N_7946,N_6736);
or U10860 (N_10860,N_7877,N_8013);
and U10861 (N_10861,N_6731,N_8541);
nand U10862 (N_10862,N_7277,N_6538);
or U10863 (N_10863,N_8388,N_7472);
or U10864 (N_10864,N_8955,N_6087);
and U10865 (N_10865,N_8929,N_7575);
and U10866 (N_10866,N_6854,N_7391);
nor U10867 (N_10867,N_6875,N_6949);
or U10868 (N_10868,N_7277,N_8533);
nor U10869 (N_10869,N_7649,N_8204);
and U10870 (N_10870,N_6441,N_7818);
xnor U10871 (N_10871,N_8050,N_7478);
xor U10872 (N_10872,N_6236,N_8582);
nand U10873 (N_10873,N_8599,N_6673);
nand U10874 (N_10874,N_8106,N_6986);
or U10875 (N_10875,N_7261,N_6722);
or U10876 (N_10876,N_6995,N_8307);
or U10877 (N_10877,N_6217,N_6913);
or U10878 (N_10878,N_8266,N_6484);
or U10879 (N_10879,N_6599,N_8058);
xnor U10880 (N_10880,N_6178,N_8968);
nor U10881 (N_10881,N_8043,N_7540);
xnor U10882 (N_10882,N_8640,N_7662);
nor U10883 (N_10883,N_6777,N_8869);
nor U10884 (N_10884,N_8482,N_6982);
or U10885 (N_10885,N_6204,N_7392);
or U10886 (N_10886,N_8101,N_8834);
and U10887 (N_10887,N_7120,N_8961);
xnor U10888 (N_10888,N_7857,N_7108);
xnor U10889 (N_10889,N_8948,N_7301);
xor U10890 (N_10890,N_7042,N_6283);
and U10891 (N_10891,N_7576,N_8690);
or U10892 (N_10892,N_7547,N_8926);
and U10893 (N_10893,N_8132,N_7822);
or U10894 (N_10894,N_8567,N_7528);
nor U10895 (N_10895,N_8495,N_6996);
xnor U10896 (N_10896,N_6370,N_6331);
xor U10897 (N_10897,N_7522,N_7533);
nand U10898 (N_10898,N_6493,N_8947);
and U10899 (N_10899,N_8595,N_8759);
nand U10900 (N_10900,N_6514,N_7601);
or U10901 (N_10901,N_6459,N_7994);
nand U10902 (N_10902,N_8477,N_6355);
or U10903 (N_10903,N_6810,N_6656);
xnor U10904 (N_10904,N_7642,N_8106);
xnor U10905 (N_10905,N_7571,N_7497);
xnor U10906 (N_10906,N_7766,N_6474);
nor U10907 (N_10907,N_7908,N_6212);
xnor U10908 (N_10908,N_8606,N_8371);
or U10909 (N_10909,N_8079,N_7967);
and U10910 (N_10910,N_7620,N_6425);
and U10911 (N_10911,N_6529,N_6587);
nand U10912 (N_10912,N_7539,N_8819);
nor U10913 (N_10913,N_8447,N_7341);
nand U10914 (N_10914,N_8990,N_8090);
nand U10915 (N_10915,N_8446,N_7716);
or U10916 (N_10916,N_6831,N_8402);
or U10917 (N_10917,N_6588,N_7502);
nor U10918 (N_10918,N_8342,N_8730);
nand U10919 (N_10919,N_8736,N_7388);
or U10920 (N_10920,N_6429,N_8427);
nand U10921 (N_10921,N_8309,N_8925);
nor U10922 (N_10922,N_7566,N_6459);
and U10923 (N_10923,N_6955,N_6005);
nor U10924 (N_10924,N_8536,N_6589);
xnor U10925 (N_10925,N_6325,N_6832);
xor U10926 (N_10926,N_6766,N_8014);
nand U10927 (N_10927,N_8881,N_7428);
or U10928 (N_10928,N_6764,N_8990);
xor U10929 (N_10929,N_7020,N_8557);
or U10930 (N_10930,N_6007,N_7372);
or U10931 (N_10931,N_6125,N_6931);
nor U10932 (N_10932,N_7385,N_8765);
nand U10933 (N_10933,N_7533,N_8309);
xor U10934 (N_10934,N_7992,N_8951);
and U10935 (N_10935,N_7720,N_8013);
xnor U10936 (N_10936,N_7621,N_8600);
nor U10937 (N_10937,N_8544,N_6564);
and U10938 (N_10938,N_8169,N_7407);
xnor U10939 (N_10939,N_8288,N_7366);
or U10940 (N_10940,N_6924,N_8373);
xor U10941 (N_10941,N_7204,N_6411);
nand U10942 (N_10942,N_6108,N_7509);
and U10943 (N_10943,N_8945,N_6798);
or U10944 (N_10944,N_8543,N_6748);
xor U10945 (N_10945,N_8495,N_7155);
nand U10946 (N_10946,N_6603,N_8273);
or U10947 (N_10947,N_7957,N_6379);
xor U10948 (N_10948,N_7458,N_6611);
xnor U10949 (N_10949,N_6339,N_7701);
and U10950 (N_10950,N_7211,N_8796);
nor U10951 (N_10951,N_6799,N_8013);
and U10952 (N_10952,N_7058,N_8908);
or U10953 (N_10953,N_6256,N_6606);
nand U10954 (N_10954,N_7851,N_6724);
or U10955 (N_10955,N_6706,N_7400);
and U10956 (N_10956,N_7797,N_6549);
or U10957 (N_10957,N_7558,N_8917);
nand U10958 (N_10958,N_8166,N_8465);
or U10959 (N_10959,N_7563,N_8466);
and U10960 (N_10960,N_8886,N_7551);
and U10961 (N_10961,N_8436,N_6396);
nor U10962 (N_10962,N_7753,N_6822);
and U10963 (N_10963,N_8267,N_6457);
and U10964 (N_10964,N_7959,N_7675);
or U10965 (N_10965,N_8627,N_8266);
xnor U10966 (N_10966,N_8693,N_6662);
nand U10967 (N_10967,N_7545,N_8292);
and U10968 (N_10968,N_6251,N_6245);
xor U10969 (N_10969,N_7052,N_8082);
or U10970 (N_10970,N_7111,N_6430);
xnor U10971 (N_10971,N_8169,N_7140);
nand U10972 (N_10972,N_8740,N_7860);
nand U10973 (N_10973,N_6537,N_8794);
and U10974 (N_10974,N_7055,N_8527);
or U10975 (N_10975,N_7158,N_7313);
and U10976 (N_10976,N_6050,N_6244);
xnor U10977 (N_10977,N_7631,N_8067);
nor U10978 (N_10978,N_8900,N_8487);
or U10979 (N_10979,N_8536,N_8524);
or U10980 (N_10980,N_7826,N_6344);
or U10981 (N_10981,N_6053,N_6955);
nor U10982 (N_10982,N_6833,N_8770);
and U10983 (N_10983,N_7433,N_7259);
and U10984 (N_10984,N_6723,N_7614);
nor U10985 (N_10985,N_6448,N_8509);
or U10986 (N_10986,N_8751,N_8879);
xor U10987 (N_10987,N_7120,N_8222);
or U10988 (N_10988,N_6518,N_6469);
xor U10989 (N_10989,N_6026,N_8846);
xor U10990 (N_10990,N_6126,N_8504);
and U10991 (N_10991,N_6445,N_8292);
nor U10992 (N_10992,N_7835,N_8247);
xnor U10993 (N_10993,N_7404,N_7753);
or U10994 (N_10994,N_6855,N_8572);
or U10995 (N_10995,N_8260,N_7300);
xnor U10996 (N_10996,N_8404,N_6367);
nand U10997 (N_10997,N_8140,N_7674);
or U10998 (N_10998,N_7244,N_6327);
or U10999 (N_10999,N_6662,N_7950);
or U11000 (N_11000,N_8500,N_6204);
nor U11001 (N_11001,N_7929,N_8138);
xnor U11002 (N_11002,N_7219,N_6822);
or U11003 (N_11003,N_8537,N_8739);
nand U11004 (N_11004,N_6067,N_7131);
or U11005 (N_11005,N_7956,N_8301);
nand U11006 (N_11006,N_6228,N_8982);
nor U11007 (N_11007,N_8333,N_8917);
xor U11008 (N_11008,N_8349,N_8375);
and U11009 (N_11009,N_6091,N_6854);
nor U11010 (N_11010,N_8981,N_8252);
nand U11011 (N_11011,N_7658,N_8871);
and U11012 (N_11012,N_6003,N_8914);
and U11013 (N_11013,N_6436,N_8129);
nand U11014 (N_11014,N_8864,N_6104);
and U11015 (N_11015,N_8064,N_7815);
nor U11016 (N_11016,N_6080,N_7805);
or U11017 (N_11017,N_6989,N_6007);
xor U11018 (N_11018,N_7104,N_6192);
xor U11019 (N_11019,N_8437,N_6576);
and U11020 (N_11020,N_7465,N_6431);
and U11021 (N_11021,N_8428,N_6619);
xnor U11022 (N_11022,N_7617,N_6696);
nor U11023 (N_11023,N_6691,N_8875);
nor U11024 (N_11024,N_6462,N_8186);
nor U11025 (N_11025,N_8700,N_8491);
xor U11026 (N_11026,N_7171,N_6674);
nand U11027 (N_11027,N_6961,N_7786);
or U11028 (N_11028,N_8150,N_6409);
nand U11029 (N_11029,N_7483,N_7723);
nand U11030 (N_11030,N_6985,N_6481);
nand U11031 (N_11031,N_6307,N_7798);
and U11032 (N_11032,N_7046,N_7179);
xor U11033 (N_11033,N_8666,N_7207);
xor U11034 (N_11034,N_8877,N_6288);
or U11035 (N_11035,N_6620,N_7951);
nand U11036 (N_11036,N_7041,N_7531);
xor U11037 (N_11037,N_8733,N_6437);
xnor U11038 (N_11038,N_7428,N_8114);
nand U11039 (N_11039,N_7805,N_8171);
nand U11040 (N_11040,N_7007,N_6300);
nand U11041 (N_11041,N_7461,N_7938);
or U11042 (N_11042,N_8484,N_7010);
and U11043 (N_11043,N_6248,N_8893);
nand U11044 (N_11044,N_8040,N_8542);
xor U11045 (N_11045,N_6155,N_7442);
xnor U11046 (N_11046,N_7003,N_6106);
nor U11047 (N_11047,N_6057,N_8909);
nand U11048 (N_11048,N_8405,N_6639);
or U11049 (N_11049,N_8759,N_7675);
and U11050 (N_11050,N_8095,N_7395);
nor U11051 (N_11051,N_7551,N_8570);
nand U11052 (N_11052,N_8728,N_7956);
nand U11053 (N_11053,N_6861,N_7628);
nand U11054 (N_11054,N_6469,N_8184);
or U11055 (N_11055,N_6942,N_8784);
and U11056 (N_11056,N_8269,N_8389);
nand U11057 (N_11057,N_7211,N_6041);
nand U11058 (N_11058,N_8219,N_7764);
nand U11059 (N_11059,N_7821,N_6913);
or U11060 (N_11060,N_8672,N_8482);
or U11061 (N_11061,N_6510,N_7354);
xnor U11062 (N_11062,N_8091,N_8782);
or U11063 (N_11063,N_7589,N_6635);
and U11064 (N_11064,N_7654,N_6894);
or U11065 (N_11065,N_6265,N_8690);
or U11066 (N_11066,N_6972,N_6985);
and U11067 (N_11067,N_7391,N_6521);
nand U11068 (N_11068,N_7401,N_7372);
or U11069 (N_11069,N_8745,N_6445);
nor U11070 (N_11070,N_6783,N_7741);
or U11071 (N_11071,N_6078,N_7482);
nor U11072 (N_11072,N_6047,N_6368);
xor U11073 (N_11073,N_6361,N_7503);
nor U11074 (N_11074,N_7210,N_6734);
nand U11075 (N_11075,N_7320,N_6569);
nand U11076 (N_11076,N_6219,N_7256);
or U11077 (N_11077,N_7130,N_7006);
nand U11078 (N_11078,N_8636,N_8465);
and U11079 (N_11079,N_6959,N_8731);
and U11080 (N_11080,N_6860,N_6079);
or U11081 (N_11081,N_8605,N_6504);
nand U11082 (N_11082,N_7301,N_6249);
and U11083 (N_11083,N_8837,N_7408);
and U11084 (N_11084,N_8272,N_6505);
or U11085 (N_11085,N_7136,N_7432);
xnor U11086 (N_11086,N_6961,N_8889);
or U11087 (N_11087,N_6550,N_7977);
or U11088 (N_11088,N_6124,N_7942);
and U11089 (N_11089,N_6513,N_8485);
xnor U11090 (N_11090,N_7090,N_8525);
nand U11091 (N_11091,N_7271,N_8475);
xnor U11092 (N_11092,N_7786,N_7448);
xnor U11093 (N_11093,N_8429,N_8219);
and U11094 (N_11094,N_6902,N_7416);
and U11095 (N_11095,N_6420,N_7658);
nand U11096 (N_11096,N_6340,N_6440);
xor U11097 (N_11097,N_6894,N_6356);
or U11098 (N_11098,N_8394,N_8790);
or U11099 (N_11099,N_8732,N_6556);
xor U11100 (N_11100,N_8801,N_6975);
nor U11101 (N_11101,N_6288,N_8926);
nand U11102 (N_11102,N_8295,N_7973);
nand U11103 (N_11103,N_7258,N_7242);
nand U11104 (N_11104,N_6632,N_7179);
or U11105 (N_11105,N_8365,N_6063);
or U11106 (N_11106,N_6968,N_8217);
or U11107 (N_11107,N_6517,N_8196);
or U11108 (N_11108,N_8268,N_8560);
nor U11109 (N_11109,N_6483,N_8165);
nor U11110 (N_11110,N_7064,N_8876);
and U11111 (N_11111,N_8910,N_8572);
and U11112 (N_11112,N_8154,N_7645);
or U11113 (N_11113,N_8733,N_7602);
or U11114 (N_11114,N_6089,N_7883);
nand U11115 (N_11115,N_7518,N_6175);
nand U11116 (N_11116,N_7715,N_6653);
or U11117 (N_11117,N_7056,N_6526);
nor U11118 (N_11118,N_8520,N_7932);
xor U11119 (N_11119,N_6453,N_6776);
or U11120 (N_11120,N_6831,N_6500);
and U11121 (N_11121,N_7992,N_8157);
nor U11122 (N_11122,N_6322,N_6200);
and U11123 (N_11123,N_7962,N_6425);
nor U11124 (N_11124,N_6800,N_7778);
nand U11125 (N_11125,N_7580,N_8335);
nand U11126 (N_11126,N_7906,N_6452);
or U11127 (N_11127,N_7417,N_6223);
or U11128 (N_11128,N_6918,N_6017);
nor U11129 (N_11129,N_7409,N_6256);
or U11130 (N_11130,N_8116,N_6336);
or U11131 (N_11131,N_8296,N_6619);
xor U11132 (N_11132,N_6208,N_8502);
and U11133 (N_11133,N_7615,N_7126);
nor U11134 (N_11134,N_8744,N_6796);
nor U11135 (N_11135,N_7668,N_8270);
or U11136 (N_11136,N_7458,N_8637);
nor U11137 (N_11137,N_6610,N_8279);
xor U11138 (N_11138,N_7618,N_7864);
nand U11139 (N_11139,N_8771,N_6216);
nand U11140 (N_11140,N_7041,N_7375);
nand U11141 (N_11141,N_8348,N_8657);
nand U11142 (N_11142,N_7413,N_7870);
and U11143 (N_11143,N_8808,N_6824);
xor U11144 (N_11144,N_7776,N_6938);
xnor U11145 (N_11145,N_7086,N_8138);
nand U11146 (N_11146,N_6344,N_8922);
and U11147 (N_11147,N_6264,N_6915);
and U11148 (N_11148,N_7936,N_7215);
or U11149 (N_11149,N_8968,N_8034);
and U11150 (N_11150,N_7558,N_8975);
nand U11151 (N_11151,N_8463,N_7397);
and U11152 (N_11152,N_7363,N_8968);
or U11153 (N_11153,N_6586,N_6222);
and U11154 (N_11154,N_7025,N_6050);
or U11155 (N_11155,N_8967,N_7278);
or U11156 (N_11156,N_8647,N_6262);
nor U11157 (N_11157,N_7425,N_7753);
and U11158 (N_11158,N_8911,N_7601);
and U11159 (N_11159,N_7904,N_7039);
or U11160 (N_11160,N_7562,N_6466);
xor U11161 (N_11161,N_8646,N_6035);
xnor U11162 (N_11162,N_7212,N_8121);
and U11163 (N_11163,N_8187,N_6982);
and U11164 (N_11164,N_7414,N_7303);
or U11165 (N_11165,N_8638,N_6116);
nand U11166 (N_11166,N_7337,N_7739);
nor U11167 (N_11167,N_8738,N_8763);
xor U11168 (N_11168,N_8511,N_7807);
and U11169 (N_11169,N_7556,N_8328);
nand U11170 (N_11170,N_7316,N_8174);
nor U11171 (N_11171,N_7690,N_6970);
nand U11172 (N_11172,N_6652,N_7747);
nand U11173 (N_11173,N_7024,N_7213);
nand U11174 (N_11174,N_6141,N_6934);
or U11175 (N_11175,N_6333,N_6754);
and U11176 (N_11176,N_7800,N_7084);
nand U11177 (N_11177,N_6481,N_7181);
nor U11178 (N_11178,N_7892,N_6181);
or U11179 (N_11179,N_8950,N_7252);
nand U11180 (N_11180,N_8967,N_8115);
nand U11181 (N_11181,N_8083,N_6998);
and U11182 (N_11182,N_6796,N_6357);
nand U11183 (N_11183,N_6708,N_8383);
xor U11184 (N_11184,N_8744,N_8440);
xnor U11185 (N_11185,N_8568,N_6561);
nand U11186 (N_11186,N_6082,N_7334);
and U11187 (N_11187,N_8339,N_6233);
and U11188 (N_11188,N_7577,N_6488);
and U11189 (N_11189,N_7482,N_6125);
nor U11190 (N_11190,N_8092,N_8940);
or U11191 (N_11191,N_7155,N_7667);
xnor U11192 (N_11192,N_8434,N_6599);
xnor U11193 (N_11193,N_7528,N_7733);
nand U11194 (N_11194,N_7026,N_6015);
or U11195 (N_11195,N_7701,N_8372);
and U11196 (N_11196,N_7618,N_8046);
or U11197 (N_11197,N_7364,N_8997);
and U11198 (N_11198,N_8696,N_6544);
nand U11199 (N_11199,N_6537,N_6860);
xor U11200 (N_11200,N_7845,N_8786);
nor U11201 (N_11201,N_7759,N_6478);
or U11202 (N_11202,N_8227,N_7685);
or U11203 (N_11203,N_6129,N_7573);
nand U11204 (N_11204,N_8771,N_6944);
or U11205 (N_11205,N_6128,N_6431);
nor U11206 (N_11206,N_6121,N_8759);
xor U11207 (N_11207,N_7931,N_7504);
nor U11208 (N_11208,N_6567,N_8632);
nand U11209 (N_11209,N_7420,N_7953);
or U11210 (N_11210,N_6243,N_8042);
nor U11211 (N_11211,N_7200,N_7208);
nor U11212 (N_11212,N_7688,N_6353);
xor U11213 (N_11213,N_7319,N_8849);
nor U11214 (N_11214,N_7550,N_7732);
xnor U11215 (N_11215,N_8810,N_7866);
nor U11216 (N_11216,N_6141,N_8696);
and U11217 (N_11217,N_7879,N_6607);
nand U11218 (N_11218,N_7362,N_7387);
nor U11219 (N_11219,N_8575,N_6741);
nand U11220 (N_11220,N_8209,N_6186);
or U11221 (N_11221,N_6413,N_7000);
or U11222 (N_11222,N_6002,N_8062);
xnor U11223 (N_11223,N_6826,N_7100);
nor U11224 (N_11224,N_8994,N_7627);
and U11225 (N_11225,N_7690,N_8696);
nand U11226 (N_11226,N_6781,N_6360);
or U11227 (N_11227,N_6257,N_6223);
xor U11228 (N_11228,N_6703,N_8759);
nand U11229 (N_11229,N_7895,N_7115);
nor U11230 (N_11230,N_6938,N_7576);
xnor U11231 (N_11231,N_7647,N_7014);
nand U11232 (N_11232,N_6270,N_6020);
and U11233 (N_11233,N_7117,N_6286);
xor U11234 (N_11234,N_7947,N_6687);
nor U11235 (N_11235,N_8607,N_6532);
or U11236 (N_11236,N_6814,N_8680);
nor U11237 (N_11237,N_7344,N_7280);
or U11238 (N_11238,N_6537,N_6980);
nor U11239 (N_11239,N_6726,N_8304);
nor U11240 (N_11240,N_7892,N_6986);
nor U11241 (N_11241,N_6785,N_6569);
xor U11242 (N_11242,N_8313,N_6787);
and U11243 (N_11243,N_8367,N_8836);
or U11244 (N_11244,N_8108,N_7960);
or U11245 (N_11245,N_7926,N_6500);
xor U11246 (N_11246,N_8766,N_8796);
or U11247 (N_11247,N_8909,N_8500);
xor U11248 (N_11248,N_7706,N_8100);
or U11249 (N_11249,N_6453,N_8295);
nand U11250 (N_11250,N_7531,N_7652);
or U11251 (N_11251,N_6325,N_6868);
xnor U11252 (N_11252,N_6549,N_6828);
xor U11253 (N_11253,N_8235,N_8573);
and U11254 (N_11254,N_7235,N_7576);
nor U11255 (N_11255,N_8027,N_8313);
xor U11256 (N_11256,N_7884,N_7155);
xor U11257 (N_11257,N_7619,N_8568);
or U11258 (N_11258,N_6020,N_8243);
xnor U11259 (N_11259,N_6327,N_8912);
nor U11260 (N_11260,N_6354,N_7300);
nand U11261 (N_11261,N_7564,N_7086);
nor U11262 (N_11262,N_6010,N_8949);
nand U11263 (N_11263,N_6188,N_7186);
xnor U11264 (N_11264,N_7064,N_8736);
nand U11265 (N_11265,N_7779,N_7022);
xnor U11266 (N_11266,N_6343,N_7038);
nand U11267 (N_11267,N_7866,N_7483);
and U11268 (N_11268,N_6750,N_7976);
and U11269 (N_11269,N_6870,N_8113);
xor U11270 (N_11270,N_7963,N_6974);
xor U11271 (N_11271,N_6751,N_8725);
xor U11272 (N_11272,N_8697,N_7640);
nor U11273 (N_11273,N_7593,N_7645);
or U11274 (N_11274,N_7715,N_8618);
nand U11275 (N_11275,N_8840,N_7973);
and U11276 (N_11276,N_8083,N_7320);
nor U11277 (N_11277,N_7402,N_6474);
xnor U11278 (N_11278,N_8367,N_6365);
and U11279 (N_11279,N_7103,N_6591);
xor U11280 (N_11280,N_6285,N_8093);
or U11281 (N_11281,N_6612,N_8589);
xnor U11282 (N_11282,N_8652,N_6839);
nor U11283 (N_11283,N_8294,N_6298);
and U11284 (N_11284,N_8197,N_8469);
and U11285 (N_11285,N_6345,N_8025);
nand U11286 (N_11286,N_6239,N_8974);
nor U11287 (N_11287,N_7265,N_6939);
nand U11288 (N_11288,N_7213,N_8092);
nand U11289 (N_11289,N_7969,N_8358);
and U11290 (N_11290,N_6126,N_8369);
xor U11291 (N_11291,N_6286,N_6830);
nand U11292 (N_11292,N_8342,N_6820);
or U11293 (N_11293,N_7530,N_7027);
nand U11294 (N_11294,N_8234,N_6315);
and U11295 (N_11295,N_7367,N_8158);
nand U11296 (N_11296,N_7358,N_7333);
and U11297 (N_11297,N_6943,N_8831);
or U11298 (N_11298,N_8198,N_6565);
nor U11299 (N_11299,N_8326,N_6639);
and U11300 (N_11300,N_7757,N_7480);
and U11301 (N_11301,N_6630,N_8521);
xnor U11302 (N_11302,N_6979,N_7676);
and U11303 (N_11303,N_8426,N_7465);
xnor U11304 (N_11304,N_7295,N_8552);
nor U11305 (N_11305,N_8014,N_8167);
nor U11306 (N_11306,N_8817,N_8837);
and U11307 (N_11307,N_8050,N_6887);
nor U11308 (N_11308,N_7527,N_8479);
xor U11309 (N_11309,N_7534,N_7244);
and U11310 (N_11310,N_7777,N_7741);
or U11311 (N_11311,N_7348,N_6571);
or U11312 (N_11312,N_7947,N_7174);
nor U11313 (N_11313,N_8994,N_7273);
xnor U11314 (N_11314,N_8048,N_7069);
and U11315 (N_11315,N_7265,N_8130);
xor U11316 (N_11316,N_7128,N_8469);
nor U11317 (N_11317,N_6138,N_6431);
nor U11318 (N_11318,N_8288,N_7279);
nor U11319 (N_11319,N_8881,N_7888);
or U11320 (N_11320,N_7304,N_7654);
and U11321 (N_11321,N_6431,N_6630);
or U11322 (N_11322,N_8903,N_7592);
or U11323 (N_11323,N_7270,N_8870);
or U11324 (N_11324,N_6072,N_6764);
nor U11325 (N_11325,N_6697,N_7336);
nand U11326 (N_11326,N_7381,N_6703);
or U11327 (N_11327,N_6753,N_6571);
nand U11328 (N_11328,N_6794,N_6932);
nor U11329 (N_11329,N_7968,N_7486);
and U11330 (N_11330,N_7455,N_8350);
nor U11331 (N_11331,N_8344,N_8582);
nor U11332 (N_11332,N_6834,N_8724);
xnor U11333 (N_11333,N_8772,N_8371);
xnor U11334 (N_11334,N_7436,N_7843);
nor U11335 (N_11335,N_7790,N_6403);
nand U11336 (N_11336,N_7046,N_6077);
or U11337 (N_11337,N_8543,N_8502);
nand U11338 (N_11338,N_6431,N_7388);
nand U11339 (N_11339,N_7271,N_6132);
nand U11340 (N_11340,N_8318,N_7521);
and U11341 (N_11341,N_6531,N_7978);
nand U11342 (N_11342,N_7657,N_8240);
nand U11343 (N_11343,N_7899,N_6479);
nand U11344 (N_11344,N_8353,N_7583);
nand U11345 (N_11345,N_8601,N_6187);
nor U11346 (N_11346,N_7401,N_6652);
and U11347 (N_11347,N_8248,N_7962);
nor U11348 (N_11348,N_8536,N_6170);
or U11349 (N_11349,N_6926,N_8515);
nor U11350 (N_11350,N_6291,N_6188);
xor U11351 (N_11351,N_7775,N_6058);
xnor U11352 (N_11352,N_6673,N_6582);
xnor U11353 (N_11353,N_6704,N_8258);
nor U11354 (N_11354,N_7031,N_8500);
xor U11355 (N_11355,N_7031,N_7653);
xnor U11356 (N_11356,N_6559,N_7251);
and U11357 (N_11357,N_7472,N_6745);
and U11358 (N_11358,N_6760,N_8315);
nor U11359 (N_11359,N_6368,N_8761);
or U11360 (N_11360,N_7432,N_7483);
nor U11361 (N_11361,N_8947,N_6389);
nand U11362 (N_11362,N_6990,N_8680);
or U11363 (N_11363,N_6621,N_6273);
and U11364 (N_11364,N_6501,N_6335);
and U11365 (N_11365,N_6459,N_7145);
xor U11366 (N_11366,N_8747,N_6729);
and U11367 (N_11367,N_8499,N_6719);
nor U11368 (N_11368,N_8449,N_8684);
or U11369 (N_11369,N_7916,N_6381);
or U11370 (N_11370,N_8682,N_8005);
nand U11371 (N_11371,N_8277,N_7005);
nor U11372 (N_11372,N_7669,N_6692);
xnor U11373 (N_11373,N_7006,N_6931);
xnor U11374 (N_11374,N_8803,N_8024);
nand U11375 (N_11375,N_8091,N_7798);
and U11376 (N_11376,N_6486,N_8242);
or U11377 (N_11377,N_6562,N_8385);
xnor U11378 (N_11378,N_6571,N_7230);
nand U11379 (N_11379,N_7995,N_6761);
nor U11380 (N_11380,N_6727,N_6844);
and U11381 (N_11381,N_8627,N_8862);
xor U11382 (N_11382,N_7009,N_6205);
or U11383 (N_11383,N_8761,N_6193);
xor U11384 (N_11384,N_8495,N_7266);
nor U11385 (N_11385,N_7800,N_8554);
nor U11386 (N_11386,N_6148,N_7183);
or U11387 (N_11387,N_6672,N_8819);
xnor U11388 (N_11388,N_8601,N_7769);
or U11389 (N_11389,N_7886,N_8098);
xnor U11390 (N_11390,N_8832,N_6686);
nor U11391 (N_11391,N_6662,N_6011);
or U11392 (N_11392,N_6218,N_7151);
nor U11393 (N_11393,N_6736,N_6750);
xor U11394 (N_11394,N_8761,N_6010);
or U11395 (N_11395,N_6976,N_6038);
or U11396 (N_11396,N_6212,N_7956);
xnor U11397 (N_11397,N_8968,N_7724);
nor U11398 (N_11398,N_7773,N_7665);
or U11399 (N_11399,N_8789,N_8122);
xnor U11400 (N_11400,N_8509,N_8029);
or U11401 (N_11401,N_6332,N_7805);
and U11402 (N_11402,N_7081,N_6324);
and U11403 (N_11403,N_7029,N_7557);
and U11404 (N_11404,N_6156,N_7907);
or U11405 (N_11405,N_8330,N_8654);
xor U11406 (N_11406,N_7231,N_6292);
and U11407 (N_11407,N_6559,N_7577);
or U11408 (N_11408,N_6091,N_8424);
and U11409 (N_11409,N_8799,N_7375);
and U11410 (N_11410,N_6800,N_7636);
and U11411 (N_11411,N_8678,N_7968);
nor U11412 (N_11412,N_6568,N_8274);
or U11413 (N_11413,N_7774,N_7790);
or U11414 (N_11414,N_6721,N_6201);
nor U11415 (N_11415,N_6226,N_8281);
nand U11416 (N_11416,N_8462,N_7868);
nor U11417 (N_11417,N_7927,N_8219);
xor U11418 (N_11418,N_6883,N_8336);
nor U11419 (N_11419,N_6774,N_7251);
or U11420 (N_11420,N_7123,N_6678);
or U11421 (N_11421,N_6436,N_7258);
xnor U11422 (N_11422,N_8171,N_6160);
or U11423 (N_11423,N_6675,N_8328);
nand U11424 (N_11424,N_8957,N_6933);
nand U11425 (N_11425,N_8964,N_7586);
xor U11426 (N_11426,N_7885,N_6707);
xnor U11427 (N_11427,N_8488,N_7215);
nand U11428 (N_11428,N_6902,N_7393);
nand U11429 (N_11429,N_7798,N_8756);
nor U11430 (N_11430,N_7659,N_7237);
or U11431 (N_11431,N_6424,N_8369);
nor U11432 (N_11432,N_8409,N_7360);
and U11433 (N_11433,N_6830,N_7311);
nor U11434 (N_11434,N_7773,N_6585);
nand U11435 (N_11435,N_6868,N_6980);
nand U11436 (N_11436,N_7140,N_8402);
nand U11437 (N_11437,N_8182,N_7366);
nor U11438 (N_11438,N_8648,N_7352);
and U11439 (N_11439,N_8288,N_8738);
nor U11440 (N_11440,N_8972,N_7903);
xnor U11441 (N_11441,N_8493,N_8788);
and U11442 (N_11442,N_6561,N_8789);
nand U11443 (N_11443,N_8671,N_6905);
and U11444 (N_11444,N_7913,N_6480);
nor U11445 (N_11445,N_7380,N_8420);
and U11446 (N_11446,N_6184,N_8893);
or U11447 (N_11447,N_8080,N_8562);
nor U11448 (N_11448,N_8781,N_7974);
xor U11449 (N_11449,N_8015,N_7752);
or U11450 (N_11450,N_7283,N_8700);
and U11451 (N_11451,N_6819,N_7070);
nand U11452 (N_11452,N_7273,N_6227);
nor U11453 (N_11453,N_8529,N_7448);
xor U11454 (N_11454,N_6920,N_7589);
and U11455 (N_11455,N_8349,N_7227);
nor U11456 (N_11456,N_6045,N_8548);
and U11457 (N_11457,N_7208,N_7738);
and U11458 (N_11458,N_7343,N_7421);
nand U11459 (N_11459,N_6737,N_6818);
and U11460 (N_11460,N_7949,N_8415);
or U11461 (N_11461,N_7710,N_6829);
nand U11462 (N_11462,N_8162,N_6653);
nor U11463 (N_11463,N_8228,N_6989);
xnor U11464 (N_11464,N_7139,N_6268);
and U11465 (N_11465,N_7104,N_6717);
and U11466 (N_11466,N_8101,N_7864);
nand U11467 (N_11467,N_7052,N_6937);
or U11468 (N_11468,N_8091,N_6634);
and U11469 (N_11469,N_6441,N_7260);
xor U11470 (N_11470,N_6192,N_6512);
and U11471 (N_11471,N_6323,N_6373);
and U11472 (N_11472,N_7033,N_8616);
and U11473 (N_11473,N_7531,N_6675);
nor U11474 (N_11474,N_6027,N_8949);
xor U11475 (N_11475,N_6733,N_7747);
or U11476 (N_11476,N_6568,N_6270);
nand U11477 (N_11477,N_8187,N_8955);
xnor U11478 (N_11478,N_6396,N_7112);
or U11479 (N_11479,N_8310,N_8366);
or U11480 (N_11480,N_7069,N_7219);
xor U11481 (N_11481,N_6456,N_7104);
nand U11482 (N_11482,N_7924,N_7474);
and U11483 (N_11483,N_7295,N_6456);
or U11484 (N_11484,N_8716,N_6592);
or U11485 (N_11485,N_7228,N_7811);
or U11486 (N_11486,N_8768,N_7687);
and U11487 (N_11487,N_7794,N_6570);
or U11488 (N_11488,N_8973,N_6984);
and U11489 (N_11489,N_6627,N_6041);
xor U11490 (N_11490,N_7418,N_6758);
and U11491 (N_11491,N_7383,N_8829);
nor U11492 (N_11492,N_6198,N_8423);
or U11493 (N_11493,N_7694,N_8368);
nor U11494 (N_11494,N_6828,N_8764);
or U11495 (N_11495,N_7994,N_7040);
nand U11496 (N_11496,N_8263,N_8319);
nand U11497 (N_11497,N_7579,N_6630);
and U11498 (N_11498,N_6560,N_7698);
and U11499 (N_11499,N_7745,N_6181);
and U11500 (N_11500,N_6636,N_6770);
xor U11501 (N_11501,N_8637,N_8168);
nand U11502 (N_11502,N_7517,N_6298);
nand U11503 (N_11503,N_8951,N_7119);
xor U11504 (N_11504,N_7959,N_6753);
nor U11505 (N_11505,N_7526,N_7720);
nor U11506 (N_11506,N_8602,N_8947);
xnor U11507 (N_11507,N_6736,N_7126);
xnor U11508 (N_11508,N_6511,N_8422);
and U11509 (N_11509,N_7288,N_7661);
nand U11510 (N_11510,N_8555,N_8341);
xnor U11511 (N_11511,N_6954,N_8203);
or U11512 (N_11512,N_6830,N_8263);
or U11513 (N_11513,N_7411,N_7530);
and U11514 (N_11514,N_8298,N_7901);
and U11515 (N_11515,N_8415,N_8064);
nor U11516 (N_11516,N_6174,N_7651);
nor U11517 (N_11517,N_7336,N_7436);
nand U11518 (N_11518,N_8694,N_6254);
nand U11519 (N_11519,N_7264,N_7329);
xnor U11520 (N_11520,N_8635,N_7641);
and U11521 (N_11521,N_6588,N_6625);
xnor U11522 (N_11522,N_7389,N_7671);
xnor U11523 (N_11523,N_8477,N_8922);
and U11524 (N_11524,N_7523,N_8068);
nor U11525 (N_11525,N_6323,N_7610);
xnor U11526 (N_11526,N_6242,N_8530);
nor U11527 (N_11527,N_7877,N_7667);
xor U11528 (N_11528,N_6876,N_6721);
nor U11529 (N_11529,N_7653,N_7243);
xor U11530 (N_11530,N_8800,N_8433);
nor U11531 (N_11531,N_7195,N_6179);
nor U11532 (N_11532,N_6651,N_6544);
or U11533 (N_11533,N_8697,N_7145);
nand U11534 (N_11534,N_7513,N_7394);
nand U11535 (N_11535,N_6714,N_8931);
and U11536 (N_11536,N_8328,N_7540);
nand U11537 (N_11537,N_8874,N_7394);
nor U11538 (N_11538,N_7029,N_6853);
xor U11539 (N_11539,N_6027,N_6415);
nor U11540 (N_11540,N_7076,N_6448);
and U11541 (N_11541,N_6984,N_6377);
or U11542 (N_11542,N_6681,N_7704);
nand U11543 (N_11543,N_8281,N_6590);
nand U11544 (N_11544,N_6389,N_8127);
nor U11545 (N_11545,N_8542,N_8917);
or U11546 (N_11546,N_8272,N_7396);
or U11547 (N_11547,N_6491,N_6892);
and U11548 (N_11548,N_7622,N_6043);
and U11549 (N_11549,N_6815,N_8519);
and U11550 (N_11550,N_8988,N_6836);
xor U11551 (N_11551,N_6951,N_7936);
and U11552 (N_11552,N_7762,N_7874);
and U11553 (N_11553,N_7390,N_6179);
and U11554 (N_11554,N_7962,N_7797);
or U11555 (N_11555,N_6106,N_7803);
xnor U11556 (N_11556,N_8483,N_8395);
nand U11557 (N_11557,N_7120,N_6191);
and U11558 (N_11558,N_6074,N_7417);
nor U11559 (N_11559,N_8739,N_8188);
and U11560 (N_11560,N_8820,N_7540);
nor U11561 (N_11561,N_6663,N_6712);
nand U11562 (N_11562,N_8841,N_8786);
nor U11563 (N_11563,N_8047,N_6348);
nand U11564 (N_11564,N_6105,N_7264);
xor U11565 (N_11565,N_6395,N_8440);
nand U11566 (N_11566,N_8480,N_8455);
xor U11567 (N_11567,N_8481,N_6218);
xnor U11568 (N_11568,N_6492,N_6338);
xor U11569 (N_11569,N_7663,N_8611);
nor U11570 (N_11570,N_8046,N_7640);
nor U11571 (N_11571,N_7609,N_6065);
and U11572 (N_11572,N_6064,N_7003);
nand U11573 (N_11573,N_8590,N_6187);
nand U11574 (N_11574,N_6315,N_7788);
or U11575 (N_11575,N_8286,N_8043);
and U11576 (N_11576,N_6071,N_7209);
or U11577 (N_11577,N_7655,N_6357);
nor U11578 (N_11578,N_6033,N_6143);
nor U11579 (N_11579,N_6575,N_8906);
nand U11580 (N_11580,N_7664,N_8607);
and U11581 (N_11581,N_6306,N_8118);
xor U11582 (N_11582,N_7610,N_6104);
or U11583 (N_11583,N_8896,N_7845);
and U11584 (N_11584,N_6290,N_6730);
or U11585 (N_11585,N_7583,N_8026);
or U11586 (N_11586,N_8666,N_6003);
nor U11587 (N_11587,N_8463,N_8115);
nand U11588 (N_11588,N_6573,N_7625);
xor U11589 (N_11589,N_6190,N_7560);
and U11590 (N_11590,N_6752,N_8766);
nor U11591 (N_11591,N_8003,N_8882);
xnor U11592 (N_11592,N_8350,N_6231);
or U11593 (N_11593,N_8916,N_8183);
or U11594 (N_11594,N_6242,N_7506);
or U11595 (N_11595,N_6927,N_6623);
or U11596 (N_11596,N_8095,N_8792);
nand U11597 (N_11597,N_8068,N_7538);
nor U11598 (N_11598,N_6430,N_6082);
or U11599 (N_11599,N_7479,N_6609);
nand U11600 (N_11600,N_6027,N_6541);
or U11601 (N_11601,N_6940,N_7194);
xnor U11602 (N_11602,N_6390,N_6421);
nand U11603 (N_11603,N_8696,N_6932);
and U11604 (N_11604,N_8212,N_8749);
and U11605 (N_11605,N_6536,N_6822);
xnor U11606 (N_11606,N_8825,N_8878);
nand U11607 (N_11607,N_6722,N_8288);
nor U11608 (N_11608,N_6759,N_8237);
nand U11609 (N_11609,N_8407,N_7622);
or U11610 (N_11610,N_8990,N_8474);
nor U11611 (N_11611,N_8819,N_8733);
nand U11612 (N_11612,N_6322,N_6149);
or U11613 (N_11613,N_8256,N_6949);
or U11614 (N_11614,N_6462,N_7672);
xnor U11615 (N_11615,N_7245,N_7404);
and U11616 (N_11616,N_8220,N_8792);
and U11617 (N_11617,N_7676,N_6429);
and U11618 (N_11618,N_8454,N_8402);
nor U11619 (N_11619,N_6172,N_8945);
xnor U11620 (N_11620,N_7713,N_7231);
and U11621 (N_11621,N_8084,N_6800);
nand U11622 (N_11622,N_7705,N_8777);
xnor U11623 (N_11623,N_7151,N_8194);
nand U11624 (N_11624,N_6350,N_8170);
nand U11625 (N_11625,N_8411,N_6630);
nand U11626 (N_11626,N_8235,N_6257);
or U11627 (N_11627,N_7741,N_8809);
or U11628 (N_11628,N_7652,N_7415);
and U11629 (N_11629,N_7363,N_6754);
nor U11630 (N_11630,N_8332,N_8051);
or U11631 (N_11631,N_7879,N_7157);
and U11632 (N_11632,N_8545,N_6981);
and U11633 (N_11633,N_6097,N_7948);
nor U11634 (N_11634,N_6430,N_8293);
xor U11635 (N_11635,N_8416,N_7135);
xor U11636 (N_11636,N_6741,N_6036);
or U11637 (N_11637,N_7232,N_6970);
and U11638 (N_11638,N_6273,N_8917);
nor U11639 (N_11639,N_6893,N_6220);
nand U11640 (N_11640,N_8624,N_7157);
nand U11641 (N_11641,N_7818,N_8024);
or U11642 (N_11642,N_6286,N_7883);
nor U11643 (N_11643,N_6302,N_7416);
nor U11644 (N_11644,N_8731,N_8468);
nand U11645 (N_11645,N_8854,N_7311);
xor U11646 (N_11646,N_6500,N_8802);
nor U11647 (N_11647,N_8262,N_8653);
and U11648 (N_11648,N_8243,N_6335);
nand U11649 (N_11649,N_6702,N_6859);
nand U11650 (N_11650,N_7135,N_6189);
or U11651 (N_11651,N_8691,N_8406);
nand U11652 (N_11652,N_8427,N_6335);
xnor U11653 (N_11653,N_8405,N_7035);
nand U11654 (N_11654,N_7266,N_8594);
nand U11655 (N_11655,N_7704,N_6223);
or U11656 (N_11656,N_7773,N_8765);
xnor U11657 (N_11657,N_7028,N_7089);
nor U11658 (N_11658,N_6352,N_8792);
xnor U11659 (N_11659,N_8399,N_6426);
nor U11660 (N_11660,N_8006,N_7324);
nor U11661 (N_11661,N_8726,N_7074);
xnor U11662 (N_11662,N_8906,N_6465);
or U11663 (N_11663,N_7581,N_6566);
nor U11664 (N_11664,N_8580,N_8878);
nor U11665 (N_11665,N_8077,N_8313);
nand U11666 (N_11666,N_7092,N_7561);
nor U11667 (N_11667,N_8792,N_7057);
or U11668 (N_11668,N_8258,N_7921);
xor U11669 (N_11669,N_6170,N_8017);
and U11670 (N_11670,N_7176,N_8192);
xnor U11671 (N_11671,N_7040,N_6456);
or U11672 (N_11672,N_7113,N_8870);
and U11673 (N_11673,N_7664,N_8851);
nor U11674 (N_11674,N_8858,N_6292);
nor U11675 (N_11675,N_8402,N_7458);
nor U11676 (N_11676,N_8809,N_7290);
or U11677 (N_11677,N_7245,N_7151);
nor U11678 (N_11678,N_6432,N_7758);
and U11679 (N_11679,N_7203,N_6057);
or U11680 (N_11680,N_7688,N_8345);
and U11681 (N_11681,N_7794,N_8751);
or U11682 (N_11682,N_6205,N_8597);
and U11683 (N_11683,N_7889,N_8522);
and U11684 (N_11684,N_8595,N_7730);
and U11685 (N_11685,N_6166,N_7550);
and U11686 (N_11686,N_6601,N_6878);
or U11687 (N_11687,N_7547,N_8896);
nor U11688 (N_11688,N_6617,N_7407);
nand U11689 (N_11689,N_8981,N_8675);
nor U11690 (N_11690,N_6509,N_7335);
xor U11691 (N_11691,N_6209,N_6979);
and U11692 (N_11692,N_6401,N_8288);
nor U11693 (N_11693,N_6823,N_7836);
nand U11694 (N_11694,N_8056,N_7712);
and U11695 (N_11695,N_7609,N_6478);
nand U11696 (N_11696,N_8054,N_6535);
or U11697 (N_11697,N_8273,N_7071);
xor U11698 (N_11698,N_7754,N_6952);
and U11699 (N_11699,N_8962,N_6352);
nor U11700 (N_11700,N_6380,N_8826);
or U11701 (N_11701,N_8987,N_7119);
xor U11702 (N_11702,N_6296,N_6108);
nand U11703 (N_11703,N_8453,N_6636);
and U11704 (N_11704,N_6405,N_8102);
or U11705 (N_11705,N_6873,N_8596);
nand U11706 (N_11706,N_7103,N_7298);
xor U11707 (N_11707,N_6754,N_6063);
nand U11708 (N_11708,N_6107,N_8337);
xnor U11709 (N_11709,N_7911,N_6941);
nor U11710 (N_11710,N_6706,N_7464);
or U11711 (N_11711,N_7553,N_6459);
or U11712 (N_11712,N_6612,N_7960);
nor U11713 (N_11713,N_6566,N_6110);
or U11714 (N_11714,N_7666,N_8114);
and U11715 (N_11715,N_7380,N_6363);
or U11716 (N_11716,N_8460,N_7660);
and U11717 (N_11717,N_6290,N_8535);
and U11718 (N_11718,N_8825,N_8307);
nand U11719 (N_11719,N_8040,N_6134);
nand U11720 (N_11720,N_6460,N_7519);
xnor U11721 (N_11721,N_6095,N_6967);
xor U11722 (N_11722,N_7264,N_7935);
and U11723 (N_11723,N_6093,N_6005);
xor U11724 (N_11724,N_7860,N_8501);
xnor U11725 (N_11725,N_7187,N_8571);
nor U11726 (N_11726,N_7208,N_6330);
xor U11727 (N_11727,N_6296,N_7045);
and U11728 (N_11728,N_6269,N_8957);
nand U11729 (N_11729,N_8775,N_6025);
nor U11730 (N_11730,N_6250,N_7724);
nor U11731 (N_11731,N_6443,N_7851);
and U11732 (N_11732,N_7050,N_8422);
or U11733 (N_11733,N_6965,N_8037);
nor U11734 (N_11734,N_7882,N_8421);
nor U11735 (N_11735,N_6732,N_8931);
or U11736 (N_11736,N_8056,N_8335);
nand U11737 (N_11737,N_6024,N_7625);
nand U11738 (N_11738,N_7924,N_7407);
and U11739 (N_11739,N_7226,N_7652);
nor U11740 (N_11740,N_6852,N_7157);
xor U11741 (N_11741,N_7373,N_8480);
and U11742 (N_11742,N_6192,N_8900);
or U11743 (N_11743,N_8545,N_8864);
nand U11744 (N_11744,N_6893,N_8999);
and U11745 (N_11745,N_7661,N_7542);
or U11746 (N_11746,N_6407,N_8429);
and U11747 (N_11747,N_7976,N_8523);
and U11748 (N_11748,N_6874,N_7186);
nor U11749 (N_11749,N_7052,N_6879);
nor U11750 (N_11750,N_6995,N_8110);
and U11751 (N_11751,N_8931,N_6842);
nand U11752 (N_11752,N_7856,N_7777);
xor U11753 (N_11753,N_8708,N_7739);
and U11754 (N_11754,N_6295,N_8085);
nor U11755 (N_11755,N_6332,N_6094);
nand U11756 (N_11756,N_8580,N_6071);
nand U11757 (N_11757,N_7185,N_6496);
nor U11758 (N_11758,N_8786,N_6356);
nor U11759 (N_11759,N_7625,N_6037);
xor U11760 (N_11760,N_8926,N_8189);
nand U11761 (N_11761,N_8005,N_8034);
and U11762 (N_11762,N_6314,N_7586);
nand U11763 (N_11763,N_6404,N_8371);
nor U11764 (N_11764,N_6151,N_7744);
or U11765 (N_11765,N_6480,N_6652);
xnor U11766 (N_11766,N_7235,N_7136);
or U11767 (N_11767,N_6481,N_7270);
or U11768 (N_11768,N_6787,N_6480);
nand U11769 (N_11769,N_8921,N_7335);
nor U11770 (N_11770,N_7770,N_8494);
nand U11771 (N_11771,N_8788,N_6621);
or U11772 (N_11772,N_7955,N_7499);
xnor U11773 (N_11773,N_6347,N_7754);
xor U11774 (N_11774,N_7606,N_7495);
nor U11775 (N_11775,N_8021,N_7707);
nor U11776 (N_11776,N_7317,N_6344);
or U11777 (N_11777,N_6368,N_8131);
xor U11778 (N_11778,N_6684,N_6643);
nor U11779 (N_11779,N_7028,N_7016);
nand U11780 (N_11780,N_8567,N_6423);
or U11781 (N_11781,N_6735,N_6729);
and U11782 (N_11782,N_6698,N_8049);
nor U11783 (N_11783,N_8586,N_7858);
nor U11784 (N_11784,N_8409,N_6427);
and U11785 (N_11785,N_7234,N_7959);
xnor U11786 (N_11786,N_6385,N_7278);
or U11787 (N_11787,N_8099,N_8745);
nor U11788 (N_11788,N_7818,N_6298);
nor U11789 (N_11789,N_7807,N_6043);
or U11790 (N_11790,N_6686,N_8058);
xnor U11791 (N_11791,N_7022,N_6775);
nand U11792 (N_11792,N_6808,N_6935);
nor U11793 (N_11793,N_8745,N_7769);
nand U11794 (N_11794,N_8586,N_8364);
and U11795 (N_11795,N_8817,N_7121);
or U11796 (N_11796,N_6147,N_6594);
or U11797 (N_11797,N_8898,N_7633);
or U11798 (N_11798,N_6381,N_7216);
nor U11799 (N_11799,N_6597,N_7640);
nand U11800 (N_11800,N_8865,N_7654);
nor U11801 (N_11801,N_7587,N_7549);
nand U11802 (N_11802,N_6361,N_7019);
or U11803 (N_11803,N_7912,N_8233);
and U11804 (N_11804,N_8195,N_7441);
or U11805 (N_11805,N_8043,N_6650);
and U11806 (N_11806,N_6767,N_6888);
xnor U11807 (N_11807,N_8774,N_8322);
and U11808 (N_11808,N_6990,N_6871);
nand U11809 (N_11809,N_6049,N_8467);
or U11810 (N_11810,N_6869,N_6115);
nand U11811 (N_11811,N_8855,N_8047);
xnor U11812 (N_11812,N_7921,N_6365);
or U11813 (N_11813,N_6490,N_8086);
nor U11814 (N_11814,N_7511,N_8458);
and U11815 (N_11815,N_6693,N_6369);
and U11816 (N_11816,N_6652,N_8031);
and U11817 (N_11817,N_7531,N_8390);
xor U11818 (N_11818,N_6284,N_7276);
xor U11819 (N_11819,N_7133,N_8639);
nand U11820 (N_11820,N_6548,N_7740);
or U11821 (N_11821,N_7692,N_8865);
or U11822 (N_11822,N_6559,N_8176);
xor U11823 (N_11823,N_7051,N_6269);
xnor U11824 (N_11824,N_8354,N_7942);
and U11825 (N_11825,N_6595,N_8042);
and U11826 (N_11826,N_8646,N_7769);
nand U11827 (N_11827,N_7980,N_6686);
nor U11828 (N_11828,N_7426,N_8522);
nand U11829 (N_11829,N_6235,N_8929);
or U11830 (N_11830,N_8641,N_6863);
and U11831 (N_11831,N_8052,N_6311);
xnor U11832 (N_11832,N_7789,N_6229);
or U11833 (N_11833,N_8745,N_7375);
and U11834 (N_11834,N_8774,N_8476);
nor U11835 (N_11835,N_8165,N_6920);
or U11836 (N_11836,N_6588,N_6575);
xnor U11837 (N_11837,N_6790,N_6952);
or U11838 (N_11838,N_6119,N_7548);
and U11839 (N_11839,N_8925,N_6722);
nor U11840 (N_11840,N_6820,N_8776);
xor U11841 (N_11841,N_6052,N_6908);
xnor U11842 (N_11842,N_6845,N_7520);
xor U11843 (N_11843,N_8622,N_8662);
xor U11844 (N_11844,N_6614,N_7778);
and U11845 (N_11845,N_7854,N_6215);
or U11846 (N_11846,N_7289,N_7394);
or U11847 (N_11847,N_6248,N_7913);
nand U11848 (N_11848,N_8984,N_6943);
nor U11849 (N_11849,N_7788,N_6388);
nor U11850 (N_11850,N_6936,N_8402);
or U11851 (N_11851,N_6260,N_7693);
or U11852 (N_11852,N_6406,N_8423);
xnor U11853 (N_11853,N_7101,N_7034);
nor U11854 (N_11854,N_7931,N_6528);
nand U11855 (N_11855,N_7720,N_8475);
nor U11856 (N_11856,N_7206,N_6204);
or U11857 (N_11857,N_6326,N_7134);
nor U11858 (N_11858,N_8755,N_7935);
or U11859 (N_11859,N_6837,N_6286);
xnor U11860 (N_11860,N_7582,N_6287);
nor U11861 (N_11861,N_6311,N_8375);
or U11862 (N_11862,N_8728,N_6735);
and U11863 (N_11863,N_6317,N_6678);
nand U11864 (N_11864,N_8460,N_6254);
and U11865 (N_11865,N_8948,N_6949);
and U11866 (N_11866,N_6100,N_8542);
and U11867 (N_11867,N_7901,N_6858);
nor U11868 (N_11868,N_6236,N_8671);
xnor U11869 (N_11869,N_6982,N_6929);
and U11870 (N_11870,N_6467,N_6703);
or U11871 (N_11871,N_8466,N_6697);
nor U11872 (N_11872,N_8695,N_6519);
nand U11873 (N_11873,N_7030,N_8270);
nand U11874 (N_11874,N_7985,N_6765);
or U11875 (N_11875,N_8855,N_6500);
nor U11876 (N_11876,N_7844,N_8184);
nand U11877 (N_11877,N_6077,N_7975);
nor U11878 (N_11878,N_8562,N_7795);
and U11879 (N_11879,N_8030,N_8772);
nand U11880 (N_11880,N_8138,N_7062);
xor U11881 (N_11881,N_8794,N_6759);
nor U11882 (N_11882,N_6147,N_8431);
nand U11883 (N_11883,N_6543,N_8882);
xnor U11884 (N_11884,N_7050,N_8595);
nor U11885 (N_11885,N_6508,N_6549);
nand U11886 (N_11886,N_6244,N_6870);
nand U11887 (N_11887,N_6412,N_7733);
nand U11888 (N_11888,N_8399,N_8698);
and U11889 (N_11889,N_6932,N_8526);
nor U11890 (N_11890,N_8178,N_7818);
and U11891 (N_11891,N_6655,N_7636);
nand U11892 (N_11892,N_8400,N_7126);
nand U11893 (N_11893,N_6313,N_6795);
and U11894 (N_11894,N_6673,N_6553);
or U11895 (N_11895,N_8130,N_6736);
xor U11896 (N_11896,N_6028,N_8326);
or U11897 (N_11897,N_7890,N_6013);
nor U11898 (N_11898,N_7683,N_7544);
nand U11899 (N_11899,N_6763,N_6453);
and U11900 (N_11900,N_8418,N_8132);
nor U11901 (N_11901,N_8399,N_6239);
and U11902 (N_11902,N_7700,N_6783);
and U11903 (N_11903,N_8688,N_6694);
nand U11904 (N_11904,N_8329,N_8505);
nand U11905 (N_11905,N_6452,N_7210);
nor U11906 (N_11906,N_6633,N_7114);
xor U11907 (N_11907,N_8765,N_8101);
and U11908 (N_11908,N_8508,N_6532);
or U11909 (N_11909,N_8051,N_6763);
and U11910 (N_11910,N_7085,N_7769);
and U11911 (N_11911,N_8850,N_8559);
nor U11912 (N_11912,N_7423,N_7485);
nand U11913 (N_11913,N_8464,N_6731);
xor U11914 (N_11914,N_7579,N_6213);
nand U11915 (N_11915,N_7761,N_7064);
xor U11916 (N_11916,N_8429,N_7996);
and U11917 (N_11917,N_7783,N_8328);
or U11918 (N_11918,N_6452,N_6349);
or U11919 (N_11919,N_7766,N_6316);
and U11920 (N_11920,N_7246,N_8619);
or U11921 (N_11921,N_6002,N_6175);
nand U11922 (N_11922,N_8760,N_6277);
nand U11923 (N_11923,N_7910,N_8403);
nand U11924 (N_11924,N_6429,N_8578);
and U11925 (N_11925,N_7464,N_7718);
nor U11926 (N_11926,N_6185,N_7875);
and U11927 (N_11927,N_8733,N_6610);
nor U11928 (N_11928,N_7145,N_8355);
nor U11929 (N_11929,N_6034,N_8315);
and U11930 (N_11930,N_7779,N_6582);
nand U11931 (N_11931,N_6498,N_8269);
xor U11932 (N_11932,N_8776,N_7793);
or U11933 (N_11933,N_6834,N_8116);
and U11934 (N_11934,N_7835,N_6866);
xor U11935 (N_11935,N_8328,N_7875);
xnor U11936 (N_11936,N_8368,N_6199);
xnor U11937 (N_11937,N_6612,N_7935);
nand U11938 (N_11938,N_7152,N_6468);
nand U11939 (N_11939,N_6629,N_8749);
nand U11940 (N_11940,N_6348,N_7404);
and U11941 (N_11941,N_6119,N_7161);
or U11942 (N_11942,N_8623,N_7761);
nor U11943 (N_11943,N_8579,N_6525);
and U11944 (N_11944,N_8714,N_6851);
nand U11945 (N_11945,N_8591,N_7574);
or U11946 (N_11946,N_8283,N_7965);
nand U11947 (N_11947,N_7505,N_8962);
and U11948 (N_11948,N_7197,N_8359);
and U11949 (N_11949,N_6379,N_6295);
xnor U11950 (N_11950,N_6198,N_8119);
nor U11951 (N_11951,N_7243,N_8223);
nor U11952 (N_11952,N_8925,N_6517);
nand U11953 (N_11953,N_7933,N_6387);
and U11954 (N_11954,N_8505,N_6731);
nor U11955 (N_11955,N_6879,N_7063);
or U11956 (N_11956,N_7327,N_8162);
xor U11957 (N_11957,N_7968,N_6192);
nand U11958 (N_11958,N_7137,N_7157);
and U11959 (N_11959,N_7688,N_6072);
nor U11960 (N_11960,N_6877,N_6843);
nor U11961 (N_11961,N_7704,N_8868);
nand U11962 (N_11962,N_7397,N_6322);
nor U11963 (N_11963,N_6807,N_8809);
nor U11964 (N_11964,N_8101,N_8588);
and U11965 (N_11965,N_7244,N_8214);
or U11966 (N_11966,N_7119,N_8027);
nand U11967 (N_11967,N_8480,N_8976);
and U11968 (N_11968,N_7602,N_7863);
xnor U11969 (N_11969,N_7347,N_6601);
xor U11970 (N_11970,N_8929,N_8190);
or U11971 (N_11971,N_6772,N_8226);
or U11972 (N_11972,N_8988,N_8955);
nand U11973 (N_11973,N_6758,N_6132);
xnor U11974 (N_11974,N_8792,N_7718);
nand U11975 (N_11975,N_8061,N_8781);
xnor U11976 (N_11976,N_6466,N_6463);
xnor U11977 (N_11977,N_7739,N_7605);
nor U11978 (N_11978,N_6476,N_7583);
and U11979 (N_11979,N_7871,N_6964);
or U11980 (N_11980,N_6792,N_8389);
xnor U11981 (N_11981,N_6855,N_8645);
or U11982 (N_11982,N_7146,N_8894);
or U11983 (N_11983,N_7655,N_6360);
nand U11984 (N_11984,N_7244,N_6495);
xnor U11985 (N_11985,N_6684,N_8707);
nor U11986 (N_11986,N_8419,N_8459);
nand U11987 (N_11987,N_8227,N_8635);
nand U11988 (N_11988,N_8412,N_8706);
xnor U11989 (N_11989,N_8648,N_6719);
and U11990 (N_11990,N_6934,N_7618);
nand U11991 (N_11991,N_7657,N_8360);
and U11992 (N_11992,N_8472,N_7349);
nor U11993 (N_11993,N_7894,N_6307);
and U11994 (N_11994,N_7317,N_7528);
or U11995 (N_11995,N_8176,N_7592);
nor U11996 (N_11996,N_6936,N_8924);
nand U11997 (N_11997,N_8170,N_7668);
nand U11998 (N_11998,N_7795,N_8511);
and U11999 (N_11999,N_7121,N_6499);
nand U12000 (N_12000,N_11493,N_9716);
and U12001 (N_12001,N_10011,N_9363);
or U12002 (N_12002,N_9864,N_10639);
xnor U12003 (N_12003,N_10718,N_9167);
nand U12004 (N_12004,N_9302,N_9830);
and U12005 (N_12005,N_9658,N_10697);
nor U12006 (N_12006,N_10229,N_10115);
nor U12007 (N_12007,N_9389,N_10520);
or U12008 (N_12008,N_10852,N_11820);
and U12009 (N_12009,N_10197,N_10965);
nand U12010 (N_12010,N_10098,N_10044);
and U12011 (N_12011,N_10861,N_11763);
nor U12012 (N_12012,N_10045,N_10300);
nor U12013 (N_12013,N_10938,N_11108);
nor U12014 (N_12014,N_10502,N_9917);
nand U12015 (N_12015,N_10326,N_10913);
and U12016 (N_12016,N_9979,N_11170);
xor U12017 (N_12017,N_11344,N_9464);
nor U12018 (N_12018,N_11421,N_11691);
nor U12019 (N_12019,N_9121,N_9843);
xor U12020 (N_12020,N_9606,N_10695);
nor U12021 (N_12021,N_10422,N_9100);
or U12022 (N_12022,N_10220,N_9504);
xnor U12023 (N_12023,N_9275,N_10734);
nand U12024 (N_12024,N_11652,N_11321);
nor U12025 (N_12025,N_11009,N_10386);
nor U12026 (N_12026,N_9184,N_11625);
nor U12027 (N_12027,N_9530,N_9962);
nand U12028 (N_12028,N_11517,N_11392);
xnor U12029 (N_12029,N_9286,N_10435);
nor U12030 (N_12030,N_9891,N_9812);
nor U12031 (N_12031,N_10963,N_10975);
xor U12032 (N_12032,N_10807,N_10318);
or U12033 (N_12033,N_10692,N_11569);
or U12034 (N_12034,N_10077,N_9294);
nand U12035 (N_12035,N_11035,N_11702);
nand U12036 (N_12036,N_10382,N_11119);
and U12037 (N_12037,N_11232,N_11315);
and U12038 (N_12038,N_11249,N_9729);
xor U12039 (N_12039,N_11647,N_10768);
nand U12040 (N_12040,N_10980,N_9905);
nor U12041 (N_12041,N_10253,N_11582);
and U12042 (N_12042,N_9300,N_10739);
nand U12043 (N_12043,N_9580,N_9863);
xnor U12044 (N_12044,N_11020,N_10612);
and U12045 (N_12045,N_10645,N_9157);
or U12046 (N_12046,N_11914,N_10978);
or U12047 (N_12047,N_10711,N_11113);
or U12048 (N_12048,N_11062,N_11649);
nand U12049 (N_12049,N_10727,N_10407);
nor U12050 (N_12050,N_11061,N_9485);
or U12051 (N_12051,N_9595,N_9524);
or U12052 (N_12052,N_9258,N_10927);
nand U12053 (N_12053,N_11380,N_9352);
nor U12054 (N_12054,N_10555,N_9357);
nor U12055 (N_12055,N_10104,N_10821);
xnor U12056 (N_12056,N_9832,N_10515);
nand U12057 (N_12057,N_10616,N_9028);
or U12058 (N_12058,N_10819,N_10730);
or U12059 (N_12059,N_11995,N_11431);
nor U12060 (N_12060,N_9124,N_10690);
nor U12061 (N_12061,N_11197,N_10689);
xnor U12062 (N_12062,N_11484,N_11561);
nor U12063 (N_12063,N_9949,N_10056);
or U12064 (N_12064,N_10346,N_10181);
and U12065 (N_12065,N_10342,N_10859);
nand U12066 (N_12066,N_10619,N_11055);
nor U12067 (N_12067,N_11362,N_10336);
xnor U12068 (N_12068,N_11048,N_10775);
and U12069 (N_12069,N_9860,N_11111);
nand U12070 (N_12070,N_10200,N_9734);
nor U12071 (N_12071,N_11879,N_10420);
nor U12072 (N_12072,N_9492,N_11328);
xor U12073 (N_12073,N_9248,N_10273);
or U12074 (N_12074,N_9410,N_9427);
and U12075 (N_12075,N_11872,N_9977);
nand U12076 (N_12076,N_10446,N_9011);
or U12077 (N_12077,N_10479,N_10554);
nor U12078 (N_12078,N_11643,N_9455);
nand U12079 (N_12079,N_9365,N_11548);
and U12080 (N_12080,N_10482,N_9088);
nand U12081 (N_12081,N_10939,N_10603);
xor U12082 (N_12082,N_11278,N_11984);
or U12083 (N_12083,N_11019,N_10150);
nand U12084 (N_12084,N_9256,N_10785);
xnor U12085 (N_12085,N_10163,N_11211);
or U12086 (N_12086,N_10125,N_9277);
nand U12087 (N_12087,N_11758,N_9975);
or U12088 (N_12088,N_10224,N_11853);
and U12089 (N_12089,N_10109,N_9325);
xor U12090 (N_12090,N_9963,N_10545);
xor U12091 (N_12091,N_11774,N_11870);
nor U12092 (N_12092,N_9204,N_11078);
nand U12093 (N_12093,N_9902,N_10086);
or U12094 (N_12094,N_9055,N_9933);
nand U12095 (N_12095,N_10982,N_9845);
xor U12096 (N_12096,N_10550,N_11951);
and U12097 (N_12097,N_11699,N_11496);
xnor U12098 (N_12098,N_9825,N_10284);
nor U12099 (N_12099,N_11830,N_10924);
nand U12100 (N_12100,N_10486,N_9487);
or U12101 (N_12101,N_10454,N_10298);
and U12102 (N_12102,N_11653,N_11961);
nand U12103 (N_12103,N_11865,N_11139);
nand U12104 (N_12104,N_10410,N_10055);
or U12105 (N_12105,N_11573,N_10989);
and U12106 (N_12106,N_10276,N_10837);
or U12107 (N_12107,N_9925,N_11129);
nor U12108 (N_12108,N_9225,N_9641);
nor U12109 (N_12109,N_11439,N_11401);
nand U12110 (N_12110,N_10018,N_11618);
nor U12111 (N_12111,N_11192,N_10042);
or U12112 (N_12112,N_11958,N_11550);
nor U12113 (N_12113,N_9445,N_11724);
or U12114 (N_12114,N_9871,N_9936);
xnor U12115 (N_12115,N_11990,N_10249);
and U12116 (N_12116,N_11179,N_11474);
nor U12117 (N_12117,N_9875,N_11148);
xnor U12118 (N_12118,N_10970,N_9746);
nor U12119 (N_12119,N_9113,N_10396);
and U12120 (N_12120,N_11755,N_10987);
nand U12121 (N_12121,N_11181,N_11571);
nor U12122 (N_12122,N_10521,N_11043);
or U12123 (N_12123,N_11521,N_11268);
and U12124 (N_12124,N_11704,N_11846);
xnor U12125 (N_12125,N_11432,N_9222);
nor U12126 (N_12126,N_10010,N_10789);
nand U12127 (N_12127,N_10823,N_10857);
and U12128 (N_12128,N_11271,N_10793);
and U12129 (N_12129,N_10904,N_10874);
or U12130 (N_12130,N_10642,N_9609);
nor U12131 (N_12131,N_10828,N_9136);
nand U12132 (N_12132,N_9235,N_11992);
or U12133 (N_12133,N_11188,N_11930);
or U12134 (N_12134,N_11174,N_11240);
xor U12135 (N_12135,N_10577,N_11359);
nand U12136 (N_12136,N_10050,N_10751);
and U12137 (N_12137,N_10031,N_9549);
or U12138 (N_12138,N_11418,N_9027);
nand U12139 (N_12139,N_10111,N_11160);
nor U12140 (N_12140,N_11650,N_11156);
nor U12141 (N_12141,N_9773,N_9638);
and U12142 (N_12142,N_11149,N_10095);
nor U12143 (N_12143,N_10879,N_11182);
nor U12144 (N_12144,N_11244,N_11054);
xnor U12145 (N_12145,N_9698,N_10663);
xor U12146 (N_12146,N_11821,N_9588);
or U12147 (N_12147,N_11497,N_10764);
nand U12148 (N_12148,N_9444,N_9061);
nor U12149 (N_12149,N_10759,N_9457);
xnor U12150 (N_12150,N_10270,N_10184);
xnor U12151 (N_12151,N_10929,N_10331);
and U12152 (N_12152,N_10911,N_10434);
nor U12153 (N_12153,N_11639,N_11023);
xnor U12154 (N_12154,N_10899,N_9318);
and U12155 (N_12155,N_10377,N_10179);
or U12156 (N_12156,N_10796,N_10441);
nor U12157 (N_12157,N_9390,N_9801);
nor U12158 (N_12158,N_11534,N_9818);
nor U12159 (N_12159,N_11030,N_10263);
or U12160 (N_12160,N_11782,N_11016);
or U12161 (N_12161,N_11620,N_11936);
xnor U12162 (N_12162,N_10745,N_9846);
xor U12163 (N_12163,N_10790,N_10091);
nor U12164 (N_12164,N_11089,N_9626);
nand U12165 (N_12165,N_11709,N_9508);
nor U12166 (N_12166,N_11124,N_9346);
xor U12167 (N_12167,N_10315,N_10824);
nand U12168 (N_12168,N_10430,N_10211);
nor U12169 (N_12169,N_10539,N_11404);
nor U12170 (N_12170,N_11634,N_10247);
nand U12171 (N_12171,N_10267,N_11388);
or U12172 (N_12172,N_10130,N_9397);
and U12173 (N_12173,N_9023,N_9896);
xor U12174 (N_12174,N_9715,N_9534);
xnor U12175 (N_12175,N_11504,N_11577);
or U12176 (N_12176,N_11415,N_10035);
nor U12177 (N_12177,N_9035,N_9705);
or U12178 (N_12178,N_11799,N_11308);
nand U12179 (N_12179,N_10912,N_11520);
or U12180 (N_12180,N_9495,N_9425);
and U12181 (N_12181,N_9998,N_9470);
and U12182 (N_12182,N_10032,N_11880);
nor U12183 (N_12183,N_9065,N_10239);
nand U12184 (N_12184,N_11045,N_10292);
or U12185 (N_12185,N_9345,N_10078);
nand U12186 (N_12186,N_11884,N_11364);
and U12187 (N_12187,N_9795,N_9141);
and U12188 (N_12188,N_10508,N_9461);
xor U12189 (N_12189,N_9146,N_11395);
nor U12190 (N_12190,N_9759,N_11233);
or U12191 (N_12191,N_9765,N_10702);
or U12192 (N_12192,N_10848,N_10934);
and U12193 (N_12193,N_10997,N_11728);
or U12194 (N_12194,N_11097,N_11437);
nand U12195 (N_12195,N_10607,N_9192);
and U12196 (N_12196,N_11658,N_10665);
nor U12197 (N_12197,N_9770,N_10002);
nor U12198 (N_12198,N_11163,N_9736);
or U12199 (N_12199,N_10408,N_9369);
nor U12200 (N_12200,N_9976,N_9964);
and U12201 (N_12201,N_9500,N_11266);
and U12202 (N_12202,N_11127,N_11340);
and U12203 (N_12203,N_9551,N_11834);
nor U12204 (N_12204,N_9719,N_10684);
and U12205 (N_12205,N_10752,N_10747);
or U12206 (N_12206,N_10058,N_10312);
or U12207 (N_12207,N_11447,N_9030);
or U12208 (N_12208,N_9611,N_9407);
and U12209 (N_12209,N_11076,N_10809);
and U12210 (N_12210,N_10835,N_9456);
nand U12211 (N_12211,N_11071,N_9331);
xnor U12212 (N_12212,N_11559,N_10503);
nand U12213 (N_12213,N_9819,N_11001);
or U12214 (N_12214,N_10631,N_10059);
nand U12215 (N_12215,N_9560,N_10514);
or U12216 (N_12216,N_10105,N_11794);
nor U12217 (N_12217,N_9873,N_9955);
or U12218 (N_12218,N_10381,N_11903);
xnor U12219 (N_12219,N_9499,N_9667);
xor U12220 (N_12220,N_10632,N_10240);
xor U12221 (N_12221,N_11736,N_9627);
nand U12222 (N_12222,N_11003,N_11463);
and U12223 (N_12223,N_10582,N_9637);
xor U12224 (N_12224,N_11205,N_11682);
or U12225 (N_12225,N_10588,N_11579);
nor U12226 (N_12226,N_11191,N_10327);
and U12227 (N_12227,N_11310,N_11049);
nand U12228 (N_12228,N_9058,N_10943);
nand U12229 (N_12229,N_9621,N_9583);
or U12230 (N_12230,N_11118,N_10216);
or U12231 (N_12231,N_11688,N_10624);
nand U12232 (N_12232,N_11341,N_11768);
nor U12233 (N_12233,N_9285,N_9233);
xnor U12234 (N_12234,N_9631,N_11263);
or U12235 (N_12235,N_10073,N_9985);
and U12236 (N_12236,N_11350,N_11087);
or U12237 (N_12237,N_10235,N_11540);
nor U12238 (N_12238,N_11370,N_9144);
or U12239 (N_12239,N_10260,N_10748);
or U12240 (N_12240,N_11706,N_9350);
nor U12241 (N_12241,N_11096,N_9243);
xor U12242 (N_12242,N_10082,N_10969);
nor U12243 (N_12243,N_10413,N_9993);
nor U12244 (N_12244,N_11151,N_10596);
nand U12245 (N_12245,N_11198,N_10760);
xor U12246 (N_12246,N_9351,N_11982);
and U12247 (N_12247,N_9909,N_10345);
nand U12248 (N_12248,N_11664,N_10783);
and U12249 (N_12249,N_9912,N_11121);
or U12250 (N_12250,N_9571,N_11812);
xor U12251 (N_12251,N_9661,N_10173);
nand U12252 (N_12252,N_10827,N_11294);
xor U12253 (N_12253,N_10391,N_10025);
nand U12254 (N_12254,N_9854,N_10255);
nand U12255 (N_12255,N_11318,N_11367);
and U12256 (N_12256,N_9249,N_10724);
nor U12257 (N_12257,N_11122,N_10708);
nor U12258 (N_12258,N_9409,N_9349);
nand U12259 (N_12259,N_11331,N_10669);
or U12260 (N_12260,N_11720,N_11464);
or U12261 (N_12261,N_10895,N_9737);
xor U12262 (N_12262,N_11874,N_9980);
nor U12263 (N_12263,N_10875,N_9572);
xor U12264 (N_12264,N_11826,N_11923);
nor U12265 (N_12265,N_11901,N_10483);
xnor U12266 (N_12266,N_10530,N_9408);
nand U12267 (N_12267,N_9198,N_10106);
nor U12268 (N_12268,N_9502,N_9344);
or U12269 (N_12269,N_9454,N_10473);
or U12270 (N_12270,N_10758,N_9991);
and U12271 (N_12271,N_10057,N_9512);
or U12272 (N_12272,N_11592,N_10769);
nand U12273 (N_12273,N_10426,N_9660);
and U12274 (N_12274,N_11539,N_11665);
nand U12275 (N_12275,N_9359,N_11802);
nor U12276 (N_12276,N_10524,N_11811);
nand U12277 (N_12277,N_10822,N_10755);
and U12278 (N_12278,N_9813,N_11337);
nor U12279 (N_12279,N_10676,N_10634);
xnor U12280 (N_12280,N_9663,N_11186);
or U12281 (N_12281,N_11717,N_9191);
nor U12282 (N_12282,N_9617,N_10121);
and U12283 (N_12283,N_9724,N_9388);
or U12284 (N_12284,N_10960,N_10876);
nor U12285 (N_12285,N_11301,N_9927);
nand U12286 (N_12286,N_9634,N_10762);
and U12287 (N_12287,N_11695,N_9155);
and U12288 (N_12288,N_10048,N_9423);
or U12289 (N_12289,N_10471,N_9266);
nand U12290 (N_12290,N_9440,N_11784);
xor U12291 (N_12291,N_9918,N_11660);
nand U12292 (N_12292,N_10074,N_9794);
or U12293 (N_12293,N_11200,N_9796);
or U12294 (N_12294,N_10818,N_11679);
and U12295 (N_12295,N_11687,N_10275);
nor U12296 (N_12296,N_11397,N_9041);
nor U12297 (N_12297,N_10604,N_10628);
or U12298 (N_12298,N_9757,N_10232);
nor U12299 (N_12299,N_11748,N_9378);
nand U12300 (N_12300,N_10404,N_9594);
nor U12301 (N_12301,N_9209,N_11265);
nor U12302 (N_12302,N_10863,N_10221);
xnor U12303 (N_12303,N_10036,N_10366);
nand U12304 (N_12304,N_9600,N_9342);
and U12305 (N_12305,N_11269,N_11937);
xor U12306 (N_12306,N_11231,N_11985);
and U12307 (N_12307,N_9134,N_10333);
xnor U12308 (N_12308,N_10262,N_11195);
and U12309 (N_12309,N_10215,N_10511);
nor U12310 (N_12310,N_10204,N_10584);
and U12311 (N_12311,N_10030,N_10124);
and U12312 (N_12312,N_9557,N_9546);
xor U12313 (N_12313,N_10449,N_10667);
nor U12314 (N_12314,N_11461,N_11317);
nor U12315 (N_12315,N_10672,N_11819);
xor U12316 (N_12316,N_11626,N_9681);
and U12317 (N_12317,N_9820,N_11435);
nor U12318 (N_12318,N_11616,N_10379);
xnor U12319 (N_12319,N_11296,N_11696);
xor U12320 (N_12320,N_11042,N_11581);
nor U12321 (N_12321,N_10506,N_11888);
nand U12322 (N_12322,N_9699,N_10172);
or U12323 (N_12323,N_11183,N_9025);
xor U12324 (N_12324,N_10349,N_11672);
nor U12325 (N_12325,N_9556,N_9511);
and U12326 (N_12326,N_10709,N_10329);
nand U12327 (N_12327,N_9029,N_9809);
and U12328 (N_12328,N_10817,N_10977);
and U12329 (N_12329,N_10617,N_9307);
or U12330 (N_12330,N_11100,N_9525);
or U12331 (N_12331,N_11628,N_11851);
or U12332 (N_12332,N_9942,N_11018);
and U12333 (N_12333,N_9089,N_10787);
and U12334 (N_12334,N_10203,N_10113);
nand U12335 (N_12335,N_10926,N_9710);
xnor U12336 (N_12336,N_9123,N_11533);
or U12337 (N_12337,N_10991,N_10870);
or U12338 (N_12338,N_11594,N_10947);
nand U12339 (N_12339,N_11661,N_11017);
nor U12340 (N_12340,N_9558,N_9672);
and U12341 (N_12341,N_9674,N_10020);
xor U12342 (N_12342,N_10626,N_11719);
and U12343 (N_12343,N_9239,N_11408);
or U12344 (N_12344,N_9568,N_11253);
or U12345 (N_12345,N_11116,N_9886);
nor U12346 (N_12346,N_10467,N_11632);
or U12347 (N_12347,N_10317,N_11630);
xor U12348 (N_12348,N_9091,N_11254);
nand U12349 (N_12349,N_10374,N_10258);
or U12350 (N_12350,N_9449,N_11613);
and U12351 (N_12351,N_9040,N_9140);
nor U12352 (N_12352,N_11899,N_10902);
and U12353 (N_12353,N_9945,N_9578);
nor U12354 (N_12354,N_9259,N_9833);
and U12355 (N_12355,N_11386,N_10551);
and U12356 (N_12356,N_9334,N_10343);
xnor U12357 (N_12357,N_10595,N_9742);
and U12358 (N_12358,N_11378,N_9154);
and U12359 (N_12359,N_10836,N_11952);
and U12360 (N_12360,N_10829,N_11508);
nand U12361 (N_12361,N_11676,N_11843);
nor U12362 (N_12362,N_9202,N_9372);
nor U12363 (N_12363,N_9236,N_10526);
xnor U12364 (N_12364,N_11742,N_10794);
xor U12365 (N_12365,N_11201,N_9007);
and U12366 (N_12366,N_10557,N_10282);
xnor U12367 (N_12367,N_11220,N_11537);
nand U12368 (N_12368,N_10928,N_11074);
xor U12369 (N_12369,N_10359,N_9644);
nand U12370 (N_12370,N_9478,N_9394);
or U12371 (N_12371,N_11471,N_10694);
nor U12372 (N_12372,N_11223,N_10311);
xor U12373 (N_12373,N_9458,N_11040);
or U12374 (N_12374,N_9547,N_11473);
nor U12375 (N_12375,N_10328,N_9989);
and U12376 (N_12376,N_11919,N_11526);
nand U12377 (N_12377,N_9778,N_10773);
or U12378 (N_12378,N_11565,N_10016);
nand U12379 (N_12379,N_11886,N_10999);
xnor U12380 (N_12380,N_10305,N_11804);
xor U12381 (N_12381,N_10459,N_11327);
nor U12382 (N_12382,N_10922,N_10443);
or U12383 (N_12383,N_10706,N_9861);
xnor U12384 (N_12384,N_9207,N_10714);
xnor U12385 (N_12385,N_9870,N_9623);
or U12386 (N_12386,N_10308,N_9185);
nand U12387 (N_12387,N_9085,N_10679);
nand U12388 (N_12388,N_11070,N_9777);
nor U12389 (N_12389,N_10309,N_11711);
and U12390 (N_12390,N_10461,N_10839);
nor U12391 (N_12391,N_10162,N_9893);
nand U12392 (N_12392,N_10820,N_10208);
and U12393 (N_12393,N_11595,N_10814);
and U12394 (N_12394,N_10039,N_11503);
nand U12395 (N_12395,N_11445,N_11123);
nor U12396 (N_12396,N_11757,N_11624);
xor U12397 (N_12397,N_9760,N_9016);
and U12398 (N_12398,N_10693,N_10715);
and U12399 (N_12399,N_11566,N_10721);
or U12400 (N_12400,N_10542,N_11409);
xor U12401 (N_12401,N_10332,N_9730);
xnor U12402 (N_12402,N_9646,N_9348);
nor U12403 (N_12403,N_9153,N_9727);
and U12404 (N_12404,N_9133,N_9094);
nand U12405 (N_12405,N_9805,N_9139);
or U12406 (N_12406,N_10842,N_11848);
and U12407 (N_12407,N_9138,N_9959);
nand U12408 (N_12408,N_10507,N_11092);
nor U12409 (N_12409,N_10257,N_10403);
xor U12410 (N_12410,N_10347,N_11155);
nor U12411 (N_12411,N_9288,N_9001);
xor U12412 (N_12412,N_9261,N_9633);
and U12413 (N_12413,N_9262,N_10637);
and U12414 (N_12414,N_9589,N_10070);
xor U12415 (N_12415,N_9045,N_10427);
nand U12416 (N_12416,N_11701,N_9567);
or U12417 (N_12417,N_9276,N_10865);
or U12418 (N_12418,N_9356,N_11286);
or U12419 (N_12419,N_11068,N_9024);
xor U12420 (N_12420,N_9829,N_11737);
xnor U12421 (N_12421,N_9043,N_9940);
xnor U12422 (N_12422,N_10571,N_9067);
nand U12423 (N_12423,N_9943,N_9740);
and U12424 (N_12424,N_9108,N_9200);
nand U12425 (N_12425,N_11259,N_9301);
or U12426 (N_12426,N_11172,N_10222);
nor U12427 (N_12427,N_11411,N_11145);
nand U12428 (N_12428,N_9518,N_10850);
nand U12429 (N_12429,N_10394,N_11966);
or U12430 (N_12430,N_10517,N_11452);
or U12431 (N_12431,N_10119,N_11668);
nand U12432 (N_12432,N_11207,N_10553);
nor U12433 (N_12433,N_10770,N_11382);
or U12434 (N_12434,N_9822,N_11239);
and U12435 (N_12435,N_10447,N_10207);
nor U12436 (N_12436,N_9319,N_9537);
or U12437 (N_12437,N_11645,N_11556);
nand U12438 (N_12438,N_11929,N_10192);
and U12439 (N_12439,N_10087,N_10581);
nand U12440 (N_12440,N_11334,N_11956);
nor U12441 (N_12441,N_10761,N_11029);
nand U12442 (N_12442,N_9939,N_9063);
xor U12443 (N_12443,N_9438,N_9280);
nand U12444 (N_12444,N_10896,N_10148);
and U12445 (N_12445,N_11322,N_11833);
or U12446 (N_12446,N_9570,N_11831);
and U12447 (N_12447,N_11470,N_9069);
nor U12448 (N_12448,N_9255,N_10500);
nor U12449 (N_12449,N_9966,N_10568);
nand U12450 (N_12450,N_11525,N_9208);
xor U12451 (N_12451,N_9037,N_10217);
or U12452 (N_12452,N_10136,N_10015);
xor U12453 (N_12453,N_11562,N_10264);
nor U12454 (N_12454,N_11863,N_9009);
and U12455 (N_12455,N_10883,N_11293);
nand U12456 (N_12456,N_10432,N_10518);
and U12457 (N_12457,N_10323,N_9230);
or U12458 (N_12458,N_11363,N_10161);
or U12459 (N_12459,N_11673,N_11304);
nor U12460 (N_12460,N_11896,N_10522);
xnor U12461 (N_12461,N_11841,N_11541);
nand U12462 (N_12462,N_9254,N_10014);
and U12463 (N_12463,N_11861,N_10310);
xnor U12464 (N_12464,N_9019,N_9102);
and U12465 (N_12465,N_9823,N_10587);
xnor U12466 (N_12466,N_9908,N_10352);
or U12467 (N_12467,N_11475,N_11277);
and U12468 (N_12468,N_9603,N_11906);
and U12469 (N_12469,N_9761,N_11967);
xor U12470 (N_12470,N_10069,N_11750);
or U12471 (N_12471,N_11636,N_9892);
and U12472 (N_12472,N_11291,N_9364);
or U12473 (N_12473,N_9756,N_9187);
nand U12474 (N_12474,N_9084,N_10765);
nand U12475 (N_12475,N_10841,N_10649);
nand U12476 (N_12476,N_9643,N_11607);
or U12477 (N_12477,N_9732,N_11777);
nor U12478 (N_12478,N_9437,N_10981);
xor U12479 (N_12479,N_9840,N_10226);
or U12480 (N_12480,N_9279,N_10831);
nand U12481 (N_12481,N_9703,N_11159);
and U12482 (N_12482,N_9450,N_11007);
nand U12483 (N_12483,N_11945,N_11491);
xor U12484 (N_12484,N_11765,N_9628);
and U12485 (N_12485,N_11545,N_11199);
nand U12486 (N_12486,N_10971,N_10849);
nand U12487 (N_12487,N_10952,N_10205);
and U12488 (N_12488,N_9189,N_11684);
xnor U12489 (N_12489,N_9278,N_11480);
xor U12490 (N_12490,N_10278,N_9622);
nor U12491 (N_12491,N_10494,N_10658);
nand U12492 (N_12492,N_9869,N_11046);
and U12493 (N_12493,N_9324,N_9771);
nand U12494 (N_12494,N_11772,N_11570);
and U12495 (N_12495,N_11938,N_11086);
xor U12496 (N_12496,N_9129,N_11084);
and U12497 (N_12497,N_11081,N_11136);
nor U12498 (N_12498,N_9416,N_9735);
nand U12499 (N_12499,N_11131,N_11776);
or U12500 (N_12500,N_9070,N_10027);
nor U12501 (N_12501,N_10277,N_9164);
or U12502 (N_12502,N_11887,N_11026);
xor U12503 (N_12503,N_11258,N_9282);
and U12504 (N_12504,N_9471,N_11756);
nand U12505 (N_12505,N_9387,N_9811);
xor U12506 (N_12506,N_11187,N_10214);
and U12507 (N_12507,N_9163,N_9402);
and U12508 (N_12508,N_11587,N_10984);
nor U12509 (N_12509,N_10102,N_9543);
nand U12510 (N_12510,N_11022,N_9206);
and U12511 (N_12511,N_10319,N_9105);
nor U12512 (N_12512,N_10877,N_10560);
xor U12513 (N_12513,N_9938,N_10139);
or U12514 (N_12514,N_11790,N_11680);
and U12515 (N_12515,N_10572,N_10122);
nand U12516 (N_12516,N_11402,N_9422);
and U12517 (N_12517,N_10579,N_9573);
nor U12518 (N_12518,N_11443,N_11735);
or U12519 (N_12519,N_10625,N_10815);
nand U12520 (N_12520,N_11109,N_10897);
nand U12521 (N_12521,N_9321,N_9034);
xor U12522 (N_12522,N_9510,N_9718);
xor U12523 (N_12523,N_9821,N_10065);
and U12524 (N_12524,N_10885,N_11662);
nor U12525 (N_12525,N_10418,N_10559);
and U12526 (N_12526,N_10930,N_10613);
nand U12527 (N_12527,N_11235,N_9054);
nor U12528 (N_12528,N_10353,N_9951);
and U12529 (N_12529,N_9816,N_11273);
nor U12530 (N_12530,N_10729,N_11492);
xnor U12531 (N_12531,N_11667,N_9311);
nor U12532 (N_12532,N_10996,N_11808);
and U12533 (N_12533,N_11456,N_10103);
or U12534 (N_12534,N_11407,N_10259);
nand U12535 (N_12535,N_11749,N_10167);
and U12536 (N_12536,N_11394,N_9283);
nand U12537 (N_12537,N_9491,N_10662);
or U12538 (N_12538,N_9156,N_11466);
or U12539 (N_12539,N_10395,N_10325);
nor U12540 (N_12540,N_9849,N_11692);
and U12541 (N_12541,N_11489,N_10160);
or U12542 (N_12542,N_11041,N_9323);
xor U12543 (N_12543,N_9711,N_10605);
or U12544 (N_12544,N_9733,N_10610);
nand U12545 (N_12545,N_9784,N_9087);
nand U12546 (N_12546,N_9649,N_11522);
nor U12547 (N_12547,N_10033,N_11824);
nor U12548 (N_12548,N_10096,N_11185);
nor U12549 (N_12549,N_11924,N_10591);
nor U12550 (N_12550,N_9316,N_10966);
xnor U12551 (N_12551,N_10241,N_11779);
xnor U12552 (N_12552,N_9057,N_10297);
and U12553 (N_12553,N_9159,N_10470);
or U12554 (N_12554,N_10338,N_9166);
and U12555 (N_12555,N_11933,N_10574);
and U12556 (N_12556,N_9150,N_9247);
nand U12557 (N_12557,N_9559,N_10512);
or U12558 (N_12558,N_11399,N_11313);
xor U12559 (N_12559,N_10199,N_10601);
or U12560 (N_12560,N_9763,N_10886);
xor U12561 (N_12561,N_11002,N_9420);
xnor U12562 (N_12562,N_10330,N_10252);
nor U12563 (N_12563,N_10633,N_11485);
xor U12564 (N_12564,N_10373,N_10402);
xor U12565 (N_12565,N_11196,N_11114);
and U12566 (N_12566,N_11528,N_11376);
nand U12567 (N_12567,N_10028,N_10387);
nor U12568 (N_12568,N_11034,N_11413);
and U12569 (N_12569,N_9050,N_11917);
xnor U12570 (N_12570,N_9447,N_10967);
nor U12571 (N_12571,N_9632,N_11446);
nor U12572 (N_12572,N_11989,N_11307);
xnor U12573 (N_12573,N_11659,N_11529);
and U12574 (N_12574,N_9047,N_10611);
or U12575 (N_12575,N_11490,N_10320);
or U12576 (N_12576,N_11789,N_10754);
or U12577 (N_12577,N_10092,N_10945);
xnor U12578 (N_12578,N_9577,N_9895);
or U12579 (N_12579,N_10398,N_11056);
or U12580 (N_12580,N_10746,N_9272);
or U12581 (N_12581,N_10012,N_10777);
or U12582 (N_12582,N_11479,N_11907);
xnor U12583 (N_12583,N_10114,N_10233);
or U12584 (N_12584,N_11614,N_9160);
xnor U12585 (N_12585,N_11733,N_9581);
or U12586 (N_12586,N_10193,N_11193);
nand U12587 (N_12587,N_11615,N_11780);
nand U12588 (N_12588,N_11707,N_11393);
or U12589 (N_12589,N_9786,N_10908);
xnor U12590 (N_12590,N_9305,N_11726);
nor U12591 (N_12591,N_9486,N_9788);
xor U12592 (N_12592,N_11970,N_9683);
xnor U12593 (N_12593,N_9368,N_9439);
or U12594 (N_12594,N_11314,N_9848);
nand U12595 (N_12595,N_9937,N_11788);
nand U12596 (N_12596,N_9553,N_9205);
or U12597 (N_12597,N_10000,N_11746);
xnor U12598 (N_12598,N_11342,N_11950);
and U12599 (N_12599,N_9971,N_10213);
nor U12600 (N_12600,N_9252,N_10866);
nor U12601 (N_12601,N_10832,N_9347);
xor U12602 (N_12602,N_10725,N_10742);
nand U12603 (N_12603,N_11530,N_10153);
and U12604 (N_12604,N_10110,N_11604);
nor U12605 (N_12605,N_10757,N_11663);
xnor U12606 (N_12606,N_9304,N_9109);
xnor U12607 (N_12607,N_9446,N_9377);
nor U12608 (N_12608,N_11453,N_10622);
or U12609 (N_12609,N_11335,N_11621);
or U12610 (N_12610,N_10266,N_10699);
nand U12611 (N_12611,N_10949,N_10914);
nand U12612 (N_12612,N_9498,N_11905);
nor U12613 (N_12613,N_11754,N_9036);
nand U12614 (N_12614,N_9629,N_10873);
xor U12615 (N_12615,N_9441,N_9921);
or U12616 (N_12616,N_10474,N_9509);
and U12617 (N_12617,N_10808,N_10844);
xor U12618 (N_12618,N_9924,N_11274);
or U12619 (N_12619,N_9493,N_11242);
nor U12620 (N_12620,N_10890,N_10008);
and U12621 (N_12621,N_10691,N_9576);
xnor U12622 (N_12622,N_11925,N_11454);
nor U12623 (N_12623,N_10918,N_11079);
nand U12624 (N_12624,N_10826,N_9853);
and U12625 (N_12625,N_9171,N_9503);
or U12626 (N_12626,N_9340,N_9618);
nor U12627 (N_12627,N_11025,N_11449);
nand U12628 (N_12628,N_9941,N_11712);
nand U12629 (N_12629,N_9292,N_9506);
nor U12630 (N_12630,N_9807,N_9290);
nor U12631 (N_12631,N_10180,N_11633);
nor U12632 (N_12632,N_11338,N_11133);
nor U12633 (N_12633,N_10548,N_10001);
nand U12634 (N_12634,N_9213,N_9953);
xor U12635 (N_12635,N_11303,N_11354);
nand U12636 (N_12636,N_10006,N_11608);
xor U12637 (N_12637,N_11931,N_11499);
xnor U12638 (N_12638,N_11311,N_10364);
nand U12639 (N_12639,N_10578,N_9268);
or U12640 (N_12640,N_9967,N_11066);
and U12641 (N_12641,N_11510,N_11527);
or U12642 (N_12642,N_9666,N_11915);
and U12643 (N_12643,N_10592,N_9907);
or U12644 (N_12644,N_10979,N_10191);
and U12645 (N_12645,N_10528,N_9417);
or U12646 (N_12646,N_11256,N_10081);
or U12647 (N_12647,N_10576,N_11883);
nand U12648 (N_12648,N_9384,N_10303);
and U12649 (N_12649,N_9062,N_9052);
and U12650 (N_12650,N_9265,N_10872);
nor U12651 (N_12651,N_10741,N_11460);
and U12652 (N_12652,N_10362,N_11889);
nand U12653 (N_12653,N_9060,N_11998);
nor U12654 (N_12654,N_11759,N_10905);
nor U12655 (N_12655,N_9597,N_10855);
xnor U12656 (N_12656,N_10439,N_10972);
or U12657 (N_12657,N_11798,N_11962);
and U12658 (N_12658,N_11854,N_11215);
or U12659 (N_12659,N_9929,N_9531);
nor U12660 (N_12660,N_9545,N_11281);
and U12661 (N_12661,N_11705,N_9079);
nand U12662 (N_12662,N_10811,N_10437);
nand U12663 (N_12663,N_11024,N_10621);
nor U12664 (N_12664,N_10901,N_10657);
xor U12665 (N_12665,N_11072,N_11146);
xnor U12666 (N_12666,N_10485,N_10392);
nand U12667 (N_12667,N_10465,N_9744);
and U12668 (N_12668,N_9026,N_11400);
xor U12669 (N_12669,N_9776,N_9170);
nand U12670 (N_12670,N_10664,N_11868);
or U12671 (N_12671,N_10942,N_10004);
nor U12672 (N_12672,N_10288,N_11973);
and U12673 (N_12673,N_10671,N_11670);
nor U12674 (N_12674,N_9590,N_9630);
or U12675 (N_12675,N_11815,N_11214);
or U12676 (N_12676,N_10295,N_11518);
nand U12677 (N_12677,N_11488,N_10302);
and U12678 (N_12678,N_11971,N_9484);
nor U12679 (N_12679,N_10128,N_9126);
xor U12680 (N_12680,N_10355,N_9619);
nor U12681 (N_12681,N_10962,N_11797);
nor U12682 (N_12682,N_9897,N_11980);
xnor U12683 (N_12683,N_11057,N_9932);
and U12684 (N_12684,N_11734,N_10806);
and U12685 (N_12685,N_11442,N_10838);
nor U12686 (N_12686,N_9930,N_10535);
nor U12687 (N_12687,N_10916,N_11270);
xor U12688 (N_12688,N_11284,N_11450);
nand U12689 (N_12689,N_10602,N_10202);
xor U12690 (N_12690,N_9883,N_10519);
nor U12691 (N_12691,N_9017,N_11006);
and U12692 (N_12692,N_11292,N_10419);
or U12693 (N_12693,N_10060,N_11631);
or U12694 (N_12694,N_11960,N_10112);
nor U12695 (N_12695,N_9260,N_9650);
nand U12696 (N_12696,N_11600,N_10615);
and U12697 (N_12697,N_11816,N_11251);
or U12698 (N_12698,N_9448,N_10290);
xnor U12699 (N_12699,N_11564,N_9743);
nand U12700 (N_12700,N_11583,N_11713);
nand U12701 (N_12701,N_10894,N_11551);
nor U12702 (N_12702,N_11678,N_9151);
or U12703 (N_12703,N_10019,N_9685);
and U12704 (N_12704,N_10740,N_10462);
xnor U12705 (N_12705,N_9122,N_10882);
xor U12706 (N_12706,N_11424,N_9973);
nor U12707 (N_12707,N_10480,N_10749);
or U12708 (N_12708,N_9591,N_9521);
and U12709 (N_12709,N_11972,N_9931);
and U12710 (N_12710,N_10932,N_10431);
and U12711 (N_12711,N_9916,N_10964);
xor U12712 (N_12712,N_9095,N_10185);
nor U12713 (N_12713,N_11532,N_9005);
nand U12714 (N_12714,N_11226,N_9839);
nand U12715 (N_12715,N_9215,N_10510);
nor U12716 (N_12716,N_10155,N_11558);
or U12717 (N_12717,N_9330,N_9353);
nand U12718 (N_12718,N_11189,N_11419);
or U12719 (N_12719,N_9398,N_9678);
or U12720 (N_12720,N_11339,N_10460);
and U12721 (N_12721,N_11352,N_11037);
nor U12722 (N_12722,N_10767,N_11374);
nor U12723 (N_12723,N_9548,N_11852);
or U12724 (N_12724,N_11036,N_9982);
nand U12725 (N_12725,N_11847,N_11646);
or U12726 (N_12726,N_11176,N_9898);
xnor U12727 (N_12727,N_10779,N_10640);
nor U12728 (N_12728,N_10763,N_9826);
or U12729 (N_12729,N_9467,N_11908);
and U12730 (N_12730,N_10244,N_9762);
and U12731 (N_12731,N_11622,N_10686);
or U12732 (N_12732,N_10380,N_10314);
nand U12733 (N_12733,N_11358,N_11429);
and U12734 (N_12734,N_11791,N_11584);
nand U12735 (N_12735,N_9783,N_10661);
nor U12736 (N_12736,N_9997,N_10477);
or U12737 (N_12737,N_10234,N_10369);
nor U12738 (N_12738,N_10778,N_10974);
and U12739 (N_12739,N_9426,N_10062);
and U12740 (N_12740,N_11147,N_10921);
or U12741 (N_12741,N_9750,N_11379);
or U12742 (N_12742,N_9599,N_11918);
xnor U12743 (N_12743,N_9804,N_10186);
and U12744 (N_12744,N_9957,N_10804);
nor U12745 (N_12745,N_9176,N_10884);
xor U12746 (N_12746,N_10478,N_11275);
xor U12747 (N_12747,N_11099,N_9128);
nand U12748 (N_12748,N_9514,N_10813);
nor U12749 (N_12749,N_10166,N_11892);
nand U12750 (N_12750,N_9162,N_10170);
nor U12751 (N_12751,N_10017,N_9598);
or U12752 (N_12752,N_10438,N_11801);
nand U12753 (N_12753,N_9038,N_9382);
xnor U12754 (N_12754,N_11422,N_11715);
nand U12755 (N_12755,N_10710,N_9114);
nor U12756 (N_12756,N_9231,N_11117);
nor U12757 (N_12757,N_11913,N_11050);
or U12758 (N_12758,N_9197,N_10948);
nor U12759 (N_12759,N_10195,N_11714);
xnor U12760 (N_12760,N_9555,N_11312);
nand U12761 (N_12761,N_9313,N_10029);
nor U12762 (N_12762,N_9722,N_10083);
xor U12763 (N_12763,N_9031,N_9954);
nor U12764 (N_12764,N_11605,N_11014);
xnor U12765 (N_12765,N_11430,N_9601);
nand U12766 (N_12766,N_10868,N_9104);
nor U12767 (N_12767,N_11289,N_9728);
nand U12768 (N_12768,N_11606,N_9469);
or U12769 (N_12769,N_10118,N_11218);
xnor U12770 (N_12770,N_9403,N_9293);
nand U12771 (N_12771,N_9701,N_10411);
xnor U12772 (N_12772,N_10569,N_11703);
nor U12773 (N_12773,N_11725,N_9550);
nand U12774 (N_12774,N_10097,N_10423);
nand U12775 (N_12775,N_11894,N_10009);
xor U12776 (N_12776,N_9186,N_10851);
and U12777 (N_12777,N_11560,N_9700);
or U12778 (N_12778,N_9175,N_10466);
nor U12779 (N_12779,N_11957,N_11428);
xnor U12780 (N_12780,N_9190,N_9179);
nor U12781 (N_12781,N_10707,N_9226);
and U12782 (N_12782,N_10149,N_10531);
or U12783 (N_12783,N_9752,N_11065);
xnor U12784 (N_12784,N_9119,N_9605);
nor U12785 (N_12785,N_10869,N_11178);
nor U12786 (N_12786,N_11455,N_9517);
and U12787 (N_12787,N_10291,N_11398);
nand U12788 (N_12788,N_11384,N_10123);
or U12789 (N_12789,N_11505,N_9911);
or U12790 (N_12790,N_11168,N_9404);
nand U12791 (N_12791,N_10005,N_11069);
xor U12792 (N_12792,N_9474,N_11623);
nand U12793 (N_12793,N_10484,N_9874);
xor U12794 (N_12794,N_10390,N_11467);
xnor U12795 (N_12795,N_11320,N_9362);
or U12796 (N_12796,N_11988,N_9987);
nand U12797 (N_12797,N_9857,N_9376);
nor U12798 (N_12798,N_9267,N_10618);
nand U12799 (N_12799,N_9798,N_11406);
nand U12800 (N_12800,N_11825,N_9552);
and U12801 (N_12801,N_9451,N_9996);
or U12802 (N_12802,N_10830,N_9078);
nand U12803 (N_12803,N_11137,N_9059);
and U12804 (N_12804,N_9831,N_10650);
xnor U12805 (N_12805,N_9465,N_9149);
and U12806 (N_12806,N_11448,N_10152);
xnor U12807 (N_12807,N_11738,N_10846);
and U12808 (N_12808,N_11955,N_11949);
nor U12809 (N_12809,N_11027,N_9968);
nand U12810 (N_12810,N_10853,N_9797);
xnor U12811 (N_12811,N_11860,N_11729);
nand U12812 (N_12812,N_9575,N_10992);
nand U12813 (N_12813,N_11800,N_11891);
nor U12814 (N_12814,N_11383,N_11864);
xnor U12815 (N_12815,N_11552,N_9533);
nand U12816 (N_12816,N_10368,N_11850);
nor U12817 (N_12817,N_9507,N_10562);
and U12818 (N_12818,N_11890,N_10492);
xor U12819 (N_12819,N_10281,N_10933);
xor U12820 (N_12820,N_9990,N_9112);
or U12821 (N_12821,N_11698,N_11325);
nor U12822 (N_12822,N_9068,N_10847);
nor U12823 (N_12823,N_9679,N_9411);
xor U12824 (N_12824,N_9371,N_10322);
and U12825 (N_12825,N_9961,N_10614);
nand U12826 (N_12826,N_9858,N_10071);
and U12827 (N_12827,N_9834,N_10146);
and U12828 (N_12828,N_9901,N_9505);
nor U12829 (N_12829,N_10703,N_10532);
or U12830 (N_12830,N_9386,N_9536);
and U12831 (N_12831,N_10643,N_10816);
xnor U12832 (N_12832,N_9008,N_11237);
xnor U12833 (N_12833,N_10134,N_10834);
or U12834 (N_12834,N_11229,N_11953);
and U12835 (N_12835,N_11839,N_9295);
and U12836 (N_12836,N_9787,N_10735);
and U12837 (N_12837,N_11814,N_9586);
nand U12838 (N_12838,N_11360,N_10704);
and U12839 (N_12839,N_9241,N_11468);
and U12840 (N_12840,N_9894,N_10646);
or U12841 (N_12841,N_11981,N_10504);
xor U12842 (N_12842,N_10862,N_11760);
xnor U12843 (N_12843,N_9039,N_10656);
nand U12844 (N_12844,N_10356,N_11225);
and U12845 (N_12845,N_9675,N_11154);
and U12846 (N_12846,N_9328,N_11213);
xor U12847 (N_12847,N_11964,N_11088);
or U12848 (N_12848,N_9528,N_9868);
xnor U12849 (N_12849,N_11637,N_10294);
and U12850 (N_12850,N_11171,N_9970);
nand U12851 (N_12851,N_10120,N_10301);
and U12852 (N_12852,N_10189,N_11090);
nor U12853 (N_12853,N_11324,N_9721);
and U12854 (N_12854,N_9476,N_9488);
nor U12855 (N_12855,N_10733,N_9434);
nor U12856 (N_12856,N_11228,N_9799);
nand U12857 (N_12857,N_9844,N_9223);
and U12858 (N_12858,N_9214,N_11916);
and U12859 (N_12859,N_9562,N_10142);
nor U12860 (N_12860,N_10780,N_11775);
or U12861 (N_12861,N_11495,N_9400);
xor U12862 (N_12862,N_10354,N_9291);
nor U12863 (N_12863,N_9707,N_11783);
xor U12864 (N_12864,N_9132,N_10361);
and U12865 (N_12865,N_11786,N_9774);
or U12866 (N_12866,N_10416,N_10367);
and U12867 (N_12867,N_11369,N_9250);
and U12868 (N_12868,N_11052,N_9817);
nor U12869 (N_12869,N_11104,N_10786);
xnor U12870 (N_12870,N_11285,N_10944);
nor U12871 (N_12871,N_10464,N_11827);
xnor U12872 (N_12872,N_10440,N_9615);
and U12873 (N_12873,N_10132,N_10475);
nor U12874 (N_12874,N_11184,N_11245);
nand U12875 (N_12875,N_11381,N_11809);
nor U12876 (N_12876,N_11762,N_10946);
nor U12877 (N_12877,N_9314,N_11837);
xor U12878 (N_12878,N_10131,N_10958);
and U12879 (N_12879,N_11366,N_10638);
nor U12880 (N_12880,N_9995,N_11433);
nand U12881 (N_12881,N_11795,N_9413);
nand U12882 (N_12882,N_10547,N_9885);
or U12883 (N_12883,N_11596,N_9147);
and U12884 (N_12884,N_10871,N_11651);
xor U12885 (N_12885,N_9118,N_11333);
or U12886 (N_12886,N_9194,N_9527);
nand U12887 (N_12887,N_10101,N_11747);
or U12888 (N_12888,N_11770,N_11013);
or U12889 (N_12889,N_9994,N_11927);
nand U12890 (N_12890,N_9810,N_9174);
or U12891 (N_12891,N_10090,N_10127);
or U12892 (N_12892,N_10797,N_11107);
xnor U12893 (N_12893,N_11862,N_9782);
and U12894 (N_12894,N_9793,N_9694);
and U12895 (N_12895,N_10756,N_11410);
xor U12896 (N_12896,N_11602,N_10705);
or U12897 (N_12897,N_10472,N_10812);
xnor U12898 (N_12898,N_11085,N_10072);
nor U12899 (N_12899,N_11716,N_9145);
xnor U12900 (N_12900,N_11175,N_11994);
nand U12901 (N_12901,N_9173,N_9785);
and U12902 (N_12902,N_11368,N_11112);
xor U12903 (N_12903,N_9483,N_10744);
nor U12904 (N_12904,N_10961,N_9432);
or U12905 (N_12905,N_11063,N_9920);
or U12906 (N_12906,N_9076,N_9042);
or U12907 (N_12907,N_11272,N_11764);
or U12908 (N_12908,N_9862,N_9106);
and U12909 (N_12909,N_9373,N_10597);
xor U12910 (N_12910,N_11377,N_11849);
nor U12911 (N_12911,N_11125,N_11752);
nand U12912 (N_12912,N_9906,N_11103);
xor U12913 (N_12913,N_11128,N_10496);
nor U12914 (N_12914,N_11416,N_10429);
or U12915 (N_12915,N_9056,N_10350);
and U12916 (N_12916,N_9274,N_9928);
xnor U12917 (N_12917,N_11015,N_10054);
nand U12918 (N_12918,N_11838,N_11330);
or U12919 (N_12919,N_11590,N_11657);
nand U12920 (N_12920,N_11666,N_11813);
and U12921 (N_12921,N_10795,N_9203);
or U12922 (N_12922,N_11543,N_9117);
or U12923 (N_12923,N_9022,N_9872);
nor U12924 (N_12924,N_10151,N_10644);
or U12925 (N_12925,N_9308,N_11610);
or U12926 (N_12926,N_10287,N_11132);
or U12927 (N_12927,N_11878,N_11599);
nand U12928 (N_12928,N_11158,N_10445);
xor U12929 (N_12929,N_10858,N_10061);
or U12930 (N_12930,N_11236,N_11297);
and U12931 (N_12931,N_11648,N_10860);
nor U12932 (N_12932,N_10585,N_11803);
or U12933 (N_12933,N_9086,N_9044);
or U12934 (N_12934,N_9664,N_10732);
or U12935 (N_12935,N_9983,N_11840);
nor U12936 (N_12936,N_9565,N_10201);
nor U12937 (N_12937,N_11162,N_11387);
xnor U12938 (N_12938,N_11778,N_11098);
nand U12939 (N_12939,N_11302,N_10998);
xor U12940 (N_12940,N_9237,N_9326);
nand U12941 (N_12941,N_10533,N_9758);
xor U12942 (N_12942,N_9642,N_9367);
or U12943 (N_12943,N_10424,N_11250);
nand U12944 (N_12944,N_10344,N_9978);
nor U12945 (N_12945,N_11140,N_9659);
and U12946 (N_12946,N_9199,N_11441);
nand U12947 (N_12947,N_9780,N_9337);
nand U12948 (N_12948,N_10457,N_9336);
or U12949 (N_12949,N_11538,N_9613);
nand U12950 (N_12950,N_11150,N_10013);
or U12951 (N_12951,N_10629,N_9299);
nor U12952 (N_12952,N_9234,N_11141);
xnor U12953 (N_12953,N_11059,N_10388);
or U12954 (N_12954,N_11486,N_11909);
or U12955 (N_12955,N_10880,N_9827);
or U12956 (N_12956,N_11144,N_10687);
nand U12957 (N_12957,N_9101,N_11494);
or U12958 (N_12958,N_9161,N_9180);
nor U12959 (N_12959,N_10231,N_10299);
or U12960 (N_12960,N_9720,N_10209);
or U12961 (N_12961,N_11942,N_9051);
and U12962 (N_12962,N_9956,N_11589);
and U12963 (N_12963,N_10743,N_9092);
xnor U12964 (N_12964,N_10590,N_10126);
nand U12965 (N_12965,N_9381,N_11873);
nor U12966 (N_12966,N_11869,N_9690);
xnor U12967 (N_12967,N_11655,N_10566);
and U12968 (N_12968,N_10495,N_10268);
nor U12969 (N_12969,N_11227,N_10782);
nor U12970 (N_12970,N_11115,N_10129);
nand U12971 (N_12971,N_10940,N_11690);
xnor U12972 (N_12972,N_10463,N_11921);
nor U12973 (N_12973,N_9329,N_9676);
xor U12974 (N_12974,N_10306,N_11021);
or U12975 (N_12975,N_9726,N_11572);
or U12976 (N_12976,N_9836,N_11968);
or U12977 (N_12977,N_11753,N_9922);
xor U12978 (N_12978,N_10393,N_9395);
xor U12979 (N_12979,N_9881,N_9653);
nand U12980 (N_12980,N_10688,N_10867);
nand U12981 (N_12981,N_9748,N_11261);
nand U12982 (N_12982,N_9934,N_10986);
nor U12983 (N_12983,N_10279,N_9366);
xnor U12984 (N_12984,N_10575,N_10973);
and U12985 (N_12985,N_10580,N_9946);
and U12986 (N_12986,N_9490,N_9481);
or U12987 (N_12987,N_9806,N_11208);
nor U12988 (N_12988,N_10750,N_10022);
nor U12989 (N_12989,N_10488,N_9723);
or U12990 (N_12990,N_11385,N_10570);
xnor U12991 (N_12991,N_9201,N_9610);
and U12992 (N_12992,N_9952,N_9779);
nand U12993 (N_12993,N_10242,N_11295);
nor U12994 (N_12994,N_9421,N_11881);
or U12995 (N_12995,N_11904,N_9677);
nor U12996 (N_12996,N_9655,N_10774);
and U12997 (N_12997,N_11469,N_10254);
and U12998 (N_12998,N_10337,N_11047);
nor U12999 (N_12999,N_10219,N_9263);
xnor U13000 (N_13000,N_9635,N_11910);
or U13001 (N_13001,N_11405,N_9012);
nor U13002 (N_13002,N_10340,N_10917);
nor U13003 (N_13003,N_10583,N_10243);
and U13004 (N_13004,N_9841,N_9284);
xnor U13005 (N_13005,N_9497,N_9981);
xor U13006 (N_13006,N_11391,N_9193);
nand U13007 (N_13007,N_10421,N_9343);
and U13008 (N_13008,N_9405,N_9668);
nor U13009 (N_13009,N_9242,N_9015);
xor U13010 (N_13010,N_10107,N_9332);
nand U13011 (N_13011,N_10909,N_9691);
or U13012 (N_13012,N_10776,N_10399);
nor U13013 (N_13013,N_9814,N_9475);
or U13014 (N_13014,N_11723,N_10476);
xor U13015 (N_13015,N_10893,N_9935);
nor U13016 (N_13016,N_9298,N_11740);
nor U13017 (N_13017,N_11744,N_11535);
nand U13018 (N_13018,N_11210,N_10138);
nand U13019 (N_13019,N_11262,N_11255);
and U13020 (N_13020,N_10864,N_11351);
nor U13021 (N_13021,N_11932,N_10549);
or U13022 (N_13022,N_9379,N_10223);
xnor U13023 (N_13023,N_9731,N_11058);
and U13024 (N_13024,N_10280,N_9972);
and U13025 (N_13025,N_11067,N_11234);
and U13026 (N_13026,N_10371,N_9686);
nand U13027 (N_13027,N_9099,N_11361);
xor U13028 (N_13028,N_11279,N_11373);
xnor U13029 (N_13029,N_9135,N_11524);
and U13030 (N_13030,N_11375,N_10137);
nand U13031 (N_13031,N_11126,N_11481);
or U13032 (N_13032,N_10677,N_9168);
nor U13033 (N_13033,N_10376,N_10037);
nor U13034 (N_13034,N_9496,N_9443);
nand U13035 (N_13035,N_9682,N_9221);
nand U13036 (N_13036,N_11010,N_9216);
and U13037 (N_13037,N_9764,N_10722);
nor U13038 (N_13038,N_9212,N_10630);
or U13039 (N_13039,N_11243,N_9066);
and U13040 (N_13040,N_10451,N_10598);
xnor U13041 (N_13041,N_10541,N_10436);
nand U13042 (N_13042,N_9320,N_11743);
or U13043 (N_13043,N_11434,N_10406);
nor U13044 (N_13044,N_9142,N_11169);
nand U13045 (N_13045,N_9219,N_10976);
or U13046 (N_13046,N_11920,N_11773);
or U13047 (N_13047,N_10143,N_9535);
or U13048 (N_13048,N_9341,N_9120);
xor U13049 (N_13049,N_11823,N_11818);
or U13050 (N_13050,N_10365,N_11031);
nor U13051 (N_13051,N_10256,N_11983);
or U13052 (N_13052,N_10183,N_10737);
or U13053 (N_13053,N_11221,N_11288);
xnor U13054 (N_13054,N_9472,N_10210);
or U13055 (N_13055,N_10481,N_10175);
or U13056 (N_13056,N_9616,N_9984);
or U13057 (N_13057,N_11135,N_11515);
nor U13058 (N_13058,N_11345,N_11822);
nor U13059 (N_13059,N_10953,N_10792);
nor U13060 (N_13060,N_11039,N_9083);
nand U13061 (N_13061,N_10505,N_11267);
nand U13062 (N_13062,N_10833,N_9851);
and U13063 (N_13063,N_9333,N_10360);
nor U13064 (N_13064,N_10417,N_9312);
and U13065 (N_13065,N_9662,N_9082);
nor U13066 (N_13066,N_11440,N_9767);
xnor U13067 (N_13067,N_10187,N_9915);
or U13068 (N_13068,N_10678,N_9354);
or U13069 (N_13069,N_11954,N_11298);
or U13070 (N_13070,N_9494,N_11241);
or U13071 (N_13071,N_11568,N_10563);
or U13072 (N_13072,N_10265,N_9670);
or U13073 (N_13073,N_11300,N_9539);
nand U13074 (N_13074,N_10455,N_10856);
xnor U13075 (N_13075,N_11194,N_10135);
nand U13076 (N_13076,N_10051,N_11991);
xnor U13077 (N_13077,N_11934,N_11247);
xor U13078 (N_13078,N_9582,N_9847);
and U13079 (N_13079,N_11554,N_10995);
xor U13080 (N_13080,N_9900,N_11693);
nand U13081 (N_13081,N_11785,N_9745);
nand U13082 (N_13082,N_9396,N_9532);
xor U13083 (N_13083,N_9232,N_11948);
nor U13084 (N_13084,N_11669,N_10384);
nor U13085 (N_13085,N_11999,N_10400);
nand U13086 (N_13086,N_10047,N_11462);
xor U13087 (N_13087,N_9986,N_11355);
and U13088 (N_13088,N_9257,N_10003);
xor U13089 (N_13089,N_9749,N_10383);
xnor U13090 (N_13090,N_11326,N_11642);
nand U13091 (N_13091,N_9824,N_10516);
and U13092 (N_13092,N_9842,N_10099);
xnor U13093 (N_13093,N_10245,N_11871);
or U13094 (N_13094,N_10165,N_9074);
nor U13095 (N_13095,N_10358,N_9903);
or U13096 (N_13096,N_11396,N_11829);
nand U13097 (N_13097,N_10458,N_11977);
nor U13098 (N_13098,N_9182,N_10919);
nand U13099 (N_13099,N_10950,N_11343);
nand U13100 (N_13100,N_10498,N_11856);
xnor U13101 (N_13101,N_10903,N_11944);
or U13102 (N_13102,N_9018,N_10728);
or U13103 (N_13103,N_9177,N_11611);
xor U13104 (N_13104,N_9835,N_10556);
and U13105 (N_13105,N_10089,N_10594);
and U13106 (N_13106,N_10100,N_10666);
nor U13107 (N_13107,N_10491,N_11876);
or U13108 (N_13108,N_10293,N_11216);
and U13109 (N_13109,N_9566,N_10983);
nand U13110 (N_13110,N_10720,N_9310);
nand U13111 (N_13111,N_11897,N_11502);
xnor U13112 (N_13112,N_9754,N_11044);
or U13113 (N_13113,N_9152,N_9431);
nand U13114 (N_13114,N_11346,N_11190);
nor U13115 (N_13115,N_11730,N_11627);
nand U13116 (N_13116,N_9960,N_11080);
nor U13117 (N_13117,N_9004,N_11542);
xnor U13118 (N_13118,N_9837,N_11349);
nand U13119 (N_13119,N_10840,N_10444);
xnor U13120 (N_13120,N_11969,N_10805);
and U13121 (N_13121,N_9739,N_9741);
xor U13122 (N_13122,N_9385,N_11603);
nor U13123 (N_13123,N_10670,N_11877);
and U13124 (N_13124,N_9564,N_11805);
and U13125 (N_13125,N_9462,N_9501);
and U13126 (N_13126,N_10726,N_10357);
nor U13127 (N_13127,N_11845,N_9689);
xnor U13128 (N_13128,N_9399,N_9271);
and U13129 (N_13129,N_11487,N_9596);
nor U13130 (N_13130,N_10212,N_11465);
nor U13131 (N_13131,N_10738,N_9000);
and U13132 (N_13132,N_10190,N_10075);
nor U13133 (N_13133,N_10227,N_11012);
or U13134 (N_13134,N_10493,N_11353);
nand U13135 (N_13135,N_10108,N_11477);
or U13136 (N_13136,N_10712,N_11574);
or U13137 (N_13137,N_10448,N_9889);
or U13138 (N_13138,N_9442,N_9137);
or U13139 (N_13139,N_9855,N_9245);
nand U13140 (N_13140,N_11586,N_10324);
nand U13141 (N_13141,N_11997,N_11858);
xnor U13142 (N_13142,N_10442,N_10923);
or U13143 (N_13143,N_10674,N_9714);
nand U13144 (N_13144,N_11975,N_11993);
nor U13145 (N_13145,N_9436,N_10843);
and U13146 (N_13146,N_10854,N_10068);
and U13147 (N_13147,N_9482,N_9355);
nor U13148 (N_13148,N_11935,N_10717);
nand U13149 (N_13149,N_9048,N_10716);
nor U13150 (N_13150,N_9887,N_10372);
nand U13151 (N_13151,N_9419,N_9309);
and U13152 (N_13152,N_10228,N_10668);
nand U13153 (N_13153,N_10236,N_11867);
or U13154 (N_13154,N_10469,N_11372);
or U13155 (N_13155,N_11576,N_11260);
and U13156 (N_13156,N_10304,N_11143);
and U13157 (N_13157,N_11371,N_11423);
nor U13158 (N_13158,N_10673,N_9080);
and U13159 (N_13159,N_10527,N_11093);
or U13160 (N_13160,N_9072,N_9639);
and U13161 (N_13161,N_9116,N_11106);
nand U13162 (N_13162,N_10117,N_9111);
nand U13163 (N_13163,N_9992,N_9585);
xor U13164 (N_13164,N_10723,N_11458);
and U13165 (N_13165,N_11222,N_11965);
xor U13166 (N_13166,N_11436,N_11028);
nor U13167 (N_13167,N_10558,N_11656);
xor U13168 (N_13168,N_11276,N_11403);
and U13169 (N_13169,N_11511,N_11926);
nand U13170 (N_13170,N_10681,N_11389);
or U13171 (N_13171,N_10652,N_10497);
nor U13172 (N_13172,N_10283,N_10409);
and U13173 (N_13173,N_11694,N_10990);
and U13174 (N_13174,N_11008,N_11219);
nand U13175 (N_13175,N_9988,N_10878);
nand U13176 (N_13176,N_11102,N_11138);
nand U13177 (N_13177,N_10171,N_10053);
xor U13178 (N_13178,N_10450,N_10937);
nor U13179 (N_13179,N_10049,N_11167);
nand U13180 (N_13180,N_11457,N_10781);
nand U13181 (N_13181,N_11617,N_10334);
and U13182 (N_13182,N_10141,N_10024);
or U13183 (N_13183,N_11523,N_9654);
nand U13184 (N_13184,N_9224,N_11557);
and U13185 (N_13185,N_11685,N_9289);
nand U13186 (N_13186,N_9693,N_9625);
nor U13187 (N_13187,N_11674,N_9671);
nor U13188 (N_13188,N_9688,N_11280);
nand U13189 (N_13189,N_9418,N_9270);
or U13190 (N_13190,N_11578,N_11911);
nor U13191 (N_13191,N_9673,N_9882);
nor U13192 (N_13192,N_11727,N_11152);
xnor U13193 (N_13193,N_10468,N_9753);
nor U13194 (N_13194,N_11501,N_11091);
nor U13195 (N_13195,N_11635,N_11507);
and U13196 (N_13196,N_11817,N_11248);
or U13197 (N_13197,N_10307,N_10898);
nand U13198 (N_13198,N_9433,N_11319);
and U13199 (N_13199,N_9747,N_9526);
nand U13200 (N_13200,N_10453,N_11005);
nand U13201 (N_13201,N_9791,N_9196);
nand U13202 (N_13202,N_9704,N_11940);
nand U13203 (N_13203,N_10600,N_9890);
nand U13204 (N_13204,N_9607,N_10955);
nand U13205 (N_13205,N_11721,N_10561);
or U13206 (N_13206,N_9867,N_9317);
or U13207 (N_13207,N_10412,N_11157);
nand U13208 (N_13208,N_11947,N_10271);
xor U13209 (N_13209,N_9542,N_9692);
and U13210 (N_13210,N_10546,N_10067);
and U13211 (N_13211,N_10627,N_11710);
and U13212 (N_13212,N_9850,N_11987);
and U13213 (N_13213,N_10064,N_10339);
or U13214 (N_13214,N_11575,N_9020);
nand U13215 (N_13215,N_11444,N_9227);
or U13216 (N_13216,N_9614,N_10925);
xor U13217 (N_13217,N_11700,N_9053);
xor U13218 (N_13218,N_10401,N_11943);
xnor U13219 (N_13219,N_10544,N_11836);
and U13220 (N_13220,N_11426,N_11893);
and U13221 (N_13221,N_11885,N_10145);
xnor U13222 (N_13222,N_11638,N_10389);
and U13223 (N_13223,N_11166,N_11996);
xor U13224 (N_13224,N_9211,N_10892);
or U13225 (N_13225,N_9246,N_9800);
and U13226 (N_13226,N_10889,N_10063);
xor U13227 (N_13227,N_9006,N_10935);
and U13228 (N_13228,N_10920,N_9064);
xor U13229 (N_13229,N_9296,N_10565);
nand U13230 (N_13230,N_10157,N_10154);
and U13231 (N_13231,N_10490,N_10147);
nor U13232 (N_13232,N_9569,N_11796);
and U13233 (N_13233,N_9253,N_10093);
nor U13234 (N_13234,N_11832,N_11283);
nor U13235 (N_13235,N_9651,N_9415);
nand U13236 (N_13236,N_11978,N_10791);
and U13237 (N_13237,N_9944,N_11177);
or U13238 (N_13238,N_9339,N_10731);
and U13239 (N_13239,N_9383,N_9281);
xor U13240 (N_13240,N_9725,N_10428);
and U13241 (N_13241,N_9453,N_9228);
nand U13242 (N_13242,N_11427,N_9098);
nand U13243 (N_13243,N_11619,N_11212);
nand U13244 (N_13244,N_9096,N_10772);
or U13245 (N_13245,N_9561,N_11974);
and U13246 (N_13246,N_9401,N_11105);
or U13247 (N_13247,N_11580,N_10285);
and U13248 (N_13248,N_11675,N_11882);
xor U13249 (N_13249,N_10701,N_10682);
nand U13250 (N_13250,N_9790,N_10713);
or U13251 (N_13251,N_10026,N_11767);
or U13252 (N_13252,N_9519,N_11514);
nand U13253 (N_13253,N_10158,N_10881);
and U13254 (N_13254,N_9926,N_11912);
or U13255 (N_13255,N_11238,N_9240);
and U13256 (N_13256,N_10606,N_10182);
xnor U13257 (N_13257,N_11004,N_9656);
nor U13258 (N_13258,N_11287,N_9238);
xnor U13259 (N_13259,N_11230,N_11553);
xor U13260 (N_13260,N_9717,N_11506);
and U13261 (N_13261,N_9636,N_9103);
nand U13262 (N_13262,N_11946,N_10269);
or U13263 (N_13263,N_11032,N_10957);
xor U13264 (N_13264,N_9169,N_9877);
nor U13265 (N_13265,N_10080,N_9172);
or U13266 (N_13266,N_10968,N_11866);
nand U13267 (N_13267,N_9899,N_11939);
nor U13268 (N_13268,N_9684,N_11567);
nor U13269 (N_13269,N_10246,N_10348);
xnor U13270 (N_13270,N_9165,N_9480);
xor U13271 (N_13271,N_9665,N_9878);
or U13272 (N_13272,N_9781,N_11438);
nand U13273 (N_13273,N_10931,N_10487);
nor U13274 (N_13274,N_11563,N_10771);
nand U13275 (N_13275,N_10801,N_11033);
and U13276 (N_13276,N_10156,N_10370);
and U13277 (N_13277,N_11498,N_11357);
nor U13278 (N_13278,N_11771,N_9755);
nor U13279 (N_13279,N_10543,N_11202);
and U13280 (N_13280,N_9188,N_11075);
nor U13281 (N_13281,N_11683,N_11900);
nor U13282 (N_13282,N_10499,N_11459);
or U13283 (N_13283,N_11082,N_10891);
xor U13284 (N_13284,N_9127,N_9766);
xor U13285 (N_13285,N_10116,N_11476);
xor U13286 (N_13286,N_10620,N_11902);
and U13287 (N_13287,N_11336,N_10218);
and U13288 (N_13288,N_11769,N_11828);
nor U13289 (N_13289,N_11203,N_9477);
nand U13290 (N_13290,N_10696,N_11513);
xnor U13291 (N_13291,N_10534,N_11482);
xnor U13292 (N_13292,N_11316,N_11051);
or U13293 (N_13293,N_10375,N_10085);
xnor U13294 (N_13294,N_9792,N_10405);
nor U13295 (N_13295,N_9838,N_10993);
or U13296 (N_13296,N_11591,N_9322);
or U13297 (N_13297,N_9523,N_10174);
nor U13298 (N_13298,N_9856,N_9244);
xor U13299 (N_13299,N_11979,N_11483);
and U13300 (N_13300,N_9375,N_11209);
nor U13301 (N_13301,N_9358,N_9608);
or U13302 (N_13302,N_11976,N_11835);
xor U13303 (N_13303,N_11751,N_11246);
nor U13304 (N_13304,N_9697,N_10523);
or U13305 (N_13305,N_11217,N_9013);
or U13306 (N_13306,N_11332,N_11793);
and U13307 (N_13307,N_10641,N_9468);
nor U13308 (N_13308,N_11928,N_11110);
nand U13309 (N_13309,N_9592,N_9584);
nor U13310 (N_13310,N_9913,N_10177);
or U13311 (N_13311,N_9370,N_9657);
nand U13312 (N_13312,N_9948,N_10188);
or U13313 (N_13313,N_10802,N_9406);
nand U13314 (N_13314,N_10985,N_10810);
nor U13315 (N_13315,N_9338,N_9217);
or U13316 (N_13316,N_10316,N_10289);
nand U13317 (N_13317,N_10043,N_9032);
and U13318 (N_13318,N_11224,N_10248);
nor U13319 (N_13319,N_11252,N_10609);
nor U13320 (N_13320,N_9264,N_11153);
nor U13321 (N_13321,N_10397,N_10654);
and U13322 (N_13322,N_11547,N_10988);
xor U13323 (N_13323,N_11739,N_9859);
xnor U13324 (N_13324,N_11173,N_10196);
nand U13325 (N_13325,N_9430,N_9515);
and U13326 (N_13326,N_9904,N_9602);
nand U13327 (N_13327,N_10286,N_9947);
nand U13328 (N_13328,N_10501,N_11689);
and U13329 (N_13329,N_10425,N_10784);
or U13330 (N_13330,N_9919,N_9593);
nand U13331 (N_13331,N_11898,N_9888);
nand U13332 (N_13332,N_10845,N_11420);
nor U13333 (N_13333,N_11299,N_10651);
or U13334 (N_13334,N_10680,N_9538);
or U13335 (N_13335,N_11180,N_11130);
xnor U13336 (N_13336,N_10915,N_10635);
and U13337 (N_13337,N_9775,N_11000);
xnor U13338 (N_13338,N_9529,N_11038);
nand U13339 (N_13339,N_11745,N_9958);
or U13340 (N_13340,N_10608,N_10007);
or U13341 (N_13341,N_11844,N_11588);
and U13342 (N_13342,N_11348,N_9540);
xor U13343 (N_13343,N_11120,N_11612);
nor U13344 (N_13344,N_9463,N_10540);
nand U13345 (N_13345,N_9435,N_11323);
and U13346 (N_13346,N_10675,N_10900);
and U13347 (N_13347,N_9414,N_9695);
xor U13348 (N_13348,N_10798,N_11875);
or U13349 (N_13349,N_9181,N_11412);
nor U13350 (N_13350,N_10951,N_9769);
nor U13351 (N_13351,N_10564,N_10552);
nand U13352 (N_13352,N_10660,N_10041);
or U13353 (N_13353,N_9489,N_9021);
and U13354 (N_13354,N_10452,N_9195);
nand U13355 (N_13355,N_11859,N_9479);
nor U13356 (N_13356,N_10159,N_11142);
or U13357 (N_13357,N_9090,N_9229);
xnor U13358 (N_13358,N_9815,N_9473);
nand U13359 (N_13359,N_9969,N_9183);
or U13360 (N_13360,N_9107,N_11516);
nor U13361 (N_13361,N_9544,N_9046);
xor U13362 (N_13362,N_11011,N_11549);
nor U13363 (N_13363,N_9049,N_9178);
or U13364 (N_13364,N_11077,N_10140);
nand U13365 (N_13365,N_10685,N_10274);
or U13366 (N_13366,N_11519,N_10094);
and U13367 (N_13367,N_9287,N_10538);
nor U13368 (N_13368,N_9412,N_11053);
nand U13369 (N_13369,N_11101,N_10225);
and U13370 (N_13370,N_10038,N_11451);
nand U13371 (N_13371,N_11857,N_9452);
nand U13372 (N_13372,N_11761,N_9303);
or U13373 (N_13373,N_9516,N_11414);
nor U13374 (N_13374,N_10959,N_11390);
nand U13375 (N_13375,N_11842,N_10168);
nand U13376 (N_13376,N_9680,N_11257);
nor U13377 (N_13377,N_9645,N_11164);
nor U13378 (N_13378,N_11741,N_10250);
xor U13379 (N_13379,N_9914,N_9950);
and U13380 (N_13380,N_9884,N_11629);
or U13381 (N_13381,N_9131,N_10176);
xnor U13382 (N_13382,N_10335,N_9143);
nor U13383 (N_13383,N_9520,N_10144);
and U13384 (N_13384,N_10272,N_11305);
or U13385 (N_13385,N_10623,N_11204);
nor U13386 (N_13386,N_10906,N_10536);
or U13387 (N_13387,N_11597,N_10433);
or U13388 (N_13388,N_10076,N_9852);
and U13389 (N_13389,N_11986,N_11732);
or U13390 (N_13390,N_11644,N_10653);
nor U13391 (N_13391,N_9640,N_9269);
or U13392 (N_13392,N_10825,N_9652);
xnor U13393 (N_13393,N_9624,N_10021);
or U13394 (N_13394,N_10321,N_9460);
or U13395 (N_13395,N_11641,N_10954);
or U13396 (N_13396,N_9158,N_10788);
and U13397 (N_13397,N_9125,N_9541);
xor U13398 (N_13398,N_10525,N_10529);
nand U13399 (N_13399,N_9866,N_11855);
and U13400 (N_13400,N_9093,N_11671);
and U13401 (N_13401,N_9097,N_11094);
and U13402 (N_13402,N_9466,N_9768);
or U13403 (N_13403,N_9130,N_11731);
xor U13404 (N_13404,N_11787,N_10133);
or U13405 (N_13405,N_10088,N_11064);
or U13406 (N_13406,N_11718,N_9429);
nor U13407 (N_13407,N_11478,N_9075);
xor U13408 (N_13408,N_9706,N_9513);
xor U13409 (N_13409,N_9392,N_11536);
or U13410 (N_13410,N_9828,N_9612);
nand U13411 (N_13411,N_9218,N_10659);
nand U13412 (N_13412,N_11546,N_9647);
and U13413 (N_13413,N_11722,N_9003);
nor U13414 (N_13414,N_9579,N_9709);
nor U13415 (N_13415,N_10599,N_10251);
or U13416 (N_13416,N_11781,N_11941);
nand U13417 (N_13417,N_9424,N_10910);
nand U13418 (N_13418,N_9713,N_11681);
nor U13419 (N_13419,N_11165,N_10766);
nor U13420 (N_13420,N_9563,N_11686);
and U13421 (N_13421,N_11531,N_10700);
nand U13422 (N_13422,N_11766,N_9999);
nand U13423 (N_13423,N_10586,N_10509);
nand U13424 (N_13424,N_10956,N_10655);
and U13425 (N_13425,N_11417,N_11472);
or U13426 (N_13426,N_9077,N_9879);
and U13427 (N_13427,N_10351,N_11365);
xnor U13428 (N_13428,N_10414,N_9273);
nor U13429 (N_13429,N_9148,N_10936);
xor U13430 (N_13430,N_10736,N_10261);
xor U13431 (N_13431,N_9033,N_10385);
xor U13432 (N_13432,N_10238,N_10647);
xor U13433 (N_13433,N_9073,N_9210);
nand U13434 (N_13434,N_9702,N_9071);
xor U13435 (N_13435,N_10888,N_10363);
xnor U13436 (N_13436,N_10994,N_11807);
nand U13437 (N_13437,N_10034,N_11309);
nand U13438 (N_13438,N_9910,N_10803);
nor U13439 (N_13439,N_9522,N_10719);
nor U13440 (N_13440,N_10513,N_10753);
xor U13441 (N_13441,N_10593,N_11512);
nand U13442 (N_13442,N_10230,N_9803);
nand U13443 (N_13443,N_11347,N_11500);
xnor U13444 (N_13444,N_9687,N_9554);
xnor U13445 (N_13445,N_10079,N_11959);
or U13446 (N_13446,N_10573,N_9604);
xor U13447 (N_13447,N_11306,N_10799);
xor U13448 (N_13448,N_9380,N_11922);
nand U13449 (N_13449,N_10313,N_10169);
or U13450 (N_13450,N_10164,N_9297);
and U13451 (N_13451,N_11810,N_10046);
xnor U13452 (N_13452,N_11555,N_9648);
xnor U13453 (N_13453,N_9459,N_11425);
nand U13454 (N_13454,N_10489,N_11264);
xnor U13455 (N_13455,N_11806,N_11134);
or U13456 (N_13456,N_11206,N_9751);
nor U13457 (N_13457,N_9712,N_11282);
nand U13458 (N_13458,N_11963,N_9251);
nand U13459 (N_13459,N_9361,N_9428);
xor U13460 (N_13460,N_10683,N_9110);
nand U13461 (N_13461,N_11060,N_10698);
nor U13462 (N_13462,N_10023,N_10415);
and U13463 (N_13463,N_10066,N_11585);
nand U13464 (N_13464,N_9014,N_11544);
nand U13465 (N_13465,N_11290,N_11677);
xnor U13466 (N_13466,N_9220,N_9923);
or U13467 (N_13467,N_10887,N_10456);
nor U13468 (N_13468,N_11356,N_9974);
or U13469 (N_13469,N_9789,N_9620);
and U13470 (N_13470,N_9808,N_10052);
and U13471 (N_13471,N_9574,N_10084);
or U13472 (N_13472,N_9696,N_9315);
and U13473 (N_13473,N_9669,N_9360);
nand U13474 (N_13474,N_9772,N_11095);
and U13475 (N_13475,N_10194,N_10206);
or U13476 (N_13476,N_9865,N_9002);
xor U13477 (N_13477,N_10648,N_10567);
or U13478 (N_13478,N_11601,N_10907);
and U13479 (N_13479,N_11792,N_11509);
and U13480 (N_13480,N_9738,N_9115);
xnor U13481 (N_13481,N_9965,N_9306);
or U13482 (N_13482,N_10296,N_9708);
nand U13483 (N_13483,N_10178,N_9374);
or U13484 (N_13484,N_11598,N_11654);
and U13485 (N_13485,N_9327,N_10378);
nand U13486 (N_13486,N_11083,N_9391);
nor U13487 (N_13487,N_9010,N_9335);
nor U13488 (N_13488,N_11708,N_11895);
nor U13489 (N_13489,N_11640,N_10237);
nand U13490 (N_13490,N_10040,N_10341);
nand U13491 (N_13491,N_10537,N_11073);
nor U13492 (N_13492,N_11329,N_9587);
and U13493 (N_13493,N_11593,N_11697);
or U13494 (N_13494,N_10636,N_9802);
and U13495 (N_13495,N_11609,N_10198);
nand U13496 (N_13496,N_9880,N_10800);
or U13497 (N_13497,N_10941,N_11161);
or U13498 (N_13498,N_10589,N_9081);
nand U13499 (N_13499,N_9876,N_9393);
nand U13500 (N_13500,N_9460,N_10243);
or U13501 (N_13501,N_9300,N_10902);
and U13502 (N_13502,N_10722,N_9831);
nand U13503 (N_13503,N_11575,N_10070);
and U13504 (N_13504,N_10616,N_10257);
and U13505 (N_13505,N_10504,N_9621);
nand U13506 (N_13506,N_11267,N_11348);
or U13507 (N_13507,N_10308,N_10400);
and U13508 (N_13508,N_10518,N_11394);
nand U13509 (N_13509,N_9082,N_10201);
and U13510 (N_13510,N_10915,N_10639);
xnor U13511 (N_13511,N_10240,N_9109);
xnor U13512 (N_13512,N_11144,N_11128);
xnor U13513 (N_13513,N_9750,N_11188);
nor U13514 (N_13514,N_10682,N_9584);
nor U13515 (N_13515,N_9274,N_11849);
or U13516 (N_13516,N_10046,N_9158);
and U13517 (N_13517,N_9788,N_9200);
and U13518 (N_13518,N_9965,N_10736);
nand U13519 (N_13519,N_11135,N_9557);
and U13520 (N_13520,N_11048,N_10794);
or U13521 (N_13521,N_10754,N_9412);
or U13522 (N_13522,N_11912,N_10817);
or U13523 (N_13523,N_10935,N_9280);
or U13524 (N_13524,N_9770,N_11990);
or U13525 (N_13525,N_9416,N_11486);
xnor U13526 (N_13526,N_11856,N_9643);
xor U13527 (N_13527,N_11195,N_10060);
xor U13528 (N_13528,N_9725,N_9757);
nand U13529 (N_13529,N_9120,N_11522);
and U13530 (N_13530,N_10285,N_11663);
and U13531 (N_13531,N_10624,N_10133);
xnor U13532 (N_13532,N_9176,N_9953);
xor U13533 (N_13533,N_10590,N_10910);
or U13534 (N_13534,N_9112,N_9962);
or U13535 (N_13535,N_9161,N_9185);
nand U13536 (N_13536,N_10265,N_11874);
xor U13537 (N_13537,N_11936,N_9369);
xor U13538 (N_13538,N_11279,N_10560);
and U13539 (N_13539,N_10758,N_9280);
or U13540 (N_13540,N_9438,N_10444);
xnor U13541 (N_13541,N_10282,N_11907);
nand U13542 (N_13542,N_10232,N_11005);
nor U13543 (N_13543,N_9819,N_11806);
nor U13544 (N_13544,N_11927,N_11946);
nand U13545 (N_13545,N_10732,N_9015);
xnor U13546 (N_13546,N_10545,N_9949);
nand U13547 (N_13547,N_10358,N_10974);
nor U13548 (N_13548,N_11597,N_11925);
xnor U13549 (N_13549,N_10234,N_11539);
and U13550 (N_13550,N_11214,N_10977);
nand U13551 (N_13551,N_9462,N_11745);
nor U13552 (N_13552,N_11397,N_10150);
nand U13553 (N_13553,N_9659,N_9079);
or U13554 (N_13554,N_10409,N_10217);
nand U13555 (N_13555,N_11785,N_9787);
nand U13556 (N_13556,N_9948,N_9535);
nor U13557 (N_13557,N_10436,N_10739);
nand U13558 (N_13558,N_11859,N_10224);
or U13559 (N_13559,N_10865,N_11103);
nor U13560 (N_13560,N_10009,N_10274);
and U13561 (N_13561,N_11527,N_9451);
xor U13562 (N_13562,N_10648,N_11323);
or U13563 (N_13563,N_9441,N_11395);
xnor U13564 (N_13564,N_9654,N_11746);
xnor U13565 (N_13565,N_11340,N_10846);
nor U13566 (N_13566,N_9306,N_10843);
nand U13567 (N_13567,N_11957,N_11655);
nor U13568 (N_13568,N_11140,N_10521);
or U13569 (N_13569,N_9438,N_11152);
nand U13570 (N_13570,N_10689,N_10034);
and U13571 (N_13571,N_11850,N_11525);
and U13572 (N_13572,N_11356,N_11388);
and U13573 (N_13573,N_11695,N_10487);
xor U13574 (N_13574,N_11756,N_11096);
nor U13575 (N_13575,N_11195,N_11651);
and U13576 (N_13576,N_11903,N_9374);
or U13577 (N_13577,N_10637,N_11990);
or U13578 (N_13578,N_11301,N_11249);
or U13579 (N_13579,N_9281,N_9340);
or U13580 (N_13580,N_10126,N_9185);
xor U13581 (N_13581,N_10441,N_9890);
xor U13582 (N_13582,N_10173,N_11990);
and U13583 (N_13583,N_11071,N_9962);
nor U13584 (N_13584,N_9663,N_9712);
xnor U13585 (N_13585,N_9559,N_10622);
nor U13586 (N_13586,N_11960,N_10074);
and U13587 (N_13587,N_9363,N_9996);
xor U13588 (N_13588,N_11796,N_10168);
nor U13589 (N_13589,N_11642,N_9470);
or U13590 (N_13590,N_9602,N_9953);
nand U13591 (N_13591,N_9727,N_11873);
or U13592 (N_13592,N_11633,N_10421);
and U13593 (N_13593,N_11510,N_9101);
nor U13594 (N_13594,N_11275,N_11968);
xnor U13595 (N_13595,N_11981,N_9964);
nand U13596 (N_13596,N_11055,N_10405);
or U13597 (N_13597,N_11388,N_11008);
xnor U13598 (N_13598,N_11947,N_11804);
nor U13599 (N_13599,N_9219,N_10267);
nor U13600 (N_13600,N_11379,N_9826);
and U13601 (N_13601,N_11395,N_11957);
or U13602 (N_13602,N_10271,N_11256);
nor U13603 (N_13603,N_11598,N_11452);
nor U13604 (N_13604,N_9110,N_10186);
nand U13605 (N_13605,N_11751,N_11636);
nor U13606 (N_13606,N_9493,N_10698);
nand U13607 (N_13607,N_10636,N_11972);
nand U13608 (N_13608,N_10776,N_10966);
and U13609 (N_13609,N_9805,N_10926);
and U13610 (N_13610,N_11555,N_11252);
or U13611 (N_13611,N_9440,N_10453);
and U13612 (N_13612,N_9333,N_9367);
or U13613 (N_13613,N_10673,N_10527);
or U13614 (N_13614,N_11968,N_11727);
nand U13615 (N_13615,N_10955,N_10487);
xnor U13616 (N_13616,N_11913,N_9748);
xnor U13617 (N_13617,N_11308,N_9903);
nand U13618 (N_13618,N_9771,N_9909);
nand U13619 (N_13619,N_11517,N_10459);
and U13620 (N_13620,N_11259,N_11889);
xnor U13621 (N_13621,N_10903,N_10426);
and U13622 (N_13622,N_10081,N_10026);
and U13623 (N_13623,N_10169,N_11736);
xor U13624 (N_13624,N_9574,N_10486);
nor U13625 (N_13625,N_9866,N_9348);
nor U13626 (N_13626,N_10021,N_9638);
nand U13627 (N_13627,N_11638,N_9738);
xnor U13628 (N_13628,N_10263,N_11850);
nor U13629 (N_13629,N_10366,N_9029);
xnor U13630 (N_13630,N_11848,N_9441);
nor U13631 (N_13631,N_10100,N_11784);
xor U13632 (N_13632,N_9000,N_9786);
nor U13633 (N_13633,N_10777,N_10118);
nand U13634 (N_13634,N_10039,N_9075);
or U13635 (N_13635,N_10738,N_11769);
or U13636 (N_13636,N_9884,N_10199);
xor U13637 (N_13637,N_11352,N_11218);
or U13638 (N_13638,N_11260,N_11203);
and U13639 (N_13639,N_10980,N_10058);
xor U13640 (N_13640,N_9195,N_11643);
nor U13641 (N_13641,N_11471,N_11968);
or U13642 (N_13642,N_11804,N_11015);
nand U13643 (N_13643,N_11911,N_10094);
xnor U13644 (N_13644,N_9629,N_9131);
nand U13645 (N_13645,N_11486,N_11166);
and U13646 (N_13646,N_10430,N_10275);
nand U13647 (N_13647,N_10467,N_11788);
nand U13648 (N_13648,N_10647,N_11512);
nand U13649 (N_13649,N_11818,N_10878);
or U13650 (N_13650,N_11667,N_10921);
and U13651 (N_13651,N_11333,N_11093);
nor U13652 (N_13652,N_11361,N_11370);
nor U13653 (N_13653,N_9080,N_10285);
nand U13654 (N_13654,N_10066,N_9424);
nor U13655 (N_13655,N_10763,N_9955);
nand U13656 (N_13656,N_11368,N_11606);
and U13657 (N_13657,N_10018,N_10608);
nor U13658 (N_13658,N_10634,N_9120);
and U13659 (N_13659,N_10781,N_11845);
and U13660 (N_13660,N_10477,N_10272);
nand U13661 (N_13661,N_11535,N_10464);
or U13662 (N_13662,N_11294,N_10402);
nand U13663 (N_13663,N_10380,N_10660);
nor U13664 (N_13664,N_9650,N_9731);
and U13665 (N_13665,N_9292,N_11439);
nor U13666 (N_13666,N_11662,N_11274);
nand U13667 (N_13667,N_9644,N_9482);
xnor U13668 (N_13668,N_11530,N_9516);
xnor U13669 (N_13669,N_11803,N_11904);
or U13670 (N_13670,N_10212,N_9562);
and U13671 (N_13671,N_9065,N_10028);
and U13672 (N_13672,N_11986,N_10225);
xor U13673 (N_13673,N_11938,N_11753);
and U13674 (N_13674,N_11146,N_10684);
nor U13675 (N_13675,N_11158,N_10290);
xor U13676 (N_13676,N_10534,N_10137);
nand U13677 (N_13677,N_9370,N_11252);
and U13678 (N_13678,N_9778,N_11751);
or U13679 (N_13679,N_11602,N_11587);
and U13680 (N_13680,N_11199,N_11854);
nand U13681 (N_13681,N_11590,N_11535);
nand U13682 (N_13682,N_10174,N_9744);
or U13683 (N_13683,N_10399,N_9804);
and U13684 (N_13684,N_9779,N_11215);
xor U13685 (N_13685,N_11839,N_10244);
and U13686 (N_13686,N_10728,N_9910);
or U13687 (N_13687,N_9344,N_11151);
or U13688 (N_13688,N_10905,N_11452);
and U13689 (N_13689,N_9198,N_11374);
xnor U13690 (N_13690,N_10758,N_9148);
nor U13691 (N_13691,N_11501,N_10930);
nand U13692 (N_13692,N_11026,N_9437);
or U13693 (N_13693,N_9577,N_10223);
and U13694 (N_13694,N_9274,N_9677);
xor U13695 (N_13695,N_9746,N_9888);
xor U13696 (N_13696,N_10254,N_10264);
nand U13697 (N_13697,N_10031,N_10017);
nor U13698 (N_13698,N_9398,N_11486);
or U13699 (N_13699,N_10005,N_9705);
nor U13700 (N_13700,N_10414,N_11892);
or U13701 (N_13701,N_10514,N_10883);
nor U13702 (N_13702,N_9600,N_9185);
or U13703 (N_13703,N_11810,N_9323);
nand U13704 (N_13704,N_10582,N_9379);
nand U13705 (N_13705,N_9114,N_9763);
and U13706 (N_13706,N_11207,N_9631);
nor U13707 (N_13707,N_9358,N_9241);
or U13708 (N_13708,N_11252,N_9238);
nand U13709 (N_13709,N_11287,N_10439);
or U13710 (N_13710,N_9102,N_10193);
nor U13711 (N_13711,N_9000,N_10523);
nor U13712 (N_13712,N_9976,N_10090);
xnor U13713 (N_13713,N_11646,N_11117);
nand U13714 (N_13714,N_10647,N_10440);
or U13715 (N_13715,N_9447,N_10520);
nand U13716 (N_13716,N_9319,N_9337);
or U13717 (N_13717,N_9211,N_9472);
and U13718 (N_13718,N_11777,N_11468);
xor U13719 (N_13719,N_9154,N_10162);
xor U13720 (N_13720,N_9655,N_9385);
nand U13721 (N_13721,N_11377,N_11080);
or U13722 (N_13722,N_9538,N_10932);
nor U13723 (N_13723,N_10576,N_10734);
or U13724 (N_13724,N_11976,N_11032);
nor U13725 (N_13725,N_10005,N_11579);
nor U13726 (N_13726,N_9049,N_11643);
nor U13727 (N_13727,N_9654,N_9540);
nor U13728 (N_13728,N_9339,N_9566);
nand U13729 (N_13729,N_11032,N_9002);
or U13730 (N_13730,N_10777,N_10080);
nor U13731 (N_13731,N_9326,N_9921);
nand U13732 (N_13732,N_10615,N_10817);
nor U13733 (N_13733,N_10099,N_11962);
nor U13734 (N_13734,N_9436,N_10436);
and U13735 (N_13735,N_9461,N_9032);
xnor U13736 (N_13736,N_11002,N_10430);
and U13737 (N_13737,N_9879,N_11939);
nand U13738 (N_13738,N_11681,N_9225);
or U13739 (N_13739,N_10045,N_9495);
and U13740 (N_13740,N_9221,N_10890);
and U13741 (N_13741,N_9275,N_9072);
nand U13742 (N_13742,N_9328,N_11811);
or U13743 (N_13743,N_9377,N_10475);
and U13744 (N_13744,N_9891,N_11385);
and U13745 (N_13745,N_9955,N_10324);
and U13746 (N_13746,N_11424,N_10070);
or U13747 (N_13747,N_11543,N_9562);
or U13748 (N_13748,N_10167,N_10380);
nor U13749 (N_13749,N_9031,N_9026);
or U13750 (N_13750,N_11476,N_11516);
nand U13751 (N_13751,N_10085,N_11166);
nor U13752 (N_13752,N_11554,N_11298);
or U13753 (N_13753,N_10636,N_11546);
xnor U13754 (N_13754,N_9009,N_11935);
nor U13755 (N_13755,N_9260,N_11670);
or U13756 (N_13756,N_9016,N_9444);
nand U13757 (N_13757,N_9018,N_9386);
or U13758 (N_13758,N_9800,N_9876);
nand U13759 (N_13759,N_11065,N_9267);
xnor U13760 (N_13760,N_10275,N_10780);
xnor U13761 (N_13761,N_9279,N_10860);
or U13762 (N_13762,N_11231,N_9920);
xnor U13763 (N_13763,N_10695,N_9396);
or U13764 (N_13764,N_10325,N_10254);
and U13765 (N_13765,N_11983,N_9995);
or U13766 (N_13766,N_10390,N_10992);
or U13767 (N_13767,N_11302,N_10582);
nor U13768 (N_13768,N_9497,N_9675);
and U13769 (N_13769,N_11558,N_11371);
nand U13770 (N_13770,N_9464,N_9247);
xnor U13771 (N_13771,N_9437,N_10600);
or U13772 (N_13772,N_11639,N_10385);
or U13773 (N_13773,N_10108,N_10403);
or U13774 (N_13774,N_9127,N_9930);
xnor U13775 (N_13775,N_10979,N_10300);
nand U13776 (N_13776,N_11233,N_9336);
and U13777 (N_13777,N_10040,N_11859);
nor U13778 (N_13778,N_11932,N_11260);
and U13779 (N_13779,N_9159,N_11336);
or U13780 (N_13780,N_10709,N_10217);
and U13781 (N_13781,N_10801,N_10854);
and U13782 (N_13782,N_11433,N_9137);
or U13783 (N_13783,N_9994,N_11206);
nor U13784 (N_13784,N_10762,N_10800);
or U13785 (N_13785,N_11864,N_10687);
or U13786 (N_13786,N_9642,N_11352);
nand U13787 (N_13787,N_10748,N_10029);
and U13788 (N_13788,N_10347,N_9588);
nor U13789 (N_13789,N_11615,N_10215);
nor U13790 (N_13790,N_11010,N_10276);
xnor U13791 (N_13791,N_11540,N_10584);
nor U13792 (N_13792,N_11271,N_9776);
nor U13793 (N_13793,N_10375,N_9926);
or U13794 (N_13794,N_11885,N_10860);
nor U13795 (N_13795,N_10933,N_11137);
and U13796 (N_13796,N_11830,N_9545);
xor U13797 (N_13797,N_11228,N_11314);
nor U13798 (N_13798,N_10720,N_11258);
xor U13799 (N_13799,N_9813,N_10761);
and U13800 (N_13800,N_9854,N_11025);
and U13801 (N_13801,N_9563,N_10164);
xor U13802 (N_13802,N_9708,N_9417);
nor U13803 (N_13803,N_10297,N_9321);
and U13804 (N_13804,N_9609,N_10702);
nand U13805 (N_13805,N_9676,N_11597);
xor U13806 (N_13806,N_9867,N_11911);
nand U13807 (N_13807,N_9972,N_11176);
and U13808 (N_13808,N_10422,N_11845);
or U13809 (N_13809,N_9493,N_10996);
nor U13810 (N_13810,N_10402,N_10285);
and U13811 (N_13811,N_11161,N_11690);
and U13812 (N_13812,N_10146,N_10905);
and U13813 (N_13813,N_9303,N_11303);
or U13814 (N_13814,N_9283,N_11147);
or U13815 (N_13815,N_10843,N_11197);
and U13816 (N_13816,N_11917,N_10980);
xnor U13817 (N_13817,N_10495,N_10648);
nor U13818 (N_13818,N_10303,N_10115);
and U13819 (N_13819,N_10266,N_11793);
nand U13820 (N_13820,N_9092,N_9524);
and U13821 (N_13821,N_9319,N_11880);
and U13822 (N_13822,N_11651,N_11627);
nor U13823 (N_13823,N_9370,N_10418);
or U13824 (N_13824,N_10877,N_11065);
nor U13825 (N_13825,N_10495,N_9236);
and U13826 (N_13826,N_9403,N_9200);
nor U13827 (N_13827,N_11756,N_10517);
and U13828 (N_13828,N_10324,N_9356);
xor U13829 (N_13829,N_10374,N_11653);
and U13830 (N_13830,N_9376,N_11526);
nand U13831 (N_13831,N_9503,N_10266);
and U13832 (N_13832,N_10640,N_9254);
nor U13833 (N_13833,N_11816,N_11703);
nand U13834 (N_13834,N_10682,N_10451);
nor U13835 (N_13835,N_9170,N_9460);
or U13836 (N_13836,N_10612,N_10471);
or U13837 (N_13837,N_11983,N_10378);
nand U13838 (N_13838,N_10114,N_11846);
nand U13839 (N_13839,N_10428,N_10634);
or U13840 (N_13840,N_11832,N_11057);
or U13841 (N_13841,N_10157,N_9979);
nor U13842 (N_13842,N_11266,N_11336);
nor U13843 (N_13843,N_9784,N_10868);
or U13844 (N_13844,N_11751,N_10435);
or U13845 (N_13845,N_11342,N_11760);
xnor U13846 (N_13846,N_9070,N_10185);
nand U13847 (N_13847,N_9817,N_9951);
or U13848 (N_13848,N_11427,N_11522);
nor U13849 (N_13849,N_11690,N_9877);
nand U13850 (N_13850,N_11859,N_9303);
or U13851 (N_13851,N_9005,N_11715);
nor U13852 (N_13852,N_9581,N_11412);
nand U13853 (N_13853,N_9717,N_9970);
or U13854 (N_13854,N_9982,N_9215);
nor U13855 (N_13855,N_10337,N_11092);
xnor U13856 (N_13856,N_10364,N_10047);
nand U13857 (N_13857,N_11244,N_11927);
nor U13858 (N_13858,N_11063,N_11684);
and U13859 (N_13859,N_10133,N_9799);
nand U13860 (N_13860,N_11716,N_11295);
nand U13861 (N_13861,N_10893,N_9630);
nor U13862 (N_13862,N_11997,N_11618);
nand U13863 (N_13863,N_10208,N_9877);
xor U13864 (N_13864,N_11233,N_11192);
or U13865 (N_13865,N_10144,N_11271);
or U13866 (N_13866,N_9735,N_9447);
or U13867 (N_13867,N_9925,N_9202);
nand U13868 (N_13868,N_9215,N_10500);
nor U13869 (N_13869,N_11678,N_11323);
and U13870 (N_13870,N_11263,N_9666);
nand U13871 (N_13871,N_11117,N_9562);
and U13872 (N_13872,N_9954,N_10975);
xnor U13873 (N_13873,N_9319,N_11525);
nor U13874 (N_13874,N_11712,N_9521);
or U13875 (N_13875,N_10807,N_9035);
nor U13876 (N_13876,N_10871,N_9907);
or U13877 (N_13877,N_9602,N_10621);
or U13878 (N_13878,N_11574,N_11375);
nor U13879 (N_13879,N_11149,N_9761);
or U13880 (N_13880,N_10990,N_10207);
nand U13881 (N_13881,N_11954,N_10380);
and U13882 (N_13882,N_10064,N_9134);
nor U13883 (N_13883,N_11548,N_10163);
nand U13884 (N_13884,N_10714,N_9445);
or U13885 (N_13885,N_10708,N_10743);
xnor U13886 (N_13886,N_10465,N_10255);
nor U13887 (N_13887,N_11816,N_11768);
nor U13888 (N_13888,N_10170,N_11408);
nand U13889 (N_13889,N_9199,N_9878);
and U13890 (N_13890,N_10052,N_9179);
xnor U13891 (N_13891,N_11952,N_9395);
nor U13892 (N_13892,N_11795,N_9879);
nor U13893 (N_13893,N_10674,N_9918);
and U13894 (N_13894,N_10203,N_9888);
nand U13895 (N_13895,N_10145,N_10535);
or U13896 (N_13896,N_9961,N_9272);
xnor U13897 (N_13897,N_10783,N_11973);
nand U13898 (N_13898,N_11736,N_10201);
nor U13899 (N_13899,N_9758,N_11554);
nand U13900 (N_13900,N_9922,N_9806);
xor U13901 (N_13901,N_11692,N_10860);
nand U13902 (N_13902,N_9442,N_10013);
or U13903 (N_13903,N_9295,N_9322);
xnor U13904 (N_13904,N_9140,N_11483);
nor U13905 (N_13905,N_9240,N_9605);
nor U13906 (N_13906,N_11127,N_10564);
nor U13907 (N_13907,N_9964,N_10876);
xor U13908 (N_13908,N_11191,N_9700);
or U13909 (N_13909,N_9254,N_10129);
xor U13910 (N_13910,N_11272,N_10554);
nor U13911 (N_13911,N_11008,N_10616);
or U13912 (N_13912,N_10619,N_10810);
nor U13913 (N_13913,N_9413,N_9810);
or U13914 (N_13914,N_10950,N_10245);
nor U13915 (N_13915,N_9539,N_11662);
nor U13916 (N_13916,N_11500,N_9270);
nand U13917 (N_13917,N_11914,N_11932);
nor U13918 (N_13918,N_10919,N_9623);
or U13919 (N_13919,N_9753,N_11401);
and U13920 (N_13920,N_11346,N_10525);
xnor U13921 (N_13921,N_10287,N_11738);
nor U13922 (N_13922,N_9789,N_10662);
xor U13923 (N_13923,N_10466,N_11730);
nor U13924 (N_13924,N_11992,N_11192);
nand U13925 (N_13925,N_10325,N_10884);
or U13926 (N_13926,N_9828,N_9806);
nand U13927 (N_13927,N_11377,N_9531);
and U13928 (N_13928,N_10469,N_11125);
or U13929 (N_13929,N_9579,N_10013);
and U13930 (N_13930,N_10337,N_9931);
or U13931 (N_13931,N_10357,N_9452);
nand U13932 (N_13932,N_11864,N_10780);
or U13933 (N_13933,N_9391,N_9999);
nor U13934 (N_13934,N_11578,N_11916);
nor U13935 (N_13935,N_10286,N_9722);
xnor U13936 (N_13936,N_10899,N_10982);
xor U13937 (N_13937,N_10427,N_9689);
nor U13938 (N_13938,N_9274,N_11569);
or U13939 (N_13939,N_10388,N_10703);
or U13940 (N_13940,N_11040,N_9426);
and U13941 (N_13941,N_9730,N_10400);
nor U13942 (N_13942,N_9533,N_11856);
xnor U13943 (N_13943,N_11206,N_10745);
nand U13944 (N_13944,N_11229,N_9037);
nand U13945 (N_13945,N_9769,N_11521);
xnor U13946 (N_13946,N_10486,N_9537);
and U13947 (N_13947,N_11566,N_10762);
or U13948 (N_13948,N_10297,N_10100);
nor U13949 (N_13949,N_9146,N_10219);
or U13950 (N_13950,N_11418,N_9077);
nand U13951 (N_13951,N_10170,N_9941);
or U13952 (N_13952,N_10619,N_9937);
and U13953 (N_13953,N_9143,N_9142);
or U13954 (N_13954,N_11569,N_11987);
xor U13955 (N_13955,N_11167,N_9352);
or U13956 (N_13956,N_11979,N_9094);
nor U13957 (N_13957,N_9190,N_11739);
nand U13958 (N_13958,N_10616,N_10121);
nand U13959 (N_13959,N_11489,N_9930);
nand U13960 (N_13960,N_10660,N_9251);
or U13961 (N_13961,N_10576,N_9387);
nand U13962 (N_13962,N_9087,N_9592);
nand U13963 (N_13963,N_11692,N_9034);
or U13964 (N_13964,N_11765,N_9569);
nor U13965 (N_13965,N_9754,N_10409);
or U13966 (N_13966,N_10259,N_9279);
nand U13967 (N_13967,N_9877,N_9885);
and U13968 (N_13968,N_10586,N_11743);
nor U13969 (N_13969,N_11884,N_10958);
xor U13970 (N_13970,N_11903,N_11753);
xor U13971 (N_13971,N_9014,N_9082);
and U13972 (N_13972,N_9822,N_10544);
and U13973 (N_13973,N_10114,N_11241);
nor U13974 (N_13974,N_11372,N_10407);
or U13975 (N_13975,N_9036,N_10081);
nand U13976 (N_13976,N_11101,N_11262);
xnor U13977 (N_13977,N_9104,N_10634);
nand U13978 (N_13978,N_11156,N_10699);
and U13979 (N_13979,N_10732,N_9383);
nand U13980 (N_13980,N_10286,N_9283);
nand U13981 (N_13981,N_11353,N_9708);
nand U13982 (N_13982,N_9067,N_11819);
and U13983 (N_13983,N_11475,N_11368);
or U13984 (N_13984,N_9498,N_11925);
and U13985 (N_13985,N_10637,N_10135);
xnor U13986 (N_13986,N_10384,N_11110);
xor U13987 (N_13987,N_9360,N_11415);
or U13988 (N_13988,N_10125,N_9299);
nand U13989 (N_13989,N_11349,N_9791);
and U13990 (N_13990,N_11110,N_10759);
nand U13991 (N_13991,N_11814,N_9576);
nand U13992 (N_13992,N_10412,N_10443);
and U13993 (N_13993,N_11858,N_11674);
or U13994 (N_13994,N_11187,N_10691);
xnor U13995 (N_13995,N_11271,N_10283);
and U13996 (N_13996,N_9005,N_10250);
or U13997 (N_13997,N_10367,N_9363);
xor U13998 (N_13998,N_9159,N_10505);
xor U13999 (N_13999,N_11061,N_9588);
and U14000 (N_14000,N_9936,N_9770);
or U14001 (N_14001,N_11279,N_9716);
nand U14002 (N_14002,N_9936,N_10955);
nand U14003 (N_14003,N_9471,N_10779);
nor U14004 (N_14004,N_11107,N_9369);
xor U14005 (N_14005,N_10563,N_9815);
nor U14006 (N_14006,N_11308,N_9827);
nand U14007 (N_14007,N_9269,N_11002);
and U14008 (N_14008,N_10572,N_11742);
or U14009 (N_14009,N_10175,N_11403);
or U14010 (N_14010,N_11728,N_9466);
or U14011 (N_14011,N_9466,N_10623);
nor U14012 (N_14012,N_9155,N_11002);
nand U14013 (N_14013,N_9639,N_10215);
and U14014 (N_14014,N_11347,N_11068);
and U14015 (N_14015,N_9894,N_11908);
or U14016 (N_14016,N_10700,N_11525);
xnor U14017 (N_14017,N_11948,N_10128);
and U14018 (N_14018,N_11993,N_9701);
and U14019 (N_14019,N_9717,N_9481);
or U14020 (N_14020,N_9135,N_11186);
nor U14021 (N_14021,N_9718,N_9068);
and U14022 (N_14022,N_11774,N_9074);
and U14023 (N_14023,N_10173,N_9769);
nand U14024 (N_14024,N_10388,N_10368);
or U14025 (N_14025,N_9915,N_9682);
xor U14026 (N_14026,N_9979,N_9190);
nor U14027 (N_14027,N_11233,N_9545);
and U14028 (N_14028,N_11384,N_11644);
and U14029 (N_14029,N_11152,N_9351);
and U14030 (N_14030,N_9295,N_11868);
xor U14031 (N_14031,N_11570,N_10954);
xor U14032 (N_14032,N_10090,N_11740);
and U14033 (N_14033,N_9442,N_10852);
or U14034 (N_14034,N_10588,N_11835);
or U14035 (N_14035,N_10379,N_11150);
and U14036 (N_14036,N_10252,N_9760);
or U14037 (N_14037,N_9636,N_10430);
and U14038 (N_14038,N_9280,N_9151);
and U14039 (N_14039,N_9555,N_9361);
nor U14040 (N_14040,N_11059,N_9769);
or U14041 (N_14041,N_10993,N_11569);
xnor U14042 (N_14042,N_10062,N_10943);
nand U14043 (N_14043,N_10175,N_9776);
nor U14044 (N_14044,N_11979,N_9590);
nor U14045 (N_14045,N_10527,N_9395);
or U14046 (N_14046,N_11176,N_11166);
or U14047 (N_14047,N_9797,N_11105);
and U14048 (N_14048,N_10554,N_10324);
nand U14049 (N_14049,N_11767,N_11709);
and U14050 (N_14050,N_11455,N_10388);
nor U14051 (N_14051,N_10672,N_10443);
or U14052 (N_14052,N_11592,N_9540);
or U14053 (N_14053,N_11117,N_10758);
and U14054 (N_14054,N_9150,N_10772);
nand U14055 (N_14055,N_11468,N_9457);
nor U14056 (N_14056,N_9682,N_11094);
nand U14057 (N_14057,N_9780,N_11207);
and U14058 (N_14058,N_10946,N_10765);
or U14059 (N_14059,N_11509,N_11076);
nand U14060 (N_14060,N_11043,N_11289);
and U14061 (N_14061,N_10990,N_10319);
nor U14062 (N_14062,N_10393,N_10987);
nor U14063 (N_14063,N_10914,N_9169);
xor U14064 (N_14064,N_9204,N_11859);
xnor U14065 (N_14065,N_9420,N_9323);
xor U14066 (N_14066,N_10289,N_10307);
or U14067 (N_14067,N_9288,N_9244);
nor U14068 (N_14068,N_10498,N_9400);
and U14069 (N_14069,N_10848,N_9525);
nor U14070 (N_14070,N_11380,N_10656);
xnor U14071 (N_14071,N_11306,N_10955);
nor U14072 (N_14072,N_10273,N_10238);
nand U14073 (N_14073,N_11630,N_11554);
nor U14074 (N_14074,N_9342,N_10884);
nand U14075 (N_14075,N_11769,N_11480);
xnor U14076 (N_14076,N_11679,N_11571);
or U14077 (N_14077,N_11356,N_11948);
or U14078 (N_14078,N_9554,N_11421);
nand U14079 (N_14079,N_11980,N_10171);
nand U14080 (N_14080,N_11528,N_10073);
nand U14081 (N_14081,N_10286,N_11547);
xnor U14082 (N_14082,N_11431,N_9972);
and U14083 (N_14083,N_10191,N_10192);
or U14084 (N_14084,N_9838,N_10697);
xor U14085 (N_14085,N_10644,N_10027);
nand U14086 (N_14086,N_10960,N_10145);
or U14087 (N_14087,N_10789,N_9758);
and U14088 (N_14088,N_10756,N_10539);
nor U14089 (N_14089,N_10709,N_10230);
xnor U14090 (N_14090,N_11534,N_10040);
nand U14091 (N_14091,N_11505,N_11966);
and U14092 (N_14092,N_10772,N_11641);
nand U14093 (N_14093,N_11830,N_11551);
nand U14094 (N_14094,N_9251,N_11888);
or U14095 (N_14095,N_10796,N_10046);
nor U14096 (N_14096,N_11159,N_9582);
and U14097 (N_14097,N_9679,N_9759);
or U14098 (N_14098,N_10229,N_11194);
and U14099 (N_14099,N_11920,N_9076);
nand U14100 (N_14100,N_11116,N_10185);
xnor U14101 (N_14101,N_10048,N_9637);
and U14102 (N_14102,N_9589,N_9502);
or U14103 (N_14103,N_10664,N_10538);
or U14104 (N_14104,N_10943,N_9036);
or U14105 (N_14105,N_10315,N_9411);
nand U14106 (N_14106,N_9576,N_10667);
xor U14107 (N_14107,N_10945,N_11893);
nand U14108 (N_14108,N_10302,N_9445);
nand U14109 (N_14109,N_9870,N_11294);
nor U14110 (N_14110,N_9346,N_10073);
nand U14111 (N_14111,N_9341,N_10614);
or U14112 (N_14112,N_11500,N_10747);
or U14113 (N_14113,N_11564,N_9602);
xor U14114 (N_14114,N_10066,N_9443);
and U14115 (N_14115,N_9285,N_9757);
or U14116 (N_14116,N_9477,N_11551);
nor U14117 (N_14117,N_9800,N_9610);
nand U14118 (N_14118,N_9036,N_11105);
and U14119 (N_14119,N_10070,N_10074);
nand U14120 (N_14120,N_10330,N_11683);
xnor U14121 (N_14121,N_9167,N_11246);
xnor U14122 (N_14122,N_11543,N_10953);
or U14123 (N_14123,N_10814,N_11351);
and U14124 (N_14124,N_11019,N_10637);
and U14125 (N_14125,N_11835,N_9315);
and U14126 (N_14126,N_11116,N_10590);
nand U14127 (N_14127,N_11546,N_10946);
nand U14128 (N_14128,N_9855,N_10348);
nand U14129 (N_14129,N_10736,N_9394);
nand U14130 (N_14130,N_10930,N_10364);
xnor U14131 (N_14131,N_10564,N_10645);
xor U14132 (N_14132,N_11953,N_9828);
nand U14133 (N_14133,N_9266,N_11416);
nand U14134 (N_14134,N_11893,N_11375);
and U14135 (N_14135,N_10891,N_9056);
or U14136 (N_14136,N_10628,N_11697);
nor U14137 (N_14137,N_10957,N_9268);
or U14138 (N_14138,N_9023,N_9425);
xor U14139 (N_14139,N_9500,N_9348);
and U14140 (N_14140,N_9016,N_10123);
nor U14141 (N_14141,N_11143,N_9564);
nor U14142 (N_14142,N_10259,N_10419);
nand U14143 (N_14143,N_9008,N_9172);
nand U14144 (N_14144,N_9402,N_11919);
nand U14145 (N_14145,N_11846,N_10888);
and U14146 (N_14146,N_10547,N_10376);
nand U14147 (N_14147,N_11396,N_10822);
nor U14148 (N_14148,N_9354,N_10907);
xor U14149 (N_14149,N_10985,N_9742);
nand U14150 (N_14150,N_10066,N_11559);
and U14151 (N_14151,N_9121,N_9777);
or U14152 (N_14152,N_10343,N_10495);
xor U14153 (N_14153,N_9682,N_11887);
nand U14154 (N_14154,N_10889,N_11735);
and U14155 (N_14155,N_11177,N_10521);
nor U14156 (N_14156,N_9838,N_11714);
nand U14157 (N_14157,N_9591,N_10567);
and U14158 (N_14158,N_10745,N_10709);
nor U14159 (N_14159,N_11216,N_11804);
nor U14160 (N_14160,N_10975,N_10587);
nor U14161 (N_14161,N_10187,N_10976);
nor U14162 (N_14162,N_11720,N_10005);
and U14163 (N_14163,N_11410,N_10966);
xnor U14164 (N_14164,N_10809,N_10263);
nand U14165 (N_14165,N_11975,N_11334);
nor U14166 (N_14166,N_11955,N_11692);
nand U14167 (N_14167,N_10235,N_9833);
nor U14168 (N_14168,N_9314,N_10146);
and U14169 (N_14169,N_11759,N_11992);
xnor U14170 (N_14170,N_11215,N_9329);
and U14171 (N_14171,N_10856,N_9759);
or U14172 (N_14172,N_10689,N_10579);
and U14173 (N_14173,N_9308,N_11049);
nand U14174 (N_14174,N_10330,N_10297);
nor U14175 (N_14175,N_10150,N_11343);
and U14176 (N_14176,N_9304,N_10589);
xor U14177 (N_14177,N_9951,N_9942);
or U14178 (N_14178,N_10431,N_11753);
xor U14179 (N_14179,N_9117,N_9655);
and U14180 (N_14180,N_9711,N_11502);
and U14181 (N_14181,N_10770,N_9157);
nand U14182 (N_14182,N_11957,N_10490);
or U14183 (N_14183,N_10507,N_11070);
or U14184 (N_14184,N_11582,N_9274);
or U14185 (N_14185,N_11899,N_11154);
nand U14186 (N_14186,N_10042,N_11284);
nand U14187 (N_14187,N_11023,N_11901);
and U14188 (N_14188,N_9829,N_10455);
nor U14189 (N_14189,N_10552,N_9218);
nand U14190 (N_14190,N_9698,N_10572);
xor U14191 (N_14191,N_10294,N_11049);
nand U14192 (N_14192,N_11107,N_11443);
xnor U14193 (N_14193,N_9192,N_10448);
nand U14194 (N_14194,N_10831,N_11543);
nand U14195 (N_14195,N_10476,N_10675);
nor U14196 (N_14196,N_11597,N_11410);
nand U14197 (N_14197,N_9783,N_11021);
nor U14198 (N_14198,N_11747,N_11098);
or U14199 (N_14199,N_10235,N_9496);
nor U14200 (N_14200,N_9248,N_9469);
and U14201 (N_14201,N_11768,N_11108);
xnor U14202 (N_14202,N_9267,N_11133);
nand U14203 (N_14203,N_9595,N_11273);
nor U14204 (N_14204,N_10377,N_10944);
nor U14205 (N_14205,N_11883,N_11716);
and U14206 (N_14206,N_9417,N_11029);
and U14207 (N_14207,N_11108,N_11835);
or U14208 (N_14208,N_9680,N_9572);
or U14209 (N_14209,N_10044,N_9324);
xnor U14210 (N_14210,N_9328,N_9127);
nor U14211 (N_14211,N_10611,N_11546);
nand U14212 (N_14212,N_9997,N_11051);
nand U14213 (N_14213,N_11896,N_10961);
nor U14214 (N_14214,N_9251,N_11859);
nand U14215 (N_14215,N_11421,N_11547);
and U14216 (N_14216,N_10527,N_10187);
nand U14217 (N_14217,N_10960,N_11380);
xnor U14218 (N_14218,N_11000,N_11601);
and U14219 (N_14219,N_10116,N_11428);
or U14220 (N_14220,N_10365,N_9214);
and U14221 (N_14221,N_10721,N_11254);
nor U14222 (N_14222,N_11707,N_9342);
and U14223 (N_14223,N_10328,N_11445);
xor U14224 (N_14224,N_9331,N_10222);
nor U14225 (N_14225,N_9361,N_11922);
xnor U14226 (N_14226,N_9980,N_9468);
xor U14227 (N_14227,N_9395,N_11267);
nor U14228 (N_14228,N_11789,N_11648);
or U14229 (N_14229,N_10256,N_11751);
nand U14230 (N_14230,N_11190,N_10477);
and U14231 (N_14231,N_9870,N_10457);
xor U14232 (N_14232,N_11041,N_9753);
nand U14233 (N_14233,N_11679,N_9811);
or U14234 (N_14234,N_11182,N_10750);
nor U14235 (N_14235,N_11023,N_11577);
xor U14236 (N_14236,N_9976,N_10992);
xnor U14237 (N_14237,N_10638,N_10121);
or U14238 (N_14238,N_11215,N_10425);
xnor U14239 (N_14239,N_9859,N_11108);
and U14240 (N_14240,N_9964,N_10311);
and U14241 (N_14241,N_11654,N_11961);
or U14242 (N_14242,N_10219,N_10524);
or U14243 (N_14243,N_11844,N_9809);
or U14244 (N_14244,N_9627,N_11941);
nand U14245 (N_14245,N_11440,N_9834);
nand U14246 (N_14246,N_11712,N_11652);
and U14247 (N_14247,N_9589,N_10675);
xor U14248 (N_14248,N_10014,N_11662);
nand U14249 (N_14249,N_9481,N_11329);
nand U14250 (N_14250,N_10727,N_10221);
nand U14251 (N_14251,N_11176,N_11706);
nor U14252 (N_14252,N_10858,N_11728);
and U14253 (N_14253,N_9743,N_10068);
xor U14254 (N_14254,N_9241,N_10476);
and U14255 (N_14255,N_10017,N_10962);
or U14256 (N_14256,N_11451,N_11159);
nor U14257 (N_14257,N_10099,N_9188);
xor U14258 (N_14258,N_11395,N_11240);
nor U14259 (N_14259,N_9499,N_10981);
and U14260 (N_14260,N_9113,N_11786);
xnor U14261 (N_14261,N_11987,N_10845);
nand U14262 (N_14262,N_9545,N_11131);
and U14263 (N_14263,N_10628,N_10802);
nor U14264 (N_14264,N_9329,N_9658);
nor U14265 (N_14265,N_11685,N_9206);
or U14266 (N_14266,N_9936,N_11200);
nand U14267 (N_14267,N_10932,N_10602);
nor U14268 (N_14268,N_10846,N_9288);
and U14269 (N_14269,N_11543,N_11298);
nand U14270 (N_14270,N_10588,N_10481);
and U14271 (N_14271,N_11675,N_10780);
or U14272 (N_14272,N_9165,N_9787);
xnor U14273 (N_14273,N_9972,N_9936);
or U14274 (N_14274,N_11769,N_11373);
xnor U14275 (N_14275,N_9422,N_10773);
and U14276 (N_14276,N_10128,N_11983);
or U14277 (N_14277,N_9320,N_10195);
and U14278 (N_14278,N_10901,N_9135);
xnor U14279 (N_14279,N_10295,N_11858);
xnor U14280 (N_14280,N_9734,N_10243);
or U14281 (N_14281,N_11251,N_10247);
nor U14282 (N_14282,N_9064,N_9854);
and U14283 (N_14283,N_10723,N_11227);
nor U14284 (N_14284,N_9627,N_10729);
and U14285 (N_14285,N_11982,N_9430);
nor U14286 (N_14286,N_10059,N_9556);
and U14287 (N_14287,N_11916,N_10849);
and U14288 (N_14288,N_9997,N_9909);
nand U14289 (N_14289,N_9142,N_11315);
xor U14290 (N_14290,N_9674,N_11895);
xor U14291 (N_14291,N_10108,N_11397);
nand U14292 (N_14292,N_10100,N_9923);
and U14293 (N_14293,N_9137,N_9029);
or U14294 (N_14294,N_9581,N_9665);
nand U14295 (N_14295,N_10525,N_11332);
and U14296 (N_14296,N_10973,N_10839);
nand U14297 (N_14297,N_9582,N_10455);
and U14298 (N_14298,N_9529,N_9567);
or U14299 (N_14299,N_11363,N_10525);
nand U14300 (N_14300,N_9835,N_11173);
or U14301 (N_14301,N_11002,N_10866);
xor U14302 (N_14302,N_10984,N_11015);
nor U14303 (N_14303,N_10050,N_9789);
nor U14304 (N_14304,N_11475,N_9860);
or U14305 (N_14305,N_10128,N_10874);
nand U14306 (N_14306,N_10118,N_9181);
xor U14307 (N_14307,N_11521,N_10689);
xor U14308 (N_14308,N_11059,N_10306);
or U14309 (N_14309,N_9294,N_9766);
or U14310 (N_14310,N_10143,N_10231);
or U14311 (N_14311,N_10071,N_9932);
nand U14312 (N_14312,N_11113,N_9096);
and U14313 (N_14313,N_9505,N_10714);
nor U14314 (N_14314,N_10072,N_11062);
xnor U14315 (N_14315,N_11240,N_11572);
and U14316 (N_14316,N_10652,N_9827);
nand U14317 (N_14317,N_9180,N_10141);
nor U14318 (N_14318,N_11963,N_9133);
nand U14319 (N_14319,N_9620,N_9498);
xnor U14320 (N_14320,N_11758,N_11222);
or U14321 (N_14321,N_11658,N_11522);
nand U14322 (N_14322,N_11212,N_10859);
nor U14323 (N_14323,N_11025,N_9216);
nand U14324 (N_14324,N_10491,N_9591);
xnor U14325 (N_14325,N_10862,N_9621);
nor U14326 (N_14326,N_9623,N_10071);
xor U14327 (N_14327,N_10386,N_11902);
and U14328 (N_14328,N_9704,N_10121);
xnor U14329 (N_14329,N_11481,N_9327);
and U14330 (N_14330,N_9835,N_10746);
nor U14331 (N_14331,N_9687,N_11917);
nand U14332 (N_14332,N_10361,N_9061);
xor U14333 (N_14333,N_11581,N_11975);
or U14334 (N_14334,N_9017,N_9100);
nor U14335 (N_14335,N_9210,N_11148);
nor U14336 (N_14336,N_9995,N_10925);
nand U14337 (N_14337,N_10690,N_11987);
xor U14338 (N_14338,N_10188,N_11219);
and U14339 (N_14339,N_11660,N_10173);
xnor U14340 (N_14340,N_10469,N_9759);
and U14341 (N_14341,N_11327,N_9222);
xor U14342 (N_14342,N_9775,N_10967);
or U14343 (N_14343,N_9668,N_11587);
or U14344 (N_14344,N_10667,N_10966);
xor U14345 (N_14345,N_9276,N_10397);
xor U14346 (N_14346,N_10091,N_9343);
and U14347 (N_14347,N_10718,N_11027);
nor U14348 (N_14348,N_10125,N_9701);
and U14349 (N_14349,N_11213,N_10153);
nor U14350 (N_14350,N_11463,N_9941);
and U14351 (N_14351,N_11453,N_10471);
xnor U14352 (N_14352,N_11447,N_9821);
and U14353 (N_14353,N_11582,N_9488);
xor U14354 (N_14354,N_10681,N_10123);
nand U14355 (N_14355,N_11290,N_9329);
nand U14356 (N_14356,N_10300,N_9872);
and U14357 (N_14357,N_9247,N_10749);
nand U14358 (N_14358,N_9682,N_9267);
nor U14359 (N_14359,N_11856,N_11452);
and U14360 (N_14360,N_11675,N_9133);
and U14361 (N_14361,N_11325,N_11850);
nand U14362 (N_14362,N_11528,N_11448);
and U14363 (N_14363,N_10023,N_9190);
xor U14364 (N_14364,N_9527,N_9067);
xor U14365 (N_14365,N_10362,N_11427);
nand U14366 (N_14366,N_10015,N_11535);
and U14367 (N_14367,N_9900,N_10341);
nand U14368 (N_14368,N_10306,N_11968);
or U14369 (N_14369,N_9362,N_9777);
nand U14370 (N_14370,N_10047,N_10979);
nor U14371 (N_14371,N_10398,N_10116);
xnor U14372 (N_14372,N_10943,N_10969);
nor U14373 (N_14373,N_10963,N_10269);
xor U14374 (N_14374,N_9308,N_9554);
nand U14375 (N_14375,N_11444,N_10125);
xor U14376 (N_14376,N_10518,N_10349);
nor U14377 (N_14377,N_10627,N_10856);
and U14378 (N_14378,N_11532,N_9965);
or U14379 (N_14379,N_11460,N_9497);
nand U14380 (N_14380,N_9528,N_11625);
xor U14381 (N_14381,N_11183,N_11757);
or U14382 (N_14382,N_9221,N_11014);
or U14383 (N_14383,N_10334,N_11107);
and U14384 (N_14384,N_11754,N_11003);
xnor U14385 (N_14385,N_9582,N_10467);
xor U14386 (N_14386,N_11981,N_11044);
or U14387 (N_14387,N_9420,N_10602);
xor U14388 (N_14388,N_9944,N_11466);
and U14389 (N_14389,N_10410,N_11882);
nor U14390 (N_14390,N_10300,N_10448);
and U14391 (N_14391,N_10172,N_10431);
nand U14392 (N_14392,N_10221,N_11740);
or U14393 (N_14393,N_9490,N_11269);
xnor U14394 (N_14394,N_10084,N_9034);
nor U14395 (N_14395,N_9039,N_10978);
nand U14396 (N_14396,N_9579,N_10091);
or U14397 (N_14397,N_9686,N_9428);
or U14398 (N_14398,N_9414,N_11730);
nor U14399 (N_14399,N_11934,N_9762);
or U14400 (N_14400,N_10170,N_11517);
or U14401 (N_14401,N_10831,N_11064);
and U14402 (N_14402,N_11846,N_10438);
xnor U14403 (N_14403,N_9997,N_10683);
nand U14404 (N_14404,N_10142,N_9138);
and U14405 (N_14405,N_10675,N_9512);
nor U14406 (N_14406,N_11032,N_11012);
or U14407 (N_14407,N_10202,N_11818);
xor U14408 (N_14408,N_11391,N_11543);
nor U14409 (N_14409,N_9613,N_9428);
xnor U14410 (N_14410,N_10520,N_10711);
and U14411 (N_14411,N_9331,N_9782);
nand U14412 (N_14412,N_10487,N_9366);
or U14413 (N_14413,N_11840,N_11634);
nor U14414 (N_14414,N_11362,N_10794);
nor U14415 (N_14415,N_10026,N_9931);
nand U14416 (N_14416,N_10903,N_11192);
xor U14417 (N_14417,N_10154,N_10083);
nor U14418 (N_14418,N_9728,N_10489);
xor U14419 (N_14419,N_11526,N_11416);
or U14420 (N_14420,N_9012,N_9930);
and U14421 (N_14421,N_11051,N_9265);
and U14422 (N_14422,N_11126,N_9031);
xor U14423 (N_14423,N_9192,N_11935);
nand U14424 (N_14424,N_9993,N_11990);
xor U14425 (N_14425,N_9768,N_10604);
xor U14426 (N_14426,N_9286,N_9797);
nand U14427 (N_14427,N_11049,N_9289);
or U14428 (N_14428,N_11861,N_10060);
or U14429 (N_14429,N_11923,N_9565);
xnor U14430 (N_14430,N_11268,N_10260);
xor U14431 (N_14431,N_9560,N_11063);
xor U14432 (N_14432,N_10926,N_11763);
nand U14433 (N_14433,N_10658,N_9844);
nor U14434 (N_14434,N_9363,N_9052);
nand U14435 (N_14435,N_11929,N_10770);
xor U14436 (N_14436,N_9888,N_10190);
and U14437 (N_14437,N_10475,N_11098);
nor U14438 (N_14438,N_10890,N_10762);
or U14439 (N_14439,N_10136,N_10413);
nor U14440 (N_14440,N_9302,N_10438);
or U14441 (N_14441,N_11313,N_10181);
nand U14442 (N_14442,N_10770,N_9257);
xor U14443 (N_14443,N_11058,N_11602);
and U14444 (N_14444,N_11536,N_10763);
or U14445 (N_14445,N_9002,N_10227);
or U14446 (N_14446,N_10123,N_10021);
xnor U14447 (N_14447,N_9594,N_9115);
or U14448 (N_14448,N_9738,N_9413);
or U14449 (N_14449,N_9020,N_11753);
nor U14450 (N_14450,N_11410,N_9769);
nand U14451 (N_14451,N_9201,N_11645);
and U14452 (N_14452,N_10826,N_10772);
or U14453 (N_14453,N_11937,N_9717);
and U14454 (N_14454,N_9142,N_10849);
and U14455 (N_14455,N_11231,N_10413);
nand U14456 (N_14456,N_11576,N_11589);
xor U14457 (N_14457,N_11922,N_11344);
nor U14458 (N_14458,N_10999,N_10559);
xnor U14459 (N_14459,N_9234,N_10206);
xor U14460 (N_14460,N_11655,N_10837);
nor U14461 (N_14461,N_9829,N_10036);
nand U14462 (N_14462,N_9590,N_11301);
and U14463 (N_14463,N_9264,N_9813);
or U14464 (N_14464,N_10232,N_11204);
xor U14465 (N_14465,N_10459,N_10739);
xnor U14466 (N_14466,N_9447,N_9241);
or U14467 (N_14467,N_9416,N_11897);
nor U14468 (N_14468,N_9725,N_10517);
or U14469 (N_14469,N_9612,N_10167);
nor U14470 (N_14470,N_9527,N_9503);
nand U14471 (N_14471,N_10181,N_11064);
nor U14472 (N_14472,N_9080,N_11015);
or U14473 (N_14473,N_11352,N_11391);
or U14474 (N_14474,N_11672,N_11741);
xor U14475 (N_14475,N_9777,N_9074);
nor U14476 (N_14476,N_9696,N_10371);
nor U14477 (N_14477,N_10393,N_10059);
nand U14478 (N_14478,N_10477,N_9049);
and U14479 (N_14479,N_9139,N_11607);
xnor U14480 (N_14480,N_10175,N_10714);
xnor U14481 (N_14481,N_11023,N_10017);
nor U14482 (N_14482,N_10812,N_10162);
or U14483 (N_14483,N_10399,N_9578);
and U14484 (N_14484,N_10238,N_11142);
xnor U14485 (N_14485,N_10369,N_11084);
nand U14486 (N_14486,N_11164,N_10597);
nand U14487 (N_14487,N_10059,N_9939);
nand U14488 (N_14488,N_9825,N_9823);
nand U14489 (N_14489,N_11167,N_11539);
nand U14490 (N_14490,N_11926,N_10114);
xor U14491 (N_14491,N_9006,N_9217);
and U14492 (N_14492,N_11813,N_11914);
xnor U14493 (N_14493,N_11932,N_9234);
nand U14494 (N_14494,N_11247,N_9026);
nor U14495 (N_14495,N_9284,N_10331);
nor U14496 (N_14496,N_9387,N_10710);
nand U14497 (N_14497,N_9266,N_11959);
nand U14498 (N_14498,N_9457,N_9025);
or U14499 (N_14499,N_9720,N_10834);
or U14500 (N_14500,N_9644,N_11480);
nor U14501 (N_14501,N_10704,N_11471);
or U14502 (N_14502,N_10739,N_9241);
and U14503 (N_14503,N_10384,N_10180);
nand U14504 (N_14504,N_9255,N_10853);
xor U14505 (N_14505,N_9534,N_9079);
nor U14506 (N_14506,N_9058,N_11451);
or U14507 (N_14507,N_10450,N_9061);
or U14508 (N_14508,N_10549,N_11194);
or U14509 (N_14509,N_9848,N_9006);
xnor U14510 (N_14510,N_11255,N_9755);
nor U14511 (N_14511,N_11314,N_11785);
and U14512 (N_14512,N_10393,N_9360);
or U14513 (N_14513,N_11064,N_9729);
xnor U14514 (N_14514,N_9400,N_9398);
and U14515 (N_14515,N_11647,N_11197);
nand U14516 (N_14516,N_9917,N_10546);
nor U14517 (N_14517,N_11224,N_10628);
nand U14518 (N_14518,N_10024,N_10767);
nor U14519 (N_14519,N_10289,N_11097);
xor U14520 (N_14520,N_11110,N_10598);
or U14521 (N_14521,N_11563,N_11442);
and U14522 (N_14522,N_9363,N_9452);
or U14523 (N_14523,N_9950,N_11742);
nand U14524 (N_14524,N_11896,N_10719);
and U14525 (N_14525,N_11486,N_10041);
xor U14526 (N_14526,N_10783,N_11539);
or U14527 (N_14527,N_10752,N_11890);
nor U14528 (N_14528,N_9117,N_10868);
nor U14529 (N_14529,N_11446,N_11134);
xor U14530 (N_14530,N_9097,N_11025);
nand U14531 (N_14531,N_11434,N_9827);
xor U14532 (N_14532,N_11729,N_10485);
or U14533 (N_14533,N_10695,N_10631);
and U14534 (N_14534,N_9455,N_11683);
and U14535 (N_14535,N_11782,N_11807);
nand U14536 (N_14536,N_9615,N_10759);
and U14537 (N_14537,N_9294,N_11511);
or U14538 (N_14538,N_10312,N_10909);
nor U14539 (N_14539,N_10258,N_11384);
nor U14540 (N_14540,N_9751,N_10822);
nor U14541 (N_14541,N_10097,N_11240);
nor U14542 (N_14542,N_10739,N_11046);
xnor U14543 (N_14543,N_11359,N_10898);
xor U14544 (N_14544,N_9856,N_11733);
or U14545 (N_14545,N_11501,N_11572);
nand U14546 (N_14546,N_11768,N_9439);
xor U14547 (N_14547,N_9489,N_9685);
xnor U14548 (N_14548,N_10872,N_9212);
nand U14549 (N_14549,N_9660,N_9161);
nand U14550 (N_14550,N_9955,N_9292);
nor U14551 (N_14551,N_10623,N_10940);
and U14552 (N_14552,N_11679,N_9484);
nand U14553 (N_14553,N_11120,N_9010);
xnor U14554 (N_14554,N_11758,N_9666);
and U14555 (N_14555,N_10106,N_9345);
xor U14556 (N_14556,N_9995,N_9348);
or U14557 (N_14557,N_9572,N_10658);
xnor U14558 (N_14558,N_11740,N_9502);
xnor U14559 (N_14559,N_10116,N_11400);
and U14560 (N_14560,N_11361,N_9291);
xor U14561 (N_14561,N_10532,N_11285);
or U14562 (N_14562,N_10469,N_11806);
xnor U14563 (N_14563,N_9273,N_11213);
nand U14564 (N_14564,N_9068,N_9898);
nor U14565 (N_14565,N_11063,N_11664);
or U14566 (N_14566,N_9564,N_11176);
or U14567 (N_14567,N_11954,N_11271);
and U14568 (N_14568,N_9244,N_11112);
and U14569 (N_14569,N_9282,N_11659);
or U14570 (N_14570,N_11414,N_11969);
nor U14571 (N_14571,N_11452,N_10149);
and U14572 (N_14572,N_9276,N_11539);
xnor U14573 (N_14573,N_10409,N_11747);
nand U14574 (N_14574,N_11413,N_11902);
nand U14575 (N_14575,N_9940,N_9942);
or U14576 (N_14576,N_11077,N_9125);
xor U14577 (N_14577,N_11595,N_9481);
nor U14578 (N_14578,N_11009,N_9386);
nand U14579 (N_14579,N_10977,N_9844);
and U14580 (N_14580,N_10708,N_11389);
or U14581 (N_14581,N_9509,N_11166);
or U14582 (N_14582,N_10020,N_10767);
and U14583 (N_14583,N_11031,N_11915);
and U14584 (N_14584,N_11976,N_10320);
or U14585 (N_14585,N_9253,N_9784);
xor U14586 (N_14586,N_9257,N_9713);
nor U14587 (N_14587,N_9643,N_9303);
or U14588 (N_14588,N_10877,N_11352);
or U14589 (N_14589,N_9975,N_9849);
nand U14590 (N_14590,N_11620,N_11778);
or U14591 (N_14591,N_11961,N_10791);
and U14592 (N_14592,N_9644,N_10902);
nor U14593 (N_14593,N_10241,N_10074);
and U14594 (N_14594,N_10365,N_9835);
nand U14595 (N_14595,N_10277,N_10310);
xor U14596 (N_14596,N_10204,N_11524);
nor U14597 (N_14597,N_11093,N_10329);
or U14598 (N_14598,N_9558,N_10549);
and U14599 (N_14599,N_9870,N_9323);
nor U14600 (N_14600,N_10818,N_11853);
and U14601 (N_14601,N_11576,N_11843);
xnor U14602 (N_14602,N_10421,N_11043);
xor U14603 (N_14603,N_9205,N_9260);
or U14604 (N_14604,N_9310,N_9040);
nor U14605 (N_14605,N_10090,N_11614);
nor U14606 (N_14606,N_10253,N_9463);
nand U14607 (N_14607,N_9482,N_9585);
xor U14608 (N_14608,N_9251,N_9403);
nand U14609 (N_14609,N_11965,N_11858);
xor U14610 (N_14610,N_11881,N_11839);
and U14611 (N_14611,N_9071,N_9291);
and U14612 (N_14612,N_11207,N_10689);
and U14613 (N_14613,N_10979,N_10380);
xor U14614 (N_14614,N_9817,N_9523);
nor U14615 (N_14615,N_11238,N_11779);
nand U14616 (N_14616,N_9838,N_9919);
nand U14617 (N_14617,N_11079,N_9772);
nand U14618 (N_14618,N_10748,N_9129);
nand U14619 (N_14619,N_10337,N_9985);
and U14620 (N_14620,N_11837,N_10204);
or U14621 (N_14621,N_10647,N_11382);
or U14622 (N_14622,N_11248,N_10870);
xnor U14623 (N_14623,N_10642,N_11494);
or U14624 (N_14624,N_10800,N_10980);
xnor U14625 (N_14625,N_10872,N_9986);
nand U14626 (N_14626,N_10207,N_11699);
and U14627 (N_14627,N_9278,N_9056);
or U14628 (N_14628,N_11769,N_10407);
xnor U14629 (N_14629,N_11179,N_10882);
nand U14630 (N_14630,N_9436,N_9600);
xor U14631 (N_14631,N_10611,N_11712);
nor U14632 (N_14632,N_11382,N_10497);
xnor U14633 (N_14633,N_9067,N_11748);
nor U14634 (N_14634,N_9169,N_10097);
nor U14635 (N_14635,N_9222,N_11817);
nor U14636 (N_14636,N_9499,N_9007);
nor U14637 (N_14637,N_11316,N_10397);
or U14638 (N_14638,N_10563,N_11367);
xnor U14639 (N_14639,N_10535,N_11212);
nor U14640 (N_14640,N_10692,N_10016);
and U14641 (N_14641,N_10743,N_11674);
and U14642 (N_14642,N_10098,N_11315);
xnor U14643 (N_14643,N_11192,N_11768);
and U14644 (N_14644,N_9958,N_9414);
nor U14645 (N_14645,N_11007,N_9316);
xor U14646 (N_14646,N_11785,N_10254);
and U14647 (N_14647,N_10870,N_10685);
nand U14648 (N_14648,N_11024,N_9132);
xor U14649 (N_14649,N_11695,N_9649);
xor U14650 (N_14650,N_9200,N_9599);
xor U14651 (N_14651,N_11818,N_10683);
or U14652 (N_14652,N_11781,N_9432);
or U14653 (N_14653,N_9846,N_11987);
nand U14654 (N_14654,N_10703,N_10644);
nand U14655 (N_14655,N_10661,N_11228);
and U14656 (N_14656,N_10835,N_9261);
xnor U14657 (N_14657,N_11851,N_10919);
xnor U14658 (N_14658,N_9779,N_9248);
nand U14659 (N_14659,N_11123,N_9165);
and U14660 (N_14660,N_10683,N_11391);
and U14661 (N_14661,N_9896,N_9522);
xnor U14662 (N_14662,N_9555,N_11123);
or U14663 (N_14663,N_9577,N_11862);
and U14664 (N_14664,N_11247,N_11745);
nand U14665 (N_14665,N_9829,N_9543);
nand U14666 (N_14666,N_10121,N_9520);
xor U14667 (N_14667,N_9875,N_11703);
and U14668 (N_14668,N_11114,N_9056);
and U14669 (N_14669,N_11980,N_11988);
or U14670 (N_14670,N_11871,N_10900);
xor U14671 (N_14671,N_10354,N_10854);
xnor U14672 (N_14672,N_10074,N_10491);
nand U14673 (N_14673,N_10860,N_11430);
nor U14674 (N_14674,N_9351,N_11065);
xnor U14675 (N_14675,N_11740,N_9400);
and U14676 (N_14676,N_9314,N_10891);
xnor U14677 (N_14677,N_11160,N_10078);
or U14678 (N_14678,N_11208,N_9211);
or U14679 (N_14679,N_11552,N_9582);
and U14680 (N_14680,N_11093,N_10837);
or U14681 (N_14681,N_11156,N_11794);
or U14682 (N_14682,N_10554,N_9037);
and U14683 (N_14683,N_11684,N_11656);
xor U14684 (N_14684,N_10093,N_11525);
nand U14685 (N_14685,N_9082,N_9667);
nand U14686 (N_14686,N_10012,N_10645);
or U14687 (N_14687,N_9363,N_11825);
xor U14688 (N_14688,N_10270,N_10081);
nand U14689 (N_14689,N_9887,N_9533);
nor U14690 (N_14690,N_10384,N_10297);
nor U14691 (N_14691,N_11640,N_10497);
xnor U14692 (N_14692,N_11511,N_10443);
and U14693 (N_14693,N_11182,N_10644);
and U14694 (N_14694,N_10757,N_9749);
xnor U14695 (N_14695,N_10749,N_9854);
nor U14696 (N_14696,N_11358,N_9091);
or U14697 (N_14697,N_10532,N_11640);
and U14698 (N_14698,N_10427,N_10279);
xor U14699 (N_14699,N_11009,N_9611);
nor U14700 (N_14700,N_9012,N_10809);
nor U14701 (N_14701,N_9746,N_10031);
nand U14702 (N_14702,N_9803,N_10064);
and U14703 (N_14703,N_11984,N_11550);
xnor U14704 (N_14704,N_9893,N_9874);
nor U14705 (N_14705,N_11218,N_11621);
xnor U14706 (N_14706,N_9435,N_9562);
nor U14707 (N_14707,N_10089,N_9141);
xor U14708 (N_14708,N_11958,N_11231);
or U14709 (N_14709,N_10998,N_10053);
nor U14710 (N_14710,N_10382,N_9315);
and U14711 (N_14711,N_9461,N_11879);
or U14712 (N_14712,N_11020,N_9385);
and U14713 (N_14713,N_11605,N_10128);
xnor U14714 (N_14714,N_11785,N_11064);
nand U14715 (N_14715,N_10723,N_11998);
nand U14716 (N_14716,N_11794,N_9082);
and U14717 (N_14717,N_10968,N_10661);
xor U14718 (N_14718,N_11466,N_11844);
or U14719 (N_14719,N_10554,N_10517);
or U14720 (N_14720,N_9434,N_10713);
nand U14721 (N_14721,N_11375,N_10910);
nand U14722 (N_14722,N_9425,N_9831);
xnor U14723 (N_14723,N_9876,N_9545);
nor U14724 (N_14724,N_10931,N_9538);
and U14725 (N_14725,N_11863,N_9799);
nand U14726 (N_14726,N_9763,N_10846);
nor U14727 (N_14727,N_10941,N_11648);
xnor U14728 (N_14728,N_11214,N_11907);
xnor U14729 (N_14729,N_11492,N_9484);
nand U14730 (N_14730,N_9678,N_11513);
nor U14731 (N_14731,N_9037,N_11665);
and U14732 (N_14732,N_9913,N_11360);
nor U14733 (N_14733,N_11367,N_11582);
xnor U14734 (N_14734,N_11228,N_11745);
and U14735 (N_14735,N_9108,N_9250);
xnor U14736 (N_14736,N_10667,N_11305);
nor U14737 (N_14737,N_10833,N_9123);
and U14738 (N_14738,N_11730,N_11849);
nor U14739 (N_14739,N_10884,N_10550);
or U14740 (N_14740,N_11480,N_10710);
or U14741 (N_14741,N_11449,N_9250);
xor U14742 (N_14742,N_10828,N_11590);
and U14743 (N_14743,N_9462,N_11698);
or U14744 (N_14744,N_10761,N_9173);
nor U14745 (N_14745,N_9756,N_11651);
nor U14746 (N_14746,N_10839,N_11838);
and U14747 (N_14747,N_11494,N_11342);
and U14748 (N_14748,N_11377,N_11686);
nand U14749 (N_14749,N_11629,N_11139);
xnor U14750 (N_14750,N_10413,N_9012);
xnor U14751 (N_14751,N_11900,N_11592);
or U14752 (N_14752,N_9174,N_9404);
xor U14753 (N_14753,N_10805,N_11092);
nor U14754 (N_14754,N_9215,N_9759);
xor U14755 (N_14755,N_11676,N_9313);
nand U14756 (N_14756,N_10929,N_10927);
or U14757 (N_14757,N_11363,N_11372);
and U14758 (N_14758,N_10909,N_11514);
or U14759 (N_14759,N_9865,N_9842);
nor U14760 (N_14760,N_10739,N_10693);
or U14761 (N_14761,N_10287,N_9573);
xor U14762 (N_14762,N_10210,N_10747);
nor U14763 (N_14763,N_11453,N_11792);
or U14764 (N_14764,N_11844,N_11567);
nor U14765 (N_14765,N_11688,N_11759);
xnor U14766 (N_14766,N_9590,N_11799);
xnor U14767 (N_14767,N_9715,N_10050);
or U14768 (N_14768,N_11167,N_10625);
xnor U14769 (N_14769,N_11033,N_11771);
nor U14770 (N_14770,N_9096,N_10801);
or U14771 (N_14771,N_9783,N_10774);
or U14772 (N_14772,N_10729,N_11622);
nor U14773 (N_14773,N_9477,N_11565);
xor U14774 (N_14774,N_10068,N_9145);
nand U14775 (N_14775,N_10170,N_11556);
or U14776 (N_14776,N_9659,N_11414);
or U14777 (N_14777,N_10672,N_9134);
xnor U14778 (N_14778,N_9941,N_10755);
nor U14779 (N_14779,N_9863,N_10421);
and U14780 (N_14780,N_11875,N_10086);
xnor U14781 (N_14781,N_9104,N_11200);
nand U14782 (N_14782,N_10133,N_11169);
and U14783 (N_14783,N_10320,N_9054);
xor U14784 (N_14784,N_11324,N_11246);
nor U14785 (N_14785,N_10241,N_9775);
nor U14786 (N_14786,N_9569,N_11002);
or U14787 (N_14787,N_9778,N_9243);
xor U14788 (N_14788,N_9352,N_11369);
and U14789 (N_14789,N_11867,N_11634);
xor U14790 (N_14790,N_11987,N_10152);
and U14791 (N_14791,N_10652,N_10955);
nand U14792 (N_14792,N_10888,N_9007);
xnor U14793 (N_14793,N_9693,N_11901);
and U14794 (N_14794,N_9511,N_11541);
and U14795 (N_14795,N_10359,N_10564);
and U14796 (N_14796,N_9476,N_11319);
or U14797 (N_14797,N_9198,N_9173);
nor U14798 (N_14798,N_11714,N_10835);
and U14799 (N_14799,N_11666,N_11554);
or U14800 (N_14800,N_9334,N_10632);
xor U14801 (N_14801,N_10934,N_11031);
or U14802 (N_14802,N_10728,N_11384);
nand U14803 (N_14803,N_9797,N_11507);
or U14804 (N_14804,N_9009,N_10569);
nand U14805 (N_14805,N_10272,N_11707);
nand U14806 (N_14806,N_9867,N_9208);
xor U14807 (N_14807,N_10368,N_10807);
and U14808 (N_14808,N_10022,N_11179);
xor U14809 (N_14809,N_10396,N_10391);
and U14810 (N_14810,N_10195,N_10480);
nor U14811 (N_14811,N_10222,N_11418);
xor U14812 (N_14812,N_9053,N_9965);
or U14813 (N_14813,N_9762,N_9276);
xor U14814 (N_14814,N_10366,N_11978);
nor U14815 (N_14815,N_10566,N_10373);
and U14816 (N_14816,N_11791,N_10304);
nand U14817 (N_14817,N_11414,N_11635);
nor U14818 (N_14818,N_11383,N_10922);
nor U14819 (N_14819,N_9602,N_9960);
and U14820 (N_14820,N_9948,N_11405);
nand U14821 (N_14821,N_11608,N_10641);
xor U14822 (N_14822,N_10808,N_11932);
nand U14823 (N_14823,N_10069,N_10911);
nand U14824 (N_14824,N_9927,N_9969);
and U14825 (N_14825,N_9135,N_10467);
nand U14826 (N_14826,N_11341,N_10111);
and U14827 (N_14827,N_11717,N_11481);
or U14828 (N_14828,N_10711,N_9353);
and U14829 (N_14829,N_11910,N_9570);
nor U14830 (N_14830,N_10626,N_9146);
nand U14831 (N_14831,N_10759,N_9177);
or U14832 (N_14832,N_11751,N_10260);
xor U14833 (N_14833,N_11294,N_11818);
xnor U14834 (N_14834,N_11464,N_10539);
and U14835 (N_14835,N_9654,N_9030);
xor U14836 (N_14836,N_10690,N_10827);
or U14837 (N_14837,N_9470,N_9023);
xnor U14838 (N_14838,N_11417,N_9261);
or U14839 (N_14839,N_11968,N_9763);
or U14840 (N_14840,N_9877,N_11013);
or U14841 (N_14841,N_9399,N_9132);
nand U14842 (N_14842,N_9019,N_11300);
or U14843 (N_14843,N_11734,N_9038);
nor U14844 (N_14844,N_9118,N_9627);
or U14845 (N_14845,N_10214,N_11449);
xnor U14846 (N_14846,N_9846,N_10403);
nand U14847 (N_14847,N_10346,N_11150);
xor U14848 (N_14848,N_9965,N_10700);
nand U14849 (N_14849,N_10126,N_10978);
nor U14850 (N_14850,N_11981,N_9591);
nand U14851 (N_14851,N_9044,N_10395);
or U14852 (N_14852,N_11162,N_10469);
xor U14853 (N_14853,N_11820,N_9261);
nand U14854 (N_14854,N_11831,N_11693);
xor U14855 (N_14855,N_9924,N_11131);
nor U14856 (N_14856,N_10281,N_9293);
and U14857 (N_14857,N_9299,N_9480);
nand U14858 (N_14858,N_11937,N_9359);
nor U14859 (N_14859,N_10423,N_11296);
nor U14860 (N_14860,N_9474,N_10941);
nor U14861 (N_14861,N_9868,N_10956);
and U14862 (N_14862,N_10165,N_9428);
nor U14863 (N_14863,N_9785,N_9815);
nand U14864 (N_14864,N_10824,N_9691);
and U14865 (N_14865,N_9103,N_9435);
or U14866 (N_14866,N_10396,N_10106);
or U14867 (N_14867,N_10711,N_9989);
and U14868 (N_14868,N_11001,N_9724);
xnor U14869 (N_14869,N_11381,N_11966);
nor U14870 (N_14870,N_10780,N_9342);
nor U14871 (N_14871,N_10471,N_9428);
nor U14872 (N_14872,N_11894,N_11336);
xor U14873 (N_14873,N_9015,N_9209);
xnor U14874 (N_14874,N_10741,N_10755);
nand U14875 (N_14875,N_9278,N_10419);
xor U14876 (N_14876,N_11786,N_9887);
nor U14877 (N_14877,N_10693,N_11595);
nand U14878 (N_14878,N_11579,N_9065);
nor U14879 (N_14879,N_11563,N_10097);
or U14880 (N_14880,N_9222,N_9395);
and U14881 (N_14881,N_11254,N_9996);
xor U14882 (N_14882,N_9943,N_10775);
nand U14883 (N_14883,N_11041,N_11181);
xnor U14884 (N_14884,N_9024,N_9956);
or U14885 (N_14885,N_9912,N_10622);
nand U14886 (N_14886,N_11667,N_9428);
nor U14887 (N_14887,N_9509,N_11089);
or U14888 (N_14888,N_9835,N_9733);
and U14889 (N_14889,N_11472,N_9780);
nor U14890 (N_14890,N_10556,N_11401);
nor U14891 (N_14891,N_10441,N_9847);
nand U14892 (N_14892,N_9778,N_11966);
nand U14893 (N_14893,N_11356,N_9725);
nor U14894 (N_14894,N_9517,N_10746);
or U14895 (N_14895,N_10695,N_11498);
nand U14896 (N_14896,N_9405,N_9016);
nand U14897 (N_14897,N_11202,N_9418);
and U14898 (N_14898,N_10542,N_9728);
nor U14899 (N_14899,N_11381,N_10515);
xor U14900 (N_14900,N_11807,N_10258);
nor U14901 (N_14901,N_9910,N_9855);
xnor U14902 (N_14902,N_10856,N_10479);
nand U14903 (N_14903,N_11036,N_10221);
xnor U14904 (N_14904,N_11831,N_11048);
nand U14905 (N_14905,N_11331,N_10770);
or U14906 (N_14906,N_10292,N_9187);
nor U14907 (N_14907,N_9621,N_10287);
xor U14908 (N_14908,N_11641,N_10057);
xor U14909 (N_14909,N_9674,N_11718);
or U14910 (N_14910,N_9149,N_11308);
or U14911 (N_14911,N_9392,N_11466);
xnor U14912 (N_14912,N_11692,N_11624);
or U14913 (N_14913,N_10153,N_10291);
and U14914 (N_14914,N_11200,N_9823);
nor U14915 (N_14915,N_9975,N_9224);
nor U14916 (N_14916,N_11099,N_10388);
nand U14917 (N_14917,N_11331,N_11158);
or U14918 (N_14918,N_10995,N_9976);
nor U14919 (N_14919,N_11505,N_10019);
and U14920 (N_14920,N_10868,N_11204);
xnor U14921 (N_14921,N_11323,N_9049);
and U14922 (N_14922,N_9367,N_9452);
nor U14923 (N_14923,N_10514,N_10310);
or U14924 (N_14924,N_11348,N_10592);
xnor U14925 (N_14925,N_10210,N_11799);
nand U14926 (N_14926,N_11154,N_10453);
or U14927 (N_14927,N_11982,N_9615);
nor U14928 (N_14928,N_9650,N_9489);
nor U14929 (N_14929,N_9270,N_9878);
nand U14930 (N_14930,N_11495,N_9577);
nand U14931 (N_14931,N_11345,N_10237);
and U14932 (N_14932,N_9302,N_9891);
nand U14933 (N_14933,N_9777,N_11952);
nor U14934 (N_14934,N_10526,N_11095);
xor U14935 (N_14935,N_11336,N_10610);
xnor U14936 (N_14936,N_10106,N_10525);
or U14937 (N_14937,N_9903,N_10407);
xor U14938 (N_14938,N_9330,N_11131);
nand U14939 (N_14939,N_10657,N_11810);
xor U14940 (N_14940,N_9524,N_9871);
or U14941 (N_14941,N_10968,N_9473);
and U14942 (N_14942,N_9187,N_9279);
or U14943 (N_14943,N_11553,N_11446);
xnor U14944 (N_14944,N_9834,N_9894);
nor U14945 (N_14945,N_10193,N_10646);
nand U14946 (N_14946,N_10048,N_9578);
nand U14947 (N_14947,N_9288,N_9307);
nand U14948 (N_14948,N_9514,N_9422);
or U14949 (N_14949,N_9801,N_10216);
or U14950 (N_14950,N_9692,N_9529);
nor U14951 (N_14951,N_11784,N_9066);
xor U14952 (N_14952,N_10348,N_9615);
nand U14953 (N_14953,N_10421,N_11837);
or U14954 (N_14954,N_9941,N_11950);
nand U14955 (N_14955,N_11651,N_10984);
nand U14956 (N_14956,N_9412,N_10862);
xor U14957 (N_14957,N_10833,N_11115);
nand U14958 (N_14958,N_10019,N_11088);
or U14959 (N_14959,N_10910,N_9967);
and U14960 (N_14960,N_9986,N_10829);
xnor U14961 (N_14961,N_11627,N_10161);
nor U14962 (N_14962,N_10622,N_10853);
and U14963 (N_14963,N_10405,N_11979);
nand U14964 (N_14964,N_9633,N_10107);
nor U14965 (N_14965,N_9302,N_11417);
or U14966 (N_14966,N_9288,N_10260);
nor U14967 (N_14967,N_9776,N_11212);
nor U14968 (N_14968,N_9668,N_9357);
and U14969 (N_14969,N_10540,N_9826);
xnor U14970 (N_14970,N_11476,N_9083);
and U14971 (N_14971,N_10394,N_9882);
or U14972 (N_14972,N_9732,N_9638);
and U14973 (N_14973,N_9343,N_11299);
nor U14974 (N_14974,N_9603,N_9859);
or U14975 (N_14975,N_9020,N_9770);
nand U14976 (N_14976,N_9525,N_10662);
or U14977 (N_14977,N_10993,N_10742);
xnor U14978 (N_14978,N_10086,N_11579);
nand U14979 (N_14979,N_11732,N_9080);
or U14980 (N_14980,N_9784,N_10805);
xnor U14981 (N_14981,N_9886,N_9061);
or U14982 (N_14982,N_11665,N_10209);
nor U14983 (N_14983,N_9316,N_10904);
nand U14984 (N_14984,N_11886,N_9259);
xor U14985 (N_14985,N_10744,N_11628);
or U14986 (N_14986,N_11836,N_11658);
xnor U14987 (N_14987,N_11562,N_11298);
and U14988 (N_14988,N_11522,N_11631);
nand U14989 (N_14989,N_10864,N_9677);
or U14990 (N_14990,N_11646,N_10087);
nand U14991 (N_14991,N_11879,N_11172);
or U14992 (N_14992,N_11147,N_11815);
nand U14993 (N_14993,N_11589,N_11901);
nand U14994 (N_14994,N_10146,N_10637);
xnor U14995 (N_14995,N_10575,N_10348);
and U14996 (N_14996,N_11258,N_10553);
or U14997 (N_14997,N_10177,N_9409);
xnor U14998 (N_14998,N_10347,N_11937);
and U14999 (N_14999,N_9272,N_9119);
nor UO_0 (O_0,N_13899,N_13982);
or UO_1 (O_1,N_14980,N_13490);
nor UO_2 (O_2,N_13848,N_14084);
nand UO_3 (O_3,N_12422,N_12447);
and UO_4 (O_4,N_12553,N_13505);
and UO_5 (O_5,N_13780,N_13748);
or UO_6 (O_6,N_14233,N_12647);
and UO_7 (O_7,N_14875,N_12194);
xnor UO_8 (O_8,N_14096,N_13768);
and UO_9 (O_9,N_14365,N_12236);
nor UO_10 (O_10,N_13511,N_12469);
and UO_11 (O_11,N_13064,N_14940);
xor UO_12 (O_12,N_12744,N_13143);
nor UO_13 (O_13,N_13335,N_14874);
or UO_14 (O_14,N_14291,N_14195);
or UO_15 (O_15,N_13433,N_14660);
xnor UO_16 (O_16,N_14804,N_12839);
or UO_17 (O_17,N_12097,N_14871);
xnor UO_18 (O_18,N_12090,N_13874);
or UO_19 (O_19,N_14974,N_12063);
xnor UO_20 (O_20,N_13018,N_14171);
or UO_21 (O_21,N_14080,N_12737);
nor UO_22 (O_22,N_12154,N_13261);
or UO_23 (O_23,N_12809,N_14077);
nor UO_24 (O_24,N_14833,N_14008);
or UO_25 (O_25,N_13041,N_12257);
or UO_26 (O_26,N_13167,N_13029);
nor UO_27 (O_27,N_14919,N_14123);
nor UO_28 (O_28,N_14458,N_13249);
nor UO_29 (O_29,N_12437,N_12598);
or UO_30 (O_30,N_14081,N_14067);
nor UO_31 (O_31,N_12901,N_14167);
or UO_32 (O_32,N_13668,N_12274);
nand UO_33 (O_33,N_12178,N_12108);
nand UO_34 (O_34,N_12416,N_13156);
nor UO_35 (O_35,N_14714,N_14961);
nor UO_36 (O_36,N_13763,N_12112);
xnor UO_37 (O_37,N_13749,N_13783);
nor UO_38 (O_38,N_14684,N_12440);
and UO_39 (O_39,N_12244,N_14633);
and UO_40 (O_40,N_13286,N_12654);
nor UO_41 (O_41,N_12894,N_14929);
nor UO_42 (O_42,N_14032,N_12708);
and UO_43 (O_43,N_14103,N_13451);
nor UO_44 (O_44,N_12045,N_13546);
or UO_45 (O_45,N_13788,N_13761);
nand UO_46 (O_46,N_14773,N_12648);
xor UO_47 (O_47,N_13195,N_12566);
nor UO_48 (O_48,N_12495,N_12327);
nor UO_49 (O_49,N_13208,N_12914);
nand UO_50 (O_50,N_14581,N_13804);
or UO_51 (O_51,N_12070,N_14055);
nor UO_52 (O_52,N_12129,N_14087);
nand UO_53 (O_53,N_13694,N_14512);
xnor UO_54 (O_54,N_13497,N_12599);
xnor UO_55 (O_55,N_14223,N_12775);
and UO_56 (O_56,N_14631,N_13627);
nand UO_57 (O_57,N_13680,N_12199);
nor UO_58 (O_58,N_13913,N_14105);
nand UO_59 (O_59,N_13199,N_14457);
and UO_60 (O_60,N_14554,N_12740);
or UO_61 (O_61,N_13098,N_13320);
and UO_62 (O_62,N_13103,N_13082);
and UO_63 (O_63,N_13206,N_12111);
or UO_64 (O_64,N_12823,N_13990);
and UO_65 (O_65,N_12197,N_13213);
and UO_66 (O_66,N_12774,N_12915);
xor UO_67 (O_67,N_14001,N_14187);
nand UO_68 (O_68,N_12237,N_12000);
xnor UO_69 (O_69,N_13328,N_14518);
or UO_70 (O_70,N_13678,N_13922);
and UO_71 (O_71,N_14686,N_12443);
or UO_72 (O_72,N_12463,N_13622);
nand UO_73 (O_73,N_12337,N_13309);
nor UO_74 (O_74,N_12867,N_14572);
xnor UO_75 (O_75,N_13608,N_14138);
xnor UO_76 (O_76,N_12816,N_12455);
or UO_77 (O_77,N_14226,N_14054);
xnor UO_78 (O_78,N_14827,N_12876);
and UO_79 (O_79,N_14030,N_14824);
nand UO_80 (O_80,N_12946,N_13991);
and UO_81 (O_81,N_12052,N_13332);
nor UO_82 (O_82,N_14320,N_12082);
nand UO_83 (O_83,N_12355,N_12672);
or UO_84 (O_84,N_12940,N_12509);
or UO_85 (O_85,N_13532,N_14795);
or UO_86 (O_86,N_14580,N_14748);
or UO_87 (O_87,N_13220,N_14786);
nand UO_88 (O_88,N_13515,N_14693);
nor UO_89 (O_89,N_13541,N_13701);
nor UO_90 (O_90,N_12342,N_13579);
and UO_91 (O_91,N_13814,N_13355);
nor UO_92 (O_92,N_12323,N_13056);
nand UO_93 (O_93,N_12214,N_12033);
nand UO_94 (O_94,N_14937,N_13354);
xor UO_95 (O_95,N_13853,N_12726);
and UO_96 (O_96,N_12467,N_12472);
or UO_97 (O_97,N_12164,N_12375);
nor UO_98 (O_98,N_12360,N_12717);
or UO_99 (O_99,N_12021,N_12427);
nor UO_100 (O_100,N_13581,N_14578);
nor UO_101 (O_101,N_14391,N_13284);
and UO_102 (O_102,N_12292,N_14606);
xor UO_103 (O_103,N_13821,N_13154);
nand UO_104 (O_104,N_12275,N_12367);
xnor UO_105 (O_105,N_12724,N_13767);
nand UO_106 (O_106,N_12736,N_13770);
or UO_107 (O_107,N_13996,N_13194);
or UO_108 (O_108,N_13023,N_14479);
nand UO_109 (O_109,N_12528,N_13402);
and UO_110 (O_110,N_12419,N_12895);
nand UO_111 (O_111,N_13221,N_12564);
nand UO_112 (O_112,N_14825,N_12067);
or UO_113 (O_113,N_13090,N_12746);
xnor UO_114 (O_114,N_13021,N_12686);
xor UO_115 (O_115,N_14037,N_12857);
nor UO_116 (O_116,N_14869,N_13462);
and UO_117 (O_117,N_13383,N_14925);
nand UO_118 (O_118,N_14627,N_14445);
or UO_119 (O_119,N_12168,N_13431);
xnor UO_120 (O_120,N_13096,N_14230);
and UO_121 (O_121,N_14299,N_14254);
or UO_122 (O_122,N_14735,N_14311);
and UO_123 (O_123,N_13429,N_12403);
xor UO_124 (O_124,N_12673,N_12372);
nand UO_125 (O_125,N_13455,N_14890);
and UO_126 (O_126,N_13440,N_12718);
and UO_127 (O_127,N_12379,N_14726);
or UO_128 (O_128,N_14115,N_12478);
nand UO_129 (O_129,N_13474,N_13258);
nor UO_130 (O_130,N_14927,N_13447);
and UO_131 (O_131,N_12976,N_13074);
nand UO_132 (O_132,N_13227,N_13902);
nand UO_133 (O_133,N_14677,N_13673);
and UO_134 (O_134,N_14489,N_12661);
and UO_135 (O_135,N_14826,N_12698);
xor UO_136 (O_136,N_14165,N_12623);
xor UO_137 (O_137,N_13507,N_13252);
nand UO_138 (O_138,N_13719,N_14352);
or UO_139 (O_139,N_14351,N_12757);
xor UO_140 (O_140,N_13285,N_12973);
or UO_141 (O_141,N_13594,N_14800);
xnor UO_142 (O_142,N_13959,N_13311);
and UO_143 (O_143,N_12691,N_12578);
nor UO_144 (O_144,N_12974,N_12295);
and UO_145 (O_145,N_12435,N_12493);
nand UO_146 (O_146,N_12822,N_13563);
or UO_147 (O_147,N_14011,N_13501);
or UO_148 (O_148,N_12605,N_12119);
nand UO_149 (O_149,N_12808,N_14500);
and UO_150 (O_150,N_13796,N_12346);
xnor UO_151 (O_151,N_13831,N_12273);
or UO_152 (O_152,N_14034,N_14889);
xnor UO_153 (O_153,N_12017,N_12653);
or UO_154 (O_154,N_12238,N_14955);
xor UO_155 (O_155,N_14375,N_14117);
nand UO_156 (O_156,N_13629,N_13560);
or UO_157 (O_157,N_12591,N_13549);
nand UO_158 (O_158,N_14136,N_14013);
nor UO_159 (O_159,N_12428,N_13747);
xor UO_160 (O_160,N_14381,N_14740);
and UO_161 (O_161,N_13260,N_14215);
nor UO_162 (O_162,N_13139,N_12968);
nor UO_163 (O_163,N_12335,N_13979);
nor UO_164 (O_164,N_12460,N_13779);
xor UO_165 (O_165,N_12999,N_12320);
nand UO_166 (O_166,N_14367,N_13508);
nor UO_167 (O_167,N_14732,N_14917);
and UO_168 (O_168,N_12415,N_12056);
nand UO_169 (O_169,N_12889,N_12036);
and UO_170 (O_170,N_13793,N_13007);
nor UO_171 (O_171,N_13245,N_14396);
or UO_172 (O_172,N_14066,N_12747);
or UO_173 (O_173,N_14569,N_14023);
nor UO_174 (O_174,N_12414,N_12870);
nor UO_175 (O_175,N_13444,N_13114);
xnor UO_176 (O_176,N_14941,N_12265);
nor UO_177 (O_177,N_13461,N_12436);
and UO_178 (O_178,N_14177,N_13215);
nor UO_179 (O_179,N_13304,N_12219);
nor UO_180 (O_180,N_14624,N_13346);
nand UO_181 (O_181,N_12312,N_13476);
and UO_182 (O_182,N_13906,N_13281);
and UO_183 (O_183,N_12583,N_13843);
nand UO_184 (O_184,N_13870,N_12719);
nor UO_185 (O_185,N_14471,N_13319);
nor UO_186 (O_186,N_12992,N_12473);
and UO_187 (O_187,N_14607,N_13127);
nor UO_188 (O_188,N_14547,N_12608);
xor UO_189 (O_189,N_14993,N_13192);
and UO_190 (O_190,N_13027,N_12484);
and UO_191 (O_191,N_14106,N_13610);
xnor UO_192 (O_192,N_14621,N_12853);
or UO_193 (O_193,N_13813,N_14611);
xor UO_194 (O_194,N_12296,N_12301);
nand UO_195 (O_195,N_14543,N_12147);
nand UO_196 (O_196,N_14027,N_12169);
and UO_197 (O_197,N_12030,N_13801);
or UO_198 (O_198,N_12878,N_14753);
and UO_199 (O_199,N_12964,N_13299);
nand UO_200 (O_200,N_14002,N_13233);
and UO_201 (O_201,N_14022,N_14112);
nor UO_202 (O_202,N_13479,N_13115);
nand UO_203 (O_203,N_14775,N_13120);
and UO_204 (O_204,N_13604,N_13720);
nand UO_205 (O_205,N_12622,N_13099);
nand UO_206 (O_206,N_12924,N_12777);
or UO_207 (O_207,N_14522,N_12303);
xor UO_208 (O_208,N_13070,N_13240);
and UO_209 (O_209,N_12184,N_13693);
or UO_210 (O_210,N_12785,N_14092);
xor UO_211 (O_211,N_13058,N_14741);
xnor UO_212 (O_212,N_14549,N_12887);
nor UO_213 (O_213,N_12015,N_13280);
xor UO_214 (O_214,N_14636,N_14082);
nor UO_215 (O_215,N_14063,N_12358);
or UO_216 (O_216,N_13205,N_13995);
or UO_217 (O_217,N_13081,N_12242);
and UO_218 (O_218,N_12179,N_13266);
nor UO_219 (O_219,N_14809,N_14987);
nand UO_220 (O_220,N_13264,N_12374);
or UO_221 (O_221,N_13956,N_13651);
xnor UO_222 (O_222,N_14563,N_12629);
and UO_223 (O_223,N_13835,N_12364);
or UO_224 (O_224,N_14959,N_13772);
nor UO_225 (O_225,N_13924,N_14407);
xnor UO_226 (O_226,N_12318,N_14279);
nor UO_227 (O_227,N_14336,N_13318);
nand UO_228 (O_228,N_14520,N_14348);
and UO_229 (O_229,N_13690,N_13002);
nand UO_230 (O_230,N_13443,N_13117);
xnor UO_231 (O_231,N_14900,N_13689);
or UO_232 (O_232,N_13411,N_12798);
nand UO_233 (O_233,N_12313,N_14615);
and UO_234 (O_234,N_14237,N_14573);
nor UO_235 (O_235,N_12165,N_13614);
xor UO_236 (O_236,N_13174,N_14628);
and UO_237 (O_237,N_12571,N_13184);
and UO_238 (O_238,N_12175,N_13055);
or UO_239 (O_239,N_12287,N_13800);
nor UO_240 (O_240,N_12211,N_12170);
and UO_241 (O_241,N_13238,N_12700);
and UO_242 (O_242,N_13438,N_14700);
nor UO_243 (O_243,N_12558,N_12347);
nor UO_244 (O_244,N_13279,N_14224);
or UO_245 (O_245,N_13527,N_14467);
or UO_246 (O_246,N_12842,N_12424);
nand UO_247 (O_247,N_13083,N_13970);
and UO_248 (O_248,N_12458,N_12250);
nor UO_249 (O_249,N_14702,N_14613);
nor UO_250 (O_250,N_12146,N_12457);
and UO_251 (O_251,N_12247,N_13726);
xnor UO_252 (O_252,N_13186,N_12567);
nand UO_253 (O_253,N_14250,N_12863);
nand UO_254 (O_254,N_14951,N_13412);
and UO_255 (O_255,N_12202,N_14413);
xnor UO_256 (O_256,N_13542,N_13927);
xor UO_257 (O_257,N_14293,N_12105);
xor UO_258 (O_258,N_14946,N_14172);
and UO_259 (O_259,N_12064,N_12779);
xnor UO_260 (O_260,N_14059,N_12961);
xnor UO_261 (O_261,N_14932,N_13562);
xnor UO_262 (O_262,N_14368,N_12134);
or UO_263 (O_263,N_14409,N_14446);
nand UO_264 (O_264,N_12204,N_13672);
and UO_265 (O_265,N_14026,N_13964);
nor UO_266 (O_266,N_14425,N_14767);
and UO_267 (O_267,N_13949,N_14160);
and UO_268 (O_268,N_12353,N_12288);
nor UO_269 (O_269,N_14745,N_14854);
or UO_270 (O_270,N_12444,N_13375);
or UO_271 (O_271,N_14733,N_14857);
xnor UO_272 (O_272,N_13528,N_13308);
and UO_273 (O_273,N_12908,N_12882);
xnor UO_274 (O_274,N_14072,N_12910);
or UO_275 (O_275,N_12299,N_13307);
xnor UO_276 (O_276,N_13535,N_14738);
xor UO_277 (O_277,N_14286,N_13269);
nand UO_278 (O_278,N_14899,N_13583);
nand UO_279 (O_279,N_12087,N_13357);
nor UO_280 (O_280,N_13567,N_12019);
nor UO_281 (O_281,N_12276,N_12307);
nor UO_282 (O_282,N_12368,N_14156);
nor UO_283 (O_283,N_12573,N_13921);
xor UO_284 (O_284,N_14596,N_12640);
xnor UO_285 (O_285,N_13519,N_13033);
and UO_286 (O_286,N_13934,N_12480);
or UO_287 (O_287,N_13773,N_13551);
or UO_288 (O_288,N_13926,N_13262);
nor UO_289 (O_289,N_14464,N_13126);
nor UO_290 (O_290,N_14670,N_12471);
or UO_291 (O_291,N_13047,N_13868);
nand UO_292 (O_292,N_14043,N_12268);
or UO_293 (O_293,N_14537,N_12084);
xor UO_294 (O_294,N_13432,N_13534);
nor UO_295 (O_295,N_12972,N_14546);
or UO_296 (O_296,N_14759,N_13645);
or UO_297 (O_297,N_14594,N_12426);
nand UO_298 (O_298,N_14124,N_13282);
or UO_299 (O_299,N_13175,N_13569);
or UO_300 (O_300,N_13172,N_14189);
xor UO_301 (O_301,N_12462,N_13166);
or UO_302 (O_302,N_13675,N_12971);
and UO_303 (O_303,N_14397,N_12406);
xor UO_304 (O_304,N_12039,N_12384);
or UO_305 (O_305,N_12389,N_13464);
nor UO_306 (O_306,N_12735,N_12217);
xnor UO_307 (O_307,N_13558,N_14360);
and UO_308 (O_308,N_12854,N_14065);
nor UO_309 (O_309,N_13891,N_13271);
xor UO_310 (O_310,N_13823,N_12913);
or UO_311 (O_311,N_13697,N_14521);
and UO_312 (O_312,N_12231,N_12262);
or UO_313 (O_313,N_12802,N_13424);
nand UO_314 (O_314,N_12118,N_14905);
and UO_315 (O_315,N_14109,N_12138);
xnor UO_316 (O_316,N_12958,N_14975);
and UO_317 (O_317,N_13035,N_13405);
or UO_318 (O_318,N_13846,N_13631);
and UO_319 (O_319,N_13553,N_14765);
and UO_320 (O_320,N_13601,N_14417);
or UO_321 (O_321,N_14325,N_12137);
or UO_322 (O_322,N_12845,N_13983);
xor UO_323 (O_323,N_13705,N_12136);
nor UO_324 (O_324,N_12044,N_12606);
and UO_325 (O_325,N_13883,N_12094);
or UO_326 (O_326,N_14829,N_13998);
or UO_327 (O_327,N_14316,N_14499);
nand UO_328 (O_328,N_12451,N_14971);
and UO_329 (O_329,N_12446,N_13592);
nand UO_330 (O_330,N_13585,N_13010);
nor UO_331 (O_331,N_12788,N_13024);
nor UO_332 (O_332,N_12912,N_14426);
and UO_333 (O_333,N_13446,N_14392);
xor UO_334 (O_334,N_14508,N_12923);
nand UO_335 (O_335,N_13756,N_13342);
or UO_336 (O_336,N_14845,N_12302);
nand UO_337 (O_337,N_13094,N_13571);
or UO_338 (O_338,N_14284,N_12615);
and UO_339 (O_339,N_12476,N_13655);
nor UO_340 (O_340,N_13231,N_13219);
and UO_341 (O_341,N_13459,N_14333);
and UO_342 (O_342,N_14968,N_14672);
and UO_343 (O_343,N_13536,N_12811);
or UO_344 (O_344,N_12651,N_13830);
and UO_345 (O_345,N_14328,N_14620);
or UO_346 (O_346,N_14872,N_13810);
and UO_347 (O_347,N_12871,N_13520);
xor UO_348 (O_348,N_12324,N_12351);
xor UO_349 (O_349,N_12429,N_14746);
nand UO_350 (O_350,N_13837,N_14754);
nand UO_351 (O_351,N_13013,N_13586);
and UO_352 (O_352,N_14398,N_12949);
nand UO_353 (O_353,N_13379,N_13646);
xnor UO_354 (O_354,N_12487,N_13591);
nor UO_355 (O_355,N_14369,N_12768);
or UO_356 (O_356,N_12167,N_12003);
nor UO_357 (O_357,N_14862,N_13677);
nor UO_358 (O_358,N_13803,N_12891);
and UO_359 (O_359,N_14793,N_14930);
and UO_360 (O_360,N_14926,N_12266);
nor UO_361 (O_361,N_12413,N_12225);
nand UO_362 (O_362,N_14093,N_14656);
nor UO_363 (O_363,N_14244,N_12470);
nand UO_364 (O_364,N_14472,N_14421);
nor UO_365 (O_365,N_12228,N_13860);
xor UO_366 (O_366,N_12208,N_13660);
and UO_367 (O_367,N_12649,N_13992);
xor UO_368 (O_368,N_14395,N_14120);
and UO_369 (O_369,N_14943,N_12297);
xor UO_370 (O_370,N_14148,N_13545);
or UO_371 (O_371,N_14129,N_12678);
nor UO_372 (O_372,N_14680,N_14557);
nand UO_373 (O_373,N_14097,N_14193);
nor UO_374 (O_374,N_13664,N_12091);
and UO_375 (O_375,N_13657,N_13742);
nor UO_376 (O_376,N_12388,N_12804);
nor UO_377 (O_377,N_12684,N_12145);
or UO_378 (O_378,N_13957,N_13089);
xnor UO_379 (O_379,N_14094,N_14590);
and UO_380 (O_380,N_12611,N_13495);
nor UO_381 (O_381,N_13104,N_12518);
xor UO_382 (O_382,N_14159,N_14222);
and UO_383 (O_383,N_14438,N_12875);
nor UO_384 (O_384,N_13313,N_12079);
or UO_385 (O_385,N_12791,N_14152);
nor UO_386 (O_386,N_13822,N_12590);
and UO_387 (O_387,N_13952,N_12069);
or UO_388 (O_388,N_12874,N_14509);
nand UO_389 (O_389,N_13514,N_12594);
nor UO_390 (O_390,N_14444,N_12319);
nand UO_391 (O_391,N_14855,N_13376);
nand UO_392 (O_392,N_12078,N_14902);
nor UO_393 (O_393,N_14238,N_14301);
nand UO_394 (O_394,N_12585,N_14588);
nand UO_395 (O_395,N_14343,N_12174);
xor UO_396 (O_396,N_14019,N_13159);
nor UO_397 (O_397,N_14642,N_12475);
xor UO_398 (O_398,N_14796,N_12340);
nor UO_399 (O_399,N_12479,N_14762);
and UO_400 (O_400,N_13297,N_13894);
nand UO_401 (O_401,N_13350,N_13059);
or UO_402 (O_402,N_14038,N_12789);
xnor UO_403 (O_403,N_13946,N_13960);
nor UO_404 (O_404,N_12710,N_13015);
xor UO_405 (O_405,N_13566,N_14527);
xnor UO_406 (O_406,N_13948,N_12113);
or UO_407 (O_407,N_12563,N_13401);
xor UO_408 (O_408,N_14272,N_14377);
and UO_409 (O_409,N_13373,N_14147);
or UO_410 (O_410,N_14653,N_13302);
nor UO_411 (O_411,N_12357,N_13873);
nor UO_412 (O_412,N_13133,N_13997);
or UO_413 (O_413,N_14675,N_14571);
or UO_414 (O_414,N_12657,N_13557);
or UO_415 (O_415,N_12356,N_14168);
and UO_416 (O_416,N_12897,N_13733);
or UO_417 (O_417,N_13574,N_12182);
nand UO_418 (O_418,N_12350,N_12284);
and UO_419 (O_419,N_12630,N_14432);
or UO_420 (O_420,N_13889,N_14655);
xor UO_421 (O_421,N_13616,N_13442);
and UO_422 (O_422,N_14057,N_12668);
nand UO_423 (O_423,N_14142,N_14047);
nor UO_424 (O_424,N_12970,N_14587);
or UO_425 (O_425,N_12127,N_13872);
nor UO_426 (O_426,N_14637,N_14814);
nor UO_427 (O_427,N_14404,N_12565);
nand UO_428 (O_428,N_13503,N_14942);
and UO_429 (O_429,N_14064,N_12742);
nor UO_430 (O_430,N_14135,N_12561);
or UO_431 (O_431,N_12612,N_12120);
or UO_432 (O_432,N_13204,N_12866);
nand UO_433 (O_433,N_13050,N_12043);
nor UO_434 (O_434,N_12507,N_13650);
or UO_435 (O_435,N_13524,N_13703);
nand UO_436 (O_436,N_12835,N_12283);
and UO_437 (O_437,N_12150,N_14918);
or UO_438 (O_438,N_13338,N_13273);
nand UO_439 (O_439,N_12362,N_13973);
xnor UO_440 (O_440,N_12054,N_13864);
or UO_441 (O_441,N_14589,N_14679);
nor UO_442 (O_442,N_12074,N_12445);
nor UO_443 (O_443,N_12492,N_14758);
xnor UO_444 (O_444,N_13125,N_13393);
or UO_445 (O_445,N_14743,N_12525);
or UO_446 (O_446,N_13955,N_12782);
xnor UO_447 (O_447,N_13169,N_14711);
nor UO_448 (O_448,N_14449,N_13102);
and UO_449 (O_449,N_14663,N_14884);
xnor UO_450 (O_450,N_12226,N_13859);
xnor UO_451 (O_451,N_13600,N_12510);
and UO_452 (O_452,N_13079,N_13950);
or UO_453 (O_453,N_13333,N_14989);
xor UO_454 (O_454,N_14950,N_12192);
nand UO_455 (O_455,N_14505,N_14648);
or UO_456 (O_456,N_13718,N_14837);
or UO_457 (O_457,N_14935,N_13316);
or UO_458 (O_458,N_12898,N_14475);
nand UO_459 (O_459,N_14225,N_14658);
nor UO_460 (O_460,N_14113,N_12125);
nand UO_461 (O_461,N_14880,N_12925);
and UO_462 (O_462,N_13044,N_14128);
nand UO_463 (O_463,N_13915,N_13106);
or UO_464 (O_464,N_13406,N_14705);
xnor UO_465 (O_465,N_12173,N_12140);
nand UO_466 (O_466,N_14789,N_12665);
and UO_467 (O_467,N_13738,N_14842);
xnor UO_468 (O_468,N_12890,N_13858);
xnor UO_469 (O_469,N_13760,N_13981);
and UO_470 (O_470,N_14896,N_14098);
xor UO_471 (O_471,N_13595,N_14209);
and UO_472 (O_472,N_13190,N_14337);
and UO_473 (O_473,N_13879,N_12233);
xnor UO_474 (O_474,N_13630,N_12821);
xor UO_475 (O_475,N_13188,N_13638);
nand UO_476 (O_476,N_14544,N_14480);
and UO_477 (O_477,N_13940,N_13931);
xor UO_478 (O_478,N_12001,N_13232);
or UO_479 (O_479,N_12819,N_12269);
nand UO_480 (O_480,N_12251,N_14843);
nor UO_481 (O_481,N_14912,N_13730);
nor UO_482 (O_482,N_14240,N_13776);
nand UO_483 (O_483,N_14056,N_12062);
nor UO_484 (O_484,N_13988,N_12050);
xnor UO_485 (O_485,N_13420,N_12489);
or UO_486 (O_486,N_13975,N_12452);
or UO_487 (O_487,N_12454,N_14778);
xor UO_488 (O_488,N_12279,N_12230);
or UO_489 (O_489,N_14983,N_14114);
and UO_490 (O_490,N_14524,N_12763);
xnor UO_491 (O_491,N_13961,N_14831);
xnor UO_492 (O_492,N_14704,N_14806);
nand UO_493 (O_493,N_13789,N_12930);
nand UO_494 (O_494,N_14771,N_14476);
nand UO_495 (O_495,N_13177,N_14374);
xor UO_496 (O_496,N_13051,N_14085);
and UO_497 (O_497,N_12341,N_13419);
or UO_498 (O_498,N_12911,N_13989);
nand UO_499 (O_499,N_14288,N_14695);
nor UO_500 (O_500,N_14703,N_14502);
or UO_501 (O_501,N_12117,N_14934);
nand UO_502 (O_502,N_14206,N_12133);
nand UO_503 (O_503,N_12213,N_12730);
or UO_504 (O_504,N_12016,N_14353);
and UO_505 (O_505,N_13494,N_13234);
nor UO_506 (O_506,N_14305,N_12688);
xnor UO_507 (O_507,N_12041,N_14747);
nand UO_508 (O_508,N_13395,N_14213);
nand UO_509 (O_509,N_14263,N_14308);
and UO_510 (O_510,N_14781,N_14635);
nand UO_511 (O_511,N_13624,N_14956);
nand UO_512 (O_512,N_14259,N_12696);
or UO_513 (O_513,N_13587,N_13603);
or UO_514 (O_514,N_14274,N_14616);
nand UO_515 (O_515,N_13588,N_14634);
nand UO_516 (O_516,N_12899,N_13118);
nand UO_517 (O_517,N_12652,N_12191);
xor UO_518 (O_518,N_14423,N_12511);
nand UO_519 (O_519,N_13529,N_14241);
or UO_520 (O_520,N_14341,N_14539);
nand UO_521 (O_521,N_13428,N_12008);
or UO_522 (O_522,N_14849,N_13135);
xnor UO_523 (O_523,N_14331,N_12773);
xor UO_524 (O_524,N_13386,N_14867);
nand UO_525 (O_525,N_12830,N_14181);
nor UO_526 (O_526,N_14349,N_14858);
and UO_527 (O_527,N_13091,N_12190);
xor UO_528 (O_528,N_12942,N_12529);
xor UO_529 (O_529,N_12643,N_12149);
nand UO_530 (O_530,N_14145,N_13016);
nor UO_531 (O_531,N_14605,N_12928);
or UO_532 (O_532,N_12088,N_12865);
nand UO_533 (O_533,N_13439,N_12670);
nand UO_534 (O_534,N_13400,N_12620);
xor UO_535 (O_535,N_14960,N_14730);
xor UO_536 (O_536,N_13815,N_13341);
and UO_537 (O_537,N_13131,N_12820);
or UO_538 (O_538,N_13214,N_12682);
and UO_539 (O_539,N_14454,N_12316);
and UO_540 (O_540,N_12267,N_12159);
and UO_541 (O_541,N_12801,N_12392);
or UO_542 (O_542,N_12627,N_14340);
nor UO_543 (O_543,N_14510,N_13809);
nor UO_544 (O_544,N_14370,N_12873);
and UO_545 (O_545,N_14086,N_12607);
or UO_546 (O_546,N_13380,N_14358);
or UO_547 (O_547,N_12979,N_12409);
nor UO_548 (O_548,N_13224,N_13530);
or UO_549 (O_549,N_12944,N_12505);
and UO_550 (O_550,N_12089,N_12642);
and UO_551 (O_551,N_13414,N_12290);
nor UO_552 (O_552,N_12704,N_12439);
nor UO_553 (O_553,N_12568,N_13715);
and UO_554 (O_554,N_14787,N_13667);
and UO_555 (O_555,N_13471,N_12246);
or UO_556 (O_556,N_14863,N_14729);
nor UO_557 (O_557,N_12646,N_13644);
or UO_558 (O_558,N_13200,N_14803);
nor UO_559 (O_559,N_12543,N_12817);
nor UO_560 (O_560,N_12697,N_13391);
nor UO_561 (O_561,N_12352,N_12706);
nor UO_562 (O_562,N_13599,N_12520);
nor UO_563 (O_563,N_12771,N_14722);
or UO_564 (O_564,N_12151,N_12760);
and UO_565 (O_565,N_13244,N_13739);
nand UO_566 (O_566,N_12883,N_14083);
or UO_567 (O_567,N_14916,N_13618);
nor UO_568 (O_568,N_14585,N_14175);
or UO_569 (O_569,N_14764,N_14070);
nor UO_570 (O_570,N_12715,N_12963);
xor UO_571 (O_571,N_14997,N_14061);
nor UO_572 (O_572,N_13303,N_13196);
and UO_573 (O_573,N_12329,N_12674);
or UO_574 (O_574,N_14736,N_13201);
or UO_575 (O_575,N_14995,N_13290);
nand UO_576 (O_576,N_12399,N_14496);
and UO_577 (O_577,N_14111,N_12592);
and UO_578 (O_578,N_12252,N_13750);
nand UO_579 (O_579,N_14931,N_14548);
xnor UO_580 (O_580,N_14785,N_13688);
nand UO_581 (O_581,N_14799,N_12609);
nor UO_582 (O_582,N_12569,N_12278);
and UO_583 (O_583,N_13832,N_14784);
xnor UO_584 (O_584,N_14761,N_12163);
nand UO_585 (O_585,N_13935,N_12795);
or UO_586 (O_586,N_14021,N_12253);
xnor UO_587 (O_587,N_14173,N_12376);
and UO_588 (O_588,N_13076,N_12556);
xnor UO_589 (O_589,N_13576,N_13017);
or UO_590 (O_590,N_12035,N_14321);
xnor UO_591 (O_591,N_12002,N_14144);
and UO_592 (O_592,N_14277,N_13769);
and UO_593 (O_593,N_14289,N_12685);
nand UO_594 (O_594,N_13203,N_13019);
and UO_595 (O_595,N_14646,N_14877);
and UO_596 (O_596,N_14095,N_13572);
nor UO_597 (O_597,N_13757,N_12548);
and UO_598 (O_598,N_14376,N_14207);
xnor UO_599 (O_599,N_14344,N_12482);
nand UO_600 (O_600,N_12282,N_13778);
and UO_601 (O_601,N_12645,N_12663);
or UO_602 (O_602,N_12433,N_14992);
xor UO_603 (O_603,N_14309,N_14319);
xor UO_604 (O_604,N_14882,N_14629);
and UO_605 (O_605,N_12378,N_14091);
or UO_606 (O_606,N_13254,N_12751);
nor UO_607 (O_607,N_13732,N_12541);
xor UO_608 (O_608,N_14155,N_13075);
xor UO_609 (O_609,N_12954,N_13144);
nand UO_610 (O_610,N_14928,N_12224);
or UO_611 (O_611,N_14078,N_14774);
nor UO_612 (O_612,N_13905,N_13817);
xnor UO_613 (O_613,N_14252,N_12420);
nand UO_614 (O_614,N_13065,N_12220);
xnor UO_615 (O_615,N_13417,N_12690);
xnor UO_616 (O_616,N_14131,N_13477);
nor UO_617 (O_617,N_13687,N_13827);
nand UO_618 (O_618,N_12806,N_12205);
xor UO_619 (O_619,N_13596,N_12098);
or UO_620 (O_620,N_14455,N_14553);
xnor UO_621 (O_621,N_13578,N_14281);
and UO_622 (O_622,N_13671,N_14887);
xor UO_623 (O_623,N_12530,N_13223);
nand UO_624 (O_624,N_12818,N_14390);
nor UO_625 (O_625,N_12631,N_12754);
nor UO_626 (O_626,N_13639,N_14772);
nor UO_627 (O_627,N_14051,N_12860);
or UO_628 (O_628,N_14262,N_14324);
nor UO_629 (O_629,N_12235,N_13216);
and UO_630 (O_630,N_12308,N_13556);
nand UO_631 (O_631,N_12832,N_14379);
or UO_632 (O_632,N_13445,N_14371);
nand UO_633 (O_633,N_14231,N_13661);
xnor UO_634 (O_634,N_12153,N_13819);
and UO_635 (O_635,N_13005,N_14534);
or UO_636 (O_636,N_14462,N_13758);
nand UO_637 (O_637,N_14180,N_14382);
and UO_638 (O_638,N_12756,N_14090);
or UO_639 (O_639,N_14116,N_13685);
nor UO_640 (O_640,N_13623,N_12586);
and UO_641 (O_641,N_13936,N_13522);
nor UO_642 (O_642,N_14640,N_12048);
and UO_643 (O_643,N_12636,N_12109);
nor UO_644 (O_644,N_14101,N_14219);
and UO_645 (O_645,N_13043,N_13971);
or UO_646 (O_646,N_13063,N_14041);
and UO_647 (O_647,N_13740,N_13032);
nand UO_648 (O_648,N_13692,N_14538);
or UO_649 (O_649,N_12933,N_14345);
or UO_650 (O_650,N_12539,N_13317);
nor UO_651 (O_651,N_13358,N_13540);
or UO_652 (O_652,N_12122,N_14126);
nor UO_653 (O_653,N_12155,N_13403);
nand UO_654 (O_654,N_12291,N_12610);
nor UO_655 (O_655,N_13647,N_14967);
nand UO_656 (O_656,N_13331,N_13628);
or UO_657 (O_657,N_14335,N_12277);
xnor UO_658 (O_658,N_13180,N_12018);
nor UO_659 (O_659,N_13036,N_13654);
xor UO_660 (O_660,N_12071,N_13759);
nand UO_661 (O_661,N_14217,N_13155);
or UO_662 (O_662,N_14561,N_12776);
xor UO_663 (O_663,N_12051,N_14984);
xnor UO_664 (O_664,N_12761,N_12330);
xor UO_665 (O_665,N_12201,N_12850);
nor UO_666 (O_666,N_12488,N_14125);
and UO_667 (O_667,N_14182,N_14253);
nand UO_668 (O_668,N_14346,N_13597);
nand UO_669 (O_669,N_13901,N_14555);
nand UO_670 (O_670,N_14551,N_13721);
and UO_671 (O_671,N_14721,N_14133);
and UO_672 (O_672,N_14604,N_12349);
nand UO_673 (O_673,N_12877,N_13734);
xnor UO_674 (O_674,N_14200,N_14493);
or UO_675 (O_675,N_14338,N_12841);
nor UO_676 (O_676,N_14052,N_14661);
nand UO_677 (O_677,N_14256,N_12900);
or UO_678 (O_678,N_14383,N_14456);
or UO_679 (O_679,N_13727,N_13362);
or UO_680 (O_680,N_13550,N_12381);
xor UO_681 (O_681,N_13724,N_12535);
xor UO_682 (O_682,N_14532,N_12542);
nand UO_683 (O_683,N_14906,N_12260);
nand UO_684 (O_684,N_14622,N_14523);
xnor UO_685 (O_685,N_12203,N_12745);
nand UO_686 (O_686,N_13633,N_13452);
and UO_687 (O_687,N_14007,N_14267);
and UO_688 (O_688,N_13001,N_13725);
and UO_689 (O_689,N_13840,N_12387);
and UO_690 (O_690,N_14750,N_12836);
xnor UO_691 (O_691,N_14535,N_13897);
and UO_692 (O_692,N_12232,N_14560);
and UO_693 (O_693,N_14313,N_14776);
xor UO_694 (O_694,N_13611,N_13965);
nor UO_695 (O_695,N_13142,N_12658);
nand UO_696 (O_696,N_12815,N_14507);
nor UO_697 (O_697,N_13009,N_14895);
and UO_698 (O_698,N_13941,N_13381);
xor UO_699 (O_699,N_12503,N_14192);
or UO_700 (O_700,N_12345,N_13669);
and UO_701 (O_701,N_13071,N_13862);
or UO_702 (O_702,N_13141,N_12662);
and UO_703 (O_703,N_12466,N_14342);
nor UO_704 (O_704,N_12948,N_12011);
nor UO_705 (O_705,N_12692,N_13893);
and UO_706 (O_706,N_14873,N_14838);
nand UO_707 (O_707,N_12065,N_14565);
and UO_708 (O_708,N_13953,N_12886);
xnor UO_709 (O_709,N_14850,N_14808);
xor UO_710 (O_710,N_14638,N_14671);
or UO_711 (O_711,N_12397,N_14861);
or UO_712 (O_712,N_14491,N_13861);
nor UO_713 (O_713,N_14162,N_13895);
nand UO_714 (O_714,N_14540,N_13348);
nor UO_715 (O_715,N_14016,N_13128);
nor UO_716 (O_716,N_14251,N_12086);
and UO_717 (O_717,N_14214,N_13782);
xnor UO_718 (O_718,N_13165,N_13301);
nand UO_719 (O_719,N_12550,N_13226);
xnor UO_720 (O_720,N_12738,N_12410);
and UO_721 (O_721,N_12254,N_13570);
or UO_722 (O_722,N_12603,N_12264);
and UO_723 (O_723,N_14593,N_14879);
nor UO_724 (O_724,N_12824,N_13824);
or UO_725 (O_725,N_14204,N_12411);
xor UO_726 (O_726,N_13658,N_12061);
nor UO_727 (O_727,N_13121,N_12896);
or UO_728 (O_728,N_13475,N_13048);
and UO_729 (O_729,N_12783,N_12042);
and UO_730 (O_730,N_13086,N_12049);
nand UO_731 (O_731,N_13841,N_14973);
and UO_732 (O_732,N_12868,N_14218);
or UO_733 (O_733,N_12023,N_13472);
xor UO_734 (O_734,N_14283,N_12261);
nor UO_735 (O_735,N_12240,N_12477);
nor UO_736 (O_736,N_13818,N_13430);
nand UO_737 (O_737,N_13160,N_12075);
xor UO_738 (O_738,N_13397,N_12846);
xor UO_739 (O_739,N_14908,N_14506);
and UO_740 (O_740,N_12432,N_14405);
nor UO_741 (O_741,N_14583,N_12936);
and UO_742 (O_742,N_14673,N_12905);
or UO_743 (O_743,N_14366,N_12083);
nand UO_744 (O_744,N_14350,N_14751);
and UO_745 (O_745,N_14482,N_14949);
xnor UO_746 (O_746,N_12941,N_13004);
xnor UO_747 (O_747,N_13662,N_13917);
or UO_748 (O_748,N_12060,N_13218);
and UO_749 (O_749,N_13367,N_14603);
nor UO_750 (O_750,N_13300,N_12750);
and UO_751 (O_751,N_12210,N_12363);
xor UO_752 (O_752,N_13288,N_14452);
or UO_753 (O_753,N_14246,N_13728);
and UO_754 (O_754,N_12540,N_14511);
nor UO_755 (O_755,N_13067,N_13878);
nand UO_756 (O_756,N_14484,N_12152);
or UO_757 (O_757,N_12864,N_14517);
nor UO_758 (O_758,N_13704,N_13937);
nand UO_759 (O_759,N_13263,N_12595);
and UO_760 (O_760,N_12012,N_13994);
nor UO_761 (O_761,N_14255,N_14836);
nand UO_762 (O_762,N_13025,N_13394);
or UO_763 (O_763,N_12046,N_13722);
or UO_764 (O_764,N_13833,N_13682);
nand UO_765 (O_765,N_12858,N_13785);
and UO_766 (O_766,N_12402,N_12259);
xnor UO_767 (O_767,N_12935,N_12453);
nand UO_768 (O_768,N_12072,N_12132);
xor UO_769 (O_769,N_12577,N_12371);
or UO_770 (O_770,N_12305,N_13385);
and UO_771 (O_771,N_12714,N_12177);
and UO_772 (O_772,N_14818,N_14292);
xnor UO_773 (O_773,N_14430,N_13857);
and UO_774 (O_774,N_14718,N_12239);
or UO_775 (O_775,N_13798,N_12066);
xnor UO_776 (O_776,N_14477,N_13235);
nor UO_777 (O_777,N_12531,N_13613);
nor UO_778 (O_778,N_13140,N_13185);
xnor UO_779 (O_779,N_13132,N_13268);
or UO_780 (O_780,N_13709,N_13110);
nand UO_781 (O_781,N_12703,N_12985);
or UO_782 (O_782,N_13648,N_12694);
xnor UO_783 (O_783,N_13521,N_14470);
or UO_784 (O_784,N_14805,N_12527);
xor UO_785 (O_785,N_14221,N_12523);
nor UO_786 (O_786,N_13353,N_14999);
nor UO_787 (O_787,N_12172,N_13531);
or UO_788 (O_788,N_13046,N_14044);
nor UO_789 (O_789,N_12570,N_14801);
xnor UO_790 (O_790,N_12759,N_14777);
or UO_791 (O_791,N_12506,N_12952);
xor UO_792 (O_792,N_12770,N_14488);
nand UO_793 (O_793,N_13084,N_13849);
nand UO_794 (O_794,N_12792,N_14782);
and UO_795 (O_795,N_12366,N_12679);
and UO_796 (O_796,N_14364,N_14362);
xor UO_797 (O_797,N_12227,N_14649);
or UO_798 (O_798,N_13296,N_14894);
or UO_799 (O_799,N_14531,N_12434);
nor UO_800 (O_800,N_12600,N_12695);
xnor UO_801 (O_801,N_13212,N_12171);
nor UO_802 (O_802,N_12513,N_12880);
or UO_803 (O_803,N_13619,N_12943);
and UO_804 (O_804,N_13339,N_14811);
nand UO_805 (O_805,N_13062,N_12810);
xor UO_806 (O_806,N_13347,N_14812);
or UO_807 (O_807,N_12336,N_13518);
or UO_808 (O_808,N_14541,N_13885);
and UO_809 (O_809,N_12289,N_14963);
nor UO_810 (O_810,N_13176,N_14048);
or UO_811 (O_811,N_12148,N_13807);
nor UO_812 (O_812,N_13670,N_12028);
nand UO_813 (O_813,N_13396,N_12144);
xnor UO_814 (O_814,N_13828,N_12637);
nor UO_815 (O_815,N_14591,N_14400);
xnor UO_816 (O_816,N_13517,N_14089);
nor UO_817 (O_817,N_12255,N_12281);
and UO_818 (O_818,N_13305,N_12978);
nor UO_819 (O_819,N_13145,N_13336);
nor UO_820 (O_820,N_14323,N_13468);
nand UO_821 (O_821,N_12731,N_13839);
nand UO_822 (O_822,N_12183,N_14387);
nand UO_823 (O_823,N_12486,N_13136);
xnor UO_824 (O_824,N_12947,N_13330);
nand UO_825 (O_825,N_13454,N_14584);
xor UO_826 (O_826,N_13918,N_14186);
or UO_827 (O_827,N_13371,N_12572);
or UO_828 (O_828,N_12998,N_13040);
nand UO_829 (O_829,N_13516,N_14878);
xor UO_830 (O_830,N_12143,N_12474);
or UO_831 (O_831,N_12602,N_14361);
nand UO_832 (O_832,N_13845,N_13134);
and UO_833 (O_833,N_12644,N_13150);
nand UO_834 (O_834,N_12085,N_13741);
or UO_835 (O_835,N_13700,N_13236);
or UO_836 (O_836,N_14760,N_12249);
xnor UO_837 (O_837,N_13707,N_12906);
nor UO_838 (O_838,N_12909,N_14731);
and UO_839 (O_839,N_14258,N_14559);
nor UO_840 (O_840,N_12559,N_14228);
nand UO_841 (O_841,N_12104,N_14923);
nor UO_842 (O_842,N_12142,N_12187);
or UO_843 (O_843,N_12332,N_14964);
xnor UO_844 (O_844,N_14137,N_12593);
and UO_845 (O_845,N_13182,N_12621);
nor UO_846 (O_846,N_14830,N_13875);
nand UO_847 (O_847,N_12650,N_12536);
nand UO_848 (O_848,N_14356,N_13635);
nor UO_849 (O_849,N_13856,N_13966);
or UO_850 (O_850,N_13974,N_14683);
and UO_851 (O_851,N_12456,N_14434);
and UO_852 (O_852,N_14828,N_12787);
nor UO_853 (O_853,N_12407,N_12720);
or UO_854 (O_854,N_13483,N_12707);
xnor UO_855 (O_855,N_14651,N_12790);
nor UO_856 (O_856,N_12160,N_14779);
or UO_857 (O_857,N_14798,N_13746);
or UO_858 (O_858,N_12081,N_12158);
nand UO_859 (O_859,N_14118,N_13496);
nor UO_860 (O_860,N_12884,N_13755);
nor UO_861 (O_861,N_12712,N_12881);
nor UO_862 (O_862,N_14676,N_12916);
nand UO_863 (O_863,N_14264,N_14389);
xnor UO_864 (O_864,N_12223,N_12448);
or UO_865 (O_865,N_14619,N_14685);
or UO_866 (O_866,N_13409,N_12579);
and UO_867 (O_867,N_12716,N_13152);
xnor UO_868 (O_868,N_13198,N_12995);
and UO_869 (O_869,N_14261,N_13976);
nand UO_870 (O_870,N_12981,N_13904);
nor UO_871 (O_871,N_14428,N_12797);
nand UO_872 (O_872,N_14644,N_14427);
or UO_873 (O_873,N_14478,N_12524);
or UO_874 (O_874,N_13222,N_12166);
or UO_875 (O_875,N_12856,N_14852);
nor UO_876 (O_876,N_13716,N_12382);
xnor UO_877 (O_877,N_14691,N_13907);
nand UO_878 (O_878,N_14525,N_13866);
xor UO_879 (O_879,N_13786,N_12006);
xor UO_880 (O_880,N_14609,N_13509);
nor UO_881 (O_881,N_14045,N_14146);
or UO_882 (O_882,N_12206,N_12953);
xnor UO_883 (O_883,N_13022,N_13298);
and UO_884 (O_884,N_12491,N_12929);
nor UO_885 (O_885,N_14897,N_14040);
and UO_886 (O_886,N_13548,N_13408);
and UO_887 (O_887,N_13467,N_13525);
nor UO_888 (O_888,N_13489,N_13456);
or UO_889 (O_889,N_13314,N_12215);
nand UO_890 (O_890,N_12982,N_12990);
xnor UO_891 (O_891,N_14717,N_14632);
nor UO_892 (O_892,N_12258,N_13179);
and UO_893 (O_893,N_12216,N_13986);
nor UO_894 (O_894,N_14678,N_13078);
or UO_895 (O_895,N_14939,N_12825);
nor UO_896 (O_896,N_14608,N_14486);
and UO_897 (O_897,N_13237,N_14208);
nand UO_898 (O_898,N_14958,N_12309);
or UO_899 (O_899,N_13243,N_14378);
or UO_900 (O_900,N_13228,N_14102);
nor UO_901 (O_901,N_13539,N_14003);
xor UO_902 (O_902,N_12997,N_14727);
nor UO_903 (O_903,N_12022,N_12829);
or UO_904 (O_904,N_13625,N_14460);
xor UO_905 (O_905,N_14848,N_13276);
xor UO_906 (O_906,N_14031,N_14790);
nor UO_907 (O_907,N_14183,N_14414);
and UO_908 (O_908,N_14339,N_12778);
nor UO_909 (O_909,N_12481,N_12270);
and UO_910 (O_910,N_14597,N_14198);
or UO_911 (O_911,N_14453,N_13107);
nand UO_912 (O_912,N_13181,N_12047);
xor UO_913 (O_913,N_14058,N_14840);
or UO_914 (O_914,N_12927,N_12844);
nand UO_915 (O_915,N_14441,N_13463);
and UO_916 (O_916,N_13500,N_12076);
xor UO_917 (O_917,N_12450,N_13093);
xor UO_918 (O_918,N_12861,N_12126);
or UO_919 (O_919,N_12110,N_14205);
nand UO_920 (O_920,N_13077,N_14914);
and UO_921 (O_921,N_13183,N_12960);
nor UO_922 (O_922,N_12057,N_14682);
nand UO_923 (O_923,N_14202,N_12124);
nor UO_924 (O_924,N_13484,N_14297);
nand UO_925 (O_925,N_13057,N_13272);
or UO_926 (O_926,N_14459,N_14742);
or UO_927 (O_927,N_14909,N_14719);
xnor UO_928 (O_928,N_14024,N_14174);
nor UO_929 (O_929,N_13762,N_13552);
nor UO_930 (O_930,N_12904,N_12656);
or UO_931 (O_931,N_12521,N_12917);
nor UO_932 (O_932,N_14954,N_13735);
nor UO_933 (O_933,N_13352,N_14139);
or UO_934 (O_934,N_14768,N_14269);
xnor UO_935 (O_935,N_13916,N_12793);
nor UO_936 (O_936,N_12512,N_14841);
xor UO_937 (O_937,N_12483,N_13425);
xnor UO_938 (O_938,N_12676,N_12584);
nor UO_939 (O_939,N_12721,N_13372);
and UO_940 (O_940,N_13577,N_12635);
nand UO_941 (O_941,N_14245,N_14610);
and UO_942 (O_942,N_12769,N_13951);
and UO_943 (O_943,N_14461,N_12504);
nor UO_944 (O_944,N_14270,N_13816);
or UO_945 (O_945,N_14248,N_13607);
xor UO_946 (O_946,N_13947,N_14903);
and UO_947 (O_947,N_13163,N_13679);
xor UO_948 (O_948,N_13049,N_14550);
xnor UO_949 (O_949,N_12141,N_14810);
nor UO_950 (O_950,N_12101,N_12156);
or UO_951 (O_951,N_14227,N_12010);
xnor UO_952 (O_952,N_12498,N_13617);
nand UO_953 (O_953,N_12711,N_12538);
nand UO_954 (O_954,N_12762,N_14938);
xor UO_955 (O_955,N_12032,N_13294);
or UO_956 (O_956,N_12814,N_12641);
nand UO_957 (O_957,N_14465,N_14976);
or UO_958 (O_958,N_12675,N_13326);
or UO_959 (O_959,N_14630,N_13968);
nand UO_960 (O_960,N_13737,N_14602);
or UO_961 (O_961,N_13854,N_13621);
xnor UO_962 (O_962,N_13389,N_13066);
nand UO_963 (O_963,N_13034,N_13932);
and UO_964 (O_964,N_14119,N_14273);
nand UO_965 (O_965,N_14957,N_14823);
xnor UO_966 (O_966,N_14986,N_13351);
nor UO_967 (O_967,N_13312,N_12373);
nor UO_968 (O_968,N_13765,N_13977);
nand UO_969 (O_969,N_14372,N_14469);
or UO_970 (O_970,N_12024,N_13323);
nor UO_971 (O_971,N_13129,N_12080);
nor UO_972 (O_972,N_13573,N_12727);
or UO_973 (O_973,N_13533,N_14108);
and UO_974 (O_974,N_13210,N_14410);
xor UO_975 (O_975,N_14668,N_14490);
xor UO_976 (O_976,N_12195,N_14994);
nor UO_977 (O_977,N_14315,N_13555);
and UO_978 (O_978,N_12855,N_12732);
xor UO_979 (O_979,N_14025,N_13207);
or UO_980 (O_980,N_14249,N_14385);
or UO_981 (O_981,N_13708,N_14359);
xor UO_982 (O_982,N_14763,N_13972);
nor UO_983 (O_983,N_12361,N_12702);
nor UO_984 (O_984,N_13925,N_14300);
or UO_985 (O_985,N_13543,N_12664);
and UO_986 (O_986,N_12121,N_12557);
nand UO_987 (O_987,N_12040,N_12544);
xnor UO_988 (O_988,N_12597,N_13148);
xnor UO_989 (O_989,N_12582,N_13674);
xor UO_990 (O_990,N_13942,N_14592);
or UO_991 (O_991,N_14723,N_12634);
or UO_992 (O_992,N_14991,N_13794);
xor UO_993 (O_993,N_14792,N_14966);
or UO_994 (O_994,N_13787,N_14536);
and UO_995 (O_995,N_14888,N_13802);
nor UO_996 (O_996,N_14612,N_13795);
nand UO_997 (O_997,N_14699,N_13421);
nor UO_998 (O_998,N_13825,N_14437);
or UO_999 (O_999,N_12991,N_13097);
nor UO_1000 (O_1000,N_12516,N_14947);
or UO_1001 (O_1001,N_12234,N_14487);
or UO_1002 (O_1002,N_13980,N_12034);
and UO_1003 (O_1003,N_12501,N_13020);
nor UO_1004 (O_1004,N_13911,N_12321);
nand UO_1005 (O_1005,N_14334,N_14197);
or UO_1006 (O_1006,N_13526,N_12689);
nor UO_1007 (O_1007,N_14614,N_12957);
or UO_1008 (O_1008,N_14278,N_14210);
xnor UO_1009 (O_1009,N_13712,N_14996);
and UO_1010 (O_1010,N_14298,N_14780);
nor UO_1011 (O_1011,N_14357,N_13247);
nor UO_1012 (O_1012,N_14435,N_12519);
and UO_1013 (O_1013,N_14659,N_12624);
nor UO_1014 (O_1014,N_12365,N_12115);
xor UO_1015 (O_1015,N_14088,N_14856);
xor UO_1016 (O_1016,N_14235,N_14839);
and UO_1017 (O_1017,N_13640,N_12945);
xnor UO_1018 (O_1018,N_13130,N_13146);
or UO_1019 (O_1019,N_12838,N_13714);
or UO_1020 (O_1020,N_12554,N_13512);
and UO_1021 (O_1021,N_14280,N_14327);
and UO_1022 (O_1022,N_14164,N_12996);
nor UO_1023 (O_1023,N_14519,N_14910);
or UO_1024 (O_1024,N_13168,N_14883);
nand UO_1025 (O_1025,N_14724,N_13384);
or UO_1026 (O_1026,N_13602,N_12263);
xnor UO_1027 (O_1027,N_13820,N_12331);
or UO_1028 (O_1028,N_14783,N_12918);
nor UO_1029 (O_1029,N_12438,N_14617);
or UO_1030 (O_1030,N_13470,N_14564);
xnor UO_1031 (O_1031,N_14817,N_13643);
nand UO_1032 (O_1032,N_14073,N_14802);
xnor UO_1033 (O_1033,N_14130,N_13026);
or UO_1034 (O_1034,N_14203,N_13774);
or UO_1035 (O_1035,N_14418,N_14697);
xnor UO_1036 (O_1036,N_14545,N_14473);
xor UO_1037 (O_1037,N_13469,N_12423);
nor UO_1038 (O_1038,N_13388,N_13178);
nand UO_1039 (O_1039,N_14515,N_14595);
and UO_1040 (O_1040,N_14196,N_13291);
nand UO_1041 (O_1041,N_14577,N_13360);
nor UO_1042 (O_1042,N_13124,N_13641);
or UO_1043 (O_1043,N_14965,N_14600);
and UO_1044 (O_1044,N_12180,N_12975);
or UO_1045 (O_1045,N_14322,N_13108);
xor UO_1046 (O_1046,N_13900,N_13978);
nor UO_1047 (O_1047,N_14158,N_14846);
or UO_1048 (O_1048,N_12986,N_13109);
nand UO_1049 (O_1049,N_14232,N_13028);
nand UO_1050 (O_1050,N_12955,N_13969);
nand UO_1051 (O_1051,N_14355,N_13538);
and UO_1052 (O_1052,N_13493,N_13100);
xnor UO_1053 (O_1053,N_14285,N_14303);
nor UO_1054 (O_1054,N_12508,N_13327);
and UO_1055 (O_1055,N_12390,N_13030);
or UO_1056 (O_1056,N_13256,N_14921);
nor UO_1057 (O_1057,N_12588,N_13967);
or UO_1058 (O_1058,N_12218,N_14239);
nor UO_1059 (O_1059,N_13851,N_13088);
or UO_1060 (O_1060,N_14669,N_14503);
nor UO_1061 (O_1061,N_12449,N_12765);
nor UO_1062 (O_1062,N_14010,N_14816);
or UO_1063 (O_1063,N_13903,N_14074);
and UO_1064 (O_1064,N_13426,N_13887);
and UO_1065 (O_1065,N_14006,N_13038);
and UO_1066 (O_1066,N_13847,N_14485);
xnor UO_1067 (O_1067,N_12311,N_13559);
or UO_1068 (O_1068,N_13229,N_14725);
xor UO_1069 (O_1069,N_14694,N_13390);
nand UO_1070 (O_1070,N_13116,N_13000);
xor UO_1071 (O_1071,N_13766,N_13441);
xor UO_1072 (O_1072,N_12131,N_12833);
nand UO_1073 (O_1073,N_14050,N_13275);
and UO_1074 (O_1074,N_13612,N_13458);
or UO_1075 (O_1075,N_14211,N_13435);
nor UO_1076 (O_1076,N_14533,N_13392);
or UO_1077 (O_1077,N_13418,N_13366);
nand UO_1078 (O_1078,N_13826,N_12139);
and UO_1079 (O_1079,N_14893,N_12013);
nand UO_1080 (O_1080,N_14665,N_12903);
and UO_1081 (O_1081,N_14179,N_14310);
or UO_1082 (O_1082,N_13217,N_12293);
nor UO_1083 (O_1083,N_12162,N_13287);
nor UO_1084 (O_1084,N_13092,N_12729);
xnor UO_1085 (O_1085,N_12562,N_12157);
or UO_1086 (O_1086,N_13255,N_12514);
nand UO_1087 (O_1087,N_14924,N_13806);
nor UO_1088 (O_1088,N_14662,N_12093);
nor UO_1089 (O_1089,N_13153,N_12619);
nand UO_1090 (O_1090,N_13871,N_13652);
nor UO_1091 (O_1091,N_12497,N_14706);
or UO_1092 (O_1092,N_14504,N_12306);
xor UO_1093 (O_1093,N_13230,N_13775);
or UO_1094 (O_1094,N_12123,N_13663);
or UO_1095 (O_1095,N_12325,N_13575);
nor UO_1096 (O_1096,N_14710,N_14451);
xor UO_1097 (O_1097,N_12980,N_14734);
and UO_1098 (O_1098,N_14716,N_14528);
and UO_1099 (O_1099,N_12764,N_13683);
xnor UO_1100 (O_1100,N_14104,N_12683);
xor UO_1101 (O_1101,N_13876,N_14598);
nand UO_1102 (O_1102,N_14212,N_14140);
nand UO_1103 (O_1103,N_13834,N_14582);
or UO_1104 (O_1104,N_14885,N_14891);
and UO_1105 (O_1105,N_14399,N_14797);
nor UO_1106 (O_1106,N_13938,N_14623);
nor UO_1107 (O_1107,N_13729,N_13615);
xor UO_1108 (O_1108,N_13466,N_14530);
nor UO_1109 (O_1109,N_12549,N_13488);
nor UO_1110 (O_1110,N_14069,N_13751);
nor UO_1111 (O_1111,N_14952,N_12626);
and UO_1112 (O_1112,N_13413,N_14985);
or UO_1113 (O_1113,N_13045,N_13457);
or UO_1114 (O_1114,N_13197,N_13506);
and UO_1115 (O_1115,N_13480,N_13731);
xnor UO_1116 (O_1116,N_12828,N_13137);
and UO_1117 (O_1117,N_13609,N_12221);
nor UO_1118 (O_1118,N_12677,N_12037);
xnor UO_1119 (O_1119,N_13158,N_14132);
xor UO_1120 (O_1120,N_14687,N_12639);
nand UO_1121 (O_1121,N_13584,N_12073);
or UO_1122 (O_1122,N_14972,N_14243);
and UO_1123 (O_1123,N_13344,N_13706);
nor UO_1124 (O_1124,N_12827,N_12813);
nand UO_1125 (O_1125,N_13523,N_14868);
or UO_1126 (O_1126,N_13486,N_14526);
nand UO_1127 (O_1127,N_13193,N_12796);
nand UO_1128 (O_1128,N_12848,N_14296);
or UO_1129 (O_1129,N_14415,N_14275);
and UO_1130 (O_1130,N_12613,N_12552);
or UO_1131 (O_1131,N_12545,N_12879);
nor UO_1132 (O_1132,N_14122,N_12271);
nand UO_1133 (O_1133,N_12705,N_13250);
xor UO_1134 (O_1134,N_13187,N_14257);
nand UO_1135 (O_1135,N_13498,N_13321);
xor UO_1136 (O_1136,N_13634,N_14657);
or UO_1137 (O_1137,N_14494,N_14977);
nor UO_1138 (O_1138,N_14881,N_13449);
nor UO_1139 (O_1139,N_12596,N_13053);
nand UO_1140 (O_1140,N_13365,N_12181);
nand UO_1141 (O_1141,N_13289,N_14157);
and UO_1142 (O_1142,N_12852,N_14042);
xor UO_1143 (O_1143,N_14990,N_12128);
xnor UO_1144 (O_1144,N_13315,N_12849);
or UO_1145 (O_1145,N_13642,N_13422);
nand UO_1146 (O_1146,N_12581,N_12546);
nor UO_1147 (O_1147,N_12993,N_14650);
nand UO_1148 (O_1148,N_14907,N_14406);
or UO_1149 (O_1149,N_12380,N_12888);
nor UO_1150 (O_1150,N_14689,N_13473);
and UO_1151 (O_1151,N_14794,N_13880);
nor UO_1152 (O_1152,N_12304,N_14306);
or UO_1153 (O_1153,N_13242,N_13283);
nor UO_1154 (O_1154,N_12533,N_12014);
or UO_1155 (O_1155,N_14005,N_12315);
or UO_1156 (O_1156,N_13069,N_14474);
or UO_1157 (O_1157,N_12459,N_13863);
nor UO_1158 (O_1158,N_14720,N_12430);
and UO_1159 (O_1159,N_13274,N_12781);
and UO_1160 (O_1160,N_14898,N_12464);
nand UO_1161 (O_1161,N_14690,N_13410);
and UO_1162 (O_1162,N_12977,N_14865);
nand UO_1163 (O_1163,N_13812,N_14944);
and UO_1164 (O_1164,N_13954,N_14265);
xnor UO_1165 (O_1165,N_13502,N_13945);
and UO_1166 (O_1166,N_14481,N_14033);
nor UO_1167 (O_1167,N_12280,N_12984);
nand UO_1168 (O_1168,N_12031,N_12580);
xor UO_1169 (O_1169,N_14737,N_14529);
nand UO_1170 (O_1170,N_13713,N_13886);
and UO_1171 (O_1171,N_13416,N_14201);
nand UO_1172 (O_1172,N_12404,N_12517);
or UO_1173 (O_1173,N_14386,N_14692);
and UO_1174 (O_1174,N_13695,N_14501);
nor UO_1175 (O_1175,N_14876,N_13564);
nor UO_1176 (O_1176,N_14151,N_12547);
or UO_1177 (O_1177,N_14988,N_12555);
or UO_1178 (O_1178,N_13363,N_14562);
nand UO_1179 (O_1179,N_12425,N_14029);
and UO_1180 (O_1180,N_13112,N_13164);
nand UO_1181 (O_1181,N_13637,N_14307);
and UO_1182 (O_1182,N_12701,N_14708);
xor UO_1183 (O_1183,N_14373,N_13914);
nand UO_1184 (O_1184,N_12396,N_14433);
nor UO_1185 (O_1185,N_12198,N_12102);
and UO_1186 (O_1186,N_12370,N_13202);
or UO_1187 (O_1187,N_12934,N_13743);
nor UO_1188 (O_1188,N_14440,N_14287);
nor UO_1189 (O_1189,N_12767,N_14920);
and UO_1190 (O_1190,N_12207,N_14314);
xor UO_1191 (O_1191,N_13399,N_13364);
or UO_1192 (O_1192,N_13877,N_13620);
and UO_1193 (O_1193,N_14282,N_13060);
nand UO_1194 (O_1194,N_13382,N_13012);
nor UO_1195 (O_1195,N_14443,N_14701);
xnor UO_1196 (O_1196,N_14568,N_13867);
nor UO_1197 (O_1197,N_13014,N_14969);
nand UO_1198 (O_1198,N_13656,N_14516);
nand UO_1199 (O_1199,N_14260,N_12417);
and UO_1200 (O_1200,N_14652,N_12826);
nor UO_1201 (O_1201,N_14892,N_13797);
xor UO_1202 (O_1202,N_14134,N_14468);
nor UO_1203 (O_1203,N_14075,N_14851);
nand UO_1204 (O_1204,N_13811,N_14028);
or UO_1205 (O_1205,N_12614,N_14822);
or UO_1206 (O_1206,N_12812,N_12989);
or UO_1207 (O_1207,N_12298,N_12485);
or UO_1208 (O_1208,N_14247,N_12604);
or UO_1209 (O_1209,N_13248,N_13448);
xor UO_1210 (O_1210,N_14576,N_14681);
xnor UO_1211 (O_1211,N_12753,N_13113);
xnor UO_1212 (O_1212,N_12405,N_13836);
and UO_1213 (O_1213,N_12851,N_13377);
xor UO_1214 (O_1214,N_12377,N_13434);
nand UO_1215 (O_1215,N_13792,N_12431);
and UO_1216 (O_1216,N_12241,N_13359);
nor UO_1217 (O_1217,N_12248,N_13537);
xnor UO_1218 (O_1218,N_14000,N_12739);
xnor UO_1219 (O_1219,N_14945,N_12669);
and UO_1220 (O_1220,N_13225,N_13838);
xor UO_1221 (O_1221,N_14170,N_13322);
nand UO_1222 (O_1222,N_13191,N_14419);
and UO_1223 (O_1223,N_14012,N_12383);
nor UO_1224 (O_1224,N_13292,N_13329);
nor UO_1225 (O_1225,N_13888,N_13277);
and UO_1226 (O_1226,N_13398,N_14236);
or UO_1227 (O_1227,N_13698,N_12418);
and UO_1228 (O_1228,N_14913,N_12969);
xnor UO_1229 (O_1229,N_12053,N_12026);
or UO_1230 (O_1230,N_12161,N_12310);
nor UO_1231 (O_1231,N_12314,N_12987);
and UO_1232 (O_1232,N_12681,N_12408);
or UO_1233 (O_1233,N_14184,N_12800);
xor UO_1234 (O_1234,N_12576,N_12490);
or UO_1235 (O_1235,N_14586,N_14643);
and UO_1236 (O_1236,N_12872,N_14185);
and UO_1237 (O_1237,N_12902,N_14575);
xor UO_1238 (O_1238,N_12400,N_12243);
nor UO_1239 (O_1239,N_12772,N_14566);
nor UO_1240 (O_1240,N_12994,N_12005);
and UO_1241 (O_1241,N_13407,N_14076);
nor UO_1242 (O_1242,N_13958,N_14832);
nor UO_1243 (O_1243,N_12465,N_13138);
and UO_1244 (O_1244,N_12758,N_13246);
and UO_1245 (O_1245,N_13119,N_14161);
and UO_1246 (O_1246,N_14411,N_13790);
or UO_1247 (O_1247,N_14036,N_13387);
and UO_1248 (O_1248,N_12922,N_12551);
nand UO_1249 (O_1249,N_13306,N_12660);
xnor UO_1250 (O_1250,N_14813,N_14807);
or UO_1251 (O_1251,N_13482,N_13850);
xor UO_1252 (O_1252,N_13095,N_14268);
and UO_1253 (O_1253,N_12938,N_13368);
nor UO_1254 (O_1254,N_14757,N_13211);
nand UO_1255 (O_1255,N_14295,N_13340);
xnor UO_1256 (O_1256,N_12741,N_14556);
xnor UO_1257 (O_1257,N_14948,N_14979);
nor UO_1258 (O_1258,N_13808,N_14216);
nor UO_1259 (O_1259,N_14639,N_13777);
or UO_1260 (O_1260,N_12193,N_12391);
or UO_1261 (O_1261,N_12092,N_14567);
or UO_1262 (O_1262,N_14498,N_14978);
and UO_1263 (O_1263,N_12461,N_14436);
nand UO_1264 (O_1264,N_14420,N_13606);
or UO_1265 (O_1265,N_13580,N_13295);
xor UO_1266 (O_1266,N_14294,N_12322);
xor UO_1267 (O_1267,N_13239,N_14601);
nor UO_1268 (O_1268,N_13944,N_12713);
nand UO_1269 (O_1269,N_13711,N_14570);
xor UO_1270 (O_1270,N_12749,N_14049);
nor UO_1271 (O_1271,N_12328,N_12722);
nand UO_1272 (O_1272,N_14422,N_13632);
nand UO_1273 (O_1273,N_14749,N_12537);
or UO_1274 (O_1274,N_12666,N_12725);
or UO_1275 (O_1275,N_12633,N_12386);
or UO_1276 (O_1276,N_13890,N_14018);
nand UO_1277 (O_1277,N_12966,N_12840);
or UO_1278 (O_1278,N_14035,N_12834);
nand UO_1279 (O_1279,N_14199,N_14715);
xor UO_1280 (O_1280,N_13744,N_12004);
and UO_1281 (O_1281,N_12502,N_12709);
nand UO_1282 (O_1282,N_12348,N_14302);
and UO_1283 (O_1283,N_14915,N_14401);
and UO_1284 (O_1284,N_13039,N_14791);
or UO_1285 (O_1285,N_12256,N_13487);
and UO_1286 (O_1286,N_14143,N_12099);
or UO_1287 (O_1287,N_12859,N_14099);
and UO_1288 (O_1288,N_12135,N_12025);
xnor UO_1289 (O_1289,N_14149,N_14962);
nor UO_1290 (O_1290,N_13805,N_12965);
or UO_1291 (O_1291,N_14429,N_13912);
nand UO_1292 (O_1292,N_13011,N_13453);
nand UO_1293 (O_1293,N_12334,N_13653);
nand UO_1294 (O_1294,N_13554,N_14688);
nand UO_1295 (O_1295,N_12937,N_14674);
nor UO_1296 (O_1296,N_13278,N_13717);
nor UO_1297 (O_1297,N_14667,N_13696);
nand UO_1298 (O_1298,N_12574,N_13930);
and UO_1299 (O_1299,N_13649,N_14766);
xor UO_1300 (O_1300,N_13699,N_13686);
nor UO_1301 (O_1301,N_12209,N_14121);
nand UO_1302 (O_1302,N_13054,N_12532);
nand UO_1303 (O_1303,N_12638,N_13349);
nand UO_1304 (O_1304,N_13565,N_13547);
and UO_1305 (O_1305,N_12847,N_14060);
nand UO_1306 (O_1306,N_12059,N_14707);
nand UO_1307 (O_1307,N_14698,N_14819);
or UO_1308 (O_1308,N_12743,N_13209);
nand UO_1309 (O_1309,N_12920,N_13437);
or UO_1310 (O_1310,N_12100,N_14394);
and UO_1311 (O_1311,N_12007,N_13745);
nor UO_1312 (O_1312,N_12601,N_12196);
nor UO_1313 (O_1313,N_14442,N_14514);
or UO_1314 (O_1314,N_14866,N_13504);
nand UO_1315 (O_1315,N_13943,N_13149);
xor UO_1316 (O_1316,N_14835,N_12212);
and UO_1317 (O_1317,N_13884,N_13791);
or UO_1318 (O_1318,N_14847,N_14492);
and UO_1319 (O_1319,N_13189,N_13626);
nand UO_1320 (O_1320,N_13465,N_12286);
or UO_1321 (O_1321,N_14853,N_13415);
nor UO_1322 (O_1322,N_13491,N_12951);
nor UO_1323 (O_1323,N_14079,N_14666);
xnor UO_1324 (O_1324,N_12038,N_13270);
and UO_1325 (O_1325,N_13460,N_12068);
or UO_1326 (O_1326,N_12526,N_12393);
or UO_1327 (O_1327,N_14709,N_13037);
nor UO_1328 (O_1328,N_14513,N_13003);
or UO_1329 (O_1329,N_14276,N_14821);
xor UO_1330 (O_1330,N_13111,N_13752);
nand UO_1331 (O_1331,N_13896,N_12369);
nand UO_1332 (O_1332,N_12401,N_13702);
nor UO_1333 (O_1333,N_14864,N_13598);
and UO_1334 (O_1334,N_12723,N_14416);
and UO_1335 (O_1335,N_14859,N_14982);
and UO_1336 (O_1336,N_14188,N_14153);
nor UO_1337 (O_1337,N_12412,N_12926);
or UO_1338 (O_1338,N_12441,N_13999);
and UO_1339 (O_1339,N_12009,N_13923);
or UO_1340 (O_1340,N_14981,N_12755);
nand UO_1341 (O_1341,N_12794,N_12116);
xor UO_1342 (O_1342,N_13499,N_13909);
and UO_1343 (O_1343,N_12522,N_13910);
nor UO_1344 (O_1344,N_13582,N_14190);
xnor UO_1345 (O_1345,N_12831,N_12272);
xnor UO_1346 (O_1346,N_12534,N_12106);
or UO_1347 (O_1347,N_13920,N_14326);
nand UO_1348 (O_1348,N_13478,N_14015);
or UO_1349 (O_1349,N_14014,N_13241);
xnor UO_1350 (O_1350,N_13324,N_12799);
nand UO_1351 (O_1351,N_13589,N_13101);
xor UO_1352 (O_1352,N_12962,N_13590);
nand UO_1353 (O_1353,N_14363,N_13605);
xnor UO_1354 (O_1354,N_12659,N_14304);
nor UO_1355 (O_1355,N_13370,N_12229);
or UO_1356 (O_1356,N_12803,N_13882);
nand UO_1357 (O_1357,N_12185,N_13984);
nand UO_1358 (O_1358,N_14380,N_13771);
xor UO_1359 (O_1359,N_13427,N_13052);
nor UO_1360 (O_1360,N_12095,N_13799);
nand UO_1361 (O_1361,N_12919,N_13593);
nor UO_1362 (O_1362,N_12096,N_13881);
and UO_1363 (O_1363,N_14625,N_14017);
or UO_1364 (O_1364,N_13659,N_14483);
xor UO_1365 (O_1365,N_12892,N_14191);
nor UO_1366 (O_1366,N_13784,N_12103);
and UO_1367 (O_1367,N_14020,N_13710);
nand UO_1368 (O_1368,N_12752,N_13267);
or UO_1369 (O_1369,N_12339,N_12862);
and UO_1370 (O_1370,N_12959,N_12200);
nand UO_1371 (O_1371,N_13962,N_13157);
nor UO_1372 (O_1372,N_12189,N_13122);
and UO_1373 (O_1373,N_14071,N_14752);
nand UO_1374 (O_1374,N_12333,N_14100);
nor UO_1375 (O_1375,N_14755,N_12617);
and UO_1376 (O_1376,N_13251,N_12843);
nand UO_1377 (O_1377,N_12468,N_13265);
nand UO_1378 (O_1378,N_14815,N_13781);
and UO_1379 (O_1379,N_12077,N_13723);
nor UO_1380 (O_1380,N_14901,N_13869);
xor UO_1381 (O_1381,N_14317,N_13993);
or UO_1382 (O_1382,N_14739,N_14330);
nor UO_1383 (O_1383,N_14466,N_13404);
or UO_1384 (O_1384,N_13963,N_12300);
nand UO_1385 (O_1385,N_13939,N_13337);
nand UO_1386 (O_1386,N_13561,N_14447);
nand UO_1387 (O_1387,N_13170,N_12560);
xnor UO_1388 (O_1388,N_12343,N_12188);
nand UO_1389 (O_1389,N_13492,N_13842);
nor UO_1390 (O_1390,N_12130,N_13684);
nor UO_1391 (O_1391,N_14998,N_12055);
or UO_1392 (O_1392,N_12687,N_14039);
nand UO_1393 (O_1393,N_14062,N_13928);
xor UO_1394 (O_1394,N_14574,N_14107);
xnor UO_1395 (O_1395,N_14194,N_13933);
nor UO_1396 (O_1396,N_13985,N_13681);
xor UO_1397 (O_1397,N_12728,N_14936);
and UO_1398 (O_1398,N_14463,N_12748);
nand UO_1399 (O_1399,N_14626,N_14242);
nor UO_1400 (O_1400,N_12869,N_14431);
or UO_1401 (O_1401,N_12029,N_14645);
nand UO_1402 (O_1402,N_13105,N_14178);
nor UO_1403 (O_1403,N_14318,N_14127);
and UO_1404 (O_1404,N_12632,N_12780);
xor UO_1405 (O_1405,N_14290,N_14860);
or UO_1406 (O_1406,N_14266,N_13865);
or UO_1407 (O_1407,N_14439,N_12499);
nor UO_1408 (O_1408,N_14150,N_13151);
and UO_1409 (O_1409,N_14922,N_12326);
or UO_1410 (O_1410,N_14756,N_12176);
xor UO_1411 (O_1411,N_13844,N_14788);
and UO_1412 (O_1412,N_13481,N_14412);
and UO_1413 (O_1413,N_13369,N_12693);
xnor UO_1414 (O_1414,N_12950,N_14388);
nor UO_1415 (O_1415,N_13666,N_14542);
and UO_1416 (O_1416,N_12885,N_12589);
or UO_1417 (O_1417,N_14450,N_13259);
or UO_1418 (O_1418,N_13378,N_14820);
and UO_1419 (O_1419,N_12442,N_14552);
or UO_1420 (O_1420,N_12921,N_14769);
or UO_1421 (O_1421,N_13513,N_12354);
xnor UO_1422 (O_1422,N_14271,N_13325);
nor UO_1423 (O_1423,N_14110,N_13691);
and UO_1424 (O_1424,N_13374,N_14347);
nand UO_1425 (O_1425,N_12618,N_14220);
nor UO_1426 (O_1426,N_13450,N_14312);
xnor UO_1427 (O_1427,N_12398,N_14154);
xnor UO_1428 (O_1428,N_12222,N_14166);
xor UO_1429 (O_1429,N_14664,N_14953);
nor UO_1430 (O_1430,N_12114,N_12931);
or UO_1431 (O_1431,N_14579,N_14495);
nand UO_1432 (O_1432,N_14599,N_13764);
nor UO_1433 (O_1433,N_12766,N_12805);
and UO_1434 (O_1434,N_12616,N_13253);
nor UO_1435 (O_1435,N_14904,N_14004);
or UO_1436 (O_1436,N_13173,N_14933);
nor UO_1437 (O_1437,N_13929,N_14448);
nand UO_1438 (O_1438,N_12628,N_13568);
nor UO_1439 (O_1439,N_13345,N_12421);
or UO_1440 (O_1440,N_12988,N_14176);
xor UO_1441 (O_1441,N_12733,N_13171);
nand UO_1442 (O_1442,N_13987,N_13736);
and UO_1443 (O_1443,N_13676,N_14558);
nand UO_1444 (O_1444,N_13293,N_12020);
and UO_1445 (O_1445,N_13068,N_14332);
or UO_1446 (O_1446,N_12671,N_14844);
xnor UO_1447 (O_1447,N_14618,N_12932);
and UO_1448 (O_1448,N_14402,N_12500);
and UO_1449 (O_1449,N_13892,N_13852);
nor UO_1450 (O_1450,N_13006,N_13665);
nor UO_1451 (O_1451,N_12027,N_12807);
nand UO_1452 (O_1452,N_12395,N_12983);
nor UO_1453 (O_1453,N_13343,N_12317);
nor UO_1454 (O_1454,N_13334,N_14911);
or UO_1455 (O_1455,N_12655,N_14163);
xnor UO_1456 (O_1456,N_13908,N_14393);
xor UO_1457 (O_1457,N_12667,N_13436);
nand UO_1458 (O_1458,N_12734,N_13423);
and UO_1459 (O_1459,N_13753,N_13147);
xnor UO_1460 (O_1460,N_12394,N_13061);
nand UO_1461 (O_1461,N_12784,N_13919);
xnor UO_1462 (O_1462,N_14068,N_14713);
and UO_1463 (O_1463,N_12907,N_12338);
xnor UO_1464 (O_1464,N_12893,N_13485);
nand UO_1465 (O_1465,N_14424,N_13073);
nand UO_1466 (O_1466,N_13162,N_13356);
nand UO_1467 (O_1467,N_12186,N_12939);
or UO_1468 (O_1468,N_12245,N_14870);
xor UO_1469 (O_1469,N_12344,N_14647);
nor UO_1470 (O_1470,N_13754,N_12359);
nor UO_1471 (O_1471,N_13257,N_12956);
nand UO_1472 (O_1472,N_13636,N_14497);
or UO_1473 (O_1473,N_14053,N_13898);
nand UO_1474 (O_1474,N_14696,N_14744);
and UO_1475 (O_1475,N_14408,N_14384);
nor UO_1476 (O_1476,N_12786,N_14712);
and UO_1477 (O_1477,N_14354,N_14654);
nand UO_1478 (O_1478,N_14009,N_13361);
xnor UO_1479 (O_1479,N_14141,N_13087);
or UO_1480 (O_1480,N_12837,N_12294);
or UO_1481 (O_1481,N_13085,N_14229);
nand UO_1482 (O_1482,N_14641,N_14403);
xnor UO_1483 (O_1483,N_12285,N_14329);
and UO_1484 (O_1484,N_12967,N_14234);
nand UO_1485 (O_1485,N_12680,N_12575);
and UO_1486 (O_1486,N_13123,N_12107);
and UO_1487 (O_1487,N_12587,N_13310);
or UO_1488 (O_1488,N_13161,N_12496);
xnor UO_1489 (O_1489,N_12385,N_13510);
and UO_1490 (O_1490,N_14046,N_13042);
nand UO_1491 (O_1491,N_12494,N_14886);
nor UO_1492 (O_1492,N_14770,N_13080);
or UO_1493 (O_1493,N_14970,N_13544);
nor UO_1494 (O_1494,N_13072,N_13829);
nor UO_1495 (O_1495,N_12625,N_14169);
xor UO_1496 (O_1496,N_14728,N_13031);
or UO_1497 (O_1497,N_14834,N_12699);
nand UO_1498 (O_1498,N_13855,N_13008);
nand UO_1499 (O_1499,N_12515,N_12058);
nor UO_1500 (O_1500,N_12398,N_13976);
and UO_1501 (O_1501,N_14265,N_13727);
nor UO_1502 (O_1502,N_13583,N_13205);
or UO_1503 (O_1503,N_14352,N_14393);
nand UO_1504 (O_1504,N_12895,N_13449);
or UO_1505 (O_1505,N_13323,N_12352);
or UO_1506 (O_1506,N_13958,N_14829);
nor UO_1507 (O_1507,N_13662,N_14114);
xnor UO_1508 (O_1508,N_13655,N_12091);
nand UO_1509 (O_1509,N_13559,N_12166);
nand UO_1510 (O_1510,N_14830,N_13746);
or UO_1511 (O_1511,N_14755,N_13865);
or UO_1512 (O_1512,N_13936,N_14283);
and UO_1513 (O_1513,N_13166,N_12678);
and UO_1514 (O_1514,N_14025,N_14205);
or UO_1515 (O_1515,N_14504,N_12349);
and UO_1516 (O_1516,N_13016,N_12020);
nor UO_1517 (O_1517,N_14732,N_13063);
nand UO_1518 (O_1518,N_14558,N_12378);
xnor UO_1519 (O_1519,N_12812,N_12233);
and UO_1520 (O_1520,N_12527,N_12005);
or UO_1521 (O_1521,N_12595,N_14887);
and UO_1522 (O_1522,N_14614,N_14546);
nand UO_1523 (O_1523,N_14126,N_12609);
xor UO_1524 (O_1524,N_14499,N_13943);
xor UO_1525 (O_1525,N_14900,N_12666);
nand UO_1526 (O_1526,N_13221,N_12491);
and UO_1527 (O_1527,N_12544,N_12086);
xnor UO_1528 (O_1528,N_12183,N_13757);
nor UO_1529 (O_1529,N_12190,N_13647);
nor UO_1530 (O_1530,N_13851,N_12649);
nor UO_1531 (O_1531,N_14289,N_12336);
or UO_1532 (O_1532,N_14458,N_14806);
nand UO_1533 (O_1533,N_14032,N_13210);
nor UO_1534 (O_1534,N_14762,N_14132);
xor UO_1535 (O_1535,N_12015,N_13685);
nand UO_1536 (O_1536,N_14081,N_13079);
and UO_1537 (O_1537,N_14700,N_13023);
and UO_1538 (O_1538,N_13939,N_12384);
and UO_1539 (O_1539,N_13414,N_13588);
xnor UO_1540 (O_1540,N_14615,N_13967);
and UO_1541 (O_1541,N_13732,N_12470);
nand UO_1542 (O_1542,N_14323,N_12296);
nor UO_1543 (O_1543,N_13144,N_14914);
or UO_1544 (O_1544,N_14183,N_12264);
nor UO_1545 (O_1545,N_13433,N_14717);
xnor UO_1546 (O_1546,N_13295,N_14362);
xnor UO_1547 (O_1547,N_14049,N_14036);
xor UO_1548 (O_1548,N_13273,N_14300);
nor UO_1549 (O_1549,N_13063,N_13012);
or UO_1550 (O_1550,N_12252,N_14125);
nor UO_1551 (O_1551,N_13784,N_14333);
nand UO_1552 (O_1552,N_14672,N_13811);
xnor UO_1553 (O_1553,N_12620,N_13972);
xnor UO_1554 (O_1554,N_12509,N_12960);
nand UO_1555 (O_1555,N_13957,N_14118);
or UO_1556 (O_1556,N_13187,N_14634);
nor UO_1557 (O_1557,N_12840,N_14252);
nand UO_1558 (O_1558,N_14841,N_12046);
and UO_1559 (O_1559,N_14975,N_14383);
or UO_1560 (O_1560,N_13019,N_12117);
nor UO_1561 (O_1561,N_13940,N_13630);
nor UO_1562 (O_1562,N_12004,N_14287);
or UO_1563 (O_1563,N_13977,N_12858);
and UO_1564 (O_1564,N_14375,N_12797);
or UO_1565 (O_1565,N_14883,N_12071);
nand UO_1566 (O_1566,N_14243,N_13456);
nand UO_1567 (O_1567,N_13587,N_13145);
nor UO_1568 (O_1568,N_14934,N_12313);
nand UO_1569 (O_1569,N_14716,N_13845);
or UO_1570 (O_1570,N_13114,N_13647);
nor UO_1571 (O_1571,N_12749,N_14722);
and UO_1572 (O_1572,N_12041,N_12028);
nand UO_1573 (O_1573,N_14573,N_14523);
nor UO_1574 (O_1574,N_14963,N_12702);
or UO_1575 (O_1575,N_12084,N_13441);
nand UO_1576 (O_1576,N_13893,N_12375);
xnor UO_1577 (O_1577,N_13685,N_12171);
or UO_1578 (O_1578,N_14769,N_12156);
and UO_1579 (O_1579,N_14701,N_12402);
nor UO_1580 (O_1580,N_12255,N_12416);
xor UO_1581 (O_1581,N_12080,N_13454);
xor UO_1582 (O_1582,N_12425,N_14775);
or UO_1583 (O_1583,N_13491,N_14924);
and UO_1584 (O_1584,N_14796,N_13668);
and UO_1585 (O_1585,N_12909,N_14247);
nor UO_1586 (O_1586,N_13619,N_12981);
or UO_1587 (O_1587,N_14733,N_12897);
xor UO_1588 (O_1588,N_12988,N_13230);
and UO_1589 (O_1589,N_14108,N_12150);
or UO_1590 (O_1590,N_12227,N_14164);
nor UO_1591 (O_1591,N_12172,N_12427);
or UO_1592 (O_1592,N_14077,N_13004);
or UO_1593 (O_1593,N_12111,N_12083);
nand UO_1594 (O_1594,N_12601,N_14613);
nor UO_1595 (O_1595,N_12494,N_12351);
xor UO_1596 (O_1596,N_12629,N_14851);
or UO_1597 (O_1597,N_13036,N_12051);
or UO_1598 (O_1598,N_12444,N_13507);
nand UO_1599 (O_1599,N_12972,N_13301);
nor UO_1600 (O_1600,N_14635,N_13961);
and UO_1601 (O_1601,N_13742,N_14742);
nand UO_1602 (O_1602,N_13338,N_13193);
or UO_1603 (O_1603,N_12709,N_13809);
xnor UO_1604 (O_1604,N_14789,N_13984);
and UO_1605 (O_1605,N_12516,N_12236);
or UO_1606 (O_1606,N_14360,N_13805);
nand UO_1607 (O_1607,N_14256,N_14849);
or UO_1608 (O_1608,N_12571,N_12863);
and UO_1609 (O_1609,N_13768,N_14180);
xnor UO_1610 (O_1610,N_14468,N_14109);
nand UO_1611 (O_1611,N_13554,N_13857);
nand UO_1612 (O_1612,N_13029,N_13832);
or UO_1613 (O_1613,N_12178,N_14222);
xnor UO_1614 (O_1614,N_12650,N_13881);
or UO_1615 (O_1615,N_12472,N_13682);
and UO_1616 (O_1616,N_14954,N_13043);
and UO_1617 (O_1617,N_13673,N_13939);
and UO_1618 (O_1618,N_12336,N_13413);
xor UO_1619 (O_1619,N_12728,N_12631);
xnor UO_1620 (O_1620,N_12933,N_13610);
or UO_1621 (O_1621,N_13349,N_14676);
xnor UO_1622 (O_1622,N_14587,N_13868);
or UO_1623 (O_1623,N_12400,N_14166);
nand UO_1624 (O_1624,N_14685,N_14035);
nand UO_1625 (O_1625,N_12767,N_12231);
xnor UO_1626 (O_1626,N_13553,N_13762);
nor UO_1627 (O_1627,N_12352,N_13096);
or UO_1628 (O_1628,N_12074,N_12552);
xnor UO_1629 (O_1629,N_12023,N_14910);
or UO_1630 (O_1630,N_14872,N_12100);
or UO_1631 (O_1631,N_14902,N_12909);
nand UO_1632 (O_1632,N_13370,N_13979);
nor UO_1633 (O_1633,N_14458,N_14474);
and UO_1634 (O_1634,N_12933,N_12996);
nand UO_1635 (O_1635,N_12294,N_14798);
or UO_1636 (O_1636,N_14836,N_12193);
and UO_1637 (O_1637,N_12455,N_12639);
nand UO_1638 (O_1638,N_13758,N_12626);
or UO_1639 (O_1639,N_13394,N_13121);
nand UO_1640 (O_1640,N_14848,N_12429);
and UO_1641 (O_1641,N_12949,N_14046);
and UO_1642 (O_1642,N_13894,N_12809);
or UO_1643 (O_1643,N_13484,N_12278);
nor UO_1644 (O_1644,N_14838,N_13027);
nand UO_1645 (O_1645,N_12262,N_13207);
nor UO_1646 (O_1646,N_14887,N_12032);
nand UO_1647 (O_1647,N_12778,N_14061);
nand UO_1648 (O_1648,N_14307,N_13524);
or UO_1649 (O_1649,N_14461,N_14631);
nand UO_1650 (O_1650,N_12393,N_12959);
nor UO_1651 (O_1651,N_14421,N_12323);
nor UO_1652 (O_1652,N_12865,N_14287);
nand UO_1653 (O_1653,N_14177,N_13253);
and UO_1654 (O_1654,N_14934,N_13581);
and UO_1655 (O_1655,N_14460,N_13210);
nor UO_1656 (O_1656,N_13006,N_14462);
xnor UO_1657 (O_1657,N_14745,N_12455);
nor UO_1658 (O_1658,N_14348,N_12493);
nand UO_1659 (O_1659,N_13926,N_12185);
nor UO_1660 (O_1660,N_14984,N_12514);
xor UO_1661 (O_1661,N_12940,N_14492);
and UO_1662 (O_1662,N_12170,N_12671);
xnor UO_1663 (O_1663,N_14567,N_13832);
and UO_1664 (O_1664,N_14315,N_14289);
or UO_1665 (O_1665,N_13034,N_13129);
nor UO_1666 (O_1666,N_14094,N_14461);
nor UO_1667 (O_1667,N_12314,N_13924);
nor UO_1668 (O_1668,N_14459,N_12146);
nor UO_1669 (O_1669,N_13742,N_12962);
nor UO_1670 (O_1670,N_13397,N_12647);
nor UO_1671 (O_1671,N_12056,N_14391);
and UO_1672 (O_1672,N_12188,N_12287);
xor UO_1673 (O_1673,N_13679,N_14512);
nand UO_1674 (O_1674,N_14663,N_12121);
nor UO_1675 (O_1675,N_13070,N_12422);
nand UO_1676 (O_1676,N_14389,N_13677);
or UO_1677 (O_1677,N_13639,N_14650);
or UO_1678 (O_1678,N_14396,N_12256);
xnor UO_1679 (O_1679,N_12754,N_14534);
and UO_1680 (O_1680,N_14142,N_14922);
or UO_1681 (O_1681,N_12977,N_14424);
nor UO_1682 (O_1682,N_12201,N_12840);
or UO_1683 (O_1683,N_13065,N_13585);
nand UO_1684 (O_1684,N_12281,N_12090);
nor UO_1685 (O_1685,N_13085,N_13676);
and UO_1686 (O_1686,N_13808,N_13889);
or UO_1687 (O_1687,N_14972,N_14767);
nand UO_1688 (O_1688,N_14211,N_13017);
or UO_1689 (O_1689,N_13556,N_14082);
and UO_1690 (O_1690,N_13061,N_14641);
or UO_1691 (O_1691,N_13703,N_12883);
and UO_1692 (O_1692,N_14417,N_13251);
or UO_1693 (O_1693,N_13494,N_14356);
xor UO_1694 (O_1694,N_13607,N_13065);
or UO_1695 (O_1695,N_14882,N_13448);
nor UO_1696 (O_1696,N_13862,N_12490);
nand UO_1697 (O_1697,N_14426,N_12206);
nor UO_1698 (O_1698,N_13776,N_12292);
or UO_1699 (O_1699,N_14164,N_14833);
nor UO_1700 (O_1700,N_13072,N_14738);
xnor UO_1701 (O_1701,N_14091,N_14315);
and UO_1702 (O_1702,N_12745,N_14499);
nor UO_1703 (O_1703,N_13827,N_13357);
or UO_1704 (O_1704,N_14344,N_13131);
and UO_1705 (O_1705,N_14613,N_14022);
nand UO_1706 (O_1706,N_14168,N_14530);
nand UO_1707 (O_1707,N_12799,N_14779);
or UO_1708 (O_1708,N_12938,N_13050);
nand UO_1709 (O_1709,N_14188,N_14177);
nand UO_1710 (O_1710,N_14536,N_14847);
xor UO_1711 (O_1711,N_12468,N_14324);
nand UO_1712 (O_1712,N_13729,N_13442);
nand UO_1713 (O_1713,N_12387,N_14195);
xnor UO_1714 (O_1714,N_14761,N_12374);
nor UO_1715 (O_1715,N_13718,N_13181);
xor UO_1716 (O_1716,N_13409,N_13566);
and UO_1717 (O_1717,N_12180,N_12312);
nand UO_1718 (O_1718,N_13155,N_12874);
or UO_1719 (O_1719,N_14961,N_12437);
or UO_1720 (O_1720,N_12374,N_12157);
nand UO_1721 (O_1721,N_12856,N_14124);
and UO_1722 (O_1722,N_13750,N_13193);
nor UO_1723 (O_1723,N_13019,N_12692);
nor UO_1724 (O_1724,N_13672,N_12176);
nor UO_1725 (O_1725,N_14253,N_14806);
or UO_1726 (O_1726,N_13613,N_13967);
nand UO_1727 (O_1727,N_14835,N_14421);
nand UO_1728 (O_1728,N_13000,N_12303);
xnor UO_1729 (O_1729,N_13720,N_14007);
xor UO_1730 (O_1730,N_12561,N_12182);
and UO_1731 (O_1731,N_14064,N_12069);
and UO_1732 (O_1732,N_13160,N_14536);
nand UO_1733 (O_1733,N_14025,N_12781);
nor UO_1734 (O_1734,N_14382,N_14773);
nand UO_1735 (O_1735,N_14490,N_14465);
and UO_1736 (O_1736,N_14773,N_13078);
nand UO_1737 (O_1737,N_12251,N_13668);
nand UO_1738 (O_1738,N_14070,N_13306);
nor UO_1739 (O_1739,N_14527,N_12677);
nor UO_1740 (O_1740,N_12886,N_14251);
nand UO_1741 (O_1741,N_12075,N_13122);
or UO_1742 (O_1742,N_14109,N_12927);
or UO_1743 (O_1743,N_14809,N_13665);
nor UO_1744 (O_1744,N_13457,N_13349);
nor UO_1745 (O_1745,N_12633,N_14455);
and UO_1746 (O_1746,N_13756,N_14456);
nand UO_1747 (O_1747,N_13001,N_13172);
or UO_1748 (O_1748,N_14870,N_12096);
nand UO_1749 (O_1749,N_12683,N_12890);
or UO_1750 (O_1750,N_12992,N_14256);
xor UO_1751 (O_1751,N_14515,N_12840);
xnor UO_1752 (O_1752,N_13577,N_13824);
nand UO_1753 (O_1753,N_12148,N_12195);
nor UO_1754 (O_1754,N_12124,N_12050);
or UO_1755 (O_1755,N_14787,N_12101);
and UO_1756 (O_1756,N_12212,N_12979);
nor UO_1757 (O_1757,N_13089,N_12317);
or UO_1758 (O_1758,N_12234,N_14520);
or UO_1759 (O_1759,N_12656,N_13077);
nor UO_1760 (O_1760,N_13397,N_14123);
or UO_1761 (O_1761,N_14206,N_13899);
or UO_1762 (O_1762,N_12301,N_14431);
nor UO_1763 (O_1763,N_12704,N_13207);
and UO_1764 (O_1764,N_12078,N_13750);
or UO_1765 (O_1765,N_12019,N_14337);
nor UO_1766 (O_1766,N_14231,N_13377);
and UO_1767 (O_1767,N_13032,N_13888);
xnor UO_1768 (O_1768,N_13333,N_14300);
nor UO_1769 (O_1769,N_14416,N_13668);
or UO_1770 (O_1770,N_13377,N_12388);
and UO_1771 (O_1771,N_14008,N_13903);
xor UO_1772 (O_1772,N_13076,N_13758);
nand UO_1773 (O_1773,N_14519,N_12069);
or UO_1774 (O_1774,N_14846,N_14303);
nand UO_1775 (O_1775,N_14012,N_14461);
xnor UO_1776 (O_1776,N_14129,N_13322);
nand UO_1777 (O_1777,N_12914,N_13921);
nand UO_1778 (O_1778,N_12061,N_12711);
xor UO_1779 (O_1779,N_13408,N_12258);
nor UO_1780 (O_1780,N_14059,N_13328);
nor UO_1781 (O_1781,N_13464,N_12061);
or UO_1782 (O_1782,N_12361,N_14455);
xnor UO_1783 (O_1783,N_13571,N_13135);
or UO_1784 (O_1784,N_14979,N_12543);
xor UO_1785 (O_1785,N_12682,N_12938);
and UO_1786 (O_1786,N_14311,N_12080);
xor UO_1787 (O_1787,N_12065,N_12817);
nand UO_1788 (O_1788,N_13866,N_14178);
nor UO_1789 (O_1789,N_12270,N_12776);
or UO_1790 (O_1790,N_14248,N_14177);
or UO_1791 (O_1791,N_14349,N_12360);
and UO_1792 (O_1792,N_14742,N_14066);
and UO_1793 (O_1793,N_14316,N_14613);
and UO_1794 (O_1794,N_12204,N_14933);
and UO_1795 (O_1795,N_12647,N_12572);
or UO_1796 (O_1796,N_12534,N_14809);
nand UO_1797 (O_1797,N_13414,N_14455);
and UO_1798 (O_1798,N_13764,N_14372);
xor UO_1799 (O_1799,N_12508,N_12817);
nand UO_1800 (O_1800,N_12532,N_12457);
and UO_1801 (O_1801,N_13620,N_12134);
or UO_1802 (O_1802,N_12315,N_13647);
nand UO_1803 (O_1803,N_12269,N_12206);
nor UO_1804 (O_1804,N_13612,N_14089);
xor UO_1805 (O_1805,N_12378,N_13698);
or UO_1806 (O_1806,N_13092,N_13556);
nand UO_1807 (O_1807,N_14727,N_12829);
xnor UO_1808 (O_1808,N_14846,N_12012);
or UO_1809 (O_1809,N_14042,N_14172);
xnor UO_1810 (O_1810,N_12435,N_12615);
xor UO_1811 (O_1811,N_14280,N_13611);
and UO_1812 (O_1812,N_13313,N_14552);
nor UO_1813 (O_1813,N_14290,N_13556);
xor UO_1814 (O_1814,N_13902,N_13812);
nand UO_1815 (O_1815,N_14797,N_13098);
nor UO_1816 (O_1816,N_14888,N_13022);
xnor UO_1817 (O_1817,N_14758,N_14858);
xnor UO_1818 (O_1818,N_12204,N_14271);
nand UO_1819 (O_1819,N_13951,N_13318);
nand UO_1820 (O_1820,N_13906,N_13775);
xor UO_1821 (O_1821,N_14305,N_13497);
xor UO_1822 (O_1822,N_14971,N_14297);
nor UO_1823 (O_1823,N_14745,N_12433);
nor UO_1824 (O_1824,N_14816,N_14806);
and UO_1825 (O_1825,N_13225,N_12463);
and UO_1826 (O_1826,N_13555,N_12427);
nor UO_1827 (O_1827,N_12802,N_14674);
nor UO_1828 (O_1828,N_12413,N_13731);
nand UO_1829 (O_1829,N_12661,N_12731);
nand UO_1830 (O_1830,N_13489,N_12674);
or UO_1831 (O_1831,N_13908,N_13180);
nor UO_1832 (O_1832,N_14696,N_14807);
or UO_1833 (O_1833,N_12153,N_12844);
and UO_1834 (O_1834,N_14046,N_14854);
and UO_1835 (O_1835,N_12683,N_14129);
nand UO_1836 (O_1836,N_12287,N_13283);
nor UO_1837 (O_1837,N_14071,N_14502);
xnor UO_1838 (O_1838,N_12728,N_14385);
xor UO_1839 (O_1839,N_12605,N_13114);
or UO_1840 (O_1840,N_12585,N_14376);
and UO_1841 (O_1841,N_12626,N_12054);
nand UO_1842 (O_1842,N_14768,N_13335);
nor UO_1843 (O_1843,N_12438,N_13217);
nand UO_1844 (O_1844,N_13762,N_13136);
or UO_1845 (O_1845,N_13436,N_13031);
or UO_1846 (O_1846,N_13361,N_12056);
or UO_1847 (O_1847,N_12081,N_14816);
nand UO_1848 (O_1848,N_13623,N_12684);
xor UO_1849 (O_1849,N_13534,N_13906);
or UO_1850 (O_1850,N_14735,N_14518);
nand UO_1851 (O_1851,N_14506,N_14471);
nand UO_1852 (O_1852,N_13261,N_13822);
and UO_1853 (O_1853,N_13281,N_13347);
and UO_1854 (O_1854,N_13898,N_12047);
and UO_1855 (O_1855,N_13845,N_14275);
nand UO_1856 (O_1856,N_13698,N_14062);
or UO_1857 (O_1857,N_13795,N_14546);
or UO_1858 (O_1858,N_14642,N_14490);
xnor UO_1859 (O_1859,N_12848,N_14896);
or UO_1860 (O_1860,N_14761,N_14977);
nor UO_1861 (O_1861,N_12361,N_14568);
xnor UO_1862 (O_1862,N_14862,N_13365);
nor UO_1863 (O_1863,N_14669,N_13902);
xnor UO_1864 (O_1864,N_14176,N_13950);
nor UO_1865 (O_1865,N_14821,N_12018);
or UO_1866 (O_1866,N_13296,N_12122);
or UO_1867 (O_1867,N_14876,N_12313);
or UO_1868 (O_1868,N_12767,N_12105);
xnor UO_1869 (O_1869,N_13468,N_13415);
nor UO_1870 (O_1870,N_14179,N_14980);
or UO_1871 (O_1871,N_14359,N_14775);
or UO_1872 (O_1872,N_12326,N_13385);
nand UO_1873 (O_1873,N_12283,N_12188);
and UO_1874 (O_1874,N_14146,N_14053);
nor UO_1875 (O_1875,N_14526,N_12397);
nor UO_1876 (O_1876,N_13638,N_12155);
and UO_1877 (O_1877,N_12594,N_13352);
xor UO_1878 (O_1878,N_12492,N_14036);
and UO_1879 (O_1879,N_12368,N_12354);
nand UO_1880 (O_1880,N_12002,N_12645);
nor UO_1881 (O_1881,N_14593,N_12576);
nor UO_1882 (O_1882,N_14047,N_12011);
and UO_1883 (O_1883,N_14125,N_12764);
xnor UO_1884 (O_1884,N_12277,N_13475);
and UO_1885 (O_1885,N_13495,N_13011);
xnor UO_1886 (O_1886,N_14594,N_12994);
nor UO_1887 (O_1887,N_12818,N_12919);
xnor UO_1888 (O_1888,N_13752,N_14333);
or UO_1889 (O_1889,N_12528,N_14901);
nand UO_1890 (O_1890,N_13183,N_13156);
xor UO_1891 (O_1891,N_13092,N_12453);
nand UO_1892 (O_1892,N_12198,N_13278);
or UO_1893 (O_1893,N_12797,N_12995);
nand UO_1894 (O_1894,N_14855,N_12219);
xnor UO_1895 (O_1895,N_12343,N_12965);
nand UO_1896 (O_1896,N_12346,N_13520);
nor UO_1897 (O_1897,N_12231,N_12449);
nand UO_1898 (O_1898,N_13111,N_14187);
xnor UO_1899 (O_1899,N_13178,N_14640);
nand UO_1900 (O_1900,N_13791,N_13878);
nor UO_1901 (O_1901,N_13159,N_14362);
or UO_1902 (O_1902,N_12106,N_12970);
xor UO_1903 (O_1903,N_14764,N_12485);
or UO_1904 (O_1904,N_14449,N_14685);
or UO_1905 (O_1905,N_13164,N_13547);
or UO_1906 (O_1906,N_14426,N_12240);
and UO_1907 (O_1907,N_12528,N_12687);
or UO_1908 (O_1908,N_13614,N_12348);
and UO_1909 (O_1909,N_12524,N_13518);
or UO_1910 (O_1910,N_12359,N_12956);
nor UO_1911 (O_1911,N_13250,N_14190);
nand UO_1912 (O_1912,N_14915,N_12779);
nand UO_1913 (O_1913,N_12586,N_14780);
or UO_1914 (O_1914,N_13832,N_14245);
nor UO_1915 (O_1915,N_14528,N_12974);
nand UO_1916 (O_1916,N_12984,N_13186);
xor UO_1917 (O_1917,N_13413,N_12406);
or UO_1918 (O_1918,N_13658,N_14119);
or UO_1919 (O_1919,N_12447,N_12061);
nand UO_1920 (O_1920,N_14951,N_14788);
or UO_1921 (O_1921,N_12059,N_12889);
and UO_1922 (O_1922,N_14087,N_13907);
xor UO_1923 (O_1923,N_14938,N_13282);
nand UO_1924 (O_1924,N_12302,N_12481);
nor UO_1925 (O_1925,N_14480,N_12221);
xor UO_1926 (O_1926,N_14928,N_12099);
xor UO_1927 (O_1927,N_12581,N_14600);
nand UO_1928 (O_1928,N_13290,N_13940);
nand UO_1929 (O_1929,N_14573,N_12589);
and UO_1930 (O_1930,N_12771,N_13493);
nor UO_1931 (O_1931,N_12703,N_12169);
nor UO_1932 (O_1932,N_14318,N_12415);
nand UO_1933 (O_1933,N_14900,N_12950);
or UO_1934 (O_1934,N_12036,N_13653);
xnor UO_1935 (O_1935,N_14653,N_14644);
or UO_1936 (O_1936,N_14727,N_12387);
nor UO_1937 (O_1937,N_12001,N_14284);
or UO_1938 (O_1938,N_12590,N_13705);
nand UO_1939 (O_1939,N_14624,N_13373);
nand UO_1940 (O_1940,N_14123,N_13361);
or UO_1941 (O_1941,N_13037,N_14660);
nand UO_1942 (O_1942,N_13206,N_14019);
nand UO_1943 (O_1943,N_12529,N_12743);
or UO_1944 (O_1944,N_12147,N_14529);
and UO_1945 (O_1945,N_14351,N_14771);
and UO_1946 (O_1946,N_12343,N_12128);
or UO_1947 (O_1947,N_13587,N_13729);
or UO_1948 (O_1948,N_12790,N_14168);
nor UO_1949 (O_1949,N_12516,N_14812);
nand UO_1950 (O_1950,N_12642,N_13843);
nor UO_1951 (O_1951,N_14762,N_14923);
and UO_1952 (O_1952,N_13313,N_12884);
or UO_1953 (O_1953,N_13255,N_12464);
nor UO_1954 (O_1954,N_12783,N_13723);
xor UO_1955 (O_1955,N_13443,N_13904);
and UO_1956 (O_1956,N_14178,N_12378);
or UO_1957 (O_1957,N_12785,N_12537);
and UO_1958 (O_1958,N_13443,N_12784);
xor UO_1959 (O_1959,N_14936,N_12242);
or UO_1960 (O_1960,N_14724,N_14146);
xnor UO_1961 (O_1961,N_13631,N_12900);
nor UO_1962 (O_1962,N_13311,N_12904);
nand UO_1963 (O_1963,N_14793,N_13798);
xor UO_1964 (O_1964,N_13760,N_12909);
and UO_1965 (O_1965,N_14043,N_14509);
xnor UO_1966 (O_1966,N_13479,N_14683);
nor UO_1967 (O_1967,N_14661,N_12750);
nand UO_1968 (O_1968,N_12940,N_14258);
nor UO_1969 (O_1969,N_12937,N_14882);
and UO_1970 (O_1970,N_14854,N_14275);
xnor UO_1971 (O_1971,N_12218,N_12736);
and UO_1972 (O_1972,N_13379,N_14422);
nand UO_1973 (O_1973,N_13871,N_14459);
xnor UO_1974 (O_1974,N_12724,N_13977);
or UO_1975 (O_1975,N_12306,N_14080);
nor UO_1976 (O_1976,N_12469,N_14285);
xor UO_1977 (O_1977,N_13398,N_13323);
nor UO_1978 (O_1978,N_13924,N_14198);
and UO_1979 (O_1979,N_14061,N_13231);
nand UO_1980 (O_1980,N_14810,N_13555);
or UO_1981 (O_1981,N_13607,N_13019);
or UO_1982 (O_1982,N_12468,N_12169);
and UO_1983 (O_1983,N_13856,N_12751);
and UO_1984 (O_1984,N_14786,N_13645);
or UO_1985 (O_1985,N_12686,N_14793);
and UO_1986 (O_1986,N_13001,N_12332);
nor UO_1987 (O_1987,N_13135,N_14264);
and UO_1988 (O_1988,N_14402,N_14909);
or UO_1989 (O_1989,N_13628,N_12881);
and UO_1990 (O_1990,N_12294,N_12508);
xor UO_1991 (O_1991,N_14897,N_13242);
or UO_1992 (O_1992,N_13564,N_14130);
or UO_1993 (O_1993,N_12507,N_12387);
nor UO_1994 (O_1994,N_13271,N_12060);
and UO_1995 (O_1995,N_14707,N_12454);
or UO_1996 (O_1996,N_12300,N_14233);
xor UO_1997 (O_1997,N_14928,N_14559);
or UO_1998 (O_1998,N_12351,N_14010);
or UO_1999 (O_1999,N_13765,N_12097);
endmodule