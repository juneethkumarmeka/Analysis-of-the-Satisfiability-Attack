module basic_750_5000_1000_2_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2503,N_2504,N_2505,N_2506,N_2507,N_2509,N_2511,N_2513,N_2514,N_2515,N_2516,N_2517,N_2519,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2537,N_2538,N_2539,N_2540,N_2541,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2571,N_2573,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2585,N_2586,N_2587,N_2589,N_2590,N_2591,N_2592,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2631,N_2632,N_2633,N_2634,N_2635,N_2637,N_2638,N_2640,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2650,N_2652,N_2654,N_2655,N_2657,N_2659,N_2662,N_2663,N_2664,N_2665,N_2667,N_2668,N_2669,N_2671,N_2672,N_2673,N_2676,N_2680,N_2681,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2702,N_2703,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2713,N_2714,N_2716,N_2717,N_2718,N_2720,N_2721,N_2722,N_2725,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2736,N_2737,N_2738,N_2739,N_2741,N_2742,N_2743,N_2744,N_2746,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2758,N_2759,N_2760,N_2761,N_2764,N_2765,N_2766,N_2767,N_2768,N_2770,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2788,N_2790,N_2791,N_2792,N_2795,N_2797,N_2798,N_2799,N_2800,N_2804,N_2805,N_2806,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2816,N_2817,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2839,N_2840,N_2841,N_2842,N_2843,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2853,N_2855,N_2856,N_2857,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2912,N_2913,N_2914,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2923,N_2924,N_2925,N_2926,N_2927,N_2929,N_2930,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2952,N_2953,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2991,N_2992,N_2993,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3012,N_3014,N_3015,N_3016,N_3019,N_3021,N_3023,N_3025,N_3026,N_3027,N_3028,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3043,N_3044,N_3045,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3068,N_3071,N_3072,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3088,N_3089,N_3092,N_3094,N_3095,N_3096,N_3097,N_3100,N_3101,N_3102,N_3103,N_3104,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3175,N_3177,N_3178,N_3180,N_3181,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3191,N_3193,N_3194,N_3195,N_3198,N_3199,N_3200,N_3202,N_3203,N_3204,N_3205,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3247,N_3248,N_3249,N_3250,N_3251,N_3253,N_3254,N_3255,N_3256,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3288,N_3289,N_3290,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3299,N_3300,N_3301,N_3302,N_3308,N_3309,N_3310,N_3311,N_3312,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3330,N_3331,N_3332,N_3334,N_3335,N_3336,N_3337,N_3340,N_3341,N_3343,N_3346,N_3347,N_3348,N_3349,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3373,N_3374,N_3375,N_3376,N_3377,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3389,N_3391,N_3392,N_3393,N_3394,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3408,N_3409,N_3411,N_3412,N_3413,N_3416,N_3418,N_3419,N_3420,N_3421,N_3422,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3435,N_3436,N_3437,N_3439,N_3440,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3449,N_3450,N_3451,N_3452,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3484,N_3485,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3513,N_3515,N_3516,N_3517,N_3518,N_3519,N_3521,N_3522,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3538,N_3539,N_3540,N_3543,N_3544,N_3545,N_3547,N_3548,N_3549,N_3551,N_3552,N_3553,N_3554,N_3556,N_3557,N_3558,N_3559,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3569,N_3570,N_3571,N_3572,N_3573,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3600,N_3601,N_3604,N_3605,N_3606,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3616,N_3617,N_3618,N_3620,N_3621,N_3622,N_3624,N_3625,N_3627,N_3628,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3638,N_3639,N_3641,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3657,N_3658,N_3659,N_3661,N_3663,N_3664,N_3665,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3691,N_3693,N_3694,N_3695,N_3696,N_3699,N_3700,N_3701,N_3703,N_3704,N_3705,N_3707,N_3708,N_3709,N_3710,N_3711,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3728,N_3729,N_3730,N_3731,N_3735,N_3736,N_3738,N_3739,N_3740,N_3741,N_3742,N_3744,N_3745,N_3746,N_3747,N_3752,N_3753,N_3754,N_3756,N_3757,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3768,N_3769,N_3773,N_3774,N_3775,N_3776,N_3777,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3792,N_3793,N_3795,N_3796,N_3800,N_3801,N_3802,N_3803,N_3805,N_3810,N_3811,N_3812,N_3813,N_3814,N_3816,N_3817,N_3818,N_3819,N_3821,N_3822,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3841,N_3842,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3857,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3867,N_3869,N_3870,N_3871,N_3872,N_3874,N_3875,N_3877,N_3878,N_3879,N_3882,N_3883,N_3884,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3905,N_3906,N_3907,N_3909,N_3910,N_3911,N_3914,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3923,N_3924,N_3925,N_3926,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3954,N_3955,N_3957,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3976,N_3978,N_3979,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4007,N_4008,N_4009,N_4010,N_4011,N_4014,N_4015,N_4016,N_4017,N_4019,N_4020,N_4021,N_4022,N_4023,N_4025,N_4026,N_4027,N_4028,N_4029,N_4031,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4041,N_4042,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4054,N_4055,N_4056,N_4057,N_4062,N_4063,N_4064,N_4066,N_4069,N_4070,N_4071,N_4072,N_4074,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4083,N_4084,N_4086,N_4087,N_4088,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4122,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4131,N_4133,N_4134,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4147,N_4148,N_4152,N_4153,N_4154,N_4156,N_4157,N_4159,N_4161,N_4163,N_4164,N_4165,N_4166,N_4167,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4189,N_4192,N_4193,N_4194,N_4195,N_4196,N_4198,N_4200,N_4201,N_4204,N_4206,N_4207,N_4208,N_4210,N_4211,N_4213,N_4214,N_4216,N_4218,N_4219,N_4220,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4230,N_4232,N_4233,N_4234,N_4235,N_4236,N_4239,N_4240,N_4242,N_4243,N_4244,N_4245,N_4246,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4265,N_4266,N_4269,N_4270,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4279,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4302,N_4303,N_4304,N_4305,N_4306,N_4308,N_4309,N_4310,N_4311,N_4313,N_4314,N_4316,N_4318,N_4320,N_4321,N_4323,N_4324,N_4325,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4344,N_4345,N_4346,N_4348,N_4349,N_4351,N_4353,N_4354,N_4355,N_4356,N_4357,N_4359,N_4361,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4374,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4385,N_4386,N_4388,N_4389,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4398,N_4399,N_4400,N_4401,N_4403,N_4404,N_4405,N_4409,N_4410,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4442,N_4443,N_4444,N_4446,N_4448,N_4449,N_4450,N_4451,N_4452,N_4455,N_4456,N_4457,N_4458,N_4459,N_4461,N_4463,N_4464,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4483,N_4484,N_4486,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4519,N_4520,N_4522,N_4523,N_4524,N_4525,N_4526,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4540,N_4541,N_4543,N_4545,N_4546,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4555,N_4556,N_4558,N_4560,N_4561,N_4563,N_4564,N_4567,N_4569,N_4570,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4595,N_4596,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4605,N_4607,N_4608,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4629,N_4630,N_4631,N_4632,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4653,N_4654,N_4655,N_4659,N_4660,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4690,N_4691,N_4692,N_4694,N_4695,N_4696,N_4697,N_4699,N_4701,N_4703,N_4704,N_4705,N_4706,N_4707,N_4709,N_4710,N_4711,N_4714,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4734,N_4735,N_4736,N_4737,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4795,N_4796,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4807,N_4808,N_4809,N_4810,N_4812,N_4814,N_4817,N_4818,N_4819,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4829,N_4830,N_4831,N_4832,N_4833,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4843,N_4845,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4856,N_4859,N_4861,N_4862,N_4863,N_4865,N_4866,N_4868,N_4869,N_4871,N_4872,N_4873,N_4874,N_4876,N_4877,N_4878,N_4879,N_4880,N_4882,N_4883,N_4884,N_4886,N_4887,N_4888,N_4889,N_4890,N_4892,N_4894,N_4895,N_4896,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4923,N_4925,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4947,N_4948,N_4949,N_4950,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4973,N_4975,N_4976,N_4977,N_4978,N_4979,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4998,N_4999;
nor U0 (N_0,In_475,In_12);
nand U1 (N_1,In_338,In_744);
nor U2 (N_2,In_720,In_204);
and U3 (N_3,In_738,In_633);
or U4 (N_4,In_657,In_733);
and U5 (N_5,In_623,In_539);
or U6 (N_6,In_5,In_134);
nand U7 (N_7,In_280,In_464);
or U8 (N_8,In_448,In_365);
or U9 (N_9,In_414,In_700);
xnor U10 (N_10,In_678,In_291);
nand U11 (N_11,In_129,In_650);
nand U12 (N_12,In_692,In_159);
or U13 (N_13,In_431,In_117);
and U14 (N_14,In_15,In_339);
nand U15 (N_15,In_285,In_284);
xnor U16 (N_16,In_606,In_385);
nand U17 (N_17,In_273,In_451);
and U18 (N_18,In_77,In_256);
nor U19 (N_19,In_579,In_468);
or U20 (N_20,In_47,In_296);
xor U21 (N_21,In_557,In_637);
or U22 (N_22,In_82,In_547);
or U23 (N_23,In_416,In_505);
nand U24 (N_24,In_149,In_211);
and U25 (N_25,In_563,In_699);
nand U26 (N_26,In_721,In_271);
and U27 (N_27,In_402,In_119);
or U28 (N_28,In_17,In_270);
nor U29 (N_29,In_694,In_519);
or U30 (N_30,In_495,In_259);
nor U31 (N_31,In_16,In_481);
nand U32 (N_32,In_329,In_364);
or U33 (N_33,In_397,In_100);
xnor U34 (N_34,In_555,In_676);
or U35 (N_35,In_455,In_80);
and U36 (N_36,In_503,In_644);
nand U37 (N_37,In_581,In_716);
nand U38 (N_38,In_244,In_366);
or U39 (N_39,In_671,In_517);
and U40 (N_40,In_321,In_81);
nand U41 (N_41,In_585,In_314);
and U42 (N_42,In_34,In_670);
xnor U43 (N_43,In_357,In_446);
nand U44 (N_44,In_293,In_132);
or U45 (N_45,In_155,In_54);
nand U46 (N_46,In_550,In_304);
and U47 (N_47,In_510,In_693);
nand U48 (N_48,In_210,In_601);
or U49 (N_49,In_660,In_69);
or U50 (N_50,In_383,In_465);
or U51 (N_51,In_595,In_661);
xor U52 (N_52,In_592,In_231);
nand U53 (N_53,In_351,In_717);
and U54 (N_54,In_695,In_347);
or U55 (N_55,In_367,In_303);
xnor U56 (N_56,In_619,In_173);
or U57 (N_57,In_118,In_102);
nor U58 (N_58,In_684,In_687);
nand U59 (N_59,In_192,In_655);
and U60 (N_60,In_86,In_126);
or U61 (N_61,In_45,In_656);
nand U62 (N_62,In_61,In_525);
or U63 (N_63,In_324,In_530);
nand U64 (N_64,In_443,In_691);
xor U65 (N_65,In_131,In_723);
nand U66 (N_66,In_35,In_197);
and U67 (N_67,In_564,In_390);
nor U68 (N_68,In_335,In_441);
or U69 (N_69,In_710,In_469);
nor U70 (N_70,In_311,In_307);
xnor U71 (N_71,In_415,In_20);
and U72 (N_72,In_609,In_728);
or U73 (N_73,In_111,In_42);
nand U74 (N_74,In_493,In_242);
and U75 (N_75,In_147,In_130);
nand U76 (N_76,In_686,In_243);
nand U77 (N_77,In_437,In_747);
or U78 (N_78,In_562,In_94);
nand U79 (N_79,In_705,In_707);
nand U80 (N_80,In_0,In_279);
nand U81 (N_81,In_158,In_306);
or U82 (N_82,In_301,In_191);
nor U83 (N_83,In_394,In_545);
and U84 (N_84,In_188,In_101);
or U85 (N_85,In_289,In_152);
nand U86 (N_86,In_590,In_355);
nand U87 (N_87,In_275,In_621);
nand U88 (N_88,In_514,In_706);
and U89 (N_89,In_583,In_486);
nand U90 (N_90,In_466,In_326);
nand U91 (N_91,In_460,In_520);
nand U92 (N_92,In_257,In_540);
nor U93 (N_93,In_309,In_327);
nor U94 (N_94,In_38,In_749);
and U95 (N_95,In_491,In_108);
nor U96 (N_96,In_630,In_429);
nand U97 (N_97,In_120,In_635);
nor U98 (N_98,In_438,In_740);
nand U99 (N_99,In_288,In_23);
nor U100 (N_100,In_229,In_263);
or U101 (N_101,In_64,In_194);
nor U102 (N_102,In_53,In_328);
xor U103 (N_103,In_167,In_235);
and U104 (N_104,In_214,In_389);
nor U105 (N_105,In_499,In_648);
and U106 (N_106,In_571,In_471);
nor U107 (N_107,In_354,In_62);
xor U108 (N_108,In_400,In_299);
or U109 (N_109,In_487,In_658);
nor U110 (N_110,In_613,In_391);
and U111 (N_111,In_315,In_654);
or U112 (N_112,In_375,In_10);
nor U113 (N_113,In_36,In_269);
or U114 (N_114,In_203,In_739);
or U115 (N_115,In_239,In_737);
nand U116 (N_116,In_578,In_382);
or U117 (N_117,In_109,In_542);
nand U118 (N_118,In_295,In_652);
or U119 (N_119,In_218,In_157);
xnor U120 (N_120,In_404,In_622);
nand U121 (N_121,In_160,In_424);
or U122 (N_122,In_513,In_711);
nor U123 (N_123,In_268,In_219);
and U124 (N_124,In_125,In_22);
and U125 (N_125,In_470,In_84);
nand U126 (N_126,In_361,In_141);
nand U127 (N_127,In_186,In_209);
or U128 (N_128,In_140,In_260);
or U129 (N_129,In_734,In_484);
nor U130 (N_130,In_228,In_206);
or U131 (N_131,In_411,In_234);
and U132 (N_132,In_169,In_39);
and U133 (N_133,In_551,In_71);
nand U134 (N_134,In_729,In_272);
or U135 (N_135,In_57,In_418);
or U136 (N_136,In_50,In_697);
and U137 (N_137,In_180,In_709);
nor U138 (N_138,In_608,In_55);
nor U139 (N_139,In_122,In_531);
nand U140 (N_140,In_2,In_392);
nor U141 (N_141,In_317,In_535);
nor U142 (N_142,In_461,In_467);
and U143 (N_143,In_735,In_316);
nand U144 (N_144,In_476,In_340);
nor U145 (N_145,In_70,In_52);
nand U146 (N_146,In_369,In_376);
or U147 (N_147,In_282,In_398);
and U148 (N_148,In_712,In_223);
and U149 (N_149,In_509,In_359);
and U150 (N_150,In_121,In_439);
or U151 (N_151,In_78,In_384);
and U152 (N_152,In_277,In_552);
nand U153 (N_153,In_485,In_640);
and U154 (N_154,In_110,In_406);
nor U155 (N_155,In_248,In_163);
nor U156 (N_156,In_453,In_27);
and U157 (N_157,In_25,In_594);
or U158 (N_158,In_628,In_156);
nor U159 (N_159,In_115,In_128);
xnor U160 (N_160,In_447,In_445);
nand U161 (N_161,In_607,In_430);
nand U162 (N_162,In_154,In_165);
and U163 (N_163,In_546,In_377);
or U164 (N_164,In_704,In_360);
nor U165 (N_165,In_106,In_488);
nand U166 (N_166,In_479,In_565);
nand U167 (N_167,In_715,In_124);
and U168 (N_168,In_745,In_220);
nand U169 (N_169,In_548,In_393);
or U170 (N_170,In_489,In_645);
and U171 (N_171,In_200,In_230);
and U172 (N_172,In_330,In_379);
nor U173 (N_173,In_341,In_216);
nor U174 (N_174,In_343,In_148);
nand U175 (N_175,In_419,In_305);
nor U176 (N_176,In_508,In_422);
nand U177 (N_177,In_472,In_620);
and U178 (N_178,In_212,In_647);
or U179 (N_179,In_629,In_420);
nor U180 (N_180,In_569,In_342);
and U181 (N_181,In_283,In_150);
nor U182 (N_182,In_249,In_176);
nand U183 (N_183,In_1,In_208);
and U184 (N_184,In_182,In_170);
or U185 (N_185,In_591,In_181);
xor U186 (N_186,In_336,In_602);
xor U187 (N_187,In_92,In_528);
nor U188 (N_188,In_127,In_185);
and U189 (N_189,In_171,In_417);
nor U190 (N_190,In_201,In_144);
or U191 (N_191,In_196,In_240);
and U192 (N_192,In_325,In_538);
or U193 (N_193,In_350,In_74);
nand U194 (N_194,In_534,In_6);
and U195 (N_195,In_164,In_589);
and U196 (N_196,In_412,In_588);
nor U197 (N_197,In_688,In_587);
nor U198 (N_198,In_673,In_99);
or U199 (N_199,In_319,In_617);
nor U200 (N_200,In_561,In_153);
nor U201 (N_201,In_261,In_444);
or U202 (N_202,In_541,In_236);
nor U203 (N_203,In_559,In_708);
and U204 (N_204,In_667,In_46);
or U205 (N_205,In_252,In_428);
xor U206 (N_206,In_213,In_237);
and U207 (N_207,In_523,In_65);
or U208 (N_208,In_643,In_241);
xor U209 (N_209,In_501,In_199);
and U210 (N_210,In_741,In_123);
or U211 (N_211,In_615,In_690);
nand U212 (N_212,In_107,In_238);
xor U213 (N_213,In_8,In_135);
nand U214 (N_214,In_674,In_205);
and U215 (N_215,In_600,In_189);
or U216 (N_216,In_586,In_462);
nand U217 (N_217,In_480,In_85);
nand U218 (N_218,In_651,In_529);
nand U219 (N_219,In_266,In_251);
xor U220 (N_220,In_427,In_677);
nand U221 (N_221,In_576,In_274);
nand U222 (N_222,In_574,In_262);
and U223 (N_223,In_222,In_533);
and U224 (N_224,In_663,In_88);
nand U225 (N_225,In_103,In_177);
xor U226 (N_226,In_675,In_627);
xor U227 (N_227,In_380,In_450);
nand U228 (N_228,In_506,In_318);
or U229 (N_229,In_41,In_454);
nand U230 (N_230,In_297,In_233);
nor U231 (N_231,In_572,In_162);
nor U232 (N_232,In_407,In_24);
nor U233 (N_233,In_40,In_685);
or U234 (N_234,In_145,In_168);
nand U235 (N_235,In_179,In_423);
and U236 (N_236,In_639,In_549);
or U237 (N_237,In_138,In_18);
or U238 (N_238,In_224,In_456);
nand U239 (N_239,In_611,In_626);
or U240 (N_240,In_386,In_308);
and U241 (N_241,In_665,In_287);
and U242 (N_242,In_313,In_136);
nor U243 (N_243,In_166,In_672);
nand U244 (N_244,In_9,In_536);
or U245 (N_245,In_312,In_458);
or U246 (N_246,In_87,In_178);
or U247 (N_247,In_421,In_436);
nand U248 (N_248,In_250,In_405);
and U249 (N_249,In_207,In_151);
nor U250 (N_250,In_48,In_51);
nand U251 (N_251,In_596,In_298);
and U252 (N_252,In_642,In_33);
nand U253 (N_253,In_76,In_526);
nor U254 (N_254,In_452,In_473);
nand U255 (N_255,In_174,In_267);
and U256 (N_256,In_133,In_659);
nor U257 (N_257,In_532,In_724);
nor U258 (N_258,In_246,In_290);
and U259 (N_259,In_597,In_703);
xnor U260 (N_260,In_527,In_477);
or U261 (N_261,In_19,In_7);
and U262 (N_262,In_334,In_730);
and U263 (N_263,In_278,In_348);
or U264 (N_264,In_175,In_255);
or U265 (N_265,In_641,In_43);
nor U266 (N_266,In_599,In_410);
or U267 (N_267,In_373,In_37);
or U268 (N_268,In_582,In_403);
nor U269 (N_269,In_666,In_96);
and U270 (N_270,In_554,In_215);
nand U271 (N_271,In_98,In_302);
xor U272 (N_272,In_49,In_112);
nor U273 (N_273,In_187,In_322);
nor U274 (N_274,In_143,In_713);
nor U275 (N_275,In_30,In_344);
nor U276 (N_276,In_413,In_634);
or U277 (N_277,In_746,In_743);
nor U278 (N_278,In_89,In_90);
nand U279 (N_279,In_396,In_32);
and U280 (N_280,In_649,In_492);
nand U281 (N_281,In_276,In_227);
nor U282 (N_282,In_368,In_668);
nor U283 (N_283,In_440,In_172);
xnor U284 (N_284,In_254,In_75);
xor U285 (N_285,In_320,In_95);
nor U286 (N_286,In_202,In_566);
and U287 (N_287,In_604,In_683);
nor U288 (N_288,In_190,In_356);
and U289 (N_289,In_732,In_13);
nor U290 (N_290,In_264,In_638);
nand U291 (N_291,In_568,In_232);
or U292 (N_292,In_605,In_378);
or U293 (N_293,In_245,In_73);
nor U294 (N_294,In_142,In_573);
and U295 (N_295,In_631,In_401);
and U296 (N_296,In_105,In_544);
and U297 (N_297,In_474,In_435);
xor U298 (N_298,In_93,In_610);
nor U299 (N_299,In_494,In_502);
and U300 (N_300,In_67,In_388);
and U301 (N_301,In_636,In_4);
or U302 (N_302,In_577,In_294);
nand U303 (N_303,In_714,In_725);
nor U304 (N_304,In_332,In_323);
nor U305 (N_305,In_58,In_727);
nand U306 (N_306,In_113,In_56);
or U307 (N_307,In_584,In_560);
nor U308 (N_308,In_116,In_247);
nor U309 (N_309,In_198,In_567);
or U310 (N_310,In_91,In_482);
or U311 (N_311,In_104,In_696);
and U312 (N_312,In_399,In_97);
or U313 (N_313,In_662,In_217);
nor U314 (N_314,In_353,In_226);
nor U315 (N_315,In_372,In_281);
or U316 (N_316,In_408,In_370);
and U317 (N_317,In_748,In_625);
and U318 (N_318,In_114,In_500);
nand U319 (N_319,In_83,In_60);
nand U320 (N_320,In_21,In_395);
nand U321 (N_321,In_183,In_346);
and U322 (N_322,In_3,In_434);
nor U323 (N_323,In_333,In_409);
nand U324 (N_324,In_345,In_603);
or U325 (N_325,In_522,In_253);
nand U326 (N_326,In_516,In_537);
or U327 (N_327,In_463,In_646);
or U328 (N_328,In_512,In_702);
or U329 (N_329,In_736,In_459);
and U330 (N_330,In_449,In_478);
and U331 (N_331,In_483,In_31);
nor U332 (N_332,In_679,In_511);
and U333 (N_333,In_349,In_504);
nand U334 (N_334,In_664,In_310);
nor U335 (N_335,In_742,In_722);
nand U336 (N_336,In_161,In_669);
or U337 (N_337,In_225,In_457);
or U338 (N_338,In_331,In_553);
nand U339 (N_339,In_300,In_575);
nor U340 (N_340,In_498,In_184);
nand U341 (N_341,In_381,In_44);
nand U342 (N_342,In_68,In_718);
and U343 (N_343,In_337,In_719);
or U344 (N_344,In_524,In_79);
and U345 (N_345,In_28,In_521);
or U346 (N_346,In_731,In_681);
and U347 (N_347,In_614,In_442);
xor U348 (N_348,In_26,In_11);
or U349 (N_349,In_698,In_653);
and U350 (N_350,In_515,In_556);
xor U351 (N_351,In_371,In_258);
xor U352 (N_352,In_432,In_374);
and U353 (N_353,In_543,In_358);
nor U354 (N_354,In_689,In_59);
nand U355 (N_355,In_580,In_490);
xor U356 (N_356,In_632,In_433);
or U357 (N_357,In_137,In_292);
or U358 (N_358,In_518,In_66);
nor U359 (N_359,In_593,In_139);
xnor U360 (N_360,In_682,In_726);
and U361 (N_361,In_497,In_286);
or U362 (N_362,In_618,In_221);
nor U363 (N_363,In_701,In_146);
nor U364 (N_364,In_363,In_29);
nor U365 (N_365,In_265,In_63);
or U366 (N_366,In_680,In_426);
xor U367 (N_367,In_14,In_425);
xnor U368 (N_368,In_193,In_362);
and U369 (N_369,In_507,In_624);
nor U370 (N_370,In_558,In_570);
or U371 (N_371,In_195,In_598);
or U372 (N_372,In_387,In_72);
nor U373 (N_373,In_352,In_616);
nand U374 (N_374,In_612,In_496);
xor U375 (N_375,In_158,In_628);
nand U376 (N_376,In_471,In_230);
xnor U377 (N_377,In_340,In_543);
nand U378 (N_378,In_497,In_191);
or U379 (N_379,In_589,In_245);
and U380 (N_380,In_453,In_600);
nand U381 (N_381,In_412,In_425);
or U382 (N_382,In_517,In_238);
or U383 (N_383,In_478,In_659);
nand U384 (N_384,In_128,In_276);
nand U385 (N_385,In_11,In_65);
and U386 (N_386,In_338,In_285);
or U387 (N_387,In_350,In_540);
or U388 (N_388,In_558,In_150);
or U389 (N_389,In_436,In_423);
and U390 (N_390,In_242,In_16);
or U391 (N_391,In_440,In_10);
nor U392 (N_392,In_399,In_253);
nor U393 (N_393,In_265,In_544);
nor U394 (N_394,In_258,In_411);
and U395 (N_395,In_373,In_326);
xnor U396 (N_396,In_688,In_337);
or U397 (N_397,In_208,In_253);
nand U398 (N_398,In_449,In_179);
or U399 (N_399,In_720,In_42);
nor U400 (N_400,In_634,In_60);
and U401 (N_401,In_191,In_612);
or U402 (N_402,In_529,In_416);
and U403 (N_403,In_623,In_411);
xnor U404 (N_404,In_234,In_121);
nor U405 (N_405,In_641,In_395);
nand U406 (N_406,In_179,In_683);
or U407 (N_407,In_203,In_139);
xor U408 (N_408,In_197,In_588);
nand U409 (N_409,In_292,In_82);
nor U410 (N_410,In_364,In_74);
nand U411 (N_411,In_473,In_646);
and U412 (N_412,In_665,In_626);
nand U413 (N_413,In_45,In_133);
or U414 (N_414,In_116,In_296);
and U415 (N_415,In_490,In_449);
nor U416 (N_416,In_105,In_537);
and U417 (N_417,In_135,In_206);
and U418 (N_418,In_398,In_74);
or U419 (N_419,In_734,In_627);
or U420 (N_420,In_749,In_170);
xor U421 (N_421,In_480,In_14);
or U422 (N_422,In_304,In_670);
nor U423 (N_423,In_603,In_334);
xor U424 (N_424,In_639,In_645);
nor U425 (N_425,In_628,In_657);
nand U426 (N_426,In_393,In_305);
and U427 (N_427,In_48,In_395);
and U428 (N_428,In_609,In_202);
xnor U429 (N_429,In_288,In_576);
or U430 (N_430,In_153,In_303);
nor U431 (N_431,In_716,In_84);
nand U432 (N_432,In_367,In_684);
nand U433 (N_433,In_559,In_340);
xnor U434 (N_434,In_363,In_36);
nand U435 (N_435,In_567,In_397);
or U436 (N_436,In_745,In_60);
nor U437 (N_437,In_517,In_323);
and U438 (N_438,In_150,In_481);
and U439 (N_439,In_512,In_310);
nand U440 (N_440,In_36,In_734);
or U441 (N_441,In_164,In_51);
and U442 (N_442,In_242,In_509);
or U443 (N_443,In_246,In_317);
nor U444 (N_444,In_402,In_563);
nor U445 (N_445,In_189,In_27);
nor U446 (N_446,In_597,In_250);
nand U447 (N_447,In_190,In_651);
nand U448 (N_448,In_663,In_214);
and U449 (N_449,In_280,In_661);
xnor U450 (N_450,In_309,In_581);
nand U451 (N_451,In_652,In_427);
and U452 (N_452,In_680,In_549);
and U453 (N_453,In_639,In_445);
nand U454 (N_454,In_554,In_184);
and U455 (N_455,In_187,In_606);
nor U456 (N_456,In_163,In_470);
or U457 (N_457,In_463,In_478);
or U458 (N_458,In_345,In_495);
nor U459 (N_459,In_387,In_242);
and U460 (N_460,In_263,In_660);
and U461 (N_461,In_507,In_186);
or U462 (N_462,In_149,In_659);
nor U463 (N_463,In_295,In_201);
nor U464 (N_464,In_600,In_451);
nor U465 (N_465,In_167,In_461);
or U466 (N_466,In_474,In_321);
or U467 (N_467,In_262,In_115);
xor U468 (N_468,In_407,In_279);
nand U469 (N_469,In_412,In_616);
xnor U470 (N_470,In_731,In_513);
xor U471 (N_471,In_251,In_471);
nand U472 (N_472,In_255,In_311);
nor U473 (N_473,In_158,In_302);
nand U474 (N_474,In_425,In_452);
and U475 (N_475,In_712,In_601);
or U476 (N_476,In_142,In_638);
and U477 (N_477,In_431,In_175);
nand U478 (N_478,In_325,In_486);
or U479 (N_479,In_17,In_740);
nand U480 (N_480,In_564,In_79);
xor U481 (N_481,In_539,In_732);
nand U482 (N_482,In_596,In_652);
nand U483 (N_483,In_378,In_15);
nor U484 (N_484,In_197,In_586);
nand U485 (N_485,In_180,In_738);
nor U486 (N_486,In_645,In_654);
or U487 (N_487,In_749,In_223);
and U488 (N_488,In_334,In_312);
and U489 (N_489,In_707,In_600);
xnor U490 (N_490,In_214,In_139);
xnor U491 (N_491,In_279,In_400);
or U492 (N_492,In_299,In_0);
or U493 (N_493,In_739,In_529);
or U494 (N_494,In_9,In_70);
xnor U495 (N_495,In_530,In_181);
nand U496 (N_496,In_503,In_307);
nor U497 (N_497,In_666,In_593);
nand U498 (N_498,In_631,In_622);
nor U499 (N_499,In_44,In_307);
nand U500 (N_500,In_200,In_521);
or U501 (N_501,In_157,In_453);
xnor U502 (N_502,In_321,In_730);
and U503 (N_503,In_489,In_300);
nor U504 (N_504,In_669,In_167);
or U505 (N_505,In_104,In_554);
nand U506 (N_506,In_599,In_577);
nand U507 (N_507,In_168,In_520);
and U508 (N_508,In_447,In_180);
xnor U509 (N_509,In_631,In_188);
nand U510 (N_510,In_551,In_221);
or U511 (N_511,In_165,In_47);
and U512 (N_512,In_261,In_488);
nor U513 (N_513,In_724,In_409);
nor U514 (N_514,In_131,In_80);
or U515 (N_515,In_109,In_58);
nor U516 (N_516,In_461,In_542);
nor U517 (N_517,In_490,In_124);
nand U518 (N_518,In_560,In_539);
nor U519 (N_519,In_17,In_275);
or U520 (N_520,In_646,In_30);
or U521 (N_521,In_356,In_199);
xnor U522 (N_522,In_38,In_34);
nand U523 (N_523,In_519,In_653);
nor U524 (N_524,In_69,In_218);
or U525 (N_525,In_134,In_617);
xor U526 (N_526,In_693,In_252);
xor U527 (N_527,In_687,In_624);
nand U528 (N_528,In_267,In_473);
nor U529 (N_529,In_224,In_200);
nor U530 (N_530,In_107,In_3);
nand U531 (N_531,In_387,In_640);
or U532 (N_532,In_431,In_495);
nand U533 (N_533,In_670,In_374);
nor U534 (N_534,In_3,In_394);
or U535 (N_535,In_182,In_615);
xor U536 (N_536,In_409,In_594);
nor U537 (N_537,In_627,In_574);
nor U538 (N_538,In_739,In_745);
and U539 (N_539,In_238,In_585);
nand U540 (N_540,In_270,In_476);
and U541 (N_541,In_663,In_510);
nor U542 (N_542,In_180,In_726);
and U543 (N_543,In_245,In_637);
xor U544 (N_544,In_359,In_287);
and U545 (N_545,In_241,In_631);
nor U546 (N_546,In_250,In_269);
and U547 (N_547,In_661,In_452);
and U548 (N_548,In_241,In_488);
or U549 (N_549,In_160,In_458);
nor U550 (N_550,In_431,In_187);
or U551 (N_551,In_403,In_624);
and U552 (N_552,In_174,In_199);
nor U553 (N_553,In_655,In_536);
nand U554 (N_554,In_109,In_280);
or U555 (N_555,In_71,In_683);
or U556 (N_556,In_49,In_238);
nand U557 (N_557,In_382,In_91);
and U558 (N_558,In_159,In_286);
or U559 (N_559,In_653,In_306);
and U560 (N_560,In_562,In_52);
nor U561 (N_561,In_77,In_214);
and U562 (N_562,In_204,In_691);
nor U563 (N_563,In_634,In_189);
nand U564 (N_564,In_243,In_16);
xnor U565 (N_565,In_368,In_715);
xor U566 (N_566,In_141,In_582);
nor U567 (N_567,In_530,In_29);
nor U568 (N_568,In_72,In_699);
or U569 (N_569,In_168,In_126);
nor U570 (N_570,In_320,In_652);
nor U571 (N_571,In_16,In_367);
nor U572 (N_572,In_557,In_296);
or U573 (N_573,In_470,In_747);
and U574 (N_574,In_67,In_616);
and U575 (N_575,In_193,In_105);
or U576 (N_576,In_614,In_661);
xor U577 (N_577,In_616,In_579);
or U578 (N_578,In_103,In_554);
and U579 (N_579,In_548,In_200);
nand U580 (N_580,In_46,In_353);
nor U581 (N_581,In_546,In_476);
nor U582 (N_582,In_252,In_31);
and U583 (N_583,In_245,In_690);
nand U584 (N_584,In_429,In_378);
nor U585 (N_585,In_559,In_317);
nand U586 (N_586,In_115,In_637);
and U587 (N_587,In_286,In_155);
nand U588 (N_588,In_580,In_727);
or U589 (N_589,In_343,In_608);
and U590 (N_590,In_73,In_242);
nor U591 (N_591,In_697,In_631);
nand U592 (N_592,In_243,In_405);
nor U593 (N_593,In_269,In_395);
or U594 (N_594,In_536,In_505);
or U595 (N_595,In_213,In_116);
and U596 (N_596,In_660,In_81);
nor U597 (N_597,In_446,In_9);
or U598 (N_598,In_640,In_477);
or U599 (N_599,In_412,In_397);
and U600 (N_600,In_37,In_504);
and U601 (N_601,In_555,In_569);
nand U602 (N_602,In_586,In_324);
nor U603 (N_603,In_382,In_161);
nor U604 (N_604,In_49,In_265);
nor U605 (N_605,In_186,In_637);
nor U606 (N_606,In_526,In_493);
nor U607 (N_607,In_688,In_630);
or U608 (N_608,In_427,In_512);
or U609 (N_609,In_18,In_63);
xnor U610 (N_610,In_149,In_54);
nor U611 (N_611,In_562,In_227);
nor U612 (N_612,In_426,In_126);
nor U613 (N_613,In_220,In_641);
and U614 (N_614,In_281,In_166);
or U615 (N_615,In_678,In_421);
and U616 (N_616,In_57,In_518);
nor U617 (N_617,In_151,In_90);
and U618 (N_618,In_655,In_665);
and U619 (N_619,In_709,In_16);
nor U620 (N_620,In_186,In_242);
and U621 (N_621,In_40,In_651);
nor U622 (N_622,In_41,In_478);
nand U623 (N_623,In_479,In_604);
or U624 (N_624,In_652,In_289);
and U625 (N_625,In_271,In_249);
or U626 (N_626,In_618,In_4);
nand U627 (N_627,In_241,In_397);
and U628 (N_628,In_468,In_577);
and U629 (N_629,In_723,In_6);
and U630 (N_630,In_594,In_41);
and U631 (N_631,In_591,In_671);
and U632 (N_632,In_309,In_272);
nor U633 (N_633,In_600,In_36);
nor U634 (N_634,In_343,In_451);
nor U635 (N_635,In_412,In_595);
nor U636 (N_636,In_304,In_212);
xor U637 (N_637,In_570,In_468);
nand U638 (N_638,In_267,In_537);
or U639 (N_639,In_359,In_342);
and U640 (N_640,In_564,In_70);
nand U641 (N_641,In_83,In_504);
nand U642 (N_642,In_30,In_148);
nand U643 (N_643,In_100,In_108);
or U644 (N_644,In_652,In_357);
nand U645 (N_645,In_6,In_541);
xor U646 (N_646,In_431,In_88);
nor U647 (N_647,In_238,In_424);
xor U648 (N_648,In_426,In_168);
nor U649 (N_649,In_714,In_41);
nor U650 (N_650,In_699,In_675);
nand U651 (N_651,In_746,In_106);
and U652 (N_652,In_222,In_568);
xor U653 (N_653,In_141,In_299);
xnor U654 (N_654,In_69,In_140);
nor U655 (N_655,In_96,In_286);
nand U656 (N_656,In_314,In_365);
xor U657 (N_657,In_146,In_643);
or U658 (N_658,In_551,In_632);
nor U659 (N_659,In_287,In_555);
and U660 (N_660,In_207,In_343);
and U661 (N_661,In_678,In_336);
or U662 (N_662,In_346,In_243);
nor U663 (N_663,In_492,In_83);
or U664 (N_664,In_629,In_477);
nor U665 (N_665,In_696,In_88);
nor U666 (N_666,In_738,In_358);
nand U667 (N_667,In_488,In_126);
and U668 (N_668,In_650,In_488);
or U669 (N_669,In_499,In_125);
and U670 (N_670,In_446,In_435);
nor U671 (N_671,In_251,In_690);
and U672 (N_672,In_532,In_24);
xnor U673 (N_673,In_315,In_424);
or U674 (N_674,In_184,In_285);
and U675 (N_675,In_401,In_180);
nand U676 (N_676,In_90,In_113);
or U677 (N_677,In_353,In_439);
nand U678 (N_678,In_344,In_125);
nand U679 (N_679,In_682,In_450);
nand U680 (N_680,In_91,In_669);
nand U681 (N_681,In_90,In_540);
and U682 (N_682,In_554,In_13);
and U683 (N_683,In_427,In_239);
and U684 (N_684,In_585,In_171);
and U685 (N_685,In_708,In_268);
and U686 (N_686,In_647,In_515);
and U687 (N_687,In_586,In_581);
and U688 (N_688,In_305,In_503);
nor U689 (N_689,In_507,In_549);
or U690 (N_690,In_399,In_261);
nand U691 (N_691,In_83,In_742);
nor U692 (N_692,In_309,In_31);
nor U693 (N_693,In_115,In_224);
nor U694 (N_694,In_302,In_418);
and U695 (N_695,In_700,In_712);
nand U696 (N_696,In_288,In_493);
nand U697 (N_697,In_136,In_358);
and U698 (N_698,In_445,In_306);
and U699 (N_699,In_528,In_738);
nor U700 (N_700,In_396,In_402);
and U701 (N_701,In_337,In_599);
and U702 (N_702,In_689,In_636);
xor U703 (N_703,In_27,In_674);
nor U704 (N_704,In_447,In_97);
xor U705 (N_705,In_477,In_597);
or U706 (N_706,In_534,In_394);
nand U707 (N_707,In_69,In_73);
nor U708 (N_708,In_199,In_583);
or U709 (N_709,In_381,In_499);
nor U710 (N_710,In_448,In_292);
or U711 (N_711,In_373,In_254);
and U712 (N_712,In_78,In_344);
or U713 (N_713,In_391,In_205);
xor U714 (N_714,In_702,In_228);
or U715 (N_715,In_466,In_256);
or U716 (N_716,In_464,In_544);
nand U717 (N_717,In_379,In_659);
nor U718 (N_718,In_3,In_407);
nor U719 (N_719,In_297,In_637);
nor U720 (N_720,In_394,In_587);
or U721 (N_721,In_363,In_59);
or U722 (N_722,In_414,In_672);
and U723 (N_723,In_543,In_573);
nor U724 (N_724,In_189,In_501);
and U725 (N_725,In_643,In_599);
nor U726 (N_726,In_324,In_475);
and U727 (N_727,In_217,In_317);
or U728 (N_728,In_585,In_301);
and U729 (N_729,In_749,In_73);
nor U730 (N_730,In_605,In_167);
or U731 (N_731,In_257,In_103);
or U732 (N_732,In_579,In_668);
and U733 (N_733,In_211,In_492);
and U734 (N_734,In_245,In_430);
and U735 (N_735,In_202,In_149);
nor U736 (N_736,In_124,In_424);
and U737 (N_737,In_620,In_686);
nor U738 (N_738,In_492,In_340);
or U739 (N_739,In_171,In_404);
nor U740 (N_740,In_437,In_208);
nand U741 (N_741,In_11,In_626);
nand U742 (N_742,In_250,In_259);
and U743 (N_743,In_409,In_692);
nor U744 (N_744,In_668,In_562);
or U745 (N_745,In_462,In_491);
nand U746 (N_746,In_585,In_311);
xor U747 (N_747,In_299,In_429);
and U748 (N_748,In_238,In_147);
or U749 (N_749,In_717,In_99);
nand U750 (N_750,In_279,In_713);
and U751 (N_751,In_512,In_153);
or U752 (N_752,In_407,In_440);
nand U753 (N_753,In_527,In_603);
nor U754 (N_754,In_676,In_487);
nand U755 (N_755,In_339,In_382);
or U756 (N_756,In_114,In_190);
and U757 (N_757,In_46,In_44);
or U758 (N_758,In_189,In_62);
or U759 (N_759,In_410,In_182);
nand U760 (N_760,In_463,In_625);
nor U761 (N_761,In_20,In_744);
xor U762 (N_762,In_407,In_16);
nand U763 (N_763,In_700,In_100);
and U764 (N_764,In_611,In_113);
or U765 (N_765,In_266,In_371);
or U766 (N_766,In_37,In_674);
nor U767 (N_767,In_266,In_669);
nor U768 (N_768,In_323,In_555);
or U769 (N_769,In_189,In_671);
nand U770 (N_770,In_58,In_201);
and U771 (N_771,In_238,In_481);
or U772 (N_772,In_423,In_294);
nand U773 (N_773,In_325,In_380);
nand U774 (N_774,In_278,In_202);
xor U775 (N_775,In_201,In_291);
nor U776 (N_776,In_411,In_103);
nor U777 (N_777,In_254,In_54);
or U778 (N_778,In_586,In_223);
nor U779 (N_779,In_197,In_640);
and U780 (N_780,In_728,In_243);
xor U781 (N_781,In_411,In_235);
and U782 (N_782,In_614,In_51);
and U783 (N_783,In_215,In_478);
and U784 (N_784,In_556,In_406);
or U785 (N_785,In_374,In_375);
or U786 (N_786,In_400,In_219);
nand U787 (N_787,In_377,In_599);
xnor U788 (N_788,In_374,In_358);
or U789 (N_789,In_458,In_298);
nand U790 (N_790,In_332,In_657);
nand U791 (N_791,In_729,In_528);
or U792 (N_792,In_147,In_371);
and U793 (N_793,In_86,In_414);
nand U794 (N_794,In_481,In_715);
or U795 (N_795,In_40,In_609);
nand U796 (N_796,In_417,In_186);
nor U797 (N_797,In_703,In_67);
nor U798 (N_798,In_127,In_507);
nand U799 (N_799,In_605,In_662);
nor U800 (N_800,In_112,In_412);
nand U801 (N_801,In_699,In_622);
or U802 (N_802,In_108,In_319);
nor U803 (N_803,In_170,In_514);
or U804 (N_804,In_650,In_280);
and U805 (N_805,In_188,In_302);
nor U806 (N_806,In_185,In_299);
nand U807 (N_807,In_119,In_39);
nand U808 (N_808,In_65,In_36);
nor U809 (N_809,In_579,In_346);
and U810 (N_810,In_112,In_189);
nor U811 (N_811,In_186,In_32);
or U812 (N_812,In_688,In_650);
nor U813 (N_813,In_0,In_171);
xnor U814 (N_814,In_231,In_264);
or U815 (N_815,In_98,In_286);
nor U816 (N_816,In_749,In_420);
or U817 (N_817,In_66,In_87);
and U818 (N_818,In_134,In_124);
or U819 (N_819,In_194,In_688);
and U820 (N_820,In_435,In_580);
or U821 (N_821,In_691,In_180);
nor U822 (N_822,In_372,In_605);
nor U823 (N_823,In_174,In_249);
nand U824 (N_824,In_162,In_180);
and U825 (N_825,In_686,In_379);
or U826 (N_826,In_675,In_648);
nor U827 (N_827,In_527,In_1);
xnor U828 (N_828,In_2,In_306);
and U829 (N_829,In_376,In_159);
and U830 (N_830,In_9,In_212);
and U831 (N_831,In_344,In_213);
xor U832 (N_832,In_370,In_499);
or U833 (N_833,In_342,In_385);
and U834 (N_834,In_374,In_97);
and U835 (N_835,In_579,In_367);
xnor U836 (N_836,In_432,In_598);
nor U837 (N_837,In_581,In_348);
or U838 (N_838,In_398,In_560);
nor U839 (N_839,In_271,In_730);
nor U840 (N_840,In_344,In_179);
or U841 (N_841,In_500,In_659);
nand U842 (N_842,In_403,In_86);
or U843 (N_843,In_662,In_127);
nor U844 (N_844,In_315,In_118);
nor U845 (N_845,In_503,In_51);
or U846 (N_846,In_447,In_38);
or U847 (N_847,In_81,In_255);
or U848 (N_848,In_84,In_213);
nor U849 (N_849,In_156,In_371);
nor U850 (N_850,In_415,In_5);
nand U851 (N_851,In_587,In_389);
and U852 (N_852,In_451,In_491);
and U853 (N_853,In_448,In_484);
and U854 (N_854,In_566,In_299);
xnor U855 (N_855,In_27,In_542);
xor U856 (N_856,In_638,In_99);
nor U857 (N_857,In_725,In_606);
or U858 (N_858,In_615,In_260);
nand U859 (N_859,In_525,In_33);
nor U860 (N_860,In_695,In_130);
and U861 (N_861,In_470,In_311);
and U862 (N_862,In_556,In_502);
nand U863 (N_863,In_490,In_519);
nor U864 (N_864,In_280,In_283);
nor U865 (N_865,In_712,In_743);
nor U866 (N_866,In_463,In_552);
nor U867 (N_867,In_442,In_368);
or U868 (N_868,In_68,In_122);
and U869 (N_869,In_41,In_705);
nand U870 (N_870,In_534,In_519);
and U871 (N_871,In_691,In_480);
nor U872 (N_872,In_298,In_385);
nand U873 (N_873,In_210,In_285);
and U874 (N_874,In_486,In_297);
nand U875 (N_875,In_143,In_626);
xor U876 (N_876,In_727,In_341);
nand U877 (N_877,In_457,In_238);
nand U878 (N_878,In_668,In_426);
nand U879 (N_879,In_489,In_30);
nor U880 (N_880,In_545,In_199);
or U881 (N_881,In_646,In_137);
and U882 (N_882,In_474,In_236);
xnor U883 (N_883,In_436,In_651);
xnor U884 (N_884,In_418,In_225);
xor U885 (N_885,In_135,In_67);
xnor U886 (N_886,In_54,In_268);
nand U887 (N_887,In_185,In_276);
xor U888 (N_888,In_420,In_345);
nand U889 (N_889,In_51,In_285);
and U890 (N_890,In_335,In_446);
nand U891 (N_891,In_53,In_519);
xor U892 (N_892,In_688,In_545);
and U893 (N_893,In_544,In_75);
nand U894 (N_894,In_671,In_31);
and U895 (N_895,In_223,In_392);
or U896 (N_896,In_749,In_628);
nand U897 (N_897,In_162,In_41);
and U898 (N_898,In_358,In_476);
and U899 (N_899,In_590,In_23);
nor U900 (N_900,In_391,In_15);
and U901 (N_901,In_249,In_204);
and U902 (N_902,In_490,In_520);
and U903 (N_903,In_30,In_597);
and U904 (N_904,In_65,In_706);
or U905 (N_905,In_647,In_150);
and U906 (N_906,In_450,In_214);
or U907 (N_907,In_400,In_143);
or U908 (N_908,In_736,In_301);
nor U909 (N_909,In_698,In_216);
nor U910 (N_910,In_706,In_170);
nand U911 (N_911,In_135,In_657);
nand U912 (N_912,In_391,In_740);
or U913 (N_913,In_41,In_474);
or U914 (N_914,In_170,In_622);
and U915 (N_915,In_51,In_77);
nor U916 (N_916,In_261,In_416);
and U917 (N_917,In_387,In_659);
xor U918 (N_918,In_592,In_524);
and U919 (N_919,In_22,In_747);
nor U920 (N_920,In_242,In_679);
xor U921 (N_921,In_168,In_323);
nor U922 (N_922,In_305,In_693);
nor U923 (N_923,In_526,In_31);
or U924 (N_924,In_642,In_395);
nand U925 (N_925,In_555,In_637);
and U926 (N_926,In_717,In_188);
or U927 (N_927,In_526,In_722);
and U928 (N_928,In_363,In_308);
nand U929 (N_929,In_547,In_313);
nor U930 (N_930,In_638,In_663);
and U931 (N_931,In_184,In_661);
nand U932 (N_932,In_471,In_19);
or U933 (N_933,In_650,In_742);
nor U934 (N_934,In_725,In_703);
nor U935 (N_935,In_715,In_625);
or U936 (N_936,In_563,In_578);
or U937 (N_937,In_269,In_117);
xnor U938 (N_938,In_611,In_99);
or U939 (N_939,In_365,In_107);
and U940 (N_940,In_716,In_635);
nor U941 (N_941,In_89,In_216);
nor U942 (N_942,In_581,In_46);
xnor U943 (N_943,In_466,In_489);
nor U944 (N_944,In_253,In_86);
xnor U945 (N_945,In_651,In_587);
or U946 (N_946,In_429,In_519);
or U947 (N_947,In_288,In_133);
nor U948 (N_948,In_719,In_67);
nand U949 (N_949,In_506,In_747);
and U950 (N_950,In_371,In_418);
or U951 (N_951,In_64,In_338);
and U952 (N_952,In_581,In_21);
and U953 (N_953,In_637,In_585);
xnor U954 (N_954,In_373,In_487);
nand U955 (N_955,In_689,In_196);
or U956 (N_956,In_82,In_277);
nor U957 (N_957,In_724,In_117);
and U958 (N_958,In_274,In_446);
and U959 (N_959,In_276,In_291);
xor U960 (N_960,In_277,In_309);
nor U961 (N_961,In_705,In_675);
and U962 (N_962,In_176,In_676);
or U963 (N_963,In_71,In_238);
and U964 (N_964,In_515,In_449);
or U965 (N_965,In_652,In_505);
nor U966 (N_966,In_297,In_743);
and U967 (N_967,In_713,In_712);
or U968 (N_968,In_227,In_733);
and U969 (N_969,In_159,In_375);
nor U970 (N_970,In_206,In_218);
nor U971 (N_971,In_55,In_56);
nor U972 (N_972,In_270,In_177);
or U973 (N_973,In_245,In_480);
or U974 (N_974,In_557,In_319);
nand U975 (N_975,In_281,In_734);
or U976 (N_976,In_189,In_14);
and U977 (N_977,In_201,In_109);
and U978 (N_978,In_136,In_740);
or U979 (N_979,In_667,In_375);
and U980 (N_980,In_121,In_244);
and U981 (N_981,In_5,In_488);
xor U982 (N_982,In_722,In_512);
and U983 (N_983,In_637,In_154);
and U984 (N_984,In_212,In_537);
and U985 (N_985,In_743,In_162);
nand U986 (N_986,In_668,In_219);
and U987 (N_987,In_331,In_176);
nand U988 (N_988,In_245,In_83);
and U989 (N_989,In_347,In_273);
or U990 (N_990,In_390,In_548);
nand U991 (N_991,In_251,In_637);
nor U992 (N_992,In_417,In_562);
or U993 (N_993,In_291,In_314);
nand U994 (N_994,In_652,In_173);
and U995 (N_995,In_446,In_353);
or U996 (N_996,In_729,In_480);
nand U997 (N_997,In_111,In_618);
xnor U998 (N_998,In_602,In_128);
nand U999 (N_999,In_674,In_391);
nand U1000 (N_1000,In_183,In_464);
nand U1001 (N_1001,In_28,In_345);
nor U1002 (N_1002,In_691,In_676);
or U1003 (N_1003,In_626,In_291);
and U1004 (N_1004,In_407,In_301);
nor U1005 (N_1005,In_352,In_487);
nor U1006 (N_1006,In_542,In_402);
nand U1007 (N_1007,In_475,In_720);
nor U1008 (N_1008,In_472,In_311);
nand U1009 (N_1009,In_550,In_667);
and U1010 (N_1010,In_139,In_134);
xor U1011 (N_1011,In_344,In_23);
and U1012 (N_1012,In_595,In_109);
nand U1013 (N_1013,In_363,In_317);
and U1014 (N_1014,In_164,In_320);
nand U1015 (N_1015,In_140,In_426);
and U1016 (N_1016,In_305,In_689);
xor U1017 (N_1017,In_156,In_212);
nor U1018 (N_1018,In_290,In_171);
nand U1019 (N_1019,In_116,In_566);
and U1020 (N_1020,In_52,In_119);
nor U1021 (N_1021,In_222,In_466);
nor U1022 (N_1022,In_330,In_147);
and U1023 (N_1023,In_739,In_239);
and U1024 (N_1024,In_446,In_407);
nor U1025 (N_1025,In_488,In_88);
nor U1026 (N_1026,In_122,In_75);
and U1027 (N_1027,In_497,In_485);
xor U1028 (N_1028,In_219,In_260);
or U1029 (N_1029,In_456,In_178);
nand U1030 (N_1030,In_717,In_266);
xnor U1031 (N_1031,In_169,In_322);
or U1032 (N_1032,In_135,In_306);
nor U1033 (N_1033,In_210,In_449);
and U1034 (N_1034,In_15,In_527);
and U1035 (N_1035,In_345,In_565);
nor U1036 (N_1036,In_159,In_429);
nor U1037 (N_1037,In_116,In_144);
nor U1038 (N_1038,In_684,In_532);
xor U1039 (N_1039,In_8,In_213);
or U1040 (N_1040,In_221,In_365);
nand U1041 (N_1041,In_570,In_14);
nand U1042 (N_1042,In_63,In_536);
nor U1043 (N_1043,In_451,In_724);
xor U1044 (N_1044,In_286,In_322);
nand U1045 (N_1045,In_380,In_693);
or U1046 (N_1046,In_235,In_193);
nand U1047 (N_1047,In_607,In_609);
xnor U1048 (N_1048,In_422,In_427);
nor U1049 (N_1049,In_71,In_275);
or U1050 (N_1050,In_275,In_117);
nor U1051 (N_1051,In_327,In_294);
and U1052 (N_1052,In_659,In_507);
nand U1053 (N_1053,In_347,In_637);
and U1054 (N_1054,In_220,In_650);
nand U1055 (N_1055,In_409,In_138);
and U1056 (N_1056,In_22,In_267);
or U1057 (N_1057,In_738,In_119);
or U1058 (N_1058,In_491,In_407);
or U1059 (N_1059,In_64,In_518);
nor U1060 (N_1060,In_368,In_18);
or U1061 (N_1061,In_521,In_151);
and U1062 (N_1062,In_257,In_679);
nor U1063 (N_1063,In_203,In_625);
or U1064 (N_1064,In_248,In_293);
nand U1065 (N_1065,In_533,In_509);
nand U1066 (N_1066,In_559,In_97);
nand U1067 (N_1067,In_732,In_501);
xor U1068 (N_1068,In_2,In_292);
or U1069 (N_1069,In_255,In_8);
or U1070 (N_1070,In_435,In_605);
nand U1071 (N_1071,In_534,In_704);
nand U1072 (N_1072,In_619,In_15);
nand U1073 (N_1073,In_209,In_281);
or U1074 (N_1074,In_507,In_612);
xor U1075 (N_1075,In_438,In_599);
nor U1076 (N_1076,In_514,In_426);
or U1077 (N_1077,In_312,In_327);
nor U1078 (N_1078,In_527,In_414);
and U1079 (N_1079,In_377,In_254);
nor U1080 (N_1080,In_69,In_156);
nor U1081 (N_1081,In_615,In_503);
and U1082 (N_1082,In_413,In_498);
or U1083 (N_1083,In_256,In_151);
and U1084 (N_1084,In_246,In_386);
or U1085 (N_1085,In_272,In_655);
xnor U1086 (N_1086,In_240,In_275);
nand U1087 (N_1087,In_188,In_332);
nand U1088 (N_1088,In_265,In_275);
nand U1089 (N_1089,In_71,In_388);
nand U1090 (N_1090,In_732,In_399);
nand U1091 (N_1091,In_1,In_494);
and U1092 (N_1092,In_648,In_693);
or U1093 (N_1093,In_50,In_710);
and U1094 (N_1094,In_687,In_147);
or U1095 (N_1095,In_165,In_498);
nand U1096 (N_1096,In_323,In_328);
or U1097 (N_1097,In_740,In_319);
xnor U1098 (N_1098,In_441,In_218);
and U1099 (N_1099,In_738,In_692);
xnor U1100 (N_1100,In_22,In_228);
and U1101 (N_1101,In_407,In_141);
xnor U1102 (N_1102,In_730,In_150);
nor U1103 (N_1103,In_3,In_43);
or U1104 (N_1104,In_415,In_505);
xor U1105 (N_1105,In_721,In_399);
nand U1106 (N_1106,In_260,In_653);
nand U1107 (N_1107,In_233,In_221);
or U1108 (N_1108,In_582,In_9);
nand U1109 (N_1109,In_27,In_675);
nand U1110 (N_1110,In_646,In_533);
nor U1111 (N_1111,In_452,In_607);
nand U1112 (N_1112,In_584,In_189);
nor U1113 (N_1113,In_594,In_522);
nand U1114 (N_1114,In_640,In_381);
or U1115 (N_1115,In_283,In_618);
or U1116 (N_1116,In_179,In_347);
or U1117 (N_1117,In_386,In_107);
or U1118 (N_1118,In_545,In_716);
and U1119 (N_1119,In_436,In_394);
or U1120 (N_1120,In_307,In_1);
nand U1121 (N_1121,In_189,In_149);
nand U1122 (N_1122,In_31,In_642);
or U1123 (N_1123,In_740,In_604);
or U1124 (N_1124,In_32,In_543);
or U1125 (N_1125,In_340,In_114);
or U1126 (N_1126,In_302,In_284);
xor U1127 (N_1127,In_556,In_248);
and U1128 (N_1128,In_563,In_455);
nand U1129 (N_1129,In_659,In_71);
and U1130 (N_1130,In_603,In_107);
xor U1131 (N_1131,In_20,In_149);
or U1132 (N_1132,In_95,In_196);
and U1133 (N_1133,In_355,In_233);
nand U1134 (N_1134,In_460,In_58);
nor U1135 (N_1135,In_32,In_213);
xor U1136 (N_1136,In_642,In_714);
nor U1137 (N_1137,In_89,In_398);
and U1138 (N_1138,In_371,In_703);
xor U1139 (N_1139,In_206,In_524);
or U1140 (N_1140,In_273,In_193);
nor U1141 (N_1141,In_573,In_110);
nand U1142 (N_1142,In_359,In_665);
or U1143 (N_1143,In_622,In_407);
and U1144 (N_1144,In_729,In_15);
or U1145 (N_1145,In_633,In_81);
nand U1146 (N_1146,In_268,In_635);
or U1147 (N_1147,In_495,In_673);
nand U1148 (N_1148,In_152,In_67);
or U1149 (N_1149,In_378,In_482);
nand U1150 (N_1150,In_745,In_25);
nor U1151 (N_1151,In_514,In_672);
or U1152 (N_1152,In_13,In_576);
nand U1153 (N_1153,In_566,In_616);
xnor U1154 (N_1154,In_268,In_599);
or U1155 (N_1155,In_525,In_573);
nor U1156 (N_1156,In_404,In_205);
and U1157 (N_1157,In_472,In_719);
nor U1158 (N_1158,In_441,In_655);
nand U1159 (N_1159,In_2,In_678);
and U1160 (N_1160,In_481,In_181);
or U1161 (N_1161,In_14,In_692);
nor U1162 (N_1162,In_613,In_575);
xnor U1163 (N_1163,In_400,In_686);
nand U1164 (N_1164,In_559,In_79);
nand U1165 (N_1165,In_55,In_216);
xor U1166 (N_1166,In_29,In_444);
or U1167 (N_1167,In_589,In_16);
and U1168 (N_1168,In_404,In_693);
nand U1169 (N_1169,In_647,In_574);
and U1170 (N_1170,In_134,In_174);
nor U1171 (N_1171,In_442,In_127);
nand U1172 (N_1172,In_73,In_144);
nor U1173 (N_1173,In_190,In_677);
and U1174 (N_1174,In_16,In_62);
nand U1175 (N_1175,In_338,In_289);
or U1176 (N_1176,In_690,In_183);
xor U1177 (N_1177,In_679,In_409);
and U1178 (N_1178,In_385,In_312);
xnor U1179 (N_1179,In_36,In_408);
and U1180 (N_1180,In_162,In_611);
nand U1181 (N_1181,In_375,In_15);
nand U1182 (N_1182,In_52,In_639);
and U1183 (N_1183,In_380,In_466);
or U1184 (N_1184,In_319,In_101);
and U1185 (N_1185,In_444,In_602);
or U1186 (N_1186,In_201,In_128);
and U1187 (N_1187,In_382,In_481);
xnor U1188 (N_1188,In_6,In_262);
and U1189 (N_1189,In_597,In_732);
nor U1190 (N_1190,In_431,In_365);
and U1191 (N_1191,In_631,In_616);
nand U1192 (N_1192,In_247,In_410);
nand U1193 (N_1193,In_524,In_0);
or U1194 (N_1194,In_608,In_338);
or U1195 (N_1195,In_473,In_557);
and U1196 (N_1196,In_201,In_494);
xnor U1197 (N_1197,In_731,In_128);
or U1198 (N_1198,In_605,In_646);
and U1199 (N_1199,In_390,In_74);
nor U1200 (N_1200,In_558,In_66);
or U1201 (N_1201,In_729,In_353);
or U1202 (N_1202,In_124,In_370);
nand U1203 (N_1203,In_493,In_681);
nor U1204 (N_1204,In_357,In_450);
nor U1205 (N_1205,In_702,In_407);
nand U1206 (N_1206,In_288,In_461);
xnor U1207 (N_1207,In_522,In_509);
or U1208 (N_1208,In_71,In_232);
xor U1209 (N_1209,In_136,In_421);
or U1210 (N_1210,In_675,In_196);
nand U1211 (N_1211,In_364,In_306);
nor U1212 (N_1212,In_676,In_633);
nand U1213 (N_1213,In_460,In_260);
nor U1214 (N_1214,In_17,In_639);
or U1215 (N_1215,In_365,In_312);
nand U1216 (N_1216,In_137,In_174);
nand U1217 (N_1217,In_53,In_317);
nor U1218 (N_1218,In_159,In_138);
or U1219 (N_1219,In_90,In_205);
nor U1220 (N_1220,In_386,In_153);
xnor U1221 (N_1221,In_310,In_217);
or U1222 (N_1222,In_328,In_473);
nor U1223 (N_1223,In_598,In_690);
and U1224 (N_1224,In_664,In_559);
nand U1225 (N_1225,In_623,In_129);
xor U1226 (N_1226,In_140,In_314);
or U1227 (N_1227,In_247,In_299);
and U1228 (N_1228,In_585,In_178);
nor U1229 (N_1229,In_737,In_683);
and U1230 (N_1230,In_212,In_569);
nor U1231 (N_1231,In_682,In_137);
or U1232 (N_1232,In_422,In_281);
nand U1233 (N_1233,In_447,In_441);
and U1234 (N_1234,In_665,In_272);
nand U1235 (N_1235,In_485,In_220);
nand U1236 (N_1236,In_230,In_368);
or U1237 (N_1237,In_184,In_242);
nor U1238 (N_1238,In_234,In_194);
nand U1239 (N_1239,In_291,In_641);
or U1240 (N_1240,In_181,In_363);
nor U1241 (N_1241,In_541,In_129);
nand U1242 (N_1242,In_683,In_552);
nand U1243 (N_1243,In_373,In_47);
nor U1244 (N_1244,In_147,In_35);
xor U1245 (N_1245,In_441,In_708);
nand U1246 (N_1246,In_226,In_152);
nor U1247 (N_1247,In_522,In_57);
and U1248 (N_1248,In_98,In_634);
nor U1249 (N_1249,In_637,In_649);
and U1250 (N_1250,In_574,In_395);
nor U1251 (N_1251,In_589,In_182);
nand U1252 (N_1252,In_378,In_29);
and U1253 (N_1253,In_450,In_165);
and U1254 (N_1254,In_8,In_612);
and U1255 (N_1255,In_394,In_468);
nor U1256 (N_1256,In_306,In_519);
nand U1257 (N_1257,In_399,In_565);
xnor U1258 (N_1258,In_413,In_504);
nor U1259 (N_1259,In_141,In_700);
or U1260 (N_1260,In_57,In_45);
and U1261 (N_1261,In_721,In_240);
and U1262 (N_1262,In_415,In_732);
nor U1263 (N_1263,In_585,In_353);
nor U1264 (N_1264,In_2,In_476);
xor U1265 (N_1265,In_433,In_541);
nand U1266 (N_1266,In_336,In_469);
xnor U1267 (N_1267,In_361,In_230);
nor U1268 (N_1268,In_360,In_220);
nand U1269 (N_1269,In_82,In_387);
nor U1270 (N_1270,In_80,In_742);
and U1271 (N_1271,In_52,In_480);
and U1272 (N_1272,In_253,In_422);
nand U1273 (N_1273,In_519,In_182);
or U1274 (N_1274,In_316,In_708);
xor U1275 (N_1275,In_478,In_156);
nor U1276 (N_1276,In_669,In_197);
and U1277 (N_1277,In_248,In_51);
and U1278 (N_1278,In_102,In_130);
nand U1279 (N_1279,In_720,In_69);
and U1280 (N_1280,In_661,In_478);
nand U1281 (N_1281,In_735,In_91);
nor U1282 (N_1282,In_647,In_659);
and U1283 (N_1283,In_118,In_458);
nor U1284 (N_1284,In_312,In_413);
or U1285 (N_1285,In_142,In_5);
and U1286 (N_1286,In_713,In_97);
or U1287 (N_1287,In_19,In_517);
xnor U1288 (N_1288,In_325,In_38);
nand U1289 (N_1289,In_449,In_251);
and U1290 (N_1290,In_358,In_607);
or U1291 (N_1291,In_129,In_109);
xnor U1292 (N_1292,In_714,In_393);
or U1293 (N_1293,In_219,In_403);
nand U1294 (N_1294,In_715,In_446);
and U1295 (N_1295,In_708,In_516);
or U1296 (N_1296,In_507,In_83);
nor U1297 (N_1297,In_682,In_65);
nor U1298 (N_1298,In_199,In_202);
nand U1299 (N_1299,In_696,In_98);
nand U1300 (N_1300,In_466,In_299);
and U1301 (N_1301,In_171,In_351);
or U1302 (N_1302,In_678,In_572);
nor U1303 (N_1303,In_658,In_98);
nor U1304 (N_1304,In_655,In_578);
nand U1305 (N_1305,In_93,In_156);
and U1306 (N_1306,In_61,In_67);
or U1307 (N_1307,In_571,In_348);
or U1308 (N_1308,In_483,In_405);
and U1309 (N_1309,In_709,In_344);
xnor U1310 (N_1310,In_729,In_547);
or U1311 (N_1311,In_266,In_357);
nand U1312 (N_1312,In_545,In_382);
and U1313 (N_1313,In_552,In_470);
nor U1314 (N_1314,In_214,In_500);
and U1315 (N_1315,In_203,In_9);
and U1316 (N_1316,In_598,In_187);
nand U1317 (N_1317,In_164,In_453);
or U1318 (N_1318,In_318,In_403);
nand U1319 (N_1319,In_444,In_176);
nor U1320 (N_1320,In_616,In_360);
nand U1321 (N_1321,In_182,In_175);
or U1322 (N_1322,In_413,In_102);
nor U1323 (N_1323,In_727,In_16);
nand U1324 (N_1324,In_63,In_538);
or U1325 (N_1325,In_178,In_448);
nor U1326 (N_1326,In_596,In_644);
nand U1327 (N_1327,In_340,In_66);
nor U1328 (N_1328,In_565,In_233);
xor U1329 (N_1329,In_263,In_267);
or U1330 (N_1330,In_544,In_37);
nand U1331 (N_1331,In_636,In_255);
nor U1332 (N_1332,In_709,In_484);
xor U1333 (N_1333,In_308,In_693);
or U1334 (N_1334,In_141,In_241);
nand U1335 (N_1335,In_103,In_375);
nor U1336 (N_1336,In_85,In_368);
or U1337 (N_1337,In_503,In_700);
and U1338 (N_1338,In_478,In_437);
nor U1339 (N_1339,In_564,In_672);
and U1340 (N_1340,In_541,In_427);
nor U1341 (N_1341,In_46,In_356);
and U1342 (N_1342,In_677,In_400);
nand U1343 (N_1343,In_623,In_600);
and U1344 (N_1344,In_656,In_378);
nand U1345 (N_1345,In_267,In_113);
nand U1346 (N_1346,In_554,In_504);
nand U1347 (N_1347,In_248,In_590);
nor U1348 (N_1348,In_127,In_652);
nor U1349 (N_1349,In_226,In_247);
or U1350 (N_1350,In_431,In_595);
nor U1351 (N_1351,In_16,In_636);
xor U1352 (N_1352,In_175,In_451);
and U1353 (N_1353,In_592,In_79);
xnor U1354 (N_1354,In_670,In_438);
nand U1355 (N_1355,In_642,In_618);
or U1356 (N_1356,In_616,In_636);
nor U1357 (N_1357,In_639,In_455);
nand U1358 (N_1358,In_498,In_708);
and U1359 (N_1359,In_188,In_656);
and U1360 (N_1360,In_321,In_496);
nand U1361 (N_1361,In_202,In_84);
nor U1362 (N_1362,In_451,In_26);
nand U1363 (N_1363,In_358,In_82);
and U1364 (N_1364,In_504,In_581);
nand U1365 (N_1365,In_462,In_317);
and U1366 (N_1366,In_17,In_228);
nor U1367 (N_1367,In_445,In_716);
nand U1368 (N_1368,In_280,In_569);
and U1369 (N_1369,In_236,In_191);
or U1370 (N_1370,In_91,In_591);
and U1371 (N_1371,In_4,In_651);
and U1372 (N_1372,In_407,In_738);
nand U1373 (N_1373,In_463,In_288);
xor U1374 (N_1374,In_217,In_689);
xnor U1375 (N_1375,In_568,In_244);
or U1376 (N_1376,In_719,In_213);
nand U1377 (N_1377,In_554,In_319);
nor U1378 (N_1378,In_248,In_503);
and U1379 (N_1379,In_155,In_633);
or U1380 (N_1380,In_665,In_494);
nor U1381 (N_1381,In_300,In_725);
nor U1382 (N_1382,In_500,In_411);
nand U1383 (N_1383,In_449,In_370);
and U1384 (N_1384,In_575,In_88);
nand U1385 (N_1385,In_166,In_359);
nor U1386 (N_1386,In_335,In_380);
or U1387 (N_1387,In_223,In_122);
nand U1388 (N_1388,In_347,In_47);
nand U1389 (N_1389,In_330,In_385);
and U1390 (N_1390,In_209,In_593);
or U1391 (N_1391,In_301,In_292);
nand U1392 (N_1392,In_513,In_577);
and U1393 (N_1393,In_439,In_270);
nor U1394 (N_1394,In_423,In_366);
xnor U1395 (N_1395,In_140,In_356);
nor U1396 (N_1396,In_614,In_334);
and U1397 (N_1397,In_109,In_43);
nand U1398 (N_1398,In_6,In_623);
or U1399 (N_1399,In_547,In_494);
xor U1400 (N_1400,In_370,In_633);
or U1401 (N_1401,In_411,In_741);
nand U1402 (N_1402,In_89,In_570);
or U1403 (N_1403,In_487,In_680);
or U1404 (N_1404,In_276,In_541);
nor U1405 (N_1405,In_645,In_641);
and U1406 (N_1406,In_11,In_247);
nand U1407 (N_1407,In_683,In_301);
nor U1408 (N_1408,In_564,In_261);
nand U1409 (N_1409,In_613,In_136);
and U1410 (N_1410,In_390,In_414);
or U1411 (N_1411,In_278,In_704);
or U1412 (N_1412,In_189,In_555);
and U1413 (N_1413,In_11,In_181);
and U1414 (N_1414,In_533,In_545);
nand U1415 (N_1415,In_711,In_147);
nor U1416 (N_1416,In_699,In_204);
nand U1417 (N_1417,In_585,In_448);
xnor U1418 (N_1418,In_746,In_390);
or U1419 (N_1419,In_215,In_279);
and U1420 (N_1420,In_203,In_638);
or U1421 (N_1421,In_614,In_734);
nor U1422 (N_1422,In_288,In_350);
and U1423 (N_1423,In_535,In_385);
or U1424 (N_1424,In_275,In_669);
nand U1425 (N_1425,In_214,In_422);
or U1426 (N_1426,In_473,In_269);
nand U1427 (N_1427,In_581,In_483);
nand U1428 (N_1428,In_269,In_246);
nand U1429 (N_1429,In_244,In_130);
nor U1430 (N_1430,In_281,In_46);
or U1431 (N_1431,In_34,In_189);
nor U1432 (N_1432,In_529,In_630);
nor U1433 (N_1433,In_678,In_240);
or U1434 (N_1434,In_76,In_53);
and U1435 (N_1435,In_203,In_385);
xnor U1436 (N_1436,In_456,In_98);
xor U1437 (N_1437,In_365,In_108);
nor U1438 (N_1438,In_171,In_153);
or U1439 (N_1439,In_747,In_580);
and U1440 (N_1440,In_623,In_272);
or U1441 (N_1441,In_735,In_729);
nor U1442 (N_1442,In_743,In_389);
or U1443 (N_1443,In_412,In_573);
nor U1444 (N_1444,In_369,In_609);
nor U1445 (N_1445,In_293,In_573);
and U1446 (N_1446,In_399,In_6);
nand U1447 (N_1447,In_466,In_114);
nor U1448 (N_1448,In_243,In_37);
or U1449 (N_1449,In_155,In_31);
or U1450 (N_1450,In_638,In_716);
nor U1451 (N_1451,In_739,In_70);
xnor U1452 (N_1452,In_601,In_130);
and U1453 (N_1453,In_554,In_633);
nand U1454 (N_1454,In_288,In_3);
nor U1455 (N_1455,In_442,In_544);
and U1456 (N_1456,In_387,In_497);
nor U1457 (N_1457,In_6,In_134);
nand U1458 (N_1458,In_568,In_639);
and U1459 (N_1459,In_672,In_589);
or U1460 (N_1460,In_234,In_2);
and U1461 (N_1461,In_188,In_405);
and U1462 (N_1462,In_356,In_509);
nor U1463 (N_1463,In_448,In_471);
and U1464 (N_1464,In_54,In_289);
or U1465 (N_1465,In_749,In_393);
nor U1466 (N_1466,In_541,In_704);
and U1467 (N_1467,In_137,In_61);
and U1468 (N_1468,In_725,In_607);
and U1469 (N_1469,In_529,In_315);
or U1470 (N_1470,In_535,In_637);
and U1471 (N_1471,In_191,In_741);
or U1472 (N_1472,In_557,In_721);
nand U1473 (N_1473,In_93,In_146);
xnor U1474 (N_1474,In_70,In_291);
or U1475 (N_1475,In_633,In_486);
or U1476 (N_1476,In_566,In_729);
nand U1477 (N_1477,In_488,In_281);
xnor U1478 (N_1478,In_662,In_422);
nor U1479 (N_1479,In_22,In_686);
and U1480 (N_1480,In_446,In_241);
nand U1481 (N_1481,In_404,In_745);
or U1482 (N_1482,In_61,In_635);
or U1483 (N_1483,In_414,In_331);
nor U1484 (N_1484,In_725,In_403);
and U1485 (N_1485,In_97,In_297);
and U1486 (N_1486,In_494,In_206);
or U1487 (N_1487,In_723,In_181);
nand U1488 (N_1488,In_662,In_469);
and U1489 (N_1489,In_291,In_292);
nor U1490 (N_1490,In_741,In_447);
nand U1491 (N_1491,In_524,In_151);
and U1492 (N_1492,In_718,In_142);
nor U1493 (N_1493,In_247,In_240);
or U1494 (N_1494,In_590,In_638);
nor U1495 (N_1495,In_224,In_155);
and U1496 (N_1496,In_174,In_290);
and U1497 (N_1497,In_245,In_569);
or U1498 (N_1498,In_15,In_658);
nor U1499 (N_1499,In_574,In_733);
nand U1500 (N_1500,In_452,In_736);
nand U1501 (N_1501,In_450,In_592);
nor U1502 (N_1502,In_53,In_585);
or U1503 (N_1503,In_527,In_199);
nand U1504 (N_1504,In_72,In_593);
nand U1505 (N_1505,In_313,In_418);
and U1506 (N_1506,In_327,In_167);
or U1507 (N_1507,In_433,In_614);
and U1508 (N_1508,In_727,In_313);
xor U1509 (N_1509,In_310,In_580);
nor U1510 (N_1510,In_306,In_223);
nand U1511 (N_1511,In_551,In_745);
nand U1512 (N_1512,In_242,In_661);
and U1513 (N_1513,In_734,In_340);
or U1514 (N_1514,In_474,In_238);
xor U1515 (N_1515,In_293,In_680);
and U1516 (N_1516,In_501,In_434);
nor U1517 (N_1517,In_202,In_728);
or U1518 (N_1518,In_253,In_632);
and U1519 (N_1519,In_545,In_705);
or U1520 (N_1520,In_542,In_271);
nand U1521 (N_1521,In_620,In_68);
xor U1522 (N_1522,In_282,In_268);
and U1523 (N_1523,In_658,In_89);
xor U1524 (N_1524,In_314,In_370);
nand U1525 (N_1525,In_125,In_732);
or U1526 (N_1526,In_357,In_89);
or U1527 (N_1527,In_531,In_737);
xnor U1528 (N_1528,In_340,In_12);
nor U1529 (N_1529,In_401,In_713);
nand U1530 (N_1530,In_34,In_275);
or U1531 (N_1531,In_592,In_217);
nor U1532 (N_1532,In_34,In_679);
and U1533 (N_1533,In_470,In_425);
nor U1534 (N_1534,In_667,In_499);
xnor U1535 (N_1535,In_487,In_301);
or U1536 (N_1536,In_749,In_330);
nand U1537 (N_1537,In_140,In_630);
xor U1538 (N_1538,In_631,In_326);
and U1539 (N_1539,In_75,In_80);
or U1540 (N_1540,In_632,In_635);
and U1541 (N_1541,In_601,In_168);
nor U1542 (N_1542,In_465,In_534);
and U1543 (N_1543,In_711,In_107);
and U1544 (N_1544,In_440,In_237);
and U1545 (N_1545,In_728,In_132);
nor U1546 (N_1546,In_621,In_73);
nor U1547 (N_1547,In_391,In_62);
and U1548 (N_1548,In_218,In_187);
and U1549 (N_1549,In_639,In_88);
or U1550 (N_1550,In_580,In_261);
xnor U1551 (N_1551,In_128,In_726);
nand U1552 (N_1552,In_473,In_347);
and U1553 (N_1553,In_699,In_67);
nor U1554 (N_1554,In_130,In_463);
nor U1555 (N_1555,In_572,In_566);
xnor U1556 (N_1556,In_148,In_240);
nand U1557 (N_1557,In_719,In_449);
and U1558 (N_1558,In_300,In_215);
or U1559 (N_1559,In_736,In_686);
and U1560 (N_1560,In_253,In_275);
and U1561 (N_1561,In_542,In_83);
xor U1562 (N_1562,In_602,In_202);
and U1563 (N_1563,In_603,In_152);
nor U1564 (N_1564,In_646,In_587);
and U1565 (N_1565,In_539,In_331);
or U1566 (N_1566,In_106,In_52);
or U1567 (N_1567,In_443,In_202);
and U1568 (N_1568,In_230,In_519);
nand U1569 (N_1569,In_550,In_610);
nand U1570 (N_1570,In_681,In_242);
or U1571 (N_1571,In_225,In_294);
xor U1572 (N_1572,In_199,In_201);
nor U1573 (N_1573,In_563,In_672);
nor U1574 (N_1574,In_199,In_279);
xor U1575 (N_1575,In_91,In_624);
and U1576 (N_1576,In_24,In_492);
nand U1577 (N_1577,In_503,In_323);
and U1578 (N_1578,In_157,In_493);
nand U1579 (N_1579,In_435,In_659);
and U1580 (N_1580,In_609,In_219);
or U1581 (N_1581,In_690,In_174);
or U1582 (N_1582,In_151,In_505);
nor U1583 (N_1583,In_297,In_190);
and U1584 (N_1584,In_390,In_681);
or U1585 (N_1585,In_664,In_38);
or U1586 (N_1586,In_444,In_204);
or U1587 (N_1587,In_670,In_5);
nor U1588 (N_1588,In_742,In_551);
xnor U1589 (N_1589,In_593,In_504);
and U1590 (N_1590,In_107,In_2);
or U1591 (N_1591,In_310,In_617);
xor U1592 (N_1592,In_421,In_345);
or U1593 (N_1593,In_541,In_618);
or U1594 (N_1594,In_227,In_338);
and U1595 (N_1595,In_147,In_286);
nand U1596 (N_1596,In_207,In_74);
or U1597 (N_1597,In_92,In_667);
nand U1598 (N_1598,In_398,In_446);
nand U1599 (N_1599,In_448,In_656);
xnor U1600 (N_1600,In_536,In_164);
and U1601 (N_1601,In_429,In_85);
nand U1602 (N_1602,In_535,In_373);
nand U1603 (N_1603,In_657,In_3);
or U1604 (N_1604,In_423,In_527);
and U1605 (N_1605,In_698,In_195);
xnor U1606 (N_1606,In_682,In_556);
or U1607 (N_1607,In_78,In_558);
nor U1608 (N_1608,In_549,In_383);
nor U1609 (N_1609,In_185,In_687);
nand U1610 (N_1610,In_277,In_95);
and U1611 (N_1611,In_335,In_576);
nor U1612 (N_1612,In_208,In_629);
and U1613 (N_1613,In_654,In_553);
and U1614 (N_1614,In_51,In_274);
and U1615 (N_1615,In_97,In_595);
nor U1616 (N_1616,In_33,In_472);
or U1617 (N_1617,In_450,In_23);
xnor U1618 (N_1618,In_398,In_659);
nor U1619 (N_1619,In_580,In_491);
nor U1620 (N_1620,In_112,In_390);
or U1621 (N_1621,In_382,In_399);
nor U1622 (N_1622,In_41,In_697);
nand U1623 (N_1623,In_499,In_582);
or U1624 (N_1624,In_81,In_552);
nand U1625 (N_1625,In_147,In_221);
nor U1626 (N_1626,In_739,In_181);
nor U1627 (N_1627,In_374,In_81);
or U1628 (N_1628,In_452,In_525);
and U1629 (N_1629,In_141,In_555);
or U1630 (N_1630,In_116,In_682);
nor U1631 (N_1631,In_646,In_286);
or U1632 (N_1632,In_405,In_328);
or U1633 (N_1633,In_32,In_551);
nor U1634 (N_1634,In_139,In_438);
nor U1635 (N_1635,In_434,In_672);
nand U1636 (N_1636,In_543,In_575);
nand U1637 (N_1637,In_538,In_11);
or U1638 (N_1638,In_529,In_470);
nor U1639 (N_1639,In_339,In_70);
and U1640 (N_1640,In_699,In_169);
and U1641 (N_1641,In_403,In_563);
nor U1642 (N_1642,In_151,In_542);
and U1643 (N_1643,In_482,In_170);
nand U1644 (N_1644,In_342,In_155);
nand U1645 (N_1645,In_97,In_717);
or U1646 (N_1646,In_9,In_734);
nor U1647 (N_1647,In_81,In_747);
and U1648 (N_1648,In_639,In_47);
nor U1649 (N_1649,In_632,In_704);
and U1650 (N_1650,In_432,In_88);
and U1651 (N_1651,In_365,In_136);
or U1652 (N_1652,In_328,In_516);
and U1653 (N_1653,In_523,In_351);
and U1654 (N_1654,In_437,In_136);
nand U1655 (N_1655,In_324,In_156);
or U1656 (N_1656,In_177,In_114);
nor U1657 (N_1657,In_177,In_389);
or U1658 (N_1658,In_693,In_488);
nand U1659 (N_1659,In_286,In_19);
or U1660 (N_1660,In_223,In_58);
or U1661 (N_1661,In_156,In_695);
nor U1662 (N_1662,In_698,In_353);
and U1663 (N_1663,In_78,In_181);
nor U1664 (N_1664,In_420,In_639);
nand U1665 (N_1665,In_623,In_437);
nor U1666 (N_1666,In_538,In_41);
nor U1667 (N_1667,In_742,In_171);
or U1668 (N_1668,In_385,In_76);
and U1669 (N_1669,In_681,In_186);
or U1670 (N_1670,In_6,In_289);
nand U1671 (N_1671,In_163,In_421);
nand U1672 (N_1672,In_557,In_215);
and U1673 (N_1673,In_431,In_116);
and U1674 (N_1674,In_11,In_676);
nand U1675 (N_1675,In_683,In_674);
nor U1676 (N_1676,In_411,In_524);
or U1677 (N_1677,In_697,In_515);
or U1678 (N_1678,In_44,In_127);
and U1679 (N_1679,In_418,In_147);
nor U1680 (N_1680,In_496,In_301);
or U1681 (N_1681,In_738,In_168);
nor U1682 (N_1682,In_16,In_278);
nor U1683 (N_1683,In_676,In_223);
or U1684 (N_1684,In_501,In_691);
and U1685 (N_1685,In_10,In_241);
nor U1686 (N_1686,In_343,In_488);
or U1687 (N_1687,In_482,In_538);
nor U1688 (N_1688,In_124,In_511);
nand U1689 (N_1689,In_100,In_537);
xor U1690 (N_1690,In_548,In_483);
nor U1691 (N_1691,In_250,In_415);
or U1692 (N_1692,In_472,In_497);
nor U1693 (N_1693,In_317,In_162);
or U1694 (N_1694,In_636,In_526);
and U1695 (N_1695,In_715,In_460);
and U1696 (N_1696,In_124,In_6);
or U1697 (N_1697,In_482,In_650);
nor U1698 (N_1698,In_563,In_203);
and U1699 (N_1699,In_659,In_281);
nand U1700 (N_1700,In_465,In_165);
nor U1701 (N_1701,In_598,In_404);
or U1702 (N_1702,In_745,In_632);
and U1703 (N_1703,In_351,In_163);
nor U1704 (N_1704,In_52,In_186);
and U1705 (N_1705,In_485,In_606);
or U1706 (N_1706,In_308,In_413);
nand U1707 (N_1707,In_46,In_105);
or U1708 (N_1708,In_312,In_174);
nand U1709 (N_1709,In_359,In_49);
and U1710 (N_1710,In_725,In_166);
nor U1711 (N_1711,In_170,In_428);
xnor U1712 (N_1712,In_342,In_106);
nor U1713 (N_1713,In_158,In_510);
or U1714 (N_1714,In_471,In_283);
nand U1715 (N_1715,In_373,In_80);
nor U1716 (N_1716,In_552,In_23);
and U1717 (N_1717,In_94,In_389);
nand U1718 (N_1718,In_33,In_77);
nor U1719 (N_1719,In_471,In_517);
and U1720 (N_1720,In_90,In_568);
xnor U1721 (N_1721,In_196,In_7);
or U1722 (N_1722,In_226,In_478);
or U1723 (N_1723,In_389,In_447);
or U1724 (N_1724,In_674,In_202);
or U1725 (N_1725,In_654,In_310);
and U1726 (N_1726,In_553,In_369);
nor U1727 (N_1727,In_89,In_86);
and U1728 (N_1728,In_538,In_152);
xnor U1729 (N_1729,In_193,In_231);
nor U1730 (N_1730,In_153,In_47);
nor U1731 (N_1731,In_31,In_505);
and U1732 (N_1732,In_181,In_660);
or U1733 (N_1733,In_138,In_312);
and U1734 (N_1734,In_501,In_313);
or U1735 (N_1735,In_30,In_383);
and U1736 (N_1736,In_471,In_484);
nor U1737 (N_1737,In_452,In_585);
nor U1738 (N_1738,In_26,In_640);
nand U1739 (N_1739,In_78,In_408);
nor U1740 (N_1740,In_337,In_26);
or U1741 (N_1741,In_114,In_369);
or U1742 (N_1742,In_511,In_408);
and U1743 (N_1743,In_132,In_199);
xnor U1744 (N_1744,In_110,In_127);
nor U1745 (N_1745,In_272,In_193);
and U1746 (N_1746,In_714,In_358);
nor U1747 (N_1747,In_726,In_436);
nor U1748 (N_1748,In_241,In_320);
xor U1749 (N_1749,In_299,In_396);
or U1750 (N_1750,In_296,In_203);
nand U1751 (N_1751,In_31,In_627);
and U1752 (N_1752,In_342,In_373);
nand U1753 (N_1753,In_270,In_134);
or U1754 (N_1754,In_727,In_425);
or U1755 (N_1755,In_258,In_322);
nand U1756 (N_1756,In_663,In_232);
nor U1757 (N_1757,In_708,In_0);
nor U1758 (N_1758,In_511,In_366);
and U1759 (N_1759,In_427,In_35);
nor U1760 (N_1760,In_372,In_147);
nor U1761 (N_1761,In_141,In_228);
and U1762 (N_1762,In_669,In_569);
nor U1763 (N_1763,In_632,In_42);
and U1764 (N_1764,In_372,In_700);
nand U1765 (N_1765,In_67,In_401);
nand U1766 (N_1766,In_363,In_132);
nand U1767 (N_1767,In_590,In_505);
or U1768 (N_1768,In_202,In_561);
xnor U1769 (N_1769,In_647,In_328);
or U1770 (N_1770,In_458,In_437);
nand U1771 (N_1771,In_194,In_17);
and U1772 (N_1772,In_123,In_5);
or U1773 (N_1773,In_558,In_435);
or U1774 (N_1774,In_728,In_245);
nor U1775 (N_1775,In_521,In_466);
nand U1776 (N_1776,In_548,In_629);
nand U1777 (N_1777,In_232,In_185);
nand U1778 (N_1778,In_640,In_34);
nand U1779 (N_1779,In_53,In_712);
nor U1780 (N_1780,In_190,In_624);
or U1781 (N_1781,In_661,In_503);
nand U1782 (N_1782,In_556,In_226);
nor U1783 (N_1783,In_51,In_396);
nand U1784 (N_1784,In_373,In_418);
xnor U1785 (N_1785,In_151,In_263);
nor U1786 (N_1786,In_539,In_438);
nor U1787 (N_1787,In_749,In_706);
or U1788 (N_1788,In_625,In_593);
nand U1789 (N_1789,In_453,In_51);
xnor U1790 (N_1790,In_374,In_637);
nor U1791 (N_1791,In_141,In_303);
nand U1792 (N_1792,In_394,In_578);
or U1793 (N_1793,In_4,In_743);
and U1794 (N_1794,In_300,In_630);
and U1795 (N_1795,In_724,In_682);
and U1796 (N_1796,In_107,In_458);
xnor U1797 (N_1797,In_672,In_550);
and U1798 (N_1798,In_550,In_463);
or U1799 (N_1799,In_690,In_645);
and U1800 (N_1800,In_113,In_174);
nor U1801 (N_1801,In_253,In_605);
xor U1802 (N_1802,In_702,In_88);
nand U1803 (N_1803,In_244,In_578);
nor U1804 (N_1804,In_307,In_512);
nand U1805 (N_1805,In_109,In_736);
nor U1806 (N_1806,In_210,In_632);
and U1807 (N_1807,In_595,In_433);
and U1808 (N_1808,In_467,In_338);
or U1809 (N_1809,In_521,In_456);
nor U1810 (N_1810,In_541,In_691);
nand U1811 (N_1811,In_205,In_680);
xnor U1812 (N_1812,In_708,In_252);
or U1813 (N_1813,In_261,In_598);
or U1814 (N_1814,In_649,In_440);
nand U1815 (N_1815,In_364,In_664);
and U1816 (N_1816,In_450,In_630);
nor U1817 (N_1817,In_416,In_541);
and U1818 (N_1818,In_386,In_521);
nand U1819 (N_1819,In_403,In_676);
nor U1820 (N_1820,In_118,In_344);
nand U1821 (N_1821,In_279,In_709);
xor U1822 (N_1822,In_401,In_614);
nand U1823 (N_1823,In_604,In_242);
or U1824 (N_1824,In_410,In_447);
nand U1825 (N_1825,In_389,In_195);
nand U1826 (N_1826,In_260,In_184);
nor U1827 (N_1827,In_43,In_208);
or U1828 (N_1828,In_161,In_551);
nand U1829 (N_1829,In_150,In_720);
nand U1830 (N_1830,In_469,In_21);
or U1831 (N_1831,In_244,In_551);
nand U1832 (N_1832,In_76,In_201);
nand U1833 (N_1833,In_304,In_466);
or U1834 (N_1834,In_162,In_567);
nand U1835 (N_1835,In_101,In_362);
nand U1836 (N_1836,In_448,In_46);
and U1837 (N_1837,In_347,In_475);
nand U1838 (N_1838,In_602,In_9);
nand U1839 (N_1839,In_413,In_108);
nor U1840 (N_1840,In_491,In_331);
xor U1841 (N_1841,In_724,In_699);
and U1842 (N_1842,In_180,In_581);
or U1843 (N_1843,In_319,In_286);
or U1844 (N_1844,In_369,In_140);
nor U1845 (N_1845,In_360,In_736);
nor U1846 (N_1846,In_236,In_697);
and U1847 (N_1847,In_609,In_645);
xnor U1848 (N_1848,In_507,In_59);
nor U1849 (N_1849,In_630,In_575);
or U1850 (N_1850,In_266,In_264);
or U1851 (N_1851,In_404,In_5);
xnor U1852 (N_1852,In_220,In_300);
or U1853 (N_1853,In_538,In_725);
and U1854 (N_1854,In_743,In_251);
and U1855 (N_1855,In_417,In_541);
nor U1856 (N_1856,In_571,In_12);
or U1857 (N_1857,In_407,In_728);
nor U1858 (N_1858,In_128,In_444);
or U1859 (N_1859,In_372,In_341);
or U1860 (N_1860,In_667,In_140);
and U1861 (N_1861,In_124,In_439);
and U1862 (N_1862,In_118,In_519);
or U1863 (N_1863,In_305,In_99);
nor U1864 (N_1864,In_168,In_749);
or U1865 (N_1865,In_117,In_294);
nand U1866 (N_1866,In_721,In_596);
or U1867 (N_1867,In_663,In_694);
nand U1868 (N_1868,In_192,In_501);
nor U1869 (N_1869,In_314,In_340);
nand U1870 (N_1870,In_84,In_422);
nand U1871 (N_1871,In_426,In_436);
nand U1872 (N_1872,In_710,In_384);
nand U1873 (N_1873,In_61,In_201);
or U1874 (N_1874,In_652,In_62);
xor U1875 (N_1875,In_222,In_239);
and U1876 (N_1876,In_290,In_74);
xor U1877 (N_1877,In_315,In_37);
or U1878 (N_1878,In_537,In_536);
nand U1879 (N_1879,In_728,In_724);
and U1880 (N_1880,In_389,In_358);
xnor U1881 (N_1881,In_389,In_357);
or U1882 (N_1882,In_453,In_670);
or U1883 (N_1883,In_449,In_616);
or U1884 (N_1884,In_477,In_321);
and U1885 (N_1885,In_520,In_147);
nor U1886 (N_1886,In_179,In_236);
nor U1887 (N_1887,In_597,In_749);
nor U1888 (N_1888,In_336,In_333);
or U1889 (N_1889,In_394,In_539);
or U1890 (N_1890,In_736,In_668);
nor U1891 (N_1891,In_75,In_705);
nor U1892 (N_1892,In_493,In_100);
xnor U1893 (N_1893,In_222,In_640);
nor U1894 (N_1894,In_519,In_441);
xnor U1895 (N_1895,In_262,In_681);
nor U1896 (N_1896,In_220,In_37);
nor U1897 (N_1897,In_387,In_626);
nand U1898 (N_1898,In_686,In_249);
nor U1899 (N_1899,In_437,In_543);
nand U1900 (N_1900,In_334,In_503);
and U1901 (N_1901,In_110,In_73);
and U1902 (N_1902,In_615,In_650);
nor U1903 (N_1903,In_184,In_204);
xnor U1904 (N_1904,In_733,In_617);
nor U1905 (N_1905,In_373,In_596);
nor U1906 (N_1906,In_5,In_685);
xnor U1907 (N_1907,In_145,In_157);
nand U1908 (N_1908,In_552,In_580);
or U1909 (N_1909,In_667,In_484);
nor U1910 (N_1910,In_334,In_530);
and U1911 (N_1911,In_141,In_601);
and U1912 (N_1912,In_387,In_625);
and U1913 (N_1913,In_345,In_381);
nand U1914 (N_1914,In_167,In_40);
or U1915 (N_1915,In_212,In_73);
or U1916 (N_1916,In_6,In_254);
and U1917 (N_1917,In_443,In_568);
xor U1918 (N_1918,In_297,In_381);
and U1919 (N_1919,In_480,In_177);
or U1920 (N_1920,In_377,In_356);
nand U1921 (N_1921,In_608,In_371);
nand U1922 (N_1922,In_359,In_440);
nand U1923 (N_1923,In_390,In_297);
nor U1924 (N_1924,In_654,In_188);
nor U1925 (N_1925,In_169,In_326);
nand U1926 (N_1926,In_217,In_471);
or U1927 (N_1927,In_736,In_93);
and U1928 (N_1928,In_16,In_47);
nor U1929 (N_1929,In_72,In_422);
nand U1930 (N_1930,In_28,In_339);
xor U1931 (N_1931,In_76,In_255);
nor U1932 (N_1932,In_655,In_443);
and U1933 (N_1933,In_10,In_579);
and U1934 (N_1934,In_627,In_477);
or U1935 (N_1935,In_232,In_251);
or U1936 (N_1936,In_43,In_620);
and U1937 (N_1937,In_105,In_625);
and U1938 (N_1938,In_28,In_555);
nand U1939 (N_1939,In_214,In_374);
or U1940 (N_1940,In_574,In_419);
nand U1941 (N_1941,In_584,In_683);
and U1942 (N_1942,In_562,In_57);
xnor U1943 (N_1943,In_702,In_743);
and U1944 (N_1944,In_655,In_230);
and U1945 (N_1945,In_586,In_697);
nor U1946 (N_1946,In_200,In_294);
or U1947 (N_1947,In_410,In_161);
nand U1948 (N_1948,In_66,In_391);
or U1949 (N_1949,In_414,In_699);
and U1950 (N_1950,In_426,In_609);
nor U1951 (N_1951,In_422,In_223);
nor U1952 (N_1952,In_698,In_663);
nand U1953 (N_1953,In_243,In_387);
nand U1954 (N_1954,In_143,In_553);
and U1955 (N_1955,In_48,In_151);
and U1956 (N_1956,In_299,In_291);
nand U1957 (N_1957,In_154,In_659);
or U1958 (N_1958,In_692,In_37);
and U1959 (N_1959,In_678,In_278);
nor U1960 (N_1960,In_580,In_211);
xor U1961 (N_1961,In_351,In_660);
and U1962 (N_1962,In_26,In_421);
nand U1963 (N_1963,In_89,In_450);
nor U1964 (N_1964,In_391,In_466);
or U1965 (N_1965,In_371,In_219);
nor U1966 (N_1966,In_296,In_353);
nor U1967 (N_1967,In_650,In_230);
nand U1968 (N_1968,In_495,In_317);
nand U1969 (N_1969,In_746,In_500);
or U1970 (N_1970,In_376,In_534);
nand U1971 (N_1971,In_150,In_152);
xnor U1972 (N_1972,In_104,In_358);
and U1973 (N_1973,In_192,In_378);
or U1974 (N_1974,In_317,In_550);
and U1975 (N_1975,In_47,In_109);
or U1976 (N_1976,In_366,In_29);
or U1977 (N_1977,In_182,In_279);
and U1978 (N_1978,In_15,In_452);
or U1979 (N_1979,In_466,In_375);
or U1980 (N_1980,In_286,In_641);
nand U1981 (N_1981,In_543,In_628);
or U1982 (N_1982,In_428,In_713);
nor U1983 (N_1983,In_513,In_149);
nand U1984 (N_1984,In_500,In_190);
and U1985 (N_1985,In_244,In_289);
and U1986 (N_1986,In_559,In_715);
and U1987 (N_1987,In_642,In_509);
nand U1988 (N_1988,In_59,In_395);
xor U1989 (N_1989,In_132,In_146);
and U1990 (N_1990,In_65,In_426);
and U1991 (N_1991,In_643,In_437);
xor U1992 (N_1992,In_681,In_460);
or U1993 (N_1993,In_190,In_315);
or U1994 (N_1994,In_735,In_665);
nor U1995 (N_1995,In_164,In_65);
and U1996 (N_1996,In_528,In_628);
or U1997 (N_1997,In_42,In_154);
or U1998 (N_1998,In_572,In_608);
or U1999 (N_1999,In_316,In_404);
nand U2000 (N_2000,In_417,In_384);
or U2001 (N_2001,In_615,In_675);
nor U2002 (N_2002,In_490,In_656);
or U2003 (N_2003,In_441,In_251);
and U2004 (N_2004,In_368,In_309);
nand U2005 (N_2005,In_703,In_464);
and U2006 (N_2006,In_619,In_634);
nor U2007 (N_2007,In_378,In_118);
xor U2008 (N_2008,In_36,In_253);
and U2009 (N_2009,In_691,In_510);
or U2010 (N_2010,In_178,In_491);
nand U2011 (N_2011,In_715,In_682);
nand U2012 (N_2012,In_254,In_430);
nand U2013 (N_2013,In_306,In_131);
xor U2014 (N_2014,In_268,In_336);
and U2015 (N_2015,In_2,In_411);
xor U2016 (N_2016,In_585,In_128);
or U2017 (N_2017,In_647,In_441);
nand U2018 (N_2018,In_318,In_138);
or U2019 (N_2019,In_333,In_472);
xnor U2020 (N_2020,In_663,In_145);
xnor U2021 (N_2021,In_466,In_332);
nand U2022 (N_2022,In_75,In_697);
and U2023 (N_2023,In_161,In_486);
nand U2024 (N_2024,In_617,In_234);
nand U2025 (N_2025,In_34,In_41);
nand U2026 (N_2026,In_387,In_623);
and U2027 (N_2027,In_47,In_648);
and U2028 (N_2028,In_134,In_647);
nor U2029 (N_2029,In_330,In_613);
nand U2030 (N_2030,In_534,In_443);
and U2031 (N_2031,In_302,In_677);
nor U2032 (N_2032,In_674,In_74);
and U2033 (N_2033,In_99,In_241);
and U2034 (N_2034,In_4,In_14);
nand U2035 (N_2035,In_582,In_40);
and U2036 (N_2036,In_172,In_479);
and U2037 (N_2037,In_60,In_295);
nor U2038 (N_2038,In_652,In_563);
and U2039 (N_2039,In_393,In_669);
nand U2040 (N_2040,In_473,In_247);
nor U2041 (N_2041,In_384,In_88);
and U2042 (N_2042,In_661,In_365);
nand U2043 (N_2043,In_242,In_533);
nor U2044 (N_2044,In_136,In_416);
or U2045 (N_2045,In_580,In_441);
and U2046 (N_2046,In_210,In_99);
or U2047 (N_2047,In_210,In_406);
nor U2048 (N_2048,In_429,In_30);
xnor U2049 (N_2049,In_484,In_339);
xnor U2050 (N_2050,In_264,In_442);
or U2051 (N_2051,In_588,In_536);
nand U2052 (N_2052,In_354,In_47);
and U2053 (N_2053,In_408,In_108);
xnor U2054 (N_2054,In_99,In_344);
nand U2055 (N_2055,In_123,In_335);
nand U2056 (N_2056,In_393,In_438);
or U2057 (N_2057,In_272,In_125);
nor U2058 (N_2058,In_441,In_423);
or U2059 (N_2059,In_493,In_80);
xnor U2060 (N_2060,In_421,In_557);
nand U2061 (N_2061,In_429,In_136);
nand U2062 (N_2062,In_702,In_310);
and U2063 (N_2063,In_68,In_186);
nor U2064 (N_2064,In_187,In_533);
or U2065 (N_2065,In_118,In_36);
nor U2066 (N_2066,In_616,In_562);
xor U2067 (N_2067,In_211,In_328);
nor U2068 (N_2068,In_126,In_724);
xnor U2069 (N_2069,In_684,In_44);
or U2070 (N_2070,In_276,In_19);
xnor U2071 (N_2071,In_26,In_297);
nand U2072 (N_2072,In_537,In_498);
or U2073 (N_2073,In_70,In_85);
or U2074 (N_2074,In_679,In_119);
xor U2075 (N_2075,In_415,In_587);
nor U2076 (N_2076,In_363,In_523);
nand U2077 (N_2077,In_58,In_316);
and U2078 (N_2078,In_460,In_103);
nor U2079 (N_2079,In_398,In_639);
or U2080 (N_2080,In_635,In_109);
nor U2081 (N_2081,In_546,In_430);
or U2082 (N_2082,In_613,In_119);
or U2083 (N_2083,In_625,In_70);
nor U2084 (N_2084,In_728,In_738);
nand U2085 (N_2085,In_12,In_48);
nand U2086 (N_2086,In_337,In_220);
and U2087 (N_2087,In_419,In_146);
nor U2088 (N_2088,In_691,In_722);
nand U2089 (N_2089,In_467,In_632);
nand U2090 (N_2090,In_82,In_187);
or U2091 (N_2091,In_431,In_34);
or U2092 (N_2092,In_704,In_266);
nand U2093 (N_2093,In_695,In_623);
and U2094 (N_2094,In_177,In_472);
nand U2095 (N_2095,In_304,In_396);
or U2096 (N_2096,In_475,In_183);
and U2097 (N_2097,In_540,In_183);
nor U2098 (N_2098,In_304,In_601);
nor U2099 (N_2099,In_482,In_52);
and U2100 (N_2100,In_454,In_407);
and U2101 (N_2101,In_26,In_71);
xor U2102 (N_2102,In_446,In_250);
nand U2103 (N_2103,In_110,In_281);
and U2104 (N_2104,In_220,In_608);
or U2105 (N_2105,In_367,In_203);
nand U2106 (N_2106,In_252,In_41);
or U2107 (N_2107,In_396,In_390);
or U2108 (N_2108,In_687,In_647);
and U2109 (N_2109,In_644,In_268);
or U2110 (N_2110,In_727,In_41);
or U2111 (N_2111,In_588,In_126);
nor U2112 (N_2112,In_597,In_540);
nor U2113 (N_2113,In_515,In_294);
xnor U2114 (N_2114,In_133,In_289);
nor U2115 (N_2115,In_248,In_469);
nand U2116 (N_2116,In_233,In_564);
or U2117 (N_2117,In_197,In_683);
nand U2118 (N_2118,In_614,In_508);
or U2119 (N_2119,In_38,In_521);
nor U2120 (N_2120,In_565,In_155);
and U2121 (N_2121,In_651,In_145);
nand U2122 (N_2122,In_49,In_646);
and U2123 (N_2123,In_185,In_34);
nor U2124 (N_2124,In_694,In_717);
nand U2125 (N_2125,In_640,In_105);
or U2126 (N_2126,In_346,In_162);
xnor U2127 (N_2127,In_585,In_28);
nand U2128 (N_2128,In_594,In_16);
nand U2129 (N_2129,In_239,In_340);
and U2130 (N_2130,In_646,In_107);
nand U2131 (N_2131,In_469,In_264);
nor U2132 (N_2132,In_106,In_559);
and U2133 (N_2133,In_571,In_177);
or U2134 (N_2134,In_39,In_695);
nor U2135 (N_2135,In_616,In_316);
or U2136 (N_2136,In_491,In_448);
nor U2137 (N_2137,In_394,In_353);
or U2138 (N_2138,In_388,In_45);
nand U2139 (N_2139,In_7,In_567);
and U2140 (N_2140,In_686,In_359);
and U2141 (N_2141,In_64,In_733);
nor U2142 (N_2142,In_474,In_152);
nor U2143 (N_2143,In_124,In_163);
and U2144 (N_2144,In_481,In_361);
nor U2145 (N_2145,In_43,In_561);
or U2146 (N_2146,In_279,In_366);
nor U2147 (N_2147,In_640,In_710);
and U2148 (N_2148,In_655,In_209);
nand U2149 (N_2149,In_667,In_302);
xor U2150 (N_2150,In_77,In_61);
nor U2151 (N_2151,In_199,In_631);
and U2152 (N_2152,In_330,In_92);
or U2153 (N_2153,In_9,In_541);
or U2154 (N_2154,In_515,In_51);
xnor U2155 (N_2155,In_602,In_516);
nor U2156 (N_2156,In_629,In_408);
nand U2157 (N_2157,In_625,In_499);
or U2158 (N_2158,In_108,In_2);
or U2159 (N_2159,In_181,In_678);
nor U2160 (N_2160,In_318,In_413);
and U2161 (N_2161,In_591,In_165);
nor U2162 (N_2162,In_369,In_200);
nand U2163 (N_2163,In_613,In_57);
or U2164 (N_2164,In_612,In_215);
nand U2165 (N_2165,In_639,In_424);
nor U2166 (N_2166,In_460,In_381);
nand U2167 (N_2167,In_419,In_616);
nor U2168 (N_2168,In_656,In_731);
or U2169 (N_2169,In_63,In_172);
or U2170 (N_2170,In_48,In_621);
nand U2171 (N_2171,In_512,In_536);
xnor U2172 (N_2172,In_475,In_663);
nor U2173 (N_2173,In_398,In_406);
and U2174 (N_2174,In_358,In_575);
or U2175 (N_2175,In_491,In_308);
or U2176 (N_2176,In_506,In_234);
nor U2177 (N_2177,In_358,In_98);
or U2178 (N_2178,In_132,In_59);
nor U2179 (N_2179,In_483,In_605);
and U2180 (N_2180,In_85,In_376);
nand U2181 (N_2181,In_458,In_97);
and U2182 (N_2182,In_625,In_202);
and U2183 (N_2183,In_20,In_129);
nand U2184 (N_2184,In_8,In_634);
and U2185 (N_2185,In_84,In_85);
nand U2186 (N_2186,In_227,In_634);
nand U2187 (N_2187,In_603,In_22);
nor U2188 (N_2188,In_692,In_336);
nand U2189 (N_2189,In_602,In_232);
nor U2190 (N_2190,In_265,In_570);
and U2191 (N_2191,In_153,In_388);
or U2192 (N_2192,In_8,In_340);
nand U2193 (N_2193,In_99,In_283);
or U2194 (N_2194,In_118,In_237);
and U2195 (N_2195,In_228,In_327);
and U2196 (N_2196,In_309,In_444);
nand U2197 (N_2197,In_552,In_729);
nor U2198 (N_2198,In_262,In_731);
and U2199 (N_2199,In_356,In_655);
nor U2200 (N_2200,In_487,In_139);
nor U2201 (N_2201,In_170,In_36);
nand U2202 (N_2202,In_77,In_54);
nor U2203 (N_2203,In_437,In_380);
and U2204 (N_2204,In_304,In_258);
nand U2205 (N_2205,In_729,In_589);
nor U2206 (N_2206,In_502,In_614);
nand U2207 (N_2207,In_444,In_324);
and U2208 (N_2208,In_507,In_64);
xor U2209 (N_2209,In_461,In_10);
nor U2210 (N_2210,In_48,In_697);
nand U2211 (N_2211,In_408,In_271);
or U2212 (N_2212,In_282,In_257);
nor U2213 (N_2213,In_556,In_729);
and U2214 (N_2214,In_309,In_646);
nor U2215 (N_2215,In_617,In_343);
or U2216 (N_2216,In_584,In_506);
nor U2217 (N_2217,In_255,In_437);
or U2218 (N_2218,In_24,In_16);
nand U2219 (N_2219,In_372,In_353);
and U2220 (N_2220,In_323,In_535);
nand U2221 (N_2221,In_56,In_573);
nand U2222 (N_2222,In_376,In_140);
nor U2223 (N_2223,In_286,In_521);
xnor U2224 (N_2224,In_292,In_621);
or U2225 (N_2225,In_733,In_262);
nand U2226 (N_2226,In_204,In_268);
and U2227 (N_2227,In_471,In_399);
nand U2228 (N_2228,In_104,In_147);
xnor U2229 (N_2229,In_522,In_427);
or U2230 (N_2230,In_558,In_110);
nor U2231 (N_2231,In_388,In_537);
xnor U2232 (N_2232,In_301,In_700);
nand U2233 (N_2233,In_211,In_708);
nor U2234 (N_2234,In_616,In_262);
xnor U2235 (N_2235,In_61,In_740);
and U2236 (N_2236,In_676,In_353);
or U2237 (N_2237,In_472,In_288);
or U2238 (N_2238,In_286,In_418);
and U2239 (N_2239,In_383,In_526);
and U2240 (N_2240,In_377,In_81);
nand U2241 (N_2241,In_142,In_199);
nor U2242 (N_2242,In_658,In_526);
nand U2243 (N_2243,In_65,In_570);
and U2244 (N_2244,In_701,In_57);
nor U2245 (N_2245,In_619,In_529);
or U2246 (N_2246,In_374,In_728);
or U2247 (N_2247,In_7,In_224);
and U2248 (N_2248,In_216,In_207);
and U2249 (N_2249,In_261,In_185);
nand U2250 (N_2250,In_477,In_219);
or U2251 (N_2251,In_70,In_172);
and U2252 (N_2252,In_42,In_329);
xor U2253 (N_2253,In_132,In_163);
xnor U2254 (N_2254,In_57,In_644);
or U2255 (N_2255,In_354,In_299);
nand U2256 (N_2256,In_500,In_596);
and U2257 (N_2257,In_516,In_506);
and U2258 (N_2258,In_629,In_67);
or U2259 (N_2259,In_526,In_94);
and U2260 (N_2260,In_284,In_274);
xnor U2261 (N_2261,In_12,In_362);
or U2262 (N_2262,In_77,In_599);
and U2263 (N_2263,In_259,In_536);
nand U2264 (N_2264,In_710,In_374);
and U2265 (N_2265,In_456,In_192);
nor U2266 (N_2266,In_354,In_386);
nand U2267 (N_2267,In_183,In_478);
nor U2268 (N_2268,In_73,In_459);
or U2269 (N_2269,In_178,In_169);
or U2270 (N_2270,In_334,In_12);
nor U2271 (N_2271,In_166,In_523);
nand U2272 (N_2272,In_743,In_85);
and U2273 (N_2273,In_541,In_93);
nor U2274 (N_2274,In_76,In_106);
nor U2275 (N_2275,In_440,In_678);
and U2276 (N_2276,In_136,In_295);
nor U2277 (N_2277,In_515,In_183);
nand U2278 (N_2278,In_417,In_247);
nand U2279 (N_2279,In_230,In_169);
and U2280 (N_2280,In_31,In_356);
nor U2281 (N_2281,In_646,In_361);
nand U2282 (N_2282,In_557,In_262);
xnor U2283 (N_2283,In_7,In_447);
xnor U2284 (N_2284,In_126,In_154);
or U2285 (N_2285,In_11,In_327);
nand U2286 (N_2286,In_79,In_365);
and U2287 (N_2287,In_414,In_519);
nand U2288 (N_2288,In_427,In_381);
nand U2289 (N_2289,In_287,In_311);
nor U2290 (N_2290,In_727,In_45);
nor U2291 (N_2291,In_424,In_731);
nand U2292 (N_2292,In_387,In_18);
nand U2293 (N_2293,In_234,In_611);
nand U2294 (N_2294,In_648,In_6);
or U2295 (N_2295,In_493,In_473);
nor U2296 (N_2296,In_197,In_27);
and U2297 (N_2297,In_246,In_8);
and U2298 (N_2298,In_381,In_566);
nand U2299 (N_2299,In_189,In_537);
and U2300 (N_2300,In_363,In_237);
or U2301 (N_2301,In_230,In_546);
nand U2302 (N_2302,In_348,In_106);
nand U2303 (N_2303,In_693,In_709);
nor U2304 (N_2304,In_510,In_416);
nor U2305 (N_2305,In_565,In_581);
nor U2306 (N_2306,In_640,In_168);
or U2307 (N_2307,In_380,In_261);
and U2308 (N_2308,In_681,In_152);
nor U2309 (N_2309,In_735,In_726);
and U2310 (N_2310,In_261,In_538);
nand U2311 (N_2311,In_628,In_168);
nand U2312 (N_2312,In_144,In_263);
nand U2313 (N_2313,In_236,In_43);
nand U2314 (N_2314,In_226,In_392);
nor U2315 (N_2315,In_706,In_412);
nor U2316 (N_2316,In_128,In_482);
nor U2317 (N_2317,In_162,In_74);
nand U2318 (N_2318,In_4,In_140);
nand U2319 (N_2319,In_251,In_679);
nor U2320 (N_2320,In_35,In_733);
nor U2321 (N_2321,In_632,In_406);
nor U2322 (N_2322,In_182,In_165);
xor U2323 (N_2323,In_96,In_737);
or U2324 (N_2324,In_55,In_209);
or U2325 (N_2325,In_605,In_57);
and U2326 (N_2326,In_236,In_376);
or U2327 (N_2327,In_480,In_142);
nand U2328 (N_2328,In_251,In_172);
or U2329 (N_2329,In_462,In_4);
and U2330 (N_2330,In_457,In_336);
nand U2331 (N_2331,In_606,In_201);
xnor U2332 (N_2332,In_435,In_501);
nor U2333 (N_2333,In_695,In_558);
nor U2334 (N_2334,In_185,In_8);
and U2335 (N_2335,In_668,In_602);
nor U2336 (N_2336,In_33,In_585);
or U2337 (N_2337,In_436,In_43);
nor U2338 (N_2338,In_465,In_572);
nand U2339 (N_2339,In_478,In_515);
and U2340 (N_2340,In_382,In_41);
nand U2341 (N_2341,In_118,In_194);
nand U2342 (N_2342,In_276,In_63);
nand U2343 (N_2343,In_276,In_653);
or U2344 (N_2344,In_202,In_302);
xnor U2345 (N_2345,In_365,In_585);
nand U2346 (N_2346,In_29,In_545);
nand U2347 (N_2347,In_394,In_101);
nand U2348 (N_2348,In_470,In_32);
nor U2349 (N_2349,In_108,In_112);
nor U2350 (N_2350,In_743,In_507);
and U2351 (N_2351,In_117,In_567);
nor U2352 (N_2352,In_605,In_107);
and U2353 (N_2353,In_360,In_440);
and U2354 (N_2354,In_332,In_672);
or U2355 (N_2355,In_600,In_55);
and U2356 (N_2356,In_393,In_627);
nor U2357 (N_2357,In_477,In_134);
and U2358 (N_2358,In_688,In_543);
and U2359 (N_2359,In_683,In_587);
and U2360 (N_2360,In_656,In_345);
xnor U2361 (N_2361,In_35,In_610);
nor U2362 (N_2362,In_732,In_687);
and U2363 (N_2363,In_161,In_257);
or U2364 (N_2364,In_494,In_504);
and U2365 (N_2365,In_441,In_611);
or U2366 (N_2366,In_172,In_341);
nand U2367 (N_2367,In_332,In_478);
nor U2368 (N_2368,In_476,In_641);
or U2369 (N_2369,In_467,In_588);
nand U2370 (N_2370,In_196,In_338);
or U2371 (N_2371,In_354,In_628);
or U2372 (N_2372,In_181,In_589);
or U2373 (N_2373,In_284,In_357);
and U2374 (N_2374,In_579,In_234);
or U2375 (N_2375,In_746,In_274);
xnor U2376 (N_2376,In_456,In_302);
nor U2377 (N_2377,In_648,In_408);
and U2378 (N_2378,In_159,In_710);
nor U2379 (N_2379,In_49,In_577);
nor U2380 (N_2380,In_692,In_517);
nor U2381 (N_2381,In_631,In_500);
nand U2382 (N_2382,In_586,In_431);
xnor U2383 (N_2383,In_322,In_253);
or U2384 (N_2384,In_348,In_601);
or U2385 (N_2385,In_314,In_359);
nand U2386 (N_2386,In_484,In_698);
nor U2387 (N_2387,In_21,In_128);
nor U2388 (N_2388,In_244,In_91);
and U2389 (N_2389,In_691,In_335);
nor U2390 (N_2390,In_551,In_142);
or U2391 (N_2391,In_475,In_21);
and U2392 (N_2392,In_633,In_28);
nor U2393 (N_2393,In_535,In_224);
nor U2394 (N_2394,In_623,In_607);
xnor U2395 (N_2395,In_555,In_134);
nor U2396 (N_2396,In_230,In_700);
and U2397 (N_2397,In_465,In_371);
xnor U2398 (N_2398,In_498,In_58);
xor U2399 (N_2399,In_172,In_155);
or U2400 (N_2400,In_335,In_339);
xnor U2401 (N_2401,In_241,In_200);
or U2402 (N_2402,In_175,In_726);
xor U2403 (N_2403,In_741,In_470);
nor U2404 (N_2404,In_577,In_297);
nor U2405 (N_2405,In_70,In_425);
nor U2406 (N_2406,In_601,In_731);
nand U2407 (N_2407,In_20,In_335);
nor U2408 (N_2408,In_185,In_564);
or U2409 (N_2409,In_108,In_512);
or U2410 (N_2410,In_98,In_234);
or U2411 (N_2411,In_706,In_159);
nand U2412 (N_2412,In_213,In_359);
nand U2413 (N_2413,In_334,In_716);
or U2414 (N_2414,In_4,In_573);
or U2415 (N_2415,In_609,In_15);
or U2416 (N_2416,In_127,In_716);
nor U2417 (N_2417,In_154,In_446);
nand U2418 (N_2418,In_688,In_209);
or U2419 (N_2419,In_42,In_212);
nand U2420 (N_2420,In_468,In_654);
or U2421 (N_2421,In_284,In_59);
nor U2422 (N_2422,In_497,In_156);
and U2423 (N_2423,In_248,In_566);
nor U2424 (N_2424,In_221,In_80);
and U2425 (N_2425,In_383,In_101);
or U2426 (N_2426,In_264,In_681);
nor U2427 (N_2427,In_602,In_219);
or U2428 (N_2428,In_70,In_502);
nor U2429 (N_2429,In_213,In_111);
and U2430 (N_2430,In_183,In_433);
xnor U2431 (N_2431,In_474,In_279);
nor U2432 (N_2432,In_516,In_464);
nand U2433 (N_2433,In_2,In_373);
nand U2434 (N_2434,In_316,In_551);
or U2435 (N_2435,In_155,In_49);
xor U2436 (N_2436,In_621,In_540);
or U2437 (N_2437,In_702,In_316);
and U2438 (N_2438,In_161,In_641);
nor U2439 (N_2439,In_209,In_376);
or U2440 (N_2440,In_678,In_395);
xnor U2441 (N_2441,In_316,In_96);
xor U2442 (N_2442,In_566,In_211);
xor U2443 (N_2443,In_135,In_451);
nor U2444 (N_2444,In_42,In_525);
nor U2445 (N_2445,In_653,In_38);
and U2446 (N_2446,In_209,In_289);
nand U2447 (N_2447,In_30,In_7);
or U2448 (N_2448,In_504,In_121);
nor U2449 (N_2449,In_742,In_627);
xnor U2450 (N_2450,In_187,In_95);
nand U2451 (N_2451,In_494,In_244);
and U2452 (N_2452,In_368,In_306);
and U2453 (N_2453,In_381,In_665);
nand U2454 (N_2454,In_343,In_265);
nand U2455 (N_2455,In_593,In_522);
nand U2456 (N_2456,In_190,In_289);
and U2457 (N_2457,In_158,In_230);
and U2458 (N_2458,In_242,In_715);
nand U2459 (N_2459,In_567,In_542);
nor U2460 (N_2460,In_518,In_1);
nor U2461 (N_2461,In_38,In_424);
and U2462 (N_2462,In_717,In_165);
nor U2463 (N_2463,In_327,In_511);
and U2464 (N_2464,In_466,In_218);
xnor U2465 (N_2465,In_557,In_588);
nor U2466 (N_2466,In_149,In_152);
nand U2467 (N_2467,In_538,In_35);
and U2468 (N_2468,In_627,In_702);
and U2469 (N_2469,In_607,In_339);
nor U2470 (N_2470,In_545,In_423);
nand U2471 (N_2471,In_381,In_173);
nor U2472 (N_2472,In_198,In_694);
xnor U2473 (N_2473,In_99,In_67);
nor U2474 (N_2474,In_274,In_508);
and U2475 (N_2475,In_491,In_164);
and U2476 (N_2476,In_568,In_613);
nand U2477 (N_2477,In_245,In_277);
nand U2478 (N_2478,In_175,In_97);
or U2479 (N_2479,In_158,In_174);
nor U2480 (N_2480,In_446,In_439);
nand U2481 (N_2481,In_674,In_608);
nor U2482 (N_2482,In_63,In_523);
or U2483 (N_2483,In_231,In_636);
xor U2484 (N_2484,In_418,In_747);
and U2485 (N_2485,In_259,In_705);
or U2486 (N_2486,In_44,In_35);
and U2487 (N_2487,In_605,In_694);
nand U2488 (N_2488,In_440,In_205);
or U2489 (N_2489,In_278,In_533);
nand U2490 (N_2490,In_658,In_34);
nor U2491 (N_2491,In_327,In_412);
nand U2492 (N_2492,In_660,In_688);
nor U2493 (N_2493,In_645,In_674);
or U2494 (N_2494,In_343,In_735);
or U2495 (N_2495,In_400,In_105);
nor U2496 (N_2496,In_207,In_745);
nor U2497 (N_2497,In_658,In_137);
or U2498 (N_2498,In_332,In_534);
nand U2499 (N_2499,In_604,In_373);
or U2500 (N_2500,N_2194,N_1666);
or U2501 (N_2501,N_423,N_1682);
or U2502 (N_2502,N_1555,N_154);
nand U2503 (N_2503,N_2030,N_113);
or U2504 (N_2504,N_1784,N_1362);
nor U2505 (N_2505,N_1859,N_2253);
or U2506 (N_2506,N_232,N_753);
and U2507 (N_2507,N_945,N_808);
nand U2508 (N_2508,N_310,N_643);
or U2509 (N_2509,N_1292,N_2338);
nand U2510 (N_2510,N_2163,N_376);
and U2511 (N_2511,N_2259,N_2183);
or U2512 (N_2512,N_1103,N_2040);
nand U2513 (N_2513,N_2246,N_2447);
xnor U2514 (N_2514,N_324,N_2132);
nand U2515 (N_2515,N_462,N_1409);
nand U2516 (N_2516,N_1965,N_2362);
nor U2517 (N_2517,N_1188,N_2022);
xor U2518 (N_2518,N_1456,N_2358);
nand U2519 (N_2519,N_800,N_522);
nand U2520 (N_2520,N_1209,N_2087);
and U2521 (N_2521,N_359,N_1667);
or U2522 (N_2522,N_569,N_1658);
nor U2523 (N_2523,N_2160,N_1909);
nand U2524 (N_2524,N_481,N_21);
or U2525 (N_2525,N_1560,N_1948);
and U2526 (N_2526,N_134,N_595);
or U2527 (N_2527,N_1049,N_693);
nor U2528 (N_2528,N_1809,N_114);
nand U2529 (N_2529,N_989,N_238);
nand U2530 (N_2530,N_1070,N_1792);
nor U2531 (N_2531,N_2366,N_952);
nor U2532 (N_2532,N_1683,N_2387);
or U2533 (N_2533,N_1819,N_1613);
or U2534 (N_2534,N_830,N_2393);
or U2535 (N_2535,N_247,N_190);
or U2536 (N_2536,N_1363,N_2279);
xnor U2537 (N_2537,N_2458,N_1435);
or U2538 (N_2538,N_672,N_1731);
xnor U2539 (N_2539,N_373,N_1836);
xor U2540 (N_2540,N_2343,N_2267);
nand U2541 (N_2541,N_2435,N_2092);
nor U2542 (N_2542,N_1801,N_1381);
and U2543 (N_2543,N_1820,N_1984);
nand U2544 (N_2544,N_1419,N_1158);
xor U2545 (N_2545,N_39,N_1214);
nand U2546 (N_2546,N_1795,N_1598);
nand U2547 (N_2547,N_2175,N_457);
or U2548 (N_2548,N_341,N_768);
and U2549 (N_2549,N_600,N_611);
and U2550 (N_2550,N_1443,N_1061);
nor U2551 (N_2551,N_2011,N_777);
nor U2552 (N_2552,N_1594,N_2446);
xor U2553 (N_2553,N_1777,N_1018);
nor U2554 (N_2554,N_1046,N_428);
and U2555 (N_2555,N_1932,N_2115);
and U2556 (N_2556,N_1229,N_202);
nor U2557 (N_2557,N_292,N_667);
nand U2558 (N_2558,N_991,N_1811);
nor U2559 (N_2559,N_529,N_1524);
and U2560 (N_2560,N_2353,N_1614);
nand U2561 (N_2561,N_1254,N_1082);
nor U2562 (N_2562,N_943,N_1601);
nand U2563 (N_2563,N_2047,N_588);
nor U2564 (N_2564,N_2309,N_120);
xor U2565 (N_2565,N_687,N_2078);
and U2566 (N_2566,N_1392,N_658);
and U2567 (N_2567,N_156,N_1734);
nor U2568 (N_2568,N_869,N_524);
or U2569 (N_2569,N_319,N_408);
and U2570 (N_2570,N_165,N_2421);
and U2571 (N_2571,N_2096,N_2328);
or U2572 (N_2572,N_1349,N_1521);
and U2573 (N_2573,N_1438,N_841);
or U2574 (N_2574,N_105,N_2373);
or U2575 (N_2575,N_1403,N_1698);
or U2576 (N_2576,N_1951,N_1036);
nand U2577 (N_2577,N_1796,N_1257);
nand U2578 (N_2578,N_819,N_2146);
nand U2579 (N_2579,N_228,N_691);
nand U2580 (N_2580,N_1330,N_850);
nor U2581 (N_2581,N_107,N_2473);
or U2582 (N_2582,N_1239,N_2382);
or U2583 (N_2583,N_990,N_161);
or U2584 (N_2584,N_1689,N_563);
or U2585 (N_2585,N_2449,N_158);
xnor U2586 (N_2586,N_1747,N_2306);
nand U2587 (N_2587,N_1370,N_1743);
and U2588 (N_2588,N_182,N_1007);
and U2589 (N_2589,N_870,N_126);
nor U2590 (N_2590,N_2125,N_110);
or U2591 (N_2591,N_723,N_2344);
or U2592 (N_2592,N_1968,N_965);
and U2593 (N_2593,N_1204,N_262);
nand U2594 (N_2594,N_1118,N_1998);
or U2595 (N_2595,N_791,N_1117);
and U2596 (N_2596,N_251,N_538);
nor U2597 (N_2597,N_245,N_720);
xnor U2598 (N_2598,N_1173,N_936);
nor U2599 (N_2599,N_1723,N_1778);
or U2600 (N_2600,N_1448,N_663);
nor U2601 (N_2601,N_1919,N_24);
nor U2602 (N_2602,N_647,N_249);
and U2603 (N_2603,N_60,N_1741);
or U2604 (N_2604,N_698,N_1423);
and U2605 (N_2605,N_1464,N_561);
or U2606 (N_2606,N_492,N_1640);
or U2607 (N_2607,N_2263,N_129);
and U2608 (N_2608,N_1926,N_555);
and U2609 (N_2609,N_179,N_1359);
or U2610 (N_2610,N_1275,N_80);
and U2611 (N_2611,N_2468,N_1800);
nand U2612 (N_2612,N_342,N_1923);
nor U2613 (N_2613,N_1293,N_52);
xor U2614 (N_2614,N_437,N_616);
or U2615 (N_2615,N_856,N_1880);
or U2616 (N_2616,N_546,N_2354);
or U2617 (N_2617,N_823,N_1181);
and U2618 (N_2618,N_1245,N_1404);
nand U2619 (N_2619,N_1288,N_2315);
nand U2620 (N_2620,N_2091,N_681);
nand U2621 (N_2621,N_1092,N_2256);
nand U2622 (N_2622,N_1621,N_1452);
and U2623 (N_2623,N_534,N_637);
and U2624 (N_2624,N_1054,N_95);
or U2625 (N_2625,N_464,N_1029);
nand U2626 (N_2626,N_2470,N_1746);
and U2627 (N_2627,N_950,N_1259);
nand U2628 (N_2628,N_515,N_1608);
xor U2629 (N_2629,N_1168,N_1852);
and U2630 (N_2630,N_1371,N_1713);
nand U2631 (N_2631,N_1765,N_1099);
nor U2632 (N_2632,N_2217,N_557);
nand U2633 (N_2633,N_1350,N_1177);
nor U2634 (N_2634,N_1261,N_350);
nand U2635 (N_2635,N_1983,N_1062);
or U2636 (N_2636,N_2498,N_2365);
or U2637 (N_2637,N_131,N_1575);
or U2638 (N_2638,N_1969,N_2227);
and U2639 (N_2639,N_2189,N_683);
nand U2640 (N_2640,N_1833,N_1664);
nand U2641 (N_2641,N_436,N_1553);
nand U2642 (N_2642,N_627,N_1896);
and U2643 (N_2643,N_2207,N_1405);
nand U2644 (N_2644,N_883,N_811);
and U2645 (N_2645,N_56,N_734);
nor U2646 (N_2646,N_178,N_1040);
and U2647 (N_2647,N_2411,N_736);
xor U2648 (N_2648,N_1749,N_893);
xnor U2649 (N_2649,N_8,N_2260);
nand U2650 (N_2650,N_2117,N_374);
nor U2651 (N_2651,N_1520,N_150);
nand U2652 (N_2652,N_2381,N_2258);
xnor U2653 (N_2653,N_826,N_1043);
or U2654 (N_2654,N_2123,N_1073);
nor U2655 (N_2655,N_15,N_807);
or U2656 (N_2656,N_1160,N_1543);
and U2657 (N_2657,N_1961,N_1633);
nand U2658 (N_2658,N_751,N_455);
or U2659 (N_2659,N_981,N_1697);
nand U2660 (N_2660,N_1059,N_2351);
and U2661 (N_2661,N_1535,N_864);
nor U2662 (N_2662,N_2109,N_2185);
and U2663 (N_2663,N_521,N_2172);
nand U2664 (N_2664,N_122,N_294);
nor U2665 (N_2665,N_1722,N_142);
or U2666 (N_2666,N_1476,N_699);
or U2667 (N_2667,N_2417,N_700);
or U2668 (N_2668,N_1990,N_2436);
nor U2669 (N_2669,N_1367,N_340);
xor U2670 (N_2670,N_1321,N_2289);
and U2671 (N_2671,N_380,N_2406);
nor U2672 (N_2672,N_1441,N_716);
nor U2673 (N_2673,N_1651,N_1055);
and U2674 (N_2674,N_2198,N_194);
and U2675 (N_2675,N_102,N_2312);
and U2676 (N_2676,N_1434,N_912);
nand U2677 (N_2677,N_1974,N_1869);
nand U2678 (N_2678,N_2340,N_470);
or U2679 (N_2679,N_388,N_2467);
xnor U2680 (N_2680,N_2089,N_419);
or U2681 (N_2681,N_2334,N_630);
or U2682 (N_2682,N_1557,N_1510);
xnor U2683 (N_2683,N_934,N_2173);
xnor U2684 (N_2684,N_103,N_325);
nand U2685 (N_2685,N_2196,N_1729);
nor U2686 (N_2686,N_2081,N_996);
or U2687 (N_2687,N_1996,N_1752);
nor U2688 (N_2688,N_1922,N_358);
or U2689 (N_2689,N_2039,N_1121);
and U2690 (N_2690,N_282,N_903);
nor U2691 (N_2691,N_2445,N_2477);
nand U2692 (N_2692,N_1324,N_977);
nor U2693 (N_2693,N_2368,N_668);
or U2694 (N_2694,N_1347,N_270);
and U2695 (N_2695,N_493,N_1562);
or U2696 (N_2696,N_1461,N_2367);
and U2697 (N_2697,N_449,N_1935);
nand U2698 (N_2698,N_2157,N_2032);
nand U2699 (N_2699,N_2300,N_1891);
nor U2700 (N_2700,N_382,N_812);
xor U2701 (N_2701,N_1774,N_1186);
nor U2702 (N_2702,N_1313,N_1477);
nor U2703 (N_2703,N_653,N_301);
nand U2704 (N_2704,N_705,N_256);
and U2705 (N_2705,N_2150,N_1439);
nor U2706 (N_2706,N_2097,N_295);
xor U2707 (N_2707,N_1766,N_1875);
nor U2708 (N_2708,N_939,N_430);
or U2709 (N_2709,N_1629,N_1114);
or U2710 (N_2710,N_1794,N_654);
nor U2711 (N_2711,N_845,N_542);
and U2712 (N_2712,N_2021,N_1033);
nor U2713 (N_2713,N_2288,N_2156);
and U2714 (N_2714,N_2184,N_1915);
and U2715 (N_2715,N_786,N_1034);
or U2716 (N_2716,N_589,N_1587);
nand U2717 (N_2717,N_1609,N_724);
nor U2718 (N_2718,N_69,N_1789);
and U2719 (N_2719,N_1041,N_1430);
and U2720 (N_2720,N_548,N_496);
xnor U2721 (N_2721,N_1767,N_2401);
nand U2722 (N_2722,N_1332,N_1652);
nand U2723 (N_2723,N_298,N_944);
and U2724 (N_2724,N_2164,N_1690);
nor U2725 (N_2725,N_2405,N_619);
nand U2726 (N_2726,N_258,N_170);
xor U2727 (N_2727,N_2178,N_2451);
or U2728 (N_2728,N_1720,N_335);
or U2729 (N_2729,N_196,N_16);
nand U2730 (N_2730,N_2273,N_1178);
nor U2731 (N_2731,N_495,N_1802);
or U2732 (N_2732,N_1377,N_396);
nand U2733 (N_2733,N_626,N_740);
and U2734 (N_2734,N_100,N_463);
or U2735 (N_2735,N_207,N_1716);
nor U2736 (N_2736,N_1316,N_1606);
xor U2737 (N_2737,N_886,N_223);
nand U2738 (N_2738,N_1374,N_1740);
and U2739 (N_2739,N_1402,N_401);
xnor U2740 (N_2740,N_2059,N_1101);
and U2741 (N_2741,N_1591,N_1110);
nand U2742 (N_2742,N_1527,N_2474);
xnor U2743 (N_2743,N_767,N_2023);
or U2744 (N_2744,N_1718,N_1270);
nor U2745 (N_2745,N_2229,N_1266);
nor U2746 (N_2746,N_1098,N_2348);
or U2747 (N_2747,N_1433,N_1876);
xor U2748 (N_2748,N_553,N_1067);
and U2749 (N_2749,N_1424,N_306);
and U2750 (N_2750,N_2107,N_584);
xnor U2751 (N_2751,N_1281,N_2031);
nor U2752 (N_2752,N_1782,N_750);
or U2753 (N_2753,N_2442,N_473);
or U2754 (N_2754,N_1821,N_1425);
and U2755 (N_2755,N_1361,N_47);
nand U2756 (N_2756,N_180,N_586);
nor U2757 (N_2757,N_565,N_2298);
or U2758 (N_2758,N_773,N_1742);
nor U2759 (N_2759,N_1907,N_1053);
nor U2760 (N_2760,N_1309,N_528);
nor U2761 (N_2761,N_1421,N_2314);
xnor U2762 (N_2762,N_1336,N_1842);
or U2763 (N_2763,N_964,N_628);
or U2764 (N_2764,N_11,N_321);
nand U2765 (N_2765,N_2018,N_549);
or U2766 (N_2766,N_2086,N_1297);
nand U2767 (N_2767,N_1908,N_1194);
and U2768 (N_2768,N_1847,N_222);
nand U2769 (N_2769,N_1903,N_1171);
or U2770 (N_2770,N_979,N_2235);
nand U2771 (N_2771,N_1963,N_1704);
nor U2772 (N_2772,N_2228,N_2119);
nand U2773 (N_2773,N_1646,N_1659);
nor U2774 (N_2774,N_1132,N_853);
nor U2775 (N_2775,N_2006,N_1516);
nand U2776 (N_2776,N_1385,N_1702);
and U2777 (N_2777,N_1661,N_1979);
nor U2778 (N_2778,N_821,N_276);
nand U2779 (N_2779,N_576,N_1016);
and U2780 (N_2780,N_897,N_1406);
nand U2781 (N_2781,N_2350,N_661);
or U2782 (N_2782,N_439,N_1502);
or U2783 (N_2783,N_422,N_562);
and U2784 (N_2784,N_1564,N_1879);
nand U2785 (N_2785,N_1576,N_928);
xnor U2786 (N_2786,N_1216,N_2280);
xor U2787 (N_2787,N_545,N_2307);
nand U2788 (N_2788,N_1170,N_2179);
and U2789 (N_2789,N_608,N_506);
or U2790 (N_2790,N_2181,N_1739);
xnor U2791 (N_2791,N_2476,N_2045);
nor U2792 (N_2792,N_948,N_313);
nand U2793 (N_2793,N_1641,N_266);
nor U2794 (N_2794,N_685,N_2310);
and U2795 (N_2795,N_101,N_1299);
nor U2796 (N_2796,N_2482,N_55);
or U2797 (N_2797,N_1351,N_2360);
or U2798 (N_2798,N_1133,N_185);
or U2799 (N_2799,N_967,N_848);
and U2800 (N_2800,N_1572,N_959);
xnor U2801 (N_2801,N_1202,N_1672);
xor U2802 (N_2802,N_1900,N_2292);
and U2803 (N_2803,N_802,N_369);
nor U2804 (N_2804,N_2054,N_1737);
xor U2805 (N_2805,N_1144,N_390);
or U2806 (N_2806,N_2322,N_1113);
and U2807 (N_2807,N_2215,N_363);
nor U2808 (N_2808,N_25,N_746);
or U2809 (N_2809,N_828,N_1655);
xnor U2810 (N_2810,N_1512,N_930);
and U2811 (N_2811,N_960,N_917);
or U2812 (N_2812,N_2294,N_2145);
or U2813 (N_2813,N_1180,N_2383);
nand U2814 (N_2814,N_138,N_1203);
and U2815 (N_2815,N_434,N_1224);
xor U2816 (N_2816,N_2187,N_1486);
and U2817 (N_2817,N_2068,N_2141);
and U2818 (N_2818,N_523,N_1289);
nand U2819 (N_2819,N_1420,N_1255);
and U2820 (N_2820,N_2297,N_1941);
xnor U2821 (N_2821,N_2004,N_629);
or U2822 (N_2822,N_797,N_2493);
and U2823 (N_2823,N_2323,N_1416);
nor U2824 (N_2824,N_919,N_938);
nor U2825 (N_2825,N_1124,N_1724);
nor U2826 (N_2826,N_7,N_925);
nand U2827 (N_2827,N_526,N_404);
nand U2828 (N_2828,N_2330,N_1952);
or U2829 (N_2829,N_448,N_308);
or U2830 (N_2830,N_764,N_1342);
nand U2831 (N_2831,N_417,N_1693);
or U2832 (N_2832,N_1943,N_2149);
xnor U2833 (N_2833,N_707,N_1584);
nor U2834 (N_2834,N_638,N_1414);
or U2835 (N_2835,N_1084,N_1389);
and U2836 (N_2836,N_2152,N_242);
or U2837 (N_2837,N_1870,N_62);
nor U2838 (N_2838,N_1408,N_484);
nor U2839 (N_2839,N_982,N_1328);
nor U2840 (N_2840,N_1000,N_1921);
nor U2841 (N_2841,N_1938,N_927);
and U2842 (N_2842,N_2035,N_835);
xnor U2843 (N_2843,N_754,N_1123);
and U2844 (N_2844,N_2240,N_2019);
and U2845 (N_2845,N_874,N_2245);
nand U2846 (N_2846,N_1278,N_1507);
or U2847 (N_2847,N_1319,N_805);
nor U2848 (N_2848,N_1858,N_2209);
nor U2849 (N_2849,N_2127,N_2203);
xor U2850 (N_2850,N_214,N_1494);
nor U2851 (N_2851,N_739,N_1413);
or U2852 (N_2852,N_1945,N_1992);
xnor U2853 (N_2853,N_508,N_353);
nor U2854 (N_2854,N_935,N_218);
and U2855 (N_2855,N_145,N_88);
nor U2856 (N_2856,N_116,N_348);
and U2857 (N_2857,N_1088,N_1586);
or U2858 (N_2858,N_1705,N_2155);
and U2859 (N_2859,N_890,N_891);
and U2860 (N_2860,N_849,N_1942);
nor U2861 (N_2861,N_1369,N_832);
nor U2862 (N_2862,N_1868,N_1872);
nor U2863 (N_2863,N_1376,N_1481);
and U2864 (N_2864,N_2250,N_984);
nor U2865 (N_2865,N_1159,N_1615);
and U2866 (N_2866,N_2494,N_591);
nor U2867 (N_2867,N_975,N_2057);
xnor U2868 (N_2868,N_1709,N_1933);
and U2869 (N_2869,N_192,N_1212);
nand U2870 (N_2870,N_143,N_1981);
or U2871 (N_2871,N_1972,N_880);
and U2872 (N_2872,N_1378,N_433);
and U2873 (N_2873,N_818,N_780);
xor U2874 (N_2874,N_2414,N_132);
and U2875 (N_2875,N_907,N_1388);
or U2876 (N_2876,N_360,N_1253);
nand U2877 (N_2877,N_1599,N_2180);
and U2878 (N_2878,N_621,N_755);
or U2879 (N_2879,N_1806,N_1544);
nor U2880 (N_2880,N_1276,N_1152);
xnor U2881 (N_2881,N_957,N_1567);
nand U2882 (N_2882,N_1597,N_625);
nand U2883 (N_2883,N_1662,N_894);
nor U2884 (N_2884,N_833,N_128);
or U2885 (N_2885,N_2176,N_1341);
nor U2886 (N_2886,N_1344,N_1617);
and U2887 (N_2887,N_487,N_533);
or U2888 (N_2888,N_1927,N_507);
xnor U2889 (N_2889,N_1860,N_947);
or U2890 (N_2890,N_2169,N_712);
or U2891 (N_2891,N_99,N_1190);
nand U2892 (N_2892,N_166,N_211);
and U2893 (N_2893,N_568,N_488);
nand U2894 (N_2894,N_689,N_642);
and U2895 (N_2895,N_1487,N_806);
or U2896 (N_2896,N_79,N_1048);
nand U2897 (N_2897,N_824,N_1220);
nor U2898 (N_2898,N_1387,N_188);
or U2899 (N_2899,N_160,N_1480);
or U2900 (N_2900,N_2038,N_109);
or U2901 (N_2901,N_420,N_167);
or U2902 (N_2902,N_1395,N_1009);
and U2903 (N_2903,N_787,N_1375);
and U2904 (N_2904,N_1338,N_415);
xor U2905 (N_2905,N_617,N_1753);
or U2906 (N_2906,N_995,N_2147);
nand U2907 (N_2907,N_680,N_253);
and U2908 (N_2908,N_351,N_778);
nor U2909 (N_2909,N_867,N_1892);
nand U2910 (N_2910,N_163,N_1014);
or U2911 (N_2911,N_1910,N_328);
or U2912 (N_2912,N_1146,N_762);
and U2913 (N_2913,N_123,N_2475);
nand U2914 (N_2914,N_2214,N_392);
or U2915 (N_2915,N_1066,N_1934);
and U2916 (N_2916,N_1138,N_547);
and U2917 (N_2917,N_774,N_599);
nor U2918 (N_2918,N_1580,N_877);
nand U2919 (N_2919,N_1322,N_2302);
nand U2920 (N_2920,N_2463,N_790);
or U2921 (N_2921,N_367,N_840);
nor U2922 (N_2922,N_862,N_2371);
and U2923 (N_2923,N_2211,N_476);
and U2924 (N_2924,N_1217,N_692);
xor U2925 (N_2925,N_1358,N_2153);
nand U2926 (N_2926,N_1714,N_879);
nand U2927 (N_2927,N_1145,N_210);
nor U2928 (N_2928,N_1,N_1468);
nand U2929 (N_2929,N_135,N_924);
nor U2930 (N_2930,N_2225,N_1240);
or U2931 (N_2931,N_1855,N_124);
and U2932 (N_2932,N_1156,N_1883);
xnor U2933 (N_2933,N_2027,N_1788);
xnor U2934 (N_2934,N_1081,N_1304);
and U2935 (N_2935,N_1356,N_26);
nand U2936 (N_2936,N_2384,N_2492);
and U2937 (N_2937,N_387,N_1256);
or U2938 (N_2938,N_1491,N_1696);
nor U2939 (N_2939,N_1492,N_1967);
or U2940 (N_2940,N_2304,N_875);
and U2941 (N_2941,N_1238,N_48);
nand U2942 (N_2942,N_594,N_861);
nor U2943 (N_2943,N_275,N_2378);
or U2944 (N_2944,N_1906,N_570);
and U2945 (N_2945,N_2299,N_908);
nand U2946 (N_2946,N_2252,N_1274);
or U2947 (N_2947,N_941,N_1712);
and U2948 (N_2948,N_651,N_648);
nand U2949 (N_2949,N_1195,N_785);
and U2950 (N_2950,N_1115,N_1807);
nand U2951 (N_2951,N_1856,N_347);
nor U2952 (N_2952,N_421,N_585);
nor U2953 (N_2953,N_2231,N_997);
nand U2954 (N_2954,N_1588,N_623);
nor U2955 (N_2955,N_104,N_1686);
nand U2956 (N_2956,N_1684,N_1277);
xnor U2957 (N_2957,N_789,N_999);
xnor U2958 (N_2958,N_1611,N_43);
or U2959 (N_2959,N_2264,N_10);
nor U2960 (N_2960,N_2379,N_299);
nor U2961 (N_2961,N_1399,N_1355);
or U2962 (N_2962,N_511,N_1104);
nor U2963 (N_2963,N_610,N_1989);
and U2964 (N_2964,N_1432,N_193);
nor U2965 (N_2965,N_2313,N_1843);
and U2966 (N_2966,N_973,N_1089);
and U2967 (N_2967,N_2266,N_516);
and U2968 (N_2968,N_2193,N_2462);
or U2969 (N_2969,N_1635,N_920);
and U2970 (N_2970,N_771,N_371);
and U2971 (N_2971,N_1340,N_277);
or U2972 (N_2972,N_1757,N_901);
nor U2973 (N_2973,N_1940,N_318);
and U2974 (N_2974,N_1947,N_2485);
xor U2975 (N_2975,N_2100,N_690);
and U2976 (N_2976,N_1565,N_2080);
and U2977 (N_2977,N_940,N_98);
and U2978 (N_2978,N_514,N_2465);
nor U2979 (N_2979,N_1444,N_168);
or U2980 (N_2980,N_682,N_587);
and U2981 (N_2981,N_23,N_283);
nand U2982 (N_2982,N_157,N_96);
nor U2983 (N_2983,N_775,N_2425);
and U2984 (N_2984,N_1023,N_1725);
nand U2985 (N_2985,N_1978,N_1519);
nor U2986 (N_2986,N_2284,N_756);
or U2987 (N_2987,N_477,N_860);
and U2988 (N_2988,N_2174,N_106);
and U2989 (N_2989,N_1727,N_1415);
or U2990 (N_2990,N_1864,N_2305);
nand U2991 (N_2991,N_913,N_1971);
nor U2992 (N_2992,N_2443,N_498);
nand U2993 (N_2993,N_1525,N_1656);
nor U2994 (N_2994,N_1244,N_1648);
nor U2995 (N_2995,N_1877,N_2254);
nand U2996 (N_2996,N_1447,N_2437);
or U2997 (N_2997,N_361,N_1808);
or U2998 (N_2998,N_2438,N_1366);
nor U2999 (N_2999,N_2095,N_851);
or U3000 (N_3000,N_87,N_618);
nor U3001 (N_3001,N_1096,N_1215);
and U3002 (N_3002,N_1083,N_1654);
nand U3003 (N_3003,N_2380,N_315);
or U3004 (N_3004,N_1632,N_933);
or U3005 (N_3005,N_1760,N_2131);
nand U3006 (N_3006,N_153,N_1065);
or U3007 (N_3007,N_326,N_813);
and U3008 (N_3008,N_1095,N_409);
or U3009 (N_3009,N_727,N_6);
xor U3010 (N_3010,N_2014,N_2165);
and U3011 (N_3011,N_2191,N_953);
nand U3012 (N_3012,N_1549,N_794);
nand U3013 (N_3013,N_2058,N_1176);
and U3014 (N_3014,N_1164,N_1057);
or U3015 (N_3015,N_1446,N_1368);
or U3016 (N_3016,N_2345,N_831);
nand U3017 (N_3017,N_1673,N_911);
or U3018 (N_3018,N_1296,N_378);
nor U3019 (N_3019,N_1738,N_1008);
or U3020 (N_3020,N_41,N_93);
and U3021 (N_3021,N_147,N_2083);
and U3022 (N_3022,N_2070,N_1312);
nor U3023 (N_3023,N_184,N_1100);
nor U3024 (N_3024,N_453,N_983);
nand U3025 (N_3025,N_1210,N_281);
nor U3026 (N_3026,N_2496,N_14);
and U3027 (N_3027,N_1895,N_2017);
xor U3028 (N_3028,N_1071,N_1848);
and U3029 (N_3029,N_1282,N_1687);
or U3030 (N_3030,N_140,N_942);
nor U3031 (N_3031,N_899,N_343);
and U3032 (N_3032,N_486,N_1364);
nand U3033 (N_3033,N_956,N_2287);
nor U3034 (N_3034,N_2008,N_923);
nor U3035 (N_3035,N_604,N_918);
or U3036 (N_3036,N_741,N_1700);
and U3037 (N_3037,N_1816,N_1745);
and U3038 (N_3038,N_1552,N_398);
or U3039 (N_3039,N_1015,N_2201);
and U3040 (N_3040,N_344,N_1701);
and U3041 (N_3041,N_2456,N_173);
xor U3042 (N_3042,N_2478,N_1691);
nor U3043 (N_3043,N_779,N_1568);
nor U3044 (N_3044,N_1068,N_2077);
nand U3045 (N_3045,N_1192,N_1668);
or U3046 (N_3046,N_1810,N_635);
nand U3047 (N_3047,N_759,N_82);
nor U3048 (N_3048,N_827,N_71);
or U3049 (N_3049,N_1024,N_2349);
and U3050 (N_3050,N_2416,N_1636);
and U3051 (N_3051,N_1284,N_1175);
and U3052 (N_3052,N_1726,N_579);
nand U3053 (N_3053,N_1286,N_1531);
or U3054 (N_3054,N_1382,N_149);
nand U3055 (N_3055,N_717,N_410);
nand U3056 (N_3056,N_537,N_490);
and U3057 (N_3057,N_505,N_2321);
nand U3058 (N_3058,N_279,N_748);
nor U3059 (N_3059,N_1812,N_447);
nand U3060 (N_3060,N_213,N_31);
nand U3061 (N_3061,N_2461,N_431);
or U3062 (N_3062,N_2223,N_1899);
nor U3063 (N_3063,N_852,N_2116);
nor U3064 (N_3064,N_384,N_1166);
xnor U3065 (N_3065,N_1853,N_1920);
nor U3066 (N_3066,N_804,N_815);
nand U3067 (N_3067,N_1897,N_2372);
and U3068 (N_3068,N_1473,N_1548);
nand U3069 (N_3069,N_1830,N_1754);
nand U3070 (N_3070,N_2093,N_1660);
nor U3071 (N_3071,N_2063,N_2234);
nand U3072 (N_3072,N_201,N_1600);
and U3073 (N_3073,N_349,N_1596);
and U3074 (N_3074,N_331,N_1189);
nor U3075 (N_3075,N_28,N_1841);
xnor U3076 (N_3076,N_2272,N_1108);
nand U3077 (N_3077,N_2082,N_1249);
xor U3078 (N_3078,N_2440,N_825);
nand U3079 (N_3079,N_2238,N_1032);
and U3080 (N_3080,N_246,N_2408);
nor U3081 (N_3081,N_882,N_2283);
or U3082 (N_3082,N_655,N_1028);
nor U3083 (N_3083,N_2212,N_1026);
and U3084 (N_3084,N_722,N_1167);
or U3085 (N_3085,N_2385,N_233);
and U3086 (N_3086,N_1703,N_702);
nand U3087 (N_3087,N_2392,N_1437);
or U3088 (N_3088,N_483,N_2355);
nand U3089 (N_3089,N_2369,N_726);
nor U3090 (N_3090,N_613,N_2177);
and U3091 (N_3091,N_1307,N_1975);
nand U3092 (N_3092,N_2143,N_1397);
nor U3093 (N_3093,N_1593,N_1861);
and U3094 (N_3094,N_554,N_1241);
or U3095 (N_3095,N_1823,N_1056);
and U3096 (N_3096,N_2419,N_578);
nand U3097 (N_3097,N_2395,N_92);
or U3098 (N_3098,N_2060,N_1574);
xnor U3099 (N_3099,N_904,N_1157);
nor U3100 (N_3100,N_1581,N_1005);
nand U3101 (N_3101,N_465,N_2277);
xnor U3102 (N_3102,N_509,N_2084);
or U3103 (N_3103,N_1125,N_1290);
and U3104 (N_3104,N_1523,N_742);
nor U3105 (N_3105,N_1187,N_776);
nand U3106 (N_3106,N_2327,N_1917);
nor U3107 (N_3107,N_302,N_974);
and U3108 (N_3108,N_1271,N_873);
nor U3109 (N_3109,N_921,N_2426);
nor U3110 (N_3110,N_293,N_1226);
and U3111 (N_3111,N_1643,N_2166);
or U3112 (N_3112,N_566,N_2010);
nand U3113 (N_3113,N_1913,N_1455);
or U3114 (N_3114,N_1205,N_1429);
nand U3115 (N_3115,N_2453,N_2110);
or U3116 (N_3116,N_1206,N_1094);
or U3117 (N_3117,N_1506,N_2200);
or U3118 (N_3118,N_972,N_1396);
nand U3119 (N_3119,N_479,N_968);
nor U3120 (N_3120,N_1551,N_543);
xnor U3121 (N_3121,N_1825,N_1208);
nand U3122 (N_3122,N_1694,N_677);
and U3123 (N_3123,N_580,N_108);
nand U3124 (N_3124,N_1463,N_30);
nand U3125 (N_3125,N_2457,N_1268);
nand U3126 (N_3126,N_1069,N_497);
xnor U3127 (N_3127,N_1243,N_1928);
nor U3128 (N_3128,N_2041,N_45);
nor U3129 (N_3129,N_272,N_847);
nor U3130 (N_3130,N_2391,N_1165);
nand U3131 (N_3131,N_2230,N_386);
or U3132 (N_3132,N_53,N_675);
nand U3133 (N_3133,N_255,N_552);
nor U3134 (N_3134,N_174,N_2337);
nor U3135 (N_3135,N_1503,N_402);
xor U3136 (N_3136,N_1193,N_1287);
nor U3137 (N_3137,N_2428,N_1962);
nand U3138 (N_3138,N_889,N_2341);
nor U3139 (N_3139,N_1736,N_650);
or U3140 (N_3140,N_1571,N_782);
nor U3141 (N_3141,N_602,N_1246);
nor U3142 (N_3142,N_994,N_1949);
or U3143 (N_3143,N_530,N_733);
and U3144 (N_3144,N_2135,N_1001);
nand U3145 (N_3145,N_2396,N_252);
nor U3146 (N_3146,N_1237,N_2422);
nand U3147 (N_3147,N_2013,N_405);
nor U3148 (N_3148,N_83,N_2167);
and U3149 (N_3149,N_2495,N_489);
nor U3150 (N_3150,N_1936,N_2265);
nand U3151 (N_3151,N_1905,N_1105);
and U3152 (N_3152,N_2318,N_426);
nor U3153 (N_3153,N_1302,N_1051);
and U3154 (N_3154,N_2226,N_2377);
and U3155 (N_3155,N_1522,N_1674);
and U3156 (N_3156,N_221,N_1779);
nor U3157 (N_3157,N_2376,N_2195);
nor U3158 (N_3158,N_624,N_391);
nand U3159 (N_3159,N_662,N_171);
and U3160 (N_3160,N_1019,N_2413);
or U3161 (N_3161,N_155,N_1207);
or U3162 (N_3162,N_237,N_327);
and U3163 (N_3163,N_1730,N_1470);
xor U3164 (N_3164,N_1323,N_1805);
nand U3165 (N_3165,N_590,N_27);
nand U3166 (N_3166,N_1865,N_1042);
or U3167 (N_3167,N_2486,N_582);
or U3168 (N_3168,N_267,N_631);
and U3169 (N_3169,N_1479,N_905);
nor U3170 (N_3170,N_356,N_1653);
xor U3171 (N_3171,N_769,N_97);
nor U3172 (N_3172,N_63,N_35);
or U3173 (N_3173,N_2316,N_148);
or U3174 (N_3174,N_2268,N_2460);
or U3175 (N_3175,N_254,N_1197);
nand U3176 (N_3176,N_393,N_708);
xor U3177 (N_3177,N_892,N_2237);
and U3178 (N_3178,N_993,N_1604);
nor U3179 (N_3179,N_614,N_1874);
nor U3180 (N_3180,N_581,N_1154);
nor U3181 (N_3181,N_1116,N_2424);
and U3182 (N_3182,N_2346,N_2398);
or U3183 (N_3183,N_531,N_316);
and U3184 (N_3184,N_1185,N_460);
or U3185 (N_3185,N_783,N_1258);
nor U3186 (N_3186,N_2037,N_1944);
xnor U3187 (N_3187,N_674,N_446);
nor U3188 (N_3188,N_2242,N_1579);
nor U3189 (N_3189,N_2003,N_969);
nand U3190 (N_3190,N_472,N_288);
nor U3191 (N_3191,N_474,N_2048);
xnor U3192 (N_3192,N_2448,N_1803);
or U3193 (N_3193,N_713,N_801);
or U3194 (N_3194,N_2130,N_1793);
nor U3195 (N_3195,N_1162,N_2455);
and U3196 (N_3196,N_536,N_743);
nor U3197 (N_3197,N_2361,N_471);
nor U3198 (N_3198,N_2454,N_1086);
nand U3199 (N_3199,N_72,N_259);
or U3200 (N_3200,N_1010,N_571);
or U3201 (N_3201,N_671,N_1151);
nor U3202 (N_3202,N_2098,N_1561);
and U3203 (N_3203,N_1398,N_2085);
nor U3204 (N_3204,N_441,N_2247);
nand U3205 (N_3205,N_721,N_715);
nand U3206 (N_3206,N_958,N_1454);
and U3207 (N_3207,N_1862,N_1744);
and U3208 (N_3208,N_1995,N_273);
nor U3209 (N_3209,N_729,N_2190);
nand U3210 (N_3210,N_837,N_858);
or U3211 (N_3211,N_440,N_1228);
and U3212 (N_3212,N_2142,N_1179);
nand U3213 (N_3213,N_1474,N_2397);
and U3214 (N_3214,N_679,N_2319);
nor U3215 (N_3215,N_1326,N_1234);
and U3216 (N_3216,N_435,N_1348);
nor U3217 (N_3217,N_1422,N_502);
and U3218 (N_3218,N_694,N_229);
nor U3219 (N_3219,N_1102,N_1300);
nor U3220 (N_3220,N_2113,N_1485);
and U3221 (N_3221,N_855,N_1556);
nor U3222 (N_3222,N_931,N_839);
and U3223 (N_3223,N_2356,N_612);
and U3224 (N_3224,N_1832,N_1269);
and U3225 (N_3225,N_598,N_1320);
nand U3226 (N_3226,N_1265,N_1846);
or U3227 (N_3227,N_70,N_2029);
nor U3228 (N_3228,N_1889,N_1924);
nor U3229 (N_3229,N_1669,N_985);
or U3230 (N_3230,N_66,N_199);
or U3231 (N_3231,N_718,N_2136);
and U3232 (N_3232,N_2274,N_763);
nor U3233 (N_3233,N_719,N_227);
or U3234 (N_3234,N_1251,N_532);
xnor U3235 (N_3235,N_1457,N_2363);
and U3236 (N_3236,N_1139,N_1699);
and U3237 (N_3237,N_645,N_2076);
nand U3238 (N_3238,N_1785,N_312);
xnor U3239 (N_3239,N_1680,N_208);
or U3240 (N_3240,N_871,N_1153);
nor U3241 (N_3241,N_1534,N_2161);
and U3242 (N_3242,N_1003,N_1657);
or U3243 (N_3243,N_2016,N_2055);
or U3244 (N_3244,N_172,N_606);
or U3245 (N_3245,N_2335,N_1025);
nand U3246 (N_3246,N_1991,N_656);
or U3247 (N_3247,N_452,N_1223);
or U3248 (N_3248,N_711,N_1465);
nor U3249 (N_3249,N_2257,N_187);
or U3250 (N_3250,N_1076,N_127);
nor U3251 (N_3251,N_141,N_2199);
and U3252 (N_3252,N_485,N_898);
or U3253 (N_3253,N_1333,N_1038);
or U3254 (N_3254,N_1143,N_250);
or U3255 (N_3255,N_459,N_1536);
nor U3256 (N_3256,N_1291,N_2034);
xnor U3257 (N_3257,N_2489,N_1140);
nor U3258 (N_3258,N_2216,N_900);
or U3259 (N_3259,N_1295,N_2009);
or U3260 (N_3260,N_67,N_368);
nand U3261 (N_3261,N_1645,N_843);
nor U3262 (N_3262,N_732,N_203);
nor U3263 (N_3263,N_1735,N_2317);
or U3264 (N_3264,N_1022,N_257);
or U3265 (N_3265,N_1623,N_263);
xnor U3266 (N_3266,N_2137,N_593);
nor U3267 (N_3267,N_2423,N_1155);
and U3268 (N_3268,N_2062,N_334);
and U3269 (N_3269,N_1528,N_962);
or U3270 (N_3270,N_2202,N_1106);
and U3271 (N_3271,N_1532,N_660);
xor U3272 (N_3272,N_1692,N_2386);
and U3273 (N_3273,N_125,N_501);
nor U3274 (N_3274,N_1314,N_2134);
nor U3275 (N_3275,N_1393,N_2472);
xnor U3276 (N_3276,N_909,N_1511);
and U3277 (N_3277,N_1970,N_1471);
nor U3278 (N_3278,N_639,N_1235);
or U3279 (N_3279,N_269,N_2464);
xnor U3280 (N_3280,N_1835,N_333);
xor U3281 (N_3281,N_2213,N_1466);
or U3282 (N_3282,N_1685,N_520);
and U3283 (N_3283,N_244,N_622);
and U3284 (N_3284,N_1925,N_2427);
or U3285 (N_3285,N_42,N_2241);
or U3286 (N_3286,N_1997,N_370);
or U3287 (N_3287,N_1573,N_1762);
or U3288 (N_3288,N_1017,N_198);
and U3289 (N_3289,N_268,N_480);
xor U3290 (N_3290,N_89,N_2430);
and U3291 (N_3291,N_1063,N_2364);
nand U3292 (N_3292,N_38,N_77);
nor U3293 (N_3293,N_271,N_829);
nand U3294 (N_3294,N_1977,N_20);
nand U3295 (N_3295,N_1436,N_1353);
or U3296 (N_3296,N_152,N_2222);
xor U3297 (N_3297,N_1849,N_2036);
and U3298 (N_3298,N_1484,N_1301);
nand U3299 (N_3299,N_1930,N_2069);
or U3300 (N_3300,N_1514,N_2159);
nand U3301 (N_3301,N_9,N_1976);
nand U3302 (N_3302,N_1751,N_929);
or U3303 (N_3303,N_1093,N_1442);
and U3304 (N_3304,N_1365,N_1770);
and U3305 (N_3305,N_541,N_1147);
nand U3306 (N_3306,N_2106,N_1515);
nor U3307 (N_3307,N_5,N_1719);
or U3308 (N_3308,N_1417,N_1822);
nor U3309 (N_3309,N_1529,N_2410);
and U3310 (N_3310,N_906,N_427);
or U3311 (N_3311,N_1247,N_987);
and U3312 (N_3312,N_226,N_1458);
nand U3313 (N_3313,N_596,N_881);
or U3314 (N_3314,N_884,N_2444);
or U3315 (N_3315,N_1431,N_1182);
xnor U3316 (N_3316,N_50,N_1126);
and U3317 (N_3317,N_383,N_264);
nand U3318 (N_3318,N_159,N_2052);
nand U3319 (N_3319,N_2270,N_1006);
nand U3320 (N_3320,N_338,N_970);
or U3321 (N_3321,N_1267,N_512);
nand U3322 (N_3322,N_795,N_117);
and U3323 (N_3323,N_1780,N_1279);
and U3324 (N_3324,N_703,N_636);
or U3325 (N_3325,N_519,N_1563);
nand U3326 (N_3326,N_1710,N_220);
nor U3327 (N_3327,N_2103,N_1390);
nor U3328 (N_3328,N_696,N_1867);
and U3329 (N_3329,N_1863,N_1866);
and U3330 (N_3330,N_1272,N_1857);
and U3331 (N_3331,N_1080,N_1957);
nor U3332 (N_3332,N_1052,N_834);
and U3333 (N_3333,N_59,N_1407);
or U3334 (N_3334,N_2071,N_2061);
nor U3335 (N_3335,N_525,N_322);
nor U3336 (N_3336,N_765,N_118);
nor U3337 (N_3337,N_2026,N_467);
nand U3338 (N_3338,N_1711,N_1937);
or U3339 (N_3339,N_2133,N_2255);
xnor U3340 (N_3340,N_2192,N_329);
or U3341 (N_3341,N_2262,N_1495);
nor U3342 (N_3342,N_352,N_1893);
and U3343 (N_3343,N_1352,N_1191);
and U3344 (N_3344,N_1817,N_2374);
or U3345 (N_3345,N_2046,N_2450);
nor U3346 (N_3346,N_1791,N_29);
nor U3347 (N_3347,N_2120,N_305);
or U3348 (N_3348,N_400,N_567);
or U3349 (N_3349,N_633,N_583);
and U3350 (N_3350,N_1035,N_1488);
nor U3351 (N_3351,N_416,N_2439);
xor U3352 (N_3352,N_413,N_1184);
xnor U3353 (N_3353,N_1334,N_1169);
nor U3354 (N_3354,N_1642,N_468);
xor U3355 (N_3355,N_2281,N_1426);
or U3356 (N_3356,N_2104,N_1317);
and U3357 (N_3357,N_2488,N_2053);
and U3358 (N_3358,N_37,N_2342);
nand U3359 (N_3359,N_770,N_2128);
and U3360 (N_3360,N_68,N_451);
nand U3361 (N_3361,N_2320,N_418);
xor U3362 (N_3362,N_466,N_564);
nor U3363 (N_3363,N_820,N_1183);
and U3364 (N_3364,N_2303,N_2065);
nand U3365 (N_3365,N_1675,N_1400);
or U3366 (N_3366,N_878,N_1929);
nand U3367 (N_3367,N_1715,N_389);
nand U3368 (N_3368,N_1950,N_1469);
and U3369 (N_3369,N_2399,N_1109);
or U3370 (N_3370,N_379,N_2433);
and U3371 (N_3371,N_1966,N_572);
or U3372 (N_3372,N_1799,N_397);
and U3373 (N_3373,N_640,N_1539);
or U3374 (N_3374,N_1622,N_592);
nor U3375 (N_3375,N_1885,N_186);
nand U3376 (N_3376,N_1263,N_1946);
and U3377 (N_3377,N_887,N_1786);
and U3378 (N_3378,N_2114,N_217);
and U3379 (N_3379,N_2295,N_1360);
nor U3380 (N_3380,N_1262,N_1882);
and U3381 (N_3381,N_752,N_1418);
or U3382 (N_3382,N_559,N_205);
and U3383 (N_3383,N_1285,N_1087);
or U3384 (N_3384,N_1959,N_2484);
or U3385 (N_3385,N_2124,N_1329);
nand U3386 (N_3386,N_13,N_206);
nand U3387 (N_3387,N_2002,N_1902);
nand U3388 (N_3388,N_2275,N_289);
nand U3389 (N_3389,N_278,N_1039);
and U3390 (N_3390,N_176,N_1401);
nor U3391 (N_3391,N_1252,N_309);
nand U3392 (N_3392,N_1518,N_1530);
and U3393 (N_3393,N_1912,N_1090);
nor U3394 (N_3394,N_94,N_2151);
and U3395 (N_3395,N_183,N_1818);
nor U3396 (N_3396,N_2325,N_1771);
or U3397 (N_3397,N_745,N_704);
or U3398 (N_3398,N_932,N_1331);
and U3399 (N_3399,N_951,N_1773);
xor U3400 (N_3400,N_2049,N_2418);
and U3401 (N_3401,N_998,N_926);
and U3402 (N_3402,N_2073,N_766);
nand U3403 (N_3403,N_1644,N_1122);
nor U3404 (N_3404,N_231,N_757);
or U3405 (N_3405,N_772,N_2042);
nand U3406 (N_3406,N_971,N_1831);
nand U3407 (N_3407,N_761,N_112);
xnor U3408 (N_3408,N_902,N_1198);
or U3409 (N_3409,N_191,N_706);
or U3410 (N_3410,N_988,N_980);
and U3411 (N_3411,N_414,N_230);
or U3412 (N_3412,N_2033,N_1112);
or U3413 (N_3413,N_1013,N_136);
and U3414 (N_3414,N_2220,N_1728);
nor U3415 (N_3415,N_1379,N_1955);
and U3416 (N_3416,N_1638,N_915);
nor U3417 (N_3417,N_2244,N_1993);
nor U3418 (N_3418,N_323,N_2249);
or U3419 (N_3419,N_2269,N_357);
nand U3420 (N_3420,N_337,N_1750);
or U3421 (N_3421,N_1678,N_317);
and U3422 (N_3422,N_551,N_1445);
and U3423 (N_3423,N_1578,N_888);
nor U3424 (N_3424,N_2497,N_1280);
and U3425 (N_3425,N_76,N_1904);
nand U3426 (N_3426,N_2290,N_442);
nor U3427 (N_3427,N_2324,N_375);
or U3428 (N_3428,N_1283,N_425);
nor U3429 (N_3429,N_836,N_2293);
nor U3430 (N_3430,N_494,N_1077);
nor U3431 (N_3431,N_1769,N_2232);
nor U3432 (N_3432,N_2248,N_2204);
nand U3433 (N_3433,N_2296,N_2236);
and U3434 (N_3434,N_2352,N_2056);
nand U3435 (N_3435,N_1346,N_1650);
or U3436 (N_3436,N_1383,N_297);
or U3437 (N_3437,N_458,N_1482);
xor U3438 (N_3438,N_1219,N_2409);
nand U3439 (N_3439,N_1345,N_1545);
or U3440 (N_3440,N_1804,N_2015);
nand U3441 (N_3441,N_339,N_1047);
nor U3442 (N_3442,N_314,N_1410);
nand U3443 (N_3443,N_36,N_688);
or U3444 (N_3444,N_1851,N_1759);
nor U3445 (N_3445,N_1839,N_364);
and U3446 (N_3446,N_2218,N_2188);
or U3447 (N_3447,N_1218,N_1002);
nor U3448 (N_3448,N_2168,N_438);
and U3449 (N_3449,N_846,N_248);
and U3450 (N_3450,N_443,N_556);
or U3451 (N_3451,N_1838,N_1663);
and U3452 (N_3452,N_1554,N_1031);
nand U3453 (N_3453,N_2000,N_986);
or U3454 (N_3454,N_445,N_1130);
or U3455 (N_3455,N_1768,N_1854);
or U3456 (N_3456,N_2390,N_1517);
or U3457 (N_3457,N_747,N_1546);
and U3458 (N_3458,N_842,N_215);
or U3459 (N_3459,N_224,N_411);
xor U3460 (N_3460,N_1449,N_714);
and U3461 (N_3461,N_1939,N_2024);
nor U3462 (N_3462,N_17,N_2001);
and U3463 (N_3463,N_539,N_1236);
nor U3464 (N_3464,N_236,N_1483);
nand U3465 (N_3465,N_1174,N_817);
nor U3466 (N_3466,N_285,N_885);
nand U3467 (N_3467,N_1315,N_177);
or U3468 (N_3468,N_32,N_1665);
or U3469 (N_3469,N_1222,N_1814);
nor U3470 (N_3470,N_503,N_2051);
and U3471 (N_3471,N_2499,N_1306);
nand U3472 (N_3472,N_1559,N_1141);
nor U3473 (N_3473,N_64,N_731);
nor U3474 (N_3474,N_664,N_1504);
nor U3475 (N_3475,N_709,N_2491);
and U3476 (N_3476,N_649,N_1453);
or U3477 (N_3477,N_399,N_1781);
nor U3478 (N_3478,N_1706,N_1624);
nand U3479 (N_3479,N_280,N_424);
and U3480 (N_3480,N_85,N_491);
or U3481 (N_3481,N_1391,N_209);
nor U3482 (N_3482,N_1305,N_2205);
and U3483 (N_3483,N_816,N_286);
or U3484 (N_3484,N_1137,N_1325);
xor U3485 (N_3485,N_1987,N_1129);
and U3486 (N_3486,N_1733,N_1097);
and U3487 (N_3487,N_676,N_469);
or U3488 (N_3488,N_615,N_151);
and U3489 (N_3489,N_2094,N_1199);
or U3490 (N_3490,N_1670,N_320);
nand U3491 (N_3491,N_910,N_550);
nand U3492 (N_3492,N_788,N_1343);
nor U3493 (N_3493,N_74,N_1763);
nor U3494 (N_3494,N_1721,N_1566);
xnor U3495 (N_3495,N_2311,N_710);
and U3496 (N_3496,N_2012,N_336);
xnor U3497 (N_3497,N_784,N_2067);
nand U3498 (N_3498,N_669,N_966);
xnor U3499 (N_3499,N_1248,N_2403);
and U3500 (N_3500,N_2210,N_1227);
xor U3501 (N_3501,N_200,N_2111);
nand U3502 (N_3502,N_2118,N_2182);
nor U3503 (N_3503,N_1649,N_865);
or U3504 (N_3504,N_2138,N_798);
nor U3505 (N_3505,N_1911,N_1339);
and U3506 (N_3506,N_1619,N_2479);
and U3507 (N_3507,N_1850,N_822);
or U3508 (N_3508,N_1956,N_1999);
nor U3509 (N_3509,N_1537,N_607);
nand U3510 (N_3510,N_1499,N_946);
nand U3511 (N_3511,N_1072,N_1060);
nor U3512 (N_3512,N_1871,N_992);
and U3513 (N_3513,N_2064,N_54);
nor U3514 (N_3514,N_1886,N_2375);
nor U3515 (N_3515,N_1878,N_1884);
nand U3516 (N_3516,N_544,N_429);
or U3517 (N_3517,N_1844,N_212);
or U3518 (N_3518,N_1813,N_362);
and U3519 (N_3519,N_1901,N_175);
and U3520 (N_3520,N_2154,N_2121);
nand U3521 (N_3521,N_1980,N_1200);
or U3522 (N_3522,N_119,N_2487);
and U3523 (N_3523,N_169,N_641);
and U3524 (N_3524,N_2099,N_2412);
and U3525 (N_3525,N_1764,N_1845);
nor U3526 (N_3526,N_2224,N_240);
xnor U3527 (N_3527,N_1679,N_2171);
or U3528 (N_3528,N_139,N_1136);
nand U3529 (N_3529,N_225,N_2329);
nand U3530 (N_3530,N_1021,N_235);
and U3531 (N_3531,N_2431,N_195);
and U3532 (N_3532,N_1075,N_58);
nor U3533 (N_3533,N_659,N_2112);
nor U3534 (N_3534,N_1440,N_1732);
or U3535 (N_3535,N_2122,N_1837);
and U3536 (N_3536,N_1127,N_838);
nor U3537 (N_3537,N_1538,N_49);
or U3538 (N_3538,N_1605,N_1756);
or U3539 (N_3539,N_1394,N_1890);
xnor U3540 (N_3540,N_2291,N_1004);
nor U3541 (N_3541,N_2088,N_1357);
nor U3542 (N_3542,N_1676,N_2394);
xnor U3543 (N_3543,N_1958,N_2158);
nand U3544 (N_3544,N_1960,N_1058);
nand U3545 (N_3545,N_2072,N_1373);
nand U3546 (N_3546,N_500,N_1776);
or U3547 (N_3547,N_2243,N_1490);
or U3548 (N_3548,N_284,N_1020);
nor U3549 (N_3549,N_1681,N_2434);
and U3550 (N_3550,N_1570,N_1931);
or U3551 (N_3551,N_1627,N_1954);
and U3552 (N_3552,N_330,N_4);
nand U3553 (N_3553,N_274,N_1824);
nor U3554 (N_3554,N_1577,N_673);
xnor U3555 (N_3555,N_372,N_1318);
and U3556 (N_3556,N_2441,N_2139);
and U3557 (N_3557,N_81,N_1973);
nand U3558 (N_3558,N_963,N_91);
and U3559 (N_3559,N_1450,N_644);
nor U3560 (N_3560,N_1460,N_1428);
or U3561 (N_3561,N_1631,N_1620);
or U3562 (N_3562,N_1327,N_2469);
nor U3563 (N_3563,N_1916,N_2148);
or U3564 (N_3564,N_291,N_234);
xor U3565 (N_3565,N_1050,N_558);
nor U3566 (N_3566,N_922,N_678);
nor U3567 (N_3567,N_33,N_916);
and U3568 (N_3568,N_1513,N_2490);
nor U3569 (N_3569,N_1616,N_2271);
and U3570 (N_3570,N_84,N_311);
xnor U3571 (N_3571,N_146,N_609);
or U3572 (N_3572,N_1585,N_2282);
and U3573 (N_3573,N_2459,N_1467);
nor U3574 (N_3574,N_2400,N_2415);
nand U3575 (N_3575,N_461,N_1505);
nor U3576 (N_3576,N_1628,N_482);
or U3577 (N_3577,N_1592,N_450);
xor U3578 (N_3578,N_2429,N_189);
and U3579 (N_3579,N_517,N_2105);
nand U3580 (N_3580,N_12,N_2388);
and U3581 (N_3581,N_738,N_1834);
nand U3582 (N_3582,N_601,N_1985);
nor U3583 (N_3583,N_1610,N_540);
nand U3584 (N_3584,N_1273,N_2025);
or U3585 (N_3585,N_854,N_1755);
and U3586 (N_3586,N_403,N_1508);
nand U3587 (N_3587,N_1827,N_1308);
and U3588 (N_3588,N_1994,N_2129);
or U3589 (N_3589,N_2239,N_949);
and U3590 (N_3590,N_1829,N_1898);
nand U3591 (N_3591,N_2044,N_1798);
nand U3592 (N_3592,N_1027,N_216);
nor U3593 (N_3593,N_1671,N_1541);
and U3594 (N_3594,N_3,N_504);
or U3595 (N_3595,N_475,N_1618);
and U3596 (N_3596,N_686,N_735);
and U3597 (N_3597,N_1085,N_1107);
and U3598 (N_3598,N_1826,N_65);
xnor U3599 (N_3599,N_1982,N_2197);
and U3600 (N_3600,N_2233,N_577);
nor U3601 (N_3601,N_1384,N_261);
and U3602 (N_3602,N_2261,N_1772);
or U3603 (N_3603,N_181,N_1840);
nand U3604 (N_3604,N_730,N_2326);
or U3605 (N_3605,N_1708,N_2483);
nand U3606 (N_3606,N_728,N_1790);
or U3607 (N_3607,N_1078,N_876);
xnor U3608 (N_3608,N_1012,N_1589);
nand U3609 (N_3609,N_814,N_1310);
or U3610 (N_3610,N_976,N_133);
nor U3611 (N_3611,N_1695,N_2219);
nor U3612 (N_3612,N_2101,N_2404);
and U3613 (N_3613,N_1354,N_2140);
nand U3614 (N_3614,N_573,N_793);
nand U3615 (N_3615,N_1569,N_657);
nand U3616 (N_3616,N_130,N_86);
nor U3617 (N_3617,N_1451,N_19);
and U3618 (N_3618,N_2251,N_385);
xor U3619 (N_3619,N_1607,N_2286);
and U3620 (N_3620,N_597,N_574);
nand U3621 (N_3621,N_1881,N_1030);
nand U3622 (N_3622,N_1707,N_1079);
and U3623 (N_3623,N_2144,N_1797);
xnor U3624 (N_3624,N_2420,N_2370);
and U3625 (N_3625,N_2347,N_1412);
and U3626 (N_3626,N_407,N_1201);
nor U3627 (N_3627,N_2108,N_1142);
nor U3628 (N_3628,N_345,N_1677);
or U3629 (N_3629,N_857,N_57);
nand U3630 (N_3630,N_670,N_2206);
or U3631 (N_3631,N_2162,N_955);
xnor U3632 (N_3632,N_1509,N_2278);
nand U3633 (N_3633,N_2,N_1478);
or U3634 (N_3634,N_1380,N_2126);
nand U3635 (N_3635,N_303,N_377);
and U3636 (N_3636,N_1761,N_2005);
nand U3637 (N_3637,N_115,N_810);
nand U3638 (N_3638,N_1493,N_1533);
nand U3639 (N_3639,N_1064,N_1748);
nor U3640 (N_3640,N_2102,N_412);
or U3641 (N_3641,N_744,N_2208);
nand U3642 (N_3642,N_395,N_1120);
and U3643 (N_3643,N_1211,N_2050);
xnor U3644 (N_3644,N_219,N_1311);
nand U3645 (N_3645,N_46,N_2090);
and U3646 (N_3646,N_1498,N_2028);
or U3647 (N_3647,N_1111,N_1637);
and U3648 (N_3648,N_381,N_2357);
nor U3649 (N_3649,N_1427,N_1630);
nand U3650 (N_3650,N_1011,N_1612);
or U3651 (N_3651,N_1590,N_1149);
nand U3652 (N_3652,N_499,N_978);
or U3653 (N_3653,N_758,N_2170);
or U3654 (N_3654,N_1472,N_162);
or U3655 (N_3655,N_241,N_603);
xnor U3656 (N_3656,N_1303,N_809);
nor U3657 (N_3657,N_1582,N_1150);
nor U3658 (N_3658,N_535,N_2480);
and U3659 (N_3659,N_1459,N_1250);
or U3660 (N_3660,N_290,N_1119);
nand U3661 (N_3661,N_792,N_1634);
nor U3662 (N_3662,N_1044,N_1775);
xor U3663 (N_3663,N_2074,N_1625);
nor U3664 (N_3664,N_34,N_1489);
or U3665 (N_3665,N_1045,N_1233);
nor U3666 (N_3666,N_1873,N_1161);
nor U3667 (N_3667,N_111,N_1172);
xor U3668 (N_3668,N_1501,N_863);
or U3669 (N_3669,N_1337,N_1894);
and U3670 (N_3670,N_1550,N_895);
and U3671 (N_3671,N_456,N_354);
nand U3672 (N_3672,N_695,N_1260);
and U3673 (N_3673,N_1411,N_2481);
nand U3674 (N_3674,N_527,N_1386);
or U3675 (N_3675,N_137,N_2359);
xor U3676 (N_3676,N_1074,N_2339);
nor U3677 (N_3677,N_1787,N_2407);
and U3678 (N_3678,N_1500,N_1815);
xnor U3679 (N_3679,N_1758,N_1828);
and U3680 (N_3680,N_666,N_2308);
xnor U3681 (N_3681,N_243,N_2276);
or U3682 (N_3682,N_2079,N_204);
or U3683 (N_3683,N_605,N_1647);
xor U3684 (N_3684,N_725,N_444);
nor U3685 (N_3685,N_18,N_510);
or U3686 (N_3686,N_866,N_1540);
and U3687 (N_3687,N_1135,N_300);
nor U3688 (N_3688,N_1264,N_265);
xor U3689 (N_3689,N_164,N_2301);
nand U3690 (N_3690,N_2389,N_914);
and U3691 (N_3691,N_1558,N_2075);
nand U3692 (N_3692,N_1037,N_1888);
and U3693 (N_3693,N_78,N_2285);
nand U3694 (N_3694,N_40,N_1547);
and U3695 (N_3695,N_121,N_260);
nand U3696 (N_3696,N_365,N_197);
xnor U3697 (N_3697,N_2466,N_1091);
xnor U3698 (N_3698,N_2007,N_1372);
or U3699 (N_3699,N_697,N_1964);
xnor U3700 (N_3700,N_760,N_1148);
nor U3701 (N_3701,N_1221,N_560);
or U3702 (N_3702,N_1462,N_652);
nor U3703 (N_3703,N_868,N_73);
nand U3704 (N_3704,N_1988,N_1717);
and U3705 (N_3705,N_2432,N_1914);
nor U3706 (N_3706,N_620,N_1688);
nand U3707 (N_3707,N_1335,N_799);
nor U3708 (N_3708,N_406,N_1602);
nand U3709 (N_3709,N_51,N_575);
nand U3710 (N_3710,N_1583,N_2332);
nor U3711 (N_3711,N_287,N_2020);
nand U3712 (N_3712,N_346,N_1986);
or U3713 (N_3713,N_844,N_1595);
nor U3714 (N_3714,N_2043,N_2066);
nor U3715 (N_3715,N_961,N_144);
xor U3716 (N_3716,N_896,N_513);
or U3717 (N_3717,N_803,N_737);
or U3718 (N_3718,N_1887,N_1603);
nor U3719 (N_3719,N_432,N_1918);
nor U3720 (N_3720,N_2471,N_2221);
or U3721 (N_3721,N_366,N_1497);
nand U3722 (N_3722,N_2336,N_1475);
nand U3723 (N_3723,N_632,N_701);
nand U3724 (N_3724,N_2452,N_1230);
xor U3725 (N_3725,N_954,N_796);
nand U3726 (N_3726,N_296,N_478);
nand U3727 (N_3727,N_684,N_1496);
nand U3728 (N_3728,N_859,N_1242);
nor U3729 (N_3729,N_646,N_518);
nand U3730 (N_3730,N_1232,N_1213);
or U3731 (N_3731,N_1953,N_44);
nor U3732 (N_3732,N_61,N_90);
xnor U3733 (N_3733,N_872,N_1294);
nand U3734 (N_3734,N_2186,N_2402);
xor U3735 (N_3735,N_307,N_1225);
and U3736 (N_3736,N_394,N_1783);
nand U3737 (N_3737,N_332,N_454);
or U3738 (N_3738,N_304,N_75);
nand U3739 (N_3739,N_665,N_1639);
nor U3740 (N_3740,N_1128,N_1131);
nand U3741 (N_3741,N_781,N_355);
or U3742 (N_3742,N_634,N_1298);
or U3743 (N_3743,N_2331,N_239);
nand U3744 (N_3744,N_1163,N_0);
and U3745 (N_3745,N_749,N_22);
nand U3746 (N_3746,N_1526,N_1542);
nand U3747 (N_3747,N_1196,N_2333);
and U3748 (N_3748,N_937,N_1231);
or U3749 (N_3749,N_1626,N_1134);
nor U3750 (N_3750,N_699,N_608);
and U3751 (N_3751,N_712,N_245);
xnor U3752 (N_3752,N_2005,N_1566);
or U3753 (N_3753,N_185,N_1513);
xnor U3754 (N_3754,N_994,N_518);
nand U3755 (N_3755,N_1447,N_1472);
nand U3756 (N_3756,N_2253,N_1112);
xor U3757 (N_3757,N_1529,N_1600);
or U3758 (N_3758,N_1131,N_2444);
nand U3759 (N_3759,N_96,N_1478);
xnor U3760 (N_3760,N_2135,N_614);
or U3761 (N_3761,N_2294,N_2412);
or U3762 (N_3762,N_1177,N_1870);
nor U3763 (N_3763,N_1221,N_1618);
and U3764 (N_3764,N_1892,N_2425);
nor U3765 (N_3765,N_2430,N_1689);
nor U3766 (N_3766,N_736,N_2465);
nor U3767 (N_3767,N_1998,N_579);
nor U3768 (N_3768,N_1149,N_1434);
and U3769 (N_3769,N_1815,N_944);
nand U3770 (N_3770,N_727,N_2094);
and U3771 (N_3771,N_1264,N_2017);
and U3772 (N_3772,N_857,N_544);
xnor U3773 (N_3773,N_753,N_1979);
and U3774 (N_3774,N_478,N_518);
or U3775 (N_3775,N_1371,N_813);
nor U3776 (N_3776,N_313,N_654);
nand U3777 (N_3777,N_1633,N_391);
nor U3778 (N_3778,N_1293,N_1565);
and U3779 (N_3779,N_1018,N_2434);
nand U3780 (N_3780,N_994,N_2425);
or U3781 (N_3781,N_539,N_2367);
xnor U3782 (N_3782,N_2359,N_927);
xnor U3783 (N_3783,N_1012,N_1363);
or U3784 (N_3784,N_1242,N_474);
nor U3785 (N_3785,N_1965,N_2326);
nor U3786 (N_3786,N_2122,N_2031);
nand U3787 (N_3787,N_795,N_816);
nor U3788 (N_3788,N_434,N_1218);
and U3789 (N_3789,N_489,N_2418);
nor U3790 (N_3790,N_683,N_2483);
and U3791 (N_3791,N_762,N_481);
and U3792 (N_3792,N_2230,N_2227);
and U3793 (N_3793,N_2408,N_1026);
or U3794 (N_3794,N_2347,N_828);
or U3795 (N_3795,N_2213,N_1792);
or U3796 (N_3796,N_672,N_765);
nand U3797 (N_3797,N_603,N_1118);
or U3798 (N_3798,N_37,N_1208);
xnor U3799 (N_3799,N_1721,N_951);
nand U3800 (N_3800,N_2311,N_2400);
and U3801 (N_3801,N_2145,N_166);
nand U3802 (N_3802,N_917,N_401);
xnor U3803 (N_3803,N_692,N_1423);
xnor U3804 (N_3804,N_572,N_1040);
xor U3805 (N_3805,N_2169,N_2222);
or U3806 (N_3806,N_467,N_1068);
nor U3807 (N_3807,N_78,N_242);
or U3808 (N_3808,N_1637,N_191);
xnor U3809 (N_3809,N_229,N_2252);
or U3810 (N_3810,N_1886,N_815);
and U3811 (N_3811,N_1670,N_756);
nor U3812 (N_3812,N_257,N_1135);
nand U3813 (N_3813,N_869,N_1151);
or U3814 (N_3814,N_210,N_895);
or U3815 (N_3815,N_2307,N_1289);
nor U3816 (N_3816,N_1489,N_853);
nor U3817 (N_3817,N_1162,N_500);
nand U3818 (N_3818,N_232,N_238);
and U3819 (N_3819,N_2217,N_929);
nand U3820 (N_3820,N_1851,N_1626);
and U3821 (N_3821,N_2238,N_565);
nor U3822 (N_3822,N_1742,N_921);
nor U3823 (N_3823,N_268,N_1914);
nor U3824 (N_3824,N_919,N_1934);
and U3825 (N_3825,N_1033,N_1063);
nand U3826 (N_3826,N_2043,N_217);
xor U3827 (N_3827,N_2288,N_108);
nor U3828 (N_3828,N_2233,N_2180);
nor U3829 (N_3829,N_1112,N_2151);
and U3830 (N_3830,N_1704,N_1037);
nor U3831 (N_3831,N_65,N_898);
nor U3832 (N_3832,N_555,N_1745);
nand U3833 (N_3833,N_2260,N_775);
nand U3834 (N_3834,N_1245,N_2088);
and U3835 (N_3835,N_974,N_1983);
or U3836 (N_3836,N_1099,N_883);
xor U3837 (N_3837,N_1648,N_1831);
or U3838 (N_3838,N_417,N_1650);
and U3839 (N_3839,N_627,N_818);
nand U3840 (N_3840,N_287,N_584);
xnor U3841 (N_3841,N_2100,N_2153);
xnor U3842 (N_3842,N_2346,N_1037);
and U3843 (N_3843,N_1853,N_1071);
nor U3844 (N_3844,N_2208,N_1922);
and U3845 (N_3845,N_2329,N_1148);
nand U3846 (N_3846,N_832,N_736);
and U3847 (N_3847,N_1039,N_368);
nor U3848 (N_3848,N_123,N_1524);
or U3849 (N_3849,N_1590,N_1847);
or U3850 (N_3850,N_160,N_535);
or U3851 (N_3851,N_1713,N_1839);
nor U3852 (N_3852,N_677,N_2147);
nor U3853 (N_3853,N_2070,N_429);
and U3854 (N_3854,N_1745,N_996);
and U3855 (N_3855,N_1546,N_2365);
or U3856 (N_3856,N_58,N_486);
or U3857 (N_3857,N_720,N_1705);
nor U3858 (N_3858,N_1635,N_2312);
xor U3859 (N_3859,N_129,N_1129);
xnor U3860 (N_3860,N_1338,N_1407);
and U3861 (N_3861,N_1980,N_1326);
or U3862 (N_3862,N_798,N_2026);
nor U3863 (N_3863,N_135,N_126);
or U3864 (N_3864,N_1192,N_705);
and U3865 (N_3865,N_1022,N_1396);
and U3866 (N_3866,N_1065,N_1503);
xor U3867 (N_3867,N_1851,N_1294);
nand U3868 (N_3868,N_1038,N_423);
nand U3869 (N_3869,N_2080,N_1879);
and U3870 (N_3870,N_1252,N_333);
nand U3871 (N_3871,N_2435,N_258);
nor U3872 (N_3872,N_330,N_1429);
nor U3873 (N_3873,N_1067,N_159);
nor U3874 (N_3874,N_1028,N_809);
nor U3875 (N_3875,N_859,N_814);
and U3876 (N_3876,N_229,N_929);
xnor U3877 (N_3877,N_844,N_657);
nand U3878 (N_3878,N_36,N_2246);
nor U3879 (N_3879,N_1178,N_1508);
nor U3880 (N_3880,N_2046,N_2289);
nor U3881 (N_3881,N_701,N_1704);
nor U3882 (N_3882,N_933,N_1610);
nor U3883 (N_3883,N_1106,N_1195);
nor U3884 (N_3884,N_1138,N_19);
xor U3885 (N_3885,N_208,N_2111);
or U3886 (N_3886,N_197,N_347);
nand U3887 (N_3887,N_247,N_2260);
or U3888 (N_3888,N_264,N_1121);
nor U3889 (N_3889,N_1218,N_1283);
xor U3890 (N_3890,N_293,N_1897);
and U3891 (N_3891,N_435,N_1382);
xnor U3892 (N_3892,N_388,N_1178);
nand U3893 (N_3893,N_535,N_1973);
nor U3894 (N_3894,N_2332,N_107);
or U3895 (N_3895,N_525,N_1717);
and U3896 (N_3896,N_54,N_149);
nand U3897 (N_3897,N_488,N_364);
nor U3898 (N_3898,N_1423,N_674);
and U3899 (N_3899,N_2109,N_1194);
or U3900 (N_3900,N_642,N_219);
or U3901 (N_3901,N_499,N_425);
and U3902 (N_3902,N_761,N_1027);
xor U3903 (N_3903,N_2230,N_711);
and U3904 (N_3904,N_1347,N_1486);
nand U3905 (N_3905,N_57,N_204);
nor U3906 (N_3906,N_1497,N_2490);
nand U3907 (N_3907,N_1107,N_1604);
or U3908 (N_3908,N_2215,N_1485);
nor U3909 (N_3909,N_1537,N_237);
nand U3910 (N_3910,N_1004,N_173);
nand U3911 (N_3911,N_2131,N_2006);
and U3912 (N_3912,N_1601,N_1235);
nor U3913 (N_3913,N_29,N_1860);
nand U3914 (N_3914,N_552,N_515);
and U3915 (N_3915,N_1346,N_539);
and U3916 (N_3916,N_942,N_811);
and U3917 (N_3917,N_1394,N_1406);
and U3918 (N_3918,N_1191,N_2254);
nand U3919 (N_3919,N_2386,N_2084);
or U3920 (N_3920,N_366,N_606);
or U3921 (N_3921,N_2119,N_604);
nor U3922 (N_3922,N_2491,N_475);
or U3923 (N_3923,N_520,N_1967);
nor U3924 (N_3924,N_1849,N_1672);
and U3925 (N_3925,N_1877,N_993);
or U3926 (N_3926,N_350,N_2084);
nand U3927 (N_3927,N_2319,N_1602);
or U3928 (N_3928,N_2453,N_83);
or U3929 (N_3929,N_2323,N_1776);
and U3930 (N_3930,N_695,N_1783);
nand U3931 (N_3931,N_122,N_1496);
and U3932 (N_3932,N_960,N_1155);
nor U3933 (N_3933,N_1888,N_1579);
or U3934 (N_3934,N_1745,N_873);
or U3935 (N_3935,N_919,N_1896);
nor U3936 (N_3936,N_270,N_437);
nand U3937 (N_3937,N_955,N_1372);
nor U3938 (N_3938,N_1263,N_2275);
nand U3939 (N_3939,N_578,N_1134);
nor U3940 (N_3940,N_1721,N_104);
or U3941 (N_3941,N_956,N_1172);
nand U3942 (N_3942,N_1712,N_146);
and U3943 (N_3943,N_504,N_1537);
nand U3944 (N_3944,N_1608,N_952);
or U3945 (N_3945,N_317,N_775);
and U3946 (N_3946,N_1092,N_1980);
or U3947 (N_3947,N_401,N_604);
nor U3948 (N_3948,N_2218,N_343);
xor U3949 (N_3949,N_1569,N_1123);
xnor U3950 (N_3950,N_1606,N_412);
or U3951 (N_3951,N_2349,N_1596);
nand U3952 (N_3952,N_510,N_2357);
nand U3953 (N_3953,N_134,N_1255);
nand U3954 (N_3954,N_672,N_1159);
nand U3955 (N_3955,N_614,N_2016);
or U3956 (N_3956,N_560,N_493);
and U3957 (N_3957,N_954,N_1192);
nand U3958 (N_3958,N_803,N_1332);
or U3959 (N_3959,N_609,N_1369);
and U3960 (N_3960,N_1708,N_1192);
or U3961 (N_3961,N_1235,N_953);
xor U3962 (N_3962,N_93,N_54);
xnor U3963 (N_3963,N_2150,N_2050);
nand U3964 (N_3964,N_990,N_1792);
nand U3965 (N_3965,N_242,N_2155);
nor U3966 (N_3966,N_214,N_893);
or U3967 (N_3967,N_349,N_267);
or U3968 (N_3968,N_24,N_1120);
and U3969 (N_3969,N_1037,N_2);
and U3970 (N_3970,N_470,N_886);
nand U3971 (N_3971,N_1326,N_525);
nor U3972 (N_3972,N_555,N_2127);
and U3973 (N_3973,N_2227,N_1360);
and U3974 (N_3974,N_1075,N_2096);
or U3975 (N_3975,N_2191,N_2413);
xnor U3976 (N_3976,N_238,N_1293);
nor U3977 (N_3977,N_410,N_245);
or U3978 (N_3978,N_1640,N_2469);
nand U3979 (N_3979,N_1998,N_1614);
and U3980 (N_3980,N_1989,N_475);
nand U3981 (N_3981,N_1906,N_65);
and U3982 (N_3982,N_2279,N_2102);
nand U3983 (N_3983,N_1554,N_221);
or U3984 (N_3984,N_70,N_282);
nor U3985 (N_3985,N_2023,N_2258);
nand U3986 (N_3986,N_323,N_1524);
nand U3987 (N_3987,N_2080,N_2409);
nor U3988 (N_3988,N_491,N_405);
or U3989 (N_3989,N_1035,N_841);
xnor U3990 (N_3990,N_1011,N_577);
nor U3991 (N_3991,N_616,N_1545);
or U3992 (N_3992,N_1386,N_1132);
nor U3993 (N_3993,N_630,N_734);
nor U3994 (N_3994,N_2114,N_2199);
or U3995 (N_3995,N_1757,N_1916);
nand U3996 (N_3996,N_2044,N_271);
nor U3997 (N_3997,N_393,N_1974);
and U3998 (N_3998,N_1189,N_1907);
and U3999 (N_3999,N_1781,N_1185);
nand U4000 (N_4000,N_891,N_1924);
nand U4001 (N_4001,N_1686,N_1745);
or U4002 (N_4002,N_1182,N_1927);
and U4003 (N_4003,N_589,N_2124);
nor U4004 (N_4004,N_780,N_1257);
and U4005 (N_4005,N_856,N_891);
nand U4006 (N_4006,N_1790,N_973);
nor U4007 (N_4007,N_586,N_885);
nor U4008 (N_4008,N_418,N_2114);
or U4009 (N_4009,N_1818,N_235);
and U4010 (N_4010,N_52,N_2123);
nand U4011 (N_4011,N_1457,N_891);
nand U4012 (N_4012,N_1585,N_2359);
and U4013 (N_4013,N_1836,N_718);
nand U4014 (N_4014,N_853,N_294);
nand U4015 (N_4015,N_399,N_448);
xnor U4016 (N_4016,N_2444,N_2347);
xor U4017 (N_4017,N_1742,N_1035);
xor U4018 (N_4018,N_582,N_1832);
or U4019 (N_4019,N_1783,N_2028);
or U4020 (N_4020,N_1221,N_588);
and U4021 (N_4021,N_171,N_305);
and U4022 (N_4022,N_190,N_1824);
and U4023 (N_4023,N_1347,N_427);
nand U4024 (N_4024,N_1617,N_1306);
or U4025 (N_4025,N_1954,N_1951);
xor U4026 (N_4026,N_1322,N_917);
or U4027 (N_4027,N_538,N_1539);
or U4028 (N_4028,N_1517,N_1478);
or U4029 (N_4029,N_433,N_420);
nand U4030 (N_4030,N_1506,N_2225);
or U4031 (N_4031,N_376,N_586);
and U4032 (N_4032,N_1305,N_1059);
and U4033 (N_4033,N_924,N_1394);
or U4034 (N_4034,N_2209,N_1046);
nand U4035 (N_4035,N_1650,N_94);
and U4036 (N_4036,N_1432,N_96);
nand U4037 (N_4037,N_2328,N_1798);
nor U4038 (N_4038,N_2250,N_731);
or U4039 (N_4039,N_2284,N_1606);
nor U4040 (N_4040,N_164,N_1092);
nand U4041 (N_4041,N_1850,N_1043);
and U4042 (N_4042,N_1098,N_537);
nand U4043 (N_4043,N_733,N_20);
and U4044 (N_4044,N_1366,N_841);
nand U4045 (N_4045,N_2489,N_2324);
nor U4046 (N_4046,N_414,N_359);
nand U4047 (N_4047,N_851,N_113);
nor U4048 (N_4048,N_1264,N_321);
nand U4049 (N_4049,N_2385,N_165);
nand U4050 (N_4050,N_179,N_246);
or U4051 (N_4051,N_62,N_2007);
nand U4052 (N_4052,N_398,N_790);
or U4053 (N_4053,N_844,N_1448);
and U4054 (N_4054,N_840,N_963);
nor U4055 (N_4055,N_437,N_830);
or U4056 (N_4056,N_1120,N_899);
nor U4057 (N_4057,N_2441,N_1830);
or U4058 (N_4058,N_1978,N_687);
nor U4059 (N_4059,N_1128,N_250);
or U4060 (N_4060,N_301,N_4);
and U4061 (N_4061,N_1788,N_1545);
and U4062 (N_4062,N_1275,N_440);
or U4063 (N_4063,N_1124,N_1388);
nand U4064 (N_4064,N_1592,N_989);
or U4065 (N_4065,N_1676,N_2482);
or U4066 (N_4066,N_1193,N_2007);
nand U4067 (N_4067,N_1737,N_100);
xor U4068 (N_4068,N_71,N_387);
or U4069 (N_4069,N_1512,N_1738);
nor U4070 (N_4070,N_2134,N_1446);
xor U4071 (N_4071,N_2491,N_970);
nor U4072 (N_4072,N_890,N_887);
and U4073 (N_4073,N_1422,N_670);
and U4074 (N_4074,N_1302,N_2294);
nor U4075 (N_4075,N_2460,N_2255);
nand U4076 (N_4076,N_2171,N_807);
nor U4077 (N_4077,N_2055,N_1099);
xor U4078 (N_4078,N_1119,N_1300);
and U4079 (N_4079,N_1492,N_312);
or U4080 (N_4080,N_1417,N_2210);
or U4081 (N_4081,N_533,N_0);
xnor U4082 (N_4082,N_385,N_1691);
or U4083 (N_4083,N_367,N_1375);
or U4084 (N_4084,N_1653,N_1264);
nand U4085 (N_4085,N_2265,N_2258);
nor U4086 (N_4086,N_195,N_916);
and U4087 (N_4087,N_2221,N_1276);
nand U4088 (N_4088,N_730,N_796);
and U4089 (N_4089,N_156,N_956);
xor U4090 (N_4090,N_549,N_2438);
or U4091 (N_4091,N_1405,N_1343);
or U4092 (N_4092,N_797,N_513);
nand U4093 (N_4093,N_2246,N_301);
or U4094 (N_4094,N_1340,N_599);
xor U4095 (N_4095,N_1941,N_377);
or U4096 (N_4096,N_2019,N_1173);
and U4097 (N_4097,N_652,N_53);
and U4098 (N_4098,N_1465,N_1181);
nand U4099 (N_4099,N_447,N_133);
nand U4100 (N_4100,N_1122,N_632);
or U4101 (N_4101,N_1729,N_499);
or U4102 (N_4102,N_804,N_1087);
or U4103 (N_4103,N_891,N_1319);
xnor U4104 (N_4104,N_330,N_2282);
nor U4105 (N_4105,N_1842,N_2068);
and U4106 (N_4106,N_752,N_372);
nor U4107 (N_4107,N_354,N_450);
and U4108 (N_4108,N_814,N_529);
and U4109 (N_4109,N_1186,N_1565);
or U4110 (N_4110,N_1287,N_1033);
xnor U4111 (N_4111,N_1477,N_1012);
xor U4112 (N_4112,N_1157,N_1048);
and U4113 (N_4113,N_1903,N_2315);
nor U4114 (N_4114,N_186,N_2291);
nand U4115 (N_4115,N_689,N_2317);
nand U4116 (N_4116,N_40,N_959);
nor U4117 (N_4117,N_1998,N_1805);
xnor U4118 (N_4118,N_55,N_1907);
and U4119 (N_4119,N_1130,N_987);
nor U4120 (N_4120,N_1318,N_263);
and U4121 (N_4121,N_1259,N_1506);
nor U4122 (N_4122,N_1458,N_231);
or U4123 (N_4123,N_1325,N_1503);
and U4124 (N_4124,N_270,N_1487);
nand U4125 (N_4125,N_668,N_1188);
nor U4126 (N_4126,N_2059,N_533);
nand U4127 (N_4127,N_665,N_2405);
xnor U4128 (N_4128,N_521,N_1729);
nor U4129 (N_4129,N_55,N_1632);
xor U4130 (N_4130,N_2209,N_1847);
or U4131 (N_4131,N_1892,N_496);
or U4132 (N_4132,N_209,N_1234);
nand U4133 (N_4133,N_343,N_420);
nor U4134 (N_4134,N_1109,N_385);
or U4135 (N_4135,N_503,N_1256);
and U4136 (N_4136,N_801,N_2211);
and U4137 (N_4137,N_1520,N_2092);
or U4138 (N_4138,N_1046,N_121);
xor U4139 (N_4139,N_1140,N_1176);
nor U4140 (N_4140,N_301,N_418);
and U4141 (N_4141,N_608,N_693);
nand U4142 (N_4142,N_2041,N_1655);
or U4143 (N_4143,N_2457,N_1535);
and U4144 (N_4144,N_220,N_2432);
nor U4145 (N_4145,N_645,N_229);
and U4146 (N_4146,N_558,N_1348);
nand U4147 (N_4147,N_2004,N_592);
or U4148 (N_4148,N_2077,N_687);
or U4149 (N_4149,N_1237,N_1607);
nand U4150 (N_4150,N_2301,N_1879);
or U4151 (N_4151,N_2298,N_663);
and U4152 (N_4152,N_2042,N_1327);
or U4153 (N_4153,N_701,N_305);
or U4154 (N_4154,N_377,N_899);
nor U4155 (N_4155,N_889,N_524);
and U4156 (N_4156,N_2167,N_648);
or U4157 (N_4157,N_2409,N_976);
or U4158 (N_4158,N_2323,N_1335);
nand U4159 (N_4159,N_819,N_632);
nor U4160 (N_4160,N_1230,N_1623);
nand U4161 (N_4161,N_1405,N_2113);
nand U4162 (N_4162,N_1411,N_1279);
or U4163 (N_4163,N_2185,N_2241);
nor U4164 (N_4164,N_72,N_987);
xnor U4165 (N_4165,N_978,N_1568);
or U4166 (N_4166,N_1089,N_1653);
or U4167 (N_4167,N_1180,N_702);
or U4168 (N_4168,N_1864,N_645);
and U4169 (N_4169,N_1165,N_160);
and U4170 (N_4170,N_638,N_1595);
and U4171 (N_4171,N_1165,N_2331);
nor U4172 (N_4172,N_1822,N_2090);
xnor U4173 (N_4173,N_1013,N_1289);
xnor U4174 (N_4174,N_592,N_2370);
nor U4175 (N_4175,N_1465,N_2183);
nor U4176 (N_4176,N_894,N_1462);
or U4177 (N_4177,N_227,N_2184);
nand U4178 (N_4178,N_1657,N_158);
or U4179 (N_4179,N_114,N_868);
nor U4180 (N_4180,N_1295,N_596);
and U4181 (N_4181,N_969,N_977);
and U4182 (N_4182,N_1116,N_691);
nand U4183 (N_4183,N_221,N_1888);
nor U4184 (N_4184,N_2073,N_1752);
nand U4185 (N_4185,N_2305,N_904);
nand U4186 (N_4186,N_2173,N_1125);
nor U4187 (N_4187,N_1611,N_1829);
xor U4188 (N_4188,N_1057,N_1563);
nor U4189 (N_4189,N_799,N_1128);
xnor U4190 (N_4190,N_461,N_2277);
nand U4191 (N_4191,N_243,N_704);
or U4192 (N_4192,N_1415,N_1562);
or U4193 (N_4193,N_1548,N_230);
or U4194 (N_4194,N_314,N_2037);
or U4195 (N_4195,N_1038,N_1282);
or U4196 (N_4196,N_943,N_999);
nor U4197 (N_4197,N_1993,N_65);
and U4198 (N_4198,N_1854,N_529);
nor U4199 (N_4199,N_2321,N_2196);
or U4200 (N_4200,N_390,N_1701);
nor U4201 (N_4201,N_1260,N_1037);
nor U4202 (N_4202,N_280,N_989);
nand U4203 (N_4203,N_1209,N_2317);
nor U4204 (N_4204,N_1936,N_542);
or U4205 (N_4205,N_312,N_2437);
and U4206 (N_4206,N_1992,N_451);
nor U4207 (N_4207,N_547,N_546);
or U4208 (N_4208,N_1156,N_2254);
nor U4209 (N_4209,N_555,N_1175);
nor U4210 (N_4210,N_604,N_1442);
nor U4211 (N_4211,N_2490,N_2226);
and U4212 (N_4212,N_16,N_1481);
nor U4213 (N_4213,N_1709,N_1218);
or U4214 (N_4214,N_1531,N_1757);
and U4215 (N_4215,N_2496,N_5);
nor U4216 (N_4216,N_241,N_452);
or U4217 (N_4217,N_738,N_2083);
nor U4218 (N_4218,N_902,N_793);
nor U4219 (N_4219,N_2127,N_1871);
nor U4220 (N_4220,N_1932,N_1529);
nor U4221 (N_4221,N_686,N_556);
nand U4222 (N_4222,N_1998,N_385);
nand U4223 (N_4223,N_1539,N_374);
or U4224 (N_4224,N_774,N_1494);
nand U4225 (N_4225,N_2231,N_1482);
and U4226 (N_4226,N_1892,N_1477);
xnor U4227 (N_4227,N_811,N_1774);
nand U4228 (N_4228,N_2059,N_1470);
or U4229 (N_4229,N_756,N_13);
nand U4230 (N_4230,N_677,N_146);
or U4231 (N_4231,N_1383,N_167);
nor U4232 (N_4232,N_2194,N_54);
nand U4233 (N_4233,N_98,N_2303);
nor U4234 (N_4234,N_2212,N_1597);
xnor U4235 (N_4235,N_63,N_928);
and U4236 (N_4236,N_1229,N_826);
or U4237 (N_4237,N_1654,N_1892);
or U4238 (N_4238,N_1285,N_2432);
and U4239 (N_4239,N_1751,N_1781);
or U4240 (N_4240,N_1518,N_40);
nand U4241 (N_4241,N_1007,N_2214);
and U4242 (N_4242,N_1268,N_1183);
nor U4243 (N_4243,N_1814,N_1329);
nand U4244 (N_4244,N_888,N_590);
nand U4245 (N_4245,N_2004,N_2128);
and U4246 (N_4246,N_55,N_2279);
nor U4247 (N_4247,N_1034,N_471);
or U4248 (N_4248,N_303,N_497);
or U4249 (N_4249,N_529,N_2445);
xnor U4250 (N_4250,N_2440,N_11);
nand U4251 (N_4251,N_608,N_199);
nor U4252 (N_4252,N_2242,N_1170);
nand U4253 (N_4253,N_131,N_2082);
or U4254 (N_4254,N_1830,N_1564);
nor U4255 (N_4255,N_333,N_406);
and U4256 (N_4256,N_489,N_1696);
nor U4257 (N_4257,N_1293,N_1931);
nand U4258 (N_4258,N_2485,N_710);
nand U4259 (N_4259,N_973,N_1755);
nand U4260 (N_4260,N_234,N_1011);
nor U4261 (N_4261,N_1799,N_1018);
or U4262 (N_4262,N_1189,N_842);
and U4263 (N_4263,N_2217,N_1121);
and U4264 (N_4264,N_1881,N_2365);
or U4265 (N_4265,N_2112,N_462);
and U4266 (N_4266,N_2218,N_325);
and U4267 (N_4267,N_202,N_1086);
and U4268 (N_4268,N_1592,N_555);
nand U4269 (N_4269,N_625,N_795);
nand U4270 (N_4270,N_494,N_2250);
nand U4271 (N_4271,N_2335,N_1445);
nor U4272 (N_4272,N_2010,N_1733);
or U4273 (N_4273,N_1354,N_282);
or U4274 (N_4274,N_887,N_881);
nand U4275 (N_4275,N_1307,N_2025);
nor U4276 (N_4276,N_1314,N_422);
or U4277 (N_4277,N_428,N_942);
and U4278 (N_4278,N_2246,N_1347);
and U4279 (N_4279,N_350,N_2031);
nand U4280 (N_4280,N_1732,N_563);
and U4281 (N_4281,N_852,N_883);
or U4282 (N_4282,N_798,N_364);
nor U4283 (N_4283,N_1305,N_2146);
nor U4284 (N_4284,N_2192,N_695);
nand U4285 (N_4285,N_1475,N_2221);
nor U4286 (N_4286,N_125,N_1050);
nand U4287 (N_4287,N_2492,N_1139);
nand U4288 (N_4288,N_2007,N_1931);
or U4289 (N_4289,N_733,N_1430);
nand U4290 (N_4290,N_1734,N_165);
and U4291 (N_4291,N_1102,N_2445);
nand U4292 (N_4292,N_224,N_1156);
and U4293 (N_4293,N_1329,N_1403);
xnor U4294 (N_4294,N_697,N_805);
nor U4295 (N_4295,N_1672,N_369);
or U4296 (N_4296,N_376,N_1038);
nor U4297 (N_4297,N_800,N_2430);
nand U4298 (N_4298,N_682,N_756);
nor U4299 (N_4299,N_1813,N_400);
or U4300 (N_4300,N_2405,N_1888);
nor U4301 (N_4301,N_1798,N_696);
xnor U4302 (N_4302,N_700,N_2003);
nor U4303 (N_4303,N_1467,N_768);
nor U4304 (N_4304,N_2154,N_789);
and U4305 (N_4305,N_270,N_924);
and U4306 (N_4306,N_1707,N_154);
nor U4307 (N_4307,N_950,N_1940);
xnor U4308 (N_4308,N_444,N_493);
or U4309 (N_4309,N_1802,N_1630);
nor U4310 (N_4310,N_1788,N_1582);
nand U4311 (N_4311,N_701,N_1748);
and U4312 (N_4312,N_795,N_1953);
nor U4313 (N_4313,N_1936,N_982);
xnor U4314 (N_4314,N_1759,N_1885);
xnor U4315 (N_4315,N_1681,N_1385);
nand U4316 (N_4316,N_203,N_2363);
xnor U4317 (N_4317,N_167,N_874);
nor U4318 (N_4318,N_2207,N_373);
nor U4319 (N_4319,N_601,N_501);
or U4320 (N_4320,N_1489,N_333);
and U4321 (N_4321,N_2067,N_785);
or U4322 (N_4322,N_2151,N_844);
xor U4323 (N_4323,N_1681,N_1048);
or U4324 (N_4324,N_1902,N_648);
xnor U4325 (N_4325,N_1369,N_1687);
nor U4326 (N_4326,N_1446,N_1613);
or U4327 (N_4327,N_1002,N_1437);
and U4328 (N_4328,N_628,N_1698);
and U4329 (N_4329,N_824,N_2461);
nor U4330 (N_4330,N_220,N_1039);
and U4331 (N_4331,N_2474,N_1135);
or U4332 (N_4332,N_1782,N_1417);
nor U4333 (N_4333,N_998,N_506);
and U4334 (N_4334,N_307,N_1619);
nand U4335 (N_4335,N_798,N_2006);
nand U4336 (N_4336,N_468,N_557);
or U4337 (N_4337,N_1176,N_1666);
nor U4338 (N_4338,N_2457,N_145);
and U4339 (N_4339,N_2336,N_602);
or U4340 (N_4340,N_1781,N_1183);
nand U4341 (N_4341,N_2159,N_1499);
nor U4342 (N_4342,N_562,N_465);
xnor U4343 (N_4343,N_2034,N_1369);
or U4344 (N_4344,N_456,N_1012);
nand U4345 (N_4345,N_476,N_2477);
or U4346 (N_4346,N_2041,N_2299);
xnor U4347 (N_4347,N_1175,N_566);
xor U4348 (N_4348,N_1806,N_827);
and U4349 (N_4349,N_2058,N_734);
or U4350 (N_4350,N_325,N_1333);
nor U4351 (N_4351,N_2444,N_903);
and U4352 (N_4352,N_1369,N_2123);
and U4353 (N_4353,N_2347,N_674);
nand U4354 (N_4354,N_753,N_981);
nand U4355 (N_4355,N_1150,N_639);
nand U4356 (N_4356,N_1995,N_2172);
and U4357 (N_4357,N_2119,N_467);
nor U4358 (N_4358,N_440,N_1398);
nor U4359 (N_4359,N_1906,N_930);
nand U4360 (N_4360,N_548,N_296);
nor U4361 (N_4361,N_152,N_1185);
and U4362 (N_4362,N_1958,N_1717);
nor U4363 (N_4363,N_1768,N_1063);
nand U4364 (N_4364,N_1096,N_799);
or U4365 (N_4365,N_1991,N_146);
nand U4366 (N_4366,N_2492,N_298);
and U4367 (N_4367,N_293,N_520);
nor U4368 (N_4368,N_2267,N_373);
and U4369 (N_4369,N_1156,N_2123);
xnor U4370 (N_4370,N_273,N_321);
nand U4371 (N_4371,N_2017,N_374);
or U4372 (N_4372,N_1359,N_1686);
or U4373 (N_4373,N_931,N_2256);
nor U4374 (N_4374,N_2034,N_2143);
and U4375 (N_4375,N_2112,N_2473);
nor U4376 (N_4376,N_1887,N_2475);
nand U4377 (N_4377,N_993,N_1392);
xnor U4378 (N_4378,N_565,N_128);
and U4379 (N_4379,N_1098,N_1532);
and U4380 (N_4380,N_1073,N_534);
and U4381 (N_4381,N_1518,N_1654);
nor U4382 (N_4382,N_872,N_1926);
nor U4383 (N_4383,N_1832,N_1633);
and U4384 (N_4384,N_1684,N_339);
nor U4385 (N_4385,N_2291,N_535);
nand U4386 (N_4386,N_301,N_1575);
nor U4387 (N_4387,N_540,N_1764);
xnor U4388 (N_4388,N_1003,N_1696);
and U4389 (N_4389,N_313,N_565);
nand U4390 (N_4390,N_2146,N_2215);
nor U4391 (N_4391,N_81,N_2294);
or U4392 (N_4392,N_916,N_1477);
xnor U4393 (N_4393,N_323,N_1757);
and U4394 (N_4394,N_2140,N_2249);
nor U4395 (N_4395,N_1536,N_2093);
and U4396 (N_4396,N_699,N_1643);
nand U4397 (N_4397,N_1879,N_1888);
xor U4398 (N_4398,N_1962,N_490);
nor U4399 (N_4399,N_2176,N_1282);
nand U4400 (N_4400,N_1370,N_2432);
nor U4401 (N_4401,N_2054,N_1978);
nor U4402 (N_4402,N_1778,N_1510);
and U4403 (N_4403,N_1389,N_2007);
nand U4404 (N_4404,N_311,N_1863);
and U4405 (N_4405,N_28,N_2338);
and U4406 (N_4406,N_2197,N_1149);
nand U4407 (N_4407,N_94,N_1623);
and U4408 (N_4408,N_1381,N_852);
or U4409 (N_4409,N_2403,N_2346);
nor U4410 (N_4410,N_1675,N_1107);
nand U4411 (N_4411,N_2446,N_2129);
or U4412 (N_4412,N_1037,N_2060);
nor U4413 (N_4413,N_311,N_720);
or U4414 (N_4414,N_193,N_2482);
and U4415 (N_4415,N_1366,N_2478);
or U4416 (N_4416,N_455,N_336);
and U4417 (N_4417,N_141,N_692);
nand U4418 (N_4418,N_2340,N_872);
or U4419 (N_4419,N_1612,N_2277);
and U4420 (N_4420,N_822,N_2318);
and U4421 (N_4421,N_1080,N_97);
nand U4422 (N_4422,N_739,N_2008);
xor U4423 (N_4423,N_1481,N_1161);
or U4424 (N_4424,N_1100,N_1538);
and U4425 (N_4425,N_1440,N_341);
or U4426 (N_4426,N_1049,N_1791);
and U4427 (N_4427,N_1282,N_946);
nand U4428 (N_4428,N_148,N_1075);
nor U4429 (N_4429,N_116,N_1726);
nand U4430 (N_4430,N_2077,N_285);
nor U4431 (N_4431,N_594,N_131);
or U4432 (N_4432,N_2334,N_1966);
xor U4433 (N_4433,N_420,N_1253);
nor U4434 (N_4434,N_128,N_447);
xnor U4435 (N_4435,N_280,N_2154);
or U4436 (N_4436,N_1972,N_855);
and U4437 (N_4437,N_1665,N_2056);
nand U4438 (N_4438,N_343,N_2248);
nand U4439 (N_4439,N_123,N_1194);
or U4440 (N_4440,N_987,N_2045);
or U4441 (N_4441,N_1623,N_474);
xor U4442 (N_4442,N_1075,N_659);
nor U4443 (N_4443,N_1694,N_721);
nor U4444 (N_4444,N_1660,N_1283);
nor U4445 (N_4445,N_973,N_2010);
xnor U4446 (N_4446,N_41,N_364);
or U4447 (N_4447,N_1111,N_1418);
nand U4448 (N_4448,N_1292,N_1584);
nor U4449 (N_4449,N_592,N_1715);
nor U4450 (N_4450,N_2211,N_2450);
nor U4451 (N_4451,N_316,N_970);
or U4452 (N_4452,N_316,N_1322);
xor U4453 (N_4453,N_1974,N_105);
or U4454 (N_4454,N_2293,N_105);
and U4455 (N_4455,N_950,N_2171);
and U4456 (N_4456,N_710,N_1899);
or U4457 (N_4457,N_69,N_1869);
and U4458 (N_4458,N_1747,N_1178);
and U4459 (N_4459,N_990,N_2154);
nor U4460 (N_4460,N_1937,N_677);
or U4461 (N_4461,N_469,N_545);
and U4462 (N_4462,N_293,N_2162);
or U4463 (N_4463,N_1738,N_2334);
and U4464 (N_4464,N_51,N_278);
and U4465 (N_4465,N_435,N_1049);
and U4466 (N_4466,N_334,N_1386);
nand U4467 (N_4467,N_1132,N_1743);
or U4468 (N_4468,N_1254,N_802);
xnor U4469 (N_4469,N_943,N_1525);
xnor U4470 (N_4470,N_2013,N_799);
nand U4471 (N_4471,N_2398,N_133);
and U4472 (N_4472,N_925,N_230);
and U4473 (N_4473,N_1816,N_1677);
nor U4474 (N_4474,N_1829,N_2071);
and U4475 (N_4475,N_53,N_892);
nor U4476 (N_4476,N_1051,N_873);
and U4477 (N_4477,N_1872,N_2364);
nor U4478 (N_4478,N_1280,N_2262);
or U4479 (N_4479,N_1506,N_1430);
or U4480 (N_4480,N_185,N_912);
nor U4481 (N_4481,N_231,N_1715);
nand U4482 (N_4482,N_1436,N_1375);
nor U4483 (N_4483,N_2115,N_2065);
xor U4484 (N_4484,N_2035,N_1265);
nand U4485 (N_4485,N_1278,N_2092);
and U4486 (N_4486,N_2333,N_1692);
nor U4487 (N_4487,N_867,N_2477);
or U4488 (N_4488,N_1590,N_503);
xnor U4489 (N_4489,N_490,N_1736);
nor U4490 (N_4490,N_1705,N_1605);
xor U4491 (N_4491,N_1715,N_1813);
nand U4492 (N_4492,N_2044,N_534);
and U4493 (N_4493,N_2113,N_2204);
and U4494 (N_4494,N_2450,N_774);
or U4495 (N_4495,N_1803,N_2115);
nand U4496 (N_4496,N_823,N_955);
nor U4497 (N_4497,N_2384,N_138);
nor U4498 (N_4498,N_979,N_2368);
nand U4499 (N_4499,N_2451,N_306);
nor U4500 (N_4500,N_984,N_1823);
and U4501 (N_4501,N_2222,N_1880);
nor U4502 (N_4502,N_830,N_1680);
nor U4503 (N_4503,N_1127,N_2046);
nor U4504 (N_4504,N_219,N_2300);
and U4505 (N_4505,N_1356,N_2475);
or U4506 (N_4506,N_1736,N_793);
nand U4507 (N_4507,N_1044,N_556);
xnor U4508 (N_4508,N_1986,N_114);
and U4509 (N_4509,N_947,N_1453);
xor U4510 (N_4510,N_1309,N_1421);
and U4511 (N_4511,N_922,N_764);
nor U4512 (N_4512,N_1674,N_1151);
or U4513 (N_4513,N_82,N_1975);
xor U4514 (N_4514,N_2020,N_423);
and U4515 (N_4515,N_1126,N_659);
nand U4516 (N_4516,N_494,N_2155);
or U4517 (N_4517,N_473,N_476);
nor U4518 (N_4518,N_70,N_1058);
xnor U4519 (N_4519,N_237,N_308);
or U4520 (N_4520,N_2201,N_396);
or U4521 (N_4521,N_351,N_355);
nor U4522 (N_4522,N_1359,N_1369);
nand U4523 (N_4523,N_1717,N_349);
or U4524 (N_4524,N_1042,N_1116);
nand U4525 (N_4525,N_1181,N_1660);
or U4526 (N_4526,N_2012,N_43);
or U4527 (N_4527,N_1967,N_2442);
and U4528 (N_4528,N_1818,N_1668);
nor U4529 (N_4529,N_974,N_1665);
nand U4530 (N_4530,N_2010,N_411);
nand U4531 (N_4531,N_173,N_1285);
and U4532 (N_4532,N_1124,N_1230);
nand U4533 (N_4533,N_795,N_728);
or U4534 (N_4534,N_1188,N_1475);
nor U4535 (N_4535,N_1199,N_496);
nor U4536 (N_4536,N_2399,N_635);
or U4537 (N_4537,N_2427,N_1506);
and U4538 (N_4538,N_1131,N_1686);
nand U4539 (N_4539,N_341,N_93);
nor U4540 (N_4540,N_682,N_2101);
nand U4541 (N_4541,N_208,N_1019);
xor U4542 (N_4542,N_1953,N_1137);
and U4543 (N_4543,N_514,N_1296);
nor U4544 (N_4544,N_954,N_583);
or U4545 (N_4545,N_1991,N_775);
or U4546 (N_4546,N_1360,N_2147);
nor U4547 (N_4547,N_2144,N_266);
nor U4548 (N_4548,N_1792,N_2363);
or U4549 (N_4549,N_1376,N_173);
nor U4550 (N_4550,N_177,N_1008);
nor U4551 (N_4551,N_724,N_872);
nand U4552 (N_4552,N_1820,N_1149);
xnor U4553 (N_4553,N_563,N_1011);
nor U4554 (N_4554,N_1899,N_1383);
and U4555 (N_4555,N_2360,N_498);
nor U4556 (N_4556,N_1172,N_1848);
or U4557 (N_4557,N_2088,N_577);
nor U4558 (N_4558,N_2057,N_846);
nor U4559 (N_4559,N_1044,N_1733);
xnor U4560 (N_4560,N_957,N_1175);
xor U4561 (N_4561,N_243,N_596);
and U4562 (N_4562,N_1854,N_1687);
or U4563 (N_4563,N_182,N_1618);
nand U4564 (N_4564,N_272,N_832);
nor U4565 (N_4565,N_584,N_1875);
nor U4566 (N_4566,N_892,N_1356);
nand U4567 (N_4567,N_1737,N_2100);
and U4568 (N_4568,N_1950,N_2233);
or U4569 (N_4569,N_1743,N_2214);
nor U4570 (N_4570,N_1024,N_1190);
and U4571 (N_4571,N_988,N_2211);
xor U4572 (N_4572,N_2135,N_364);
nor U4573 (N_4573,N_1180,N_1647);
nor U4574 (N_4574,N_1543,N_2407);
or U4575 (N_4575,N_1044,N_340);
or U4576 (N_4576,N_1220,N_403);
or U4577 (N_4577,N_845,N_1693);
and U4578 (N_4578,N_1587,N_1578);
nor U4579 (N_4579,N_2404,N_1426);
and U4580 (N_4580,N_278,N_2177);
nand U4581 (N_4581,N_1978,N_2083);
and U4582 (N_4582,N_103,N_210);
nand U4583 (N_4583,N_559,N_1234);
and U4584 (N_4584,N_135,N_1793);
or U4585 (N_4585,N_870,N_1199);
or U4586 (N_4586,N_78,N_694);
nor U4587 (N_4587,N_330,N_196);
nand U4588 (N_4588,N_1696,N_642);
xnor U4589 (N_4589,N_309,N_260);
nor U4590 (N_4590,N_345,N_1927);
and U4591 (N_4591,N_2070,N_1366);
nor U4592 (N_4592,N_1767,N_1152);
and U4593 (N_4593,N_1977,N_1122);
nor U4594 (N_4594,N_2223,N_181);
nor U4595 (N_4595,N_1735,N_2310);
and U4596 (N_4596,N_1333,N_139);
and U4597 (N_4597,N_775,N_778);
and U4598 (N_4598,N_2132,N_2110);
nor U4599 (N_4599,N_609,N_1080);
or U4600 (N_4600,N_1362,N_219);
and U4601 (N_4601,N_719,N_2026);
and U4602 (N_4602,N_1094,N_1366);
nor U4603 (N_4603,N_607,N_2291);
and U4604 (N_4604,N_2303,N_1537);
nand U4605 (N_4605,N_1019,N_963);
nand U4606 (N_4606,N_2300,N_466);
nor U4607 (N_4607,N_1527,N_116);
nand U4608 (N_4608,N_172,N_1538);
or U4609 (N_4609,N_288,N_80);
nand U4610 (N_4610,N_1344,N_1476);
nor U4611 (N_4611,N_2222,N_408);
and U4612 (N_4612,N_1259,N_2294);
nand U4613 (N_4613,N_1975,N_1638);
and U4614 (N_4614,N_1472,N_559);
nand U4615 (N_4615,N_749,N_1511);
xnor U4616 (N_4616,N_1456,N_1307);
nand U4617 (N_4617,N_480,N_2300);
and U4618 (N_4618,N_24,N_425);
nand U4619 (N_4619,N_2047,N_2469);
nand U4620 (N_4620,N_1131,N_679);
or U4621 (N_4621,N_2012,N_616);
and U4622 (N_4622,N_1574,N_2139);
and U4623 (N_4623,N_1122,N_1665);
or U4624 (N_4624,N_522,N_1960);
and U4625 (N_4625,N_1700,N_666);
nor U4626 (N_4626,N_757,N_955);
nand U4627 (N_4627,N_743,N_278);
nor U4628 (N_4628,N_1530,N_483);
and U4629 (N_4629,N_1502,N_1027);
nand U4630 (N_4630,N_873,N_2053);
nor U4631 (N_4631,N_2467,N_2044);
and U4632 (N_4632,N_1602,N_1106);
nor U4633 (N_4633,N_87,N_2329);
nor U4634 (N_4634,N_1519,N_2289);
nor U4635 (N_4635,N_2336,N_2178);
or U4636 (N_4636,N_729,N_250);
and U4637 (N_4637,N_1549,N_1393);
and U4638 (N_4638,N_1905,N_1806);
nand U4639 (N_4639,N_2207,N_935);
or U4640 (N_4640,N_1288,N_780);
or U4641 (N_4641,N_114,N_2345);
nand U4642 (N_4642,N_1080,N_1944);
or U4643 (N_4643,N_2456,N_57);
or U4644 (N_4644,N_1867,N_1458);
nor U4645 (N_4645,N_325,N_933);
nor U4646 (N_4646,N_989,N_1608);
nor U4647 (N_4647,N_1025,N_260);
xor U4648 (N_4648,N_906,N_2239);
or U4649 (N_4649,N_1313,N_2487);
or U4650 (N_4650,N_1996,N_2113);
nand U4651 (N_4651,N_2381,N_289);
and U4652 (N_4652,N_2176,N_592);
and U4653 (N_4653,N_1938,N_806);
nand U4654 (N_4654,N_2036,N_1974);
and U4655 (N_4655,N_279,N_2081);
and U4656 (N_4656,N_1305,N_2389);
and U4657 (N_4657,N_1989,N_336);
nand U4658 (N_4658,N_1095,N_842);
and U4659 (N_4659,N_397,N_463);
nand U4660 (N_4660,N_1580,N_2118);
and U4661 (N_4661,N_2160,N_1705);
nand U4662 (N_4662,N_2103,N_519);
nor U4663 (N_4663,N_1322,N_1655);
nand U4664 (N_4664,N_341,N_360);
and U4665 (N_4665,N_1918,N_152);
nor U4666 (N_4666,N_831,N_1360);
or U4667 (N_4667,N_563,N_272);
nor U4668 (N_4668,N_1065,N_1684);
or U4669 (N_4669,N_345,N_1358);
or U4670 (N_4670,N_403,N_1689);
xor U4671 (N_4671,N_231,N_510);
and U4672 (N_4672,N_2473,N_1942);
and U4673 (N_4673,N_1968,N_13);
nor U4674 (N_4674,N_790,N_518);
and U4675 (N_4675,N_1897,N_2215);
nor U4676 (N_4676,N_1780,N_1748);
or U4677 (N_4677,N_2153,N_1879);
and U4678 (N_4678,N_1573,N_867);
nor U4679 (N_4679,N_275,N_752);
nor U4680 (N_4680,N_216,N_1120);
and U4681 (N_4681,N_456,N_171);
nor U4682 (N_4682,N_651,N_1984);
nor U4683 (N_4683,N_2005,N_2470);
nor U4684 (N_4684,N_1208,N_285);
and U4685 (N_4685,N_446,N_1964);
nand U4686 (N_4686,N_1619,N_1280);
or U4687 (N_4687,N_2259,N_1265);
nand U4688 (N_4688,N_1732,N_1953);
and U4689 (N_4689,N_356,N_237);
nand U4690 (N_4690,N_1646,N_101);
nand U4691 (N_4691,N_1733,N_512);
and U4692 (N_4692,N_849,N_1685);
or U4693 (N_4693,N_1454,N_674);
nor U4694 (N_4694,N_535,N_2398);
nand U4695 (N_4695,N_963,N_1983);
nor U4696 (N_4696,N_385,N_2137);
nand U4697 (N_4697,N_403,N_1024);
or U4698 (N_4698,N_980,N_1711);
or U4699 (N_4699,N_1553,N_1514);
nand U4700 (N_4700,N_1958,N_1242);
and U4701 (N_4701,N_1315,N_535);
and U4702 (N_4702,N_885,N_272);
or U4703 (N_4703,N_845,N_2192);
nor U4704 (N_4704,N_1306,N_757);
xor U4705 (N_4705,N_1947,N_112);
or U4706 (N_4706,N_1606,N_688);
or U4707 (N_4707,N_2421,N_2088);
nand U4708 (N_4708,N_276,N_1004);
and U4709 (N_4709,N_2261,N_256);
nand U4710 (N_4710,N_1127,N_1327);
nand U4711 (N_4711,N_474,N_2430);
nor U4712 (N_4712,N_879,N_1171);
nand U4713 (N_4713,N_221,N_1754);
and U4714 (N_4714,N_2149,N_1465);
and U4715 (N_4715,N_749,N_2033);
and U4716 (N_4716,N_2343,N_1462);
and U4717 (N_4717,N_1023,N_1111);
xnor U4718 (N_4718,N_1366,N_2333);
nor U4719 (N_4719,N_307,N_92);
nor U4720 (N_4720,N_583,N_75);
and U4721 (N_4721,N_330,N_1930);
nor U4722 (N_4722,N_2041,N_1063);
nor U4723 (N_4723,N_2149,N_1073);
or U4724 (N_4724,N_1986,N_1558);
and U4725 (N_4725,N_2447,N_1558);
nor U4726 (N_4726,N_1544,N_1161);
nand U4727 (N_4727,N_378,N_2181);
nand U4728 (N_4728,N_981,N_2271);
and U4729 (N_4729,N_514,N_1355);
nor U4730 (N_4730,N_1017,N_1502);
or U4731 (N_4731,N_1781,N_1665);
xor U4732 (N_4732,N_1425,N_1226);
nand U4733 (N_4733,N_1732,N_619);
nand U4734 (N_4734,N_634,N_1523);
and U4735 (N_4735,N_1152,N_1947);
nor U4736 (N_4736,N_993,N_95);
and U4737 (N_4737,N_2024,N_403);
xor U4738 (N_4738,N_1767,N_1493);
nor U4739 (N_4739,N_1941,N_431);
or U4740 (N_4740,N_406,N_727);
nand U4741 (N_4741,N_115,N_2110);
and U4742 (N_4742,N_1303,N_1052);
nor U4743 (N_4743,N_1360,N_637);
nand U4744 (N_4744,N_1879,N_890);
nand U4745 (N_4745,N_1019,N_1305);
xor U4746 (N_4746,N_2178,N_1707);
or U4747 (N_4747,N_2206,N_1000);
or U4748 (N_4748,N_1368,N_2264);
nand U4749 (N_4749,N_2417,N_2172);
xor U4750 (N_4750,N_1358,N_2334);
or U4751 (N_4751,N_862,N_1810);
nor U4752 (N_4752,N_1455,N_590);
nor U4753 (N_4753,N_537,N_2292);
and U4754 (N_4754,N_1319,N_2158);
or U4755 (N_4755,N_544,N_1759);
nor U4756 (N_4756,N_574,N_245);
xor U4757 (N_4757,N_1904,N_866);
nand U4758 (N_4758,N_2434,N_2052);
nor U4759 (N_4759,N_1743,N_2168);
xnor U4760 (N_4760,N_2143,N_2308);
nor U4761 (N_4761,N_2057,N_2287);
nand U4762 (N_4762,N_296,N_379);
and U4763 (N_4763,N_742,N_2494);
nand U4764 (N_4764,N_1355,N_2405);
nand U4765 (N_4765,N_1150,N_433);
xor U4766 (N_4766,N_1236,N_1225);
and U4767 (N_4767,N_2492,N_2136);
or U4768 (N_4768,N_874,N_787);
and U4769 (N_4769,N_402,N_1901);
nand U4770 (N_4770,N_1705,N_332);
nand U4771 (N_4771,N_390,N_2414);
or U4772 (N_4772,N_1238,N_537);
nand U4773 (N_4773,N_1879,N_555);
nand U4774 (N_4774,N_572,N_292);
and U4775 (N_4775,N_747,N_274);
nand U4776 (N_4776,N_1315,N_2488);
nor U4777 (N_4777,N_2127,N_1013);
and U4778 (N_4778,N_960,N_1904);
and U4779 (N_4779,N_1497,N_8);
nand U4780 (N_4780,N_157,N_619);
and U4781 (N_4781,N_2243,N_2112);
nand U4782 (N_4782,N_1306,N_2266);
xnor U4783 (N_4783,N_1012,N_1681);
and U4784 (N_4784,N_1198,N_1693);
and U4785 (N_4785,N_2486,N_1658);
and U4786 (N_4786,N_470,N_46);
nor U4787 (N_4787,N_1538,N_2143);
and U4788 (N_4788,N_2182,N_1013);
or U4789 (N_4789,N_221,N_254);
and U4790 (N_4790,N_1867,N_2304);
and U4791 (N_4791,N_353,N_1695);
or U4792 (N_4792,N_1239,N_396);
nor U4793 (N_4793,N_1774,N_1787);
and U4794 (N_4794,N_1033,N_1755);
or U4795 (N_4795,N_1781,N_96);
nand U4796 (N_4796,N_2480,N_1397);
or U4797 (N_4797,N_1593,N_130);
nand U4798 (N_4798,N_829,N_173);
nand U4799 (N_4799,N_1499,N_1498);
and U4800 (N_4800,N_1024,N_94);
nand U4801 (N_4801,N_152,N_28);
and U4802 (N_4802,N_1257,N_1775);
or U4803 (N_4803,N_1555,N_2128);
and U4804 (N_4804,N_1944,N_2323);
nor U4805 (N_4805,N_203,N_296);
nor U4806 (N_4806,N_1799,N_2443);
or U4807 (N_4807,N_1974,N_1121);
nand U4808 (N_4808,N_373,N_289);
nand U4809 (N_4809,N_686,N_2486);
and U4810 (N_4810,N_1246,N_1842);
and U4811 (N_4811,N_394,N_2292);
or U4812 (N_4812,N_126,N_430);
and U4813 (N_4813,N_1719,N_2246);
and U4814 (N_4814,N_144,N_871);
nor U4815 (N_4815,N_930,N_1000);
nand U4816 (N_4816,N_1203,N_852);
nor U4817 (N_4817,N_1020,N_1872);
nand U4818 (N_4818,N_214,N_1948);
nor U4819 (N_4819,N_1991,N_557);
or U4820 (N_4820,N_1384,N_1124);
nand U4821 (N_4821,N_2156,N_411);
nor U4822 (N_4822,N_2044,N_1738);
or U4823 (N_4823,N_855,N_1633);
nor U4824 (N_4824,N_1113,N_790);
or U4825 (N_4825,N_1409,N_170);
or U4826 (N_4826,N_1804,N_1275);
xor U4827 (N_4827,N_323,N_2441);
or U4828 (N_4828,N_132,N_525);
xor U4829 (N_4829,N_158,N_352);
nor U4830 (N_4830,N_1060,N_2433);
nor U4831 (N_4831,N_527,N_2189);
and U4832 (N_4832,N_1106,N_536);
nor U4833 (N_4833,N_261,N_398);
nor U4834 (N_4834,N_1950,N_566);
nor U4835 (N_4835,N_273,N_1746);
and U4836 (N_4836,N_800,N_2079);
and U4837 (N_4837,N_1200,N_1318);
nand U4838 (N_4838,N_2432,N_1420);
xor U4839 (N_4839,N_1602,N_490);
nand U4840 (N_4840,N_1288,N_123);
or U4841 (N_4841,N_256,N_2314);
xnor U4842 (N_4842,N_658,N_496);
nand U4843 (N_4843,N_2054,N_1279);
nor U4844 (N_4844,N_1131,N_2401);
nand U4845 (N_4845,N_57,N_1478);
nor U4846 (N_4846,N_1916,N_638);
nand U4847 (N_4847,N_1973,N_1381);
nand U4848 (N_4848,N_449,N_2192);
nand U4849 (N_4849,N_1574,N_845);
xor U4850 (N_4850,N_360,N_460);
and U4851 (N_4851,N_1063,N_1602);
nand U4852 (N_4852,N_388,N_464);
and U4853 (N_4853,N_1125,N_2366);
nor U4854 (N_4854,N_1340,N_1831);
and U4855 (N_4855,N_1871,N_2061);
nand U4856 (N_4856,N_44,N_56);
nor U4857 (N_4857,N_748,N_2427);
and U4858 (N_4858,N_750,N_1177);
and U4859 (N_4859,N_1580,N_629);
nor U4860 (N_4860,N_2164,N_1368);
nor U4861 (N_4861,N_1790,N_1732);
or U4862 (N_4862,N_715,N_1495);
nor U4863 (N_4863,N_2133,N_420);
xnor U4864 (N_4864,N_722,N_1549);
and U4865 (N_4865,N_1445,N_2435);
and U4866 (N_4866,N_219,N_1576);
and U4867 (N_4867,N_1728,N_2058);
nor U4868 (N_4868,N_123,N_1219);
and U4869 (N_4869,N_2087,N_1382);
or U4870 (N_4870,N_344,N_1383);
nand U4871 (N_4871,N_2229,N_850);
nor U4872 (N_4872,N_1394,N_41);
nand U4873 (N_4873,N_300,N_2449);
or U4874 (N_4874,N_1415,N_688);
nor U4875 (N_4875,N_422,N_1430);
or U4876 (N_4876,N_402,N_2348);
nor U4877 (N_4877,N_1265,N_1648);
nor U4878 (N_4878,N_1573,N_2198);
or U4879 (N_4879,N_1105,N_819);
nand U4880 (N_4880,N_1368,N_1444);
xor U4881 (N_4881,N_1878,N_2390);
or U4882 (N_4882,N_1355,N_2057);
xor U4883 (N_4883,N_1692,N_2452);
and U4884 (N_4884,N_899,N_20);
nor U4885 (N_4885,N_145,N_2139);
xor U4886 (N_4886,N_1447,N_491);
nor U4887 (N_4887,N_2436,N_2032);
nor U4888 (N_4888,N_670,N_861);
nand U4889 (N_4889,N_2052,N_33);
nor U4890 (N_4890,N_1831,N_1723);
nand U4891 (N_4891,N_2358,N_1785);
or U4892 (N_4892,N_1237,N_509);
and U4893 (N_4893,N_995,N_1315);
and U4894 (N_4894,N_197,N_1808);
nor U4895 (N_4895,N_395,N_119);
nor U4896 (N_4896,N_622,N_1342);
and U4897 (N_4897,N_2417,N_629);
nor U4898 (N_4898,N_891,N_2278);
nor U4899 (N_4899,N_100,N_1825);
nand U4900 (N_4900,N_497,N_2433);
or U4901 (N_4901,N_1769,N_2440);
or U4902 (N_4902,N_1796,N_293);
and U4903 (N_4903,N_292,N_1110);
and U4904 (N_4904,N_1570,N_283);
and U4905 (N_4905,N_410,N_1902);
or U4906 (N_4906,N_421,N_1957);
and U4907 (N_4907,N_2190,N_1256);
nand U4908 (N_4908,N_669,N_1969);
nand U4909 (N_4909,N_2489,N_1383);
and U4910 (N_4910,N_555,N_1414);
and U4911 (N_4911,N_2064,N_2229);
and U4912 (N_4912,N_449,N_1453);
or U4913 (N_4913,N_1268,N_1923);
nand U4914 (N_4914,N_2429,N_267);
and U4915 (N_4915,N_2132,N_1277);
or U4916 (N_4916,N_479,N_469);
and U4917 (N_4917,N_500,N_351);
and U4918 (N_4918,N_1170,N_370);
or U4919 (N_4919,N_2198,N_1990);
and U4920 (N_4920,N_1088,N_1035);
nand U4921 (N_4921,N_306,N_1554);
nand U4922 (N_4922,N_1992,N_557);
and U4923 (N_4923,N_752,N_2002);
or U4924 (N_4924,N_1754,N_1739);
nand U4925 (N_4925,N_1700,N_1204);
and U4926 (N_4926,N_237,N_966);
or U4927 (N_4927,N_2101,N_720);
nand U4928 (N_4928,N_615,N_1997);
and U4929 (N_4929,N_1322,N_1133);
and U4930 (N_4930,N_2321,N_1250);
xor U4931 (N_4931,N_1134,N_770);
nand U4932 (N_4932,N_866,N_1381);
and U4933 (N_4933,N_1660,N_250);
and U4934 (N_4934,N_1116,N_372);
nor U4935 (N_4935,N_2207,N_172);
nor U4936 (N_4936,N_2182,N_723);
and U4937 (N_4937,N_453,N_805);
or U4938 (N_4938,N_1721,N_2163);
nand U4939 (N_4939,N_597,N_749);
and U4940 (N_4940,N_1632,N_1114);
and U4941 (N_4941,N_1782,N_1497);
or U4942 (N_4942,N_312,N_513);
nand U4943 (N_4943,N_228,N_1335);
or U4944 (N_4944,N_2493,N_2237);
and U4945 (N_4945,N_1050,N_1130);
nand U4946 (N_4946,N_1984,N_1427);
nor U4947 (N_4947,N_2485,N_209);
and U4948 (N_4948,N_1040,N_1287);
or U4949 (N_4949,N_465,N_2060);
nand U4950 (N_4950,N_1407,N_1488);
xor U4951 (N_4951,N_353,N_1144);
xor U4952 (N_4952,N_2260,N_929);
or U4953 (N_4953,N_2242,N_1831);
and U4954 (N_4954,N_2132,N_5);
and U4955 (N_4955,N_425,N_1323);
and U4956 (N_4956,N_2479,N_1338);
or U4957 (N_4957,N_1458,N_367);
xnor U4958 (N_4958,N_337,N_2345);
nand U4959 (N_4959,N_2267,N_1584);
nand U4960 (N_4960,N_910,N_1785);
xnor U4961 (N_4961,N_129,N_1133);
nor U4962 (N_4962,N_288,N_218);
nand U4963 (N_4963,N_1024,N_365);
or U4964 (N_4964,N_2240,N_492);
nand U4965 (N_4965,N_365,N_114);
nand U4966 (N_4966,N_1954,N_2173);
nand U4967 (N_4967,N_1467,N_878);
or U4968 (N_4968,N_1712,N_2207);
nand U4969 (N_4969,N_271,N_2295);
nand U4970 (N_4970,N_1434,N_1379);
nor U4971 (N_4971,N_1163,N_272);
nand U4972 (N_4972,N_886,N_534);
or U4973 (N_4973,N_1455,N_1480);
and U4974 (N_4974,N_1113,N_1287);
nor U4975 (N_4975,N_2144,N_1574);
or U4976 (N_4976,N_253,N_883);
and U4977 (N_4977,N_204,N_1496);
nor U4978 (N_4978,N_1272,N_486);
nand U4979 (N_4979,N_0,N_1405);
and U4980 (N_4980,N_2351,N_1165);
xnor U4981 (N_4981,N_697,N_1940);
nand U4982 (N_4982,N_2384,N_2086);
or U4983 (N_4983,N_267,N_2119);
xor U4984 (N_4984,N_2061,N_923);
nand U4985 (N_4985,N_1270,N_338);
xnor U4986 (N_4986,N_1901,N_1335);
or U4987 (N_4987,N_319,N_1165);
nor U4988 (N_4988,N_619,N_2240);
and U4989 (N_4989,N_237,N_1414);
and U4990 (N_4990,N_1208,N_757);
nor U4991 (N_4991,N_826,N_2133);
and U4992 (N_4992,N_102,N_921);
or U4993 (N_4993,N_32,N_528);
nand U4994 (N_4994,N_977,N_2196);
and U4995 (N_4995,N_2035,N_1010);
nor U4996 (N_4996,N_1755,N_2424);
xor U4997 (N_4997,N_1461,N_2477);
or U4998 (N_4998,N_716,N_1542);
or U4999 (N_4999,N_322,N_2332);
and UO_0 (O_0,N_2947,N_4523);
or UO_1 (O_1,N_3440,N_2597);
nor UO_2 (O_2,N_3399,N_3286);
nand UO_3 (O_3,N_4239,N_3976);
nand UO_4 (O_4,N_3364,N_3485);
or UO_5 (O_5,N_3401,N_4910);
and UO_6 (O_6,N_4791,N_2506);
nor UO_7 (O_7,N_4431,N_2626);
or UO_8 (O_8,N_2808,N_4770);
and UO_9 (O_9,N_3175,N_4766);
or UO_10 (O_10,N_2635,N_3841);
nand UO_11 (O_11,N_4584,N_3847);
or UO_12 (O_12,N_4850,N_4599);
nor UO_13 (O_13,N_4180,N_3747);
and UO_14 (O_14,N_4939,N_2696);
nor UO_15 (O_15,N_3562,N_3040);
xor UO_16 (O_16,N_3231,N_3373);
nand UO_17 (O_17,N_3000,N_4484);
or UO_18 (O_18,N_3452,N_4423);
nand UO_19 (O_19,N_3187,N_4588);
or UO_20 (O_20,N_2685,N_3234);
nand UO_21 (O_21,N_3548,N_3676);
nor UO_22 (O_22,N_3059,N_3796);
xor UO_23 (O_23,N_4646,N_3775);
nand UO_24 (O_24,N_3597,N_3051);
and UO_25 (O_25,N_3592,N_3119);
nor UO_26 (O_26,N_3294,N_3803);
nor UO_27 (O_27,N_4847,N_3773);
nand UO_28 (O_28,N_4624,N_4051);
and UO_29 (O_29,N_4244,N_3316);
nor UO_30 (O_30,N_4611,N_4610);
and UO_31 (O_31,N_3354,N_3682);
nand UO_32 (O_32,N_3470,N_4540);
or UO_33 (O_33,N_3355,N_3383);
and UO_34 (O_34,N_4530,N_4962);
and UO_35 (O_35,N_2828,N_3198);
or UO_36 (O_36,N_4020,N_2902);
nand UO_37 (O_37,N_3244,N_3828);
nand UO_38 (O_38,N_4196,N_4178);
and UO_39 (O_39,N_4859,N_4603);
and UO_40 (O_40,N_2981,N_2933);
and UO_41 (O_41,N_4339,N_2997);
or UO_42 (O_42,N_3295,N_2982);
and UO_43 (O_43,N_3025,N_4459);
and UO_44 (O_44,N_3638,N_2629);
nor UO_45 (O_45,N_3115,N_3929);
nor UO_46 (O_46,N_3117,N_4331);
or UO_47 (O_47,N_3118,N_3239);
nor UO_48 (O_48,N_2721,N_3782);
nand UO_49 (O_49,N_4376,N_2925);
nor UO_50 (O_50,N_4042,N_3691);
nand UO_51 (O_51,N_3268,N_3785);
nand UO_52 (O_52,N_4849,N_2729);
and UO_53 (O_53,N_3150,N_4574);
nand UO_54 (O_54,N_3265,N_4297);
or UO_55 (O_55,N_4425,N_3685);
nand UO_56 (O_56,N_3739,N_4455);
nand UO_57 (O_57,N_4966,N_3821);
nand UO_58 (O_58,N_4077,N_2523);
or UO_59 (O_59,N_4729,N_3648);
nand UO_60 (O_60,N_2539,N_3177);
or UO_61 (O_61,N_3420,N_4450);
nand UO_62 (O_62,N_4685,N_2672);
and UO_63 (O_63,N_4979,N_4295);
nand UO_64 (O_64,N_4991,N_4404);
or UO_65 (O_65,N_3126,N_3524);
and UO_66 (O_66,N_2516,N_2863);
nand UO_67 (O_67,N_4678,N_3570);
xor UO_68 (O_68,N_4653,N_4461);
and UO_69 (O_69,N_4413,N_2515);
or UO_70 (O_70,N_2664,N_3971);
or UO_71 (O_71,N_2877,N_3990);
nor UO_72 (O_72,N_2594,N_3802);
or UO_73 (O_73,N_3078,N_2600);
and UO_74 (O_74,N_4107,N_4561);
nor UO_75 (O_75,N_4590,N_4345);
and UO_76 (O_76,N_3887,N_4694);
and UO_77 (O_77,N_3180,N_3409);
nor UO_78 (O_78,N_3549,N_3003);
nand UO_79 (O_79,N_3630,N_3893);
and UO_80 (O_80,N_2561,N_3478);
xnor UO_81 (O_81,N_3708,N_3359);
and UO_82 (O_82,N_4395,N_4935);
nand UO_83 (O_83,N_4741,N_3004);
and UO_84 (O_84,N_3272,N_3700);
nor UO_85 (O_85,N_4274,N_3266);
and UO_86 (O_86,N_3973,N_3002);
nor UO_87 (O_87,N_4056,N_3680);
nor UO_88 (O_88,N_4570,N_4469);
nor UO_89 (O_89,N_4756,N_3728);
nand UO_90 (O_90,N_3001,N_2827);
and UO_91 (O_91,N_4473,N_3015);
nor UO_92 (O_92,N_3972,N_3979);
nand UO_93 (O_93,N_2811,N_2768);
and UO_94 (O_94,N_3139,N_4704);
xor UO_95 (O_95,N_2904,N_3308);
xnor UO_96 (O_96,N_4688,N_4466);
nand UO_97 (O_97,N_4116,N_3085);
or UO_98 (O_98,N_3593,N_4999);
nand UO_99 (O_99,N_4591,N_3859);
or UO_100 (O_100,N_3269,N_3717);
nor UO_101 (O_101,N_4533,N_3169);
nor UO_102 (O_102,N_4169,N_3507);
nand UO_103 (O_103,N_4737,N_3695);
and UO_104 (O_104,N_3835,N_2610);
xor UO_105 (O_105,N_3038,N_4818);
nand UO_106 (O_106,N_4998,N_2607);
xnor UO_107 (O_107,N_3616,N_2874);
or UO_108 (O_108,N_4228,N_2957);
nor UO_109 (O_109,N_3931,N_3170);
xor UO_110 (O_110,N_4234,N_4201);
or UO_111 (O_111,N_4153,N_4213);
nor UO_112 (O_112,N_4257,N_3543);
or UO_113 (O_113,N_3678,N_4028);
or UO_114 (O_114,N_3419,N_3299);
nor UO_115 (O_115,N_3503,N_2631);
nand UO_116 (O_116,N_3960,N_2673);
nor UO_117 (O_117,N_3263,N_3766);
or UO_118 (O_118,N_2545,N_3787);
and UO_119 (O_119,N_2972,N_3309);
or UO_120 (O_120,N_3982,N_4699);
nand UO_121 (O_121,N_3076,N_3948);
nor UO_122 (O_122,N_3249,N_3243);
nand UO_123 (O_123,N_4906,N_3911);
or UO_124 (O_124,N_2782,N_3356);
nor UO_125 (O_125,N_3584,N_4863);
nand UO_126 (O_126,N_3844,N_4072);
xor UO_127 (O_127,N_3995,N_2973);
nand UO_128 (O_128,N_4672,N_3050);
nand UO_129 (O_129,N_4601,N_3544);
and UO_130 (O_130,N_4825,N_4335);
nand UO_131 (O_131,N_4856,N_2718);
and UO_132 (O_132,N_3944,N_4417);
xor UO_133 (O_133,N_2855,N_3932);
and UO_134 (O_134,N_3620,N_2544);
or UO_135 (O_135,N_2533,N_4074);
nor UO_136 (O_136,N_4255,N_4023);
nor UO_137 (O_137,N_2839,N_3462);
nand UO_138 (O_138,N_4617,N_4005);
or UO_139 (O_139,N_2659,N_3573);
nor UO_140 (O_140,N_3293,N_2963);
xnor UO_141 (O_141,N_3558,N_3063);
or UO_142 (O_142,N_2567,N_3255);
nor UO_143 (O_143,N_3846,N_4101);
nand UO_144 (O_144,N_4782,N_4958);
nor UO_145 (O_145,N_2730,N_3923);
and UO_146 (O_146,N_3569,N_3675);
nand UO_147 (O_147,N_4876,N_2714);
or UO_148 (O_148,N_3242,N_3661);
nor UO_149 (O_149,N_4292,N_2707);
or UO_150 (O_150,N_3610,N_3435);
and UO_151 (O_151,N_4615,N_3830);
or UO_152 (O_152,N_4754,N_2527);
xnor UO_153 (O_153,N_4304,N_3635);
nor UO_154 (O_154,N_2873,N_4551);
nand UO_155 (O_155,N_4720,N_3826);
nand UO_156 (O_156,N_3007,N_3288);
and UO_157 (O_157,N_2754,N_2623);
and UO_158 (O_158,N_3371,N_4515);
nor UO_159 (O_159,N_3508,N_2841);
or UO_160 (O_160,N_4318,N_2896);
nor UO_161 (O_161,N_4341,N_3056);
or UO_162 (O_162,N_3860,N_4671);
and UO_163 (O_163,N_4240,N_4711);
nand UO_164 (O_164,N_4186,N_3071);
nand UO_165 (O_165,N_2781,N_4346);
nor UO_166 (O_166,N_3331,N_3969);
nand UO_167 (O_167,N_4717,N_4029);
and UO_168 (O_168,N_4002,N_4984);
nor UO_169 (O_169,N_3457,N_2643);
nand UO_170 (O_170,N_4916,N_2736);
or UO_171 (O_171,N_3403,N_4682);
or UO_172 (O_172,N_2554,N_4157);
or UO_173 (O_173,N_3133,N_3416);
nand UO_174 (O_174,N_4128,N_3504);
nand UO_175 (O_175,N_4495,N_3235);
and UO_176 (O_176,N_2573,N_4506);
xor UO_177 (O_177,N_3824,N_3587);
xnor UO_178 (O_178,N_3800,N_3250);
nand UO_179 (O_179,N_2865,N_4989);
or UO_180 (O_180,N_3657,N_3928);
or UO_181 (O_181,N_2847,N_2753);
or UO_182 (O_182,N_3358,N_2761);
and UO_183 (O_183,N_4263,N_4171);
xor UO_184 (O_184,N_4369,N_4275);
nor UO_185 (O_185,N_4325,N_3653);
and UO_186 (O_186,N_2602,N_4882);
nand UO_187 (O_187,N_3023,N_4626);
nor UO_188 (O_188,N_3527,N_4415);
nand UO_189 (O_189,N_3382,N_4456);
nand UO_190 (O_190,N_2612,N_3389);
xnor UO_191 (O_191,N_2823,N_4793);
nand UO_192 (O_192,N_2652,N_3694);
nand UO_193 (O_193,N_4027,N_2927);
or UO_194 (O_194,N_4161,N_3121);
and UO_195 (O_195,N_3127,N_2857);
or UO_196 (O_196,N_2870,N_4868);
nor UO_197 (O_197,N_4154,N_3545);
nor UO_198 (O_198,N_3429,N_4819);
and UO_199 (O_199,N_3336,N_3431);
or UO_200 (O_200,N_2799,N_4892);
nor UO_201 (O_201,N_4422,N_3892);
nand UO_202 (O_202,N_3745,N_4805);
or UO_203 (O_203,N_4826,N_4973);
nor UO_204 (O_204,N_4017,N_4982);
nand UO_205 (O_205,N_3353,N_4098);
nor UO_206 (O_206,N_3159,N_3940);
nor UO_207 (O_207,N_4602,N_4903);
or UO_208 (O_208,N_4249,N_2627);
nand UO_209 (O_209,N_4477,N_2722);
or UO_210 (O_210,N_2587,N_3408);
or UO_211 (O_211,N_4443,N_4189);
xnor UO_212 (O_212,N_4481,N_3714);
and UO_213 (O_213,N_4195,N_4931);
nand UO_214 (O_214,N_2919,N_4000);
or UO_215 (O_215,N_4299,N_2646);
nor UO_216 (O_216,N_2813,N_4814);
nor UO_217 (O_217,N_3274,N_4514);
nand UO_218 (O_218,N_4250,N_4949);
and UO_219 (O_219,N_2867,N_4645);
and UO_220 (O_220,N_3109,N_4894);
and UO_221 (O_221,N_2632,N_4086);
nand UO_222 (O_222,N_3258,N_4357);
or UO_223 (O_223,N_4727,N_3757);
nand UO_224 (O_224,N_3848,N_4662);
and UO_225 (O_225,N_3722,N_3191);
nor UO_226 (O_226,N_3377,N_4505);
nor UO_227 (O_227,N_4684,N_4963);
and UO_228 (O_228,N_3565,N_4802);
and UO_229 (O_229,N_4489,N_3161);
nor UO_230 (O_230,N_2598,N_2864);
and UO_231 (O_231,N_3376,N_4066);
or UO_232 (O_232,N_3646,N_3060);
nand UO_233 (O_233,N_4651,N_3622);
or UO_234 (O_234,N_3564,N_2738);
nand UO_235 (O_235,N_3780,N_3172);
nand UO_236 (O_236,N_2592,N_4761);
and UO_237 (O_237,N_4546,N_4332);
and UO_238 (O_238,N_4091,N_4730);
nand UO_239 (O_239,N_3985,N_3380);
nor UO_240 (O_240,N_3451,N_3264);
or UO_241 (O_241,N_2688,N_2540);
nand UO_242 (O_242,N_2535,N_3477);
nand UO_243 (O_243,N_2778,N_4719);
nand UO_244 (O_244,N_4801,N_2577);
nor UO_245 (O_245,N_3128,N_2500);
nor UO_246 (O_246,N_3260,N_3934);
and UO_247 (O_247,N_3862,N_3559);
nand UO_248 (O_248,N_4955,N_3341);
xor UO_249 (O_249,N_3918,N_4140);
or UO_250 (O_250,N_4736,N_4479);
and UO_251 (O_251,N_3783,N_3647);
xnor UO_252 (O_252,N_4279,N_4796);
nand UO_253 (O_253,N_4104,N_3351);
or UO_254 (O_254,N_3164,N_3540);
nand UO_255 (O_255,N_2880,N_3491);
nand UO_256 (O_256,N_4598,N_3202);
or UO_257 (O_257,N_4444,N_4888);
and UO_258 (O_258,N_3340,N_4642);
xor UO_259 (O_259,N_2750,N_4663);
nand UO_260 (O_260,N_4647,N_2765);
and UO_261 (O_261,N_4272,N_4789);
and UO_262 (O_262,N_3954,N_4368);
nand UO_263 (O_263,N_3097,N_3701);
and UO_264 (O_264,N_3208,N_2650);
and UO_265 (O_265,N_4695,N_4529);
and UO_266 (O_266,N_3488,N_3777);
xnor UO_267 (O_267,N_4131,N_3883);
xor UO_268 (O_268,N_3151,N_4759);
and UO_269 (O_269,N_4179,N_4344);
or UO_270 (O_270,N_3209,N_3396);
nand UO_271 (O_271,N_4057,N_4364);
nand UO_272 (O_272,N_4970,N_4775);
or UO_273 (O_273,N_3831,N_4941);
or UO_274 (O_274,N_3686,N_3241);
nor UO_275 (O_275,N_4690,N_3039);
nand UO_276 (O_276,N_4224,N_4528);
nand UO_277 (O_277,N_4048,N_3450);
nand UO_278 (O_278,N_3178,N_4437);
or UO_279 (O_279,N_2929,N_2556);
or UO_280 (O_280,N_3947,N_4391);
and UO_281 (O_281,N_3480,N_3437);
nand UO_282 (O_282,N_3838,N_3962);
nor UO_283 (O_283,N_3320,N_3334);
and UO_284 (O_284,N_4115,N_4831);
and UO_285 (O_285,N_2713,N_3595);
xor UO_286 (O_286,N_3103,N_3009);
nor UO_287 (O_287,N_2755,N_3612);
or UO_288 (O_288,N_3924,N_4619);
and UO_289 (O_289,N_4094,N_4940);
nor UO_290 (O_290,N_4184,N_3219);
nand UO_291 (O_291,N_3158,N_4078);
nor UO_292 (O_292,N_3987,N_4822);
nand UO_293 (O_293,N_2595,N_3301);
nor UO_294 (O_294,N_2657,N_3400);
nand UO_295 (O_295,N_2611,N_4836);
nand UO_296 (O_296,N_3724,N_4933);
nand UO_297 (O_297,N_3754,N_3075);
xor UO_298 (O_298,N_4258,N_4714);
or UO_299 (O_299,N_4366,N_3456);
nand UO_300 (O_300,N_4083,N_3774);
nor UO_301 (O_301,N_3606,N_4767);
and UO_302 (O_302,N_2824,N_4992);
nand UO_303 (O_303,N_3955,N_2862);
or UO_304 (O_304,N_4309,N_3365);
or UO_305 (O_305,N_3825,N_3270);
or UO_306 (O_306,N_4961,N_4348);
nor UO_307 (O_307,N_3237,N_3679);
nor UO_308 (O_308,N_2748,N_4266);
or UO_309 (O_309,N_4434,N_4093);
and UO_310 (O_310,N_4036,N_4220);
or UO_311 (O_311,N_3909,N_3671);
or UO_312 (O_312,N_2836,N_2926);
nor UO_313 (O_313,N_3515,N_3643);
and UO_314 (O_314,N_4035,N_4286);
or UO_315 (O_315,N_4669,N_4001);
nor UO_316 (O_316,N_2835,N_3140);
nor UO_317 (O_317,N_3910,N_2654);
nand UO_318 (O_318,N_4890,N_3742);
nand UO_319 (O_319,N_4486,N_3813);
or UO_320 (O_320,N_3965,N_4928);
and UO_321 (O_321,N_2842,N_4480);
nand UO_322 (O_322,N_2790,N_3027);
nand UO_323 (O_323,N_3262,N_2565);
or UO_324 (O_324,N_3654,N_4648);
xnor UO_325 (O_325,N_2558,N_2949);
or UO_326 (O_326,N_3089,N_4952);
nor UO_327 (O_327,N_2940,N_2804);
nand UO_328 (O_328,N_2944,N_2642);
or UO_329 (O_329,N_3945,N_3510);
and UO_330 (O_330,N_4136,N_4981);
nand UO_331 (O_331,N_4751,N_4526);
or UO_332 (O_332,N_2662,N_4269);
xnor UO_333 (O_333,N_4956,N_3556);
nor UO_334 (O_334,N_2965,N_3311);
or UO_335 (O_335,N_3836,N_2897);
nor UO_336 (O_336,N_2909,N_4111);
nand UO_337 (O_337,N_3966,N_4866);
nand UO_338 (O_338,N_2681,N_3233);
and UO_339 (O_339,N_4954,N_4996);
or UO_340 (O_340,N_2559,N_2993);
and UO_341 (O_341,N_3368,N_3669);
nor UO_342 (O_342,N_4914,N_3132);
xor UO_343 (O_343,N_3080,N_2560);
or UO_344 (O_344,N_4778,N_2737);
or UO_345 (O_345,N_3874,N_2970);
nor UO_346 (O_346,N_3937,N_4632);
or UO_347 (O_347,N_3432,N_3705);
or UO_348 (O_348,N_4105,N_4768);
and UO_349 (O_349,N_3522,N_3094);
xor UO_350 (O_350,N_3086,N_3729);
or UO_351 (O_351,N_4385,N_3551);
or UO_352 (O_352,N_2817,N_3963);
nand UO_353 (O_353,N_2775,N_4677);
nor UO_354 (O_354,N_2814,N_3122);
or UO_355 (O_355,N_3226,N_2934);
nand UO_356 (O_356,N_4636,N_3650);
nor UO_357 (O_357,N_2859,N_4510);
nor UO_358 (O_358,N_3484,N_4338);
nand UO_359 (O_359,N_4681,N_4124);
nor UO_360 (O_360,N_3044,N_2758);
and UO_361 (O_361,N_4303,N_3949);
nand UO_362 (O_362,N_4328,N_3232);
and UO_363 (O_363,N_3604,N_3247);
nand UO_364 (O_364,N_3261,N_4354);
nand UO_365 (O_365,N_3867,N_3845);
or UO_366 (O_366,N_3789,N_2534);
nand UO_367 (O_367,N_4592,N_4830);
or UO_368 (O_368,N_2885,N_2923);
and UO_369 (O_369,N_4333,N_3853);
or UO_370 (O_370,N_4745,N_2668);
nand UO_371 (O_371,N_4080,N_4493);
nand UO_372 (O_372,N_2751,N_3411);
nand UO_373 (O_373,N_4589,N_3591);
nand UO_374 (O_374,N_2525,N_4428);
and UO_375 (O_375,N_3525,N_3238);
and UO_376 (O_376,N_2964,N_4710);
or UO_377 (O_377,N_4942,N_3625);
nor UO_378 (O_378,N_3687,N_3901);
nor UO_379 (O_379,N_3917,N_3302);
or UO_380 (O_380,N_2952,N_4064);
nand UO_381 (O_381,N_4463,N_4090);
and UO_382 (O_382,N_3200,N_3215);
nor UO_383 (O_383,N_4904,N_4500);
xor UO_384 (O_384,N_4120,N_3902);
nand UO_385 (O_385,N_3123,N_3008);
nor UO_386 (O_386,N_2887,N_2797);
nor UO_387 (O_387,N_4291,N_3125);
and UO_388 (O_388,N_3849,N_4810);
or UO_389 (O_389,N_3493,N_4494);
and UO_390 (O_390,N_2695,N_3921);
or UO_391 (O_391,N_4630,N_3218);
and UO_392 (O_392,N_3895,N_3459);
nand UO_393 (O_393,N_4401,N_2955);
nand UO_394 (O_394,N_4932,N_4638);
or UO_395 (O_395,N_2505,N_3188);
nand UO_396 (O_396,N_4635,N_3370);
or UO_397 (O_397,N_3322,N_2546);
or UO_398 (O_398,N_4483,N_3026);
nor UO_399 (O_399,N_3195,N_4372);
and UO_400 (O_400,N_4427,N_3781);
xnor UO_401 (O_401,N_4321,N_4242);
and UO_402 (O_402,N_4913,N_3518);
nand UO_403 (O_403,N_3055,N_3586);
or UO_404 (O_404,N_2849,N_4887);
nand UO_405 (O_405,N_3624,N_3444);
or UO_406 (O_406,N_2942,N_4655);
nor UO_407 (O_407,N_4467,N_4314);
nand UO_408 (O_408,N_3271,N_4509);
nand UO_409 (O_409,N_3222,N_3585);
or UO_410 (O_410,N_3108,N_2744);
or UO_411 (O_411,N_2741,N_3445);
nor UO_412 (O_412,N_2900,N_4837);
nor UO_413 (O_413,N_2557,N_4840);
or UO_414 (O_414,N_4585,N_4270);
nor UO_415 (O_415,N_3903,N_3290);
and UO_416 (O_416,N_4284,N_3731);
nand UO_417 (O_417,N_2513,N_3552);
and UO_418 (O_418,N_3865,N_2547);
nand UO_419 (O_419,N_3300,N_4612);
xor UO_420 (O_420,N_4790,N_3827);
nor UO_421 (O_421,N_4545,N_2640);
nor UO_422 (O_422,N_3553,N_4785);
nor UO_423 (O_423,N_4686,N_2571);
nand UO_424 (O_424,N_4993,N_3422);
and UO_425 (O_425,N_4734,N_3014);
nor UO_426 (O_426,N_3330,N_2579);
and UO_427 (O_427,N_2663,N_3795);
nand UO_428 (O_428,N_2671,N_4508);
nand UO_429 (O_429,N_3916,N_3938);
nor UO_430 (O_430,N_3683,N_2907);
nand UO_431 (O_431,N_3043,N_3779);
or UO_432 (O_432,N_3439,N_4679);
and UO_433 (O_433,N_4400,N_3284);
nor UO_434 (O_434,N_4394,N_4138);
nor UO_435 (O_435,N_4616,N_3919);
and UO_436 (O_436,N_3428,N_4022);
or UO_437 (O_437,N_4055,N_2935);
xor UO_438 (O_438,N_3863,N_4310);
nand UO_439 (O_439,N_4564,N_3583);
and UO_440 (O_440,N_4550,N_2503);
nor UO_441 (O_441,N_3621,N_4502);
xnor UO_442 (O_442,N_3224,N_2731);
or UO_443 (O_443,N_3332,N_4621);
nand UO_444 (O_444,N_2984,N_3538);
xor UO_445 (O_445,N_2903,N_4722);
or UO_446 (O_446,N_3479,N_3850);
and UO_447 (O_447,N_4488,N_4037);
and UO_448 (O_448,N_3424,N_3083);
nand UO_449 (O_449,N_3032,N_2834);
nor UO_450 (O_450,N_2517,N_4389);
nand UO_451 (O_451,N_3216,N_3379);
and UO_452 (O_452,N_4735,N_4577);
xor UO_453 (O_453,N_4746,N_3461);
and UO_454 (O_454,N_4884,N_3761);
and UO_455 (O_455,N_2912,N_2734);
xor UO_456 (O_456,N_2840,N_3230);
nand UO_457 (O_457,N_3699,N_3010);
xor UO_458 (O_458,N_4232,N_4225);
and UO_459 (O_459,N_4968,N_4365);
and UO_460 (O_460,N_4281,N_3942);
nor UO_461 (O_461,N_4631,N_3837);
xnor UO_462 (O_462,N_4779,N_2609);
xnor UO_463 (O_463,N_4311,N_4760);
and UO_464 (O_464,N_4853,N_4869);
nand UO_465 (O_465,N_4824,N_3596);
and UO_466 (O_466,N_2531,N_4472);
and UO_467 (O_467,N_2910,N_3582);
and UO_468 (O_468,N_4896,N_3617);
and UO_469 (O_469,N_3511,N_2868);
nand UO_470 (O_470,N_2522,N_2569);
nor UO_471 (O_471,N_2888,N_3474);
or UO_472 (O_472,N_4758,N_3709);
nor UO_473 (O_473,N_3163,N_3433);
xor UO_474 (O_474,N_4889,N_4011);
nor UO_475 (O_475,N_4675,N_3869);
xor UO_476 (O_476,N_2788,N_2705);
xor UO_477 (O_477,N_4773,N_4327);
or UO_478 (O_478,N_3282,N_4676);
nand UO_479 (O_479,N_4330,N_3328);
xor UO_480 (O_480,N_3651,N_3088);
nor UO_481 (O_481,N_3240,N_2959);
or UO_482 (O_482,N_3412,N_3213);
or UO_483 (O_483,N_4165,N_4755);
nor UO_484 (O_484,N_3152,N_2978);
or UO_485 (O_485,N_4762,N_2881);
and UO_486 (O_486,N_3186,N_4555);
nor UO_487 (O_487,N_2645,N_2792);
nor UO_488 (O_488,N_3532,N_3149);
xnor UO_489 (O_489,N_4953,N_3248);
or UO_490 (O_490,N_4219,N_3374);
or UO_491 (O_491,N_4944,N_3335);
and UO_492 (O_492,N_3978,N_3114);
or UO_493 (O_493,N_2783,N_4233);
and UO_494 (O_494,N_3786,N_2953);
nor UO_495 (O_495,N_4426,N_3812);
nand UO_496 (O_496,N_4895,N_3505);
nand UO_497 (O_497,N_4947,N_4227);
nand UO_498 (O_498,N_3259,N_2625);
nand UO_499 (O_499,N_2774,N_2717);
nand UO_500 (O_500,N_2605,N_4393);
and UO_501 (O_501,N_2591,N_4381);
and UO_502 (O_502,N_2861,N_4458);
xnor UO_503 (O_503,N_2908,N_4798);
and UO_504 (O_504,N_4063,N_3214);
or UO_505 (O_505,N_3193,N_3663);
nor UO_506 (O_506,N_2791,N_4919);
nor UO_507 (O_507,N_3494,N_2895);
xnor UO_508 (O_508,N_3707,N_4424);
and UO_509 (O_509,N_4367,N_3759);
or UO_510 (O_510,N_3130,N_3832);
or UO_511 (O_511,N_2615,N_3468);
and UO_512 (O_512,N_4723,N_2687);
or UO_513 (O_513,N_4106,N_3068);
or UO_514 (O_514,N_4039,N_4674);
nand UO_515 (O_515,N_3983,N_2618);
or UO_516 (O_516,N_4691,N_3513);
or UO_517 (O_517,N_3058,N_4313);
and UO_518 (O_518,N_3730,N_3436);
nor UO_519 (O_519,N_3716,N_3427);
and UO_520 (O_520,N_2582,N_2967);
and UO_521 (O_521,N_4222,N_3413);
and UO_522 (O_522,N_4670,N_4118);
xnor UO_523 (O_523,N_3402,N_3659);
or UO_524 (O_524,N_2992,N_4541);
and UO_525 (O_525,N_3021,N_2962);
nor UO_526 (O_526,N_3740,N_3886);
nor UO_527 (O_527,N_3418,N_4809);
xnor UO_528 (O_528,N_2892,N_4041);
or UO_529 (O_529,N_4380,N_4377);
nor UO_530 (O_530,N_4911,N_4277);
nor UO_531 (O_531,N_2749,N_4595);
nand UO_532 (O_532,N_4148,N_2590);
xnor UO_533 (O_533,N_3136,N_2538);
nor UO_534 (O_534,N_2568,N_4848);
nand UO_535 (O_535,N_3711,N_4938);
xnor UO_536 (O_536,N_2697,N_3818);
nor UO_537 (O_537,N_2689,N_4696);
or UO_538 (O_538,N_4192,N_4871);
nand UO_539 (O_539,N_4701,N_4977);
nand UO_540 (O_540,N_2716,N_3475);
or UO_541 (O_541,N_3430,N_3644);
or UO_542 (O_542,N_2832,N_3534);
nand UO_543 (O_543,N_4742,N_3404);
nor UO_544 (O_544,N_3166,N_3012);
and UO_545 (O_545,N_4851,N_3857);
xor UO_546 (O_546,N_4496,N_4019);
or UO_547 (O_547,N_4862,N_3684);
or UO_548 (O_548,N_4300,N_2530);
and UO_549 (O_549,N_3720,N_3822);
nor UO_550 (O_550,N_3472,N_4917);
xnor UO_551 (O_551,N_4260,N_3636);
or UO_552 (O_552,N_4936,N_3131);
nor UO_553 (O_553,N_3765,N_3633);
or UO_554 (O_554,N_4925,N_2882);
and UO_555 (O_555,N_4289,N_4034);
and UO_556 (O_556,N_2543,N_3968);
nand UO_557 (O_557,N_2739,N_3933);
nand UO_558 (O_558,N_2779,N_2733);
nand UO_559 (O_559,N_4100,N_4659);
xnor UO_560 (O_560,N_4198,N_2760);
or UO_561 (O_561,N_4290,N_3710);
nor UO_562 (O_562,N_3337,N_4532);
nand UO_563 (O_563,N_4079,N_3096);
or UO_564 (O_564,N_3984,N_3253);
nor UO_565 (O_565,N_2566,N_3381);
nor UO_566 (O_566,N_4668,N_4600);
nand UO_567 (O_567,N_2898,N_4503);
and UO_568 (O_568,N_3890,N_3605);
or UO_569 (O_569,N_4572,N_4433);
or UO_570 (O_570,N_2770,N_4558);
or UO_571 (O_571,N_3744,N_4446);
and UO_572 (O_572,N_3279,N_3421);
or UO_573 (O_573,N_2720,N_4464);
nor UO_574 (O_574,N_3769,N_3563);
nand UO_575 (O_575,N_3611,N_4639);
or UO_576 (O_576,N_2541,N_3171);
or UO_577 (O_577,N_3851,N_2946);
xnor UO_578 (O_578,N_4141,N_2869);
and UO_579 (O_579,N_4236,N_3111);
nor UO_580 (O_580,N_4605,N_3704);
or UO_581 (O_581,N_4845,N_3572);
or UO_582 (O_582,N_2939,N_4945);
nor UO_583 (O_583,N_4008,N_4772);
and UO_584 (O_584,N_4294,N_3397);
nand UO_585 (O_585,N_3142,N_4703);
nand UO_586 (O_586,N_4692,N_4660);
nor UO_587 (O_587,N_4971,N_3106);
and UO_588 (O_588,N_3784,N_3639);
or UO_589 (O_589,N_2528,N_3324);
nand UO_590 (O_590,N_3613,N_2777);
xor UO_591 (O_591,N_3327,N_4084);
xor UO_592 (O_592,N_2956,N_4905);
and UO_593 (O_593,N_4108,N_3137);
nor UO_594 (O_594,N_3318,N_3167);
or UO_595 (O_595,N_3509,N_2507);
nand UO_596 (O_596,N_3879,N_2725);
nor UO_597 (O_597,N_4799,N_4320);
nor UO_598 (O_598,N_3528,N_3506);
and UO_599 (O_599,N_4095,N_4167);
or UO_600 (O_600,N_4243,N_2648);
nand UO_601 (O_601,N_4622,N_4586);
nand UO_602 (O_602,N_4490,N_4316);
xor UO_603 (O_603,N_4371,N_4623);
and UO_604 (O_604,N_4957,N_4519);
and UO_605 (O_605,N_4047,N_3571);
nand UO_606 (O_606,N_3229,N_4499);
and UO_607 (O_607,N_2866,N_3203);
and UO_608 (O_608,N_3464,N_2930);
xnor UO_609 (O_609,N_4861,N_3256);
and UO_610 (O_610,N_2647,N_2693);
nand UO_611 (O_611,N_4832,N_2971);
or UO_612 (O_612,N_3455,N_3531);
or UO_613 (O_613,N_2698,N_3576);
or UO_614 (O_614,N_3319,N_2968);
nor UO_615 (O_615,N_3566,N_4504);
and UO_616 (O_616,N_4581,N_3157);
and UO_617 (O_617,N_2532,N_2694);
or UO_618 (O_618,N_2987,N_3516);
or UO_619 (O_619,N_4579,N_3499);
or UO_620 (O_620,N_2798,N_4918);
and UO_621 (O_621,N_4803,N_4172);
or UO_622 (O_622,N_4780,N_3763);
and UO_623 (O_623,N_2846,N_2894);
nand UO_624 (O_624,N_2966,N_4392);
nand UO_625 (O_625,N_4731,N_3665);
nand UO_626 (O_626,N_2938,N_4436);
and UO_627 (O_627,N_4787,N_4908);
nor UO_628 (O_628,N_3810,N_4182);
nand UO_629 (O_629,N_3842,N_4757);
nand UO_630 (O_630,N_2950,N_4031);
nand UO_631 (O_631,N_3884,N_2786);
nand UO_632 (O_632,N_3489,N_3062);
nor UO_633 (O_633,N_2860,N_3153);
and UO_634 (O_634,N_3715,N_4673);
nor UO_635 (O_635,N_3321,N_4370);
and UO_636 (O_636,N_3228,N_3079);
xnor UO_637 (O_637,N_4578,N_2710);
or UO_638 (O_638,N_4743,N_4353);
nand UO_639 (O_639,N_3100,N_3957);
and UO_640 (O_640,N_4833,N_3974);
nand UO_641 (O_641,N_4930,N_3577);
nand UO_642 (O_642,N_2829,N_2691);
or UO_643 (O_643,N_3323,N_2856);
nor UO_644 (O_644,N_3391,N_3875);
nand UO_645 (O_645,N_3053,N_3460);
nand UO_646 (O_646,N_2551,N_3988);
or UO_647 (O_647,N_3914,N_3471);
and UO_648 (O_648,N_2816,N_3964);
and UO_649 (O_649,N_4983,N_4582);
nand UO_650 (O_650,N_4769,N_4126);
nand UO_651 (O_651,N_3618,N_3072);
or UO_652 (O_652,N_4812,N_3632);
or UO_653 (O_653,N_2936,N_3031);
and UO_654 (O_654,N_3343,N_4230);
nand UO_655 (O_655,N_2977,N_4248);
nor UO_656 (O_656,N_4927,N_3598);
and UO_657 (O_657,N_4210,N_4276);
xnor UO_658 (O_658,N_3575,N_4183);
nor UO_659 (O_659,N_4929,N_4643);
xor UO_660 (O_660,N_3254,N_2853);
nor UO_661 (O_661,N_2604,N_3476);
and UO_662 (O_662,N_4697,N_4985);
nand UO_663 (O_663,N_2680,N_4596);
or UO_664 (O_664,N_2948,N_3519);
nor UO_665 (O_665,N_2837,N_4262);
and UO_666 (O_666,N_4535,N_4340);
xor UO_667 (O_667,N_4517,N_4403);
nor UO_668 (O_668,N_3725,N_4516);
nor UO_669 (O_669,N_4117,N_3501);
or UO_670 (O_670,N_4664,N_4620);
and UO_671 (O_671,N_2638,N_3861);
and UO_672 (O_672,N_4145,N_3833);
and UO_673 (O_673,N_2621,N_3463);
nand UO_674 (O_674,N_2552,N_2619);
and UO_675 (O_675,N_2879,N_4943);
nand UO_676 (O_676,N_2686,N_3281);
or UO_677 (O_677,N_3217,N_3220);
nand UO_678 (O_678,N_4122,N_4491);
xnor UO_679 (O_679,N_3764,N_4567);
nand UO_680 (O_680,N_4254,N_3891);
and UO_681 (O_681,N_4163,N_2913);
or UO_682 (O_682,N_4497,N_3326);
and UO_683 (O_683,N_3092,N_2850);
and UO_684 (O_684,N_3045,N_4637);
or UO_685 (O_685,N_4457,N_2756);
or UO_686 (O_686,N_4823,N_3184);
nor UO_687 (O_687,N_3498,N_2914);
and UO_688 (O_688,N_4950,N_4410);
nor UO_689 (O_689,N_4886,N_4214);
and UO_690 (O_690,N_3693,N_4800);
nand UO_691 (O_691,N_4181,N_4774);
or UO_692 (O_692,N_3943,N_3173);
or UO_693 (O_693,N_3273,N_4246);
nand UO_694 (O_694,N_4522,N_2690);
and UO_695 (O_695,N_2809,N_3645);
and UO_696 (O_696,N_3183,N_4206);
and UO_697 (O_697,N_4680,N_4498);
or UO_698 (O_698,N_4087,N_4994);
nor UO_699 (O_699,N_2684,N_4476);
nand UO_700 (O_700,N_4204,N_2889);
and UO_701 (O_701,N_3325,N_3211);
nand UO_702 (O_702,N_4004,N_3817);
and UO_703 (O_703,N_3970,N_4038);
or UO_704 (O_704,N_4419,N_4902);
nand UO_705 (O_705,N_2773,N_3447);
and UO_706 (O_706,N_4471,N_3144);
nand UO_707 (O_707,N_4174,N_4724);
and UO_708 (O_708,N_3871,N_3996);
nor UO_709 (O_709,N_3899,N_4226);
nor UO_710 (O_710,N_4396,N_3449);
or UO_711 (O_711,N_4070,N_3278);
nand UO_712 (O_712,N_3941,N_2711);
nor UO_713 (O_713,N_4959,N_4139);
and UO_714 (O_714,N_3189,N_3194);
nor UO_715 (O_715,N_4096,N_4194);
nand UO_716 (O_716,N_3882,N_3578);
xnor UO_717 (O_717,N_4349,N_3855);
nand UO_718 (O_718,N_2886,N_3628);
or UO_719 (O_719,N_3112,N_2875);
nand UO_720 (O_720,N_4492,N_3362);
or UO_721 (O_721,N_4650,N_4543);
and UO_722 (O_722,N_3386,N_4877);
and UO_723 (O_723,N_4049,N_3939);
xnor UO_724 (O_724,N_4355,N_3713);
or UO_725 (O_725,N_4156,N_4102);
nand UO_726 (O_726,N_4556,N_4134);
and UO_727 (O_727,N_4166,N_4552);
or UO_728 (O_728,N_3998,N_3829);
and UO_729 (O_729,N_2637,N_2822);
and UO_730 (O_730,N_4513,N_4573);
or UO_731 (O_731,N_3223,N_3664);
or UO_732 (O_732,N_3497,N_3703);
xnor UO_733 (O_733,N_4649,N_3352);
nand UO_734 (O_734,N_3719,N_3162);
nor UO_735 (O_735,N_3627,N_3608);
xor UO_736 (O_736,N_2819,N_4707);
or UO_737 (O_737,N_4306,N_2989);
nor UO_738 (O_738,N_4920,N_4416);
nand UO_739 (O_739,N_3561,N_3065);
nor UO_740 (O_740,N_2537,N_3061);
or UO_741 (O_741,N_3517,N_3181);
nor UO_742 (O_742,N_3357,N_2708);
and UO_743 (O_743,N_4361,N_4026);
nand UO_744 (O_744,N_4580,N_3375);
or UO_745 (O_745,N_3811,N_2564);
nor UO_746 (O_746,N_2669,N_4342);
nor UO_747 (O_747,N_4666,N_3688);
nand UO_748 (O_748,N_3992,N_4607);
nor UO_749 (O_749,N_4625,N_4817);
or UO_750 (O_750,N_2613,N_2683);
nand UO_751 (O_751,N_3084,N_3134);
and UO_752 (O_752,N_2937,N_4208);
or UO_753 (O_753,N_3143,N_2655);
nand UO_754 (O_754,N_4252,N_4854);
and UO_755 (O_755,N_3057,N_3107);
and UO_756 (O_756,N_4560,N_2519);
nor UO_757 (O_757,N_3533,N_2985);
nand UO_758 (O_758,N_2905,N_4728);
or UO_759 (O_759,N_3539,N_2764);
nor UO_760 (O_760,N_4009,N_4753);
xnor UO_761 (O_761,N_2979,N_4438);
or UO_762 (O_762,N_4583,N_4872);
and UO_763 (O_763,N_3801,N_2825);
or UO_764 (O_764,N_3907,N_2702);
and UO_765 (O_765,N_4409,N_4351);
or UO_766 (O_766,N_3369,N_4164);
and UO_767 (O_767,N_2581,N_4878);
nand UO_768 (O_768,N_3361,N_4273);
nor UO_769 (O_769,N_3292,N_2617);
nor UO_770 (O_770,N_4451,N_4747);
nor UO_771 (O_771,N_2608,N_3384);
and UO_772 (O_772,N_4608,N_3834);
xnor UO_773 (O_773,N_3129,N_3752);
xnor UO_774 (O_774,N_2986,N_3064);
nand UO_775 (O_775,N_3101,N_4784);
nand UO_776 (O_776,N_4114,N_4245);
and UO_777 (O_777,N_3104,N_4398);
nor UO_778 (O_778,N_4412,N_4525);
nor UO_779 (O_779,N_3458,N_4654);
or UO_780 (O_780,N_4448,N_4405);
nor UO_781 (O_781,N_2784,N_4470);
and UO_782 (O_782,N_3492,N_4133);
and UO_783 (O_783,N_4718,N_3994);
and UO_784 (O_784,N_4975,N_4531);
nor UO_785 (O_785,N_4071,N_3925);
or UO_786 (O_786,N_4125,N_2843);
nand UO_787 (O_787,N_3036,N_3926);
and UO_788 (O_788,N_3735,N_4706);
or UO_789 (O_789,N_4159,N_4629);
nand UO_790 (O_790,N_4211,N_3888);
nand UO_791 (O_791,N_4808,N_3756);
nand UO_792 (O_792,N_2586,N_2920);
or UO_793 (O_793,N_4142,N_2601);
or UO_794 (O_794,N_4923,N_2509);
and UO_795 (O_795,N_2549,N_3614);
and UO_796 (O_796,N_3877,N_3681);
nor UO_797 (O_797,N_2562,N_2805);
nor UO_798 (O_798,N_3993,N_3110);
nand UO_799 (O_799,N_3082,N_4575);
nand UO_800 (O_800,N_2795,N_3753);
nor UO_801 (O_801,N_4879,N_3041);
and UO_802 (O_802,N_4829,N_3581);
and UO_803 (O_803,N_4119,N_2624);
nor UO_804 (O_804,N_3870,N_2550);
xnor UO_805 (O_805,N_3897,N_3049);
nand UO_806 (O_806,N_2830,N_3019);
and UO_807 (O_807,N_3312,N_4374);
nand UO_808 (O_808,N_4750,N_4253);
nor UO_809 (O_809,N_2699,N_4112);
nor UO_810 (O_810,N_2752,N_4025);
nor UO_811 (O_811,N_4788,N_4804);
or UO_812 (O_812,N_4054,N_3889);
nor UO_813 (O_813,N_2732,N_4435);
or UO_814 (O_814,N_2906,N_4305);
and UO_815 (O_815,N_3793,N_3442);
nand UO_816 (O_816,N_4170,N_4549);
nor UO_817 (O_817,N_4014,N_2644);
xor UO_818 (O_818,N_4641,N_2524);
xor UO_819 (O_819,N_4256,N_3641);
nor UO_820 (O_820,N_4752,N_2514);
and UO_821 (O_821,N_2585,N_4323);
nand UO_822 (O_822,N_3347,N_4175);
xnor UO_823 (O_823,N_3473,N_4912);
or UO_824 (O_824,N_4021,N_2999);
nor UO_825 (O_825,N_3245,N_2820);
or UO_826 (O_826,N_3658,N_4143);
or UO_827 (O_827,N_4050,N_3792);
or UO_828 (O_828,N_4524,N_4147);
and UO_829 (O_829,N_4185,N_3805);
or UO_830 (O_830,N_4838,N_4827);
nand UO_831 (O_831,N_4129,N_3741);
nor UO_832 (O_832,N_4329,N_3185);
xor UO_833 (O_833,N_3905,N_2700);
or UO_834 (O_834,N_4285,N_4900);
nand UO_835 (O_835,N_4749,N_2851);
or UO_836 (O_836,N_4414,N_2960);
nand UO_837 (O_837,N_4990,N_4193);
or UO_838 (O_838,N_4109,N_3652);
or UO_839 (O_839,N_3898,N_4792);
nand UO_840 (O_840,N_4880,N_4379);
xor UO_841 (O_841,N_2871,N_2917);
or UO_842 (O_842,N_3168,N_4296);
xnor UO_843 (O_843,N_3392,N_4667);
nor UO_844 (O_844,N_4356,N_2980);
nor UO_845 (O_845,N_2766,N_2800);
nor UO_846 (O_846,N_4978,N_2995);
nand UO_847 (O_847,N_3394,N_3609);
nor UO_848 (O_848,N_3689,N_4288);
nand UO_849 (O_849,N_3490,N_4144);
xor UO_850 (O_850,N_4874,N_4726);
or UO_851 (O_851,N_3135,N_4569);
nor UO_852 (O_852,N_4934,N_2616);
and UO_853 (O_853,N_2893,N_3738);
nand UO_854 (O_854,N_3872,N_4298);
nor UO_855 (O_855,N_4865,N_3467);
or UO_856 (O_856,N_3006,N_2958);
or UO_857 (O_857,N_4501,N_2634);
nor UO_858 (O_858,N_4748,N_2596);
nor UO_859 (O_859,N_4937,N_2831);
and UO_860 (O_860,N_3580,N_3205);
nor UO_861 (O_861,N_3946,N_4282);
and UO_862 (O_862,N_3037,N_3210);
nor UO_863 (O_863,N_3852,N_3035);
or UO_864 (O_864,N_3634,N_2706);
nor UO_865 (O_865,N_3398,N_2884);
or UO_866 (O_866,N_4015,N_2555);
or UO_867 (O_867,N_2943,N_4593);
nor UO_868 (O_868,N_3267,N_2599);
nor UO_869 (O_869,N_4099,N_2975);
or UO_870 (O_870,N_4388,N_3236);
nor UO_871 (O_871,N_4010,N_3864);
nor UO_872 (O_872,N_3028,N_4137);
and UO_873 (O_873,N_4430,N_4076);
and UO_874 (O_874,N_4334,N_3649);
and UO_875 (O_875,N_4534,N_4777);
and UO_876 (O_876,N_4613,N_4763);
nand UO_877 (O_877,N_3776,N_4964);
or UO_878 (O_878,N_3289,N_4003);
xnor UO_879 (O_879,N_4665,N_4852);
nor UO_880 (O_880,N_2821,N_3212);
and UO_881 (O_881,N_4783,N_3280);
xnor UO_882 (O_882,N_3991,N_4103);
and UO_883 (O_883,N_4614,N_3935);
or UO_884 (O_884,N_3199,N_2901);
nor UO_885 (O_885,N_2998,N_2924);
xor UO_886 (O_886,N_2606,N_4378);
nand UO_887 (O_887,N_2526,N_3102);
nand UO_888 (O_888,N_3466,N_3285);
nor UO_889 (O_889,N_4883,N_4127);
nand UO_890 (O_890,N_3878,N_3034);
nor UO_891 (O_891,N_3961,N_3631);
nand UO_892 (O_892,N_2848,N_3762);
and UO_893 (O_893,N_2628,N_3589);
nor UO_894 (O_894,N_3723,N_3124);
nand UO_895 (O_895,N_3385,N_3054);
xnor UO_896 (O_896,N_3095,N_4449);
xnor UO_897 (O_897,N_4948,N_2576);
nor UO_898 (O_898,N_4097,N_3997);
xnor UO_899 (O_899,N_4744,N_3148);
nand UO_900 (O_900,N_4967,N_4921);
or UO_901 (O_901,N_4965,N_4969);
or UO_902 (O_902,N_3367,N_3349);
nor UO_903 (O_903,N_3600,N_3986);
nor UO_904 (O_904,N_3601,N_3141);
and UO_905 (O_905,N_4986,N_2932);
and UO_906 (O_906,N_3502,N_3310);
or UO_907 (O_907,N_4843,N_3900);
and UO_908 (O_908,N_3529,N_3393);
and UO_909 (O_909,N_2504,N_3074);
nand UO_910 (O_910,N_3283,N_3999);
xnor UO_911 (O_911,N_2746,N_3920);
or UO_912 (O_912,N_4207,N_3165);
or UO_913 (O_913,N_2921,N_4293);
nor UO_914 (O_914,N_2983,N_2709);
nand UO_915 (O_915,N_4399,N_2812);
nand UO_916 (O_916,N_4152,N_2589);
nor UO_917 (O_917,N_4835,N_2742);
and UO_918 (O_918,N_3469,N_3696);
nor UO_919 (O_919,N_4062,N_4873);
or UO_920 (O_920,N_4511,N_3526);
nor UO_921 (O_921,N_4216,N_3077);
nor UO_922 (O_922,N_4587,N_3116);
nand UO_923 (O_923,N_4081,N_4807);
nand UO_924 (O_924,N_3594,N_4265);
or UO_925 (O_925,N_3500,N_2622);
or UO_926 (O_926,N_4336,N_4363);
or UO_927 (O_927,N_3277,N_3588);
nor UO_928 (O_928,N_3052,N_2743);
nand UO_929 (O_929,N_2667,N_3814);
nand UO_930 (O_930,N_3854,N_3554);
and UO_931 (O_931,N_3950,N_3896);
nor UO_932 (O_932,N_2876,N_4709);
and UO_933 (O_933,N_4386,N_3906);
xor UO_934 (O_934,N_2620,N_3005);
nor UO_935 (O_935,N_4553,N_3033);
or UO_936 (O_936,N_2991,N_2845);
nand UO_937 (O_937,N_4033,N_2776);
or UO_938 (O_938,N_3348,N_3221);
xnor UO_939 (O_939,N_2899,N_3579);
nor UO_940 (O_940,N_4235,N_3746);
nand UO_941 (O_941,N_3677,N_4302);
nand UO_942 (O_942,N_3819,N_3788);
nor UO_943 (O_943,N_3296,N_2918);
and UO_944 (O_944,N_4113,N_4976);
and UO_945 (O_945,N_2703,N_4781);
nor UO_946 (O_946,N_4548,N_3547);
and UO_947 (O_947,N_4223,N_3366);
or UO_948 (O_948,N_4915,N_2916);
nor UO_949 (O_949,N_2878,N_3066);
nor UO_950 (O_950,N_4007,N_3718);
and UO_951 (O_951,N_4987,N_2945);
or UO_952 (O_952,N_4683,N_4907);
or UO_953 (O_953,N_3317,N_3521);
nand UO_954 (O_954,N_2988,N_4429);
nor UO_955 (O_955,N_3016,N_2810);
nor UO_956 (O_956,N_2548,N_4337);
and UO_957 (O_957,N_4721,N_3530);
nor UO_958 (O_958,N_4442,N_4512);
and UO_959 (O_959,N_3426,N_2833);
and UO_960 (O_960,N_3930,N_4200);
or UO_961 (O_961,N_2785,N_2511);
and UO_962 (O_962,N_4283,N_3726);
nand UO_963 (O_963,N_2961,N_4308);
nand UO_964 (O_964,N_2890,N_3297);
and UO_965 (O_965,N_3674,N_4563);
nor UO_966 (O_966,N_4771,N_2974);
or UO_967 (O_967,N_2580,N_4901);
or UO_968 (O_968,N_3670,N_4452);
nor UO_969 (O_969,N_2996,N_3736);
xor UO_970 (O_970,N_4418,N_4764);
and UO_971 (O_971,N_4839,N_4259);
and UO_972 (O_972,N_3405,N_2578);
nor UO_973 (O_973,N_3446,N_4173);
xor UO_974 (O_974,N_4218,N_4359);
xor UO_975 (O_975,N_4576,N_3204);
xnor UO_976 (O_976,N_4088,N_3275);
and UO_977 (O_977,N_4705,N_2553);
nand UO_978 (O_978,N_4634,N_4261);
or UO_979 (O_979,N_3768,N_3363);
nand UO_980 (O_980,N_4795,N_2767);
or UO_981 (O_981,N_4324,N_4909);
or UO_982 (O_982,N_2826,N_3496);
or UO_983 (O_983,N_2529,N_2665);
or UO_984 (O_984,N_3251,N_4468);
and UO_985 (O_985,N_2759,N_4640);
nand UO_986 (O_986,N_3557,N_3225);
nand UO_987 (O_987,N_3535,N_4251);
nor UO_988 (O_988,N_4439,N_3672);
and UO_989 (O_989,N_2633,N_4016);
or UO_990 (O_990,N_3481,N_3346);
nand UO_991 (O_991,N_3443,N_3081);
or UO_992 (O_992,N_4995,N_4046);
and UO_993 (O_993,N_4520,N_4687);
nor UO_994 (O_994,N_3160,N_4478);
nand UO_995 (O_995,N_2676,N_2806);
nor UO_996 (O_996,N_3673,N_3816);
nor UO_997 (O_997,N_3721,N_2501);
nand UO_998 (O_998,N_4092,N_3760);
nand UO_999 (O_999,N_4069,N_3425);
endmodule