module basic_5000_50000_5000_100_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
nand U0 (N_0,In_3608,In_2424);
or U1 (N_1,In_1091,In_2855);
and U2 (N_2,In_590,In_355);
and U3 (N_3,In_4569,In_3960);
or U4 (N_4,In_1905,In_2690);
or U5 (N_5,In_4050,In_2850);
xor U6 (N_6,In_3340,In_4890);
xor U7 (N_7,In_817,In_190);
or U8 (N_8,In_267,In_3638);
or U9 (N_9,In_3202,In_3426);
nand U10 (N_10,In_3856,In_2396);
or U11 (N_11,In_4754,In_2819);
xor U12 (N_12,In_3434,In_3447);
nand U13 (N_13,In_1391,In_3565);
and U14 (N_14,In_1356,In_137);
and U15 (N_15,In_3509,In_2746);
or U16 (N_16,In_483,In_3584);
nand U17 (N_17,In_1815,In_3421);
nor U18 (N_18,In_1267,In_4028);
xnor U19 (N_19,In_163,In_3508);
or U20 (N_20,In_2081,In_444);
nand U21 (N_21,In_2146,In_348);
nor U22 (N_22,In_2452,In_1529);
nor U23 (N_23,In_2769,In_618);
nand U24 (N_24,In_2135,In_143);
nand U25 (N_25,In_656,In_3236);
xor U26 (N_26,In_2817,In_3140);
and U27 (N_27,In_2831,In_138);
and U28 (N_28,In_2536,In_4611);
and U29 (N_29,In_4186,In_186);
xnor U30 (N_30,In_2744,In_4632);
nand U31 (N_31,In_1710,In_431);
nand U32 (N_32,In_4282,In_1385);
nor U33 (N_33,In_4230,In_2941);
nor U34 (N_34,In_241,In_3010);
and U35 (N_35,In_95,In_103);
nor U36 (N_36,In_4730,In_4276);
xnor U37 (N_37,In_2267,In_4659);
xnor U38 (N_38,In_3862,In_4289);
and U39 (N_39,In_10,In_819);
nor U40 (N_40,In_666,In_4597);
nand U41 (N_41,In_787,In_1641);
nand U42 (N_42,In_4766,In_4897);
xnor U43 (N_43,In_1266,In_2039);
and U44 (N_44,In_823,In_4059);
xor U45 (N_45,In_1310,In_4279);
or U46 (N_46,In_3507,In_1024);
or U47 (N_47,In_1735,In_1164);
xor U48 (N_48,In_721,In_2698);
or U49 (N_49,In_4086,In_3323);
or U50 (N_50,In_2503,In_2712);
or U51 (N_51,In_2641,In_4937);
or U52 (N_52,In_3785,In_958);
and U53 (N_53,In_4198,In_928);
nand U54 (N_54,In_3188,In_685);
xnor U55 (N_55,In_1280,In_3939);
xnor U56 (N_56,In_2372,In_852);
nand U57 (N_57,In_3320,In_556);
nor U58 (N_58,In_3784,In_3662);
xnor U59 (N_59,In_1471,In_1054);
nand U60 (N_60,In_3714,In_3838);
xor U61 (N_61,In_1602,In_3471);
or U62 (N_62,In_3542,In_1698);
and U63 (N_63,In_3123,In_408);
nand U64 (N_64,In_1574,In_2936);
or U65 (N_65,In_1006,In_2437);
and U66 (N_66,In_2117,In_460);
or U67 (N_67,In_2700,In_251);
nand U68 (N_68,In_3115,In_4610);
xor U69 (N_69,In_2799,In_4345);
nor U70 (N_70,In_1975,In_2792);
xnor U71 (N_71,In_3489,In_1742);
nor U72 (N_72,In_1775,In_2741);
and U73 (N_73,In_1493,In_719);
nor U74 (N_74,In_2136,In_2518);
xor U75 (N_75,In_2779,In_1963);
xnor U76 (N_76,In_1565,In_2269);
xnor U77 (N_77,In_2894,In_1635);
nand U78 (N_78,In_1467,In_2865);
and U79 (N_79,In_3443,In_932);
nor U80 (N_80,In_600,In_3316);
xor U81 (N_81,In_1432,In_3514);
or U82 (N_82,In_4614,In_689);
and U83 (N_83,In_4633,In_2988);
nor U84 (N_84,In_1382,In_136);
or U85 (N_85,In_114,In_2705);
and U86 (N_86,In_2410,In_151);
or U87 (N_87,In_257,In_2350);
and U88 (N_88,In_2376,In_1025);
xnor U89 (N_89,In_341,In_1509);
and U90 (N_90,In_651,In_2533);
nor U91 (N_91,In_4933,In_1611);
nand U92 (N_92,In_4110,In_1640);
nand U93 (N_93,In_4999,In_2360);
nor U94 (N_94,In_2822,In_829);
nor U95 (N_95,In_1646,In_1496);
nand U96 (N_96,In_3603,In_526);
and U97 (N_97,In_3308,In_1904);
nor U98 (N_98,In_3619,In_3522);
nor U99 (N_99,In_1053,In_3184);
nor U100 (N_100,In_1805,In_3494);
and U101 (N_101,In_4780,In_3807);
xor U102 (N_102,In_436,In_248);
and U103 (N_103,In_1533,In_4243);
nand U104 (N_104,In_3228,In_4866);
xnor U105 (N_105,In_2137,In_4562);
or U106 (N_106,In_2706,In_3457);
nand U107 (N_107,In_2930,In_2613);
nor U108 (N_108,In_1293,In_3212);
nand U109 (N_109,In_3691,In_2009);
or U110 (N_110,In_2773,In_1260);
nor U111 (N_111,In_1198,In_111);
nor U112 (N_112,In_2266,In_1779);
or U113 (N_113,In_1044,In_3346);
nor U114 (N_114,In_1552,In_4818);
and U115 (N_115,In_2633,In_2928);
nand U116 (N_116,In_1365,In_4468);
xor U117 (N_117,In_1057,In_3690);
and U118 (N_118,In_4719,In_4770);
and U119 (N_119,In_3131,In_4070);
nand U120 (N_120,In_3710,In_2995);
and U121 (N_121,In_43,In_1477);
and U122 (N_122,In_4386,In_3347);
xnor U123 (N_123,In_2456,In_1516);
nand U124 (N_124,In_3640,In_2260);
nor U125 (N_125,In_4959,In_1678);
nor U126 (N_126,In_3128,In_453);
and U127 (N_127,In_2497,In_1060);
or U128 (N_128,In_4406,In_1911);
or U129 (N_129,In_1107,In_4126);
and U130 (N_130,In_755,In_998);
nand U131 (N_131,In_4760,In_402);
nor U132 (N_132,In_4969,In_1498);
nor U133 (N_133,In_1560,In_734);
or U134 (N_134,In_3334,In_2723);
and U135 (N_135,In_4254,In_3549);
or U136 (N_136,In_621,In_4602);
or U137 (N_137,In_3221,In_4922);
xnor U138 (N_138,In_450,In_292);
nand U139 (N_139,In_469,In_354);
xnor U140 (N_140,In_978,In_4784);
xnor U141 (N_141,In_4416,In_3553);
and U142 (N_142,In_997,In_2823);
xnor U143 (N_143,In_1416,In_652);
or U144 (N_144,In_1576,In_2202);
nand U145 (N_145,In_3313,In_497);
nand U146 (N_146,In_2176,In_4255);
or U147 (N_147,In_1328,In_3365);
nor U148 (N_148,In_3962,In_724);
nand U149 (N_149,In_2205,In_2843);
nand U150 (N_150,In_4878,In_1544);
xor U151 (N_151,In_2010,In_3296);
nor U152 (N_152,In_69,In_869);
nand U153 (N_153,In_4278,In_278);
and U154 (N_154,In_1118,In_1426);
xor U155 (N_155,In_1605,In_4608);
nand U156 (N_156,In_1231,In_4049);
xor U157 (N_157,In_1294,In_4400);
or U158 (N_158,In_3915,In_3525);
or U159 (N_159,In_650,In_2460);
and U160 (N_160,In_767,In_2362);
and U161 (N_161,In_206,In_533);
or U162 (N_162,In_617,In_2032);
nor U163 (N_163,In_921,In_783);
nor U164 (N_164,In_1396,In_2236);
xor U165 (N_165,In_2183,In_3423);
or U166 (N_166,In_889,In_4164);
and U167 (N_167,In_4607,In_3956);
nand U168 (N_168,In_313,In_4415);
xnor U169 (N_169,In_282,In_2774);
nor U170 (N_170,In_4167,In_488);
nor U171 (N_171,In_4735,In_630);
nand U172 (N_172,In_2025,In_4862);
nand U173 (N_173,In_19,In_2945);
nand U174 (N_174,In_3275,In_141);
nor U175 (N_175,In_713,In_841);
nor U176 (N_176,In_4674,In_3586);
or U177 (N_177,In_993,In_4020);
or U178 (N_178,In_4554,In_4239);
and U179 (N_179,In_2444,In_3581);
xnor U180 (N_180,In_3240,In_3921);
nor U181 (N_181,In_2534,In_644);
xor U182 (N_182,In_1829,In_2653);
xnor U183 (N_183,In_1411,In_4767);
xnor U184 (N_184,In_4551,In_204);
or U185 (N_185,In_3612,In_4687);
xor U186 (N_186,In_16,In_1189);
nor U187 (N_187,In_4797,In_105);
nand U188 (N_188,In_4713,In_1526);
or U189 (N_189,In_3108,In_688);
or U190 (N_190,In_3961,In_4355);
xnor U191 (N_191,In_3247,In_3720);
xor U192 (N_192,In_4162,In_3940);
nor U193 (N_193,In_4982,In_1114);
or U194 (N_194,In_4302,In_559);
nor U195 (N_195,In_2834,In_385);
nand U196 (N_196,In_2419,In_2873);
and U197 (N_197,In_1128,In_1451);
nor U198 (N_198,In_4156,In_34);
and U199 (N_199,In_2191,In_4348);
nor U200 (N_200,In_3367,In_3609);
nand U201 (N_201,In_2824,In_711);
nor U202 (N_202,In_2639,In_4138);
and U203 (N_203,In_3933,In_4773);
and U204 (N_204,In_2898,In_1138);
nand U205 (N_205,In_2599,In_3162);
nor U206 (N_206,In_4710,In_326);
xnor U207 (N_207,In_4353,In_980);
xnor U208 (N_208,In_890,In_981);
or U209 (N_209,In_4361,In_3481);
xor U210 (N_210,In_794,In_2859);
and U211 (N_211,In_1400,In_866);
nand U212 (N_212,In_4160,In_4108);
or U213 (N_213,In_3526,In_2286);
and U214 (N_214,In_4616,In_1219);
and U215 (N_215,In_2273,In_4413);
nand U216 (N_216,In_2073,In_948);
xnor U217 (N_217,In_1836,In_3756);
and U218 (N_218,In_1570,In_632);
xor U219 (N_219,In_4084,In_4599);
and U220 (N_220,In_1322,In_1239);
nor U221 (N_221,In_761,In_303);
nor U222 (N_222,In_4526,In_3976);
nand U223 (N_223,In_3882,In_4171);
or U224 (N_224,In_641,In_1992);
or U225 (N_225,In_2595,In_1140);
nand U226 (N_226,In_506,In_4005);
xor U227 (N_227,In_1547,In_3178);
nand U228 (N_228,In_4716,In_1369);
nand U229 (N_229,In_75,In_1756);
nand U230 (N_230,In_3519,In_3105);
nand U231 (N_231,In_120,In_1700);
and U232 (N_232,In_2777,In_2933);
xnor U233 (N_233,In_4354,In_716);
nor U234 (N_234,In_918,In_2131);
or U235 (N_235,In_3918,In_4204);
and U236 (N_236,In_3250,In_3501);
and U237 (N_237,In_1275,In_2203);
nor U238 (N_238,In_4566,In_1677);
xor U239 (N_239,In_2416,In_1345);
xnor U240 (N_240,In_2495,In_4407);
xnor U241 (N_241,In_3706,In_912);
nor U242 (N_242,In_4728,In_1865);
xnor U243 (N_243,In_458,In_4657);
nor U244 (N_244,In_41,In_2681);
xor U245 (N_245,In_3657,In_4494);
nand U246 (N_246,In_1619,In_4304);
nor U247 (N_247,In_4264,In_4341);
or U248 (N_248,In_1931,In_1352);
and U249 (N_249,In_1309,In_2907);
xor U250 (N_250,In_315,In_3021);
nor U251 (N_251,In_2526,In_3763);
nor U252 (N_252,In_2544,In_2757);
or U253 (N_253,In_557,In_788);
nand U254 (N_254,In_1845,In_2324);
xnor U255 (N_255,In_4115,In_2151);
and U256 (N_256,In_4845,In_4805);
or U257 (N_257,In_4135,In_1305);
and U258 (N_258,In_1981,In_2130);
and U259 (N_259,In_1683,In_3822);
or U260 (N_260,In_4246,In_1609);
xor U261 (N_261,In_319,In_4478);
nand U262 (N_262,In_3222,In_3545);
or U263 (N_263,In_887,In_3911);
and U264 (N_264,In_4638,In_2059);
nor U265 (N_265,In_3794,In_2714);
and U266 (N_266,In_3739,In_4751);
xor U267 (N_267,In_35,In_476);
and U268 (N_268,In_2562,In_1510);
nand U269 (N_269,In_4768,In_1826);
nor U270 (N_270,In_2300,In_1495);
nor U271 (N_271,In_1887,In_2138);
or U272 (N_272,In_1221,In_1991);
xor U273 (N_273,In_3576,In_2354);
nand U274 (N_274,In_4842,In_2910);
nor U275 (N_275,In_2106,In_4944);
xnor U276 (N_276,In_3186,In_4124);
nor U277 (N_277,In_4427,In_2606);
nand U278 (N_278,In_1508,In_994);
and U279 (N_279,In_1146,In_3209);
nor U280 (N_280,In_2481,In_959);
and U281 (N_281,In_2790,In_2249);
xor U282 (N_282,In_3227,In_3206);
nor U283 (N_283,In_2048,In_4455);
and U284 (N_284,In_1183,In_4507);
or U285 (N_285,In_1787,In_627);
and U286 (N_286,In_448,In_2594);
or U287 (N_287,In_3554,In_2543);
xnor U288 (N_288,In_4462,In_3727);
nand U289 (N_289,In_3183,In_1951);
and U290 (N_290,In_1843,In_3799);
or U291 (N_291,In_2222,In_3414);
xor U292 (N_292,In_3042,In_2540);
or U293 (N_293,In_2689,In_1789);
or U294 (N_294,In_2529,In_4884);
or U295 (N_295,In_3895,In_4463);
and U296 (N_296,In_1979,In_862);
nand U297 (N_297,In_2221,In_771);
and U298 (N_298,In_4233,In_536);
and U299 (N_299,In_2,In_2208);
and U300 (N_300,In_570,In_3622);
xnor U301 (N_301,In_1078,In_4756);
nand U302 (N_302,In_1846,In_1831);
xor U303 (N_303,In_1001,In_4652);
or U304 (N_304,In_4109,In_1792);
or U305 (N_305,In_4506,In_2923);
nand U306 (N_306,In_2539,In_3465);
nand U307 (N_307,In_4803,In_3145);
xnor U308 (N_308,In_2507,In_2825);
xor U309 (N_309,In_4496,In_2631);
or U310 (N_310,In_1390,In_1714);
and U311 (N_311,In_2403,In_23);
xor U312 (N_312,In_917,In_3666);
or U313 (N_313,In_4612,In_3480);
nand U314 (N_314,In_4972,In_3003);
and U315 (N_315,In_2244,In_2601);
xnor U316 (N_316,In_343,In_813);
xnor U317 (N_317,In_2772,In_3842);
and U318 (N_318,In_2967,In_2782);
nor U319 (N_319,In_65,In_272);
and U320 (N_320,In_2281,In_1359);
xnor U321 (N_321,In_3122,In_4667);
and U322 (N_322,In_1050,In_1423);
nor U323 (N_323,In_4159,In_188);
and U324 (N_324,In_773,In_2007);
or U325 (N_325,In_1254,In_432);
nand U326 (N_326,In_2493,In_323);
xnor U327 (N_327,In_4572,In_3033);
xor U328 (N_328,In_1632,In_522);
or U329 (N_329,In_759,In_1850);
nor U330 (N_330,In_4880,In_4338);
or U331 (N_331,In_4130,In_2345);
xnor U332 (N_332,In_3328,In_3969);
nor U333 (N_333,In_3332,In_2869);
nand U334 (N_334,In_940,In_3451);
nand U335 (N_335,In_3502,In_676);
or U336 (N_336,In_3047,In_4517);
nor U337 (N_337,In_4078,In_4236);
or U338 (N_338,In_3823,In_992);
and U339 (N_339,In_853,In_4270);
and U340 (N_340,In_1671,In_4337);
and U341 (N_341,In_1172,In_4305);
nand U342 (N_342,In_4465,In_733);
and U343 (N_343,In_4700,In_3172);
or U344 (N_344,In_646,In_2490);
nor U345 (N_345,In_578,In_1367);
or U346 (N_346,In_1580,In_3161);
nor U347 (N_347,In_612,In_159);
xor U348 (N_348,In_3179,In_2876);
nor U349 (N_349,In_4769,In_990);
or U350 (N_350,In_3056,In_705);
xnor U351 (N_351,In_4792,In_461);
or U352 (N_352,In_4692,In_3635);
xnor U353 (N_353,In_1776,In_3664);
or U354 (N_354,In_49,In_4214);
xor U355 (N_355,In_1675,In_1893);
and U356 (N_356,In_433,In_1956);
or U357 (N_357,In_3417,In_1950);
or U358 (N_358,In_1241,In_2820);
xor U359 (N_359,In_3401,In_1966);
and U360 (N_360,In_2813,In_674);
xor U361 (N_361,In_3231,In_1766);
and U362 (N_362,In_3620,In_4013);
nor U363 (N_363,In_1317,In_1729);
xnor U364 (N_364,In_2242,In_389);
nand U365 (N_365,In_2499,In_1105);
or U366 (N_366,In_4177,In_1666);
nand U367 (N_367,In_1651,In_735);
nand U368 (N_368,In_2101,In_4613);
or U369 (N_369,In_1561,In_4539);
or U370 (N_370,In_3454,In_4336);
and U371 (N_371,In_423,In_4402);
or U372 (N_372,In_454,In_1825);
nand U373 (N_373,In_3389,In_2178);
and U374 (N_374,In_407,In_134);
or U375 (N_375,In_342,In_1937);
and U376 (N_376,In_3039,In_4707);
nor U377 (N_377,In_254,In_2323);
nor U378 (N_378,In_1397,In_4048);
nand U379 (N_379,In_3374,In_1066);
xor U380 (N_380,In_4826,In_4442);
xnor U381 (N_381,In_3448,In_3134);
and U382 (N_382,In_2798,In_2441);
nand U383 (N_383,In_834,In_4588);
and U384 (N_384,In_210,In_833);
or U385 (N_385,In_4584,In_4870);
xnor U386 (N_386,In_1456,In_4887);
nand U387 (N_387,In_4394,In_1233);
or U388 (N_388,In_2246,In_1100);
nand U389 (N_389,In_1569,In_2949);
xor U390 (N_390,In_2683,In_173);
nor U391 (N_391,In_723,In_1163);
nand U392 (N_392,In_117,In_3770);
xor U393 (N_393,In_2089,In_1627);
and U394 (N_394,In_1412,In_1301);
and U395 (N_395,In_4180,In_3653);
nand U396 (N_396,In_2768,In_440);
xnor U397 (N_397,In_2062,In_1444);
or U398 (N_398,In_1747,In_808);
nor U399 (N_399,In_2198,In_1143);
nand U400 (N_400,In_1351,In_2127);
or U401 (N_401,In_4795,In_3017);
nand U402 (N_402,In_968,In_939);
nor U403 (N_403,In_979,In_2730);
nor U404 (N_404,In_2915,In_2278);
xnor U405 (N_405,In_2346,In_2450);
nand U406 (N_406,In_1144,In_4957);
xnor U407 (N_407,In_987,In_2318);
nand U408 (N_408,In_371,In_1448);
or U409 (N_409,In_4099,In_1974);
and U410 (N_410,In_3588,In_2144);
nor U411 (N_411,In_2567,In_1798);
xnor U412 (N_412,In_4489,In_2214);
or U413 (N_413,In_4663,In_1554);
xor U414 (N_414,In_1119,In_4450);
and U415 (N_415,In_4547,In_302);
and U416 (N_416,In_3251,In_2268);
nand U417 (N_417,In_4064,In_4891);
xor U418 (N_418,In_4971,In_2672);
and U419 (N_419,In_2015,In_677);
nor U420 (N_420,In_1654,In_1549);
nor U421 (N_421,In_2100,In_4798);
xnor U422 (N_422,In_2721,In_2114);
or U423 (N_423,In_1475,In_4476);
nand U424 (N_424,In_1834,In_1377);
and U425 (N_425,In_1030,In_743);
xnor U426 (N_426,In_2245,In_2951);
or U427 (N_427,In_1088,In_4623);
xnor U428 (N_428,In_2868,In_2412);
and U429 (N_429,In_263,In_2454);
and U430 (N_430,In_1381,In_3254);
nor U431 (N_431,In_2167,In_765);
or U432 (N_432,In_20,In_1122);
and U433 (N_433,In_931,In_2522);
nand U434 (N_434,In_4231,In_2250);
and U435 (N_435,In_452,In_2057);
xnor U436 (N_436,In_3440,In_3210);
and U437 (N_437,In_3307,In_256);
xnor U438 (N_438,In_4347,In_2337);
xnor U439 (N_439,In_101,In_3955);
nor U440 (N_440,In_851,In_4913);
and U441 (N_441,In_3865,In_1469);
or U442 (N_442,In_3686,In_1511);
or U443 (N_443,In_3602,In_3436);
and U444 (N_444,In_2406,In_2916);
nor U445 (N_445,In_3632,In_3817);
or U446 (N_446,In_1197,In_1212);
xnor U447 (N_447,In_4038,In_1206);
nand U448 (N_448,In_4412,In_242);
xnor U449 (N_449,In_1773,In_3875);
nor U450 (N_450,In_886,In_3267);
and U451 (N_451,In_338,In_509);
xnor U452 (N_452,In_4002,In_2760);
or U453 (N_453,In_171,In_523);
nand U454 (N_454,In_3990,In_915);
nand U455 (N_455,In_160,In_3833);
nor U456 (N_456,In_1909,In_3740);
and U457 (N_457,In_2931,In_1967);
xnor U458 (N_458,In_4640,In_3778);
nor U459 (N_459,In_4024,In_347);
and U460 (N_460,In_1658,In_1315);
nand U461 (N_461,In_2299,In_2033);
or U462 (N_462,In_3319,In_3894);
nor U463 (N_463,In_3182,In_3618);
nor U464 (N_464,In_538,In_4989);
nor U465 (N_465,In_2909,In_792);
nor U466 (N_466,In_3928,In_2733);
nand U467 (N_467,In_905,In_4704);
or U468 (N_468,In_4154,In_217);
nand U469 (N_469,In_1620,In_700);
and U470 (N_470,In_1919,In_1917);
nand U471 (N_471,In_2758,In_2778);
and U472 (N_472,In_1108,In_1249);
nand U473 (N_473,In_2603,In_4234);
and U474 (N_474,In_2806,In_659);
and U475 (N_475,In_1803,In_757);
or U476 (N_476,In_3353,In_2084);
or U477 (N_477,In_1923,In_468);
nor U478 (N_478,In_2475,In_1325);
or U479 (N_479,In_3351,In_3280);
or U480 (N_480,In_2867,In_304);
and U481 (N_481,In_2703,In_655);
or U482 (N_482,In_4820,In_4399);
xor U483 (N_483,In_769,In_265);
and U484 (N_484,In_1817,In_3107);
or U485 (N_485,In_2431,In_2027);
nor U486 (N_486,In_286,In_1856);
nand U487 (N_487,In_1970,In_4294);
nand U488 (N_488,In_2469,In_119);
nor U489 (N_489,In_4834,In_180);
or U490 (N_490,In_1430,In_4827);
nor U491 (N_491,In_3287,In_1501);
or U492 (N_492,In_4209,In_1154);
and U493 (N_493,In_2036,In_2750);
nor U494 (N_494,In_3747,In_4945);
nor U495 (N_495,In_1871,In_3821);
nand U496 (N_496,In_3949,In_4314);
and U497 (N_497,In_1320,In_1600);
xor U498 (N_498,In_4895,In_520);
and U499 (N_499,In_24,In_2808);
nand U500 (N_500,In_3117,In_3764);
nor U501 (N_501,In_2491,In_668);
nor U502 (N_502,In_1866,In_4954);
and U503 (N_503,N_361,In_1420);
or U504 (N_504,In_3390,In_3410);
and U505 (N_505,In_4740,N_486);
nand U506 (N_506,In_3780,In_191);
or U507 (N_507,In_2216,In_1614);
xor U508 (N_508,In_1425,In_3458);
nor U509 (N_509,In_2893,In_2776);
nand U510 (N_510,In_4853,In_1152);
nor U511 (N_511,N_492,In_1763);
nand U512 (N_512,In_4096,In_3286);
or U513 (N_513,In_1199,In_972);
and U514 (N_514,N_452,In_3812);
or U515 (N_515,In_3387,In_1897);
nand U516 (N_516,In_2516,In_2224);
xnor U517 (N_517,In_398,In_4921);
or U518 (N_518,In_4137,In_4097);
and U519 (N_519,In_517,In_3593);
nor U520 (N_520,N_394,In_1655);
or U521 (N_521,In_3036,In_3980);
and U522 (N_522,In_1159,In_2593);
nand U523 (N_523,In_2133,In_2125);
and U524 (N_524,In_665,In_3592);
nand U525 (N_525,In_3297,In_3293);
nor U526 (N_526,In_4565,In_906);
and U527 (N_527,In_3364,N_156);
or U528 (N_528,In_3026,In_3382);
nand U529 (N_529,In_2752,In_3246);
xnor U530 (N_530,In_1665,In_1914);
or U531 (N_531,In_687,In_3672);
xnor U532 (N_532,In_1797,In_3897);
or U533 (N_533,In_1335,In_4684);
xor U534 (N_534,In_4723,N_95);
xnor U535 (N_535,In_4793,In_1592);
or U536 (N_536,N_333,In_3627);
or U537 (N_537,In_1071,In_1104);
xor U538 (N_538,In_1059,In_1403);
xor U539 (N_539,In_2743,N_183);
nand U540 (N_540,In_1383,N_310);
or U541 (N_541,In_4825,In_4935);
nand U542 (N_542,In_3786,In_2029);
nand U543 (N_543,In_2122,In_2139);
nor U544 (N_544,N_65,In_929);
nor U545 (N_545,N_197,In_4936);
nor U546 (N_546,In_4576,In_4357);
and U547 (N_547,In_4747,In_1236);
xor U548 (N_548,In_54,In_810);
xor U549 (N_549,In_4470,In_1760);
nand U550 (N_550,In_1141,N_493);
and U551 (N_551,In_3652,In_1685);
nor U552 (N_552,In_2807,In_4283);
nor U553 (N_553,In_214,In_1821);
nor U554 (N_554,In_64,In_3085);
xor U555 (N_555,In_4017,In_871);
and U556 (N_556,In_1872,In_786);
or U557 (N_557,In_564,In_4074);
and U558 (N_558,In_1689,In_3896);
and U559 (N_559,In_964,In_4377);
and U560 (N_560,In_199,In_3159);
xor U561 (N_561,In_599,In_746);
xnor U562 (N_562,In_4435,In_2425);
nand U563 (N_563,In_4106,N_54);
and U564 (N_564,In_1842,In_1388);
xor U565 (N_565,In_3864,N_84);
and U566 (N_566,In_1321,In_74);
xnor U567 (N_567,In_4089,In_4525);
and U568 (N_568,In_4788,In_3826);
nand U569 (N_569,In_4371,In_3314);
xnor U570 (N_570,In_613,In_1173);
and U571 (N_571,N_114,In_4188);
or U572 (N_572,In_3067,In_2240);
xor U573 (N_573,In_684,In_4646);
and U574 (N_574,N_313,In_2314);
nand U575 (N_575,N_134,N_247);
nand U576 (N_576,In_619,In_2646);
nand U577 (N_577,In_568,In_3291);
nand U578 (N_578,In_4604,In_1830);
xor U579 (N_579,In_3080,In_366);
and U580 (N_580,In_3304,In_4032);
nor U581 (N_581,In_975,In_508);
and U582 (N_582,In_631,In_2241);
nand U583 (N_583,N_8,In_2005);
nand U584 (N_584,N_132,In_3646);
nor U585 (N_585,In_1470,In_4829);
or U586 (N_586,In_726,In_3762);
nand U587 (N_587,In_4102,In_424);
xnor U588 (N_588,In_1000,N_334);
xnor U589 (N_589,In_4310,N_281);
and U590 (N_590,In_2063,In_4317);
nor U591 (N_591,In_2537,N_145);
nor U592 (N_592,In_2579,In_3616);
or U593 (N_593,In_3531,In_3376);
or U594 (N_594,In_2879,In_1838);
and U595 (N_595,In_146,In_4141);
or U596 (N_596,N_437,In_447);
and U597 (N_597,In_4469,In_1704);
nand U598 (N_598,In_2767,In_4518);
nor U599 (N_599,In_4202,In_2982);
xnor U600 (N_600,In_4744,In_184);
and U601 (N_601,In_1521,In_2677);
or U602 (N_602,In_3359,In_3474);
and U603 (N_603,In_4648,In_403);
nand U604 (N_604,In_1777,In_828);
and U605 (N_605,In_3559,In_4147);
nor U606 (N_606,In_4093,In_3759);
or U607 (N_607,In_832,In_2675);
and U608 (N_608,In_4567,In_66);
nand U609 (N_609,N_424,In_3906);
nand U610 (N_610,In_4152,In_4852);
nand U611 (N_611,In_4281,In_3204);
or U612 (N_612,In_877,In_390);
nor U613 (N_613,N_320,In_44);
nand U614 (N_614,In_1978,In_4063);
xor U615 (N_615,In_3634,N_202);
nand U616 (N_616,In_643,N_60);
or U617 (N_617,In_3975,In_3851);
nand U618 (N_618,In_1527,In_3798);
nor U619 (N_619,In_3405,In_3560);
xnor U620 (N_620,In_1386,In_2940);
nand U621 (N_621,In_109,In_1042);
nand U622 (N_622,In_4656,In_1617);
nor U623 (N_623,In_361,In_4015);
and U624 (N_624,In_758,In_1537);
and U625 (N_625,In_1618,N_309);
or U626 (N_626,In_1701,In_2748);
or U627 (N_627,In_3877,In_3802);
nand U628 (N_628,In_693,N_421);
xor U629 (N_629,In_574,In_2816);
nor U630 (N_630,In_4929,In_3089);
nor U631 (N_631,In_2657,In_2612);
and U632 (N_632,In_2258,In_2981);
or U633 (N_633,In_3109,In_220);
and U634 (N_634,In_2996,In_708);
xnor U635 (N_635,In_3621,In_463);
xor U636 (N_636,In_123,In_2280);
nor U637 (N_637,In_2973,In_3841);
nor U638 (N_638,In_554,N_354);
and U639 (N_639,In_558,N_237);
or U640 (N_640,In_3805,In_2332);
or U641 (N_641,In_1092,In_4535);
nand U642 (N_642,In_4531,In_3148);
xor U643 (N_643,In_3965,In_4333);
nand U644 (N_644,In_2908,In_473);
nand U645 (N_645,N_126,In_3556);
and U646 (N_646,In_3708,In_4018);
and U647 (N_647,In_3370,In_3312);
nand U648 (N_648,In_1543,N_458);
xnor U649 (N_649,In_2699,N_75);
nand U650 (N_650,In_4908,In_1679);
and U651 (N_651,N_399,In_1348);
nand U652 (N_652,N_242,In_2553);
nand U653 (N_653,In_1243,In_3288);
nand U654 (N_654,N_77,In_2038);
or U655 (N_655,In_3104,In_2731);
or U656 (N_656,In_4387,In_3331);
xnor U657 (N_657,In_4358,In_4107);
nor U658 (N_658,In_3472,In_953);
nor U659 (N_659,In_3669,In_514);
or U660 (N_660,In_295,In_961);
and U661 (N_661,In_2991,In_924);
nor U662 (N_662,In_4490,In_1041);
or U663 (N_663,In_4651,In_2458);
and U664 (N_664,N_101,In_4023);
nor U665 (N_665,In_2079,In_3281);
xor U666 (N_666,In_4332,In_4695);
and U667 (N_667,In_334,In_2311);
xnor U668 (N_668,In_30,In_893);
and U669 (N_669,In_1907,In_2448);
or U670 (N_670,In_3278,In_2581);
nand U671 (N_671,In_4380,In_1375);
nor U672 (N_672,In_89,In_2900);
nand U673 (N_673,In_1182,In_2917);
nand U674 (N_674,In_1827,In_1156);
nor U675 (N_675,In_4085,N_178);
nor U676 (N_676,In_1045,N_187);
or U677 (N_677,N_208,In_246);
nor U678 (N_678,In_2795,In_3165);
or U679 (N_679,In_1790,N_124);
or U680 (N_680,In_3881,In_957);
nand U681 (N_681,In_4056,In_4157);
xor U682 (N_682,In_2296,In_3904);
xor U683 (N_683,In_1488,In_2740);
nor U684 (N_684,In_2473,In_4869);
and U685 (N_685,In_4438,In_39);
and U686 (N_686,In_1928,In_275);
nand U687 (N_687,In_3277,N_418);
nand U688 (N_688,In_1648,In_1036);
xnor U689 (N_689,In_3538,In_3573);
nand U690 (N_690,In_4585,In_2651);
and U691 (N_691,In_4091,In_475);
and U692 (N_692,In_4098,In_942);
nand U693 (N_693,In_2605,N_0);
xor U694 (N_694,In_445,In_2190);
xor U695 (N_695,In_1215,In_4393);
nand U696 (N_696,In_2693,N_28);
or U697 (N_697,In_2694,N_312);
or U698 (N_698,In_3518,N_56);
nand U699 (N_699,In_3876,In_547);
xnor U700 (N_700,In_2417,In_647);
and U701 (N_701,In_4743,In_3399);
or U702 (N_702,N_22,In_3091);
or U703 (N_703,In_1946,In_850);
nor U704 (N_704,In_2756,In_2863);
and U705 (N_705,N_63,In_4175);
and U706 (N_706,N_469,In_1246);
and U707 (N_707,In_3847,In_1170);
and U708 (N_708,In_831,In_1597);
xor U709 (N_709,In_3610,In_3350);
or U710 (N_710,In_82,In_4212);
xnor U711 (N_711,In_1064,In_1296);
nand U712 (N_712,In_3343,In_2521);
or U713 (N_713,In_3818,In_1194);
or U714 (N_714,In_1427,In_3546);
nand U715 (N_715,In_2189,In_1709);
or U716 (N_716,In_367,In_1720);
nand U717 (N_717,In_1568,In_1466);
nand U718 (N_718,In_1028,In_2301);
and U719 (N_719,In_1067,N_276);
nand U720 (N_720,N_284,In_3330);
or U721 (N_721,In_2835,N_467);
or U722 (N_722,In_310,In_3333);
nor U723 (N_723,In_1270,In_3946);
or U724 (N_724,In_2556,N_321);
nand U725 (N_725,In_4299,In_3595);
and U726 (N_726,In_2906,N_191);
nor U727 (N_727,In_569,In_4452);
nand U728 (N_728,In_2277,In_923);
and U729 (N_729,In_4830,In_4280);
nor U730 (N_730,In_2370,N_104);
and U731 (N_731,In_406,In_2897);
nand U732 (N_732,In_3217,In_2275);
nand U733 (N_733,N_31,In_4620);
or U734 (N_734,In_4191,In_1015);
xor U735 (N_735,In_4121,In_3728);
nor U736 (N_736,In_1265,In_2832);
or U737 (N_737,In_4542,In_48);
or U738 (N_738,In_207,In_2418);
nor U739 (N_739,In_4595,In_4155);
and U740 (N_740,In_3880,In_3643);
nor U741 (N_741,In_96,In_966);
nand U742 (N_742,In_1409,In_1884);
and U743 (N_743,N_441,In_1047);
xnor U744 (N_744,In_4315,In_2520);
or U745 (N_745,In_4850,In_1002);
xnor U746 (N_746,In_870,In_4069);
and U747 (N_747,In_1901,In_3208);
nor U748 (N_748,In_2252,In_1354);
nand U749 (N_749,In_3783,In_1875);
xor U750 (N_750,In_3773,In_3816);
and U751 (N_751,In_4082,In_2075);
nand U752 (N_752,In_2389,In_1358);
and U753 (N_753,In_147,In_678);
nand U754 (N_754,N_70,In_4323);
nor U755 (N_755,In_2561,In_4919);
nor U756 (N_756,In_4079,In_4247);
nor U757 (N_757,In_1482,In_3504);
xor U758 (N_758,In_76,In_3890);
nor U759 (N_759,In_954,In_2132);
or U760 (N_760,In_3582,N_302);
nor U761 (N_761,In_1288,In_1308);
nor U762 (N_762,N_78,In_2530);
and U763 (N_763,In_1935,N_393);
xnor U764 (N_764,N_263,In_4628);
and U765 (N_765,In_694,In_781);
nand U766 (N_766,N_476,In_3776);
nand U767 (N_767,In_4232,In_3052);
or U768 (N_768,In_1731,In_269);
nor U769 (N_769,In_1333,In_4654);
nand U770 (N_770,In_93,In_4007);
or U771 (N_771,In_301,In_3840);
xor U772 (N_772,In_2402,In_3930);
nor U773 (N_773,In_703,In_3378);
nor U774 (N_774,In_4516,In_2400);
xor U775 (N_775,In_227,In_439);
nor U776 (N_776,In_3478,In_639);
xor U777 (N_777,In_2614,In_809);
nor U778 (N_778,In_3827,In_1669);
nor U779 (N_779,In_4984,In_1407);
nand U780 (N_780,In_2366,In_3503);
and U781 (N_781,In_790,N_87);
nand U782 (N_782,In_2302,N_29);
and U783 (N_783,In_2145,In_142);
nand U784 (N_784,In_4257,In_1638);
xor U785 (N_785,In_4942,In_2165);
or U786 (N_786,In_2598,In_1429);
xor U787 (N_787,In_750,In_2211);
and U788 (N_788,In_4080,In_1244);
nor U789 (N_789,In_1589,N_294);
and U790 (N_790,In_2842,In_3985);
nand U791 (N_791,In_1784,In_3007);
xor U792 (N_792,In_1220,N_158);
xnor U793 (N_793,In_1101,N_420);
xor U794 (N_794,In_4001,In_4466);
and U795 (N_795,In_3945,In_2615);
nor U796 (N_796,In_1663,In_2035);
xnor U797 (N_797,In_2946,In_4440);
nand U798 (N_798,In_115,In_309);
xnor U799 (N_799,In_1222,In_2156);
nor U800 (N_800,N_379,In_799);
or U801 (N_801,In_1439,In_2026);
xor U802 (N_802,In_1818,In_1973);
and U803 (N_803,In_3771,In_11);
nor U804 (N_804,In_4072,In_401);
and U805 (N_805,In_2621,In_2173);
nand U806 (N_806,In_3513,In_573);
and U807 (N_807,In_4749,In_4375);
xnor U808 (N_808,In_2472,In_1268);
xor U809 (N_809,In_3997,In_560);
nor U810 (N_810,In_2116,N_224);
or U811 (N_811,In_255,In_3216);
nand U812 (N_812,In_3547,In_1953);
nand U813 (N_813,In_756,N_274);
and U814 (N_814,In_1932,In_4308);
or U815 (N_815,In_3355,In_1298);
nor U816 (N_816,In_3397,In_782);
nor U817 (N_817,In_4817,In_2328);
or U818 (N_818,In_1755,N_305);
nand U819 (N_819,N_154,In_4448);
and U820 (N_820,N_336,In_4181);
nand U821 (N_821,N_218,In_1769);
and U822 (N_822,In_166,In_2749);
and U823 (N_823,In_1595,In_1196);
nor U824 (N_824,In_4066,In_3059);
and U825 (N_825,In_1505,In_1939);
and U826 (N_826,In_3101,In_1535);
or U827 (N_827,In_2295,In_1955);
or U828 (N_828,In_3373,In_4801);
and U829 (N_829,In_94,In_4993);
nor U830 (N_830,In_4813,N_91);
xnor U831 (N_831,In_1035,In_150);
and U832 (N_832,In_1076,In_1876);
nand U833 (N_833,N_71,In_3599);
nand U834 (N_834,In_4814,In_2891);
nor U835 (N_835,In_2021,In_3927);
or U836 (N_836,In_1380,N_26);
nand U837 (N_837,In_967,In_4927);
xor U838 (N_838,In_2578,In_4746);
xnor U839 (N_839,In_154,In_4621);
or U840 (N_840,In_3006,In_634);
and U841 (N_841,In_2588,In_2179);
nand U842 (N_842,N_248,In_4883);
or U843 (N_843,In_731,In_4176);
xor U844 (N_844,In_4859,In_1151);
nand U845 (N_845,In_3995,In_3742);
nand U846 (N_846,In_59,In_2685);
and U847 (N_847,In_800,In_399);
xnor U848 (N_848,In_4764,N_227);
or U849 (N_849,In_3071,In_308);
or U850 (N_850,In_3983,N_174);
or U851 (N_851,In_1113,In_299);
nor U852 (N_852,In_1734,In_2398);
xor U853 (N_853,In_2060,In_1849);
xnor U854 (N_854,In_3860,In_3068);
xor U855 (N_855,In_4580,In_4391);
nor U856 (N_856,In_3699,In_37);
nor U857 (N_857,In_4414,In_904);
and U858 (N_858,N_352,In_2947);
and U859 (N_859,In_3259,In_2420);
xnor U860 (N_860,In_2932,In_4025);
xnor U861 (N_861,In_4051,In_914);
xor U862 (N_862,In_4660,In_4335);
or U863 (N_863,In_1491,In_4515);
nor U864 (N_864,In_2596,In_648);
xor U865 (N_865,In_3279,In_2564);
and U866 (N_866,In_2987,In_4389);
or U867 (N_867,In_1455,N_246);
and U868 (N_868,In_4519,In_3023);
nand U869 (N_869,In_2408,In_1558);
nor U870 (N_870,In_4318,In_1761);
nand U871 (N_871,In_3993,In_3611);
or U872 (N_872,In_1711,In_4824);
or U873 (N_873,In_1473,In_3066);
or U874 (N_874,In_3292,In_4187);
or U875 (N_875,In_2736,In_3722);
and U876 (N_876,In_4058,In_2968);
xnor U877 (N_877,In_2052,In_2972);
and U878 (N_878,In_4708,In_1707);
nor U879 (N_879,In_3982,In_2629);
xor U880 (N_880,In_1494,In_4968);
nand U881 (N_881,In_3413,N_364);
and U882 (N_882,In_2797,In_3781);
and U883 (N_883,In_4504,In_2435);
nand U884 (N_884,In_4799,In_854);
xnor U885 (N_885,N_259,In_1809);
nor U886 (N_886,In_1264,In_1942);
and U887 (N_887,In_1290,In_4832);
xor U888 (N_888,In_1251,In_4815);
or U889 (N_889,In_2313,In_237);
xnor U890 (N_890,In_1868,N_359);
xnor U891 (N_891,In_3072,In_4867);
nand U892 (N_892,In_2927,In_4150);
or U893 (N_893,In_4559,In_314);
and U894 (N_894,In_4594,In_2197);
nand U895 (N_895,In_3038,N_353);
nor U896 (N_896,In_512,In_2812);
or U897 (N_897,In_1770,In_1441);
and U898 (N_898,In_1116,In_4360);
nor U899 (N_899,In_1748,In_4409);
nand U900 (N_900,In_2957,In_3958);
or U901 (N_901,In_4166,In_2283);
nand U902 (N_902,N_323,In_2502);
and U903 (N_903,In_4388,In_3226);
or U904 (N_904,In_2168,In_1474);
xnor U905 (N_905,N_59,In_4596);
and U906 (N_906,N_157,In_1022);
and U907 (N_907,In_986,In_2674);
nor U908 (N_908,In_4201,In_1598);
nand U909 (N_909,In_3568,In_4433);
and U910 (N_910,In_2804,In_1631);
nor U911 (N_911,In_1664,In_4351);
nand U912 (N_912,In_4865,In_2708);
or U913 (N_913,In_565,In_2838);
nand U914 (N_914,In_2525,N_434);
nor U915 (N_915,In_3908,In_4758);
xnor U916 (N_916,In_2912,In_4843);
xor U917 (N_917,In_1179,In_2506);
nand U918 (N_918,In_2620,N_413);
and U919 (N_919,In_3425,N_299);
nand U920 (N_920,In_4037,In_4949);
or U921 (N_921,In_827,In_3570);
and U922 (N_922,In_2886,In_1459);
nand U923 (N_923,In_3486,In_1702);
nand U924 (N_924,In_927,In_4511);
nand U925 (N_925,In_804,In_1224);
or U926 (N_926,In_216,In_1879);
and U927 (N_927,In_3988,In_1739);
xnor U928 (N_928,In_797,In_2976);
nand U929 (N_929,In_4851,In_2872);
xor U930 (N_930,In_1010,In_486);
or U931 (N_931,In_2524,N_325);
nor U932 (N_932,In_2340,In_2377);
nor U933 (N_933,In_3153,In_946);
nand U934 (N_934,In_484,N_288);
nor U935 (N_935,In_2881,In_4404);
nor U936 (N_936,In_2583,In_279);
nand U937 (N_937,In_3160,N_24);
xnor U938 (N_938,In_2517,In_2006);
nand U939 (N_939,In_3484,In_3707);
nand U940 (N_940,In_4706,In_2943);
nor U941 (N_941,In_2914,In_1480);
and U942 (N_942,In_2892,In_3412);
and U943 (N_943,In_1216,In_2597);
or U944 (N_944,In_4653,In_1771);
nand U945 (N_945,In_2926,N_220);
or U946 (N_946,In_4571,In_3076);
nand U947 (N_947,N_74,N_88);
or U948 (N_948,In_4249,In_727);
nor U949 (N_949,In_3083,In_4185);
nor U950 (N_950,In_3814,In_686);
or U951 (N_951,In_2766,In_3155);
or U952 (N_952,In_4131,In_594);
and U953 (N_953,N_184,In_4671);
and U954 (N_954,In_3127,In_2954);
nor U955 (N_955,In_4505,In_1339);
xor U956 (N_956,In_3429,In_1848);
nand U957 (N_957,In_98,In_196);
and U958 (N_958,In_4275,In_3073);
and U959 (N_959,In_911,N_159);
or U960 (N_960,In_2285,In_1622);
nor U961 (N_961,In_633,In_3380);
or U962 (N_962,In_1612,In_610);
and U963 (N_963,In_208,In_2140);
nor U964 (N_964,In_1074,In_3935);
xor U965 (N_965,In_4312,In_2904);
and U966 (N_966,In_4044,In_394);
nand U967 (N_967,In_930,In_3232);
nand U968 (N_968,In_4248,In_1744);
nor U969 (N_969,In_2338,In_2462);
nand U970 (N_970,In_3614,In_702);
and U971 (N_971,In_3163,In_1719);
xnor U972 (N_972,In_4235,In_1517);
and U973 (N_973,In_1272,In_3613);
nor U974 (N_974,In_878,In_480);
or U975 (N_975,In_58,In_4772);
and U976 (N_976,In_1257,In_3852);
and U977 (N_977,In_4190,N_327);
nor U978 (N_978,In_2531,N_222);
or U979 (N_979,In_365,N_447);
xnor U980 (N_980,In_2072,In_1413);
nor U981 (N_981,In_798,In_2064);
and U982 (N_982,In_4587,In_4664);
and U983 (N_983,In_4408,In_3651);
nor U984 (N_984,N_103,In_858);
xnor U985 (N_985,In_845,N_135);
and U986 (N_986,In_4178,In_2702);
and U987 (N_987,In_3637,In_2960);
xor U988 (N_988,In_1185,In_4144);
xnor U989 (N_989,In_4174,In_487);
xnor U990 (N_990,In_4846,In_4685);
nor U991 (N_991,In_3726,In_3536);
and U992 (N_992,N_366,In_2883);
and U993 (N_993,In_3255,In_1645);
nor U994 (N_994,In_321,In_3663);
nand U995 (N_995,In_985,In_1393);
nand U996 (N_996,In_2438,In_1518);
xor U997 (N_997,In_4894,N_76);
or U998 (N_998,N_72,N_387);
nand U999 (N_999,In_377,In_1765);
nor U1000 (N_1000,In_4888,In_2801);
xnor U1001 (N_1001,N_507,N_602);
xor U1002 (N_1002,In_2575,In_3393);
and U1003 (N_1003,In_943,In_1691);
nor U1004 (N_1004,In_4298,In_2992);
and U1005 (N_1005,In_135,In_418);
and U1006 (N_1006,N_279,In_283);
xor U1007 (N_1007,In_3658,N_572);
or U1008 (N_1008,In_2107,In_3564);
nor U1009 (N_1009,In_1512,In_3150);
xnor U1010 (N_1010,In_4714,In_2002);
or U1011 (N_1011,In_649,In_4434);
and U1012 (N_1012,In_4771,In_3442);
xnor U1013 (N_1013,In_235,In_1009);
and U1014 (N_1014,In_609,N_565);
nand U1015 (N_1015,In_3719,In_3205);
xnor U1016 (N_1016,In_2169,N_35);
and U1017 (N_1017,In_1063,In_3467);
or U1018 (N_1018,In_3419,N_482);
or U1019 (N_1019,In_2853,In_1261);
or U1020 (N_1020,In_1718,In_4964);
nor U1021 (N_1021,N_825,In_1874);
and U1022 (N_1022,N_123,N_376);
xor U1023 (N_1023,In_2161,N_658);
or U1024 (N_1024,In_546,In_3269);
nor U1025 (N_1025,In_2984,In_926);
or U1026 (N_1026,In_2963,In_3724);
and U1027 (N_1027,In_78,In_297);
xnor U1028 (N_1028,N_317,In_894);
nor U1029 (N_1029,N_589,N_289);
or U1030 (N_1030,In_863,In_2093);
or U1031 (N_1031,In_4256,N_335);
and U1032 (N_1032,In_45,In_4483);
nor U1033 (N_1033,In_2918,In_580);
nand U1034 (N_1034,In_1642,In_1661);
nand U1035 (N_1035,N_386,In_1634);
nor U1036 (N_1036,In_3914,N_721);
and U1037 (N_1037,In_1479,N_932);
nor U1038 (N_1038,N_580,In_3506);
or U1039 (N_1039,In_4334,N_109);
xor U1040 (N_1040,In_1331,In_4384);
xor U1041 (N_1041,In_3697,In_4782);
or U1042 (N_1042,In_1896,In_222);
nand U1043 (N_1043,In_4570,N_908);
nor U1044 (N_1044,N_793,In_3093);
or U1045 (N_1045,In_984,In_2925);
nor U1046 (N_1046,In_1235,In_380);
or U1047 (N_1047,N_596,In_4454);
nor U1048 (N_1048,In_51,In_884);
and U1049 (N_1049,In_4947,In_1903);
nor U1050 (N_1050,In_811,In_2310);
or U1051 (N_1051,In_2509,In_1852);
and U1052 (N_1052,In_3952,In_2298);
nor U1053 (N_1053,In_1086,In_2793);
nor U1054 (N_1054,In_2652,In_3530);
or U1055 (N_1055,N_553,In_3942);
or U1056 (N_1056,N_117,N_375);
nor U1057 (N_1057,In_4876,In_1061);
nand U1058 (N_1058,In_4577,In_2428);
xnor U1059 (N_1059,In_1214,In_3681);
or U1060 (N_1060,In_2663,In_2054);
nor U1061 (N_1061,In_2542,In_3970);
or U1062 (N_1062,In_1457,In_2827);
nand U1063 (N_1063,In_1485,N_951);
xor U1064 (N_1064,In_46,In_3305);
nand U1065 (N_1065,In_2153,In_2985);
xor U1066 (N_1066,In_1075,In_1371);
xnor U1067 (N_1067,In_1252,In_3300);
nor U1068 (N_1068,In_1730,In_434);
or U1069 (N_1069,In_3803,In_3828);
or U1070 (N_1070,In_3339,In_4675);
nand U1071 (N_1071,In_2157,In_233);
xor U1072 (N_1072,In_1795,In_244);
nand U1073 (N_1073,In_3242,In_239);
or U1074 (N_1074,In_2361,N_976);
xnor U1075 (N_1075,In_1330,N_570);
nor U1076 (N_1076,In_3696,In_784);
and U1077 (N_1077,In_3459,In_2878);
xnor U1078 (N_1078,In_2443,In_1436);
xor U1079 (N_1079,In_2289,In_4366);
or U1080 (N_1080,In_4218,N_346);
xnor U1081 (N_1081,In_1548,In_4457);
nand U1082 (N_1082,N_755,In_1124);
xnor U1083 (N_1083,In_4701,In_1079);
xnor U1084 (N_1084,In_121,In_280);
and U1085 (N_1085,In_1453,In_2109);
nor U1086 (N_1086,In_3001,In_2174);
and U1087 (N_1087,In_33,In_264);
xor U1088 (N_1088,In_1142,In_638);
and U1089 (N_1089,N_945,In_2574);
or U1090 (N_1090,In_3605,N_552);
xnor U1091 (N_1091,In_748,In_2053);
xnor U1092 (N_1092,In_1794,In_260);
and U1093 (N_1093,In_3360,In_2640);
and U1094 (N_1094,In_1326,N_678);
xor U1095 (N_1095,In_3948,In_4429);
or U1096 (N_1096,In_3926,N_769);
xnor U1097 (N_1097,In_2171,N_133);
nand U1098 (N_1098,In_2937,In_3811);
nand U1099 (N_1099,In_2030,In_2679);
and U1100 (N_1100,In_4263,In_3885);
nand U1101 (N_1101,N_556,N_702);
nor U1102 (N_1102,In_268,N_495);
nand U1103 (N_1103,N_498,In_2635);
and U1104 (N_1104,In_3257,In_2572);
nand U1105 (N_1105,In_4903,In_1814);
xnor U1106 (N_1106,In_4681,In_4683);
nand U1107 (N_1107,In_1989,In_412);
or U1108 (N_1108,N_894,In_1394);
xnor U1109 (N_1109,N_213,In_2636);
and U1110 (N_1110,N_752,In_3607);
xnor U1111 (N_1111,N_261,In_3853);
xor U1112 (N_1112,In_3121,In_3363);
or U1113 (N_1113,In_3916,In_4113);
xor U1114 (N_1114,N_371,In_507);
nor U1115 (N_1115,In_1277,In_4609);
nor U1116 (N_1116,In_2780,In_3510);
and U1117 (N_1117,In_3934,N_228);
xnor U1118 (N_1118,N_669,In_3244);
xnor U1119 (N_1119,In_3989,In_4035);
xor U1120 (N_1120,In_2392,In_1768);
and U1121 (N_1121,N_245,In_1811);
and U1122 (N_1122,In_4579,In_2188);
nand U1123 (N_1123,N_508,In_3539);
or U1124 (N_1124,In_1542,In_3352);
nor U1125 (N_1125,In_4296,In_1556);
xnor U1126 (N_1126,N_646,In_1262);
and U1127 (N_1127,In_4858,In_3290);
xor U1128 (N_1128,In_1353,In_382);
or U1129 (N_1129,In_4027,In_3034);
xnor U1130 (N_1130,In_3452,In_2217);
and U1131 (N_1131,In_2558,N_645);
nand U1132 (N_1132,In_4437,In_815);
xor U1133 (N_1133,In_1997,In_3103);
xor U1134 (N_1134,In_4514,N_445);
or U1135 (N_1135,In_3402,In_970);
and U1136 (N_1136,N_582,N_782);
and U1137 (N_1137,In_2123,In_2083);
or U1138 (N_1138,N_953,N_931);
nand U1139 (N_1139,In_3943,In_582);
and U1140 (N_1140,In_328,In_1936);
nor U1141 (N_1141,In_3655,In_608);
nand U1142 (N_1142,N_277,In_3069);
and U1143 (N_1143,In_1998,In_1984);
and U1144 (N_1144,In_3263,In_2150);
and U1145 (N_1145,N_874,In_3149);
nand U1146 (N_1146,In_1332,N_980);
nor U1147 (N_1147,N_637,N_758);
or U1148 (N_1148,In_673,In_742);
nor U1149 (N_1149,In_194,In_3061);
xor U1150 (N_1150,In_2474,In_2858);
or U1151 (N_1151,In_1193,In_4882);
xor U1152 (N_1152,In_4385,In_1583);
nand U1153 (N_1153,In_2624,In_3215);
and U1154 (N_1154,N_69,In_1740);
nor U1155 (N_1155,N_865,In_597);
nand U1156 (N_1156,In_4836,In_4211);
and U1157 (N_1157,In_1808,In_4193);
or U1158 (N_1158,N_648,In_2355);
or U1159 (N_1159,N_107,In_935);
nand U1160 (N_1160,In_491,In_2378);
or U1161 (N_1161,N_783,In_4673);
xor U1162 (N_1162,In_2476,In_4914);
and U1163 (N_1163,In_221,In_837);
nand U1164 (N_1164,In_3959,In_3552);
xnor U1165 (N_1165,In_3567,In_4291);
and U1166 (N_1166,In_1637,In_3142);
and U1167 (N_1167,In_2047,In_2655);
nand U1168 (N_1168,In_3487,In_4352);
nand U1169 (N_1169,N_164,In_3135);
or U1170 (N_1170,N_282,N_649);
and U1171 (N_1171,In_3492,N_296);
or U1172 (N_1172,N_778,In_4120);
and U1173 (N_1173,In_4095,N_64);
nor U1174 (N_1174,In_3704,In_3800);
nor U1175 (N_1175,N_693,N_868);
or U1176 (N_1176,In_289,In_2571);
or U1177 (N_1177,In_3515,N_146);
and U1178 (N_1178,In_3028,In_1657);
and U1179 (N_1179,In_1424,In_3491);
xor U1180 (N_1180,N_401,In_1085);
nor U1181 (N_1181,In_2513,N_855);
xnor U1182 (N_1182,In_4060,In_2077);
nand U1183 (N_1183,In_3986,In_2978);
or U1184 (N_1184,In_3418,N_160);
xor U1185 (N_1185,In_3114,In_616);
or U1186 (N_1186,In_795,In_796);
nor U1187 (N_1187,In_1013,In_3688);
or U1188 (N_1188,In_542,In_1847);
or U1189 (N_1189,N_768,N_230);
or U1190 (N_1190,In_1796,N_776);
xor U1191 (N_1191,In_4639,In_1670);
nand U1192 (N_1192,In_1659,In_1958);
and U1193 (N_1193,In_3979,In_4625);
or U1194 (N_1194,In_3396,In_2453);
nor U1195 (N_1195,N_362,In_1837);
or U1196 (N_1196,N_256,In_195);
nor U1197 (N_1197,In_1746,In_4521);
xnor U1198 (N_1198,In_4809,In_2019);
nor U1199 (N_1199,In_2058,In_1832);
xor U1200 (N_1200,In_1,In_276);
or U1201 (N_1201,In_3324,In_4368);
and U1202 (N_1202,N_925,In_4125);
nand U1203 (N_1203,N_316,In_2147);
or U1204 (N_1204,N_521,In_824);
or U1205 (N_1205,N_443,In_4241);
or U1206 (N_1206,In_1191,In_637);
nand U1207 (N_1207,In_2254,N_883);
xor U1208 (N_1208,In_4627,In_3253);
xnor U1209 (N_1209,In_4854,In_3485);
or U1210 (N_1210,N_538,In_3175);
nor U1211 (N_1211,In_3446,In_4219);
xnor U1212 (N_1212,N_674,In_3386);
or U1213 (N_1213,In_4778,In_3843);
or U1214 (N_1214,In_4800,In_2770);
or U1215 (N_1215,N_704,In_1490);
or U1216 (N_1216,In_2414,In_3858);
nand U1217 (N_1217,In_1625,In_305);
and U1218 (N_1218,In_3964,In_2848);
nor U1219 (N_1219,In_2619,In_4831);
nand U1220 (N_1220,In_1145,In_722);
xnor U1221 (N_1221,In_4222,In_162);
or U1222 (N_1222,N_501,In_3116);
xnor U1223 (N_1223,In_3746,In_1780);
and U1224 (N_1224,N_682,In_1577);
nor U1225 (N_1225,In_3598,In_3064);
and U1226 (N_1226,N_952,In_2604);
nand U1227 (N_1227,N_941,In_3078);
xor U1228 (N_1228,In_2447,In_3344);
and U1229 (N_1229,N_808,In_4934);
xnor U1230 (N_1230,In_4346,In_1982);
and U1231 (N_1231,N_684,In_2343);
xnor U1232 (N_1232,N_142,In_4951);
and U1233 (N_1233,In_974,In_2962);
or U1234 (N_1234,In_4424,In_3057);
nand U1235 (N_1235,In_963,In_636);
nand U1236 (N_1236,N_219,N_638);
nand U1237 (N_1237,In_3218,In_840);
or U1238 (N_1238,N_603,In_1690);
nand U1239 (N_1239,In_391,In_2461);
nor U1240 (N_1240,In_70,In_3561);
nand U1241 (N_1241,N_878,N_185);
xnor U1242 (N_1242,In_258,In_3583);
nand U1243 (N_1243,In_4229,N_770);
or U1244 (N_1244,In_4877,N_446);
nand U1245 (N_1245,In_3527,N_3);
or U1246 (N_1246,In_3015,In_1204);
xnor U1247 (N_1247,N_650,In_2687);
nand U1248 (N_1248,In_2616,N_427);
and U1249 (N_1249,In_3888,In_4536);
xnor U1250 (N_1250,In_4917,N_829);
nand U1251 (N_1251,In_936,In_1754);
and U1252 (N_1252,In_3661,In_3953);
or U1253 (N_1253,In_4383,N_36);
or U1254 (N_1254,In_4992,In_3562);
nor U1255 (N_1255,In_462,In_4806);
nor U1256 (N_1256,In_3624,N_623);
and U1257 (N_1257,N_83,In_4998);
nand U1258 (N_1258,N_821,In_2011);
nand U1259 (N_1259,In_477,In_3112);
and U1260 (N_1260,In_1149,In_1988);
xor U1261 (N_1261,In_2803,N_817);
nand U1262 (N_1262,In_3753,In_4331);
or U1263 (N_1263,N_924,In_4428);
nor U1264 (N_1264,In_2024,N_677);
xnor U1265 (N_1265,In_2056,In_2480);
and U1266 (N_1266,In_1238,N_680);
or U1267 (N_1267,N_194,In_925);
nand U1268 (N_1268,In_4544,In_71);
nor U1269 (N_1269,In_4977,In_318);
nor U1270 (N_1270,In_356,In_3541);
xnor U1271 (N_1271,N_557,In_368);
nor U1272 (N_1272,In_577,In_2660);
or U1273 (N_1273,In_1532,N_751);
xnor U1274 (N_1274,In_4216,In_2358);
or U1275 (N_1275,In_2980,In_4512);
nor U1276 (N_1276,In_3499,N_45);
xnor U1277 (N_1277,N_992,In_2929);
or U1278 (N_1278,In_413,In_4586);
nor U1279 (N_1279,In_4983,In_1027);
nor U1280 (N_1280,N_732,N_216);
nor U1281 (N_1281,In_1741,In_175);
nor U1282 (N_1282,N_754,In_252);
or U1283 (N_1283,In_2565,In_4555);
or U1284 (N_1284,N_57,In_4573);
or U1285 (N_1285,In_2339,In_3671);
and U1286 (N_1286,In_1355,In_1449);
and U1287 (N_1287,In_2046,N_707);
nor U1288 (N_1288,In_4487,In_1023);
nand U1289 (N_1289,In_2381,In_0);
and U1290 (N_1290,In_1959,In_1502);
xnor U1291 (N_1291,In_778,N_459);
nand U1292 (N_1292,In_3673,In_1158);
xnor U1293 (N_1293,In_4481,In_2477);
xnor U1294 (N_1294,In_1209,In_4477);
nand U1295 (N_1295,In_2673,In_1229);
nor U1296 (N_1296,N_79,In_3810);
nor U1297 (N_1297,N_806,In_3366);
xor U1298 (N_1298,N_568,In_4492);
xor U1299 (N_1299,In_2163,In_3734);
or U1300 (N_1300,In_409,N_47);
or U1301 (N_1301,N_696,In_4990);
nand U1302 (N_1302,In_1364,In_2557);
nand U1303 (N_1303,N_489,In_2257);
xnor U1304 (N_1304,In_1898,In_2317);
nand U1305 (N_1305,In_3505,In_3223);
xor U1306 (N_1306,In_1546,In_2263);
nor U1307 (N_1307,In_1833,In_4134);
nor U1308 (N_1308,In_397,N_882);
nor U1309 (N_1309,N_620,In_140);
nand U1310 (N_1310,In_989,In_435);
nor U1311 (N_1311,In_4533,In_1106);
nand U1312 (N_1312,In_2648,In_1980);
nand U1313 (N_1313,In_1131,N_290);
xor U1314 (N_1314,In_1506,N_238);
or U1315 (N_1315,In_4582,In_709);
xnor U1316 (N_1316,In_1037,In_2701);
nand U1317 (N_1317,In_2788,In_1721);
and U1318 (N_1318,In_2031,In_4734);
and U1319 (N_1319,In_2212,In_3268);
or U1320 (N_1320,In_2950,In_2638);
xnor U1321 (N_1321,In_1083,In_1550);
nor U1322 (N_1322,In_273,In_1759);
or U1323 (N_1323,In_4145,In_575);
xor U1324 (N_1324,N_254,In_4192);
nor U1325 (N_1325,N_626,In_937);
and U1326 (N_1326,In_4092,In_3020);
xnor U1327 (N_1327,N_796,In_2684);
nor U1328 (N_1328,In_110,N_186);
or U1329 (N_1329,In_3957,In_4021);
or U1330 (N_1330,In_1082,In_4647);
nand U1331 (N_1331,In_2837,In_2977);
or U1332 (N_1332,N_176,In_4593);
nand U1333 (N_1333,N_913,In_4396);
or U1334 (N_1334,In_1920,N_900);
nor U1335 (N_1335,In_2288,N_496);
nand U1336 (N_1336,In_2401,N_928);
and U1337 (N_1337,In_3589,In_4898);
and U1338 (N_1338,In_3758,In_2650);
and U1339 (N_1339,N_655,In_3476);
xor U1340 (N_1340,In_601,In_1134);
nor U1341 (N_1341,In_1208,In_701);
or U1342 (N_1342,In_3139,In_2487);
or U1343 (N_1343,N_833,N_473);
or U1344 (N_1344,N_298,In_1431);
xnor U1345 (N_1345,In_1169,In_3168);
xor U1346 (N_1346,In_3654,In_683);
and U1347 (N_1347,N_971,In_2580);
and U1348 (N_1348,In_3859,In_4889);
nand U1349 (N_1349,In_2704,N_193);
or U1350 (N_1350,N_547,In_3041);
nand U1351 (N_1351,In_2105,In_780);
or U1352 (N_1352,In_4911,In_501);
and U1353 (N_1353,In_149,In_3645);
or U1354 (N_1354,N_408,In_4173);
xnor U1355 (N_1355,In_122,In_2003);
nand U1356 (N_1356,In_1049,In_4987);
nor U1357 (N_1357,In_2380,In_3867);
nor U1358 (N_1358,N_699,In_3427);
xor U1359 (N_1359,In_1242,In_576);
nor U1360 (N_1360,In_3384,N_98);
nand U1361 (N_1361,In_3224,N_903);
xor U1362 (N_1362,In_3051,N_66);
xnor U1363 (N_1363,In_113,In_2920);
nor U1364 (N_1364,In_3999,N_382);
and U1365 (N_1365,In_2716,In_2637);
xor U1366 (N_1366,In_3735,N_80);
xnor U1367 (N_1367,In_3173,In_1211);
or U1368 (N_1368,In_52,N_936);
xnor U1369 (N_1369,In_1889,In_4787);
nor U1370 (N_1370,In_253,In_3025);
or U1371 (N_1371,In_4039,In_2067);
and U1372 (N_1372,In_1504,In_4563);
nor U1373 (N_1373,In_4720,In_2847);
or U1374 (N_1374,In_1895,In_4014);
and U1375 (N_1375,In_620,In_3211);
nor U1376 (N_1376,N_827,In_2118);
or U1377 (N_1377,In_3963,In_944);
and U1378 (N_1378,In_4370,In_3709);
xor U1379 (N_1379,In_1357,In_3563);
or U1380 (N_1380,In_4094,In_2718);
nand U1381 (N_1381,In_4796,In_3432);
nor U1382 (N_1382,In_4905,In_3889);
nand U1383 (N_1383,In_4022,N_111);
and U1384 (N_1384,N_42,N_801);
nand U1385 (N_1385,In_4900,N_836);
and U1386 (N_1386,In_2219,In_2040);
and U1387 (N_1387,In_3532,In_72);
nand U1388 (N_1388,In_2625,N_449);
nand U1389 (N_1389,In_1799,In_4844);
nand U1390 (N_1390,In_1947,In_3733);
nand U1391 (N_1391,In_2764,In_2814);
nor U1392 (N_1392,In_4322,In_1160);
nand U1393 (N_1393,In_4776,N_810);
nor U1394 (N_1394,In_2261,In_4374);
nand U1395 (N_1395,In_3392,In_2353);
nand U1396 (N_1396,In_481,In_4510);
nor U1397 (N_1397,In_2195,In_581);
nand U1398 (N_1398,In_493,In_4054);
nor U1399 (N_1399,In_2374,N_444);
nand U1400 (N_1400,In_2308,In_4912);
or U1401 (N_1401,N_58,N_9);
and U1402 (N_1402,In_1157,In_3214);
or U1403 (N_1403,N_389,N_43);
and U1404 (N_1404,In_3084,In_907);
or U1405 (N_1405,In_1250,N_625);
nand U1406 (N_1406,In_1125,In_1584);
and U1407 (N_1407,In_4955,In_2489);
xnor U1408 (N_1408,In_2983,In_3372);
xnor U1409 (N_1409,N_472,In_2391);
or U1410 (N_1410,In_2688,In_4321);
xor U1411 (N_1411,In_1410,In_1370);
and U1412 (N_1412,In_2076,In_521);
nand U1413 (N_1413,In_3415,In_1003);
xor U1414 (N_1414,In_296,In_3498);
or U1415 (N_1415,In_3711,In_3717);
and U1416 (N_1416,In_2643,In_353);
nor U1417 (N_1417,In_4418,In_524);
or U1418 (N_1418,In_2523,N_687);
or U1419 (N_1419,In_243,In_1681);
or U1420 (N_1420,In_3689,In_2023);
and U1421 (N_1421,N_799,In_4342);
nor U1422 (N_1422,In_4122,In_661);
nor U1423 (N_1423,In_4205,In_2969);
nor U1424 (N_1424,N_815,In_1695);
nand U1425 (N_1425,In_228,In_2407);
xor U1426 (N_1426,In_3718,In_57);
nand U1427 (N_1427,In_3475,In_330);
or U1428 (N_1428,N_667,In_2121);
xor U1429 (N_1429,In_635,In_2113);
nand U1430 (N_1430,In_2939,In_3523);
and U1431 (N_1431,N_940,In_1468);
xnor U1432 (N_1432,In_1971,In_1564);
or U1433 (N_1433,N_504,N_93);
and U1434 (N_1434,In_4444,In_3737);
xor U1435 (N_1435,In_3910,In_4425);
nor U1436 (N_1436,In_1801,In_1910);
nand U1437 (N_1437,In_1376,In_231);
nand U1438 (N_1438,In_4431,In_1112);
or U1439 (N_1439,N_138,N_962);
nand U1440 (N_1440,In_4601,In_1888);
nand U1441 (N_1441,N_169,N_115);
nand U1442 (N_1442,In_1285,In_3670);
and U1443 (N_1443,N_351,In_2535);
nor U1444 (N_1444,In_1295,In_4636);
xnor U1445 (N_1445,In_4841,In_2538);
nor U1446 (N_1446,In_2128,In_1644);
xnor U1447 (N_1447,In_161,N_909);
nor U1448 (N_1448,In_505,In_4857);
nand U1449 (N_1449,In_4789,N_23);
nor U1450 (N_1450,In_3276,In_4445);
nor U1451 (N_1451,In_2239,In_4043);
nand U1452 (N_1452,In_2065,In_3377);
xor U1453 (N_1453,In_3535,In_1586);
or U1454 (N_1454,In_3996,In_55);
nor U1455 (N_1455,In_4981,In_3716);
and U1456 (N_1456,N_562,N_760);
and U1457 (N_1457,In_1034,In_1840);
or U1458 (N_1458,N_870,In_4405);
and U1459 (N_1459,N_867,In_340);
and U1460 (N_1460,In_2628,In_1126);
nand U1461 (N_1461,N_468,In_238);
nand U1462 (N_1462,In_4910,In_4319);
nand U1463 (N_1463,In_4819,In_1155);
nand U1464 (N_1464,In_3466,In_4503);
and U1465 (N_1465,In_3846,In_4183);
or U1466 (N_1466,N_690,In_456);
nand U1467 (N_1467,In_596,In_1752);
nor U1468 (N_1468,In_764,In_531);
xor U1469 (N_1469,In_4960,N_991);
nand U1470 (N_1470,In_293,In_373);
nor U1471 (N_1471,In_1389,In_2626);
or U1472 (N_1472,In_4689,N_676);
and U1473 (N_1473,In_3063,In_3824);
xor U1474 (N_1474,N_241,In_3037);
xor U1475 (N_1475,In_1804,N_947);
xor U1476 (N_1476,In_2209,In_2091);
and U1477 (N_1477,In_183,In_1749);
nand U1478 (N_1478,In_133,In_525);
and U1479 (N_1479,N_558,In_3713);
nor U1480 (N_1480,In_3177,In_3745);
nand U1481 (N_1481,In_2566,N_966);
nand U1482 (N_1482,In_1111,In_3873);
or U1483 (N_1483,N_594,In_1559);
nand U1484 (N_1484,In_4855,In_3590);
and U1485 (N_1485,N_942,In_4010);
nor U1486 (N_1486,In_1130,In_529);
xor U1487 (N_1487,In_2465,N_997);
nand U1488 (N_1488,N_125,In_4460);
nand U1489 (N_1489,In_4600,In_2986);
nand U1490 (N_1490,In_4901,In_1717);
xnor U1491 (N_1491,In_3775,In_4267);
or U1492 (N_1492,In_4678,N_128);
nand U1493 (N_1493,In_2371,In_4967);
xnor U1494 (N_1494,In_4293,In_2875);
nor U1495 (N_1495,In_3088,In_12);
and U1496 (N_1496,In_2099,In_1650);
nand U1497 (N_1497,N_983,In_4624);
and U1498 (N_1498,In_3095,In_3086);
nand U1499 (N_1499,In_290,In_3035);
xnor U1500 (N_1500,In_4274,In_4458);
nand U1501 (N_1501,In_2830,N_1086);
nand U1502 (N_1502,In_189,N_1264);
nand U1503 (N_1503,N_614,In_1020);
nand U1504 (N_1504,In_1269,N_1090);
xnor U1505 (N_1505,N_1222,N_532);
or U1506 (N_1506,N_131,N_200);
nor U1507 (N_1507,In_3120,N_338);
nand U1508 (N_1508,N_1339,In_4227);
nand U1509 (N_1509,In_4668,N_802);
or U1510 (N_1510,N_225,N_654);
or U1511 (N_1511,N_689,In_104);
nor U1512 (N_1512,N_534,N_843);
nor U1513 (N_1513,N_844,N_1462);
nand U1514 (N_1514,In_3626,N_1192);
and U1515 (N_1515,N_1356,In_4268);
nor U1516 (N_1516,N_1459,N_1220);
nand U1517 (N_1517,N_919,In_1384);
and U1518 (N_1518,N_896,In_2303);
xnor U1519 (N_1519,In_1626,In_2809);
or U1520 (N_1520,N_1396,N_1053);
nand U1521 (N_1521,In_1476,In_381);
or U1522 (N_1522,N_129,In_1129);
nand U1523 (N_1523,N_1335,In_223);
nand U1524 (N_1524,N_943,In_192);
or U1525 (N_1525,In_3170,N_1385);
and U1526 (N_1526,In_1948,N_264);
and U1527 (N_1527,In_1186,In_3097);
or U1528 (N_1528,In_1758,In_2305);
nand U1529 (N_1529,N_1226,In_2671);
and U1530 (N_1530,N_824,In_3488);
nand U1531 (N_1531,In_3712,In_591);
nor U1532 (N_1532,In_1772,In_653);
or U1533 (N_1533,In_2560,In_1881);
nor U1534 (N_1534,In_4642,N_1398);
or U1535 (N_1535,In_4930,In_2955);
and U1536 (N_1536,In_1892,N_502);
and U1537 (N_1537,In_294,In_3087);
nor U1538 (N_1538,N_1415,N_196);
nor U1539 (N_1539,In_4046,N_127);
nand U1540 (N_1540,In_4739,In_3012);
nand U1541 (N_1541,N_201,N_790);
and U1542 (N_1542,N_1293,In_2102);
nand U1543 (N_1543,In_3835,In_3111);
xnor U1544 (N_1544,In_2956,N_1369);
and U1545 (N_1545,In_2786,In_1762);
and U1546 (N_1546,N_412,In_1933);
nand U1547 (N_1547,In_1890,In_2609);
xnor U1548 (N_1548,N_438,In_3978);
or U1549 (N_1549,N_1237,In_3938);
nand U1550 (N_1550,N_856,In_4557);
nand U1551 (N_1551,In_3138,In_4423);
nor U1552 (N_1552,In_2966,N_1471);
and U1553 (N_1553,N_510,In_4343);
xnor U1554 (N_1554,In_4493,In_4119);
or U1555 (N_1555,N_748,In_3941);
or U1556 (N_1556,In_4896,N_1382);
or U1557 (N_1557,In_3381,In_4495);
and U1558 (N_1558,In_3152,In_4217);
nand U1559 (N_1559,In_4208,In_1192);
and U1560 (N_1560,In_2104,In_3772);
nor U1561 (N_1561,In_4067,In_1649);
and U1562 (N_1562,N_528,N_1418);
nor U1563 (N_1563,In_2496,In_1764);
nor U1564 (N_1564,N_506,N_636);
and U1565 (N_1565,In_1090,In_4631);
nand U1566 (N_1566,In_1408,N_1067);
nand U1567 (N_1567,In_2810,In_1853);
nor U1568 (N_1568,N_189,N_1158);
nor U1569 (N_1569,In_2844,In_4974);
or U1570 (N_1570,In_4324,In_3375);
and U1571 (N_1571,In_973,N_1492);
or U1572 (N_1572,In_3879,In_2397);
xnor U1573 (N_1573,In_47,In_2411);
and U1574 (N_1574,N_1243,In_3725);
nand U1575 (N_1575,In_496,In_1987);
nand U1576 (N_1576,In_3266,In_3348);
or U1577 (N_1577,N_118,In_1667);
xnor U1578 (N_1578,In_872,In_1417);
and U1579 (N_1579,In_4774,In_3137);
xnor U1580 (N_1580,In_320,N_954);
or U1581 (N_1581,N_948,N_820);
or U1582 (N_1582,In_3260,In_1880);
nand U1583 (N_1583,In_2186,N_577);
and U1584 (N_1584,In_3575,In_1127);
nand U1585 (N_1585,In_3849,In_2470);
xor U1586 (N_1586,In_1864,In_1213);
xnor U1587 (N_1587,N_1172,In_359);
nand U1588 (N_1588,In_1395,In_2220);
nand U1589 (N_1589,In_3700,In_1885);
nand U1590 (N_1590,In_7,In_4956);
xnor U1591 (N_1591,N_233,In_4546);
xor U1592 (N_1592,In_2134,In_2632);
or U1593 (N_1593,In_1433,In_3923);
and U1594 (N_1594,In_1099,In_421);
nor U1595 (N_1595,In_1178,In_1575);
xnor U1596 (N_1596,In_395,In_3198);
xnor U1597 (N_1597,N_257,N_415);
xor U1598 (N_1598,In_2911,In_4985);
nor U1599 (N_1599,In_534,N_860);
xor U1600 (N_1600,In_3395,In_1610);
nor U1601 (N_1601,In_2745,In_2882);
or U1602 (N_1602,In_3977,In_2467);
and U1603 (N_1603,In_4835,N_915);
nand U1604 (N_1604,In_4273,N_410);
nor U1605 (N_1605,In_1857,N_1412);
and U1606 (N_1606,In_1793,N_712);
nor U1607 (N_1607,In_1647,N_380);
nor U1608 (N_1608,In_2709,N_1112);
nand U1609 (N_1609,N_977,N_1397);
and U1610 (N_1610,In_4978,N_832);
xor U1611 (N_1611,In_3473,In_1591);
nor U1612 (N_1612,N_1239,In_503);
xor U1613 (N_1613,N_1413,In_3954);
and U1614 (N_1614,In_3441,N_429);
or U1615 (N_1615,N_240,In_4356);
nor U1616 (N_1616,In_2511,N_544);
and U1617 (N_1617,N_1159,In_2439);
xor U1618 (N_1618,In_4148,In_211);
or U1619 (N_1619,In_3315,N_872);
nand U1620 (N_1620,N_515,In_3302);
or U1621 (N_1621,N_130,N_1177);
xor U1622 (N_1622,In_3199,N_377);
nand U1623 (N_1623,In_4179,In_4105);
nand U1624 (N_1624,In_4534,N_1267);
nor U1625 (N_1625,In_2069,In_4520);
xnor U1626 (N_1626,In_2938,N_639);
or U1627 (N_1627,N_523,In_1995);
xnor U1628 (N_1628,In_952,In_2642);
xor U1629 (N_1629,N_293,N_1355);
xor U1630 (N_1630,In_4251,In_2457);
nand U1631 (N_1631,In_859,In_492);
or U1632 (N_1632,In_2042,In_2840);
and U1633 (N_1633,In_3029,N_461);
nor U1634 (N_1634,In_4221,N_1031);
xnor U1635 (N_1635,In_219,In_3090);
nor U1636 (N_1636,N_205,In_2384);
and U1637 (N_1637,In_3731,In_3197);
nor U1638 (N_1638,N_901,In_1715);
or U1639 (N_1639,N_345,N_1449);
or U1640 (N_1640,N_1149,N_607);
nand U1641 (N_1641,In_1021,In_3094);
or U1642 (N_1642,In_1582,In_3883);
nand U1643 (N_1643,In_3321,In_1289);
nand U1644 (N_1644,In_2326,In_479);
xor U1645 (N_1645,In_2445,In_2504);
and U1646 (N_1646,In_3898,N_1277);
nand U1647 (N_1647,In_4765,In_1274);
and U1648 (N_1648,In_4513,In_1536);
and U1649 (N_1649,In_4168,In_2590);
or U1650 (N_1650,In_1442,In_2365);
nor U1651 (N_1651,In_2230,In_4456);
nand U1652 (N_1652,In_2715,N_426);
xnor U1653 (N_1653,N_1423,N_300);
or U1654 (N_1654,In_1097,In_3558);
or U1655 (N_1655,In_1303,In_3050);
nand U1656 (N_1656,In_3500,In_4196);
and U1657 (N_1657,In_4938,N_1371);
and U1658 (N_1658,N_44,N_404);
nor U1659 (N_1659,N_822,In_225);
xnor U1660 (N_1660,In_2312,N_1332);
xor U1661 (N_1661,N_311,In_4485);
xnor U1662 (N_1662,N_223,N_503);
nand U1663 (N_1663,N_1163,In_4034);
nand U1664 (N_1664,In_80,N_1093);
xor U1665 (N_1665,In_951,In_1462);
nor U1666 (N_1666,N_1170,In_3642);
nor U1667 (N_1667,In_1175,In_1727);
xnor U1668 (N_1668,N_1141,In_1026);
nor U1669 (N_1669,In_2815,N_531);
and U1670 (N_1670,In_4401,In_1464);
xor U1671 (N_1671,N_1051,N_270);
nor U1672 (N_1672,In_1304,In_3668);
nor U1673 (N_1673,In_3317,In_1696);
and U1674 (N_1674,N_537,In_2088);
or U1675 (N_1675,In_4419,In_3680);
and U1676 (N_1676,N_332,In_4053);
and U1677 (N_1677,In_1976,In_3848);
nand U1678 (N_1678,N_779,N_794);
xnor U1679 (N_1679,N_374,In_849);
nor U1680 (N_1680,N_1127,In_1557);
and U1681 (N_1681,In_1585,In_331);
nand U1682 (N_1682,In_3379,In_1965);
and U1683 (N_1683,In_4821,In_1688);
xnor U1684 (N_1684,In_4104,N_358);
nor U1685 (N_1685,In_1374,N_212);
xnor U1686 (N_1686,In_1497,In_3158);
nand U1687 (N_1687,N_543,N_365);
and U1688 (N_1688,In_2515,In_3265);
xor U1689 (N_1689,In_2000,In_4127);
nand U1690 (N_1690,N_392,In_3765);
and U1691 (N_1691,N_905,N_1054);
and U1692 (N_1692,In_3171,In_17);
or U1693 (N_1693,In_2818,In_3572);
xnor U1694 (N_1694,In_3839,In_3113);
xor U1695 (N_1695,In_3834,In_2180);
or U1696 (N_1696,In_1481,In_1225);
xnor U1697 (N_1697,In_1541,N_119);
xor U1698 (N_1698,In_200,In_2108);
xor U1699 (N_1699,In_3815,In_193);
nand U1700 (N_1700,In_572,In_1093);
nor U1701 (N_1701,N_1359,N_400);
nand U1702 (N_1702,N_1061,In_3482);
xor U1703 (N_1703,In_3408,In_615);
or U1704 (N_1704,In_2667,N_1231);
nor U1705 (N_1705,N_1255,N_1399);
and U1706 (N_1706,N_564,In_537);
nor U1707 (N_1707,In_3005,In_4823);
and U1708 (N_1708,N_858,In_1954);
and U1709 (N_1709,In_4140,In_2142);
nand U1710 (N_1710,N_269,In_1139);
nand U1711 (N_1711,In_2959,In_2085);
xnor U1712 (N_1712,In_2727,N_1368);
nand U1713 (N_1713,In_1590,In_4915);
or U1714 (N_1714,N_1358,N_405);
xor U1715 (N_1715,In_307,N_416);
and U1716 (N_1716,In_212,In_2585);
nand U1717 (N_1717,In_949,In_2229);
xor U1718 (N_1718,In_3790,In_457);
nand U1719 (N_1719,N_599,In_375);
xor U1720 (N_1720,In_1058,In_4965);
nor U1721 (N_1721,In_3174,N_475);
nor U1722 (N_1722,In_3271,N_1084);
nand U1723 (N_1723,N_1370,In_4376);
nor U1724 (N_1724,N_771,N_1183);
nor U1725 (N_1725,In_513,In_1190);
and U1726 (N_1726,In_1463,In_3905);
xor U1727 (N_1727,In_3769,In_1069);
or U1728 (N_1728,N_1169,N_168);
xor U1729 (N_1729,In_3796,In_386);
and U1730 (N_1730,N_1401,In_3144);
and U1731 (N_1731,N_1227,In_2344);
xor U1732 (N_1732,In_2243,N_481);
or U1733 (N_1733,In_1921,In_1120);
xor U1734 (N_1734,In_4849,In_420);
or U1735 (N_1735,In_1258,In_3460);
or U1736 (N_1736,N_1121,N_1033);
nand U1737 (N_1737,In_4553,N_272);
or U1738 (N_1738,In_360,In_518);
nand U1739 (N_1739,In_3987,In_2017);
nand U1740 (N_1740,In_1687,N_329);
nor U1741 (N_1741,In_1343,In_2119);
or U1742 (N_1742,In_2395,In_2696);
nor U1743 (N_1743,In_2608,In_988);
xor U1744 (N_1744,In_4617,In_2532);
and U1745 (N_1745,N_921,N_1039);
nand U1746 (N_1746,In_31,N_1016);
and U1747 (N_1747,In_2196,N_226);
xor U1748 (N_1748,In_1121,In_2658);
or U1749 (N_1749,N_1034,In_3285);
nor U1750 (N_1750,N_306,In_4262);
nand U1751 (N_1751,In_2781,N_1354);
xnor U1752 (N_1752,N_343,In_364);
nand U1753 (N_1753,In_2187,In_2720);
xnor U1754 (N_1754,In_388,N_555);
nor U1755 (N_1755,In_2686,N_1353);
nand U1756 (N_1756,N_1457,In_2546);
or U1757 (N_1757,In_3406,In_2670);
xor U1758 (N_1758,N_287,In_2238);
nor U1759 (N_1759,In_3439,In_2044);
and U1760 (N_1760,N_1338,In_4578);
and U1761 (N_1761,In_4031,In_3757);
nor U1762 (N_1762,In_803,N_955);
nor U1763 (N_1763,N_756,In_2120);
and U1764 (N_1764,In_3082,In_2430);
or U1765 (N_1765,N_337,N_106);
nor U1766 (N_1766,In_467,In_4215);
or U1767 (N_1767,In_3371,In_3282);
nand U1768 (N_1768,In_3968,In_4785);
xnor U1769 (N_1769,In_3468,N_1325);
xnor U1770 (N_1770,In_459,In_2573);
nand U1771 (N_1771,In_4240,In_215);
and U1772 (N_1772,N_706,In_1089);
nand U1773 (N_1773,N_569,N_830);
and U1774 (N_1774,N_1087,In_1869);
nor U1775 (N_1775,In_4670,In_3929);
xor U1776 (N_1776,N_673,N_1210);
or U1777 (N_1777,In_1960,In_2255);
xnor U1778 (N_1778,In_2213,N_179);
nor U1779 (N_1779,N_1225,N_411);
or U1780 (N_1780,N_1156,In_2363);
nand U1781 (N_1781,N_99,In_2751);
xnor U1782 (N_1782,In_2550,In_3920);
nor U1783 (N_1783,N_644,In_3404);
or U1784 (N_1784,In_3252,In_2501);
nand U1785 (N_1785,In_3684,N_304);
nor U1786 (N_1786,In_25,In_1943);
nand U1787 (N_1787,In_2096,In_3901);
nor U1788 (N_1788,In_3143,In_873);
nor U1789 (N_1789,In_4680,N_1060);
or U1790 (N_1790,In_4509,N_33);
nand U1791 (N_1791,In_4011,In_3648);
or U1792 (N_1792,N_462,N_7);
or U1793 (N_1793,In_2836,In_4741);
xnor U1794 (N_1794,In_442,N_1345);
nand U1795 (N_1795,In_801,N_713);
or U1796 (N_1796,In_1630,N_1167);
or U1797 (N_1797,In_4991,In_1694);
or U1798 (N_1798,In_4726,In_2375);
nand U1799 (N_1799,In_4694,In_812);
nor U1800 (N_1800,N_499,N_854);
nor U1801 (N_1801,N_747,In_3629);
nand U1802 (N_1802,N_1019,N_460);
xor U1803 (N_1803,In_3256,In_3337);
nor U1804 (N_1804,N_1063,In_4381);
nor U1805 (N_1805,In_2856,In_4750);
nor U1806 (N_1806,N_1433,In_913);
and U1807 (N_1807,N_430,N_1321);
xnor U1808 (N_1808,N_454,N_1253);
and U1809 (N_1809,N_853,In_1906);
xnor U1810 (N_1810,In_4549,In_4359);
or U1811 (N_1811,In_2423,In_654);
or U1812 (N_1812,N_920,In_3284);
and U1813 (N_1813,In_991,In_4872);
or U1814 (N_1814,In_3656,In_691);
nand U1815 (N_1815,In_4411,In_2519);
or U1816 (N_1816,In_4245,In_4733);
nand U1817 (N_1817,In_718,In_3463);
and U1818 (N_1818,In_2551,In_2321);
nand U1819 (N_1819,In_2763,In_185);
or U1820 (N_1820,In_464,In_1256);
and U1821 (N_1821,N_41,In_4779);
and U1822 (N_1822,In_4828,In_1421);
and U1823 (N_1823,N_322,N_1299);
and U1824 (N_1824,N_500,In_2971);
and U1825 (N_1825,In_888,In_2755);
and U1826 (N_1826,In_2432,In_1422);
xor U1827 (N_1827,N_1250,In_2568);
nor U1828 (N_1828,N_1326,In_1708);
xor U1829 (N_1829,In_1346,In_1253);
and U1830 (N_1830,In_2802,N_20);
xnor U1831 (N_1831,N_581,In_1929);
nor U1832 (N_1832,N_1197,N_630);
nand U1833 (N_1833,In_1703,In_126);
nand U1834 (N_1834,In_754,In_4111);
or U1835 (N_1835,N_841,In_312);
xnor U1836 (N_1836,In_4699,In_1499);
nor U1837 (N_1837,In_1011,N_1188);
nand U1838 (N_1838,In_945,N_372);
xor U1839 (N_1839,In_4364,In_4522);
and U1840 (N_1840,N_819,In_4441);
nor U1841 (N_1841,In_2623,In_3031);
or U1842 (N_1842,In_4447,N_1404);
or U1843 (N_1843,N_402,In_3264);
nor U1844 (N_1844,In_3555,In_898);
and U1845 (N_1845,In_2232,In_349);
nor U1846 (N_1846,N_1296,N_1107);
or U1847 (N_1847,In_4777,In_2828);
or U1848 (N_1848,In_4530,In_579);
nor U1849 (N_1849,N_1373,In_3336);
and U1850 (N_1850,In_4410,N_1070);
and U1851 (N_1851,N_16,N_1273);
or U1852 (N_1852,In_158,In_4285);
nor U1853 (N_1853,In_4658,N_722);
nand U1854 (N_1854,In_4369,N_396);
and U1855 (N_1855,N_731,In_2404);
and U1856 (N_1856,In_2095,In_372);
and U1857 (N_1857,In_2953,In_2270);
nand U1858 (N_1858,In_3385,N_341);
or U1859 (N_1859,In_4941,In_1070);
and U1860 (N_1860,In_1563,In_3461);
and U1861 (N_1861,In_3233,In_1201);
nor U1862 (N_1862,In_3428,N_879);
and U1863 (N_1863,In_4073,In_27);
nand U1864 (N_1864,In_1555,N_1182);
nand U1865 (N_1865,In_3797,In_4970);
or U1866 (N_1866,In_658,N_17);
xor U1867 (N_1867,In_3857,In_4339);
nand U1868 (N_1868,In_2710,N_324);
nand U1869 (N_1869,In_3483,In_1969);
xor U1870 (N_1870,In_3294,In_2233);
xor U1871 (N_1871,In_881,N_840);
nor U1872 (N_1872,In_1726,In_2292);
nand U1873 (N_1873,In_2351,In_2884);
or U1874 (N_1874,N_1035,In_3013);
and U1875 (N_1875,In_3027,In_429);
xnor U1876 (N_1876,In_4003,N_1244);
xor U1877 (N_1877,N_136,In_1168);
or U1878 (N_1878,N_1286,In_4300);
nor U1879 (N_1879,In_1226,N_1317);
xor U1880 (N_1880,In_3455,In_2482);
and U1881 (N_1881,N_1337,In_1994);
nor U1882 (N_1882,In_1227,N_530);
nand U1883 (N_1883,N_477,In_552);
xnor U1884 (N_1884,In_3971,N_1146);
nor U1885 (N_1885,N_1258,In_1056);
and U1886 (N_1886,N_367,In_2849);
or U1887 (N_1887,In_4158,In_4488);
or U1888 (N_1888,In_148,In_995);
xor U1889 (N_1889,N_235,N_1302);
and U1890 (N_1890,In_4029,In_3650);
nor U1891 (N_1891,In_370,N_786);
xnor U1892 (N_1892,In_4811,In_1177);
and U1893 (N_1893,N_52,In_2569);
xor U1894 (N_1894,In_549,In_490);
and U1895 (N_1895,In_2206,In_3043);
nand U1896 (N_1896,In_4288,In_4808);
xnor U1897 (N_1897,In_602,N_695);
nand U1898 (N_1898,In_4472,N_857);
xor U1899 (N_1899,N_188,In_4665);
xor U1900 (N_1900,In_4669,In_3248);
or U1901 (N_1901,N_249,N_1360);
nor U1902 (N_1902,In_1863,In_3129);
or U1903 (N_1903,N_470,In_740);
and U1904 (N_1904,In_1110,In_3409);
nand U1905 (N_1905,In_3917,N_1110);
and U1906 (N_1906,N_798,In_306);
nand U1907 (N_1907,In_938,In_3368);
nand U1908 (N_1908,N_629,In_604);
and U1909 (N_1909,In_3793,In_1176);
nand U1910 (N_1910,In_1302,In_2247);
xor U1911 (N_1911,In_327,N_791);
or U1912 (N_1912,N_1007,In_1571);
and U1913 (N_1913,N_1123,N_1466);
xnor U1914 (N_1914,In_595,In_84);
nor U1915 (N_1915,In_3721,In_1137);
or U1916 (N_1916,In_466,N_1435);
and U1917 (N_1917,In_880,In_426);
nor U1918 (N_1918,N_480,N_916);
or U1919 (N_1919,In_3243,N_1128);
nand U1920 (N_1920,In_3151,N_784);
xor U1921 (N_1921,N_850,In_1051);
nor U1922 (N_1922,In_825,N_765);
xnor U1923 (N_1923,N_1460,In_3574);
and U1924 (N_1924,In_2570,N_812);
nor U1925 (N_1925,N_1021,In_392);
or U1926 (N_1926,In_2478,In_1934);
nand U1927 (N_1927,In_3403,In_2584);
nand U1928 (N_1928,N_1234,N_339);
and U1929 (N_1929,In_3806,In_3356);
or U1930 (N_1930,In_4537,In_1406);
xnor U1931 (N_1931,In_2753,In_4116);
xor U1932 (N_1932,In_1062,In_2589);
xor U1933 (N_1933,N_527,In_1115);
nor U1934 (N_1934,In_606,N_1327);
xor U1935 (N_1935,In_4953,In_485);
nor U1936 (N_1936,N_982,In_3871);
xor U1937 (N_1937,In_4997,In_3580);
or U1938 (N_1938,N_1477,In_4328);
xor U1939 (N_1939,In_4090,N_1464);
nand U1940 (N_1940,In_181,N_1486);
nor U1941 (N_1941,N_912,In_2218);
xnor U1942 (N_1942,In_4591,N_1083);
xnor U1943 (N_1943,In_3974,N_513);
or U1944 (N_1944,In_3675,In_1324);
xor U1945 (N_1945,In_3201,N_398);
or U1946 (N_1946,N_1095,N_598);
nand U1947 (N_1947,N_342,In_2993);
nand U1948 (N_1948,In_739,In_1938);
xnor U1949 (N_1949,N_1322,In_1043);
nand U1950 (N_1950,In_1340,In_4077);
xnor U1951 (N_1951,In_2854,In_747);
nand U1952 (N_1952,In_1588,N_847);
nand U1953 (N_1953,In_4136,In_4940);
xnor U1954 (N_1954,In_2028,N_683);
or U1955 (N_1955,In_3516,In_2055);
and U1956 (N_1956,In_2661,N_30);
xor U1957 (N_1957,In_4184,In_511);
nor U1958 (N_1958,In_2347,In_3495);
xor U1959 (N_1959,N_207,In_261);
and U1960 (N_1960,In_4838,N_105);
nor U1961 (N_1961,N_642,In_2896);
xnor U1962 (N_1962,In_3169,N_1303);
nor U1963 (N_1963,In_4848,N_1406);
nor U1964 (N_1964,In_4868,In_2541);
xnor U1965 (N_1965,N_1272,In_1098);
nand U1966 (N_1966,N_967,In_860);
nor U1967 (N_1967,In_1579,N_848);
or U1968 (N_1968,In_3534,In_1327);
nor U1969 (N_1969,N_665,N_1044);
nand U1970 (N_1970,N_153,In_1314);
or U1971 (N_1971,In_2997,In_1245);
or U1972 (N_1972,N_615,N_1440);
or U1973 (N_1973,In_2466,N_964);
xnor U1974 (N_1974,In_3261,N_1014);
xor U1975 (N_1975,In_1404,N_551);
nor U1976 (N_1976,N_1100,In_2775);
or U1977 (N_1977,N_1268,In_640);
and U1978 (N_1978,In_1445,In_3136);
or U1979 (N_1979,N_1281,N_1394);
xnor U1980 (N_1980,N_561,In_2902);
nand U1981 (N_1981,In_3702,N_1498);
xor U1982 (N_1982,N_110,N_612);
and U1983 (N_1983,In_3014,In_2611);
nor U1984 (N_1984,In_2068,In_1344);
xor U1985 (N_1985,N_1193,N_659);
nand U1986 (N_1986,In_1633,In_4497);
nor U1987 (N_1987,N_1297,In_3660);
xor U1988 (N_1988,In_1350,In_2492);
and U1989 (N_1989,In_2857,In_3861);
nor U1990 (N_1990,N_675,In_956);
and U1991 (N_1991,N_838,In_2018);
or U1992 (N_1992,N_520,In_4645);
xnor U1993 (N_1993,In_2713,In_2811);
nand U1994 (N_1994,In_1337,In_92);
nand U1995 (N_1995,In_2885,In_3325);
and U1996 (N_1996,N_1161,N_1386);
xnor U1997 (N_1997,In_3695,N_1147);
nor U1998 (N_1998,In_2864,N_1022);
and U1999 (N_1999,N_1262,In_4839);
and U2000 (N_2000,In_2103,N_1576);
and U2001 (N_2001,N_1470,N_1687);
or U2002 (N_2002,In_259,In_1007);
xor U2003 (N_2003,In_443,In_1084);
nor U2004 (N_2004,In_3024,In_4325);
nand U2005 (N_2005,In_1195,N_463);
nor U2006 (N_2006,In_3289,N_1826);
and U2007 (N_2007,In_4258,In_2607);
or U2008 (N_2008,N_1426,N_250);
nand U2009 (N_2009,N_1455,N_1521);
nand U2010 (N_2010,In_4822,N_837);
or U2011 (N_2011,N_1768,In_2647);
nor U2012 (N_2012,In_3433,In_1259);
xnor U2013 (N_2013,N_1181,N_162);
nor U2014 (N_2014,N_1740,N_1764);
and U2015 (N_2015,In_3587,N_1407);
or U2016 (N_2016,N_1391,In_3729);
xnor U2017 (N_2017,In_232,In_4864);
nor U2018 (N_2018,In_2319,In_874);
xor U2019 (N_2019,N_1165,In_3600);
nand U2020 (N_2020,In_4129,N_1940);
or U2021 (N_2021,N_1289,N_1658);
xor U2022 (N_2022,N_1381,In_1018);
nand U2023 (N_2023,In_2468,In_1450);
or U2024 (N_2024,N_1806,In_588);
or U2025 (N_2025,N_842,In_83);
and U2026 (N_2026,In_2627,N_149);
nand U2027 (N_2027,In_4722,N_1876);
or U2028 (N_2028,In_2287,N_618);
nand U2029 (N_2029,In_2094,N_1);
nor U2030 (N_2030,N_1164,In_662);
or U2031 (N_2031,N_1730,In_891);
xor U2032 (N_2032,In_896,In_1573);
xor U2033 (N_2033,In_3044,In_4143);
and U2034 (N_2034,N_40,In_976);
and U2035 (N_2035,In_77,In_941);
nand U2036 (N_2036,In_607,In_1523);
xor U2037 (N_2037,N_1856,N_807);
or U2038 (N_2038,In_430,N_643);
or U2039 (N_2039,N_927,In_3322);
or U2040 (N_2040,In_1447,In_4966);
or U2041 (N_2041,In_2737,N_1364);
xor U2042 (N_2042,In_2999,In_4250);
or U2043 (N_2043,In_1167,In_4326);
or U2044 (N_2044,N_1285,In_1918);
xnor U2045 (N_2045,In_2871,N_1746);
nor U2046 (N_2046,N_960,In_670);
nand U2047 (N_2047,N_1976,In_3092);
nand U2048 (N_2048,N_1300,In_2471);
nor U2049 (N_2049,In_4643,N_1079);
nand U2050 (N_2050,In_3327,In_2315);
xor U2051 (N_2051,In_4189,N_1504);
nor U2052 (N_2052,N_314,In_3994);
and U2053 (N_2053,In_2225,N_1424);
nand U2054 (N_2054,In_4350,N_1995);
nand U2055 (N_2055,N_1047,N_1632);
nor U2056 (N_2056,In_2576,In_2234);
nor U2057 (N_2057,In_2942,In_1492);
nor U2058 (N_2058,In_100,N_1130);
or U2059 (N_2059,N_1291,In_4574);
or U2060 (N_2060,In_876,In_38);
and U2061 (N_2061,In_374,In_1851);
and U2062 (N_2062,In_4950,N_679);
xor U2063 (N_2063,In_3913,N_1994);
nor U2064 (N_2064,In_1705,N_579);
nor U2065 (N_2065,N_1133,N_661);
xor U2066 (N_2066,In_324,N_39);
nor U2067 (N_2067,In_1437,N_1062);
nand U2068 (N_2068,N_518,N_512);
xnor U2069 (N_2069,N_1419,N_1254);
xor U2070 (N_2070,N_893,N_344);
or U2071 (N_2071,N_759,N_21);
nand U2072 (N_2072,In_351,In_3694);
xnor U2073 (N_2073,N_1665,N_1114);
nor U2074 (N_2074,In_415,N_1582);
or U2075 (N_2075,In_3445,In_899);
or U2076 (N_2076,In_3416,N_1821);
xnor U2077 (N_2077,In_696,In_1900);
xnor U2078 (N_2078,N_923,N_1065);
nor U2079 (N_2079,In_3870,N_1585);
or U2080 (N_2080,N_1417,N_1933);
and U2081 (N_2081,In_4426,N_635);
or U2082 (N_2082,In_2464,N_1096);
xor U2083 (N_2083,In_1785,N_866);
nor U2084 (N_2084,N_1895,N_1789);
and U2085 (N_2085,In_885,In_2327);
xor U2086 (N_2086,In_2253,N_1514);
nand U2087 (N_2087,In_3674,In_879);
and U2088 (N_2088,In_3220,N_1979);
nor U2089 (N_2089,In_1613,In_337);
xnor U2090 (N_2090,In_1033,N_1827);
nand U2091 (N_2091,N_1923,N_1804);
xnor U2092 (N_2092,N_911,In_3075);
nand U2093 (N_2093,N_1784,N_1620);
nor U2094 (N_2094,N_1761,N_1372);
or U2095 (N_2095,In_527,In_1993);
nand U2096 (N_2096,N_1515,In_2762);
nand U2097 (N_2097,In_3299,N_1965);
and U2098 (N_2098,N_708,N_535);
nor U2099 (N_2099,N_1522,N_1815);
and U2100 (N_2100,N_591,In_2008);
and U2101 (N_2101,In_4432,In_4810);
nor U2102 (N_2102,In_720,N_1403);
xor U2103 (N_2103,N_211,N_112);
xor U2104 (N_2104,N_1675,In_2545);
nand U2105 (N_2105,N_1796,In_3306);
xnor U2106 (N_2106,In_3354,In_2862);
nand U2107 (N_2107,N_1377,In_1048);
and U2108 (N_2108,In_584,In_18);
xnor U2109 (N_2109,N_1558,N_688);
and U2110 (N_2110,In_2271,In_1813);
nor U2111 (N_2111,In_1109,In_287);
or U2112 (N_2112,In_692,In_500);
xnor U2113 (N_2113,In_4213,N_1140);
or U2114 (N_2114,N_1313,N_1357);
xnor U2115 (N_2115,In_1587,In_2422);
xnor U2116 (N_2116,N_1411,In_4948);
or U2117 (N_2117,N_1544,N_1853);
nand U2118 (N_2118,In_1515,N_904);
xor U2119 (N_2119,N_100,In_791);
nand U2120 (N_2120,N_1727,In_1123);
nand U2121 (N_2121,N_1894,In_2184);
or U2122 (N_2122,N_1688,N_1877);
nand U2123 (N_2123,In_332,N_1975);
nor U2124 (N_2124,In_622,N_1307);
or U2125 (N_2125,N_1429,In_3677);
or U2126 (N_2126,In_2066,In_592);
nor U2127 (N_2127,In_3167,In_539);
nor U2128 (N_2128,In_170,In_2669);
and U2129 (N_2129,N_283,In_1716);
nor U2130 (N_2130,N_1101,N_700);
xor U2131 (N_2131,In_2860,N_1126);
nand U2132 (N_2132,In_1454,In_3597);
nor U2133 (N_2133,N_139,N_356);
nand U2134 (N_2134,In_3585,N_559);
nand U2135 (N_2135,N_11,In_1415);
and U2136 (N_2136,N_663,N_150);
nand U2137 (N_2137,N_357,In_682);
or U2138 (N_2138,N_1918,N_1342);
or U2139 (N_2139,In_861,N_1160);
or U2140 (N_2140,In_2829,In_247);
xor U2141 (N_2141,N_571,In_3761);
xnor U2142 (N_2142,N_1667,In_4265);
xnor U2143 (N_2143,N_1409,In_2210);
or U2144 (N_2144,N_1568,N_1997);
xnor U2145 (N_2145,In_762,In_3453);
nand U2146 (N_2146,N_777,N_956);
and U2147 (N_2147,N_453,In_1524);
or U2148 (N_2148,In_3311,In_168);
xnor U2149 (N_2149,N_1605,N_548);
xor U2150 (N_2150,In_611,In_2483);
or U2151 (N_2151,N_1931,N_1179);
and U2152 (N_2152,N_61,In_1472);
xnor U2153 (N_2153,N_2,In_4390);
xnor U2154 (N_2154,N_1596,N_1343);
xnor U2155 (N_2155,In_4292,In_144);
nor U2156 (N_2156,N_1314,In_3237);
and U2157 (N_2157,In_4019,In_1162);
xor U2158 (N_2158,N_524,In_4075);
nor U2159 (N_2159,In_277,In_4149);
nand U2160 (N_2160,In_545,In_2383);
and U2161 (N_2161,N_1472,In_3874);
xnor U2162 (N_2162,N_729,In_3273);
or U2163 (N_2163,In_21,In_680);
xor U2164 (N_2164,In_112,In_1360);
and U2165 (N_2165,In_1133,N_1991);
nor U2166 (N_2166,In_4837,In_3836);
xor U2167 (N_2167,N_1276,In_4996);
or U2168 (N_2168,In_669,N_788);
or U2169 (N_2169,N_1910,In_2833);
xor U2170 (N_2170,In_3450,In_3049);
xor U2171 (N_2171,N_1134,In_4899);
nor U2172 (N_2172,N_497,N_1878);
or U2173 (N_2173,N_979,In_2664);
or U2174 (N_2174,In_1603,In_3947);
or U2175 (N_2175,In_2207,N_573);
nor U2176 (N_2176,N_1046,N_1673);
nand U2177 (N_2177,In_1419,In_36);
xnor U2178 (N_2178,In_3591,In_4009);
xnor U2179 (N_2179,N_1430,In_4958);
nand U2180 (N_2180,N_1136,In_4228);
and U2181 (N_2181,N_576,In_1990);
xnor U2182 (N_2182,In_1985,In_369);
nand U2183 (N_2183,In_1927,In_3540);
xor U2184 (N_2184,N_1287,N_13);
or U2185 (N_2185,N_407,N_409);
or U2186 (N_2186,In_2111,In_3730);
xor U2187 (N_2187,In_1621,In_2924);
or U2188 (N_2188,N_958,N_1494);
nor U2189 (N_2189,In_346,In_4622);
xor U2190 (N_2190,In_4373,N_1150);
nor U2191 (N_2191,In_339,N_1703);
nand U2192 (N_2192,In_2148,N_575);
nor U2193 (N_2193,In_3349,In_2341);
xnor U2194 (N_2194,In_3435,In_56);
nand U2195 (N_2195,N_749,In_2309);
nor U2196 (N_2196,In_3813,In_4000);
nor U2197 (N_2197,In_3203,In_2479);
xnor U2198 (N_2198,In_2680,N_1733);
or U2199 (N_2199,N_1772,N_1759);
or U2200 (N_2200,N_1950,In_4372);
or U2201 (N_2201,N_536,In_4128);
nor U2202 (N_2202,N_85,In_4261);
xor U2203 (N_2203,N_1509,N_1581);
nand U2204 (N_2204,N_1078,N_944);
and U2205 (N_2205,In_1135,N_681);
nand U2206 (N_2206,N_1787,In_3533);
xnor U2207 (N_2207,N_567,In_835);
nor U2208 (N_2208,N_38,N_742);
nor U2209 (N_2209,In_3521,In_3899);
nor U2210 (N_2210,In_839,N_466);
xnor U2211 (N_2211,N_1056,N_1816);
and U2212 (N_2212,In_4100,In_4398);
nor U2213 (N_2213,In_1507,In_4655);
or U2214 (N_2214,In_3792,In_3511);
or U2215 (N_2215,In_502,In_1065);
nor U2216 (N_2216,In_3944,In_1165);
xnor U2217 (N_2217,In_3190,In_882);
xnor U2218 (N_2218,In_4453,N_1870);
or U2219 (N_2219,In_4861,N_330);
nand U2220 (N_2220,N_1109,In_1174);
nand U2221 (N_2221,N_1819,In_2754);
nand U2222 (N_2222,In_2162,N_1375);
xnor U2223 (N_2223,N_621,N_1448);
nor U2224 (N_2224,In_548,In_1306);
nor U2225 (N_2225,N_1664,In_1188);
or U2226 (N_2226,In_2322,In_3074);
xor U2227 (N_2227,N_484,In_1596);
xnor U2228 (N_2228,In_3497,In_437);
xor U2229 (N_2229,N_1461,In_4397);
nor U2230 (N_2230,In_3054,In_2739);
nor U2231 (N_2231,In_3789,In_2200);
nor U2232 (N_2232,In_4071,In_1237);
and U2233 (N_2233,N_935,In_2979);
nor U2234 (N_2234,In_4340,N_1000);
nand U2235 (N_2235,N_265,N_1648);
nand U2236 (N_2236,In_405,In_4272);
nor U2237 (N_2237,N_1844,N_1122);
xor U2238 (N_2238,N_1905,In_847);
nor U2239 (N_2239,N_1185,N_1017);
and U2240 (N_2240,N_813,N_1964);
or U2241 (N_2241,In_2251,In_2610);
nor U2242 (N_2242,In_4172,In_3630);
nor U2243 (N_2243,N_1495,In_725);
and U2244 (N_2244,N_215,In_4592);
xor U2245 (N_2245,In_3801,N_761);
xor U2246 (N_2246,In_202,In_846);
and U2247 (N_2247,N_1252,In_1248);
nor U2248 (N_2248,In_3782,In_4731);
and U2249 (N_2249,In_3667,In_3891);
xor U2250 (N_2250,In_3032,In_4139);
nor U2251 (N_2251,In_2307,N_1713);
nor U2252 (N_2252,In_3358,In_3189);
or U2253 (N_2253,In_2049,In_156);
and U2254 (N_2254,In_2071,N_998);
and U2255 (N_2255,In_2964,N_488);
xnor U2256 (N_2256,N_1794,N_1348);
xnor U2257 (N_2257,N_1295,N_585);
nor U2258 (N_2258,In_3238,In_751);
nand U2259 (N_2259,N_969,In_3394);
nor U2260 (N_2260,In_2587,N_578);
nand U2261 (N_2261,In_715,In_593);
and U2262 (N_2262,In_8,N_1981);
xor U2263 (N_2263,In_4629,In_1925);
xor U2264 (N_2264,In_1200,N_1198);
nor U2265 (N_2265,N_697,N_1436);
nor U2266 (N_2266,In_182,N_251);
nor U2267 (N_2267,In_3633,In_1629);
and U2268 (N_2268,N_509,In_396);
nand U2269 (N_2269,N_116,In_3601);
nand U2270 (N_2270,In_1334,In_4676);
nor U2271 (N_2271,N_727,In_2436);
nand U2272 (N_2272,N_1683,In_2001);
xnor U2273 (N_2273,N_1584,N_780);
nand U2274 (N_2274,In_2508,In_1722);
or U2275 (N_2275,N_1384,N_1690);
or U2276 (N_2276,In_3388,In_1915);
nor U2277 (N_2277,In_4083,N_1630);
xor U2278 (N_2278,N_926,In_4210);
xor U2279 (N_2279,N_403,In_1401);
nor U2280 (N_2280,In_1341,In_1081);
nor U2281 (N_2281,In_441,N_1028);
and U2282 (N_2282,N_1175,N_711);
and U2283 (N_2283,In_826,In_4550);
or U2284 (N_2284,N_1723,In_586);
nand U2285 (N_2285,N_1833,In_2291);
nor U2286 (N_2286,N_1601,In_2413);
and U2287 (N_2287,N_1487,N_1315);
or U2288 (N_2288,In_1839,N_262);
nand U2289 (N_2289,N_995,In_4879);
nand U2290 (N_2290,N_1592,In_2794);
nand U2291 (N_2291,In_345,In_1578);
nor U2292 (N_2292,In_1553,In_176);
xnor U2293 (N_2293,N_229,In_1908);
or U2294 (N_2294,N_1037,In_4875);
and U2295 (N_2295,N_1996,N_1465);
nand U2296 (N_2296,In_1278,N_1376);
nor U2297 (N_2297,In_4916,In_3863);
xnor U2298 (N_2298,In_3422,N_1240);
or U2299 (N_2299,N_959,In_164);
nor U2300 (N_2300,In_3479,N_1771);
xnor U2301 (N_2301,In_4101,N_1319);
xnor U2302 (N_2302,In_1968,In_4378);
xnor U2303 (N_2303,In_1682,N_1685);
and U2304 (N_2304,In_1387,N_1104);
and U2305 (N_2305,N_1670,In_1693);
xnor U2306 (N_2306,N_775,N_1071);
or U2307 (N_2307,In_2022,In_4081);
and U2308 (N_2308,In_4538,In_62);
nand U2309 (N_2309,N_1753,In_1223);
xor U2310 (N_2310,N_397,In_67);
and U2311 (N_2311,In_1668,In_3617);
or U2312 (N_2312,N_1556,N_887);
xor U2313 (N_2313,In_667,N_1682);
nor U2314 (N_2314,N_1891,N_1414);
or U2315 (N_2315,In_4568,In_2306);
nand U2316 (N_2316,N_963,In_4994);
nor U2317 (N_2317,In_3543,N_990);
or U2318 (N_2318,In_2555,In_4484);
nand U2319 (N_2319,In_3118,In_1311);
or U2320 (N_2320,N_652,In_1873);
xnor U2321 (N_2321,N_1043,N_1500);
nand U2322 (N_2322,N_1290,N_391);
xnor U2323 (N_2323,N_348,N_203);
nor U2324 (N_2324,In_3100,In_3008);
nand U2325 (N_2325,N_1720,N_1346);
and U2326 (N_2326,In_1725,In_3241);
nand U2327 (N_2327,In_422,N_1052);
or U2328 (N_2328,In_4561,In_2112);
or U2329 (N_2329,N_795,N_1453);
xor U2330 (N_2330,In_4242,In_187);
nor U2331 (N_2331,N_1005,N_1441);
and U2332 (N_2332,In_3009,In_848);
and U2333 (N_2333,N_1069,In_3125);
xor U2334 (N_2334,In_362,N_217);
and U2335 (N_2335,N_1773,N_1294);
and U2336 (N_2336,N_803,N_1945);
nor U2337 (N_2337,N_1949,In_2262);
or U2338 (N_2338,In_1438,In_4804);
or U2339 (N_2339,N_1824,N_1712);
or U2340 (N_2340,N_628,In_2989);
nand U2341 (N_2341,In_2429,In_2369);
and U2342 (N_2342,N_1209,N_1151);
or U2343 (N_2343,N_198,N_1978);
or U2344 (N_2344,N_1219,N_1864);
and U2345 (N_2345,N_347,In_2618);
and U2346 (N_2346,N_1939,In_875);
nor U2347 (N_2347,In_2697,In_1184);
nor U2348 (N_2348,In_3362,N_1484);
xor U2349 (N_2349,In_2297,N_37);
nand U2350 (N_2350,In_2228,In_2227);
xor U2351 (N_2351,N_1334,N_1587);
nor U2352 (N_2352,In_1323,In_3892);
or U2353 (N_2353,In_3631,N_871);
nor U2354 (N_2354,In_2759,In_4499);
nor U2355 (N_2355,In_363,In_1743);
nand U2356 (N_2356,In_901,In_1855);
nand U2357 (N_2357,In_3470,In_1207);
nor U2358 (N_2358,In_53,N_1218);
and U2359 (N_2359,N_517,In_567);
xor U2360 (N_2360,In_2665,In_4738);
nand U2361 (N_2361,In_1686,In_3922);
nor U2362 (N_2362,In_4812,N_1248);
nand U2363 (N_2363,N_1744,N_1999);
and U2364 (N_2364,N_1742,In_4790);
and U2365 (N_2365,N_957,N_1721);
or U2366 (N_2366,In_1029,N_1378);
or U2367 (N_2367,In_4721,In_1073);
and U2368 (N_2368,In_629,N_725);
nand U2369 (N_2369,In_4976,N_863);
nor U2370 (N_2370,In_2787,N_1711);
xnor U2371 (N_2371,In_3685,In_271);
xnor U2372 (N_2372,N_1363,In_1823);
and U2373 (N_2373,In_240,N_1597);
nand U2374 (N_2374,In_1342,In_2592);
nand U2375 (N_2375,N_1088,N_1518);
xnor U2376 (N_2376,N_1668,In_198);
xor U2377 (N_2377,In_449,N_1850);
xnor U2378 (N_2378,In_1095,In_4874);
nor U2379 (N_2379,N_1908,In_249);
xor U2380 (N_2380,N_258,N_1442);
nand U2381 (N_2381,N_1001,N_1801);
nor U2382 (N_2382,N_474,In_1820);
nand U2383 (N_2383,In_603,N_593);
nand U2384 (N_2384,In_4682,In_3124);
nor U2385 (N_2385,N_121,N_175);
and U2386 (N_2386,N_845,N_1452);
nand U2387 (N_2387,In_3604,In_2600);
nor U2388 (N_2388,N_1880,In_1483);
xor U2389 (N_2389,N_1956,In_3342);
xor U2390 (N_2390,N_1861,N_12);
nor U2391 (N_2391,In_4287,N_1038);
nor U2392 (N_2392,In_499,In_3950);
and U2393 (N_2393,N_46,N_388);
nor U2394 (N_2394,In_3844,N_390);
nand U2395 (N_2395,In_3283,In_3682);
xor U2396 (N_2396,In_1205,N_1511);
nor U2397 (N_2397,In_1733,N_1117);
nand U2398 (N_2398,In_1566,In_3048);
nor U2399 (N_2399,N_1013,In_1902);
nor U2400 (N_2400,N_542,N_1271);
nand U2401 (N_2401,N_432,In_1031);
nor U2402 (N_2402,In_2160,N_505);
and U2403 (N_2403,N_1233,In_909);
or U2404 (N_2404,In_672,N_787);
nand U2405 (N_2405,In_3200,N_846);
and U2406 (N_2406,In_3683,In_4558);
nor U2407 (N_2407,In_376,In_1673);
and U2408 (N_2408,In_3065,N_906);
nor U2409 (N_2409,In_1132,N_1915);
xnor U2410 (N_2410,N_1885,N_1211);
and U2411 (N_2411,In_1446,In_4762);
or U2412 (N_2412,N_1390,In_753);
or U2413 (N_2413,In_1247,In_455);
or U2414 (N_2414,N_34,In_1440);
xnor U2415 (N_2415,In_1604,N_739);
nor U2416 (N_2416,In_2874,N_1657);
xnor U2417 (N_2417,N_1217,In_4662);
xor U2418 (N_2418,In_1922,In_4146);
xor U2419 (N_2419,N_166,N_1913);
xnor U2420 (N_2420,N_1431,N_1681);
xor U2421 (N_2421,N_1637,In_3855);
and U2422 (N_2422,In_3229,N_1843);
xor U2423 (N_2423,N_435,In_2602);
or U2424 (N_2424,In_3130,N_938);
nand U2425 (N_2425,In_2393,N_1311);
xnor U2426 (N_2426,In_1012,N_1040);
xor U2427 (N_2427,In_73,In_3326);
nor U2428 (N_2428,In_2505,In_965);
xnor U2429 (N_2429,In_4508,In_1338);
nor U2430 (N_2430,In_4199,N_686);
and U2431 (N_2431,N_1957,N_1579);
nor U2432 (N_2432,In_4260,N_1612);
nor U2433 (N_2433,In_2846,N_204);
or U2434 (N_2434,In_1593,N_895);
nor U2435 (N_2435,In_4103,N_209);
and U2436 (N_2436,In_843,In_555);
xnor U2437 (N_2437,In_2336,In_2549);
xnor U2438 (N_2438,In_4807,In_2717);
nor U2439 (N_2439,In_2890,N_595);
and U2440 (N_2440,In_4349,N_152);
nand U2441 (N_2441,N_1476,In_3703);
nor U2442 (N_2442,N_151,N_143);
or U2443 (N_2443,In_4745,In_61);
or U2444 (N_2444,N_1458,In_1736);
xnor U2445 (N_2445,In_3529,In_107);
xor U2446 (N_2446,In_2548,In_2998);
xor U2447 (N_2447,In_675,In_4439);
and U2448 (N_2448,In_543,In_2845);
nor U2449 (N_2449,In_730,In_2020);
or U2450 (N_2450,In_3431,N_613);
nor U2451 (N_2451,In_4619,In_2841);
nand U2452 (N_2452,In_1080,N_763);
nor U2453 (N_2453,N_831,In_3274);
nand U2454 (N_2454,N_869,In_2678);
or U2455 (N_2455,N_1099,N_1473);
xor U2456 (N_2456,N_698,In_738);
nor U2457 (N_2457,N_917,N_720);
and U2458 (N_2458,In_3903,In_1816);
nor U2459 (N_2459,N_525,N_1676);
and U2460 (N_2460,In_236,In_1723);
or U2461 (N_2461,In_4923,N_253);
or U2462 (N_2462,N_1186,N_588);
and U2463 (N_2463,N_970,In_1487);
nand U2464 (N_2464,In_2965,In_1750);
nand U2465 (N_2465,N_1480,N_308);
nand U2466 (N_2466,N_318,N_929);
nor U2467 (N_2467,N_560,N_1199);
nor U2468 (N_2468,N_1444,N_1526);
or U2469 (N_2469,In_2771,In_1263);
nand U2470 (N_2470,In_438,In_4724);
nor U2471 (N_2471,In_3981,In_1999);
and U2472 (N_2472,In_728,In_2405);
xor U2473 (N_2473,N_1562,N_286);
xnor U2474 (N_2474,N_1520,N_1366);
nor U2475 (N_2475,N_1874,In_4277);
nor U2476 (N_2476,N_1756,In_3180);
and U2477 (N_2477,In_3738,N_1224);
or U2478 (N_2478,N_987,N_1573);
xor U2479 (N_2479,N_753,In_4860);
nor U2480 (N_2480,In_5,N_1741);
nor U2481 (N_2481,N_1566,In_2199);
nor U2482 (N_2482,In_4436,In_2349);
nand U2483 (N_2483,In_4307,N_1595);
and U2484 (N_2484,N_1651,N_1828);
nand U2485 (N_2485,In_130,N_733);
or U2486 (N_2486,N_1732,N_1752);
xor U2487 (N_2487,N_1661,In_4417);
nor U2488 (N_2488,N_417,N_1848);
nand U2489 (N_2489,N_1481,N_902);
and U2490 (N_2490,In_1930,In_4112);
and U2491 (N_2491,N_601,N_1572);
or U2492 (N_2492,In_830,In_566);
and U2493 (N_2493,N_328,N_1867);
or U2494 (N_2494,In_2041,In_88);
or U2495 (N_2495,In_1102,N_1505);
and U2496 (N_2496,In_3909,N_692);
nor U2497 (N_2497,N_738,N_701);
or U2498 (N_2498,N_1026,In_4446);
nand U2499 (N_2499,In_1913,N_597);
xor U2500 (N_2500,N_2380,N_2091);
xor U2501 (N_2501,N_2218,In_3070);
or U2502 (N_2502,In_3750,N_1972);
or U2503 (N_2503,N_2493,N_1671);
and U2504 (N_2504,In_2691,N_1858);
xnor U2505 (N_2505,N_892,N_2174);
nor U2506 (N_2506,In_4973,In_2256);
xor U2507 (N_2507,N_809,In_3018);
or U2508 (N_2508,In_571,In_704);
xor U2509 (N_2509,N_1875,In_865);
nand U2510 (N_2510,In_2141,In_732);
and U2511 (N_2511,In_106,In_1014);
and U2512 (N_2512,N_2242,N_1947);
nor U2513 (N_2513,N_1537,In_1072);
or U2514 (N_2514,N_1943,In_414);
or U2515 (N_2515,In_3820,N_2093);
xnor U2516 (N_2516,N_1696,N_1184);
nand U2517 (N_2517,N_2187,In_504);
and U2518 (N_2518,In_2426,In_4316);
or U2519 (N_2519,In_4939,N_1619);
nor U2520 (N_2520,In_1147,N_1707);
and U2521 (N_2521,N_1901,In_4271);
nor U2522 (N_2522,In_97,N_922);
nor U2523 (N_2523,In_922,In_2512);
nor U2524 (N_2524,In_2192,N_1812);
nand U2525 (N_2525,In_561,In_3141);
nor U2526 (N_2526,In_494,In_4635);
or U2527 (N_2527,N_703,In_1428);
xor U2528 (N_2528,N_2128,N_2280);
xor U2529 (N_2529,In_1624,N_2312);
and U2530 (N_2530,In_1486,N_1882);
nand U2531 (N_2531,N_2463,N_1529);
and U2532 (N_2532,In_2284,In_3524);
nor U2533 (N_2533,N_2176,In_645);
and U2534 (N_2534,In_4395,N_2193);
and U2535 (N_2535,In_4528,N_1745);
nor U2536 (N_2536,N_2215,N_1578);
nand U2537 (N_2537,In_124,N_1259);
nand U2538 (N_2538,In_1287,In_2728);
nor U2539 (N_2539,In_776,In_515);
and U2540 (N_2540,N_2374,N_1896);
or U2541 (N_2541,In_2274,In_2952);
and U2542 (N_2542,N_2346,N_2070);
nand U2543 (N_2543,N_1600,N_395);
nor U2544 (N_2544,N_974,In_1392);
nand U2545 (N_2545,In_983,N_2278);
nand U2546 (N_2546,N_2137,In_4618);
xor U2547 (N_2547,N_2240,N_2032);
nor U2548 (N_2548,In_4705,N_1655);
nand U2549 (N_2549,In_768,In_2290);
nor U2550 (N_2550,In_4709,N_2205);
nor U2551 (N_2551,N_2260,N_2490);
and U2552 (N_2552,N_2298,N_2394);
and U2553 (N_2553,N_1541,In_1405);
or U2554 (N_2554,N_864,N_2057);
nor U2555 (N_2555,N_610,In_4311);
or U2556 (N_2556,N_1284,In_3741);
or U2557 (N_2557,In_4583,N_2387);
xnor U2558 (N_2558,N_2049,In_2645);
xor U2559 (N_2559,In_4033,N_566);
or U2560 (N_2560,N_660,In_4552);
nor U2561 (N_2561,N_1012,N_2173);
and U2562 (N_2562,N_1936,N_2252);
nor U2563 (N_2563,In_1017,In_1040);
and U2564 (N_2564,In_4479,N_53);
nand U2565 (N_2565,N_292,N_2189);
and U2566 (N_2566,In_2901,In_3925);
nand U2567 (N_2567,In_1996,N_1766);
nor U2568 (N_2568,N_2063,In_1316);
or U2569 (N_2569,N_2067,In_167);
xnor U2570 (N_2570,In_1983,In_209);
nand U2571 (N_2571,In_1639,N_1726);
xnor U2572 (N_2572,N_1205,N_2229);
xor U2573 (N_2573,In_3774,In_3249);
or U2574 (N_2574,In_1161,In_1608);
xor U2575 (N_2575,N_2248,In_962);
or U2576 (N_2576,N_716,In_4379);
nor U2577 (N_2577,N_1075,In_774);
nor U2578 (N_2578,In_2330,In_2630);
nand U2579 (N_2579,N_1015,In_2761);
xor U2580 (N_2580,In_3,N_2324);
nor U2581 (N_2581,N_1469,In_2514);
or U2582 (N_2582,N_1246,In_419);
or U2583 (N_2583,N_2207,In_2921);
nand U2584 (N_2584,N_1714,In_1117);
or U2585 (N_2585,N_406,N_2097);
nor U2586 (N_2586,N_823,In_465);
nor U2587 (N_2587,In_108,In_2528);
nor U2588 (N_2588,In_1724,N_1841);
and U2589 (N_2589,In_2342,N_2227);
and U2590 (N_2590,N_2078,N_165);
nor U2591 (N_2591,In_2944,In_707);
nand U2592 (N_2592,In_4781,N_1770);
nand U2593 (N_2593,N_1195,In_472);
or U2594 (N_2594,N_1030,N_797);
or U2595 (N_2595,N_1310,In_4752);
nand U2596 (N_2596,In_3676,In_2201);
xnor U2597 (N_2597,In_4459,In_2143);
and U2598 (N_2598,N_656,N_180);
and U2599 (N_2599,N_2188,N_1641);
and U2600 (N_2600,N_1320,In_3119);
nor U2601 (N_2601,N_1591,N_2133);
xor U2602 (N_2602,N_51,In_3951);
or U2603 (N_2603,In_2272,N_2251);
or U2604 (N_2604,N_331,N_1157);
nand U2605 (N_2605,N_1168,N_285);
nor U2606 (N_2606,N_2041,N_1545);
xnor U2607 (N_2607,N_1645,N_1032);
and U2608 (N_2608,N_120,In_752);
nor U2609 (N_2609,In_3369,In_3893);
nand U2610 (N_2610,N_1846,In_4030);
xnor U2611 (N_2611,N_1847,N_1074);
xor U2612 (N_2612,In_2154,N_1059);
xor U2613 (N_2613,N_1911,N_1340);
xor U2614 (N_2614,In_2591,N_1178);
nor U2615 (N_2615,N_1020,N_2117);
xor U2616 (N_2616,N_1538,N_1798);
and U2617 (N_2617,N_1762,N_1737);
xor U2618 (N_2618,N_1102,N_1115);
or U2619 (N_2619,In_2090,N_1135);
and U2620 (N_2620,N_2022,N_1836);
or U2621 (N_2621,In_3361,N_2443);
nand U2622 (N_2622,N_2023,N_2393);
nand U2623 (N_2623,In_3053,N_2226);
and U2624 (N_2624,N_2196,N_2337);
and U2625 (N_2625,N_2124,N_2050);
nand U2626 (N_2626,N_2429,N_1702);
or U2627 (N_2627,N_1539,N_18);
or U2628 (N_2628,In_4560,N_1223);
nor U2629 (N_2629,N_1842,In_2662);
or U2630 (N_2630,N_2462,N_195);
and U2631 (N_2631,N_2291,N_2434);
and U2632 (N_2632,N_1973,N_2367);
and U2633 (N_2633,In_729,In_1362);
or U2634 (N_2634,N_2234,N_746);
nor U2635 (N_2635,In_950,In_4365);
nand U2636 (N_2636,In_1581,N_1089);
and U2637 (N_2637,N_82,N_647);
xor U2638 (N_2638,N_2481,In_1319);
nand U2639 (N_2639,N_1018,N_2164);
xnor U2640 (N_2640,In_2050,N_1919);
xor U2641 (N_2641,N_2457,In_4904);
nor U2642 (N_2642,N_2142,In_2735);
nand U2643 (N_2643,In_3245,N_464);
nand U2644 (N_2644,N_1298,In_32);
xnor U2645 (N_2645,N_94,N_1951);
xor U2646 (N_2646,In_4430,N_2114);
and U2647 (N_2647,N_1230,N_2213);
or U2648 (N_2648,In_3391,N_1245);
nand U2649 (N_2649,In_262,N_1750);
xnor U2650 (N_2650,In_213,In_3016);
and U2651 (N_2651,In_4548,N_1719);
or U2652 (N_2652,N_1410,N_1507);
nand U2653 (N_2653,In_4118,N_2175);
nor U2654 (N_2654,In_605,In_1281);
and U2655 (N_2655,N_1912,In_2659);
xor U2656 (N_2656,N_1143,N_657);
or U2657 (N_2657,In_1286,N_1475);
or U2658 (N_2658,N_1599,N_2012);
nand U2659 (N_2659,In_2899,N_724);
or U2660 (N_2660,N_2224,In_132);
or U2661 (N_2661,In_284,In_814);
nand U2662 (N_2662,N_1791,N_448);
nor U2663 (N_2663,N_975,N_744);
and U2664 (N_2664,In_3628,N_1263);
nor U2665 (N_2665,In_4672,N_190);
xor U2666 (N_2666,N_886,In_3383);
nor U2667 (N_2667,In_1443,In_4686);
nand U2668 (N_2668,N_1897,N_1288);
or U2669 (N_2669,In_4301,In_1166);
nand U2670 (N_2670,N_1543,In_2877);
or U2671 (N_2671,N_1451,In_3341);
and U2672 (N_2672,N_378,N_2305);
nor U2673 (N_2673,In_174,In_2500);
nand U2674 (N_2674,N_2344,N_1715);
xor U2675 (N_2675,In_1972,N_2343);
nand U2676 (N_2676,In_2329,In_802);
and U2677 (N_2677,N_2151,In_2577);
xor U2678 (N_2678,N_1330,N_2382);
and U2679 (N_2679,N_2345,In_4529);
xor U2680 (N_2680,In_3623,In_4482);
nor U2681 (N_2681,In_2719,N_2211);
xnor U2682 (N_2682,N_2220,N_2470);
and U2683 (N_2683,N_1380,In_2074);
nor U2684 (N_2684,In_714,N_1517);
xor U2685 (N_2685,N_550,In_532);
and U2686 (N_2686,N_633,N_2058);
xnor U2687 (N_2687,N_1650,In_626);
or U2688 (N_2688,N_1704,N_1660);
or U2689 (N_2689,N_2399,In_4290);
nand U2690 (N_2690,In_4757,N_370);
nand U2691 (N_2691,N_2292,N_737);
nand U2692 (N_2692,In_4151,N_740);
and U2693 (N_2693,N_1493,In_4892);
and U2694 (N_2694,In_336,In_3493);
or U2695 (N_2695,In_1944,N_1623);
nand U2696 (N_2696,In_699,N_425);
nor U2697 (N_2697,N_2182,N_1328);
and U2698 (N_2698,N_1680,In_152);
or U2699 (N_2699,In_1363,N_172);
and U2700 (N_2700,In_2791,N_978);
and U2701 (N_2701,In_3081,N_1004);
or U2702 (N_2702,In_551,N_2168);
nor U2703 (N_2703,In_1519,N_2009);
nand U2704 (N_2704,In_1153,N_2007);
or U2705 (N_2705,In_1230,N_2149);
nand U2706 (N_2706,In_2385,N_1488);
or U2707 (N_2707,In_393,N_490);
or U2708 (N_2708,In_1210,In_681);
nand U2709 (N_2709,In_2990,N_859);
nand U2710 (N_2710,N_1834,N_1649);
and U2711 (N_2711,In_868,N_50);
xnor U2712 (N_2712,N_1269,In_4688);
nor U2713 (N_2713,In_2325,In_1055);
or U2714 (N_2714,N_1958,In_3884);
or U2715 (N_2715,In_165,N_170);
nand U2716 (N_2716,N_880,N_726);
and U2717 (N_2717,N_604,N_2243);
and U2718 (N_2718,In_2800,In_4491);
nand U2719 (N_2719,N_1174,In_3195);
xor U2720 (N_2720,In_4856,N_2018);
nand U2721 (N_2721,In_3748,In_1520);
or U2722 (N_2722,N_1967,N_167);
xnor U2723 (N_2723,In_157,N_2362);
xnor U2724 (N_2724,In_3791,N_2126);
or U2725 (N_2725,In_2484,In_3698);
and U2726 (N_2726,N_1722,N_2452);
xor U2727 (N_2727,In_1136,In_1861);
nand U2728 (N_2728,In_281,In_1068);
nand U2729 (N_2729,In_1150,N_1610);
nor U2730 (N_2730,N_1204,In_3225);
nand U2731 (N_2731,N_1490,N_2025);
and U2732 (N_2732,N_2237,In_4474);
nor U2733 (N_2733,N_834,N_2144);
nor U2734 (N_2734,N_1608,In_4871);
or U2735 (N_2735,In_4540,N_1024);
nor U2736 (N_2736,In_4641,N_2424);
nor U2737 (N_2737,N_2301,In_4783);
nor U2738 (N_2738,In_3146,N_2316);
xor U2739 (N_2739,N_1144,In_128);
nor U2740 (N_2740,N_1446,N_2271);
nor U2741 (N_2741,N_1962,In_63);
xnor U2742 (N_2742,In_387,N_2307);
or U2743 (N_2743,In_2442,In_4902);
and U2744 (N_2744,N_1588,N_1983);
xnor U2745 (N_2745,In_60,In_1870);
nand U2746 (N_2746,N_2360,N_2254);
xor U2747 (N_2747,N_2136,N_2386);
and U2748 (N_2748,In_793,N_1839);
nand U2749 (N_2749,In_2765,N_2303);
and U2750 (N_2750,N_811,N_2259);
xnor U2751 (N_2751,In_2446,N_2486);
nand U2752 (N_2752,In_3022,In_4133);
nor U2753 (N_2753,N_1042,In_125);
nand U2754 (N_2754,In_2164,In_3647);
and U2755 (N_2755,In_818,N_1755);
nor U2756 (N_2756,In_821,N_2270);
xor U2757 (N_2757,N_1316,N_2069);
nor U2758 (N_2758,In_3329,N_360);
or U2759 (N_2759,N_1247,In_3295);
nand U2760 (N_2760,N_2160,N_1009);
or U2761 (N_2761,In_1841,N_1963);
or U2762 (N_2762,N_2236,In_1806);
xor U2763 (N_2763,In_2386,In_3831);
or U2764 (N_2764,N_182,In_218);
nor U2765 (N_2765,N_2198,N_2066);
nand U2766 (N_2766,N_2036,N_2406);
xnor U2767 (N_2767,In_3154,N_1280);
xor U2768 (N_2768,In_3011,In_2129);
and U2769 (N_2769,N_2427,In_541);
nand U2770 (N_2770,In_1347,N_999);
xor U2771 (N_2771,N_1561,N_2170);
nor U2772 (N_2772,In_1862,N_97);
nand U2773 (N_2773,N_939,N_1832);
nor U2774 (N_2774,In_642,N_1306);
nor U2775 (N_2775,In_4737,N_1076);
nor U2776 (N_2776,In_3272,In_1674);
and U2777 (N_2777,In_4041,N_985);
nand U2778 (N_2778,In_4269,In_425);
nand U2779 (N_2779,N_1395,In_3967);
and U2780 (N_2780,N_1527,N_2461);
nand U2781 (N_2781,In_4362,N_1304);
and U2782 (N_2782,N_1362,N_173);
xor U2783 (N_2783,N_1392,N_1795);
nor U2784 (N_2784,N_2001,N_1729);
and U2785 (N_2785,In_4541,N_1575);
nor U2786 (N_2786,N_1808,N_2059);
nor U2787 (N_2787,N_2274,In_3768);
or U2788 (N_2788,In_3102,N_627);
nor U2789 (N_2789,N_839,N_2055);
or U2790 (N_2790,In_623,N_1697);
or U2791 (N_2791,In_1615,In_934);
nor U2792 (N_2792,In_3407,In_1791);
nand U2793 (N_2793,In_3000,In_3079);
nand U2794 (N_2794,In_79,N_1341);
or U2795 (N_2795,In_4816,In_4068);
nand U2796 (N_2796,In_1297,In_1077);
or U2797 (N_2797,In_3310,N_1139);
or U2798 (N_2798,N_1010,N_171);
and U2799 (N_2799,N_574,N_1305);
and U2800 (N_2800,In_2789,N_1238);
xnor U2801 (N_2801,N_2300,N_1862);
or U2802 (N_2802,In_1858,N_1132);
xor U2803 (N_2803,N_968,N_90);
or U2804 (N_2804,N_666,In_2682);
xnor U2805 (N_2805,N_1213,N_1105);
or U2806 (N_2806,N_1872,In_1891);
xor U2807 (N_2807,In_1732,N_2389);
and U2808 (N_2808,In_3469,In_910);
and U2809 (N_2809,In_2356,In_1986);
and U2810 (N_2810,N_1583,N_1614);
or U2811 (N_2811,N_1516,N_297);
or U2812 (N_2812,In_2070,In_657);
and U2813 (N_2813,In_3779,N_2492);
xnor U2814 (N_2814,In_614,N_946);
nor U2815 (N_2815,N_1547,In_2276);
or U2816 (N_2816,N_2006,N_1027);
nand U2817 (N_2817,In_3301,In_1810);
nand U2818 (N_2818,N_2112,In_2185);
and U2819 (N_2819,N_583,N_1924);
nand U2820 (N_2820,In_3551,N_934);
and U2821 (N_2821,In_2656,In_4132);
and U2822 (N_2822,N_1265,In_4924);
nor U2823 (N_2823,N_2159,In_2747);
nand U2824 (N_2824,N_2003,N_1309);
and U2825 (N_2825,N_89,N_1985);
nand U2826 (N_2826,N_1347,In_1300);
nand U2827 (N_2827,N_1092,N_1854);
nor U2828 (N_2828,N_25,N_1029);
xnor U2829 (N_2829,N_1274,N_781);
or U2830 (N_2830,In_4422,N_1928);
or U2831 (N_2831,N_828,In_4344);
or U2832 (N_2832,In_4057,In_530);
xor U2833 (N_2833,In_1616,In_3099);
or U2834 (N_2834,In_4634,In_1607);
nand U2835 (N_2835,N_885,N_1736);
nor U2836 (N_2836,N_1138,N_1508);
and U2837 (N_2837,N_1778,N_260);
and U2838 (N_2838,N_2437,N_303);
or U2839 (N_2839,N_1003,N_1119);
and U2840 (N_2840,N_494,N_2079);
nor U2841 (N_2841,In_139,N_1767);
xor U2842 (N_2842,In_820,In_3517);
nand U2843 (N_2843,In_2110,In_4885);
nand U2844 (N_2844,N_1831,In_3825);
nand U2845 (N_2845,N_147,N_1162);
xnor U2846 (N_2846,In_1819,N_55);
or U2847 (N_2847,N_710,N_876);
nor U2848 (N_2848,N_1594,N_1946);
nor U2849 (N_2849,N_2138,In_1005);
nor U2850 (N_2850,In_4153,N_2314);
nand U2851 (N_2851,N_1718,N_989);
nand U2852 (N_2852,N_1937,In_2415);
or U2853 (N_2853,In_1916,In_350);
and U2854 (N_2854,N_986,N_632);
or U2855 (N_2855,In_3641,N_1171);
and U2856 (N_2856,In_1778,In_1418);
xnor U2857 (N_2857,N_27,In_864);
or U2858 (N_2858,N_1499,N_239);
or U2859 (N_2859,In_4421,In_3819);
nand U2860 (N_2860,In_3596,N_993);
and U2861 (N_2861,N_606,N_1698);
nor U2862 (N_2862,N_800,In_3936);
and U2863 (N_2863,In_285,In_710);
nor U2864 (N_2864,N_1324,N_315);
or U2865 (N_2865,In_2459,N_1148);
and U2866 (N_2866,N_2405,N_1483);
nand U2867 (N_2867,N_2204,N_1725);
nand U2868 (N_2868,In_2994,In_1551);
nand U2869 (N_2869,In_1924,N_826);
xnor U2870 (N_2870,N_1152,In_4920);
xnor U2871 (N_2871,N_2435,In_4076);
or U2872 (N_2872,N_2439,In_977);
nand U2873 (N_2873,N_163,N_619);
or U2874 (N_2874,N_2454,N_2141);
or U2875 (N_2875,N_2482,In_2919);
nor U2876 (N_2876,In_4052,In_2455);
xor U2877 (N_2877,In_2726,N_2092);
nor U2878 (N_2878,In_1601,N_2351);
nand U2879 (N_2879,N_2135,N_1502);
nand U2880 (N_2880,N_2371,N_2155);
or U2881 (N_2881,N_81,In_1291);
and U2882 (N_2882,In_4893,N_877);
xor U2883 (N_2883,In_3235,In_1032);
and U2884 (N_2884,N_1564,In_857);
or U2885 (N_2885,N_1445,N_2401);
or U2886 (N_2886,N_2201,N_350);
nand U2887 (N_2887,N_144,N_1120);
nand U2888 (N_2888,In_4575,N_1953);
nand U2889 (N_2889,N_1352,In_4523);
xor U2890 (N_2890,In_4564,In_2223);
nand U2891 (N_2891,In_118,N_2448);
and U2892 (N_2892,In_3777,N_1822);
xor U2893 (N_2893,In_836,N_2217);
nand U2894 (N_2894,In_1656,N_1374);
nor U2895 (N_2895,In_2215,N_1036);
or U2896 (N_2896,In_2434,N_631);
or U2897 (N_2897,In_1706,N_2258);
or U2898 (N_2898,In_3045,In_3665);
nand U2899 (N_2899,In_2821,In_563);
and U2900 (N_2900,N_1191,N_694);
nand U2901 (N_2901,N_2426,In_4363);
or U2902 (N_2902,N_2390,In_3751);
xor U2903 (N_2903,In_516,In_2373);
xor U2904 (N_2904,In_3919,N_1849);
nand U2905 (N_2905,N_1769,In_1180);
xor U2906 (N_2906,N_1898,N_1993);
and U2907 (N_2907,N_280,N_1621);
or U2908 (N_2908,In_3678,N_984);
and U2909 (N_2909,N_545,N_2180);
and U2910 (N_2910,In_4946,In_3578);
nand U2911 (N_2911,N_709,N_2499);
nand U2912 (N_2912,N_1235,In_2934);
or U2913 (N_2913,N_244,N_2322);
nand U2914 (N_2914,N_529,N_1008);
nor U2915 (N_2915,N_2031,In_1788);
and U2916 (N_2916,N_2246,In_1307);
nor U2917 (N_2917,N_2422,In_3566);
xor U2918 (N_2918,N_2140,N_1057);
and U2919 (N_2919,In_4330,N_745);
xor U2920 (N_2920,N_1793,In_1202);
or U2921 (N_2921,N_2458,N_1838);
nor U2922 (N_2922,N_1173,N_2048);
nor U2923 (N_2923,N_2397,N_1845);
nand U2924 (N_2924,In_660,N_757);
xnor U2925 (N_2925,N_2121,N_373);
or U2926 (N_2926,In_3464,N_2479);
or U2927 (N_2927,In_4042,N_1774);
and U2928 (N_2928,N_2200,In_1867);
nand U2929 (N_2929,N_2099,N_907);
nand U2930 (N_2930,N_2261,N_2445);
xnor U2931 (N_2931,In_1273,In_1500);
nor U2932 (N_2932,In_2399,N_1425);
nor U2933 (N_2933,In_169,N_1550);
xnor U2934 (N_2934,N_1642,In_1802);
or U2935 (N_2935,N_1589,N_2146);
nand U2936 (N_2936,N_1113,In_2649);
or U2937 (N_2937,N_785,N_2192);
nor U2938 (N_2938,In_625,In_42);
nor U2939 (N_2939,In_446,N_1350);
and U2940 (N_2940,N_181,In_664);
or U2941 (N_2941,N_450,In_712);
xor U2942 (N_2942,In_3438,In_1283);
or U2943 (N_2943,N_1840,N_1506);
and U2944 (N_2944,In_2013,N_587);
or U2945 (N_2945,N_1631,N_1236);
xor U2946 (N_2946,N_1776,In_1860);
nor U2947 (N_2947,In_205,N_2328);
nand U2948 (N_2948,N_2013,In_1398);
xnor U2949 (N_2949,In_335,In_2729);
nand U2950 (N_2950,In_91,In_288);
xnor U2951 (N_2951,N_2318,N_1530);
or U2952 (N_2952,N_381,N_617);
xnor U2953 (N_2953,N_1888,N_1292);
and U2954 (N_2954,N_2161,N_2177);
nand U2955 (N_2955,N_1626,In_1318);
or U2956 (N_2956,N_2491,N_2206);
and U2957 (N_2957,In_4748,N_2239);
xor U2958 (N_2958,N_2127,N_1064);
and U2959 (N_2959,In_4194,N_2487);
and U2960 (N_2960,N_1929,N_670);
xnor U2961 (N_2961,In_1783,N_1782);
and U2962 (N_2962,In_1737,N_1497);
nand U2963 (N_2963,In_266,N_1695);
xor U2964 (N_2964,In_404,N_2497);
and U2965 (N_2965,N_2235,N_1153);
nand U2966 (N_2966,In_1941,In_4061);
or U2967 (N_2967,N_2378,In_806);
xnor U2968 (N_2968,N_1408,In_2124);
or U2969 (N_2969,N_273,N_1549);
nor U2970 (N_2970,N_2108,N_1129);
nand U2971 (N_2971,In_471,N_2413);
and U2972 (N_2972,In_2182,In_3701);
nor U2973 (N_2973,N_2368,In_2440);
nand U2974 (N_2974,In_3577,N_2281);
nor U2975 (N_2975,N_1830,N_1496);
nor U2976 (N_2976,In_1964,In_1894);
and U2977 (N_2977,N_1155,N_1041);
xor U2978 (N_2978,N_1137,In_2170);
or U2979 (N_2979,N_2165,In_4590);
or U2980 (N_2980,In_1878,In_145);
xnor U2981 (N_2981,In_3098,N_1785);
nor U2982 (N_2982,In_4626,N_1094);
and U2983 (N_2983,N_719,N_2431);
xnor U2984 (N_2984,In_2707,N_301);
nor U2985 (N_2985,In_3449,In_4284);
xnor U2986 (N_2986,N_2433,In_2654);
and U2987 (N_2987,In_1886,N_1693);
xnor U2988 (N_2988,N_2407,N_1301);
and U2989 (N_2989,N_773,N_2375);
and U2990 (N_2990,N_2162,In_2004);
and U2991 (N_2991,In_4244,N_122);
nor U2992 (N_2992,N_2202,N_2317);
xor U2993 (N_2993,In_1399,N_1835);
and U2994 (N_2994,N_1434,In_4715);
nand U2995 (N_2995,N_2219,N_141);
and U2996 (N_2996,N_2145,In_2889);
or U2997 (N_2997,In_3219,In_2582);
nand U2998 (N_2998,N_1705,N_1653);
or U2999 (N_2999,N_2080,N_433);
and U3000 (N_3000,In_1882,In_4696);
or U3001 (N_3001,N_1206,N_2432);
nand U3002 (N_3002,In_4220,In_4238);
nor U3003 (N_3003,In_3456,In_378);
or U3004 (N_3004,N_2501,N_1270);
xnor U3005 (N_3005,N_835,N_2005);
and U3006 (N_3006,In_1103,In_3544);
and U3007 (N_3007,N_2071,N_1813);
nor U3008 (N_3008,N_485,N_1551);
or U3009 (N_3009,N_2053,N_2617);
nor U3010 (N_3010,N_2853,In_4467);
nor U3011 (N_3011,N_2552,N_2489);
nand U3012 (N_3012,N_2509,In_1562);
xnor U3013 (N_3013,N_2599,In_1623);
xnor U3014 (N_3014,N_2150,N_2264);
xnor U3015 (N_3015,In_4928,In_785);
or U3016 (N_3016,N_2040,N_2785);
nand U3017 (N_3017,N_2788,N_2113);
and U3018 (N_3018,N_2132,N_2321);
xnor U3019 (N_3019,In_3795,N_1593);
nand U3020 (N_3020,N_1811,N_2925);
and U3021 (N_3021,In_4473,N_1636);
or U3022 (N_3022,N_148,N_1909);
nor U3023 (N_3023,In_4223,N_1886);
or U3024 (N_3024,N_2034,In_3002);
nand U3025 (N_3025,In_903,In_3912);
nand U3026 (N_3026,In_2734,N_2868);
or U3027 (N_3027,N_491,N_1118);
and U3028 (N_3028,N_849,N_774);
or U3029 (N_3029,N_1781,N_653);
nor U3030 (N_3030,N_741,N_2083);
nand U3031 (N_3031,N_2544,N_2762);
or U3032 (N_3032,N_2793,In_155);
xor U3033 (N_3033,N_2833,In_1218);
xor U3034 (N_3034,N_2611,In_3760);
xnor U3035 (N_3035,N_1438,N_2471);
xnor U3036 (N_3036,In_1460,N_2425);
nor U3037 (N_3037,In_2367,N_2646);
nor U3038 (N_3038,N_1662,In_760);
xor U3039 (N_3039,In_1312,In_3808);
and U3040 (N_3040,In_4918,N_1050);
or U3041 (N_3041,N_2550,N_2802);
and U3042 (N_3042,In_2676,N_2967);
nor U3043 (N_3043,N_232,N_2981);
nand U3044 (N_3044,N_1482,N_2598);
xor U3045 (N_3045,N_6,In_3062);
nor U3046 (N_3046,N_1917,N_1098);
nor U3047 (N_3047,In_4763,N_2073);
nor U3048 (N_3048,N_2849,In_4182);
nand U3049 (N_3049,N_2883,N_2784);
nand U3050 (N_3050,N_2705,N_2203);
and U3051 (N_3051,N_2383,N_1792);
nor U3052 (N_3052,In_3196,N_2115);
or U3053 (N_3053,In_1812,N_2233);
nand U3054 (N_3054,N_1921,N_2392);
and U3055 (N_3055,In_4980,N_2731);
xor U3056 (N_3056,N_2696,N_1992);
xor U3057 (N_3057,In_2498,In_535);
xor U3058 (N_3058,N_2912,In_379);
nor U3059 (N_3059,N_1728,N_2366);
nor U3060 (N_3060,N_2299,N_616);
or U3061 (N_3061,N_861,In_2368);
or U3062 (N_3062,N_113,N_252);
or U3063 (N_3063,N_2964,N_1708);
or U3064 (N_3064,N_2736,In_1148);
nor U3065 (N_3065,N_2570,N_1351);
xor U3066 (N_3066,In_4451,N_2484);
or U3067 (N_3067,N_1716,N_2993);
nor U3068 (N_3068,In_996,N_2249);
xor U3069 (N_3069,In_4661,N_1647);
nor U3070 (N_3070,N_155,In_3213);
nor U3071 (N_3071,In_4471,In_3303);
or U3072 (N_3072,N_1249,In_3571);
nand U3073 (N_3073,N_2922,In_29);
and U3074 (N_3074,N_1868,N_2814);
xnor U3075 (N_3075,N_2038,In_2692);
and U3076 (N_3076,N_1691,N_2692);
or U3077 (N_3077,In_1692,In_3230);
or U3078 (N_3078,N_2208,N_805);
and U3079 (N_3079,N_221,In_4309);
nand U3080 (N_3080,N_2363,N_2972);
and U3081 (N_3081,N_717,N_2860);
nand U3082 (N_3082,N_1025,N_2988);
or U3083 (N_3083,In_4114,N_1145);
xor U3084 (N_3084,In_1489,In_2970);
nor U3085 (N_3085,In_1757,N_2285);
or U3086 (N_3086,In_2390,N_1684);
nor U3087 (N_3087,N_368,In_417);
nor U3088 (N_3088,N_1692,In_1538);
nor U3089 (N_3089,N_2540,In_400);
nor U3090 (N_3090,N_2952,N_487);
xor U3091 (N_3091,N_1817,N_1903);
nand U3092 (N_3092,N_949,In_3477);
xnor U3093 (N_3093,N_1881,N_1570);
or U3094 (N_3094,N_267,In_1284);
nand U3095 (N_3095,In_4753,N_2396);
nand U3096 (N_3096,N_1863,N_1893);
nand U3097 (N_3097,In_85,In_2870);
xor U3098 (N_3098,In_1217,N_2805);
or U3099 (N_3099,In_663,N_1176);
nand U3100 (N_3100,In_1373,N_1533);
nor U3101 (N_3101,N_2908,N_1125);
and U3102 (N_3102,In_919,N_2667);
and U3103 (N_3103,N_442,N_2962);
xor U3104 (N_3104,N_2546,N_2467);
xor U3105 (N_3105,In_1672,In_1786);
nand U3106 (N_3106,In_2237,In_2159);
and U3107 (N_3107,In_4392,In_4313);
or U3108 (N_3108,N_2670,In_203);
xor U3109 (N_3109,N_1103,In_2851);
nor U3110 (N_3110,In_2494,In_2826);
nand U3111 (N_3111,N_137,In_3766);
xnor U3112 (N_3112,N_2863,N_2715);
nand U3113 (N_3113,In_1949,N_2530);
or U3114 (N_3114,N_1503,N_2772);
nor U3115 (N_3115,N_1548,N_2098);
nand U3116 (N_3116,In_4693,In_2158);
xor U3117 (N_3117,N_2593,N_2075);
and U3118 (N_3118,In_1016,N_1512);
or U3119 (N_3119,N_1906,N_2920);
nor U3120 (N_3120,In_4703,N_2899);
nand U3121 (N_3121,N_2185,N_2904);
or U3122 (N_3122,In_1676,N_2975);
xor U3123 (N_3123,N_2585,N_2787);
nor U3124 (N_3124,N_1256,In_2014);
or U3125 (N_3125,N_2376,In_2078);
nand U3126 (N_3126,N_2516,N_1799);
nor U3127 (N_3127,N_1196,N_2669);
nand U3128 (N_3128,N_2283,N_1926);
and U3129 (N_3129,In_4736,N_2845);
xnor U3130 (N_3130,N_519,N_2276);
nand U3131 (N_3131,In_226,N_2342);
xnor U3132 (N_3132,N_2028,N_2721);
or U3133 (N_3133,In_1854,N_1073);
nor U3134 (N_3134,N_2587,In_26);
and U3135 (N_3135,In_4026,N_1775);
xor U3136 (N_3136,N_73,N_2197);
and U3137 (N_3137,In_4524,N_1777);
xnor U3138 (N_3138,N_2797,N_1214);
and U3139 (N_3139,N_2974,N_2567);
xor U3140 (N_3140,In_1052,N_2895);
or U3141 (N_3141,In_1299,N_2184);
or U3142 (N_3142,In_844,N_2228);
nor U3143 (N_3143,In_1282,N_2723);
xor U3144 (N_3144,In_2166,In_971);
xor U3145 (N_3145,N_2968,In_1745);
xnor U3146 (N_3146,In_3185,In_3687);
or U3147 (N_3147,N_1749,N_2500);
and U3148 (N_3148,N_2029,N_1606);
nor U3149 (N_3149,N_2522,In_671);
nor U3150 (N_3150,N_414,N_889);
and U3151 (N_3151,N_2679,N_2296);
nor U3152 (N_3152,In_1255,In_2235);
nand U3153 (N_3153,In_4266,N_2404);
or U3154 (N_3154,N_2813,N_2494);
nor U3155 (N_3155,In_4761,N_2986);
nor U3156 (N_3156,N_1739,N_2976);
and U3157 (N_3157,N_1699,N_2866);
or U3158 (N_3158,In_3496,N_2523);
nand U3159 (N_3159,N_275,In_2887);
xor U3160 (N_3160,In_3164,In_4480);
or U3161 (N_3161,N_62,N_2095);
nand U3162 (N_3162,N_2400,In_745);
and U3163 (N_3163,N_2379,N_1365);
nor U3164 (N_3164,In_902,In_4598);
nor U3165 (N_3165,In_3754,N_2790);
xnor U3166 (N_3166,N_1889,N_1646);
xor U3167 (N_3167,N_2623,In_789);
nor U3168 (N_3168,In_4,N_1023);
nand U3169 (N_3169,N_1251,In_1461);
or U3170 (N_3170,In_6,In_2722);
nor U3171 (N_3171,In_3755,In_856);
nand U3172 (N_3172,N_2143,N_2819);
xnor U3173 (N_3173,N_2823,N_2302);
nand U3174 (N_3174,N_814,N_2893);
xnor U3175 (N_3175,In_2695,N_2537);
or U3176 (N_3176,N_2998,N_2183);
nand U3177 (N_3177,In_1859,In_2264);
nor U3178 (N_3178,N_2584,N_2100);
nor U3179 (N_3179,In_4759,N_2637);
xor U3180 (N_3180,In_2784,In_428);
and U3181 (N_3181,In_358,In_4963);
and U3182 (N_3182,N_1111,N_2672);
xor U3183 (N_3183,In_40,N_2938);
nor U3184 (N_3184,In_1751,In_4725);
xor U3185 (N_3185,In_1800,In_28);
or U3186 (N_3186,N_2120,N_1751);
and U3187 (N_3187,In_1525,N_965);
or U3188 (N_3188,In_737,N_2903);
nand U3189 (N_3189,N_2655,N_2122);
nand U3190 (N_3190,N_2882,In_805);
xnor U3191 (N_3191,In_4690,In_311);
or U3192 (N_3192,N_2571,In_3636);
and U3193 (N_3193,N_2464,N_2331);
or U3194 (N_3194,In_2409,N_767);
and U3195 (N_3195,In_4979,In_2527);
nand U3196 (N_3196,In_2711,N_2410);
nand U3197 (N_3197,In_908,In_2861);
and U3198 (N_3198,N_2693,In_4306);
nand U3199 (N_3199,N_1613,N_2735);
or U3200 (N_3200,N_2110,In_3723);
nand U3201 (N_3201,In_3147,In_2382);
nor U3202 (N_3202,In_1313,N_1323);
and U3203 (N_3203,In_528,In_4581);
nor U3204 (N_3204,N_2712,In_4637);
xor U3205 (N_3205,N_2644,N_1329);
nor U3206 (N_3206,N_2888,N_2408);
and U3207 (N_3207,N_1580,In_3132);
xor U3208 (N_3208,In_1945,N_2711);
or U3209 (N_3209,In_1684,In_1008);
or U3210 (N_3210,In_2785,N_32);
and U3211 (N_3211,N_1154,N_1598);
nor U3212 (N_3212,N_2087,N_2290);
and U3213 (N_3213,N_2871,N_2760);
xor U3214 (N_3214,N_718,N_340);
xor U3215 (N_3215,N_2106,N_2514);
or U3216 (N_3216,N_2773,N_2953);
or U3217 (N_3217,In_333,N_1447);
nor U3218 (N_3218,In_4197,In_2115);
nand U3219 (N_3219,In_816,N_2653);
and U3220 (N_3220,N_873,N_2701);
or U3221 (N_3221,N_804,In_4543);
nand U3222 (N_3222,N_2783,N_1478);
nand U3223 (N_3223,N_2245,N_2680);
or U3224 (N_3224,N_2844,N_2734);
nor U3225 (N_3225,N_2527,In_1465);
nand U3226 (N_3226,In_2320,N_2104);
nand U3227 (N_3227,N_1968,N_2751);
nand U3228 (N_3228,N_2830,N_1387);
and U3229 (N_3229,N_1187,N_1884);
nand U3230 (N_3230,In_4006,N_2348);
or U3231 (N_3231,N_743,N_2398);
or U3232 (N_3232,N_2534,In_2034);
nand U3233 (N_3233,N_2662,N_2627);
nand U3234 (N_3234,N_102,N_2223);
nor U3235 (N_3235,N_2654,In_4327);
or U3236 (N_3236,In_3345,N_422);
or U3237 (N_3237,N_2119,N_2284);
nand U3238 (N_3238,N_1524,N_2914);
nor U3239 (N_3239,N_1542,N_2297);
nand U3240 (N_3240,N_1986,In_3679);
and U3241 (N_3241,N_1420,In_766);
nand U3242 (N_3242,N_2985,N_2743);
xnor U3243 (N_3243,N_2488,N_465);
xor U3244 (N_3244,N_2977,In_4630);
nand U3245 (N_3245,In_1539,N_1615);
or U3246 (N_3246,N_2327,In_4909);
and U3247 (N_3247,N_2107,In_2725);
or U3248 (N_3248,N_2513,N_1640);
xor U3249 (N_3249,In_2488,In_2563);
nor U3250 (N_3250,N_2081,N_1200);
or U3251 (N_3251,N_2532,N_1066);
or U3252 (N_3252,N_2958,N_2665);
xor U3253 (N_3253,N_2940,In_300);
nor U3254 (N_3254,In_2193,In_1606);
or U3255 (N_3255,N_2566,N_1523);
nand U3256 (N_3256,N_1677,In_4501);
nor U3257 (N_3257,N_1914,N_2365);
xor U3258 (N_3258,In_4065,N_2313);
nand U3259 (N_3259,N_605,N_994);
xnor U3260 (N_3260,N_2836,N_852);
or U3261 (N_3261,N_439,N_15);
and U3262 (N_3262,N_2915,N_937);
and U3263 (N_3263,N_2862,N_2878);
nand U3264 (N_3264,N_1344,N_2238);
nand U3265 (N_3265,N_1402,N_278);
and U3266 (N_3266,In_960,N_2061);
nand U3267 (N_3267,In_4833,In_177);
or U3268 (N_3268,N_2700,N_2626);
nand U3269 (N_3269,N_1859,In_322);
xor U3270 (N_3270,In_4237,In_1240);
or U3271 (N_3271,N_1618,N_2084);
xor U3272 (N_3272,N_728,N_1212);
nand U3273 (N_3273,N_355,In_9);
and U3274 (N_3274,In_2839,N_2864);
or U3275 (N_3275,In_2547,N_1559);
xor U3276 (N_3276,In_3019,N_2776);
or U3277 (N_3277,In_1545,N_92);
or U3278 (N_3278,N_2588,N_2478);
and U3279 (N_3279,N_897,N_2498);
or U3280 (N_3280,N_1393,N_2742);
nand U3281 (N_3281,In_1528,N_2822);
nand U3282 (N_3282,In_2231,N_2068);
or U3283 (N_3283,In_3744,In_4702);
nor U3284 (N_3284,N_2917,N_961);
xnor U3285 (N_3285,In_3060,N_1866);
nand U3286 (N_3286,N_2035,N_2775);
nor U3287 (N_3287,N_2948,N_2641);
and U3288 (N_3288,In_3548,In_245);
xor U3289 (N_3289,N_1479,N_2051);
xnor U3290 (N_3290,N_1081,N_2231);
and U3291 (N_3291,N_2449,In_3868);
nand U3292 (N_3292,N_2607,N_2130);
and U3293 (N_3293,N_1800,N_2898);
nor U3294 (N_3294,In_3606,In_3788);
or U3295 (N_3295,N_2555,In_116);
nand U3296 (N_3296,N_2656,N_2329);
nand U3297 (N_3297,N_2503,N_2749);
and U3298 (N_3298,In_4047,N_1308);
xnor U3299 (N_3299,In_1828,In_3615);
nor U3300 (N_3300,N_2651,In_2051);
nor U3301 (N_3301,N_2726,In_695);
nand U3302 (N_3302,In_2152,N_1984);
or U3303 (N_3303,In_325,N_1180);
nand U3304 (N_3304,N_2817,N_1780);
or U3305 (N_3305,In_1366,N_2782);
xor U3306 (N_3306,N_2999,N_634);
nor U3307 (N_3307,N_1747,In_763);
nand U3308 (N_3308,N_2850,In_3830);
xnor U3309 (N_3309,N_1011,In_2204);
and U3310 (N_3310,N_2524,N_2447);
and U3311 (N_3311,N_2791,N_884);
nor U3312 (N_3312,N_2916,N_2690);
or U3313 (N_3313,In_1977,N_2733);
and U3314 (N_3314,In_2427,In_3705);
and U3315 (N_3315,In_4224,N_1388);
nand U3316 (N_3316,In_86,N_2596);
nand U3317 (N_3317,N_478,N_2529);
and U3318 (N_3318,N_2014,N_2416);
and U3319 (N_3319,N_2412,In_1336);
nand U3320 (N_3320,N_2535,N_1938);
nand U3321 (N_3321,N_1855,N_2932);
nand U3322 (N_3322,N_295,N_918);
and U3323 (N_3323,N_1349,N_1228);
xor U3324 (N_3324,In_3809,N_2777);
nand U3325 (N_3325,N_664,N_1604);
or U3326 (N_3326,N_1232,N_2984);
xor U3327 (N_3327,N_1055,N_1405);
xnor U3328 (N_3328,N_2913,N_2295);
nand U3329 (N_3329,In_3569,N_2897);
nand U3330 (N_3330,N_1068,N_1955);
or U3331 (N_3331,In_50,N_1638);
nor U3332 (N_3332,N_1803,In_1279);
xor U3333 (N_3333,N_888,N_2592);
or U3334 (N_3334,N_2622,In_4649);
xnor U3335 (N_3335,In_2644,N_2876);
or U3336 (N_3336,N_2877,N_2941);
xor U3337 (N_3337,N_1627,N_2456);
nor U3338 (N_3338,In_1824,N_1706);
xor U3339 (N_3339,N_851,In_4717);
nor U3340 (N_3340,In_3191,In_201);
nand U3341 (N_3341,In_2082,In_1349);
nand U3342 (N_3342,N_2919,In_4732);
nand U3343 (N_3343,N_2472,N_231);
and U3344 (N_3344,N_899,In_2331);
nand U3345 (N_3345,In_3886,N_2798);
and U3346 (N_3346,N_1900,N_2027);
nor U3347 (N_3347,N_1871,N_2357);
or U3348 (N_3348,N_2635,N_2147);
nand U3349 (N_3349,In_3258,In_1530);
xnor U3350 (N_3350,N_1890,In_1271);
and U3351 (N_3351,N_1432,N_2178);
nand U3352 (N_3352,In_3869,In_4943);
nor U3353 (N_3353,N_1166,N_2638);
and U3354 (N_3354,N_2792,In_4367);
and U3355 (N_3355,N_2710,N_2157);
and U3356 (N_3356,N_2786,N_483);
xnor U3357 (N_3357,In_3318,N_2323);
xor U3358 (N_3358,N_1763,N_2575);
nor U3359 (N_3359,N_2589,N_2603);
xor U3360 (N_3360,N_1797,N_1519);
nor U3361 (N_3361,N_2828,N_1124);
nor U3362 (N_3362,In_153,N_2094);
nand U3363 (N_3363,N_1261,In_4698);
xnor U3364 (N_3364,N_67,N_2483);
nor U3365 (N_3365,In_4925,N_1989);
nand U3366 (N_3366,In_3767,N_735);
nor U3367 (N_3367,N_1333,N_2309);
nor U3368 (N_3368,N_2230,In_68);
nand U3369 (N_3369,N_2673,N_2310);
xor U3370 (N_3370,N_96,N_2842);
nand U3371 (N_3371,N_2163,In_3030);
xnor U3372 (N_3372,In_3594,N_1809);
or U3373 (N_3373,N_2758,N_2841);
xor U3374 (N_3374,In_2248,N_2745);
or U3375 (N_3375,N_2466,N_2222);
nor U3376 (N_3376,In_3077,N_2856);
and U3377 (N_3377,N_1942,N_2924);
or U3378 (N_3378,N_1810,N_1818);
and U3379 (N_3379,In_1926,In_897);
and U3380 (N_3380,N_2334,In_2975);
or U3381 (N_3381,N_2105,In_2449);
nand U3382 (N_3382,N_210,N_2960);
or U3383 (N_3383,N_2821,N_1944);
nor U3384 (N_3384,In_179,In_775);
nand U3385 (N_3385,N_540,N_2340);
nand U3386 (N_3386,N_2854,N_2096);
nand U3387 (N_3387,In_131,In_4606);
nor U3388 (N_3388,In_4004,In_3715);
nor U3389 (N_3389,In_1379,In_1883);
nor U3390 (N_3390,N_2610,N_2918);
or U3391 (N_3391,N_1669,N_2704);
and U3392 (N_3392,N_2417,In_3309);
and U3393 (N_3393,N_1694,N_1603);
or U3394 (N_3394,In_234,N_2728);
and U3395 (N_3395,In_3520,In_2783);
and U3396 (N_3396,In_589,In_2913);
nand U3397 (N_3397,N_2440,N_326);
and U3398 (N_3398,In_4464,N_2294);
nand U3399 (N_3399,N_624,In_4062);
or U3400 (N_3400,In_4532,N_86);
or U3401 (N_3401,In_717,N_2551);
or U3402 (N_3402,In_855,In_770);
nand U3403 (N_3403,N_2825,In_172);
nand U3404 (N_3404,N_2591,In_585);
and U3405 (N_3405,In_2080,N_2754);
and U3406 (N_3406,In_2364,N_456);
nand U3407 (N_3407,N_2255,N_1748);
or U3408 (N_3408,N_2811,N_2549);
and U3409 (N_3409,In_4206,N_2737);
nor U3410 (N_3410,N_451,In_1540);
nor U3411 (N_3411,N_2156,N_2939);
and U3412 (N_3412,N_533,N_2597);
and U3413 (N_3413,N_2469,In_3166);
or U3414 (N_3414,N_2713,In_895);
xnor U3415 (N_3415,N_2476,N_2263);
nor U3416 (N_3416,In_4881,In_2061);
nand U3417 (N_3417,In_4382,N_2875);
xnor U3418 (N_3418,N_2045,N_2545);
or U3419 (N_3419,In_624,In_1181);
or U3420 (N_3420,N_2563,N_2531);
and U3421 (N_3421,N_2352,N_48);
nand U3422 (N_3422,N_2043,N_2547);
and U3423 (N_3423,N_2647,N_2929);
nor U3424 (N_3424,N_1961,N_440);
nand U3425 (N_3425,In_1484,In_697);
xor U3426 (N_3426,N_2216,In_628);
or U3427 (N_3427,N_1807,N_266);
or U3428 (N_3428,N_1567,N_1557);
nand U3429 (N_3429,N_2562,N_1427);
or U3430 (N_3430,N_1540,N_2455);
and U3431 (N_3431,N_2370,N_2990);
nand U3432 (N_3432,N_2037,N_640);
and U3433 (N_3433,In_2388,In_1232);
xnor U3434 (N_3434,N_2801,N_1278);
and U3435 (N_3435,N_2616,In_298);
or U3436 (N_3436,N_2746,N_2518);
nand U3437 (N_3437,In_4055,In_4207);
and U3438 (N_3438,In_3512,N_2768);
xor U3439 (N_3439,N_1709,In_1378);
xor U3440 (N_3440,N_2839,In_2554);
nor U3441 (N_3441,In_2016,N_2441);
or U3442 (N_3442,In_2935,In_4036);
or U3443 (N_3443,N_2558,In_920);
or U3444 (N_3444,N_2568,N_2629);
nor U3445 (N_3445,N_2602,N_4);
nand U3446 (N_3446,N_2718,In_3752);
and U3447 (N_3447,In_3693,In_1599);
nor U3448 (N_3448,In_3192,N_2649);
and U3449 (N_3449,N_2016,N_1920);
and U3450 (N_3450,In_1329,In_4742);
nor U3451 (N_3451,In_4644,In_2451);
or U3452 (N_3452,N_2902,In_4500);
and U3453 (N_3453,N_2987,N_2601);
xor U3454 (N_3454,In_4906,N_2256);
xnor U3455 (N_3455,In_4907,In_2172);
and U3456 (N_3456,N_1678,N_762);
xor U3457 (N_3457,N_1241,N_2496);
nand U3458 (N_3458,In_4165,N_764);
nand U3459 (N_3459,N_2694,N_554);
nor U3460 (N_3460,In_270,N_1674);
nand U3461 (N_3461,N_2428,N_2900);
and U3462 (N_3462,N_1622,N_1002);
or U3463 (N_3463,N_2660,In_2903);
or U3464 (N_3464,N_2576,N_2744);
nand U3465 (N_3465,N_2859,N_1525);
xnor U3466 (N_3466,N_1279,N_2326);
nor U3467 (N_3467,In_807,In_2012);
xnor U3468 (N_3468,N_140,N_734);
nand U3469 (N_3469,N_2042,N_1367);
xor U3470 (N_3470,N_950,In_2880);
nand U3471 (N_3471,N_2046,In_1435);
or U3472 (N_3472,In_3262,In_4711);
nand U3473 (N_3473,N_2799,N_2890);
and U3474 (N_3474,N_2172,N_1927);
and U3475 (N_3475,N_2214,N_2901);
or U3476 (N_3476,In_3437,N_2582);
nor U3477 (N_3477,N_192,In_3181);
nor U3478 (N_3478,In_4691,N_730);
and U3479 (N_3479,N_2966,N_1805);
nand U3480 (N_3480,N_2659,N_2411);
or U3481 (N_3481,N_2764,N_2004);
nand U3482 (N_3482,In_4320,N_2804);
xnor U3483 (N_3483,N_2279,N_2420);
and U3484 (N_3484,In_2348,N_2191);
nand U3485 (N_3485,In_3900,N_2684);
xnor U3486 (N_3486,N_2624,N_2800);
or U3487 (N_3487,N_609,In_13);
nor U3488 (N_3488,N_2195,N_973);
or U3489 (N_3489,N_2019,N_319);
nor U3490 (N_3490,N_1851,N_2349);
nand U3491 (N_3491,N_2959,In_1478);
nand U3492 (N_3492,In_4169,N_2148);
nand U3493 (N_3493,N_1554,N_2970);
nand U3494 (N_3494,N_383,N_2158);
and U3495 (N_3495,N_2826,N_2306);
and U3496 (N_3496,N_1644,In_3411);
nor U3497 (N_3497,In_4087,N_1611);
and U3498 (N_3498,N_2572,In_867);
nor U3499 (N_3499,N_2210,N_881);
and U3500 (N_3500,N_3272,N_3103);
nor U3501 (N_3501,N_2983,In_1534);
xor U3502 (N_3502,In_3845,N_2979);
xnor U3503 (N_3503,In_3239,N_1242);
and U3504 (N_3504,N_1400,In_1781);
xor U3505 (N_3505,In_3850,N_2687);
nand U3506 (N_3506,N_3177,N_1743);
nor U3507 (N_3507,N_3291,N_3243);
and U3508 (N_3508,In_3902,N_271);
and U3509 (N_3509,In_2622,N_2671);
or U3510 (N_3510,N_3132,N_3256);
and U3511 (N_3511,N_1857,N_2884);
nor U3512 (N_3512,In_3557,N_1536);
or U3513 (N_3513,N_1077,N_1535);
nor U3514 (N_3514,N_1934,N_2474);
and U3515 (N_3515,N_3047,N_3153);
or U3516 (N_3516,N_2444,N_2846);
and U3517 (N_3517,N_2102,N_3097);
and U3518 (N_3518,N_3368,N_1987);
nor U3519 (N_3519,In_474,In_4117);
nand U3520 (N_3520,N_2539,In_4863);
nor U3521 (N_3521,In_3907,N_1229);
nor U3522 (N_3522,In_3804,In_1276);
and U3523 (N_3523,In_583,N_3310);
nor U3524 (N_3524,N_2840,N_3483);
xor U3525 (N_3525,N_1788,N_3266);
xor U3526 (N_3526,N_2831,N_2000);
or U3527 (N_3527,N_3000,N_1571);
nor U3528 (N_3528,N_243,N_3052);
or U3529 (N_3529,In_427,N_3349);
nor U3530 (N_3530,N_3444,N_2139);
or U3531 (N_3531,In_3004,N_3484);
nand U3532 (N_3532,In_982,In_4252);
nand U3533 (N_3533,In_2387,N_3090);
nor U3534 (N_3534,N_2869,In_1522);
nor U3535 (N_3535,N_1633,N_3123);
nand U3536 (N_3536,N_3425,N_3059);
or U3537 (N_3537,N_2994,N_2194);
and U3538 (N_3538,N_3355,N_49);
nor U3539 (N_3539,N_3406,N_2969);
xnor U3540 (N_3540,N_608,In_3878);
nand U3541 (N_3541,In_4986,N_3273);
nand U3542 (N_3542,N_1085,N_1625);
xnor U3543 (N_3543,N_2675,N_2928);
xnor U3544 (N_3544,N_1049,N_2752);
and U3545 (N_3545,In_4475,In_969);
and U3546 (N_3546,N_1814,In_1767);
nand U3547 (N_3547,N_2528,N_2691);
nand U3548 (N_3548,N_3270,N_3175);
nor U3549 (N_3549,N_3361,N_3146);
nor U3550 (N_3550,N_3176,N_600);
and U3551 (N_3551,In_2037,N_3427);
or U3552 (N_3552,N_3204,N_816);
nor U3553 (N_3553,In_4329,N_2851);
nand U3554 (N_3554,N_2056,N_584);
or U3555 (N_3555,N_3110,N_436);
and U3556 (N_3556,N_3397,In_3444);
xor U3557 (N_3557,N_2560,N_3317);
xor U3558 (N_3558,N_3241,In_822);
nand U3559 (N_3559,N_3297,In_2086);
or U3560 (N_3560,N_255,N_2757);
nor U3561 (N_3561,N_2973,N_2738);
nand U3562 (N_3562,N_2288,In_4791);
nor U3563 (N_3563,N_3018,N_1450);
nand U3564 (N_3564,N_3140,N_590);
nand U3565 (N_3565,N_3464,In_3743);
nand U3566 (N_3566,N_766,N_2681);
or U3567 (N_3567,N_3049,N_2590);
nor U3568 (N_3568,In_1046,N_2010);
and U3569 (N_3569,N_2473,N_715);
or U3570 (N_3570,N_3390,N_2887);
xnor U3571 (N_3571,In_4679,N_3084);
xnor U3572 (N_3572,N_3324,N_2933);
and U3573 (N_3573,N_1952,N_3445);
xor U3574 (N_3574,In_1572,N_3334);
nor U3575 (N_3575,N_1266,N_2855);
and U3576 (N_3576,In_2958,N_3400);
or U3577 (N_3577,In_1940,In_352);
or U3578 (N_3578,N_3008,In_3046);
nand U3579 (N_3579,In_4443,In_3176);
nor U3580 (N_3580,N_3353,N_3325);
nand U3581 (N_3581,N_3498,N_3127);
xor U3582 (N_3582,N_3031,N_3025);
nor U3583 (N_3583,N_685,N_2391);
xor U3584 (N_3584,In_2485,In_3357);
and U3585 (N_3585,N_3195,N_2507);
xnor U3586 (N_3586,N_546,N_3448);
or U3587 (N_3587,N_3231,N_2824);
and U3588 (N_3588,N_3007,N_3299);
xor U3589 (N_3589,N_2658,In_4926);
nor U3590 (N_3590,N_3451,In_3937);
nand U3591 (N_3591,N_1428,N_1565);
nor U3592 (N_3592,N_3450,In_3932);
and U3593 (N_3593,N_2372,In_197);
or U3594 (N_3594,In_3058,N_2361);
and U3595 (N_3595,In_1636,N_1221);
xor U3596 (N_3596,N_3333,In_4802);
nor U3597 (N_3597,In_744,N_2770);
or U3598 (N_3598,N_3122,N_1930);
nand U3599 (N_3599,N_1443,N_3398);
and U3600 (N_3600,N_2525,In_1594);
and U3601 (N_3601,In_2265,N_2706);
and U3602 (N_3602,N_2957,N_3149);
and U3603 (N_3603,N_3165,In_2087);
and U3604 (N_3604,N_2350,N_2364);
or U3605 (N_3605,N_1883,N_1710);
and U3606 (N_3606,N_3315,N_3262);
xor U3607 (N_3607,N_2553,N_3306);
and U3608 (N_3608,N_2475,In_883);
xnor U3609 (N_3609,N_3279,N_2678);
or U3610 (N_3610,N_3494,N_2950);
nand U3611 (N_3611,N_2724,N_3305);
or U3612 (N_3612,N_2543,N_2807);
xor U3613 (N_3613,N_3106,N_3252);
or U3614 (N_3614,N_3147,In_1753);
nor U3615 (N_3615,N_1959,N_3042);
nand U3616 (N_3616,In_2961,N_2273);
and U3617 (N_3617,N_2886,N_2911);
nand U3618 (N_3618,N_586,N_3330);
nor U3619 (N_3619,N_2460,N_3160);
or U3620 (N_3620,In_3055,N_1361);
nand U3621 (N_3621,N_2837,N_1207);
xor U3622 (N_3622,N_3293,N_206);
and U3623 (N_3623,In_2294,In_2617);
xnor U3624 (N_3624,In_478,N_2419);
nand U3625 (N_3625,N_1988,In_3528);
or U3626 (N_3626,N_455,N_3274);
xnor U3627 (N_3627,In_1697,N_2809);
and U3628 (N_3628,N_3166,N_2838);
or U3629 (N_3629,N_2820,N_3189);
and U3630 (N_3630,N_1977,N_2997);
or U3631 (N_3631,N_2221,N_2930);
or U3632 (N_3632,N_750,N_1932);
xnor U3633 (N_3633,In_3490,In_1628);
or U3634 (N_3634,In_3732,N_2594);
xnor U3635 (N_3635,N_2209,N_2580);
xnor U3636 (N_3636,In_1662,In_2586);
or U3637 (N_3637,N_2319,N_2926);
nor U3638 (N_3638,N_1899,N_2755);
nor U3639 (N_3639,N_3346,N_1080);
or U3640 (N_3640,N_2894,N_2388);
and U3641 (N_3641,N_1421,N_651);
and U3642 (N_3642,In_1962,N_2872);
nand U3643 (N_3643,N_3081,In_3550);
and U3644 (N_3644,N_3462,N_3225);
or U3645 (N_3645,In_250,In_3692);
and U3646 (N_3646,N_772,N_2289);
and U3647 (N_3647,N_2695,In_1228);
nor U3648 (N_3648,N_1555,N_3321);
or U3649 (N_3649,N_2502,In_4603);
or U3650 (N_3650,N_3229,In_1452);
or U3651 (N_3651,N_2315,N_3436);
and U3652 (N_3652,N_3207,N_2065);
xor U3653 (N_3653,N_3303,N_3212);
and U3654 (N_3654,N_3275,N_2336);
nor U3655 (N_3655,N_972,N_2881);
nor U3656 (N_3656,N_3050,N_3242);
and U3657 (N_3657,N_2116,N_549);
nor U3658 (N_3658,In_2359,N_3170);
xnor U3659 (N_3659,N_2167,N_2613);
nor U3660 (N_3660,N_2753,N_672);
xnor U3661 (N_3661,In_291,In_2905);
and U3662 (N_3662,N_2865,N_2335);
nor U3663 (N_3663,N_3470,N_3214);
and U3664 (N_3664,N_2942,In_22);
xnor U3665 (N_3665,N_1590,In_2304);
xnor U3666 (N_3666,N_2077,N_2794);
xor U3667 (N_3667,N_3120,In_1514);
or U3668 (N_3668,N_1629,N_1966);
nand U3669 (N_3669,N_2090,N_2536);
nor U3670 (N_3670,N_2111,N_3351);
xnor U3671 (N_3671,N_3496,In_3194);
nor U3672 (N_3672,N_236,N_2808);
xor U3673 (N_3673,In_2149,In_2352);
and U3674 (N_3674,N_1860,In_4303);
and U3675 (N_3675,N_2293,N_268);
nor U3676 (N_3676,N_3269,In_4995);
and U3677 (N_3677,N_1189,N_2829);
nor U3678 (N_3678,In_2732,N_3327);
and U3679 (N_3679,N_1097,N_3020);
nor U3680 (N_3680,N_1663,N_2103);
and U3681 (N_3681,N_3191,N_2640);
or U3682 (N_3682,N_419,N_3283);
or U3683 (N_3683,N_3278,N_2946);
or U3684 (N_3684,N_1602,In_892);
or U3685 (N_3685,N_3341,N_3485);
nand U3686 (N_3686,N_1202,N_2722);
and U3687 (N_3687,N_2512,N_2668);
and U3688 (N_3688,N_2906,N_3366);
or U3689 (N_3689,N_2630,N_2578);
and U3690 (N_3690,N_2579,N_3245);
or U3691 (N_3691,N_3104,N_1635);
nor U3692 (N_3692,N_2674,In_4161);
nor U3693 (N_3693,In_3973,N_3064);
nor U3694 (N_3694,N_3412,N_3173);
nor U3695 (N_3695,N_3157,N_1639);
nor U3696 (N_3696,N_1757,N_2320);
and U3697 (N_3697,N_3186,N_3460);
xnor U3698 (N_3698,N_3258,N_1852);
nand U3699 (N_3699,In_4163,N_2088);
or U3700 (N_3700,N_1925,N_1491);
nand U3701 (N_3701,N_3216,N_3159);
nand U3702 (N_3702,N_2727,N_2131);
nor U3703 (N_3703,In_357,N_3061);
xor U3704 (N_3704,N_1628,N_1760);
nand U3705 (N_3705,N_3232,N_2848);
and U3706 (N_3706,In_2092,In_4755);
nor U3707 (N_3707,N_2621,N_3088);
or U3708 (N_3708,N_671,N_3392);
or U3709 (N_3709,N_3251,In_736);
and U3710 (N_3710,In_1038,N_3155);
nor U3711 (N_3711,N_1552,N_1190);
nor U3712 (N_3712,N_1974,N_2781);
nand U3713 (N_3713,In_470,N_1617);
and U3714 (N_3714,N_875,N_3004);
xor U3715 (N_3715,N_2796,In_2559);
nor U3716 (N_3716,N_3280,N_3197);
xnor U3717 (N_3717,In_3832,N_1510);
xnor U3718 (N_3718,N_3046,In_1513);
nor U3719 (N_3719,N_3376,N_3210);
xor U3720 (N_3720,N_3023,N_3309);
xor U3721 (N_3721,N_3092,N_3383);
nor U3722 (N_3722,N_2720,In_933);
or U3723 (N_3723,N_1108,N_2244);
and U3724 (N_3724,N_3362,N_3402);
and U3725 (N_3725,N_2414,N_1758);
xnor U3726 (N_3726,N_2286,N_3203);
nor U3727 (N_3727,N_2729,N_862);
and U3728 (N_3728,N_789,N_3235);
nand U3729 (N_3729,N_3429,N_2989);
nand U3730 (N_3730,N_1941,N_2698);
or U3731 (N_3731,In_2394,N_3220);
xnor U3732 (N_3732,N_2765,N_1532);
and U3733 (N_3733,In_4486,N_1837);
xnor U3734 (N_3734,N_291,N_2943);
and U3735 (N_3735,N_3240,N_563);
or U3736 (N_3736,N_3365,In_3837);
nand U3737 (N_3737,N_622,N_3183);
or U3738 (N_3738,N_2663,N_3480);
nand U3739 (N_3739,N_19,N_3224);
nor U3740 (N_3740,In_3398,In_344);
xor U3741 (N_3741,In_1835,In_2194);
nor U3742 (N_3742,N_3410,N_3345);
nand U3743 (N_3743,In_3659,N_3393);
and U3744 (N_3744,N_3083,N_2438);
and U3745 (N_3745,N_1879,N_3218);
nand U3746 (N_3746,N_3077,N_2971);
and U3747 (N_3747,N_3294,N_2756);
and U3748 (N_3748,In_587,N_2633);
xor U3749 (N_3749,In_2866,N_3385);
and U3750 (N_3750,In_4123,N_2936);
and U3751 (N_3751,N_2625,N_3072);
xnor U3752 (N_3752,N_3449,N_1672);
and U3753 (N_3753,N_2686,In_562);
nand U3754 (N_3754,In_3866,N_3128);
or U3755 (N_3755,N_1275,N_1935);
or U3756 (N_3756,N_3371,In_955);
nor U3757 (N_3757,N_2628,N_3111);
nand U3758 (N_3758,N_1045,N_3417);
nand U3759 (N_3759,In_1531,In_4203);
and U3760 (N_3760,In_4873,N_2604);
nand U3761 (N_3761,N_1820,N_662);
and U3762 (N_3762,In_4931,N_3172);
xor U3763 (N_3763,N_1383,N_3405);
and U3764 (N_3764,N_2418,N_3078);
and U3765 (N_3765,N_2612,N_3079);
and U3766 (N_3766,In_772,In_4962);
and U3767 (N_3767,N_2909,In_1699);
nor U3768 (N_3768,N_2620,N_1513);
xnor U3769 (N_3769,N_3359,N_2683);
xor U3770 (N_3770,N_2381,N_3388);
and U3771 (N_3771,N_3347,In_1234);
or U3772 (N_3772,N_1616,N_1379);
nor U3773 (N_3773,N_3307,N_3377);
xor U3774 (N_3774,N_3384,N_5);
and U3775 (N_3775,In_3133,N_3136);
nand U3776 (N_3776,In_1952,N_2559);
or U3777 (N_3777,N_68,In_15);
and U3778 (N_3778,In_4697,N_2282);
and U3779 (N_3779,N_3162,N_3441);
nand U3780 (N_3780,N_3141,N_2169);
or U3781 (N_3781,N_2661,N_2858);
and U3782 (N_3782,In_2043,In_1877);
or U3783 (N_3783,N_1652,N_2885);
xnor U3784 (N_3784,N_2874,N_3174);
nand U3785 (N_3785,N_3364,N_3156);
or U3786 (N_3786,N_3434,N_3073);
xnor U3787 (N_3787,In_3193,N_2325);
or U3788 (N_3788,N_3193,In_498);
or U3789 (N_3789,N_3472,N_3169);
xnor U3790 (N_3790,In_2666,In_1087);
and U3791 (N_3791,N_3205,N_2358);
nand U3792 (N_3792,N_2676,In_2357);
xor U3793 (N_3793,N_1456,N_1336);
nand U3794 (N_3794,N_3063,N_3014);
xnor U3795 (N_3795,In_679,N_3414);
and U3796 (N_3796,N_2789,N_2636);
or U3797 (N_3797,N_3338,N_3311);
nand U3798 (N_3798,N_2719,N_3053);
and U3799 (N_3799,N_2556,N_471);
or U3800 (N_3800,N_3350,N_2810);
or U3801 (N_3801,N_2181,In_544);
nand U3802 (N_3802,In_2259,N_3129);
nand U3803 (N_3803,N_369,In_1899);
nand U3804 (N_3804,N_3213,N_2991);
xor U3805 (N_3805,In_3400,N_2947);
or U3806 (N_3806,N_2017,N_3463);
or U3807 (N_3807,In_4195,N_3342);
xnor U3808 (N_3808,N_1574,N_2708);
nor U3809 (N_3809,In_1660,N_2750);
nand U3810 (N_3810,N_3244,N_2664);
nor U3811 (N_3811,N_1654,N_3043);
nand U3812 (N_3812,N_3194,N_3154);
nor U3813 (N_3813,N_2423,N_1948);
or U3814 (N_3814,N_3239,N_3301);
nor U3815 (N_3815,N_2332,In_410);
and U3816 (N_3816,N_1006,N_3328);
and U3817 (N_3817,N_3488,N_2677);
and U3818 (N_3818,N_1607,In_3887);
nand U3819 (N_3819,N_2186,N_3200);
nand U3820 (N_3820,N_2779,N_2072);
or U3821 (N_3821,In_4142,In_2974);
and U3822 (N_3822,N_3487,N_3001);
nor U3823 (N_3823,N_1389,N_3363);
xor U3824 (N_3824,N_2480,N_2763);
and U3825 (N_3825,In_2098,N_3479);
or U3826 (N_3826,N_3304,N_3456);
or U3827 (N_3827,N_3357,N_2225);
nand U3828 (N_3828,N_3011,N_3192);
nand U3829 (N_3829,In_1653,N_423);
and U3830 (N_3830,In_2126,In_384);
nor U3831 (N_3831,N_2123,N_3062);
or U3832 (N_3832,N_2485,In_178);
or U3833 (N_3833,N_161,In_1957);
xor U3834 (N_3834,N_1717,N_2896);
and U3835 (N_3835,In_2097,In_127);
and U3836 (N_3836,N_3439,In_3462);
nand U3837 (N_3837,N_514,N_3045);
nor U3838 (N_3838,N_3179,N_792);
nand U3839 (N_3839,N_691,N_2857);
nor U3840 (N_3840,N_3421,N_3379);
and U3841 (N_3841,N_2730,N_2506);
or U3842 (N_3842,N_3424,N_3055);
xor U3843 (N_3843,N_3284,N_3437);
xor U3844 (N_3844,N_3477,N_1907);
and U3845 (N_3845,N_2341,N_3408);
nor U3846 (N_3846,N_2771,In_4545);
nand U3847 (N_3847,N_1689,N_3308);
nand U3848 (N_3848,N_3211,In_383);
nand U3849 (N_3849,N_3331,N_3482);
nor U3850 (N_3850,In_3424,N_2951);
and U3851 (N_3851,N_2436,In_1652);
and U3852 (N_3852,N_2815,N_3407);
or U3853 (N_3853,N_10,N_3233);
xnor U3854 (N_3854,N_3428,N_1312);
nor U3855 (N_3855,N_3152,N_363);
and U3856 (N_3856,In_777,N_2277);
xor U3857 (N_3857,In_3639,N_2615);
and U3858 (N_3858,N_2648,In_4718);
nor U3859 (N_3859,N_1873,N_3348);
or U3860 (N_3860,In_224,N_2992);
or U3861 (N_3861,N_2330,N_3339);
nand U3862 (N_3862,In_3984,N_3457);
xor U3863 (N_3863,N_2795,N_2709);
nor U3864 (N_3864,N_2652,N_3182);
and U3865 (N_3865,N_2780,In_2742);
nand U3866 (N_3866,N_3234,N_3322);
nand U3867 (N_3867,In_3579,In_4045);
nor U3868 (N_3868,N_3459,N_2026);
nor U3869 (N_3869,N_3490,N_2702);
or U3870 (N_3870,In_553,N_3292);
and U3871 (N_3871,N_2538,In_1004);
xor U3872 (N_3872,N_2333,N_1724);
and U3873 (N_3873,N_2510,N_3486);
nand U3874 (N_3874,N_2002,N_3119);
xnor U3875 (N_3875,N_2965,N_3034);
and U3876 (N_3876,N_2403,N_3048);
or U3877 (N_3877,N_3277,N_2961);
nor U3878 (N_3878,In_706,N_3319);
nor U3879 (N_3879,N_3185,N_2495);
nand U3880 (N_3880,N_3121,In_698);
nand U3881 (N_3881,N_3109,N_234);
xnor U3882 (N_3882,N_3184,N_2129);
and U3883 (N_3883,N_3264,In_3924);
xor U3884 (N_3884,N_3481,In_4932);
nor U3885 (N_3885,N_3202,N_2253);
and U3886 (N_3886,N_3150,N_3003);
or U3887 (N_3887,N_3188,N_2618);
nand U3888 (N_3888,N_3474,In_3207);
and U3889 (N_3889,In_598,N_1416);
nor U3890 (N_3890,N_3074,In_2279);
xnor U3891 (N_3891,N_3344,N_1960);
nor U3892 (N_3892,In_4712,N_2052);
nor U3893 (N_3893,In_3298,In_4253);
xnor U3894 (N_3894,In_2738,In_1961);
or U3895 (N_3895,N_1779,In_741);
xor U3896 (N_3896,N_2021,In_1774);
nand U3897 (N_3897,N_1260,In_2796);
xor U3898 (N_3898,N_3391,N_2980);
and U3899 (N_3899,In_1292,N_2595);
nand U3900 (N_3900,N_3295,N_3312);
xnor U3901 (N_3901,N_2262,N_1331);
nand U3902 (N_3902,N_3337,N_2963);
xor U3903 (N_3903,N_1865,N_2689);
and U3904 (N_3904,N_1982,N_3468);
or U3905 (N_3905,N_479,N_2504);
xor U3906 (N_3906,In_4589,N_3375);
nor U3907 (N_3907,N_1577,N_3029);
and U3908 (N_3908,In_2668,In_1822);
nor U3909 (N_3909,N_3215,In_81);
nor U3910 (N_3910,In_4727,N_2606);
nor U3911 (N_3911,N_3067,N_3367);
xor U3912 (N_3912,N_3475,N_1203);
or U3913 (N_3913,N_910,N_2265);
nand U3914 (N_3914,N_3221,In_4200);
or U3915 (N_3915,In_102,N_3380);
nor U3916 (N_3916,In_1361,N_1586);
and U3917 (N_3917,N_3006,N_3017);
nor U3918 (N_3918,N_2945,N_3249);
and U3919 (N_3919,N_3164,In_3991);
xor U3920 (N_3920,N_2954,N_3161);
or U3921 (N_3921,N_3035,N_349);
xor U3922 (N_3922,N_3080,N_2047);
xor U3923 (N_3923,In_510,In_1712);
xor U3924 (N_3924,In_540,N_914);
nand U3925 (N_3925,N_1563,N_3466);
nand U3926 (N_3926,N_1954,In_4297);
nand U3927 (N_3927,N_3453,N_2033);
and U3928 (N_3928,N_2152,In_4170);
nor U3929 (N_3929,In_4403,N_2812);
xnor U3930 (N_3930,N_2232,N_3458);
and U3931 (N_3931,In_3157,N_3431);
xnor U3932 (N_3932,N_2511,N_3396);
xor U3933 (N_3933,N_1990,N_3028);
or U3934 (N_3934,N_714,N_3171);
nand U3935 (N_3935,N_3208,N_2153);
or U3936 (N_3936,N_3302,N_1738);
and U3937 (N_3937,N_2725,N_2415);
or U3938 (N_3938,N_3144,N_516);
xor U3939 (N_3939,N_1643,N_1686);
or U3940 (N_3940,N_2062,N_3187);
nor U3941 (N_3941,N_3354,N_2377);
nor U3942 (N_3942,N_3142,In_2045);
or U3943 (N_3943,N_3300,N_3019);
xnor U3944 (N_3944,In_2948,N_3255);
and U3945 (N_3945,N_2561,N_1656);
nor U3946 (N_3946,N_2074,N_2861);
nand U3947 (N_3947,In_2888,In_4952);
or U3948 (N_3948,In_1807,In_2226);
nor U3949 (N_3949,N_2430,N_2089);
xnor U3950 (N_3950,N_2044,N_3237);
or U3951 (N_3951,N_3442,In_4259);
and U3952 (N_3952,N_1468,N_898);
or U3953 (N_3953,In_495,In_1203);
and U3954 (N_3954,N_2250,N_2643);
nand U3955 (N_3955,In_4840,N_526);
and U3956 (N_3956,In_2293,N_818);
nand U3957 (N_3957,N_1106,N_3411);
nand U3958 (N_3958,N_3126,N_2011);
nor U3959 (N_3959,N_2541,N_3260);
xor U3960 (N_3960,N_3296,N_1869);
nor U3961 (N_3961,N_1082,In_900);
nor U3962 (N_3962,In_274,N_2384);
nor U3963 (N_3963,N_2477,N_2212);
and U3964 (N_3964,N_3009,N_996);
xnor U3965 (N_3965,N_3489,N_2707);
and U3966 (N_3966,N_2892,N_3394);
xor U3967 (N_3967,N_2927,N_3130);
xor U3968 (N_3968,N_385,In_1680);
or U3969 (N_3969,N_2517,N_2459);
xor U3970 (N_3970,N_14,N_2347);
nor U3971 (N_3971,N_2020,N_3452);
and U3972 (N_3972,N_723,In_999);
and U3973 (N_3973,N_3426,N_2179);
xor U3974 (N_3974,In_3972,In_4498);
nor U3975 (N_3975,N_1116,N_2657);
nand U3976 (N_3976,N_3087,N_2565);
and U3977 (N_3977,N_2015,N_2085);
nand U3978 (N_3978,N_1969,N_3473);
nor U3979 (N_3979,N_2682,N_2818);
or U3980 (N_3980,N_2688,N_1754);
nor U3981 (N_3981,In_3644,In_3625);
xnor U3982 (N_3982,N_2421,N_3263);
or U3983 (N_3983,N_2373,N_2269);
or U3984 (N_3984,N_1467,N_3024);
or U3985 (N_3985,N_2955,N_2039);
or U3986 (N_3986,N_3281,In_1643);
and U3987 (N_3987,In_2175,N_3413);
or U3988 (N_3988,In_1372,In_3649);
nand U3989 (N_3989,N_3422,N_3158);
xnor U3990 (N_3990,In_1844,In_3096);
and U3991 (N_3991,In_4729,N_3432);
xor U3992 (N_3992,N_3114,N_3247);
and U3993 (N_3993,N_3420,N_214);
nor U3994 (N_3994,N_3069,N_3015);
or U3995 (N_3995,In_1096,N_2257);
and U3996 (N_3996,N_3198,N_2631);
and U3997 (N_3997,N_3356,N_1072);
nand U3998 (N_3998,N_3492,N_1216);
or U3999 (N_3999,N_3201,N_2166);
and U4000 (N_4000,N_3707,N_3094);
xor U4001 (N_4001,N_3855,In_3537);
and U4002 (N_4002,N_3757,N_3131);
and U4003 (N_4003,N_3822,N_3814);
xnor U4004 (N_4004,N_3373,N_3401);
and U4005 (N_4005,N_3977,N_3892);
xor U4006 (N_4006,N_3726,N_3527);
nand U4007 (N_4007,N_2944,N_2934);
and U4008 (N_4008,N_3719,N_2109);
or U4009 (N_4009,In_316,N_3285);
xnor U4010 (N_4010,N_3749,N_3639);
nand U4011 (N_4011,N_3467,N_3641);
xor U4012 (N_4012,In_4775,N_3980);
nor U4013 (N_4013,N_891,N_2778);
and U4014 (N_4014,In_4666,N_2583);
or U4015 (N_4015,N_2714,N_3271);
or U4016 (N_4016,N_3525,N_2442);
and U4017 (N_4017,N_3543,N_3950);
nor U4018 (N_4018,N_3932,N_1501);
nor U4019 (N_4019,N_3013,N_2766);
nor U4020 (N_4020,N_3044,N_2521);
nand U4021 (N_4021,N_3858,N_3756);
nor U4022 (N_4022,N_3578,N_3972);
or U4023 (N_4023,N_3801,N_2609);
nand U4024 (N_4024,In_2155,N_3706);
nand U4025 (N_4025,N_3872,N_1215);
xnor U4026 (N_4026,In_1402,N_3603);
nand U4027 (N_4027,N_3725,N_3314);
xnor U4028 (N_4028,In_550,N_3139);
and U4029 (N_4029,N_2054,N_3512);
and U4030 (N_4030,In_3854,N_3638);
nor U4031 (N_4031,N_3824,N_988);
nand U4032 (N_4032,In_1912,N_3290);
xnor U4033 (N_4033,N_3605,N_3723);
and U4034 (N_4034,N_2880,N_3538);
and U4035 (N_4035,N_3879,N_3982);
nor U4036 (N_4036,N_2949,N_2338);
or U4037 (N_4037,N_2716,N_3672);
xor U4038 (N_4038,N_2870,N_2982);
nand U4039 (N_4039,In_482,N_3926);
nand U4040 (N_4040,N_3923,N_522);
nand U4041 (N_4041,N_3419,N_3771);
nor U4042 (N_4042,N_3447,N_3415);
nor U4043 (N_4043,N_3082,N_2827);
xor U4044 (N_4044,N_1634,N_3608);
nand U4045 (N_4045,N_3657,N_3236);
and U4046 (N_4046,N_3039,N_2468);
nor U4047 (N_4047,N_3542,N_3907);
and U4048 (N_4048,In_3829,N_3884);
or U4049 (N_4049,N_3724,N_2076);
nor U4050 (N_4050,N_3920,N_3071);
or U4051 (N_4051,N_3500,N_2685);
xor U4052 (N_4052,N_3763,N_2024);
nor U4053 (N_4053,N_2581,N_3145);
or U4054 (N_4054,N_1734,N_3807);
xnor U4055 (N_4055,N_3808,N_3886);
nand U4056 (N_4056,N_3526,N_3108);
nor U4057 (N_4057,N_3577,N_2739);
or U4058 (N_4058,N_3993,N_3611);
and U4059 (N_4059,N_1091,N_2847);
and U4060 (N_4060,N_3117,In_4449);
or U4061 (N_4061,N_3839,N_3943);
nand U4062 (N_4062,N_3718,In_1458);
or U4063 (N_4063,N_3919,In_229);
or U4064 (N_4064,N_2554,N_2978);
nand U4065 (N_4065,N_3734,N_736);
nand U4066 (N_4066,N_3747,N_3927);
xnor U4067 (N_4067,N_2241,N_2767);
nor U4068 (N_4068,N_1463,N_3694);
xor U4069 (N_4069,N_2564,N_3115);
and U4070 (N_4070,N_3768,N_3508);
nand U4071 (N_4071,N_2450,N_3287);
or U4072 (N_4072,N_3931,In_2634);
xor U4073 (N_4073,In_2177,N_3507);
nor U4074 (N_4074,N_3991,N_2154);
nor U4075 (N_4075,In_2316,N_3791);
nor U4076 (N_4076,N_3032,N_1474);
and U4077 (N_4077,N_3645,N_3329);
and U4078 (N_4078,N_2548,N_3717);
nand U4079 (N_4079,N_3873,N_3648);
or U4080 (N_4080,N_3866,N_2586);
xor U4081 (N_4081,N_890,N_1534);
nor U4082 (N_4082,N_3947,N_3930);
nand U4083 (N_4083,N_3504,N_3515);
and U4084 (N_4084,N_3495,N_1679);
and U4085 (N_4085,N_3836,N_3575);
nand U4086 (N_4086,N_3381,N_3819);
xor U4087 (N_4087,In_489,N_1257);
and U4088 (N_4088,N_1970,N_3286);
or U4089 (N_4089,N_3701,N_2803);
and U4090 (N_4090,N_3568,N_3086);
nand U4091 (N_4091,N_3929,In_3040);
nor U4092 (N_4092,N_3995,N_3606);
nor U4093 (N_4093,N_3758,N_3942);
or U4094 (N_4094,N_3652,N_2569);
nand U4095 (N_4095,N_3833,N_3849);
nor U4096 (N_4096,N_3689,N_3874);
and U4097 (N_4097,N_3904,N_3613);
or U4098 (N_4098,N_3567,N_3861);
nand U4099 (N_4099,N_2642,In_2724);
nor U4100 (N_4100,N_3906,N_3697);
nor U4101 (N_4101,N_3850,N_3206);
and U4102 (N_4102,N_3248,N_3683);
and U4103 (N_4103,N_3985,N_2369);
nand U4104 (N_4104,N_2748,N_1783);
nand U4105 (N_4105,In_4008,N_3016);
xnor U4106 (N_4106,N_3959,N_3829);
nor U4107 (N_4107,In_2335,N_3091);
or U4108 (N_4108,N_3790,N_3826);
nand U4109 (N_4109,N_3118,N_3880);
xor U4110 (N_4110,N_3102,N_3783);
nor U4111 (N_4111,N_1701,N_3591);
or U4112 (N_4112,N_3702,In_3430);
nor U4113 (N_4113,N_2717,N_3076);
nand U4114 (N_4114,N_3934,N_3877);
and U4115 (N_4115,N_1922,N_3894);
nand U4116 (N_4116,N_3478,In_3126);
nor U4117 (N_4117,N_2995,N_3622);
nor U4118 (N_4118,N_3497,N_3743);
xnor U4119 (N_4119,N_3668,N_3893);
nor U4120 (N_4120,N_3085,In_779);
nand U4121 (N_4121,N_3674,N_3416);
nand U4122 (N_4122,N_3853,N_3782);
nand U4123 (N_4123,N_1560,N_384);
nor U4124 (N_4124,N_3534,N_3586);
or U4125 (N_4125,N_3644,N_2697);
nand U4126 (N_4126,N_3860,N_3228);
xor U4127 (N_4127,N_3635,N_3797);
or U4128 (N_4128,N_3530,N_3340);
xnor U4129 (N_4129,N_3925,In_2922);
or U4130 (N_4130,N_3804,N_1546);
nor U4131 (N_4131,N_3780,N_3762);
nand U4132 (N_4132,N_2542,In_3998);
nor U4133 (N_4133,N_2907,N_1283);
or U4134 (N_4134,N_2268,N_3318);
nor U4135 (N_4135,N_2557,N_3838);
and U4136 (N_4136,N_1998,N_3666);
and U4137 (N_4137,In_3335,In_2181);
or U4138 (N_4138,N_3038,In_947);
nor U4139 (N_4139,N_3572,N_3370);
xnor U4140 (N_4140,N_3125,In_129);
nor U4141 (N_4141,N_3036,N_1887);
or U4142 (N_4142,N_3899,N_1058);
and U4143 (N_4143,N_2666,In_2421);
xnor U4144 (N_4144,N_3969,N_3253);
nor U4145 (N_4145,N_3446,N_2574);
nand U4146 (N_4146,N_3592,N_3659);
or U4147 (N_4147,N_3222,In_690);
xor U4148 (N_4148,In_2334,N_307);
nor U4149 (N_4149,In_4615,N_3835);
or U4150 (N_4150,N_3820,N_3057);
nand U4151 (N_4151,In_842,N_3951);
nor U4152 (N_4152,N_3806,N_3955);
and U4153 (N_4153,N_3522,N_3787);
or U4154 (N_4154,N_3505,In_4988);
nor U4155 (N_4155,N_3089,N_3915);
or U4156 (N_4156,N_1916,N_3455);
nor U4157 (N_4157,In_749,N_2931);
and U4158 (N_4158,N_2064,N_3957);
or U4159 (N_4159,N_1048,N_3547);
nand U4160 (N_4160,N_3358,N_1437);
nand U4161 (N_4161,N_3946,N_1553);
xor U4162 (N_4162,N_3544,N_3715);
and U4163 (N_4163,N_3733,N_3753);
nor U4164 (N_4164,N_3945,N_3561);
nand U4165 (N_4165,N_2134,N_3845);
and U4166 (N_4166,N_3068,N_2247);
or U4167 (N_4167,N_3903,N_3750);
nand U4168 (N_4168,N_3935,N_3887);
or U4169 (N_4169,N_3751,In_1368);
or U4170 (N_4170,N_3979,N_3852);
or U4171 (N_4171,N_3552,N_2359);
nand U4172 (N_4172,N_3630,N_3748);
nor U4173 (N_4173,N_3682,N_2889);
xnor U4174 (N_4174,N_3914,N_3802);
and U4175 (N_4175,N_3772,N_3623);
or U4176 (N_4176,N_3559,N_3847);
or U4177 (N_4177,In_90,N_3560);
or U4178 (N_4178,N_3848,N_3499);
and U4179 (N_4179,N_3545,N_3695);
and U4180 (N_4180,N_3974,N_3054);
nor U4181 (N_4181,N_3716,N_3897);
nand U4182 (N_4182,N_1735,N_3620);
nand U4183 (N_4183,N_3937,N_1282);
or U4184 (N_4184,N_3967,N_2816);
or U4185 (N_4185,N_3994,N_3138);
and U4186 (N_4186,N_3386,N_3961);
and U4187 (N_4187,N_511,N_3604);
nand U4188 (N_4188,N_2605,N_611);
nand U4189 (N_4189,N_3827,N_3677);
nor U4190 (N_4190,In_3156,N_3895);
or U4191 (N_4191,N_3335,N_3889);
and U4192 (N_4192,N_3789,N_3369);
xnor U4193 (N_4193,N_3601,N_3589);
xnor U4194 (N_4194,N_3040,N_3776);
nand U4195 (N_4195,N_3939,N_3012);
xor U4196 (N_4196,N_3135,N_3865);
and U4197 (N_4197,N_3834,N_2867);
nor U4198 (N_4198,N_3382,N_3964);
and U4199 (N_4199,N_3066,N_3662);
xnor U4200 (N_4200,N_3840,N_3681);
xnor U4201 (N_4201,N_3105,In_4225);
nand U4202 (N_4202,N_1892,N_3151);
nor U4203 (N_4203,N_3988,N_3760);
and U4204 (N_4204,N_3730,N_3583);
and U4205 (N_4205,N_3268,In_4886);
or U4206 (N_4206,N_3767,N_3493);
nor U4207 (N_4207,N_3209,N_3531);
xor U4208 (N_4208,N_3774,N_3905);
and U4209 (N_4209,In_519,N_3680);
or U4210 (N_4210,N_2834,N_3403);
nand U4211 (N_4211,N_3773,N_3671);
nor U4212 (N_4212,N_2519,N_3658);
nor U4213 (N_4213,N_3911,N_3986);
nand U4214 (N_4214,N_3343,N_3217);
xor U4215 (N_4215,N_3882,N_2619);
and U4216 (N_4216,N_2446,N_3056);
and U4217 (N_4217,N_3821,N_3825);
nand U4218 (N_4218,N_3815,N_3617);
or U4219 (N_4219,N_2353,N_3673);
nand U4220 (N_4220,In_4295,N_3711);
nand U4221 (N_4221,N_3871,N_3709);
xnor U4222 (N_4222,N_3952,N_2747);
nand U4223 (N_4223,N_3558,N_3738);
nand U4224 (N_4224,In_14,N_3588);
xnor U4225 (N_4225,N_3779,N_3777);
nand U4226 (N_4226,N_3571,N_2577);
or U4227 (N_4227,N_3863,N_3374);
nor U4228 (N_4228,N_2339,N_3631);
or U4229 (N_4229,N_2356,N_3954);
and U4230 (N_4230,N_3846,N_3703);
or U4231 (N_4231,N_2732,N_2275);
and U4232 (N_4232,N_3557,N_2451);
nand U4233 (N_4233,N_3554,N_3704);
and U4234 (N_4234,In_1039,N_3352);
or U4235 (N_4235,In_1171,N_3614);
nand U4236 (N_4236,N_3913,N_3597);
nor U4237 (N_4237,N_2632,N_3841);
nor U4238 (N_4238,N_3667,N_1823);
xnor U4239 (N_4239,N_592,N_3698);
nor U4240 (N_4240,N_3649,In_2510);
nor U4241 (N_4241,N_3831,N_3816);
and U4242 (N_4242,N_3813,N_3803);
nand U4243 (N_4243,N_3800,N_1569);
and U4244 (N_4244,N_2873,N_1208);
nor U4245 (N_4245,N_3653,N_3868);
or U4246 (N_4246,In_4420,In_4677);
xnor U4247 (N_4247,N_3565,N_3033);
or U4248 (N_4248,N_3574,N_3888);
or U4249 (N_4249,N_3070,N_3885);
or U4250 (N_4250,N_3095,N_3851);
and U4251 (N_4251,N_3984,N_3745);
nor U4252 (N_4252,N_3727,N_2355);
nor U4253 (N_4253,In_416,N_3731);
xor U4254 (N_4254,In_916,N_3687);
and U4255 (N_4255,N_457,N_3693);
xor U4256 (N_4256,N_2614,In_1567);
or U4257 (N_4257,N_3647,N_3518);
xor U4258 (N_4258,N_3143,N_3099);
nor U4259 (N_4259,N_3678,N_3736);
or U4260 (N_4260,N_3965,N_3864);
and U4261 (N_4261,N_3842,N_3968);
nor U4262 (N_4262,N_3786,N_3612);
xor U4263 (N_4263,N_3699,In_1019);
and U4264 (N_4264,N_3587,N_1700);
and U4265 (N_4265,N_3519,N_3795);
nand U4266 (N_4266,N_3710,N_2526);
and U4267 (N_4267,In_2895,N_1980);
or U4268 (N_4268,N_3532,N_3646);
or U4269 (N_4269,N_2008,N_3320);
nor U4270 (N_4270,N_3997,N_3940);
nand U4271 (N_4271,N_3562,N_3627);
and U4272 (N_4272,N_3948,N_3223);
or U4273 (N_4273,N_2060,In_1503);
and U4274 (N_4274,N_2921,N_3267);
xor U4275 (N_4275,N_3975,N_3190);
xor U4276 (N_4276,N_3844,N_3060);
or U4277 (N_4277,N_3632,N_2402);
xor U4278 (N_4278,N_3590,N_2910);
or U4279 (N_4279,N_3675,N_3941);
nor U4280 (N_4280,In_4286,N_3908);
and U4281 (N_4281,N_3506,N_3963);
and U4282 (N_4282,N_1904,N_3517);
nand U4283 (N_4283,N_3409,N_2354);
and U4284 (N_4284,In_4502,N_3389);
xor U4285 (N_4285,N_3430,N_3521);
nand U4286 (N_4286,N_3642,N_3423);
nand U4287 (N_4287,In_411,N_981);
or U4288 (N_4288,N_2171,N_3817);
and U4289 (N_4289,N_3785,N_3744);
nand U4290 (N_4290,N_1201,N_3573);
or U4291 (N_4291,N_3539,N_3818);
or U4292 (N_4292,N_3238,N_3372);
xnor U4293 (N_4293,N_2573,N_3759);
or U4294 (N_4294,N_2267,N_3005);
and U4295 (N_4295,N_3163,N_3433);
or U4296 (N_4296,N_1624,N_3541);
nand U4297 (N_4297,In_3872,N_1829);
nand U4298 (N_4298,N_3133,N_3598);
and U4299 (N_4299,N_3584,N_3728);
and U4300 (N_4300,N_3708,N_3134);
or U4301 (N_4301,N_3788,N_428);
and U4302 (N_4302,N_3944,In_3992);
or U4303 (N_4303,N_2650,N_3418);
nor U4304 (N_4304,N_1318,N_3685);
and U4305 (N_4305,N_3962,In_87);
nand U4306 (N_4306,N_3621,N_3679);
xnor U4307 (N_4307,N_3051,N_3570);
xor U4308 (N_4308,N_3246,N_3476);
and U4309 (N_4309,N_3501,N_3336);
xor U4310 (N_4310,N_3065,N_2287);
and U4311 (N_4311,N_2639,N_3812);
xnor U4312 (N_4312,In_4040,In_3966);
and U4313 (N_4313,N_3404,N_3998);
and U4314 (N_4314,N_3058,N_3761);
and U4315 (N_4315,N_3624,N_3999);
or U4316 (N_4316,N_1531,In_1434);
and U4317 (N_4317,N_3075,N_3684);
xor U4318 (N_4318,N_3721,N_1485);
or U4319 (N_4319,N_1825,N_3784);
and U4320 (N_4320,N_3890,N_3378);
xor U4321 (N_4321,In_4016,N_3026);
xnor U4322 (N_4322,N_3949,N_3933);
nor U4323 (N_4323,In_4088,N_3282);
nor U4324 (N_4324,In_329,N_3981);
xor U4325 (N_4325,N_3265,N_2272);
nand U4326 (N_4326,N_3775,N_3180);
and U4327 (N_4327,N_3626,N_3528);
nand U4328 (N_4328,N_3690,N_1666);
nor U4329 (N_4329,In_4786,N_2634);
or U4330 (N_4330,N_3737,N_3660);
nor U4331 (N_4331,N_2505,N_3615);
or U4332 (N_4332,N_3101,N_3196);
or U4333 (N_4333,N_3637,N_541);
nor U4334 (N_4334,In_2805,N_3830);
nor U4335 (N_4335,N_2759,N_3781);
xnor U4336 (N_4336,N_3435,N_3520);
xnor U4337 (N_4337,N_2308,N_2879);
xnor U4338 (N_4338,N_3799,N_1659);
nand U4339 (N_4339,N_3705,N_3655);
nand U4340 (N_4340,N_3870,In_3736);
nor U4341 (N_4341,N_641,In_4605);
nand U4342 (N_4342,N_199,N_3664);
nor U4343 (N_4343,N_3862,N_3510);
nand U4344 (N_4344,N_2645,In_1713);
nand U4345 (N_4345,N_3891,N_3516);
xnor U4346 (N_4346,N_3700,N_3794);
or U4347 (N_4347,N_3918,N_3564);
and U4348 (N_4348,N_2409,N_3902);
and U4349 (N_4349,N_930,N_3523);
or U4350 (N_4350,N_3729,N_3107);
nand U4351 (N_4351,N_3002,N_3529);
nor U4352 (N_4352,N_3769,N_3688);
and U4353 (N_4353,N_3298,N_3966);
and U4354 (N_4354,In_2486,N_2515);
or U4355 (N_4355,In_1414,In_3420);
nor U4356 (N_4356,N_3656,N_3770);
xnor U4357 (N_4357,In_3270,N_1422);
nand U4358 (N_4358,N_3654,N_3313);
nor U4359 (N_4359,In_2852,N_108);
nand U4360 (N_4360,N_3555,N_3580);
nor U4361 (N_4361,N_3765,N_3585);
or U4362 (N_4362,N_2937,N_3696);
xor U4363 (N_4363,N_3535,N_2923);
xnor U4364 (N_4364,N_3854,N_1790);
and U4365 (N_4365,N_3805,N_2703);
nand U4366 (N_4366,N_3167,N_3650);
and U4367 (N_4367,In_1094,N_3938);
or U4368 (N_4368,N_3796,In_451);
xor U4369 (N_4369,N_3629,N_3978);
xor U4370 (N_4370,N_3970,N_3250);
nor U4371 (N_4371,N_1802,N_3148);
xnor U4372 (N_4372,N_3823,N_3576);
nor U4373 (N_4373,N_3843,In_4556);
nor U4374 (N_4374,N_2699,N_2395);
xnor U4375 (N_4375,N_2453,N_3469);
and U4376 (N_4376,N_2311,N_3973);
nor U4377 (N_4377,N_3524,N_3503);
or U4378 (N_4378,N_3602,N_3692);
nor U4379 (N_4379,N_3289,N_3778);
nor U4380 (N_4380,N_3168,N_3599);
xor U4381 (N_4381,N_2385,N_3878);
nor U4382 (N_4382,N_3828,N_3566);
or U4383 (N_4383,N_3387,N_3640);
nand U4384 (N_4384,N_3625,N_3022);
nand U4385 (N_4385,N_3491,N_3593);
or U4386 (N_4386,N_3634,In_4794);
xnor U4387 (N_4387,N_3199,N_3956);
and U4388 (N_4388,N_3832,N_3764);
nor U4389 (N_4389,N_3596,N_3226);
xnor U4390 (N_4390,In_317,N_3867);
or U4391 (N_4391,In_3106,N_3792);
xor U4392 (N_4392,N_177,N_3579);
or U4393 (N_4393,In_1738,N_3259);
or U4394 (N_4394,N_3513,N_1131);
or U4395 (N_4395,N_2843,N_3910);
xnor U4396 (N_4396,N_2199,N_3595);
and U4397 (N_4397,N_3712,N_3766);
nor U4398 (N_4398,N_3619,N_2600);
nor U4399 (N_4399,N_1902,N_3537);
nor U4400 (N_4400,N_2740,In_4226);
nor U4401 (N_4401,N_3837,N_3609);
xor U4402 (N_4402,N_3230,N_3316);
nand U4403 (N_4403,N_3713,N_3027);
xor U4404 (N_4404,N_3663,N_1439);
and U4405 (N_4405,N_3720,In_2552);
and U4406 (N_4406,N_3509,In_4975);
nand U4407 (N_4407,N_3752,In_4527);
and U4408 (N_4408,N_3746,N_2832);
nor U4409 (N_4409,N_3556,N_3922);
or U4410 (N_4410,N_3581,In_230);
nand U4411 (N_4411,N_3548,N_2835);
or U4412 (N_4412,N_3928,N_3219);
nand U4413 (N_4413,N_3686,N_3628);
and U4414 (N_4414,N_3607,In_2282);
and U4415 (N_4415,N_3633,In_99);
nor U4416 (N_4416,N_3178,N_3881);
xor U4417 (N_4417,N_3987,N_3563);
or U4418 (N_4418,N_3732,N_3533);
and U4419 (N_4419,N_3569,N_3514);
or U4420 (N_4420,N_3360,N_3021);
or U4421 (N_4421,N_2996,N_3582);
nor U4422 (N_4422,N_1528,In_3749);
nor U4423 (N_4423,N_3100,N_431);
and U4424 (N_4424,N_933,N_2030);
nor U4425 (N_4425,N_3332,N_2852);
or U4426 (N_4426,In_4961,N_3960);
nand U4427 (N_4427,N_3551,N_1609);
nand U4428 (N_4428,N_3793,N_3618);
nand U4429 (N_4429,N_3440,N_3857);
nand U4430 (N_4430,N_3755,N_3096);
nor U4431 (N_4431,N_3616,N_3181);
nand U4432 (N_4432,N_1142,N_3971);
and U4433 (N_4433,N_3989,N_3990);
or U4434 (N_4434,N_705,N_2806);
and U4435 (N_4435,N_3809,N_3983);
nand U4436 (N_4436,N_3976,N_2304);
and U4437 (N_4437,N_2533,N_3869);
nand U4438 (N_4438,N_3288,N_3276);
nor U4439 (N_4439,In_4012,N_539);
nand U4440 (N_4440,N_1731,N_3461);
nor U4441 (N_4441,N_3471,N_3010);
xnor U4442 (N_4442,N_2118,N_3261);
xor U4443 (N_4443,N_3912,N_3399);
and U4444 (N_4444,N_3113,N_3921);
nor U4445 (N_4445,N_3665,N_3992);
nor U4446 (N_4446,N_1765,N_2086);
and U4447 (N_4447,N_3936,N_3443);
nor U4448 (N_4448,N_1194,N_2508);
and U4449 (N_4449,N_3600,N_3996);
nor U4450 (N_4450,N_3594,N_3546);
nor U4451 (N_4451,N_668,N_2465);
xor U4452 (N_4452,N_3856,N_3714);
nand U4453 (N_4453,N_3916,N_3550);
nand U4454 (N_4454,N_3735,N_3722);
nand U4455 (N_4455,N_1971,N_3676);
or U4456 (N_4456,N_3227,N_3740);
nand U4457 (N_4457,In_4650,N_1786);
nand U4458 (N_4458,N_3395,N_3553);
nor U4459 (N_4459,N_3549,N_3124);
nor U4460 (N_4460,N_2741,N_3636);
nand U4461 (N_4461,N_3811,N_3536);
nor U4462 (N_4462,N_3454,N_3661);
xor U4463 (N_4463,N_3112,N_3326);
nand U4464 (N_4464,In_2463,N_3438);
and U4465 (N_4465,N_2125,N_3511);
xor U4466 (N_4466,N_3875,N_2101);
and U4467 (N_4467,N_3754,N_2520);
nand U4468 (N_4468,N_2190,N_3691);
xor U4469 (N_4469,N_2891,N_3900);
nor U4470 (N_4470,N_3030,In_3787);
or U4471 (N_4471,N_3465,N_2769);
or U4472 (N_4472,N_3643,In_1728);
xor U4473 (N_4473,N_3909,N_2774);
and U4474 (N_4474,N_1454,N_2608);
xor U4475 (N_4475,N_3093,N_3742);
xnor U4476 (N_4476,N_3898,N_3651);
nand U4477 (N_4477,N_2761,In_4461);
xor U4478 (N_4478,N_3741,In_2379);
nand U4479 (N_4479,N_3859,In_3931);
and U4480 (N_4480,In_3110,In_2433);
or U4481 (N_4481,In_3234,N_1489);
nor U4482 (N_4482,N_3670,In_3187);
nand U4483 (N_4483,N_3810,In_1782);
xnor U4484 (N_4484,N_3540,N_3901);
nand U4485 (N_4485,N_3257,N_3502);
and U4486 (N_4486,N_2082,N_2956);
xor U4487 (N_4487,N_3739,N_2935);
and U4488 (N_4488,N_3323,In_4847);
xnor U4489 (N_4489,N_3798,In_3338);
nand U4490 (N_4490,N_3137,N_3098);
nand U4491 (N_4491,N_3116,In_838);
nand U4492 (N_4492,N_3917,N_3876);
nand U4493 (N_4493,N_3669,N_2266);
nand U4494 (N_4494,N_3896,N_3610);
or U4495 (N_4495,N_3883,N_3254);
or U4496 (N_4496,N_2905,N_3953);
or U4497 (N_4497,N_3037,In_2333);
or U4498 (N_4498,In_1187,N_3924);
or U4499 (N_4499,N_3041,N_3958);
and U4500 (N_4500,N_4494,N_4290);
and U4501 (N_4501,N_4133,N_4135);
or U4502 (N_4502,N_4274,N_4374);
nor U4503 (N_4503,N_4238,N_4292);
and U4504 (N_4504,N_4472,N_4232);
and U4505 (N_4505,N_4195,N_4394);
nor U4506 (N_4506,N_4301,N_4400);
or U4507 (N_4507,N_4036,N_4181);
nor U4508 (N_4508,N_4032,N_4372);
xor U4509 (N_4509,N_4276,N_4266);
xnor U4510 (N_4510,N_4401,N_4157);
xor U4511 (N_4511,N_4114,N_4188);
xor U4512 (N_4512,N_4461,N_4065);
nand U4513 (N_4513,N_4490,N_4087);
xor U4514 (N_4514,N_4284,N_4489);
nor U4515 (N_4515,N_4414,N_4345);
xnor U4516 (N_4516,N_4075,N_4039);
or U4517 (N_4517,N_4265,N_4491);
nand U4518 (N_4518,N_4455,N_4434);
nor U4519 (N_4519,N_4154,N_4331);
xor U4520 (N_4520,N_4193,N_4362);
and U4521 (N_4521,N_4113,N_4287);
xnor U4522 (N_4522,N_4302,N_4366);
nor U4523 (N_4523,N_4001,N_4465);
xor U4524 (N_4524,N_4022,N_4380);
xor U4525 (N_4525,N_4391,N_4239);
and U4526 (N_4526,N_4277,N_4329);
nand U4527 (N_4527,N_4241,N_4267);
or U4528 (N_4528,N_4378,N_4348);
and U4529 (N_4529,N_4125,N_4144);
nand U4530 (N_4530,N_4078,N_4256);
and U4531 (N_4531,N_4020,N_4245);
and U4532 (N_4532,N_4364,N_4286);
and U4533 (N_4533,N_4420,N_4224);
and U4534 (N_4534,N_4102,N_4385);
and U4535 (N_4535,N_4467,N_4179);
and U4536 (N_4536,N_4294,N_4407);
xor U4537 (N_4537,N_4166,N_4246);
nand U4538 (N_4538,N_4327,N_4080);
or U4539 (N_4539,N_4200,N_4190);
nor U4540 (N_4540,N_4122,N_4459);
and U4541 (N_4541,N_4419,N_4340);
xor U4542 (N_4542,N_4137,N_4388);
or U4543 (N_4543,N_4470,N_4175);
nor U4544 (N_4544,N_4332,N_4250);
xor U4545 (N_4545,N_4253,N_4230);
and U4546 (N_4546,N_4478,N_4344);
or U4547 (N_4547,N_4151,N_4397);
nand U4548 (N_4548,N_4028,N_4084);
nand U4549 (N_4549,N_4138,N_4269);
nand U4550 (N_4550,N_4280,N_4229);
or U4551 (N_4551,N_4043,N_4361);
or U4552 (N_4552,N_4052,N_4254);
nand U4553 (N_4553,N_4127,N_4251);
and U4554 (N_4554,N_4259,N_4024);
nand U4555 (N_4555,N_4118,N_4466);
nand U4556 (N_4556,N_4320,N_4007);
or U4557 (N_4557,N_4424,N_4045);
nor U4558 (N_4558,N_4315,N_4487);
xnor U4559 (N_4559,N_4437,N_4475);
nand U4560 (N_4560,N_4330,N_4359);
xor U4561 (N_4561,N_4495,N_4121);
and U4562 (N_4562,N_4449,N_4021);
nor U4563 (N_4563,N_4334,N_4077);
xor U4564 (N_4564,N_4070,N_4025);
nand U4565 (N_4565,N_4221,N_4278);
xnor U4566 (N_4566,N_4396,N_4428);
or U4567 (N_4567,N_4268,N_4196);
nand U4568 (N_4568,N_4283,N_4126);
nand U4569 (N_4569,N_4417,N_4341);
nor U4570 (N_4570,N_4353,N_4231);
and U4571 (N_4571,N_4053,N_4199);
and U4572 (N_4572,N_4066,N_4148);
or U4573 (N_4573,N_4046,N_4129);
xnor U4574 (N_4574,N_4103,N_4497);
nand U4575 (N_4575,N_4393,N_4104);
nand U4576 (N_4576,N_4369,N_4281);
or U4577 (N_4577,N_4422,N_4123);
or U4578 (N_4578,N_4333,N_4152);
or U4579 (N_4579,N_4346,N_4255);
nand U4580 (N_4580,N_4155,N_4371);
nor U4581 (N_4581,N_4107,N_4017);
and U4582 (N_4582,N_4197,N_4463);
xor U4583 (N_4583,N_4379,N_4016);
and U4584 (N_4584,N_4390,N_4462);
xnor U4585 (N_4585,N_4468,N_4061);
nand U4586 (N_4586,N_4404,N_4498);
and U4587 (N_4587,N_4355,N_4082);
xnor U4588 (N_4588,N_4005,N_4435);
nand U4589 (N_4589,N_4178,N_4090);
nand U4590 (N_4590,N_4034,N_4186);
nand U4591 (N_4591,N_4406,N_4479);
nand U4592 (N_4592,N_4048,N_4068);
nand U4593 (N_4593,N_4009,N_4173);
and U4594 (N_4594,N_4235,N_4314);
nor U4595 (N_4595,N_4297,N_4260);
and U4596 (N_4596,N_4206,N_4365);
or U4597 (N_4597,N_4325,N_4111);
xnor U4598 (N_4598,N_4421,N_4044);
xor U4599 (N_4599,N_4358,N_4003);
nand U4600 (N_4600,N_4030,N_4023);
or U4601 (N_4601,N_4306,N_4183);
nor U4602 (N_4602,N_4316,N_4432);
nor U4603 (N_4603,N_4049,N_4147);
nand U4604 (N_4604,N_4480,N_4405);
or U4605 (N_4605,N_4242,N_4000);
nor U4606 (N_4606,N_4142,N_4444);
and U4607 (N_4607,N_4354,N_4370);
or U4608 (N_4608,N_4488,N_4376);
nor U4609 (N_4609,N_4027,N_4457);
nor U4610 (N_4610,N_4072,N_4403);
xnor U4611 (N_4611,N_4120,N_4425);
xnor U4612 (N_4612,N_4011,N_4496);
nor U4613 (N_4613,N_4201,N_4038);
or U4614 (N_4614,N_4062,N_4060);
nor U4615 (N_4615,N_4088,N_4450);
xnor U4616 (N_4616,N_4211,N_4454);
nor U4617 (N_4617,N_4473,N_4236);
and U4618 (N_4618,N_4109,N_4054);
xor U4619 (N_4619,N_4476,N_4202);
or U4620 (N_4620,N_4431,N_4240);
and U4621 (N_4621,N_4499,N_4485);
or U4622 (N_4622,N_4213,N_4446);
and U4623 (N_4623,N_4483,N_4416);
xnor U4624 (N_4624,N_4311,N_4015);
nor U4625 (N_4625,N_4033,N_4227);
and U4626 (N_4626,N_4338,N_4386);
and U4627 (N_4627,N_4096,N_4336);
or U4628 (N_4628,N_4140,N_4203);
xnor U4629 (N_4629,N_4168,N_4207);
and U4630 (N_4630,N_4149,N_4041);
and U4631 (N_4631,N_4318,N_4050);
and U4632 (N_4632,N_4212,N_4409);
or U4633 (N_4633,N_4351,N_4309);
or U4634 (N_4634,N_4426,N_4289);
nor U4635 (N_4635,N_4436,N_4098);
and U4636 (N_4636,N_4387,N_4170);
xnor U4637 (N_4637,N_4460,N_4051);
xor U4638 (N_4638,N_4055,N_4014);
nand U4639 (N_4639,N_4439,N_4363);
and U4640 (N_4640,N_4071,N_4161);
nand U4641 (N_4641,N_4411,N_4132);
xor U4642 (N_4642,N_4136,N_4441);
or U4643 (N_4643,N_4130,N_4382);
nand U4644 (N_4644,N_4493,N_4368);
xor U4645 (N_4645,N_4205,N_4139);
or U4646 (N_4646,N_4398,N_4218);
and U4647 (N_4647,N_4299,N_4063);
and U4648 (N_4648,N_4128,N_4057);
xnor U4649 (N_4649,N_4134,N_4313);
xor U4650 (N_4650,N_4019,N_4321);
nand U4651 (N_4651,N_4037,N_4418);
and U4652 (N_4652,N_4208,N_4383);
or U4653 (N_4653,N_4189,N_4198);
and U4654 (N_4654,N_4384,N_4176);
nand U4655 (N_4655,N_4429,N_4300);
nand U4656 (N_4656,N_4004,N_4328);
xor U4657 (N_4657,N_4180,N_4097);
and U4658 (N_4658,N_4288,N_4124);
or U4659 (N_4659,N_4002,N_4101);
xor U4660 (N_4660,N_4094,N_4258);
or U4661 (N_4661,N_4308,N_4415);
nand U4662 (N_4662,N_4225,N_4184);
xnor U4663 (N_4663,N_4215,N_4185);
xnor U4664 (N_4664,N_4326,N_4408);
or U4665 (N_4665,N_4492,N_4367);
and U4666 (N_4666,N_4099,N_4165);
nand U4667 (N_4667,N_4167,N_4305);
xor U4668 (N_4668,N_4249,N_4091);
and U4669 (N_4669,N_4026,N_4262);
or U4670 (N_4670,N_4047,N_4226);
or U4671 (N_4671,N_4443,N_4412);
or U4672 (N_4672,N_4145,N_4319);
nor U4673 (N_4673,N_4076,N_4360);
nor U4674 (N_4674,N_4484,N_4270);
nand U4675 (N_4675,N_4056,N_4059);
and U4676 (N_4676,N_4273,N_4430);
nor U4677 (N_4677,N_4086,N_4452);
nand U4678 (N_4678,N_4263,N_4293);
and U4679 (N_4679,N_4008,N_4357);
nand U4680 (N_4680,N_4162,N_4217);
nand U4681 (N_4681,N_4304,N_4447);
nand U4682 (N_4682,N_4095,N_4191);
nor U4683 (N_4683,N_4337,N_4083);
or U4684 (N_4684,N_4486,N_4010);
nand U4685 (N_4685,N_4303,N_4433);
nand U4686 (N_4686,N_4058,N_4194);
xor U4687 (N_4687,N_4464,N_4013);
nor U4688 (N_4688,N_4481,N_4285);
xor U4689 (N_4689,N_4335,N_4381);
nand U4690 (N_4690,N_4233,N_4413);
or U4691 (N_4691,N_4192,N_4018);
or U4692 (N_4692,N_4150,N_4115);
or U4693 (N_4693,N_4110,N_4146);
and U4694 (N_4694,N_4423,N_4307);
and U4695 (N_4695,N_4343,N_4172);
and U4696 (N_4696,N_4223,N_4377);
xor U4697 (N_4697,N_4279,N_4324);
and U4698 (N_4698,N_4356,N_4216);
nor U4699 (N_4699,N_4141,N_4042);
and U4700 (N_4700,N_4117,N_4244);
nor U4701 (N_4701,N_4156,N_4474);
nand U4702 (N_4702,N_4085,N_4074);
nor U4703 (N_4703,N_4272,N_4092);
or U4704 (N_4704,N_4106,N_4153);
or U4705 (N_4705,N_4456,N_4160);
and U4706 (N_4706,N_4410,N_4228);
and U4707 (N_4707,N_4252,N_4310);
or U4708 (N_4708,N_4291,N_4112);
and U4709 (N_4709,N_4108,N_4312);
and U4710 (N_4710,N_4035,N_4375);
and U4711 (N_4711,N_4261,N_4298);
xor U4712 (N_4712,N_4089,N_4445);
nand U4713 (N_4713,N_4073,N_4012);
xor U4714 (N_4714,N_4159,N_4079);
and U4715 (N_4715,N_4006,N_4322);
nand U4716 (N_4716,N_4204,N_4442);
xnor U4717 (N_4717,N_4222,N_4257);
nand U4718 (N_4718,N_4214,N_4093);
and U4719 (N_4719,N_4177,N_4296);
nand U4720 (N_4720,N_4116,N_4402);
or U4721 (N_4721,N_4248,N_4347);
nand U4722 (N_4722,N_4282,N_4349);
nand U4723 (N_4723,N_4339,N_4187);
nand U4724 (N_4724,N_4243,N_4342);
xor U4725 (N_4725,N_4163,N_4234);
nand U4726 (N_4726,N_4482,N_4174);
and U4727 (N_4727,N_4040,N_4295);
nand U4728 (N_4728,N_4399,N_4373);
or U4729 (N_4729,N_4158,N_4119);
nand U4730 (N_4730,N_4237,N_4264);
nand U4731 (N_4731,N_4143,N_4451);
nand U4732 (N_4732,N_4440,N_4100);
nand U4733 (N_4733,N_4323,N_4395);
nor U4734 (N_4734,N_4164,N_4438);
nor U4735 (N_4735,N_4427,N_4219);
nand U4736 (N_4736,N_4069,N_4031);
or U4737 (N_4737,N_4105,N_4275);
nand U4738 (N_4738,N_4352,N_4350);
nor U4739 (N_4739,N_4081,N_4171);
and U4740 (N_4740,N_4271,N_4210);
nor U4741 (N_4741,N_4064,N_4182);
and U4742 (N_4742,N_4453,N_4448);
nor U4743 (N_4743,N_4067,N_4471);
xnor U4744 (N_4744,N_4469,N_4220);
xnor U4745 (N_4745,N_4389,N_4317);
or U4746 (N_4746,N_4458,N_4247);
and U4747 (N_4747,N_4392,N_4131);
xor U4748 (N_4748,N_4477,N_4169);
nand U4749 (N_4749,N_4029,N_4209);
and U4750 (N_4750,N_4312,N_4365);
or U4751 (N_4751,N_4107,N_4082);
xnor U4752 (N_4752,N_4019,N_4141);
and U4753 (N_4753,N_4286,N_4125);
xnor U4754 (N_4754,N_4444,N_4030);
xor U4755 (N_4755,N_4090,N_4205);
or U4756 (N_4756,N_4103,N_4029);
nor U4757 (N_4757,N_4062,N_4122);
nand U4758 (N_4758,N_4149,N_4264);
or U4759 (N_4759,N_4251,N_4496);
nor U4760 (N_4760,N_4496,N_4346);
nand U4761 (N_4761,N_4279,N_4328);
or U4762 (N_4762,N_4220,N_4105);
and U4763 (N_4763,N_4499,N_4008);
nand U4764 (N_4764,N_4082,N_4087);
nand U4765 (N_4765,N_4446,N_4031);
or U4766 (N_4766,N_4038,N_4224);
xor U4767 (N_4767,N_4233,N_4062);
or U4768 (N_4768,N_4480,N_4207);
xor U4769 (N_4769,N_4462,N_4119);
or U4770 (N_4770,N_4139,N_4288);
and U4771 (N_4771,N_4439,N_4383);
nand U4772 (N_4772,N_4150,N_4323);
xor U4773 (N_4773,N_4303,N_4178);
nor U4774 (N_4774,N_4470,N_4477);
nor U4775 (N_4775,N_4458,N_4310);
nand U4776 (N_4776,N_4096,N_4461);
nand U4777 (N_4777,N_4438,N_4235);
or U4778 (N_4778,N_4032,N_4430);
nand U4779 (N_4779,N_4416,N_4496);
nor U4780 (N_4780,N_4362,N_4492);
nand U4781 (N_4781,N_4187,N_4477);
or U4782 (N_4782,N_4011,N_4376);
or U4783 (N_4783,N_4214,N_4084);
nand U4784 (N_4784,N_4469,N_4129);
and U4785 (N_4785,N_4087,N_4405);
xor U4786 (N_4786,N_4466,N_4150);
nor U4787 (N_4787,N_4491,N_4016);
or U4788 (N_4788,N_4333,N_4206);
nor U4789 (N_4789,N_4188,N_4226);
nand U4790 (N_4790,N_4431,N_4151);
nor U4791 (N_4791,N_4211,N_4214);
nor U4792 (N_4792,N_4381,N_4113);
and U4793 (N_4793,N_4224,N_4344);
nor U4794 (N_4794,N_4450,N_4068);
and U4795 (N_4795,N_4405,N_4225);
and U4796 (N_4796,N_4494,N_4387);
nor U4797 (N_4797,N_4368,N_4356);
or U4798 (N_4798,N_4311,N_4477);
and U4799 (N_4799,N_4153,N_4375);
nand U4800 (N_4800,N_4266,N_4071);
or U4801 (N_4801,N_4166,N_4172);
xor U4802 (N_4802,N_4167,N_4365);
or U4803 (N_4803,N_4247,N_4249);
nor U4804 (N_4804,N_4264,N_4250);
nor U4805 (N_4805,N_4259,N_4255);
nor U4806 (N_4806,N_4106,N_4334);
or U4807 (N_4807,N_4175,N_4154);
xor U4808 (N_4808,N_4286,N_4051);
and U4809 (N_4809,N_4327,N_4061);
xor U4810 (N_4810,N_4129,N_4340);
and U4811 (N_4811,N_4481,N_4495);
nor U4812 (N_4812,N_4124,N_4406);
and U4813 (N_4813,N_4369,N_4450);
or U4814 (N_4814,N_4414,N_4231);
and U4815 (N_4815,N_4173,N_4330);
nor U4816 (N_4816,N_4356,N_4318);
and U4817 (N_4817,N_4294,N_4199);
or U4818 (N_4818,N_4157,N_4444);
nand U4819 (N_4819,N_4204,N_4378);
nand U4820 (N_4820,N_4493,N_4201);
nor U4821 (N_4821,N_4030,N_4403);
nor U4822 (N_4822,N_4387,N_4067);
or U4823 (N_4823,N_4085,N_4353);
xor U4824 (N_4824,N_4422,N_4082);
and U4825 (N_4825,N_4023,N_4206);
and U4826 (N_4826,N_4108,N_4430);
and U4827 (N_4827,N_4007,N_4151);
xnor U4828 (N_4828,N_4185,N_4262);
nor U4829 (N_4829,N_4075,N_4056);
xor U4830 (N_4830,N_4459,N_4238);
xnor U4831 (N_4831,N_4018,N_4156);
nor U4832 (N_4832,N_4461,N_4064);
and U4833 (N_4833,N_4203,N_4239);
and U4834 (N_4834,N_4093,N_4097);
nor U4835 (N_4835,N_4475,N_4077);
xnor U4836 (N_4836,N_4440,N_4341);
or U4837 (N_4837,N_4322,N_4091);
or U4838 (N_4838,N_4297,N_4412);
and U4839 (N_4839,N_4049,N_4463);
or U4840 (N_4840,N_4382,N_4027);
nand U4841 (N_4841,N_4407,N_4432);
or U4842 (N_4842,N_4138,N_4286);
nand U4843 (N_4843,N_4332,N_4094);
or U4844 (N_4844,N_4088,N_4366);
and U4845 (N_4845,N_4240,N_4341);
xor U4846 (N_4846,N_4455,N_4458);
xor U4847 (N_4847,N_4453,N_4057);
xnor U4848 (N_4848,N_4478,N_4366);
nand U4849 (N_4849,N_4357,N_4024);
xnor U4850 (N_4850,N_4454,N_4276);
xor U4851 (N_4851,N_4450,N_4431);
nor U4852 (N_4852,N_4200,N_4346);
nor U4853 (N_4853,N_4461,N_4307);
and U4854 (N_4854,N_4058,N_4167);
nand U4855 (N_4855,N_4434,N_4397);
or U4856 (N_4856,N_4484,N_4321);
or U4857 (N_4857,N_4089,N_4309);
or U4858 (N_4858,N_4083,N_4080);
and U4859 (N_4859,N_4361,N_4138);
or U4860 (N_4860,N_4339,N_4348);
nand U4861 (N_4861,N_4010,N_4101);
nor U4862 (N_4862,N_4395,N_4390);
and U4863 (N_4863,N_4067,N_4461);
xnor U4864 (N_4864,N_4238,N_4117);
nor U4865 (N_4865,N_4143,N_4446);
nand U4866 (N_4866,N_4280,N_4142);
or U4867 (N_4867,N_4072,N_4336);
and U4868 (N_4868,N_4241,N_4354);
nand U4869 (N_4869,N_4311,N_4226);
xnor U4870 (N_4870,N_4489,N_4267);
nand U4871 (N_4871,N_4430,N_4384);
and U4872 (N_4872,N_4158,N_4360);
xnor U4873 (N_4873,N_4340,N_4039);
or U4874 (N_4874,N_4038,N_4187);
or U4875 (N_4875,N_4036,N_4204);
nand U4876 (N_4876,N_4453,N_4441);
or U4877 (N_4877,N_4410,N_4442);
or U4878 (N_4878,N_4104,N_4466);
and U4879 (N_4879,N_4270,N_4316);
nor U4880 (N_4880,N_4325,N_4490);
and U4881 (N_4881,N_4133,N_4014);
xor U4882 (N_4882,N_4399,N_4278);
nor U4883 (N_4883,N_4142,N_4211);
nand U4884 (N_4884,N_4312,N_4263);
xor U4885 (N_4885,N_4179,N_4034);
or U4886 (N_4886,N_4126,N_4419);
nand U4887 (N_4887,N_4209,N_4464);
nor U4888 (N_4888,N_4051,N_4442);
and U4889 (N_4889,N_4476,N_4221);
nor U4890 (N_4890,N_4338,N_4365);
xnor U4891 (N_4891,N_4466,N_4438);
and U4892 (N_4892,N_4078,N_4405);
and U4893 (N_4893,N_4419,N_4130);
nor U4894 (N_4894,N_4439,N_4267);
or U4895 (N_4895,N_4291,N_4399);
or U4896 (N_4896,N_4084,N_4436);
xnor U4897 (N_4897,N_4038,N_4177);
nor U4898 (N_4898,N_4466,N_4430);
xnor U4899 (N_4899,N_4183,N_4099);
nand U4900 (N_4900,N_4026,N_4486);
xor U4901 (N_4901,N_4151,N_4444);
nor U4902 (N_4902,N_4094,N_4139);
or U4903 (N_4903,N_4356,N_4076);
nand U4904 (N_4904,N_4104,N_4229);
nand U4905 (N_4905,N_4451,N_4183);
and U4906 (N_4906,N_4476,N_4423);
nor U4907 (N_4907,N_4444,N_4014);
and U4908 (N_4908,N_4061,N_4141);
or U4909 (N_4909,N_4025,N_4398);
xor U4910 (N_4910,N_4201,N_4155);
and U4911 (N_4911,N_4109,N_4433);
nand U4912 (N_4912,N_4279,N_4189);
or U4913 (N_4913,N_4185,N_4444);
xor U4914 (N_4914,N_4288,N_4310);
and U4915 (N_4915,N_4358,N_4216);
nor U4916 (N_4916,N_4169,N_4325);
nand U4917 (N_4917,N_4494,N_4257);
and U4918 (N_4918,N_4381,N_4001);
and U4919 (N_4919,N_4432,N_4308);
nor U4920 (N_4920,N_4495,N_4452);
or U4921 (N_4921,N_4285,N_4453);
or U4922 (N_4922,N_4058,N_4155);
nor U4923 (N_4923,N_4141,N_4480);
nor U4924 (N_4924,N_4375,N_4104);
and U4925 (N_4925,N_4357,N_4095);
xnor U4926 (N_4926,N_4323,N_4160);
nand U4927 (N_4927,N_4253,N_4050);
nor U4928 (N_4928,N_4085,N_4162);
xnor U4929 (N_4929,N_4054,N_4208);
or U4930 (N_4930,N_4010,N_4144);
nand U4931 (N_4931,N_4266,N_4190);
and U4932 (N_4932,N_4412,N_4089);
nand U4933 (N_4933,N_4178,N_4323);
or U4934 (N_4934,N_4246,N_4096);
and U4935 (N_4935,N_4158,N_4285);
and U4936 (N_4936,N_4038,N_4393);
xor U4937 (N_4937,N_4073,N_4440);
nor U4938 (N_4938,N_4165,N_4002);
nand U4939 (N_4939,N_4456,N_4448);
and U4940 (N_4940,N_4305,N_4387);
or U4941 (N_4941,N_4466,N_4122);
or U4942 (N_4942,N_4101,N_4400);
xnor U4943 (N_4943,N_4379,N_4295);
and U4944 (N_4944,N_4170,N_4311);
or U4945 (N_4945,N_4092,N_4373);
nand U4946 (N_4946,N_4213,N_4373);
xnor U4947 (N_4947,N_4288,N_4145);
or U4948 (N_4948,N_4253,N_4197);
nor U4949 (N_4949,N_4013,N_4101);
nand U4950 (N_4950,N_4270,N_4364);
and U4951 (N_4951,N_4272,N_4384);
and U4952 (N_4952,N_4135,N_4088);
or U4953 (N_4953,N_4052,N_4427);
and U4954 (N_4954,N_4489,N_4269);
nor U4955 (N_4955,N_4406,N_4472);
and U4956 (N_4956,N_4422,N_4427);
nand U4957 (N_4957,N_4139,N_4321);
nor U4958 (N_4958,N_4153,N_4324);
nand U4959 (N_4959,N_4095,N_4249);
xnor U4960 (N_4960,N_4205,N_4259);
and U4961 (N_4961,N_4170,N_4314);
xor U4962 (N_4962,N_4303,N_4358);
nand U4963 (N_4963,N_4423,N_4181);
xnor U4964 (N_4964,N_4219,N_4014);
or U4965 (N_4965,N_4059,N_4025);
xor U4966 (N_4966,N_4117,N_4090);
xnor U4967 (N_4967,N_4159,N_4196);
or U4968 (N_4968,N_4124,N_4303);
xnor U4969 (N_4969,N_4112,N_4166);
or U4970 (N_4970,N_4337,N_4300);
or U4971 (N_4971,N_4057,N_4242);
or U4972 (N_4972,N_4194,N_4176);
nor U4973 (N_4973,N_4175,N_4219);
or U4974 (N_4974,N_4409,N_4116);
nand U4975 (N_4975,N_4017,N_4340);
xor U4976 (N_4976,N_4370,N_4394);
nor U4977 (N_4977,N_4144,N_4322);
xnor U4978 (N_4978,N_4089,N_4429);
xor U4979 (N_4979,N_4025,N_4237);
nor U4980 (N_4980,N_4443,N_4452);
and U4981 (N_4981,N_4333,N_4008);
nor U4982 (N_4982,N_4012,N_4196);
nor U4983 (N_4983,N_4019,N_4144);
and U4984 (N_4984,N_4060,N_4067);
xnor U4985 (N_4985,N_4465,N_4486);
nand U4986 (N_4986,N_4453,N_4384);
nor U4987 (N_4987,N_4094,N_4005);
xor U4988 (N_4988,N_4186,N_4057);
xor U4989 (N_4989,N_4231,N_4018);
or U4990 (N_4990,N_4222,N_4237);
nor U4991 (N_4991,N_4285,N_4484);
nand U4992 (N_4992,N_4068,N_4015);
or U4993 (N_4993,N_4238,N_4249);
and U4994 (N_4994,N_4157,N_4236);
or U4995 (N_4995,N_4337,N_4173);
nor U4996 (N_4996,N_4201,N_4435);
and U4997 (N_4997,N_4208,N_4076);
nand U4998 (N_4998,N_4338,N_4102);
nor U4999 (N_4999,N_4437,N_4398);
nor U5000 (N_5000,N_4606,N_4557);
and U5001 (N_5001,N_4724,N_4643);
xnor U5002 (N_5002,N_4753,N_4586);
nand U5003 (N_5003,N_4978,N_4782);
nor U5004 (N_5004,N_4936,N_4554);
nand U5005 (N_5005,N_4989,N_4892);
and U5006 (N_5006,N_4846,N_4979);
nor U5007 (N_5007,N_4534,N_4904);
nor U5008 (N_5008,N_4794,N_4925);
nor U5009 (N_5009,N_4560,N_4821);
xnor U5010 (N_5010,N_4746,N_4877);
and U5011 (N_5011,N_4768,N_4897);
and U5012 (N_5012,N_4712,N_4820);
or U5013 (N_5013,N_4668,N_4720);
nor U5014 (N_5014,N_4818,N_4604);
or U5015 (N_5015,N_4515,N_4552);
nand U5016 (N_5016,N_4541,N_4881);
nor U5017 (N_5017,N_4832,N_4628);
nor U5018 (N_5018,N_4775,N_4690);
or U5019 (N_5019,N_4784,N_4520);
nor U5020 (N_5020,N_4933,N_4975);
nand U5021 (N_5021,N_4519,N_4516);
nor U5022 (N_5022,N_4537,N_4996);
nor U5023 (N_5023,N_4607,N_4710);
xnor U5024 (N_5024,N_4596,N_4658);
or U5025 (N_5025,N_4684,N_4635);
nor U5026 (N_5026,N_4632,N_4859);
nor U5027 (N_5027,N_4957,N_4953);
nand U5028 (N_5028,N_4540,N_4647);
or U5029 (N_5029,N_4807,N_4799);
or U5030 (N_5030,N_4808,N_4886);
and U5031 (N_5031,N_4717,N_4816);
or U5032 (N_5032,N_4719,N_4793);
or U5033 (N_5033,N_4714,N_4967);
and U5034 (N_5034,N_4751,N_4815);
or U5035 (N_5035,N_4650,N_4580);
nor U5036 (N_5036,N_4899,N_4599);
and U5037 (N_5037,N_4943,N_4698);
or U5038 (N_5038,N_4913,N_4814);
and U5039 (N_5039,N_4907,N_4765);
and U5040 (N_5040,N_4574,N_4518);
xor U5041 (N_5041,N_4842,N_4863);
nor U5042 (N_5042,N_4920,N_4506);
xor U5043 (N_5043,N_4721,N_4940);
and U5044 (N_5044,N_4976,N_4785);
or U5045 (N_5045,N_4556,N_4734);
xor U5046 (N_5046,N_4740,N_4778);
or U5047 (N_5047,N_4739,N_4622);
nor U5048 (N_5048,N_4876,N_4588);
nand U5049 (N_5049,N_4583,N_4522);
xnor U5050 (N_5050,N_4864,N_4855);
xor U5051 (N_5051,N_4509,N_4745);
or U5052 (N_5052,N_4912,N_4566);
and U5053 (N_5053,N_4969,N_4732);
nand U5054 (N_5054,N_4570,N_4893);
xor U5055 (N_5055,N_4946,N_4743);
xnor U5056 (N_5056,N_4994,N_4601);
nor U5057 (N_5057,N_4590,N_4931);
nor U5058 (N_5058,N_4707,N_4699);
nand U5059 (N_5059,N_4733,N_4619);
nand U5060 (N_5060,N_4795,N_4676);
xnor U5061 (N_5061,N_4910,N_4669);
nand U5062 (N_5062,N_4553,N_4838);
nand U5063 (N_5063,N_4986,N_4981);
or U5064 (N_5064,N_4623,N_4716);
and U5065 (N_5065,N_4626,N_4791);
nand U5066 (N_5066,N_4923,N_4504);
nor U5067 (N_5067,N_4921,N_4835);
or U5068 (N_5068,N_4559,N_4919);
and U5069 (N_5069,N_4510,N_4853);
and U5070 (N_5070,N_4866,N_4589);
nor U5071 (N_5071,N_4900,N_4535);
nor U5072 (N_5072,N_4857,N_4550);
xnor U5073 (N_5073,N_4750,N_4823);
nor U5074 (N_5074,N_4687,N_4639);
or U5075 (N_5075,N_4591,N_4939);
and U5076 (N_5076,N_4871,N_4645);
xor U5077 (N_5077,N_4575,N_4844);
nand U5078 (N_5078,N_4971,N_4651);
and U5079 (N_5079,N_4567,N_4679);
and U5080 (N_5080,N_4674,N_4803);
or U5081 (N_5081,N_4954,N_4972);
nor U5082 (N_5082,N_4705,N_4729);
xnor U5083 (N_5083,N_4621,N_4744);
nor U5084 (N_5084,N_4722,N_4860);
xnor U5085 (N_5085,N_4701,N_4648);
nor U5086 (N_5086,N_4914,N_4505);
and U5087 (N_5087,N_4999,N_4526);
nand U5088 (N_5088,N_4528,N_4598);
xnor U5089 (N_5089,N_4749,N_4761);
and U5090 (N_5090,N_4563,N_4602);
or U5091 (N_5091,N_4875,N_4568);
nor U5092 (N_5092,N_4571,N_4500);
nor U5093 (N_5093,N_4836,N_4896);
nand U5094 (N_5094,N_4547,N_4796);
and U5095 (N_5095,N_4851,N_4608);
or U5096 (N_5096,N_4735,N_4984);
or U5097 (N_5097,N_4883,N_4817);
and U5098 (N_5098,N_4858,N_4810);
nor U5099 (N_5099,N_4538,N_4726);
or U5100 (N_5100,N_4878,N_4507);
and U5101 (N_5101,N_4809,N_4680);
or U5102 (N_5102,N_4891,N_4683);
xnor U5103 (N_5103,N_4661,N_4671);
nand U5104 (N_5104,N_4703,N_4546);
and U5105 (N_5105,N_4675,N_4630);
nand U5106 (N_5106,N_4789,N_4812);
nand U5107 (N_5107,N_4802,N_4828);
and U5108 (N_5108,N_4955,N_4508);
or U5109 (N_5109,N_4764,N_4781);
and U5110 (N_5110,N_4711,N_4523);
and U5111 (N_5111,N_4987,N_4786);
or U5112 (N_5112,N_4531,N_4542);
nand U5113 (N_5113,N_4642,N_4646);
xnor U5114 (N_5114,N_4502,N_4677);
and U5115 (N_5115,N_4682,N_4985);
or U5116 (N_5116,N_4673,N_4543);
or U5117 (N_5117,N_4718,N_4854);
or U5118 (N_5118,N_4941,N_4843);
nand U5119 (N_5119,N_4804,N_4663);
or U5120 (N_5120,N_4991,N_4767);
and U5121 (N_5121,N_4533,N_4728);
nor U5122 (N_5122,N_4551,N_4565);
or U5123 (N_5123,N_4884,N_4655);
and U5124 (N_5124,N_4800,N_4656);
nand U5125 (N_5125,N_4742,N_4937);
or U5126 (N_5126,N_4968,N_4654);
and U5127 (N_5127,N_4613,N_4696);
or U5128 (N_5128,N_4956,N_4766);
nor U5129 (N_5129,N_4944,N_4916);
xnor U5130 (N_5130,N_4770,N_4562);
or U5131 (N_5131,N_4620,N_4529);
nor U5132 (N_5132,N_4527,N_4947);
xor U5133 (N_5133,N_4521,N_4624);
nand U5134 (N_5134,N_4592,N_4911);
or U5135 (N_5135,N_4572,N_4548);
and U5136 (N_5136,N_4597,N_4934);
or U5137 (N_5137,N_4792,N_4805);
nor U5138 (N_5138,N_4888,N_4839);
xor U5139 (N_5139,N_4513,N_4609);
nor U5140 (N_5140,N_4715,N_4530);
nand U5141 (N_5141,N_4983,N_4688);
and U5142 (N_5142,N_4640,N_4852);
or U5143 (N_5143,N_4737,N_4889);
or U5144 (N_5144,N_4617,N_4625);
nor U5145 (N_5145,N_4961,N_4549);
and U5146 (N_5146,N_4774,N_4880);
xnor U5147 (N_5147,N_4992,N_4723);
and U5148 (N_5148,N_4569,N_4948);
and U5149 (N_5149,N_4539,N_4694);
xnor U5150 (N_5150,N_4762,N_4702);
or U5151 (N_5151,N_4906,N_4747);
xnor U5152 (N_5152,N_4993,N_4678);
or U5153 (N_5153,N_4874,N_4659);
nor U5154 (N_5154,N_4612,N_4926);
or U5155 (N_5155,N_4605,N_4790);
xnor U5156 (N_5156,N_4706,N_4869);
nor U5157 (N_5157,N_4657,N_4930);
or U5158 (N_5158,N_4833,N_4771);
nor U5159 (N_5159,N_4966,N_4872);
or U5160 (N_5160,N_4890,N_4545);
or U5161 (N_5161,N_4564,N_4801);
nand U5162 (N_5162,N_4798,N_4660);
or U5163 (N_5163,N_4614,N_4780);
xor U5164 (N_5164,N_4631,N_4561);
xnor U5165 (N_5165,N_4511,N_4665);
or U5166 (N_5166,N_4995,N_4756);
nor U5167 (N_5167,N_4662,N_4901);
nand U5168 (N_5168,N_4629,N_4555);
nor U5169 (N_5169,N_4962,N_4887);
or U5170 (N_5170,N_4587,N_4709);
nor U5171 (N_5171,N_4963,N_4776);
xnor U5172 (N_5172,N_4693,N_4917);
nand U5173 (N_5173,N_4932,N_4725);
nor U5174 (N_5174,N_4870,N_4637);
nor U5175 (N_5175,N_4600,N_4686);
xnor U5176 (N_5176,N_4970,N_4865);
nand U5177 (N_5177,N_4514,N_4848);
xor U5178 (N_5178,N_4692,N_4819);
xnor U5179 (N_5179,N_4670,N_4806);
xnor U5180 (N_5180,N_4689,N_4627);
or U5181 (N_5181,N_4708,N_4672);
and U5182 (N_5182,N_4649,N_4691);
and U5183 (N_5183,N_4695,N_4980);
xor U5184 (N_5184,N_4831,N_4856);
or U5185 (N_5185,N_4731,N_4952);
xnor U5186 (N_5186,N_4681,N_4641);
or U5187 (N_5187,N_4964,N_4634);
and U5188 (N_5188,N_4501,N_4697);
nand U5189 (N_5189,N_4595,N_4861);
nand U5190 (N_5190,N_4763,N_4700);
nand U5191 (N_5191,N_4945,N_4951);
nor U5192 (N_5192,N_4594,N_4584);
and U5193 (N_5193,N_4990,N_4997);
xnor U5194 (N_5194,N_4847,N_4593);
nand U5195 (N_5195,N_4950,N_4895);
nand U5196 (N_5196,N_4615,N_4811);
xnor U5197 (N_5197,N_4636,N_4576);
nand U5198 (N_5198,N_4611,N_4908);
xor U5199 (N_5199,N_4827,N_4524);
nand U5200 (N_5200,N_4736,N_4845);
nand U5201 (N_5201,N_4942,N_4758);
xor U5202 (N_5202,N_4777,N_4965);
and U5203 (N_5203,N_4824,N_4525);
or U5204 (N_5204,N_4582,N_4924);
nand U5205 (N_5205,N_4653,N_4929);
nand U5206 (N_5206,N_4652,N_4579);
nand U5207 (N_5207,N_4894,N_4503);
and U5208 (N_5208,N_4581,N_4713);
and U5209 (N_5209,N_4915,N_4935);
nand U5210 (N_5210,N_4837,N_4850);
or U5211 (N_5211,N_4664,N_4960);
nand U5212 (N_5212,N_4769,N_4873);
nor U5213 (N_5213,N_4829,N_4813);
xor U5214 (N_5214,N_4759,N_4902);
or U5215 (N_5215,N_4685,N_4959);
xor U5216 (N_5216,N_4644,N_4666);
nor U5217 (N_5217,N_4949,N_4773);
nor U5218 (N_5218,N_4862,N_4974);
nor U5219 (N_5219,N_4879,N_4822);
nand U5220 (N_5220,N_4973,N_4573);
and U5221 (N_5221,N_4841,N_4928);
xnor U5222 (N_5222,N_4977,N_4885);
nor U5223 (N_5223,N_4849,N_4760);
nor U5224 (N_5224,N_4536,N_4834);
xor U5225 (N_5225,N_4603,N_4638);
or U5226 (N_5226,N_4905,N_4741);
or U5227 (N_5227,N_4610,N_4585);
nand U5228 (N_5228,N_4667,N_4797);
nand U5229 (N_5229,N_4922,N_4788);
and U5230 (N_5230,N_4633,N_4730);
nand U5231 (N_5231,N_4772,N_4958);
nor U5232 (N_5232,N_4988,N_4577);
or U5233 (N_5233,N_4909,N_4618);
xor U5234 (N_5234,N_4754,N_4578);
nor U5235 (N_5235,N_4898,N_4918);
or U5236 (N_5236,N_4826,N_4938);
or U5237 (N_5237,N_4738,N_4927);
nor U5238 (N_5238,N_4830,N_4748);
nand U5239 (N_5239,N_4517,N_4882);
nand U5240 (N_5240,N_4868,N_4752);
nor U5241 (N_5241,N_4998,N_4512);
or U5242 (N_5242,N_4755,N_4727);
nor U5243 (N_5243,N_4704,N_4787);
nor U5244 (N_5244,N_4903,N_4867);
nand U5245 (N_5245,N_4558,N_4783);
xnor U5246 (N_5246,N_4757,N_4840);
xor U5247 (N_5247,N_4532,N_4616);
nor U5248 (N_5248,N_4779,N_4544);
nand U5249 (N_5249,N_4982,N_4825);
xnor U5250 (N_5250,N_4505,N_4649);
xor U5251 (N_5251,N_4585,N_4928);
nand U5252 (N_5252,N_4502,N_4938);
nor U5253 (N_5253,N_4833,N_4957);
nand U5254 (N_5254,N_4634,N_4751);
and U5255 (N_5255,N_4944,N_4921);
nor U5256 (N_5256,N_4696,N_4596);
xnor U5257 (N_5257,N_4934,N_4641);
nand U5258 (N_5258,N_4991,N_4774);
or U5259 (N_5259,N_4517,N_4644);
xor U5260 (N_5260,N_4623,N_4781);
or U5261 (N_5261,N_4693,N_4829);
or U5262 (N_5262,N_4616,N_4526);
nor U5263 (N_5263,N_4517,N_4858);
or U5264 (N_5264,N_4857,N_4682);
or U5265 (N_5265,N_4913,N_4787);
xor U5266 (N_5266,N_4929,N_4735);
xor U5267 (N_5267,N_4595,N_4667);
and U5268 (N_5268,N_4620,N_4778);
and U5269 (N_5269,N_4922,N_4929);
nor U5270 (N_5270,N_4601,N_4517);
xor U5271 (N_5271,N_4910,N_4556);
xnor U5272 (N_5272,N_4816,N_4964);
or U5273 (N_5273,N_4564,N_4947);
xor U5274 (N_5274,N_4584,N_4940);
nand U5275 (N_5275,N_4974,N_4853);
and U5276 (N_5276,N_4851,N_4729);
and U5277 (N_5277,N_4504,N_4619);
nor U5278 (N_5278,N_4752,N_4953);
nor U5279 (N_5279,N_4681,N_4922);
or U5280 (N_5280,N_4590,N_4752);
xnor U5281 (N_5281,N_4858,N_4851);
nor U5282 (N_5282,N_4721,N_4556);
or U5283 (N_5283,N_4719,N_4888);
xor U5284 (N_5284,N_4896,N_4663);
xnor U5285 (N_5285,N_4649,N_4573);
nand U5286 (N_5286,N_4663,N_4915);
nor U5287 (N_5287,N_4629,N_4675);
or U5288 (N_5288,N_4695,N_4629);
nand U5289 (N_5289,N_4580,N_4982);
nand U5290 (N_5290,N_4847,N_4864);
xnor U5291 (N_5291,N_4831,N_4636);
or U5292 (N_5292,N_4957,N_4783);
xor U5293 (N_5293,N_4955,N_4877);
nand U5294 (N_5294,N_4823,N_4594);
nand U5295 (N_5295,N_4628,N_4947);
nand U5296 (N_5296,N_4615,N_4568);
and U5297 (N_5297,N_4536,N_4981);
nand U5298 (N_5298,N_4908,N_4606);
xor U5299 (N_5299,N_4774,N_4922);
nand U5300 (N_5300,N_4744,N_4558);
and U5301 (N_5301,N_4678,N_4741);
xor U5302 (N_5302,N_4554,N_4786);
nand U5303 (N_5303,N_4693,N_4834);
or U5304 (N_5304,N_4531,N_4977);
nor U5305 (N_5305,N_4919,N_4804);
or U5306 (N_5306,N_4584,N_4629);
nor U5307 (N_5307,N_4720,N_4900);
or U5308 (N_5308,N_4685,N_4724);
xor U5309 (N_5309,N_4675,N_4517);
or U5310 (N_5310,N_4791,N_4862);
xor U5311 (N_5311,N_4938,N_4854);
nor U5312 (N_5312,N_4576,N_4824);
xor U5313 (N_5313,N_4968,N_4924);
and U5314 (N_5314,N_4528,N_4956);
or U5315 (N_5315,N_4902,N_4876);
nor U5316 (N_5316,N_4999,N_4993);
xor U5317 (N_5317,N_4920,N_4646);
or U5318 (N_5318,N_4908,N_4619);
or U5319 (N_5319,N_4604,N_4556);
or U5320 (N_5320,N_4680,N_4819);
and U5321 (N_5321,N_4992,N_4932);
or U5322 (N_5322,N_4984,N_4516);
xnor U5323 (N_5323,N_4597,N_4886);
nor U5324 (N_5324,N_4585,N_4612);
and U5325 (N_5325,N_4609,N_4598);
or U5326 (N_5326,N_4602,N_4680);
and U5327 (N_5327,N_4726,N_4642);
nor U5328 (N_5328,N_4736,N_4518);
and U5329 (N_5329,N_4704,N_4872);
or U5330 (N_5330,N_4628,N_4617);
nor U5331 (N_5331,N_4624,N_4535);
and U5332 (N_5332,N_4537,N_4890);
xor U5333 (N_5333,N_4700,N_4751);
and U5334 (N_5334,N_4514,N_4839);
nor U5335 (N_5335,N_4764,N_4520);
and U5336 (N_5336,N_4888,N_4964);
nor U5337 (N_5337,N_4946,N_4582);
xnor U5338 (N_5338,N_4671,N_4789);
or U5339 (N_5339,N_4703,N_4567);
or U5340 (N_5340,N_4822,N_4706);
or U5341 (N_5341,N_4825,N_4947);
or U5342 (N_5342,N_4999,N_4664);
xnor U5343 (N_5343,N_4806,N_4857);
and U5344 (N_5344,N_4510,N_4664);
nor U5345 (N_5345,N_4893,N_4723);
nor U5346 (N_5346,N_4992,N_4964);
nor U5347 (N_5347,N_4644,N_4565);
or U5348 (N_5348,N_4634,N_4965);
nand U5349 (N_5349,N_4778,N_4855);
xor U5350 (N_5350,N_4970,N_4815);
and U5351 (N_5351,N_4913,N_4736);
nor U5352 (N_5352,N_4597,N_4684);
xnor U5353 (N_5353,N_4551,N_4922);
xor U5354 (N_5354,N_4762,N_4565);
nand U5355 (N_5355,N_4552,N_4935);
or U5356 (N_5356,N_4749,N_4977);
or U5357 (N_5357,N_4519,N_4668);
nand U5358 (N_5358,N_4821,N_4931);
and U5359 (N_5359,N_4610,N_4675);
nor U5360 (N_5360,N_4795,N_4978);
or U5361 (N_5361,N_4677,N_4528);
and U5362 (N_5362,N_4678,N_4649);
nor U5363 (N_5363,N_4996,N_4504);
xor U5364 (N_5364,N_4856,N_4623);
xnor U5365 (N_5365,N_4581,N_4886);
nor U5366 (N_5366,N_4901,N_4669);
nand U5367 (N_5367,N_4803,N_4810);
nor U5368 (N_5368,N_4632,N_4892);
nor U5369 (N_5369,N_4963,N_4608);
or U5370 (N_5370,N_4813,N_4766);
or U5371 (N_5371,N_4707,N_4574);
nor U5372 (N_5372,N_4551,N_4661);
nand U5373 (N_5373,N_4596,N_4868);
nand U5374 (N_5374,N_4578,N_4847);
xnor U5375 (N_5375,N_4645,N_4608);
xnor U5376 (N_5376,N_4562,N_4918);
or U5377 (N_5377,N_4899,N_4789);
xnor U5378 (N_5378,N_4760,N_4500);
xor U5379 (N_5379,N_4698,N_4681);
nand U5380 (N_5380,N_4621,N_4523);
nor U5381 (N_5381,N_4926,N_4560);
nor U5382 (N_5382,N_4818,N_4830);
and U5383 (N_5383,N_4655,N_4974);
nor U5384 (N_5384,N_4946,N_4599);
or U5385 (N_5385,N_4511,N_4849);
nor U5386 (N_5386,N_4530,N_4978);
nand U5387 (N_5387,N_4657,N_4729);
xor U5388 (N_5388,N_4729,N_4689);
nand U5389 (N_5389,N_4724,N_4623);
nand U5390 (N_5390,N_4758,N_4995);
nor U5391 (N_5391,N_4816,N_4577);
xor U5392 (N_5392,N_4989,N_4703);
and U5393 (N_5393,N_4617,N_4522);
and U5394 (N_5394,N_4934,N_4662);
and U5395 (N_5395,N_4834,N_4868);
xor U5396 (N_5396,N_4760,N_4698);
or U5397 (N_5397,N_4547,N_4742);
and U5398 (N_5398,N_4936,N_4631);
and U5399 (N_5399,N_4586,N_4515);
nand U5400 (N_5400,N_4813,N_4978);
and U5401 (N_5401,N_4808,N_4550);
nand U5402 (N_5402,N_4825,N_4852);
and U5403 (N_5403,N_4954,N_4824);
or U5404 (N_5404,N_4786,N_4581);
nor U5405 (N_5405,N_4862,N_4980);
nor U5406 (N_5406,N_4648,N_4956);
nor U5407 (N_5407,N_4828,N_4749);
or U5408 (N_5408,N_4772,N_4512);
nor U5409 (N_5409,N_4953,N_4787);
xor U5410 (N_5410,N_4513,N_4724);
nor U5411 (N_5411,N_4717,N_4851);
xnor U5412 (N_5412,N_4641,N_4968);
xnor U5413 (N_5413,N_4513,N_4686);
xnor U5414 (N_5414,N_4832,N_4769);
or U5415 (N_5415,N_4979,N_4862);
and U5416 (N_5416,N_4757,N_4786);
or U5417 (N_5417,N_4734,N_4862);
nor U5418 (N_5418,N_4665,N_4845);
nor U5419 (N_5419,N_4531,N_4699);
nor U5420 (N_5420,N_4962,N_4579);
and U5421 (N_5421,N_4745,N_4653);
nand U5422 (N_5422,N_4991,N_4919);
xnor U5423 (N_5423,N_4862,N_4825);
or U5424 (N_5424,N_4803,N_4745);
nand U5425 (N_5425,N_4889,N_4501);
or U5426 (N_5426,N_4933,N_4747);
nor U5427 (N_5427,N_4593,N_4911);
or U5428 (N_5428,N_4834,N_4639);
nand U5429 (N_5429,N_4986,N_4761);
nor U5430 (N_5430,N_4873,N_4871);
or U5431 (N_5431,N_4562,N_4787);
nand U5432 (N_5432,N_4705,N_4617);
nor U5433 (N_5433,N_4750,N_4968);
nand U5434 (N_5434,N_4575,N_4790);
nand U5435 (N_5435,N_4687,N_4788);
or U5436 (N_5436,N_4707,N_4927);
xnor U5437 (N_5437,N_4576,N_4801);
or U5438 (N_5438,N_4807,N_4630);
and U5439 (N_5439,N_4874,N_4855);
nand U5440 (N_5440,N_4906,N_4976);
nand U5441 (N_5441,N_4821,N_4549);
or U5442 (N_5442,N_4657,N_4944);
and U5443 (N_5443,N_4634,N_4799);
xnor U5444 (N_5444,N_4964,N_4972);
and U5445 (N_5445,N_4703,N_4956);
nor U5446 (N_5446,N_4837,N_4677);
or U5447 (N_5447,N_4778,N_4944);
nand U5448 (N_5448,N_4528,N_4622);
and U5449 (N_5449,N_4657,N_4523);
nor U5450 (N_5450,N_4917,N_4722);
nand U5451 (N_5451,N_4520,N_4878);
xor U5452 (N_5452,N_4657,N_4785);
nor U5453 (N_5453,N_4861,N_4820);
and U5454 (N_5454,N_4679,N_4889);
xnor U5455 (N_5455,N_4650,N_4585);
xor U5456 (N_5456,N_4717,N_4679);
xor U5457 (N_5457,N_4725,N_4815);
and U5458 (N_5458,N_4793,N_4787);
nand U5459 (N_5459,N_4972,N_4658);
and U5460 (N_5460,N_4841,N_4953);
or U5461 (N_5461,N_4791,N_4707);
nor U5462 (N_5462,N_4727,N_4827);
xnor U5463 (N_5463,N_4939,N_4554);
xor U5464 (N_5464,N_4807,N_4722);
nand U5465 (N_5465,N_4686,N_4805);
or U5466 (N_5466,N_4897,N_4856);
or U5467 (N_5467,N_4636,N_4897);
and U5468 (N_5468,N_4921,N_4729);
or U5469 (N_5469,N_4567,N_4558);
or U5470 (N_5470,N_4941,N_4987);
or U5471 (N_5471,N_4525,N_4652);
nand U5472 (N_5472,N_4979,N_4710);
and U5473 (N_5473,N_4509,N_4537);
nand U5474 (N_5474,N_4961,N_4581);
nor U5475 (N_5475,N_4810,N_4744);
xor U5476 (N_5476,N_4864,N_4614);
nand U5477 (N_5477,N_4513,N_4507);
xnor U5478 (N_5478,N_4802,N_4552);
and U5479 (N_5479,N_4558,N_4759);
xnor U5480 (N_5480,N_4923,N_4986);
and U5481 (N_5481,N_4805,N_4520);
and U5482 (N_5482,N_4855,N_4594);
xnor U5483 (N_5483,N_4685,N_4738);
and U5484 (N_5484,N_4894,N_4681);
nand U5485 (N_5485,N_4697,N_4776);
nand U5486 (N_5486,N_4804,N_4869);
nor U5487 (N_5487,N_4667,N_4758);
or U5488 (N_5488,N_4669,N_4525);
nand U5489 (N_5489,N_4900,N_4979);
and U5490 (N_5490,N_4713,N_4874);
and U5491 (N_5491,N_4819,N_4542);
or U5492 (N_5492,N_4950,N_4672);
or U5493 (N_5493,N_4537,N_4670);
or U5494 (N_5494,N_4858,N_4803);
and U5495 (N_5495,N_4631,N_4953);
xor U5496 (N_5496,N_4590,N_4988);
and U5497 (N_5497,N_4622,N_4814);
and U5498 (N_5498,N_4769,N_4544);
xor U5499 (N_5499,N_4672,N_4671);
xnor U5500 (N_5500,N_5307,N_5391);
and U5501 (N_5501,N_5454,N_5445);
nor U5502 (N_5502,N_5011,N_5443);
and U5503 (N_5503,N_5424,N_5235);
nand U5504 (N_5504,N_5249,N_5263);
or U5505 (N_5505,N_5029,N_5300);
and U5506 (N_5506,N_5134,N_5272);
nand U5507 (N_5507,N_5057,N_5299);
nor U5508 (N_5508,N_5356,N_5339);
nor U5509 (N_5509,N_5210,N_5415);
nand U5510 (N_5510,N_5350,N_5075);
and U5511 (N_5511,N_5026,N_5146);
or U5512 (N_5512,N_5083,N_5425);
or U5513 (N_5513,N_5191,N_5273);
nor U5514 (N_5514,N_5481,N_5251);
xnor U5515 (N_5515,N_5274,N_5010);
nand U5516 (N_5516,N_5022,N_5393);
or U5517 (N_5517,N_5015,N_5061);
nor U5518 (N_5518,N_5384,N_5007);
and U5519 (N_5519,N_5448,N_5138);
nand U5520 (N_5520,N_5326,N_5483);
nor U5521 (N_5521,N_5180,N_5330);
nor U5522 (N_5522,N_5184,N_5056);
and U5523 (N_5523,N_5091,N_5468);
or U5524 (N_5524,N_5258,N_5209);
and U5525 (N_5525,N_5136,N_5471);
and U5526 (N_5526,N_5489,N_5141);
nor U5527 (N_5527,N_5065,N_5216);
nand U5528 (N_5528,N_5198,N_5036);
or U5529 (N_5529,N_5004,N_5375);
nand U5530 (N_5530,N_5123,N_5392);
nor U5531 (N_5531,N_5475,N_5217);
and U5532 (N_5532,N_5155,N_5067);
nand U5533 (N_5533,N_5130,N_5094);
and U5534 (N_5534,N_5179,N_5016);
nor U5535 (N_5535,N_5243,N_5494);
nor U5536 (N_5536,N_5014,N_5257);
nand U5537 (N_5537,N_5117,N_5051);
nor U5538 (N_5538,N_5341,N_5319);
nor U5539 (N_5539,N_5360,N_5416);
nand U5540 (N_5540,N_5335,N_5387);
nand U5541 (N_5541,N_5252,N_5241);
xnor U5542 (N_5542,N_5266,N_5012);
or U5543 (N_5543,N_5255,N_5149);
nand U5544 (N_5544,N_5098,N_5054);
or U5545 (N_5545,N_5477,N_5156);
or U5546 (N_5546,N_5143,N_5163);
xnor U5547 (N_5547,N_5039,N_5400);
nand U5548 (N_5548,N_5364,N_5491);
nor U5549 (N_5549,N_5177,N_5275);
and U5550 (N_5550,N_5355,N_5286);
xor U5551 (N_5551,N_5204,N_5404);
or U5552 (N_5552,N_5162,N_5322);
xor U5553 (N_5553,N_5315,N_5159);
and U5554 (N_5554,N_5103,N_5020);
and U5555 (N_5555,N_5389,N_5467);
nor U5556 (N_5556,N_5426,N_5394);
xnor U5557 (N_5557,N_5456,N_5239);
xor U5558 (N_5558,N_5301,N_5213);
and U5559 (N_5559,N_5174,N_5278);
and U5560 (N_5560,N_5265,N_5259);
xnor U5561 (N_5561,N_5462,N_5076);
nand U5562 (N_5562,N_5151,N_5329);
xnor U5563 (N_5563,N_5345,N_5316);
xnor U5564 (N_5564,N_5085,N_5003);
or U5565 (N_5565,N_5225,N_5199);
xor U5566 (N_5566,N_5107,N_5142);
and U5567 (N_5567,N_5070,N_5451);
nand U5568 (N_5568,N_5376,N_5305);
nand U5569 (N_5569,N_5154,N_5227);
nand U5570 (N_5570,N_5441,N_5063);
or U5571 (N_5571,N_5488,N_5205);
nand U5572 (N_5572,N_5127,N_5059);
nor U5573 (N_5573,N_5066,N_5337);
and U5574 (N_5574,N_5385,N_5458);
and U5575 (N_5575,N_5325,N_5452);
nand U5576 (N_5576,N_5013,N_5000);
nand U5577 (N_5577,N_5450,N_5058);
and U5578 (N_5578,N_5062,N_5473);
and U5579 (N_5579,N_5183,N_5147);
xor U5580 (N_5580,N_5101,N_5407);
or U5581 (N_5581,N_5294,N_5303);
nor U5582 (N_5582,N_5422,N_5268);
or U5583 (N_5583,N_5285,N_5292);
nand U5584 (N_5584,N_5283,N_5246);
or U5585 (N_5585,N_5403,N_5112);
nor U5586 (N_5586,N_5476,N_5449);
and U5587 (N_5587,N_5436,N_5496);
nand U5588 (N_5588,N_5055,N_5254);
and U5589 (N_5589,N_5229,N_5412);
or U5590 (N_5590,N_5419,N_5269);
or U5591 (N_5591,N_5228,N_5120);
xor U5592 (N_5592,N_5485,N_5038);
xor U5593 (N_5593,N_5124,N_5069);
xnor U5594 (N_5594,N_5190,N_5108);
nand U5595 (N_5595,N_5318,N_5344);
nand U5596 (N_5596,N_5109,N_5349);
and U5597 (N_5597,N_5406,N_5290);
and U5598 (N_5598,N_5171,N_5167);
nand U5599 (N_5599,N_5173,N_5359);
nand U5600 (N_5600,N_5367,N_5092);
nand U5601 (N_5601,N_5238,N_5245);
xor U5602 (N_5602,N_5479,N_5281);
or U5603 (N_5603,N_5145,N_5081);
nand U5604 (N_5604,N_5095,N_5487);
xor U5605 (N_5605,N_5202,N_5409);
xor U5606 (N_5606,N_5032,N_5370);
nand U5607 (N_5607,N_5442,N_5043);
nor U5608 (N_5608,N_5362,N_5279);
nor U5609 (N_5609,N_5405,N_5484);
and U5610 (N_5610,N_5161,N_5432);
or U5611 (N_5611,N_5386,N_5037);
nor U5612 (N_5612,N_5333,N_5313);
nand U5613 (N_5613,N_5267,N_5495);
nor U5614 (N_5614,N_5165,N_5181);
xor U5615 (N_5615,N_5347,N_5086);
and U5616 (N_5616,N_5122,N_5447);
and U5617 (N_5617,N_5129,N_5474);
and U5618 (N_5618,N_5052,N_5089);
nor U5619 (N_5619,N_5320,N_5044);
nand U5620 (N_5620,N_5050,N_5200);
xnor U5621 (N_5621,N_5352,N_5201);
and U5622 (N_5622,N_5296,N_5433);
or U5623 (N_5623,N_5308,N_5332);
nor U5624 (N_5624,N_5264,N_5446);
or U5625 (N_5625,N_5087,N_5242);
and U5626 (N_5626,N_5035,N_5371);
nand U5627 (N_5627,N_5206,N_5097);
or U5628 (N_5628,N_5119,N_5157);
or U5629 (N_5629,N_5460,N_5293);
or U5630 (N_5630,N_5490,N_5472);
xor U5631 (N_5631,N_5169,N_5423);
nand U5632 (N_5632,N_5455,N_5324);
and U5633 (N_5633,N_5250,N_5223);
and U5634 (N_5634,N_5497,N_5378);
or U5635 (N_5635,N_5176,N_5461);
nand U5636 (N_5636,N_5030,N_5018);
nor U5637 (N_5637,N_5334,N_5288);
xnor U5638 (N_5638,N_5168,N_5253);
nor U5639 (N_5639,N_5492,N_5377);
nand U5640 (N_5640,N_5459,N_5395);
nor U5641 (N_5641,N_5187,N_5219);
xor U5642 (N_5642,N_5233,N_5144);
xor U5643 (N_5643,N_5295,N_5006);
and U5644 (N_5644,N_5312,N_5357);
xnor U5645 (N_5645,N_5017,N_5369);
nand U5646 (N_5646,N_5121,N_5438);
xor U5647 (N_5647,N_5256,N_5033);
xnor U5648 (N_5648,N_5160,N_5499);
xnor U5649 (N_5649,N_5178,N_5222);
xor U5650 (N_5650,N_5262,N_5192);
and U5651 (N_5651,N_5373,N_5457);
xor U5652 (N_5652,N_5388,N_5466);
and U5653 (N_5653,N_5126,N_5413);
nor U5654 (N_5654,N_5166,N_5374);
or U5655 (N_5655,N_5444,N_5398);
nor U5656 (N_5656,N_5019,N_5150);
and U5657 (N_5657,N_5368,N_5282);
nand U5658 (N_5658,N_5310,N_5417);
nand U5659 (N_5659,N_5270,N_5153);
nor U5660 (N_5660,N_5224,N_5226);
xor U5661 (N_5661,N_5137,N_5088);
xor U5662 (N_5662,N_5193,N_5077);
and U5663 (N_5663,N_5351,N_5287);
or U5664 (N_5664,N_5340,N_5480);
nand U5665 (N_5665,N_5203,N_5005);
xor U5666 (N_5666,N_5042,N_5336);
xnor U5667 (N_5667,N_5093,N_5072);
and U5668 (N_5668,N_5429,N_5402);
nor U5669 (N_5669,N_5410,N_5453);
and U5670 (N_5670,N_5148,N_5140);
xor U5671 (N_5671,N_5164,N_5354);
and U5672 (N_5672,N_5431,N_5133);
nand U5673 (N_5673,N_5185,N_5236);
and U5674 (N_5674,N_5358,N_5113);
nor U5675 (N_5675,N_5064,N_5317);
nand U5676 (N_5676,N_5421,N_5197);
nand U5677 (N_5677,N_5323,N_5182);
nor U5678 (N_5678,N_5464,N_5118);
nor U5679 (N_5679,N_5234,N_5220);
or U5680 (N_5680,N_5208,N_5170);
or U5681 (N_5681,N_5414,N_5115);
or U5682 (N_5682,N_5306,N_5309);
xnor U5683 (N_5683,N_5172,N_5175);
and U5684 (N_5684,N_5071,N_5125);
or U5685 (N_5685,N_5248,N_5048);
and U5686 (N_5686,N_5049,N_5260);
xor U5687 (N_5687,N_5399,N_5397);
nor U5688 (N_5688,N_5261,N_5232);
or U5689 (N_5689,N_5338,N_5280);
nand U5690 (N_5690,N_5365,N_5139);
xor U5691 (N_5691,N_5478,N_5396);
and U5692 (N_5692,N_5498,N_5348);
and U5693 (N_5693,N_5240,N_5114);
nor U5694 (N_5694,N_5411,N_5331);
xor U5695 (N_5695,N_5132,N_5372);
and U5696 (N_5696,N_5023,N_5289);
nor U5697 (N_5697,N_5244,N_5096);
nor U5698 (N_5698,N_5040,N_5045);
and U5699 (N_5699,N_5298,N_5382);
xor U5700 (N_5700,N_5218,N_5008);
and U5701 (N_5701,N_5230,N_5434);
nand U5702 (N_5702,N_5221,N_5346);
nand U5703 (N_5703,N_5440,N_5024);
or U5704 (N_5704,N_5408,N_5100);
xnor U5705 (N_5705,N_5090,N_5053);
and U5706 (N_5706,N_5214,N_5231);
or U5707 (N_5707,N_5437,N_5034);
or U5708 (N_5708,N_5366,N_5079);
nor U5709 (N_5709,N_5041,N_5194);
nand U5710 (N_5710,N_5435,N_5401);
xnor U5711 (N_5711,N_5073,N_5002);
or U5712 (N_5712,N_5428,N_5189);
nor U5713 (N_5713,N_5271,N_5084);
or U5714 (N_5714,N_5276,N_5363);
nor U5715 (N_5715,N_5135,N_5128);
nand U5716 (N_5716,N_5379,N_5482);
xnor U5717 (N_5717,N_5284,N_5031);
and U5718 (N_5718,N_5099,N_5342);
nand U5719 (N_5719,N_5297,N_5247);
or U5720 (N_5720,N_5463,N_5418);
xnor U5721 (N_5721,N_5469,N_5211);
and U5722 (N_5722,N_5493,N_5328);
and U5723 (N_5723,N_5237,N_5420);
and U5724 (N_5724,N_5074,N_5047);
and U5725 (N_5725,N_5327,N_5470);
and U5726 (N_5726,N_5188,N_5361);
or U5727 (N_5727,N_5430,N_5082);
and U5728 (N_5728,N_5311,N_5116);
nor U5729 (N_5729,N_5105,N_5046);
nor U5730 (N_5730,N_5080,N_5001);
nor U5731 (N_5731,N_5131,N_5302);
xor U5732 (N_5732,N_5353,N_5186);
nor U5733 (N_5733,N_5277,N_5343);
and U5734 (N_5734,N_5106,N_5021);
nor U5735 (N_5735,N_5028,N_5304);
or U5736 (N_5736,N_5465,N_5060);
nor U5737 (N_5737,N_5439,N_5078);
and U5738 (N_5738,N_5025,N_5207);
nor U5739 (N_5739,N_5195,N_5027);
or U5740 (N_5740,N_5102,N_5427);
nand U5741 (N_5741,N_5111,N_5196);
xor U5742 (N_5742,N_5381,N_5104);
nor U5743 (N_5743,N_5383,N_5152);
nand U5744 (N_5744,N_5212,N_5158);
nand U5745 (N_5745,N_5486,N_5215);
and U5746 (N_5746,N_5068,N_5110);
and U5747 (N_5747,N_5390,N_5009);
and U5748 (N_5748,N_5314,N_5291);
and U5749 (N_5749,N_5321,N_5380);
nor U5750 (N_5750,N_5144,N_5320);
nor U5751 (N_5751,N_5281,N_5422);
and U5752 (N_5752,N_5120,N_5424);
xnor U5753 (N_5753,N_5007,N_5065);
or U5754 (N_5754,N_5184,N_5360);
or U5755 (N_5755,N_5399,N_5485);
nor U5756 (N_5756,N_5006,N_5281);
or U5757 (N_5757,N_5380,N_5095);
nand U5758 (N_5758,N_5313,N_5303);
or U5759 (N_5759,N_5121,N_5186);
and U5760 (N_5760,N_5256,N_5227);
or U5761 (N_5761,N_5018,N_5339);
and U5762 (N_5762,N_5272,N_5114);
nor U5763 (N_5763,N_5421,N_5426);
or U5764 (N_5764,N_5243,N_5324);
nor U5765 (N_5765,N_5280,N_5254);
nand U5766 (N_5766,N_5176,N_5444);
nor U5767 (N_5767,N_5013,N_5269);
nor U5768 (N_5768,N_5259,N_5375);
or U5769 (N_5769,N_5452,N_5393);
nand U5770 (N_5770,N_5161,N_5353);
xor U5771 (N_5771,N_5240,N_5040);
nor U5772 (N_5772,N_5440,N_5463);
and U5773 (N_5773,N_5146,N_5311);
nand U5774 (N_5774,N_5067,N_5410);
nor U5775 (N_5775,N_5182,N_5200);
nand U5776 (N_5776,N_5107,N_5036);
nand U5777 (N_5777,N_5316,N_5079);
nor U5778 (N_5778,N_5258,N_5224);
or U5779 (N_5779,N_5406,N_5184);
or U5780 (N_5780,N_5383,N_5357);
nand U5781 (N_5781,N_5335,N_5295);
and U5782 (N_5782,N_5052,N_5411);
and U5783 (N_5783,N_5167,N_5237);
nor U5784 (N_5784,N_5052,N_5124);
or U5785 (N_5785,N_5041,N_5423);
and U5786 (N_5786,N_5475,N_5107);
or U5787 (N_5787,N_5342,N_5416);
nand U5788 (N_5788,N_5108,N_5235);
nor U5789 (N_5789,N_5009,N_5469);
xor U5790 (N_5790,N_5184,N_5201);
nand U5791 (N_5791,N_5347,N_5191);
xor U5792 (N_5792,N_5490,N_5353);
and U5793 (N_5793,N_5187,N_5070);
nor U5794 (N_5794,N_5359,N_5166);
nand U5795 (N_5795,N_5107,N_5033);
nand U5796 (N_5796,N_5280,N_5261);
xnor U5797 (N_5797,N_5039,N_5474);
and U5798 (N_5798,N_5413,N_5372);
or U5799 (N_5799,N_5070,N_5293);
xor U5800 (N_5800,N_5210,N_5254);
nor U5801 (N_5801,N_5164,N_5338);
nor U5802 (N_5802,N_5194,N_5411);
nor U5803 (N_5803,N_5274,N_5147);
xor U5804 (N_5804,N_5129,N_5405);
xnor U5805 (N_5805,N_5204,N_5276);
nand U5806 (N_5806,N_5260,N_5417);
nand U5807 (N_5807,N_5393,N_5468);
and U5808 (N_5808,N_5057,N_5398);
xor U5809 (N_5809,N_5036,N_5308);
nor U5810 (N_5810,N_5077,N_5365);
nand U5811 (N_5811,N_5022,N_5263);
nand U5812 (N_5812,N_5458,N_5242);
nor U5813 (N_5813,N_5372,N_5095);
or U5814 (N_5814,N_5461,N_5422);
nor U5815 (N_5815,N_5085,N_5186);
and U5816 (N_5816,N_5382,N_5101);
nand U5817 (N_5817,N_5077,N_5470);
nand U5818 (N_5818,N_5374,N_5234);
nor U5819 (N_5819,N_5421,N_5107);
nor U5820 (N_5820,N_5417,N_5148);
nand U5821 (N_5821,N_5186,N_5206);
xor U5822 (N_5822,N_5354,N_5188);
and U5823 (N_5823,N_5195,N_5242);
and U5824 (N_5824,N_5321,N_5383);
nand U5825 (N_5825,N_5244,N_5414);
nor U5826 (N_5826,N_5225,N_5176);
xor U5827 (N_5827,N_5211,N_5398);
nand U5828 (N_5828,N_5492,N_5079);
and U5829 (N_5829,N_5074,N_5293);
and U5830 (N_5830,N_5122,N_5120);
and U5831 (N_5831,N_5334,N_5381);
nor U5832 (N_5832,N_5220,N_5327);
or U5833 (N_5833,N_5140,N_5435);
nor U5834 (N_5834,N_5023,N_5433);
xnor U5835 (N_5835,N_5123,N_5214);
and U5836 (N_5836,N_5362,N_5070);
or U5837 (N_5837,N_5186,N_5132);
or U5838 (N_5838,N_5329,N_5483);
nor U5839 (N_5839,N_5162,N_5200);
nand U5840 (N_5840,N_5077,N_5033);
xor U5841 (N_5841,N_5064,N_5394);
xor U5842 (N_5842,N_5177,N_5394);
nand U5843 (N_5843,N_5380,N_5151);
xnor U5844 (N_5844,N_5303,N_5219);
or U5845 (N_5845,N_5084,N_5472);
nand U5846 (N_5846,N_5060,N_5035);
or U5847 (N_5847,N_5371,N_5309);
and U5848 (N_5848,N_5012,N_5190);
or U5849 (N_5849,N_5425,N_5396);
xor U5850 (N_5850,N_5145,N_5157);
or U5851 (N_5851,N_5264,N_5415);
nand U5852 (N_5852,N_5154,N_5041);
or U5853 (N_5853,N_5424,N_5404);
xor U5854 (N_5854,N_5273,N_5177);
nor U5855 (N_5855,N_5343,N_5475);
xnor U5856 (N_5856,N_5222,N_5342);
and U5857 (N_5857,N_5291,N_5458);
nand U5858 (N_5858,N_5212,N_5370);
or U5859 (N_5859,N_5167,N_5353);
or U5860 (N_5860,N_5130,N_5113);
nand U5861 (N_5861,N_5474,N_5484);
and U5862 (N_5862,N_5488,N_5011);
nand U5863 (N_5863,N_5093,N_5430);
xor U5864 (N_5864,N_5267,N_5247);
nor U5865 (N_5865,N_5122,N_5108);
nand U5866 (N_5866,N_5405,N_5193);
or U5867 (N_5867,N_5216,N_5198);
nor U5868 (N_5868,N_5273,N_5063);
and U5869 (N_5869,N_5340,N_5275);
and U5870 (N_5870,N_5498,N_5294);
nand U5871 (N_5871,N_5389,N_5385);
nor U5872 (N_5872,N_5235,N_5373);
xnor U5873 (N_5873,N_5379,N_5064);
nor U5874 (N_5874,N_5442,N_5245);
nand U5875 (N_5875,N_5394,N_5168);
nor U5876 (N_5876,N_5025,N_5030);
nand U5877 (N_5877,N_5180,N_5216);
or U5878 (N_5878,N_5392,N_5420);
xnor U5879 (N_5879,N_5142,N_5303);
nor U5880 (N_5880,N_5008,N_5248);
and U5881 (N_5881,N_5422,N_5388);
nand U5882 (N_5882,N_5481,N_5003);
and U5883 (N_5883,N_5121,N_5252);
or U5884 (N_5884,N_5385,N_5279);
nand U5885 (N_5885,N_5132,N_5330);
nand U5886 (N_5886,N_5424,N_5076);
xnor U5887 (N_5887,N_5344,N_5124);
or U5888 (N_5888,N_5034,N_5156);
nand U5889 (N_5889,N_5186,N_5081);
nand U5890 (N_5890,N_5163,N_5236);
nor U5891 (N_5891,N_5051,N_5355);
xor U5892 (N_5892,N_5352,N_5462);
and U5893 (N_5893,N_5345,N_5237);
xor U5894 (N_5894,N_5450,N_5106);
nor U5895 (N_5895,N_5494,N_5186);
nor U5896 (N_5896,N_5036,N_5067);
nand U5897 (N_5897,N_5484,N_5124);
and U5898 (N_5898,N_5288,N_5011);
nand U5899 (N_5899,N_5289,N_5428);
nor U5900 (N_5900,N_5405,N_5390);
or U5901 (N_5901,N_5148,N_5220);
and U5902 (N_5902,N_5176,N_5333);
nand U5903 (N_5903,N_5138,N_5204);
xor U5904 (N_5904,N_5113,N_5306);
xnor U5905 (N_5905,N_5338,N_5213);
nand U5906 (N_5906,N_5275,N_5348);
nor U5907 (N_5907,N_5237,N_5416);
and U5908 (N_5908,N_5462,N_5300);
nor U5909 (N_5909,N_5070,N_5279);
and U5910 (N_5910,N_5238,N_5301);
nand U5911 (N_5911,N_5123,N_5106);
and U5912 (N_5912,N_5320,N_5215);
and U5913 (N_5913,N_5180,N_5066);
or U5914 (N_5914,N_5196,N_5239);
nor U5915 (N_5915,N_5378,N_5341);
and U5916 (N_5916,N_5219,N_5186);
xnor U5917 (N_5917,N_5354,N_5237);
and U5918 (N_5918,N_5238,N_5052);
and U5919 (N_5919,N_5256,N_5479);
nor U5920 (N_5920,N_5289,N_5473);
xor U5921 (N_5921,N_5183,N_5188);
xor U5922 (N_5922,N_5279,N_5137);
or U5923 (N_5923,N_5085,N_5349);
and U5924 (N_5924,N_5458,N_5181);
and U5925 (N_5925,N_5051,N_5227);
nor U5926 (N_5926,N_5193,N_5441);
and U5927 (N_5927,N_5496,N_5283);
or U5928 (N_5928,N_5287,N_5058);
xnor U5929 (N_5929,N_5365,N_5402);
nand U5930 (N_5930,N_5455,N_5169);
or U5931 (N_5931,N_5059,N_5454);
nor U5932 (N_5932,N_5010,N_5136);
xnor U5933 (N_5933,N_5415,N_5387);
xnor U5934 (N_5934,N_5283,N_5435);
or U5935 (N_5935,N_5125,N_5210);
and U5936 (N_5936,N_5449,N_5202);
nand U5937 (N_5937,N_5422,N_5487);
xnor U5938 (N_5938,N_5062,N_5217);
xor U5939 (N_5939,N_5114,N_5026);
nor U5940 (N_5940,N_5437,N_5465);
nor U5941 (N_5941,N_5425,N_5162);
nand U5942 (N_5942,N_5253,N_5212);
xor U5943 (N_5943,N_5237,N_5023);
and U5944 (N_5944,N_5253,N_5088);
nor U5945 (N_5945,N_5242,N_5086);
nand U5946 (N_5946,N_5419,N_5232);
and U5947 (N_5947,N_5384,N_5118);
nand U5948 (N_5948,N_5494,N_5420);
and U5949 (N_5949,N_5300,N_5474);
nor U5950 (N_5950,N_5194,N_5060);
or U5951 (N_5951,N_5261,N_5014);
xor U5952 (N_5952,N_5385,N_5074);
nand U5953 (N_5953,N_5118,N_5418);
nand U5954 (N_5954,N_5269,N_5122);
nand U5955 (N_5955,N_5189,N_5498);
nand U5956 (N_5956,N_5456,N_5059);
nor U5957 (N_5957,N_5074,N_5154);
xnor U5958 (N_5958,N_5209,N_5265);
xor U5959 (N_5959,N_5435,N_5082);
xor U5960 (N_5960,N_5117,N_5208);
or U5961 (N_5961,N_5036,N_5236);
nor U5962 (N_5962,N_5303,N_5442);
nand U5963 (N_5963,N_5443,N_5366);
xnor U5964 (N_5964,N_5272,N_5130);
xor U5965 (N_5965,N_5419,N_5422);
xor U5966 (N_5966,N_5467,N_5116);
xnor U5967 (N_5967,N_5271,N_5169);
and U5968 (N_5968,N_5368,N_5425);
xor U5969 (N_5969,N_5450,N_5155);
and U5970 (N_5970,N_5439,N_5236);
xnor U5971 (N_5971,N_5009,N_5199);
nand U5972 (N_5972,N_5178,N_5074);
nor U5973 (N_5973,N_5337,N_5392);
nor U5974 (N_5974,N_5084,N_5450);
and U5975 (N_5975,N_5472,N_5056);
nand U5976 (N_5976,N_5160,N_5123);
xnor U5977 (N_5977,N_5139,N_5395);
nor U5978 (N_5978,N_5417,N_5370);
nand U5979 (N_5979,N_5327,N_5234);
xnor U5980 (N_5980,N_5437,N_5317);
or U5981 (N_5981,N_5055,N_5169);
or U5982 (N_5982,N_5477,N_5303);
and U5983 (N_5983,N_5176,N_5258);
or U5984 (N_5984,N_5133,N_5310);
xor U5985 (N_5985,N_5302,N_5035);
nand U5986 (N_5986,N_5041,N_5336);
xnor U5987 (N_5987,N_5348,N_5189);
xor U5988 (N_5988,N_5103,N_5418);
and U5989 (N_5989,N_5457,N_5417);
and U5990 (N_5990,N_5268,N_5252);
nor U5991 (N_5991,N_5036,N_5070);
xor U5992 (N_5992,N_5188,N_5195);
and U5993 (N_5993,N_5443,N_5209);
nand U5994 (N_5994,N_5296,N_5400);
xnor U5995 (N_5995,N_5311,N_5258);
nor U5996 (N_5996,N_5350,N_5334);
or U5997 (N_5997,N_5240,N_5246);
and U5998 (N_5998,N_5071,N_5388);
xnor U5999 (N_5999,N_5471,N_5055);
nand U6000 (N_6000,N_5521,N_5834);
nor U6001 (N_6001,N_5662,N_5961);
nand U6002 (N_6002,N_5808,N_5588);
xnor U6003 (N_6003,N_5875,N_5667);
nand U6004 (N_6004,N_5764,N_5511);
nor U6005 (N_6005,N_5619,N_5715);
and U6006 (N_6006,N_5753,N_5746);
and U6007 (N_6007,N_5786,N_5925);
and U6008 (N_6008,N_5773,N_5682);
xnor U6009 (N_6009,N_5514,N_5729);
nor U6010 (N_6010,N_5986,N_5696);
nand U6011 (N_6011,N_5972,N_5651);
nor U6012 (N_6012,N_5541,N_5754);
or U6013 (N_6013,N_5862,N_5719);
and U6014 (N_6014,N_5692,N_5607);
nand U6015 (N_6015,N_5706,N_5893);
and U6016 (N_6016,N_5681,N_5683);
xor U6017 (N_6017,N_5830,N_5907);
and U6018 (N_6018,N_5740,N_5699);
or U6019 (N_6019,N_5852,N_5517);
nand U6020 (N_6020,N_5843,N_5707);
or U6021 (N_6021,N_5798,N_5570);
nand U6022 (N_6022,N_5680,N_5591);
nand U6023 (N_6023,N_5794,N_5540);
or U6024 (N_6024,N_5886,N_5596);
nor U6025 (N_6025,N_5948,N_5861);
and U6026 (N_6026,N_5985,N_5880);
or U6027 (N_6027,N_5913,N_5927);
or U6028 (N_6028,N_5530,N_5509);
nor U6029 (N_6029,N_5640,N_5974);
nor U6030 (N_6030,N_5997,N_5564);
nand U6031 (N_6031,N_5603,N_5663);
nor U6032 (N_6032,N_5917,N_5725);
nor U6033 (N_6033,N_5668,N_5868);
and U6034 (N_6034,N_5982,N_5847);
nand U6035 (N_6035,N_5557,N_5935);
and U6036 (N_6036,N_5835,N_5929);
and U6037 (N_6037,N_5920,N_5826);
nor U6038 (N_6038,N_5831,N_5535);
nand U6039 (N_6039,N_5946,N_5547);
xor U6040 (N_6040,N_5989,N_5818);
nand U6041 (N_6041,N_5936,N_5626);
xor U6042 (N_6042,N_5632,N_5611);
or U6043 (N_6043,N_5995,N_5965);
xnor U6044 (N_6044,N_5750,N_5730);
or U6045 (N_6045,N_5556,N_5685);
xor U6046 (N_6046,N_5949,N_5859);
and U6047 (N_6047,N_5615,N_5751);
nand U6048 (N_6048,N_5693,N_5860);
nand U6049 (N_6049,N_5960,N_5910);
and U6050 (N_6050,N_5973,N_5940);
nor U6051 (N_6051,N_5804,N_5643);
nand U6052 (N_6052,N_5784,N_5792);
xnor U6053 (N_6053,N_5785,N_5791);
nor U6054 (N_6054,N_5977,N_5669);
nor U6055 (N_6055,N_5676,N_5656);
and U6056 (N_6056,N_5655,N_5904);
and U6057 (N_6057,N_5871,N_5919);
or U6058 (N_6058,N_5677,N_5811);
nand U6059 (N_6059,N_5762,N_5618);
nor U6060 (N_6060,N_5513,N_5857);
nor U6061 (N_6061,N_5775,N_5614);
and U6062 (N_6062,N_5848,N_5672);
and U6063 (N_6063,N_5781,N_5993);
xor U6064 (N_6064,N_5686,N_5788);
nand U6065 (N_6065,N_5878,N_5900);
nand U6066 (N_6066,N_5732,N_5620);
nor U6067 (N_6067,N_5648,N_5534);
xor U6068 (N_6068,N_5756,N_5539);
and U6069 (N_6069,N_5806,N_5964);
or U6070 (N_6070,N_5994,N_5906);
nand U6071 (N_6071,N_5572,N_5810);
xor U6072 (N_6072,N_5687,N_5864);
xor U6073 (N_6073,N_5518,N_5931);
or U6074 (N_6074,N_5567,N_5969);
nor U6075 (N_6075,N_5749,N_5923);
and U6076 (N_6076,N_5771,N_5722);
or U6077 (N_6077,N_5512,N_5876);
nand U6078 (N_6078,N_5823,N_5665);
nor U6079 (N_6079,N_5580,N_5629);
nand U6080 (N_6080,N_5579,N_5758);
or U6081 (N_6081,N_5795,N_5704);
nor U6082 (N_6082,N_5627,N_5592);
nand U6083 (N_6083,N_5884,N_5744);
or U6084 (N_6084,N_5500,N_5538);
and U6085 (N_6085,N_5713,N_5622);
and U6086 (N_6086,N_5799,N_5597);
and U6087 (N_6087,N_5559,N_5621);
xor U6088 (N_6088,N_5610,N_5658);
or U6089 (N_6089,N_5849,N_5650);
nand U6090 (N_6090,N_5515,N_5708);
and U6091 (N_6091,N_5828,N_5703);
nand U6092 (N_6092,N_5877,N_5737);
nor U6093 (N_6093,N_5934,N_5602);
xor U6094 (N_6094,N_5714,N_5856);
xor U6095 (N_6095,N_5743,N_5953);
or U6096 (N_6096,N_5999,N_5624);
or U6097 (N_6097,N_5780,N_5970);
nor U6098 (N_6098,N_5782,N_5987);
nand U6099 (N_6099,N_5630,N_5723);
or U6100 (N_6100,N_5727,N_5959);
xor U6101 (N_6101,N_5901,N_5678);
nor U6102 (N_6102,N_5976,N_5554);
nor U6103 (N_6103,N_5613,N_5594);
and U6104 (N_6104,N_5947,N_5585);
or U6105 (N_6105,N_5608,N_5590);
nor U6106 (N_6106,N_5657,N_5821);
and U6107 (N_6107,N_5523,N_5674);
xnor U6108 (N_6108,N_5598,N_5646);
or U6109 (N_6109,N_5930,N_5951);
nor U6110 (N_6110,N_5863,N_5774);
and U6111 (N_6111,N_5816,N_5957);
nor U6112 (N_6112,N_5770,N_5736);
nor U6113 (N_6113,N_5752,N_5503);
nand U6114 (N_6114,N_5533,N_5855);
and U6115 (N_6115,N_5832,N_5548);
nor U6116 (N_6116,N_5637,N_5605);
or U6117 (N_6117,N_5793,N_5724);
nand U6118 (N_6118,N_5928,N_5805);
and U6119 (N_6119,N_5894,N_5998);
or U6120 (N_6120,N_5545,N_5887);
nand U6121 (N_6121,N_5892,N_5652);
or U6122 (N_6122,N_5996,N_5659);
xor U6123 (N_6123,N_5566,N_5845);
nor U6124 (N_6124,N_5642,N_5881);
or U6125 (N_6125,N_5552,N_5772);
and U6126 (N_6126,N_5698,N_5765);
xor U6127 (N_6127,N_5889,N_5909);
xor U6128 (N_6128,N_5939,N_5531);
nand U6129 (N_6129,N_5833,N_5790);
and U6130 (N_6130,N_5874,N_5838);
xnor U6131 (N_6131,N_5654,N_5702);
nand U6132 (N_6132,N_5546,N_5731);
and U6133 (N_6133,N_5979,N_5578);
xor U6134 (N_6134,N_5763,N_5912);
xnor U6135 (N_6135,N_5631,N_5918);
nor U6136 (N_6136,N_5922,N_5644);
nor U6137 (N_6137,N_5748,N_5755);
and U6138 (N_6138,N_5924,N_5568);
nor U6139 (N_6139,N_5670,N_5593);
nor U6140 (N_6140,N_5543,N_5779);
xnor U6141 (N_6141,N_5841,N_5710);
nand U6142 (N_6142,N_5777,N_5549);
xnor U6143 (N_6143,N_5522,N_5757);
xor U6144 (N_6144,N_5633,N_5943);
nand U6145 (N_6145,N_5839,N_5589);
and U6146 (N_6146,N_5526,N_5963);
or U6147 (N_6147,N_5885,N_5536);
or U6148 (N_6148,N_5814,N_5563);
and U6149 (N_6149,N_5802,N_5575);
nor U6150 (N_6150,N_5569,N_5600);
nand U6151 (N_6151,N_5898,N_5520);
xor U6152 (N_6152,N_5769,N_5691);
xnor U6153 (N_6153,N_5797,N_5721);
and U6154 (N_6154,N_5609,N_5911);
nand U6155 (N_6155,N_5690,N_5890);
nor U6156 (N_6156,N_5873,N_5689);
xnor U6157 (N_6157,N_5954,N_5776);
or U6158 (N_6158,N_5945,N_5504);
nor U6159 (N_6159,N_5720,N_5870);
nand U6160 (N_6160,N_5617,N_5697);
and U6161 (N_6161,N_5616,N_5813);
nor U6162 (N_6162,N_5941,N_5837);
nand U6163 (N_6163,N_5915,N_5623);
xor U6164 (N_6164,N_5789,N_5846);
nor U6165 (N_6165,N_5711,N_5747);
or U6166 (N_6166,N_5738,N_5636);
xor U6167 (N_6167,N_5506,N_5502);
nand U6168 (N_6168,N_5801,N_5952);
nand U6169 (N_6169,N_5967,N_5525);
nor U6170 (N_6170,N_5807,N_5741);
xnor U6171 (N_6171,N_5942,N_5641);
nand U6172 (N_6172,N_5815,N_5825);
and U6173 (N_6173,N_5718,N_5679);
nand U6174 (N_6174,N_5990,N_5955);
and U6175 (N_6175,N_5767,N_5992);
and U6176 (N_6176,N_5537,N_5867);
nand U6177 (N_6177,N_5712,N_5604);
or U6178 (N_6178,N_5958,N_5684);
and U6179 (N_6179,N_5968,N_5778);
and U6180 (N_6180,N_5980,N_5984);
nor U6181 (N_6181,N_5817,N_5734);
nor U6182 (N_6182,N_5975,N_5950);
and U6183 (N_6183,N_5660,N_5649);
and U6184 (N_6184,N_5638,N_5803);
nor U6185 (N_6185,N_5854,N_5571);
and U6186 (N_6186,N_5819,N_5879);
and U6187 (N_6187,N_5991,N_5516);
nand U6188 (N_6188,N_5664,N_5824);
nor U6189 (N_6189,N_5760,N_5944);
nand U6190 (N_6190,N_5921,N_5587);
nor U6191 (N_6191,N_5739,N_5584);
and U6192 (N_6192,N_5606,N_5836);
or U6193 (N_6193,N_5796,N_5905);
nor U6194 (N_6194,N_5524,N_5695);
nor U6195 (N_6195,N_5544,N_5601);
nor U6196 (N_6196,N_5895,N_5519);
or U6197 (N_6197,N_5717,N_5899);
or U6198 (N_6198,N_5812,N_5716);
or U6199 (N_6199,N_5705,N_5896);
and U6200 (N_6200,N_5562,N_5822);
xor U6201 (N_6201,N_5565,N_5745);
nand U6202 (N_6202,N_5661,N_5787);
nor U6203 (N_6203,N_5865,N_5573);
nor U6204 (N_6204,N_5561,N_5625);
nor U6205 (N_6205,N_5555,N_5783);
nor U6206 (N_6206,N_5527,N_5529);
or U6207 (N_6207,N_5914,N_5532);
and U6208 (N_6208,N_5688,N_5891);
xor U6209 (N_6209,N_5932,N_5827);
and U6210 (N_6210,N_5842,N_5595);
nand U6211 (N_6211,N_5908,N_5505);
xnor U6212 (N_6212,N_5673,N_5766);
xnor U6213 (N_6213,N_5851,N_5528);
nand U6214 (N_6214,N_5872,N_5666);
and U6215 (N_6215,N_5768,N_5574);
nand U6216 (N_6216,N_5553,N_5709);
and U6217 (N_6217,N_5510,N_5694);
nor U6218 (N_6218,N_5844,N_5675);
nand U6219 (N_6219,N_5586,N_5820);
nor U6220 (N_6220,N_5866,N_5560);
nor U6221 (N_6221,N_5853,N_5903);
nand U6222 (N_6222,N_5628,N_5761);
xor U6223 (N_6223,N_5869,N_5971);
or U6224 (N_6224,N_5926,N_5700);
nand U6225 (N_6225,N_5726,N_5988);
and U6226 (N_6226,N_5581,N_5882);
or U6227 (N_6227,N_5653,N_5829);
or U6228 (N_6228,N_5883,N_5542);
nand U6229 (N_6229,N_5759,N_5634);
xor U6230 (N_6230,N_5551,N_5508);
and U6231 (N_6231,N_5647,N_5981);
and U6232 (N_6232,N_5962,N_5966);
or U6233 (N_6233,N_5933,N_5916);
xor U6234 (N_6234,N_5635,N_5558);
nand U6235 (N_6235,N_5850,N_5612);
nand U6236 (N_6236,N_5583,N_5809);
or U6237 (N_6237,N_5897,N_5800);
nand U6238 (N_6238,N_5888,N_5902);
nor U6239 (N_6239,N_5501,N_5937);
nor U6240 (N_6240,N_5576,N_5728);
xnor U6241 (N_6241,N_5978,N_5735);
and U6242 (N_6242,N_5938,N_5550);
or U6243 (N_6243,N_5507,N_5956);
and U6244 (N_6244,N_5858,N_5645);
nand U6245 (N_6245,N_5840,N_5701);
and U6246 (N_6246,N_5582,N_5983);
nor U6247 (N_6247,N_5639,N_5599);
nor U6248 (N_6248,N_5577,N_5671);
nor U6249 (N_6249,N_5733,N_5742);
or U6250 (N_6250,N_5721,N_5695);
nand U6251 (N_6251,N_5984,N_5601);
nor U6252 (N_6252,N_5956,N_5541);
nand U6253 (N_6253,N_5520,N_5676);
nor U6254 (N_6254,N_5812,N_5701);
or U6255 (N_6255,N_5724,N_5559);
or U6256 (N_6256,N_5846,N_5562);
nand U6257 (N_6257,N_5819,N_5731);
or U6258 (N_6258,N_5953,N_5501);
and U6259 (N_6259,N_5774,N_5717);
xor U6260 (N_6260,N_5871,N_5679);
nand U6261 (N_6261,N_5980,N_5900);
nor U6262 (N_6262,N_5558,N_5717);
xor U6263 (N_6263,N_5523,N_5582);
nand U6264 (N_6264,N_5856,N_5592);
xor U6265 (N_6265,N_5504,N_5871);
nand U6266 (N_6266,N_5827,N_5833);
nand U6267 (N_6267,N_5958,N_5874);
nand U6268 (N_6268,N_5665,N_5888);
xor U6269 (N_6269,N_5737,N_5727);
nand U6270 (N_6270,N_5745,N_5569);
nor U6271 (N_6271,N_5571,N_5763);
nor U6272 (N_6272,N_5975,N_5801);
nor U6273 (N_6273,N_5517,N_5962);
or U6274 (N_6274,N_5702,N_5557);
or U6275 (N_6275,N_5785,N_5959);
nand U6276 (N_6276,N_5753,N_5854);
or U6277 (N_6277,N_5514,N_5896);
nand U6278 (N_6278,N_5899,N_5647);
nor U6279 (N_6279,N_5782,N_5678);
xnor U6280 (N_6280,N_5594,N_5813);
xnor U6281 (N_6281,N_5602,N_5838);
and U6282 (N_6282,N_5930,N_5728);
and U6283 (N_6283,N_5766,N_5633);
xor U6284 (N_6284,N_5537,N_5752);
nor U6285 (N_6285,N_5902,N_5727);
or U6286 (N_6286,N_5980,N_5642);
nor U6287 (N_6287,N_5699,N_5559);
nand U6288 (N_6288,N_5792,N_5913);
nand U6289 (N_6289,N_5699,N_5653);
or U6290 (N_6290,N_5703,N_5761);
nor U6291 (N_6291,N_5562,N_5727);
and U6292 (N_6292,N_5548,N_5918);
or U6293 (N_6293,N_5506,N_5869);
nand U6294 (N_6294,N_5756,N_5628);
nor U6295 (N_6295,N_5929,N_5836);
or U6296 (N_6296,N_5657,N_5723);
nand U6297 (N_6297,N_5596,N_5892);
or U6298 (N_6298,N_5689,N_5626);
nor U6299 (N_6299,N_5836,N_5961);
nor U6300 (N_6300,N_5863,N_5525);
or U6301 (N_6301,N_5703,N_5635);
nor U6302 (N_6302,N_5844,N_5721);
nand U6303 (N_6303,N_5576,N_5908);
and U6304 (N_6304,N_5892,N_5853);
nand U6305 (N_6305,N_5884,N_5818);
nor U6306 (N_6306,N_5980,N_5825);
or U6307 (N_6307,N_5518,N_5858);
nor U6308 (N_6308,N_5782,N_5900);
or U6309 (N_6309,N_5661,N_5986);
nand U6310 (N_6310,N_5841,N_5526);
and U6311 (N_6311,N_5984,N_5832);
nor U6312 (N_6312,N_5784,N_5851);
nand U6313 (N_6313,N_5518,N_5814);
nor U6314 (N_6314,N_5984,N_5986);
xor U6315 (N_6315,N_5891,N_5563);
or U6316 (N_6316,N_5681,N_5858);
xnor U6317 (N_6317,N_5985,N_5821);
or U6318 (N_6318,N_5961,N_5978);
nand U6319 (N_6319,N_5763,N_5536);
xnor U6320 (N_6320,N_5623,N_5849);
xnor U6321 (N_6321,N_5792,N_5985);
nand U6322 (N_6322,N_5632,N_5662);
or U6323 (N_6323,N_5736,N_5943);
nor U6324 (N_6324,N_5851,N_5618);
nor U6325 (N_6325,N_5579,N_5808);
and U6326 (N_6326,N_5813,N_5967);
nand U6327 (N_6327,N_5782,N_5700);
nand U6328 (N_6328,N_5681,N_5560);
or U6329 (N_6329,N_5752,N_5663);
nor U6330 (N_6330,N_5986,N_5819);
and U6331 (N_6331,N_5604,N_5801);
and U6332 (N_6332,N_5875,N_5895);
or U6333 (N_6333,N_5755,N_5759);
xnor U6334 (N_6334,N_5778,N_5613);
or U6335 (N_6335,N_5739,N_5803);
or U6336 (N_6336,N_5850,N_5770);
nor U6337 (N_6337,N_5568,N_5739);
and U6338 (N_6338,N_5593,N_5858);
or U6339 (N_6339,N_5724,N_5954);
nand U6340 (N_6340,N_5727,N_5893);
nand U6341 (N_6341,N_5799,N_5986);
nand U6342 (N_6342,N_5783,N_5989);
and U6343 (N_6343,N_5581,N_5752);
nor U6344 (N_6344,N_5849,N_5744);
and U6345 (N_6345,N_5693,N_5781);
or U6346 (N_6346,N_5659,N_5530);
and U6347 (N_6347,N_5866,N_5510);
or U6348 (N_6348,N_5778,N_5690);
xnor U6349 (N_6349,N_5897,N_5778);
or U6350 (N_6350,N_5990,N_5515);
and U6351 (N_6351,N_5666,N_5564);
nand U6352 (N_6352,N_5770,N_5768);
xnor U6353 (N_6353,N_5935,N_5848);
or U6354 (N_6354,N_5916,N_5893);
nand U6355 (N_6355,N_5581,N_5739);
or U6356 (N_6356,N_5941,N_5598);
nor U6357 (N_6357,N_5794,N_5801);
nand U6358 (N_6358,N_5553,N_5875);
nand U6359 (N_6359,N_5838,N_5614);
and U6360 (N_6360,N_5789,N_5689);
and U6361 (N_6361,N_5749,N_5598);
xnor U6362 (N_6362,N_5666,N_5594);
and U6363 (N_6363,N_5860,N_5949);
nor U6364 (N_6364,N_5935,N_5518);
nand U6365 (N_6365,N_5793,N_5565);
nand U6366 (N_6366,N_5813,N_5953);
nor U6367 (N_6367,N_5539,N_5585);
or U6368 (N_6368,N_5536,N_5615);
xor U6369 (N_6369,N_5606,N_5852);
nor U6370 (N_6370,N_5753,N_5668);
nor U6371 (N_6371,N_5646,N_5511);
and U6372 (N_6372,N_5738,N_5708);
and U6373 (N_6373,N_5529,N_5940);
and U6374 (N_6374,N_5707,N_5569);
nor U6375 (N_6375,N_5624,N_5637);
or U6376 (N_6376,N_5983,N_5973);
nor U6377 (N_6377,N_5724,N_5524);
nor U6378 (N_6378,N_5535,N_5969);
and U6379 (N_6379,N_5873,N_5634);
xnor U6380 (N_6380,N_5719,N_5794);
and U6381 (N_6381,N_5878,N_5999);
or U6382 (N_6382,N_5810,N_5897);
and U6383 (N_6383,N_5885,N_5707);
nor U6384 (N_6384,N_5679,N_5613);
and U6385 (N_6385,N_5774,N_5809);
nor U6386 (N_6386,N_5729,N_5996);
nand U6387 (N_6387,N_5610,N_5985);
and U6388 (N_6388,N_5765,N_5952);
or U6389 (N_6389,N_5836,N_5870);
and U6390 (N_6390,N_5658,N_5685);
or U6391 (N_6391,N_5899,N_5956);
xor U6392 (N_6392,N_5575,N_5543);
xnor U6393 (N_6393,N_5890,N_5704);
and U6394 (N_6394,N_5835,N_5814);
xnor U6395 (N_6395,N_5653,N_5787);
xnor U6396 (N_6396,N_5680,N_5748);
nand U6397 (N_6397,N_5626,N_5655);
nor U6398 (N_6398,N_5812,N_5624);
nand U6399 (N_6399,N_5910,N_5629);
nand U6400 (N_6400,N_5861,N_5869);
xnor U6401 (N_6401,N_5774,N_5951);
xor U6402 (N_6402,N_5704,N_5901);
and U6403 (N_6403,N_5673,N_5681);
and U6404 (N_6404,N_5603,N_5521);
xnor U6405 (N_6405,N_5837,N_5798);
and U6406 (N_6406,N_5631,N_5629);
xnor U6407 (N_6407,N_5808,N_5506);
or U6408 (N_6408,N_5835,N_5648);
xor U6409 (N_6409,N_5740,N_5775);
xnor U6410 (N_6410,N_5704,N_5973);
nor U6411 (N_6411,N_5935,N_5770);
nor U6412 (N_6412,N_5647,N_5934);
or U6413 (N_6413,N_5595,N_5943);
nand U6414 (N_6414,N_5899,N_5846);
nand U6415 (N_6415,N_5668,N_5835);
xor U6416 (N_6416,N_5598,N_5570);
and U6417 (N_6417,N_5893,N_5918);
and U6418 (N_6418,N_5934,N_5859);
or U6419 (N_6419,N_5684,N_5740);
and U6420 (N_6420,N_5542,N_5834);
and U6421 (N_6421,N_5635,N_5793);
and U6422 (N_6422,N_5896,N_5629);
or U6423 (N_6423,N_5891,N_5972);
and U6424 (N_6424,N_5877,N_5887);
nor U6425 (N_6425,N_5822,N_5813);
and U6426 (N_6426,N_5710,N_5942);
or U6427 (N_6427,N_5811,N_5585);
and U6428 (N_6428,N_5759,N_5606);
nor U6429 (N_6429,N_5814,N_5903);
and U6430 (N_6430,N_5910,N_5683);
xnor U6431 (N_6431,N_5500,N_5684);
and U6432 (N_6432,N_5667,N_5691);
or U6433 (N_6433,N_5825,N_5552);
or U6434 (N_6434,N_5764,N_5842);
nor U6435 (N_6435,N_5577,N_5711);
or U6436 (N_6436,N_5533,N_5964);
and U6437 (N_6437,N_5650,N_5740);
nand U6438 (N_6438,N_5811,N_5839);
xor U6439 (N_6439,N_5664,N_5846);
nor U6440 (N_6440,N_5788,N_5854);
xnor U6441 (N_6441,N_5692,N_5870);
or U6442 (N_6442,N_5858,N_5784);
nand U6443 (N_6443,N_5641,N_5574);
xnor U6444 (N_6444,N_5915,N_5996);
nand U6445 (N_6445,N_5840,N_5581);
nor U6446 (N_6446,N_5705,N_5524);
or U6447 (N_6447,N_5813,N_5532);
or U6448 (N_6448,N_5935,N_5853);
nor U6449 (N_6449,N_5708,N_5887);
and U6450 (N_6450,N_5596,N_5550);
nand U6451 (N_6451,N_5588,N_5750);
nand U6452 (N_6452,N_5571,N_5695);
xor U6453 (N_6453,N_5763,N_5645);
nor U6454 (N_6454,N_5970,N_5526);
or U6455 (N_6455,N_5867,N_5954);
nor U6456 (N_6456,N_5828,N_5589);
xor U6457 (N_6457,N_5785,N_5932);
nor U6458 (N_6458,N_5727,N_5946);
or U6459 (N_6459,N_5994,N_5511);
xor U6460 (N_6460,N_5604,N_5739);
xnor U6461 (N_6461,N_5631,N_5821);
xnor U6462 (N_6462,N_5886,N_5612);
and U6463 (N_6463,N_5752,N_5723);
or U6464 (N_6464,N_5996,N_5753);
or U6465 (N_6465,N_5607,N_5579);
and U6466 (N_6466,N_5571,N_5504);
xor U6467 (N_6467,N_5868,N_5917);
nor U6468 (N_6468,N_5960,N_5571);
xor U6469 (N_6469,N_5813,N_5516);
nor U6470 (N_6470,N_5810,N_5648);
xnor U6471 (N_6471,N_5952,N_5915);
nand U6472 (N_6472,N_5561,N_5591);
and U6473 (N_6473,N_5764,N_5520);
xor U6474 (N_6474,N_5749,N_5990);
and U6475 (N_6475,N_5520,N_5652);
nand U6476 (N_6476,N_5732,N_5644);
nor U6477 (N_6477,N_5667,N_5989);
xor U6478 (N_6478,N_5990,N_5555);
xor U6479 (N_6479,N_5858,N_5788);
nor U6480 (N_6480,N_5543,N_5770);
and U6481 (N_6481,N_5550,N_5743);
xor U6482 (N_6482,N_5848,N_5763);
or U6483 (N_6483,N_5815,N_5967);
xor U6484 (N_6484,N_5648,N_5783);
xor U6485 (N_6485,N_5857,N_5554);
and U6486 (N_6486,N_5968,N_5676);
xor U6487 (N_6487,N_5967,N_5796);
xnor U6488 (N_6488,N_5719,N_5731);
nor U6489 (N_6489,N_5597,N_5523);
nor U6490 (N_6490,N_5550,N_5539);
xor U6491 (N_6491,N_5755,N_5627);
xnor U6492 (N_6492,N_5702,N_5959);
or U6493 (N_6493,N_5792,N_5631);
or U6494 (N_6494,N_5803,N_5833);
and U6495 (N_6495,N_5891,N_5633);
or U6496 (N_6496,N_5914,N_5944);
or U6497 (N_6497,N_5828,N_5872);
nand U6498 (N_6498,N_5739,N_5623);
nor U6499 (N_6499,N_5686,N_5995);
nor U6500 (N_6500,N_6358,N_6190);
or U6501 (N_6501,N_6443,N_6131);
xor U6502 (N_6502,N_6000,N_6044);
nand U6503 (N_6503,N_6430,N_6300);
or U6504 (N_6504,N_6294,N_6041);
xnor U6505 (N_6505,N_6462,N_6260);
or U6506 (N_6506,N_6224,N_6450);
xnor U6507 (N_6507,N_6246,N_6075);
nand U6508 (N_6508,N_6205,N_6267);
xor U6509 (N_6509,N_6315,N_6382);
or U6510 (N_6510,N_6001,N_6432);
or U6511 (N_6511,N_6411,N_6169);
nor U6512 (N_6512,N_6365,N_6182);
nand U6513 (N_6513,N_6008,N_6475);
nand U6514 (N_6514,N_6407,N_6334);
nand U6515 (N_6515,N_6363,N_6264);
and U6516 (N_6516,N_6184,N_6291);
nor U6517 (N_6517,N_6012,N_6188);
xor U6518 (N_6518,N_6123,N_6158);
nand U6519 (N_6519,N_6074,N_6192);
nand U6520 (N_6520,N_6311,N_6157);
nor U6521 (N_6521,N_6455,N_6293);
and U6522 (N_6522,N_6354,N_6189);
and U6523 (N_6523,N_6346,N_6035);
nor U6524 (N_6524,N_6233,N_6400);
nor U6525 (N_6525,N_6499,N_6017);
or U6526 (N_6526,N_6173,N_6488);
or U6527 (N_6527,N_6042,N_6060);
and U6528 (N_6528,N_6222,N_6471);
nand U6529 (N_6529,N_6329,N_6433);
xnor U6530 (N_6530,N_6243,N_6106);
xor U6531 (N_6531,N_6024,N_6410);
xnor U6532 (N_6532,N_6419,N_6467);
xnor U6533 (N_6533,N_6491,N_6439);
nand U6534 (N_6534,N_6061,N_6402);
or U6535 (N_6535,N_6238,N_6466);
xnor U6536 (N_6536,N_6193,N_6463);
xor U6537 (N_6537,N_6219,N_6468);
and U6538 (N_6538,N_6047,N_6235);
nand U6539 (N_6539,N_6226,N_6498);
xor U6540 (N_6540,N_6054,N_6062);
xor U6541 (N_6541,N_6453,N_6357);
nand U6542 (N_6542,N_6483,N_6280);
nor U6543 (N_6543,N_6025,N_6415);
nand U6544 (N_6544,N_6253,N_6112);
and U6545 (N_6545,N_6201,N_6016);
xnor U6546 (N_6546,N_6218,N_6163);
xnor U6547 (N_6547,N_6091,N_6442);
nand U6548 (N_6548,N_6341,N_6274);
xnor U6549 (N_6549,N_6141,N_6362);
and U6550 (N_6550,N_6405,N_6456);
or U6551 (N_6551,N_6109,N_6277);
nand U6552 (N_6552,N_6327,N_6162);
nor U6553 (N_6553,N_6428,N_6107);
nand U6554 (N_6554,N_6139,N_6104);
nand U6555 (N_6555,N_6322,N_6198);
nand U6556 (N_6556,N_6252,N_6132);
and U6557 (N_6557,N_6090,N_6420);
nor U6558 (N_6558,N_6036,N_6495);
nand U6559 (N_6559,N_6383,N_6261);
and U6560 (N_6560,N_6019,N_6371);
xnor U6561 (N_6561,N_6368,N_6221);
or U6562 (N_6562,N_6323,N_6231);
and U6563 (N_6563,N_6404,N_6406);
nor U6564 (N_6564,N_6375,N_6048);
nor U6565 (N_6565,N_6345,N_6077);
nor U6566 (N_6566,N_6178,N_6101);
and U6567 (N_6567,N_6318,N_6305);
and U6568 (N_6568,N_6389,N_6349);
nand U6569 (N_6569,N_6333,N_6129);
nor U6570 (N_6570,N_6076,N_6203);
or U6571 (N_6571,N_6046,N_6356);
xor U6572 (N_6572,N_6195,N_6223);
nand U6573 (N_6573,N_6236,N_6102);
nand U6574 (N_6574,N_6103,N_6339);
and U6575 (N_6575,N_6239,N_6241);
and U6576 (N_6576,N_6031,N_6342);
nand U6577 (N_6577,N_6004,N_6066);
and U6578 (N_6578,N_6210,N_6181);
xnor U6579 (N_6579,N_6388,N_6056);
and U6580 (N_6580,N_6474,N_6172);
xor U6581 (N_6581,N_6020,N_6321);
nor U6582 (N_6582,N_6299,N_6118);
and U6583 (N_6583,N_6023,N_6229);
or U6584 (N_6584,N_6209,N_6298);
xnor U6585 (N_6585,N_6331,N_6426);
and U6586 (N_6586,N_6207,N_6372);
or U6587 (N_6587,N_6282,N_6204);
xor U6588 (N_6588,N_6175,N_6458);
xnor U6589 (N_6589,N_6228,N_6137);
xor U6590 (N_6590,N_6465,N_6401);
xnor U6591 (N_6591,N_6324,N_6065);
or U6592 (N_6592,N_6496,N_6427);
and U6593 (N_6593,N_6134,N_6251);
or U6594 (N_6594,N_6257,N_6119);
xor U6595 (N_6595,N_6418,N_6220);
and U6596 (N_6596,N_6494,N_6069);
nand U6597 (N_6597,N_6304,N_6288);
and U6598 (N_6598,N_6308,N_6146);
xor U6599 (N_6599,N_6459,N_6088);
and U6600 (N_6600,N_6399,N_6217);
or U6601 (N_6601,N_6492,N_6227);
nand U6602 (N_6602,N_6307,N_6050);
or U6603 (N_6603,N_6270,N_6097);
nor U6604 (N_6604,N_6285,N_6234);
and U6605 (N_6605,N_6170,N_6258);
and U6606 (N_6606,N_6249,N_6472);
or U6607 (N_6607,N_6350,N_6026);
nor U6608 (N_6608,N_6166,N_6271);
or U6609 (N_6609,N_6040,N_6437);
and U6610 (N_6610,N_6049,N_6167);
nor U6611 (N_6611,N_6160,N_6216);
or U6612 (N_6612,N_6150,N_6142);
or U6613 (N_6613,N_6164,N_6151);
xor U6614 (N_6614,N_6336,N_6072);
or U6615 (N_6615,N_6087,N_6063);
nor U6616 (N_6616,N_6117,N_6148);
nand U6617 (N_6617,N_6337,N_6099);
or U6618 (N_6618,N_6423,N_6068);
or U6619 (N_6619,N_6259,N_6010);
or U6620 (N_6620,N_6018,N_6032);
nand U6621 (N_6621,N_6125,N_6133);
nor U6622 (N_6622,N_6449,N_6470);
nor U6623 (N_6623,N_6376,N_6457);
nand U6624 (N_6624,N_6309,N_6037);
xnor U6625 (N_6625,N_6461,N_6344);
nand U6626 (N_6626,N_6168,N_6355);
and U6627 (N_6627,N_6155,N_6444);
xnor U6628 (N_6628,N_6295,N_6185);
and U6629 (N_6629,N_6263,N_6250);
nor U6630 (N_6630,N_6211,N_6165);
xor U6631 (N_6631,N_6409,N_6071);
nand U6632 (N_6632,N_6335,N_6454);
or U6633 (N_6633,N_6265,N_6292);
or U6634 (N_6634,N_6338,N_6394);
nand U6635 (N_6635,N_6197,N_6115);
nor U6636 (N_6636,N_6413,N_6002);
and U6637 (N_6637,N_6176,N_6180);
xor U6638 (N_6638,N_6098,N_6484);
or U6639 (N_6639,N_6244,N_6384);
xnor U6640 (N_6640,N_6473,N_6398);
nor U6641 (N_6641,N_6124,N_6378);
nand U6642 (N_6642,N_6199,N_6385);
xor U6643 (N_6643,N_6396,N_6092);
nand U6644 (N_6644,N_6445,N_6177);
nand U6645 (N_6645,N_6248,N_6128);
or U6646 (N_6646,N_6397,N_6353);
or U6647 (N_6647,N_6007,N_6225);
nor U6648 (N_6648,N_6441,N_6127);
and U6649 (N_6649,N_6014,N_6395);
or U6650 (N_6650,N_6206,N_6369);
nand U6651 (N_6651,N_6370,N_6108);
nand U6652 (N_6652,N_6464,N_6469);
nand U6653 (N_6653,N_6183,N_6306);
nand U6654 (N_6654,N_6200,N_6380);
or U6655 (N_6655,N_6301,N_6414);
or U6656 (N_6656,N_6312,N_6144);
nor U6657 (N_6657,N_6240,N_6290);
nor U6658 (N_6658,N_6424,N_6269);
and U6659 (N_6659,N_6482,N_6254);
nand U6660 (N_6660,N_6029,N_6256);
or U6661 (N_6661,N_6296,N_6094);
or U6662 (N_6662,N_6143,N_6320);
nand U6663 (N_6663,N_6045,N_6078);
xnor U6664 (N_6664,N_6493,N_6212);
xor U6665 (N_6665,N_6003,N_6171);
xnor U6666 (N_6666,N_6314,N_6232);
xnor U6667 (N_6667,N_6057,N_6360);
xnor U6668 (N_6668,N_6276,N_6051);
nor U6669 (N_6669,N_6245,N_6079);
or U6670 (N_6670,N_6489,N_6110);
nand U6671 (N_6671,N_6479,N_6093);
nor U6672 (N_6672,N_6043,N_6325);
xor U6673 (N_6673,N_6120,N_6438);
and U6674 (N_6674,N_6135,N_6281);
or U6675 (N_6675,N_6343,N_6303);
xnor U6676 (N_6676,N_6302,N_6242);
and U6677 (N_6677,N_6081,N_6147);
and U6678 (N_6678,N_6352,N_6435);
xor U6679 (N_6679,N_6310,N_6237);
nor U6680 (N_6680,N_6408,N_6392);
or U6681 (N_6681,N_6287,N_6340);
xor U6682 (N_6682,N_6390,N_6191);
or U6683 (N_6683,N_6215,N_6196);
nor U6684 (N_6684,N_6089,N_6015);
nand U6685 (N_6685,N_6359,N_6422);
xor U6686 (N_6686,N_6161,N_6366);
and U6687 (N_6687,N_6431,N_6214);
or U6688 (N_6688,N_6393,N_6297);
nand U6689 (N_6689,N_6027,N_6053);
xor U6690 (N_6690,N_6417,N_6033);
or U6691 (N_6691,N_6332,N_6403);
nor U6692 (N_6692,N_6064,N_6154);
nor U6693 (N_6693,N_6011,N_6425);
or U6694 (N_6694,N_6364,N_6497);
xnor U6695 (N_6695,N_6286,N_6289);
xnor U6696 (N_6696,N_6095,N_6159);
and U6697 (N_6697,N_6429,N_6179);
xor U6698 (N_6698,N_6412,N_6052);
nor U6699 (N_6699,N_6138,N_6085);
nand U6700 (N_6700,N_6202,N_6194);
xnor U6701 (N_6701,N_6275,N_6476);
and U6702 (N_6702,N_6446,N_6013);
or U6703 (N_6703,N_6230,N_6436);
xnor U6704 (N_6704,N_6096,N_6114);
nand U6705 (N_6705,N_6028,N_6039);
nor U6706 (N_6706,N_6121,N_6313);
nor U6707 (N_6707,N_6113,N_6174);
and U6708 (N_6708,N_6122,N_6373);
or U6709 (N_6709,N_6481,N_6213);
xor U6710 (N_6710,N_6480,N_6105);
and U6711 (N_6711,N_6416,N_6319);
xnor U6712 (N_6712,N_6367,N_6006);
xor U6713 (N_6713,N_6059,N_6247);
nor U6714 (N_6714,N_6374,N_6130);
or U6715 (N_6715,N_6283,N_6272);
or U6716 (N_6716,N_6421,N_6030);
nand U6717 (N_6717,N_6284,N_6434);
xor U6718 (N_6718,N_6485,N_6326);
or U6719 (N_6719,N_6022,N_6361);
xnor U6720 (N_6720,N_6034,N_6086);
or U6721 (N_6721,N_6268,N_6153);
nand U6722 (N_6722,N_6316,N_6391);
or U6723 (N_6723,N_6070,N_6278);
nand U6724 (N_6724,N_6381,N_6084);
nor U6725 (N_6725,N_6116,N_6058);
nor U6726 (N_6726,N_6186,N_6149);
xnor U6727 (N_6727,N_6486,N_6387);
nor U6728 (N_6728,N_6208,N_6080);
or U6729 (N_6729,N_6273,N_6126);
nand U6730 (N_6730,N_6082,N_6005);
or U6731 (N_6731,N_6347,N_6083);
nor U6732 (N_6732,N_6152,N_6490);
nor U6733 (N_6733,N_6448,N_6145);
xor U6734 (N_6734,N_6451,N_6351);
xor U6735 (N_6735,N_6330,N_6452);
and U6736 (N_6736,N_6317,N_6262);
nor U6737 (N_6737,N_6156,N_6478);
nor U6738 (N_6738,N_6279,N_6440);
nand U6739 (N_6739,N_6266,N_6255);
nand U6740 (N_6740,N_6055,N_6460);
or U6741 (N_6741,N_6038,N_6348);
xnor U6742 (N_6742,N_6100,N_6009);
xnor U6743 (N_6743,N_6021,N_6136);
nor U6744 (N_6744,N_6377,N_6067);
and U6745 (N_6745,N_6187,N_6111);
xor U6746 (N_6746,N_6487,N_6477);
nand U6747 (N_6747,N_6140,N_6379);
xnor U6748 (N_6748,N_6073,N_6328);
and U6749 (N_6749,N_6386,N_6447);
xnor U6750 (N_6750,N_6076,N_6411);
or U6751 (N_6751,N_6015,N_6126);
or U6752 (N_6752,N_6499,N_6420);
nor U6753 (N_6753,N_6375,N_6024);
or U6754 (N_6754,N_6163,N_6170);
and U6755 (N_6755,N_6461,N_6207);
xnor U6756 (N_6756,N_6054,N_6143);
nor U6757 (N_6757,N_6220,N_6182);
or U6758 (N_6758,N_6235,N_6076);
xnor U6759 (N_6759,N_6287,N_6187);
nand U6760 (N_6760,N_6063,N_6196);
nor U6761 (N_6761,N_6176,N_6478);
nor U6762 (N_6762,N_6189,N_6100);
or U6763 (N_6763,N_6108,N_6086);
nand U6764 (N_6764,N_6476,N_6292);
nor U6765 (N_6765,N_6267,N_6156);
nand U6766 (N_6766,N_6081,N_6224);
or U6767 (N_6767,N_6403,N_6307);
nand U6768 (N_6768,N_6001,N_6174);
xor U6769 (N_6769,N_6446,N_6437);
xor U6770 (N_6770,N_6265,N_6240);
or U6771 (N_6771,N_6436,N_6225);
or U6772 (N_6772,N_6394,N_6137);
xnor U6773 (N_6773,N_6257,N_6324);
or U6774 (N_6774,N_6043,N_6414);
xor U6775 (N_6775,N_6476,N_6008);
nor U6776 (N_6776,N_6366,N_6228);
and U6777 (N_6777,N_6243,N_6148);
xnor U6778 (N_6778,N_6173,N_6001);
and U6779 (N_6779,N_6060,N_6455);
nor U6780 (N_6780,N_6290,N_6060);
nor U6781 (N_6781,N_6268,N_6393);
nor U6782 (N_6782,N_6447,N_6126);
nand U6783 (N_6783,N_6251,N_6113);
nand U6784 (N_6784,N_6453,N_6427);
and U6785 (N_6785,N_6340,N_6226);
nand U6786 (N_6786,N_6281,N_6424);
nand U6787 (N_6787,N_6266,N_6402);
nor U6788 (N_6788,N_6038,N_6149);
or U6789 (N_6789,N_6431,N_6157);
nand U6790 (N_6790,N_6472,N_6308);
and U6791 (N_6791,N_6197,N_6292);
xor U6792 (N_6792,N_6403,N_6051);
nand U6793 (N_6793,N_6305,N_6005);
nor U6794 (N_6794,N_6153,N_6376);
and U6795 (N_6795,N_6201,N_6308);
nand U6796 (N_6796,N_6270,N_6430);
or U6797 (N_6797,N_6096,N_6107);
and U6798 (N_6798,N_6010,N_6015);
xnor U6799 (N_6799,N_6158,N_6138);
xnor U6800 (N_6800,N_6366,N_6093);
nor U6801 (N_6801,N_6266,N_6018);
nor U6802 (N_6802,N_6074,N_6459);
xor U6803 (N_6803,N_6137,N_6365);
and U6804 (N_6804,N_6423,N_6307);
nor U6805 (N_6805,N_6102,N_6430);
nand U6806 (N_6806,N_6177,N_6380);
nor U6807 (N_6807,N_6202,N_6375);
and U6808 (N_6808,N_6489,N_6117);
and U6809 (N_6809,N_6016,N_6251);
and U6810 (N_6810,N_6153,N_6234);
nand U6811 (N_6811,N_6408,N_6187);
nor U6812 (N_6812,N_6249,N_6223);
and U6813 (N_6813,N_6119,N_6142);
or U6814 (N_6814,N_6265,N_6172);
or U6815 (N_6815,N_6405,N_6079);
or U6816 (N_6816,N_6462,N_6062);
xor U6817 (N_6817,N_6375,N_6429);
nand U6818 (N_6818,N_6137,N_6499);
and U6819 (N_6819,N_6113,N_6435);
and U6820 (N_6820,N_6476,N_6449);
nand U6821 (N_6821,N_6165,N_6434);
nand U6822 (N_6822,N_6091,N_6173);
or U6823 (N_6823,N_6232,N_6076);
xor U6824 (N_6824,N_6443,N_6117);
nand U6825 (N_6825,N_6176,N_6141);
and U6826 (N_6826,N_6038,N_6283);
nand U6827 (N_6827,N_6321,N_6274);
and U6828 (N_6828,N_6215,N_6111);
nor U6829 (N_6829,N_6177,N_6379);
xor U6830 (N_6830,N_6024,N_6422);
or U6831 (N_6831,N_6456,N_6109);
or U6832 (N_6832,N_6331,N_6286);
nor U6833 (N_6833,N_6175,N_6124);
nand U6834 (N_6834,N_6472,N_6419);
and U6835 (N_6835,N_6272,N_6053);
or U6836 (N_6836,N_6370,N_6011);
nor U6837 (N_6837,N_6174,N_6094);
or U6838 (N_6838,N_6142,N_6028);
nand U6839 (N_6839,N_6489,N_6219);
nor U6840 (N_6840,N_6077,N_6043);
nand U6841 (N_6841,N_6452,N_6152);
nor U6842 (N_6842,N_6251,N_6105);
nand U6843 (N_6843,N_6419,N_6235);
xor U6844 (N_6844,N_6223,N_6190);
and U6845 (N_6845,N_6404,N_6023);
xnor U6846 (N_6846,N_6439,N_6051);
or U6847 (N_6847,N_6208,N_6359);
xor U6848 (N_6848,N_6071,N_6391);
nor U6849 (N_6849,N_6206,N_6032);
nand U6850 (N_6850,N_6116,N_6160);
and U6851 (N_6851,N_6309,N_6082);
or U6852 (N_6852,N_6465,N_6270);
xnor U6853 (N_6853,N_6249,N_6321);
xnor U6854 (N_6854,N_6327,N_6256);
and U6855 (N_6855,N_6356,N_6108);
and U6856 (N_6856,N_6030,N_6308);
or U6857 (N_6857,N_6215,N_6358);
xor U6858 (N_6858,N_6377,N_6241);
xnor U6859 (N_6859,N_6101,N_6241);
and U6860 (N_6860,N_6019,N_6204);
nor U6861 (N_6861,N_6028,N_6407);
xor U6862 (N_6862,N_6385,N_6286);
or U6863 (N_6863,N_6273,N_6253);
nand U6864 (N_6864,N_6273,N_6482);
and U6865 (N_6865,N_6337,N_6227);
nand U6866 (N_6866,N_6063,N_6108);
or U6867 (N_6867,N_6178,N_6354);
or U6868 (N_6868,N_6066,N_6405);
nand U6869 (N_6869,N_6071,N_6324);
nand U6870 (N_6870,N_6159,N_6016);
xor U6871 (N_6871,N_6256,N_6076);
nand U6872 (N_6872,N_6377,N_6437);
and U6873 (N_6873,N_6002,N_6075);
and U6874 (N_6874,N_6289,N_6151);
or U6875 (N_6875,N_6346,N_6032);
xor U6876 (N_6876,N_6210,N_6004);
nor U6877 (N_6877,N_6007,N_6140);
nor U6878 (N_6878,N_6170,N_6190);
or U6879 (N_6879,N_6223,N_6139);
nand U6880 (N_6880,N_6067,N_6018);
xor U6881 (N_6881,N_6228,N_6404);
xor U6882 (N_6882,N_6130,N_6039);
nor U6883 (N_6883,N_6273,N_6048);
nand U6884 (N_6884,N_6367,N_6385);
nand U6885 (N_6885,N_6401,N_6423);
xnor U6886 (N_6886,N_6138,N_6317);
and U6887 (N_6887,N_6346,N_6462);
xnor U6888 (N_6888,N_6455,N_6360);
xor U6889 (N_6889,N_6180,N_6004);
xnor U6890 (N_6890,N_6010,N_6277);
nor U6891 (N_6891,N_6492,N_6211);
nor U6892 (N_6892,N_6012,N_6251);
or U6893 (N_6893,N_6311,N_6193);
or U6894 (N_6894,N_6148,N_6476);
xnor U6895 (N_6895,N_6381,N_6151);
xnor U6896 (N_6896,N_6070,N_6188);
and U6897 (N_6897,N_6061,N_6212);
nand U6898 (N_6898,N_6069,N_6320);
or U6899 (N_6899,N_6175,N_6498);
nand U6900 (N_6900,N_6416,N_6214);
or U6901 (N_6901,N_6392,N_6426);
or U6902 (N_6902,N_6114,N_6039);
or U6903 (N_6903,N_6099,N_6410);
nand U6904 (N_6904,N_6100,N_6484);
nand U6905 (N_6905,N_6289,N_6433);
or U6906 (N_6906,N_6442,N_6305);
xnor U6907 (N_6907,N_6129,N_6205);
xor U6908 (N_6908,N_6087,N_6261);
or U6909 (N_6909,N_6038,N_6421);
or U6910 (N_6910,N_6101,N_6291);
or U6911 (N_6911,N_6279,N_6329);
and U6912 (N_6912,N_6182,N_6419);
or U6913 (N_6913,N_6026,N_6094);
nand U6914 (N_6914,N_6019,N_6148);
nor U6915 (N_6915,N_6051,N_6347);
and U6916 (N_6916,N_6431,N_6249);
xnor U6917 (N_6917,N_6391,N_6105);
nor U6918 (N_6918,N_6413,N_6427);
xnor U6919 (N_6919,N_6367,N_6415);
or U6920 (N_6920,N_6464,N_6030);
xor U6921 (N_6921,N_6224,N_6004);
nor U6922 (N_6922,N_6113,N_6227);
or U6923 (N_6923,N_6495,N_6174);
nor U6924 (N_6924,N_6398,N_6115);
and U6925 (N_6925,N_6222,N_6047);
and U6926 (N_6926,N_6405,N_6462);
nand U6927 (N_6927,N_6399,N_6104);
nor U6928 (N_6928,N_6298,N_6465);
nand U6929 (N_6929,N_6246,N_6448);
nand U6930 (N_6930,N_6407,N_6457);
or U6931 (N_6931,N_6326,N_6362);
and U6932 (N_6932,N_6142,N_6470);
or U6933 (N_6933,N_6099,N_6128);
and U6934 (N_6934,N_6131,N_6476);
nand U6935 (N_6935,N_6229,N_6474);
and U6936 (N_6936,N_6108,N_6381);
and U6937 (N_6937,N_6346,N_6343);
and U6938 (N_6938,N_6334,N_6134);
xnor U6939 (N_6939,N_6443,N_6402);
and U6940 (N_6940,N_6219,N_6477);
nand U6941 (N_6941,N_6414,N_6283);
or U6942 (N_6942,N_6214,N_6034);
nand U6943 (N_6943,N_6393,N_6010);
nand U6944 (N_6944,N_6478,N_6262);
nand U6945 (N_6945,N_6363,N_6250);
xnor U6946 (N_6946,N_6439,N_6245);
or U6947 (N_6947,N_6237,N_6233);
or U6948 (N_6948,N_6090,N_6307);
or U6949 (N_6949,N_6245,N_6277);
nand U6950 (N_6950,N_6188,N_6078);
nand U6951 (N_6951,N_6426,N_6149);
or U6952 (N_6952,N_6468,N_6185);
nand U6953 (N_6953,N_6175,N_6100);
and U6954 (N_6954,N_6291,N_6067);
nor U6955 (N_6955,N_6156,N_6172);
xnor U6956 (N_6956,N_6374,N_6070);
nor U6957 (N_6957,N_6302,N_6401);
xor U6958 (N_6958,N_6239,N_6206);
or U6959 (N_6959,N_6128,N_6056);
nor U6960 (N_6960,N_6163,N_6367);
or U6961 (N_6961,N_6087,N_6155);
or U6962 (N_6962,N_6363,N_6314);
or U6963 (N_6963,N_6474,N_6029);
nor U6964 (N_6964,N_6015,N_6215);
nor U6965 (N_6965,N_6043,N_6052);
and U6966 (N_6966,N_6243,N_6367);
nand U6967 (N_6967,N_6019,N_6143);
nor U6968 (N_6968,N_6408,N_6004);
nand U6969 (N_6969,N_6391,N_6049);
nor U6970 (N_6970,N_6219,N_6295);
nand U6971 (N_6971,N_6308,N_6098);
or U6972 (N_6972,N_6262,N_6373);
and U6973 (N_6973,N_6205,N_6431);
or U6974 (N_6974,N_6081,N_6182);
or U6975 (N_6975,N_6441,N_6442);
xor U6976 (N_6976,N_6293,N_6389);
and U6977 (N_6977,N_6082,N_6054);
and U6978 (N_6978,N_6371,N_6136);
and U6979 (N_6979,N_6367,N_6474);
nand U6980 (N_6980,N_6292,N_6426);
and U6981 (N_6981,N_6111,N_6084);
nand U6982 (N_6982,N_6218,N_6100);
and U6983 (N_6983,N_6225,N_6122);
nand U6984 (N_6984,N_6183,N_6217);
and U6985 (N_6985,N_6445,N_6072);
or U6986 (N_6986,N_6156,N_6253);
xnor U6987 (N_6987,N_6267,N_6236);
or U6988 (N_6988,N_6354,N_6467);
nand U6989 (N_6989,N_6407,N_6411);
nor U6990 (N_6990,N_6398,N_6227);
and U6991 (N_6991,N_6254,N_6271);
nor U6992 (N_6992,N_6356,N_6092);
nand U6993 (N_6993,N_6063,N_6168);
and U6994 (N_6994,N_6287,N_6277);
and U6995 (N_6995,N_6393,N_6349);
or U6996 (N_6996,N_6470,N_6112);
nor U6997 (N_6997,N_6476,N_6491);
nand U6998 (N_6998,N_6256,N_6290);
or U6999 (N_6999,N_6127,N_6312);
nor U7000 (N_7000,N_6661,N_6613);
xor U7001 (N_7001,N_6500,N_6952);
and U7002 (N_7002,N_6847,N_6505);
nand U7003 (N_7003,N_6854,N_6979);
xor U7004 (N_7004,N_6717,N_6513);
xor U7005 (N_7005,N_6758,N_6512);
nor U7006 (N_7006,N_6750,N_6808);
nand U7007 (N_7007,N_6871,N_6940);
nor U7008 (N_7008,N_6776,N_6915);
and U7009 (N_7009,N_6747,N_6653);
nand U7010 (N_7010,N_6627,N_6650);
nand U7011 (N_7011,N_6815,N_6555);
nand U7012 (N_7012,N_6752,N_6777);
nor U7013 (N_7013,N_6635,N_6867);
xnor U7014 (N_7014,N_6954,N_6936);
and U7015 (N_7015,N_6972,N_6585);
and U7016 (N_7016,N_6942,N_6925);
nor U7017 (N_7017,N_6764,N_6903);
xor U7018 (N_7018,N_6901,N_6893);
xnor U7019 (N_7019,N_6977,N_6608);
or U7020 (N_7020,N_6599,N_6892);
or U7021 (N_7021,N_6514,N_6891);
or U7022 (N_7022,N_6624,N_6506);
and U7023 (N_7023,N_6600,N_6788);
or U7024 (N_7024,N_6589,N_6987);
and U7025 (N_7025,N_6885,N_6775);
or U7026 (N_7026,N_6736,N_6767);
and U7027 (N_7027,N_6673,N_6548);
xnor U7028 (N_7028,N_6651,N_6643);
or U7029 (N_7029,N_6913,N_6830);
xnor U7030 (N_7030,N_6878,N_6601);
xor U7031 (N_7031,N_6754,N_6545);
and U7032 (N_7032,N_6943,N_6981);
and U7033 (N_7033,N_6700,N_6879);
or U7034 (N_7034,N_6660,N_6578);
nand U7035 (N_7035,N_6911,N_6848);
nor U7036 (N_7036,N_6739,N_6862);
and U7037 (N_7037,N_6733,N_6836);
and U7038 (N_7038,N_6725,N_6897);
xnor U7039 (N_7039,N_6706,N_6762);
and U7040 (N_7040,N_6611,N_6922);
or U7041 (N_7041,N_6842,N_6645);
nand U7042 (N_7042,N_6807,N_6692);
or U7043 (N_7043,N_6821,N_6993);
and U7044 (N_7044,N_6746,N_6701);
nand U7045 (N_7045,N_6953,N_6753);
nand U7046 (N_7046,N_6856,N_6667);
nand U7047 (N_7047,N_6845,N_6539);
and U7048 (N_7048,N_6959,N_6697);
or U7049 (N_7049,N_6751,N_6877);
nor U7050 (N_7050,N_6914,N_6960);
and U7051 (N_7051,N_6982,N_6898);
and U7052 (N_7052,N_6518,N_6698);
nand U7053 (N_7053,N_6694,N_6799);
nor U7054 (N_7054,N_6617,N_6742);
nor U7055 (N_7055,N_6865,N_6973);
and U7056 (N_7056,N_6787,N_6622);
nor U7057 (N_7057,N_6986,N_6850);
nor U7058 (N_7058,N_6665,N_6675);
or U7059 (N_7059,N_6681,N_6996);
nand U7060 (N_7060,N_6729,N_6592);
or U7061 (N_7061,N_6559,N_6588);
xnor U7062 (N_7062,N_6712,N_6796);
or U7063 (N_7063,N_6623,N_6679);
nand U7064 (N_7064,N_6540,N_6721);
nor U7065 (N_7065,N_6918,N_6929);
nor U7066 (N_7066,N_6519,N_6958);
or U7067 (N_7067,N_6761,N_6546);
nand U7068 (N_7068,N_6630,N_6510);
xor U7069 (N_7069,N_6833,N_6997);
nand U7070 (N_7070,N_6688,N_6772);
nand U7071 (N_7071,N_6852,N_6858);
xnor U7072 (N_7072,N_6726,N_6838);
nor U7073 (N_7073,N_6813,N_6535);
nor U7074 (N_7074,N_6794,N_6577);
xnor U7075 (N_7075,N_6648,N_6655);
nor U7076 (N_7076,N_6875,N_6948);
or U7077 (N_7077,N_6702,N_6735);
nor U7078 (N_7078,N_6992,N_6832);
and U7079 (N_7079,N_6872,N_6517);
and U7080 (N_7080,N_6586,N_6610);
nand U7081 (N_7081,N_6649,N_6839);
nor U7082 (N_7082,N_6511,N_6770);
nor U7083 (N_7083,N_6637,N_6786);
or U7084 (N_7084,N_6731,N_6704);
or U7085 (N_7085,N_6907,N_6890);
nand U7086 (N_7086,N_6967,N_6825);
nand U7087 (N_7087,N_6722,N_6990);
nor U7088 (N_7088,N_6521,N_6531);
nor U7089 (N_7089,N_6846,N_6920);
xnor U7090 (N_7090,N_6905,N_6949);
and U7091 (N_7091,N_6743,N_6507);
or U7092 (N_7092,N_6590,N_6549);
nand U7093 (N_7093,N_6989,N_6522);
and U7094 (N_7094,N_6502,N_6909);
xor U7095 (N_7095,N_6887,N_6889);
or U7096 (N_7096,N_6557,N_6961);
nand U7097 (N_7097,N_6594,N_6689);
nand U7098 (N_7098,N_6652,N_6827);
or U7099 (N_7099,N_6841,N_6816);
nand U7100 (N_7100,N_6537,N_6857);
xnor U7101 (N_7101,N_6570,N_6738);
nor U7102 (N_7102,N_6644,N_6716);
or U7103 (N_7103,N_6680,N_6760);
nor U7104 (N_7104,N_6790,N_6672);
xnor U7105 (N_7105,N_6793,N_6619);
xnor U7106 (N_7106,N_6873,N_6520);
or U7107 (N_7107,N_6656,N_6542);
nor U7108 (N_7108,N_6950,N_6902);
xor U7109 (N_7109,N_6646,N_6945);
nor U7110 (N_7110,N_6628,N_6564);
xor U7111 (N_7111,N_6525,N_6550);
nand U7112 (N_7112,N_6809,N_6921);
and U7113 (N_7113,N_6598,N_6917);
and U7114 (N_7114,N_6806,N_6639);
or U7115 (N_7115,N_6554,N_6558);
nand U7116 (N_7116,N_6626,N_6625);
or U7117 (N_7117,N_6831,N_6844);
xor U7118 (N_7118,N_6884,N_6551);
nor U7119 (N_7119,N_6713,N_6855);
nor U7120 (N_7120,N_6863,N_6591);
nand U7121 (N_7121,N_6965,N_6869);
nand U7122 (N_7122,N_6523,N_6524);
nand U7123 (N_7123,N_6533,N_6923);
nor U7124 (N_7124,N_6781,N_6937);
or U7125 (N_7125,N_6640,N_6971);
and U7126 (N_7126,N_6593,N_6998);
nand U7127 (N_7127,N_6866,N_6853);
nor U7128 (N_7128,N_6868,N_6620);
nor U7129 (N_7129,N_6552,N_6924);
and U7130 (N_7130,N_6707,N_6566);
nor U7131 (N_7131,N_6562,N_6976);
nand U7132 (N_7132,N_6941,N_6951);
and U7133 (N_7133,N_6730,N_6603);
nand U7134 (N_7134,N_6567,N_6536);
or U7135 (N_7135,N_6759,N_6723);
nand U7136 (N_7136,N_6840,N_6974);
xnor U7137 (N_7137,N_6851,N_6740);
nand U7138 (N_7138,N_6561,N_6933);
xnor U7139 (N_7139,N_6744,N_6718);
and U7140 (N_7140,N_6538,N_6828);
nor U7141 (N_7141,N_6876,N_6978);
or U7142 (N_7142,N_6789,N_6768);
xor U7143 (N_7143,N_6607,N_6931);
or U7144 (N_7144,N_6671,N_6774);
and U7145 (N_7145,N_6573,N_6529);
or U7146 (N_7146,N_6532,N_6810);
nor U7147 (N_7147,N_6835,N_6677);
xor U7148 (N_7148,N_6727,N_6666);
xnor U7149 (N_7149,N_6970,N_6882);
xor U7150 (N_7150,N_6800,N_6817);
nand U7151 (N_7151,N_6843,N_6896);
nor U7152 (N_7152,N_6894,N_6895);
nor U7153 (N_7153,N_6629,N_6888);
nand U7154 (N_7154,N_6528,N_6811);
nor U7155 (N_7155,N_6597,N_6690);
xnor U7156 (N_7156,N_6957,N_6930);
and U7157 (N_7157,N_6568,N_6544);
and U7158 (N_7158,N_6955,N_6691);
xnor U7159 (N_7159,N_6822,N_6814);
xnor U7160 (N_7160,N_6820,N_6926);
and U7161 (N_7161,N_6994,N_6596);
nand U7162 (N_7162,N_6874,N_6859);
nand U7163 (N_7163,N_6633,N_6670);
or U7164 (N_7164,N_6612,N_6734);
or U7165 (N_7165,N_6720,N_6964);
nand U7166 (N_7166,N_6654,N_6501);
xnor U7167 (N_7167,N_6695,N_6966);
and U7168 (N_7168,N_6693,N_6678);
or U7169 (N_7169,N_6543,N_6985);
xnor U7170 (N_7170,N_6826,N_6582);
nor U7171 (N_7171,N_6969,N_6860);
xnor U7172 (N_7172,N_6527,N_6580);
and U7173 (N_7173,N_6780,N_6946);
or U7174 (N_7174,N_6968,N_6980);
nor U7175 (N_7175,N_6685,N_6906);
or U7176 (N_7176,N_6636,N_6638);
or U7177 (N_7177,N_6728,N_6908);
and U7178 (N_7178,N_6984,N_6687);
nand U7179 (N_7179,N_6668,N_6824);
and U7180 (N_7180,N_6745,N_6516);
xor U7181 (N_7181,N_6900,N_6797);
xor U7182 (N_7182,N_6615,N_6932);
and U7183 (N_7183,N_6834,N_6703);
nand U7184 (N_7184,N_6662,N_6642);
nand U7185 (N_7185,N_6579,N_6604);
xor U7186 (N_7186,N_6515,N_6837);
and U7187 (N_7187,N_6975,N_6609);
or U7188 (N_7188,N_6556,N_6983);
or U7189 (N_7189,N_6696,N_6686);
xor U7190 (N_7190,N_6802,N_6783);
nand U7191 (N_7191,N_6553,N_6880);
nand U7192 (N_7192,N_6618,N_6769);
or U7193 (N_7193,N_6805,N_6583);
xor U7194 (N_7194,N_6748,N_6616);
nor U7195 (N_7195,N_6503,N_6883);
nand U7196 (N_7196,N_6711,N_6658);
nor U7197 (N_7197,N_6910,N_6547);
and U7198 (N_7198,N_6504,N_6795);
nor U7199 (N_7199,N_6664,N_6741);
and U7200 (N_7200,N_6714,N_6676);
xnor U7201 (N_7201,N_6999,N_6939);
and U7202 (N_7202,N_6763,N_6732);
xor U7203 (N_7203,N_6715,N_6563);
xor U7204 (N_7204,N_6757,N_6791);
nor U7205 (N_7205,N_6614,N_6634);
nand U7206 (N_7206,N_6509,N_6779);
nand U7207 (N_7207,N_6581,N_6935);
or U7208 (N_7208,N_6773,N_6621);
and U7209 (N_7209,N_6541,N_6881);
nand U7210 (N_7210,N_6803,N_6756);
xnor U7211 (N_7211,N_6899,N_6595);
xnor U7212 (N_7212,N_6904,N_6684);
nor U7213 (N_7213,N_6699,N_6919);
nand U7214 (N_7214,N_6765,N_6705);
and U7215 (N_7215,N_6916,N_6801);
xor U7216 (N_7216,N_6606,N_6576);
and U7217 (N_7217,N_6560,N_6708);
nor U7218 (N_7218,N_6755,N_6778);
or U7219 (N_7219,N_6962,N_6647);
nand U7220 (N_7220,N_6819,N_6737);
nor U7221 (N_7221,N_6572,N_6912);
nor U7222 (N_7222,N_6766,N_6938);
nand U7223 (N_7223,N_6927,N_6657);
nand U7224 (N_7224,N_6864,N_6571);
or U7225 (N_7225,N_6575,N_6792);
xor U7226 (N_7226,N_6818,N_6632);
xnor U7227 (N_7227,N_6988,N_6956);
nand U7228 (N_7228,N_6641,N_6928);
xor U7229 (N_7229,N_6823,N_6674);
nand U7230 (N_7230,N_6812,N_6569);
and U7231 (N_7231,N_6719,N_6602);
nand U7232 (N_7232,N_6782,N_6829);
nand U7233 (N_7233,N_6995,N_6631);
nor U7234 (N_7234,N_6870,N_6771);
nor U7235 (N_7235,N_6530,N_6710);
or U7236 (N_7236,N_6724,N_6508);
or U7237 (N_7237,N_6663,N_6534);
xnor U7238 (N_7238,N_6934,N_6784);
xnor U7239 (N_7239,N_6574,N_6659);
and U7240 (N_7240,N_6749,N_6804);
or U7241 (N_7241,N_6849,N_6587);
and U7242 (N_7242,N_6991,N_6526);
or U7243 (N_7243,N_6963,N_6709);
nand U7244 (N_7244,N_6683,N_6785);
nor U7245 (N_7245,N_6947,N_6682);
nand U7246 (N_7246,N_6944,N_6861);
or U7247 (N_7247,N_6584,N_6565);
nand U7248 (N_7248,N_6886,N_6605);
and U7249 (N_7249,N_6798,N_6669);
xnor U7250 (N_7250,N_6969,N_6982);
nand U7251 (N_7251,N_6692,N_6905);
or U7252 (N_7252,N_6746,N_6749);
xor U7253 (N_7253,N_6731,N_6932);
xnor U7254 (N_7254,N_6810,N_6669);
nand U7255 (N_7255,N_6677,N_6772);
nor U7256 (N_7256,N_6947,N_6973);
and U7257 (N_7257,N_6577,N_6640);
nand U7258 (N_7258,N_6691,N_6650);
or U7259 (N_7259,N_6788,N_6512);
nor U7260 (N_7260,N_6637,N_6829);
or U7261 (N_7261,N_6724,N_6947);
and U7262 (N_7262,N_6892,N_6797);
or U7263 (N_7263,N_6804,N_6611);
nor U7264 (N_7264,N_6651,N_6568);
or U7265 (N_7265,N_6848,N_6619);
or U7266 (N_7266,N_6688,N_6727);
or U7267 (N_7267,N_6697,N_6552);
nand U7268 (N_7268,N_6909,N_6611);
nor U7269 (N_7269,N_6880,N_6872);
nor U7270 (N_7270,N_6888,N_6568);
nand U7271 (N_7271,N_6506,N_6761);
or U7272 (N_7272,N_6850,N_6871);
nor U7273 (N_7273,N_6553,N_6930);
and U7274 (N_7274,N_6845,N_6570);
or U7275 (N_7275,N_6850,N_6714);
and U7276 (N_7276,N_6793,N_6783);
and U7277 (N_7277,N_6530,N_6769);
xor U7278 (N_7278,N_6938,N_6508);
xnor U7279 (N_7279,N_6627,N_6500);
xnor U7280 (N_7280,N_6697,N_6977);
xnor U7281 (N_7281,N_6557,N_6968);
and U7282 (N_7282,N_6795,N_6973);
nor U7283 (N_7283,N_6743,N_6871);
or U7284 (N_7284,N_6547,N_6960);
xor U7285 (N_7285,N_6771,N_6817);
nand U7286 (N_7286,N_6809,N_6788);
nand U7287 (N_7287,N_6943,N_6932);
nor U7288 (N_7288,N_6898,N_6583);
xnor U7289 (N_7289,N_6903,N_6875);
or U7290 (N_7290,N_6870,N_6577);
nor U7291 (N_7291,N_6904,N_6956);
and U7292 (N_7292,N_6542,N_6541);
nor U7293 (N_7293,N_6720,N_6835);
nand U7294 (N_7294,N_6529,N_6596);
or U7295 (N_7295,N_6987,N_6945);
and U7296 (N_7296,N_6987,N_6952);
nand U7297 (N_7297,N_6684,N_6626);
or U7298 (N_7298,N_6948,N_6930);
nor U7299 (N_7299,N_6705,N_6731);
nand U7300 (N_7300,N_6840,N_6533);
or U7301 (N_7301,N_6866,N_6771);
nor U7302 (N_7302,N_6696,N_6733);
and U7303 (N_7303,N_6529,N_6977);
nand U7304 (N_7304,N_6750,N_6966);
nand U7305 (N_7305,N_6924,N_6889);
or U7306 (N_7306,N_6587,N_6829);
xor U7307 (N_7307,N_6923,N_6651);
xor U7308 (N_7308,N_6786,N_6671);
nand U7309 (N_7309,N_6995,N_6683);
xnor U7310 (N_7310,N_6866,N_6712);
nand U7311 (N_7311,N_6727,N_6586);
nor U7312 (N_7312,N_6581,N_6535);
xnor U7313 (N_7313,N_6609,N_6775);
xnor U7314 (N_7314,N_6983,N_6610);
and U7315 (N_7315,N_6973,N_6620);
nand U7316 (N_7316,N_6991,N_6950);
or U7317 (N_7317,N_6743,N_6982);
and U7318 (N_7318,N_6652,N_6596);
xor U7319 (N_7319,N_6946,N_6977);
and U7320 (N_7320,N_6777,N_6740);
or U7321 (N_7321,N_6678,N_6971);
nand U7322 (N_7322,N_6798,N_6793);
or U7323 (N_7323,N_6906,N_6750);
and U7324 (N_7324,N_6673,N_6944);
or U7325 (N_7325,N_6644,N_6753);
nand U7326 (N_7326,N_6881,N_6917);
xor U7327 (N_7327,N_6619,N_6852);
xnor U7328 (N_7328,N_6557,N_6879);
or U7329 (N_7329,N_6730,N_6809);
and U7330 (N_7330,N_6682,N_6510);
nor U7331 (N_7331,N_6519,N_6817);
nor U7332 (N_7332,N_6558,N_6519);
xnor U7333 (N_7333,N_6510,N_6920);
or U7334 (N_7334,N_6588,N_6537);
nand U7335 (N_7335,N_6579,N_6501);
or U7336 (N_7336,N_6764,N_6693);
nor U7337 (N_7337,N_6779,N_6581);
nor U7338 (N_7338,N_6967,N_6933);
or U7339 (N_7339,N_6938,N_6875);
xor U7340 (N_7340,N_6704,N_6784);
nor U7341 (N_7341,N_6955,N_6932);
nand U7342 (N_7342,N_6535,N_6790);
nor U7343 (N_7343,N_6976,N_6802);
and U7344 (N_7344,N_6777,N_6614);
or U7345 (N_7345,N_6929,N_6800);
nor U7346 (N_7346,N_6659,N_6754);
xor U7347 (N_7347,N_6517,N_6912);
nand U7348 (N_7348,N_6748,N_6747);
nor U7349 (N_7349,N_6532,N_6505);
xnor U7350 (N_7350,N_6758,N_6837);
nor U7351 (N_7351,N_6728,N_6559);
nor U7352 (N_7352,N_6614,N_6621);
nor U7353 (N_7353,N_6612,N_6909);
or U7354 (N_7354,N_6945,N_6537);
nand U7355 (N_7355,N_6951,N_6639);
nand U7356 (N_7356,N_6866,N_6944);
and U7357 (N_7357,N_6727,N_6525);
nand U7358 (N_7358,N_6742,N_6532);
or U7359 (N_7359,N_6567,N_6946);
or U7360 (N_7360,N_6795,N_6774);
and U7361 (N_7361,N_6609,N_6987);
nand U7362 (N_7362,N_6813,N_6790);
nor U7363 (N_7363,N_6997,N_6928);
or U7364 (N_7364,N_6758,N_6605);
and U7365 (N_7365,N_6988,N_6548);
and U7366 (N_7366,N_6612,N_6939);
and U7367 (N_7367,N_6924,N_6682);
nand U7368 (N_7368,N_6709,N_6873);
and U7369 (N_7369,N_6590,N_6741);
xnor U7370 (N_7370,N_6792,N_6893);
and U7371 (N_7371,N_6914,N_6872);
nand U7372 (N_7372,N_6610,N_6772);
nand U7373 (N_7373,N_6956,N_6747);
nor U7374 (N_7374,N_6928,N_6653);
nor U7375 (N_7375,N_6560,N_6518);
or U7376 (N_7376,N_6715,N_6513);
xor U7377 (N_7377,N_6614,N_6561);
nand U7378 (N_7378,N_6621,N_6680);
nor U7379 (N_7379,N_6936,N_6999);
or U7380 (N_7380,N_6666,N_6767);
nor U7381 (N_7381,N_6813,N_6690);
or U7382 (N_7382,N_6700,N_6897);
nor U7383 (N_7383,N_6745,N_6721);
and U7384 (N_7384,N_6667,N_6852);
nand U7385 (N_7385,N_6514,N_6699);
or U7386 (N_7386,N_6904,N_6858);
nand U7387 (N_7387,N_6652,N_6921);
and U7388 (N_7388,N_6772,N_6605);
or U7389 (N_7389,N_6698,N_6688);
nand U7390 (N_7390,N_6937,N_6544);
nor U7391 (N_7391,N_6583,N_6835);
nor U7392 (N_7392,N_6545,N_6673);
or U7393 (N_7393,N_6622,N_6628);
nor U7394 (N_7394,N_6643,N_6712);
or U7395 (N_7395,N_6500,N_6890);
or U7396 (N_7396,N_6789,N_6650);
nand U7397 (N_7397,N_6620,N_6925);
nand U7398 (N_7398,N_6931,N_6534);
xor U7399 (N_7399,N_6543,N_6655);
and U7400 (N_7400,N_6638,N_6595);
nor U7401 (N_7401,N_6878,N_6571);
xor U7402 (N_7402,N_6832,N_6626);
or U7403 (N_7403,N_6738,N_6582);
xnor U7404 (N_7404,N_6642,N_6790);
nand U7405 (N_7405,N_6512,N_6886);
xor U7406 (N_7406,N_6761,N_6782);
nand U7407 (N_7407,N_6513,N_6708);
nor U7408 (N_7408,N_6569,N_6529);
xnor U7409 (N_7409,N_6962,N_6930);
or U7410 (N_7410,N_6948,N_6641);
nand U7411 (N_7411,N_6564,N_6671);
xor U7412 (N_7412,N_6690,N_6534);
nand U7413 (N_7413,N_6862,N_6909);
nand U7414 (N_7414,N_6567,N_6671);
or U7415 (N_7415,N_6939,N_6824);
or U7416 (N_7416,N_6674,N_6888);
nor U7417 (N_7417,N_6872,N_6989);
and U7418 (N_7418,N_6852,N_6905);
xnor U7419 (N_7419,N_6896,N_6849);
xor U7420 (N_7420,N_6756,N_6644);
and U7421 (N_7421,N_6520,N_6566);
xor U7422 (N_7422,N_6591,N_6623);
nor U7423 (N_7423,N_6697,N_6696);
or U7424 (N_7424,N_6800,N_6509);
and U7425 (N_7425,N_6966,N_6709);
nor U7426 (N_7426,N_6765,N_6754);
or U7427 (N_7427,N_6944,N_6528);
nand U7428 (N_7428,N_6802,N_6995);
xnor U7429 (N_7429,N_6636,N_6777);
or U7430 (N_7430,N_6959,N_6717);
or U7431 (N_7431,N_6641,N_6909);
nor U7432 (N_7432,N_6547,N_6663);
nand U7433 (N_7433,N_6682,N_6706);
nand U7434 (N_7434,N_6756,N_6885);
nand U7435 (N_7435,N_6942,N_6676);
xor U7436 (N_7436,N_6591,N_6665);
nand U7437 (N_7437,N_6917,N_6566);
and U7438 (N_7438,N_6796,N_6879);
xnor U7439 (N_7439,N_6630,N_6857);
nand U7440 (N_7440,N_6539,N_6883);
nor U7441 (N_7441,N_6994,N_6584);
or U7442 (N_7442,N_6565,N_6818);
xor U7443 (N_7443,N_6939,N_6699);
or U7444 (N_7444,N_6816,N_6583);
nand U7445 (N_7445,N_6632,N_6953);
and U7446 (N_7446,N_6808,N_6619);
nand U7447 (N_7447,N_6906,N_6930);
nand U7448 (N_7448,N_6849,N_6800);
or U7449 (N_7449,N_6965,N_6523);
xor U7450 (N_7450,N_6732,N_6618);
nor U7451 (N_7451,N_6849,N_6660);
nor U7452 (N_7452,N_6650,N_6790);
and U7453 (N_7453,N_6562,N_6665);
nor U7454 (N_7454,N_6847,N_6740);
nor U7455 (N_7455,N_6695,N_6944);
xor U7456 (N_7456,N_6678,N_6714);
nor U7457 (N_7457,N_6819,N_6563);
or U7458 (N_7458,N_6847,N_6722);
nor U7459 (N_7459,N_6507,N_6930);
and U7460 (N_7460,N_6703,N_6956);
nand U7461 (N_7461,N_6976,N_6676);
and U7462 (N_7462,N_6906,N_6873);
xor U7463 (N_7463,N_6792,N_6623);
or U7464 (N_7464,N_6703,N_6728);
or U7465 (N_7465,N_6504,N_6586);
nor U7466 (N_7466,N_6789,N_6728);
or U7467 (N_7467,N_6993,N_6646);
or U7468 (N_7468,N_6929,N_6746);
nor U7469 (N_7469,N_6623,N_6948);
or U7470 (N_7470,N_6505,N_6790);
xor U7471 (N_7471,N_6749,N_6748);
and U7472 (N_7472,N_6985,N_6726);
nand U7473 (N_7473,N_6868,N_6812);
or U7474 (N_7474,N_6550,N_6534);
or U7475 (N_7475,N_6679,N_6605);
nand U7476 (N_7476,N_6911,N_6847);
and U7477 (N_7477,N_6919,N_6609);
or U7478 (N_7478,N_6587,N_6728);
xnor U7479 (N_7479,N_6672,N_6512);
and U7480 (N_7480,N_6535,N_6972);
nand U7481 (N_7481,N_6863,N_6524);
nor U7482 (N_7482,N_6859,N_6976);
xor U7483 (N_7483,N_6643,N_6767);
nand U7484 (N_7484,N_6824,N_6606);
nand U7485 (N_7485,N_6795,N_6946);
xnor U7486 (N_7486,N_6921,N_6773);
nand U7487 (N_7487,N_6752,N_6729);
nand U7488 (N_7488,N_6801,N_6931);
and U7489 (N_7489,N_6529,N_6730);
and U7490 (N_7490,N_6598,N_6965);
or U7491 (N_7491,N_6904,N_6652);
xnor U7492 (N_7492,N_6580,N_6641);
nor U7493 (N_7493,N_6667,N_6560);
and U7494 (N_7494,N_6501,N_6525);
nand U7495 (N_7495,N_6852,N_6560);
nor U7496 (N_7496,N_6677,N_6528);
or U7497 (N_7497,N_6699,N_6556);
and U7498 (N_7498,N_6539,N_6729);
and U7499 (N_7499,N_6742,N_6857);
nor U7500 (N_7500,N_7188,N_7157);
nand U7501 (N_7501,N_7449,N_7498);
and U7502 (N_7502,N_7235,N_7306);
xor U7503 (N_7503,N_7073,N_7028);
nor U7504 (N_7504,N_7411,N_7171);
xnor U7505 (N_7505,N_7030,N_7489);
xnor U7506 (N_7506,N_7197,N_7384);
nor U7507 (N_7507,N_7420,N_7187);
nand U7508 (N_7508,N_7365,N_7205);
nor U7509 (N_7509,N_7457,N_7417);
and U7510 (N_7510,N_7275,N_7447);
nand U7511 (N_7511,N_7196,N_7353);
nand U7512 (N_7512,N_7361,N_7139);
and U7513 (N_7513,N_7122,N_7403);
or U7514 (N_7514,N_7112,N_7283);
and U7515 (N_7515,N_7305,N_7439);
nand U7516 (N_7516,N_7227,N_7085);
and U7517 (N_7517,N_7102,N_7047);
nor U7518 (N_7518,N_7321,N_7001);
nor U7519 (N_7519,N_7100,N_7156);
nand U7520 (N_7520,N_7201,N_7036);
xor U7521 (N_7521,N_7468,N_7237);
nor U7522 (N_7522,N_7229,N_7163);
xor U7523 (N_7523,N_7445,N_7425);
nand U7524 (N_7524,N_7183,N_7109);
and U7525 (N_7525,N_7376,N_7071);
nor U7526 (N_7526,N_7140,N_7180);
nor U7527 (N_7527,N_7477,N_7082);
nand U7528 (N_7528,N_7089,N_7147);
or U7529 (N_7529,N_7342,N_7162);
and U7530 (N_7530,N_7459,N_7209);
nand U7531 (N_7531,N_7350,N_7182);
or U7532 (N_7532,N_7255,N_7118);
nand U7533 (N_7533,N_7474,N_7159);
and U7534 (N_7534,N_7366,N_7007);
nor U7535 (N_7535,N_7479,N_7000);
or U7536 (N_7536,N_7079,N_7240);
or U7537 (N_7537,N_7480,N_7331);
nor U7538 (N_7538,N_7228,N_7189);
xor U7539 (N_7539,N_7055,N_7057);
or U7540 (N_7540,N_7370,N_7110);
nand U7541 (N_7541,N_7203,N_7127);
or U7542 (N_7542,N_7276,N_7048);
xor U7543 (N_7543,N_7388,N_7026);
nand U7544 (N_7544,N_7216,N_7263);
nand U7545 (N_7545,N_7052,N_7031);
nor U7546 (N_7546,N_7322,N_7400);
and U7547 (N_7547,N_7021,N_7387);
nor U7548 (N_7548,N_7349,N_7446);
and U7549 (N_7549,N_7485,N_7016);
and U7550 (N_7550,N_7272,N_7310);
xor U7551 (N_7551,N_7015,N_7087);
xor U7552 (N_7552,N_7280,N_7393);
or U7553 (N_7553,N_7409,N_7222);
or U7554 (N_7554,N_7399,N_7499);
nand U7555 (N_7555,N_7179,N_7098);
xnor U7556 (N_7556,N_7101,N_7287);
and U7557 (N_7557,N_7012,N_7492);
xor U7558 (N_7558,N_7056,N_7105);
or U7559 (N_7559,N_7076,N_7049);
nor U7560 (N_7560,N_7160,N_7313);
xor U7561 (N_7561,N_7435,N_7029);
and U7562 (N_7562,N_7017,N_7174);
nand U7563 (N_7563,N_7264,N_7300);
xnor U7564 (N_7564,N_7067,N_7151);
or U7565 (N_7565,N_7131,N_7330);
nand U7566 (N_7566,N_7362,N_7319);
or U7567 (N_7567,N_7221,N_7438);
or U7568 (N_7568,N_7194,N_7359);
and U7569 (N_7569,N_7153,N_7311);
and U7570 (N_7570,N_7486,N_7185);
and U7571 (N_7571,N_7422,N_7238);
and U7572 (N_7572,N_7317,N_7066);
nor U7573 (N_7573,N_7195,N_7137);
nand U7574 (N_7574,N_7234,N_7011);
xor U7575 (N_7575,N_7148,N_7415);
or U7576 (N_7576,N_7441,N_7009);
or U7577 (N_7577,N_7471,N_7404);
and U7578 (N_7578,N_7285,N_7249);
nor U7579 (N_7579,N_7394,N_7230);
xnor U7580 (N_7580,N_7382,N_7368);
nand U7581 (N_7581,N_7242,N_7419);
or U7582 (N_7582,N_7466,N_7129);
or U7583 (N_7583,N_7490,N_7142);
nor U7584 (N_7584,N_7429,N_7337);
nand U7585 (N_7585,N_7473,N_7476);
nand U7586 (N_7586,N_7274,N_7440);
and U7587 (N_7587,N_7080,N_7236);
or U7588 (N_7588,N_7231,N_7309);
nor U7589 (N_7589,N_7020,N_7006);
or U7590 (N_7590,N_7223,N_7314);
nor U7591 (N_7591,N_7053,N_7124);
xor U7592 (N_7592,N_7482,N_7074);
nor U7593 (N_7593,N_7024,N_7428);
xor U7594 (N_7594,N_7130,N_7186);
xor U7595 (N_7595,N_7348,N_7025);
and U7596 (N_7596,N_7450,N_7093);
and U7597 (N_7597,N_7347,N_7323);
and U7598 (N_7598,N_7418,N_7041);
nand U7599 (N_7599,N_7448,N_7345);
nor U7600 (N_7600,N_7005,N_7010);
xnor U7601 (N_7601,N_7412,N_7068);
xnor U7602 (N_7602,N_7246,N_7308);
nand U7603 (N_7603,N_7371,N_7161);
and U7604 (N_7604,N_7072,N_7108);
and U7605 (N_7605,N_7135,N_7475);
xnor U7606 (N_7606,N_7051,N_7256);
nand U7607 (N_7607,N_7250,N_7279);
nand U7608 (N_7608,N_7232,N_7324);
and U7609 (N_7609,N_7431,N_7369);
nand U7610 (N_7610,N_7455,N_7251);
or U7611 (N_7611,N_7270,N_7291);
or U7612 (N_7612,N_7225,N_7226);
xor U7613 (N_7613,N_7396,N_7217);
or U7614 (N_7614,N_7367,N_7451);
nand U7615 (N_7615,N_7248,N_7060);
nor U7616 (N_7616,N_7470,N_7289);
nor U7617 (N_7617,N_7346,N_7019);
xor U7618 (N_7618,N_7304,N_7106);
nor U7619 (N_7619,N_7293,N_7042);
or U7620 (N_7620,N_7332,N_7372);
xnor U7621 (N_7621,N_7063,N_7261);
nor U7622 (N_7622,N_7004,N_7172);
nor U7623 (N_7623,N_7084,N_7046);
and U7624 (N_7624,N_7333,N_7117);
and U7625 (N_7625,N_7318,N_7401);
or U7626 (N_7626,N_7436,N_7344);
nand U7627 (N_7627,N_7043,N_7104);
or U7628 (N_7628,N_7444,N_7290);
nor U7629 (N_7629,N_7266,N_7136);
xnor U7630 (N_7630,N_7096,N_7391);
or U7631 (N_7631,N_7430,N_7335);
and U7632 (N_7632,N_7247,N_7037);
nor U7633 (N_7633,N_7132,N_7107);
xnor U7634 (N_7634,N_7325,N_7395);
nand U7635 (N_7635,N_7058,N_7038);
or U7636 (N_7636,N_7111,N_7408);
nand U7637 (N_7637,N_7421,N_7336);
nand U7638 (N_7638,N_7214,N_7297);
xor U7639 (N_7639,N_7352,N_7478);
xor U7640 (N_7640,N_7464,N_7392);
or U7641 (N_7641,N_7390,N_7040);
nand U7642 (N_7642,N_7032,N_7341);
and U7643 (N_7643,N_7168,N_7152);
xor U7644 (N_7644,N_7339,N_7095);
and U7645 (N_7645,N_7113,N_7302);
nor U7646 (N_7646,N_7364,N_7062);
nor U7647 (N_7647,N_7167,N_7338);
nand U7648 (N_7648,N_7181,N_7045);
nor U7649 (N_7649,N_7363,N_7134);
nand U7650 (N_7650,N_7259,N_7407);
or U7651 (N_7651,N_7061,N_7257);
or U7652 (N_7652,N_7427,N_7375);
and U7653 (N_7653,N_7312,N_7343);
nand U7654 (N_7654,N_7078,N_7269);
xnor U7655 (N_7655,N_7398,N_7402);
or U7656 (N_7656,N_7299,N_7145);
or U7657 (N_7657,N_7410,N_7383);
nand U7658 (N_7658,N_7380,N_7433);
or U7659 (N_7659,N_7386,N_7358);
and U7660 (N_7660,N_7355,N_7220);
and U7661 (N_7661,N_7483,N_7158);
and U7662 (N_7662,N_7405,N_7044);
nor U7663 (N_7663,N_7138,N_7200);
or U7664 (N_7664,N_7496,N_7090);
nand U7665 (N_7665,N_7146,N_7334);
nand U7666 (N_7666,N_7059,N_7092);
xor U7667 (N_7667,N_7193,N_7245);
xnor U7668 (N_7668,N_7469,N_7281);
xor U7669 (N_7669,N_7003,N_7088);
xor U7670 (N_7670,N_7170,N_7277);
and U7671 (N_7671,N_7065,N_7284);
or U7672 (N_7672,N_7144,N_7351);
and U7673 (N_7673,N_7219,N_7320);
nand U7674 (N_7674,N_7099,N_7303);
xor U7675 (N_7675,N_7199,N_7260);
nand U7676 (N_7676,N_7416,N_7206);
nand U7677 (N_7677,N_7120,N_7125);
and U7678 (N_7678,N_7215,N_7452);
or U7679 (N_7679,N_7064,N_7211);
nor U7680 (N_7680,N_7443,N_7212);
and U7681 (N_7681,N_7273,N_7022);
and U7682 (N_7682,N_7296,N_7002);
nand U7683 (N_7683,N_7115,N_7282);
and U7684 (N_7684,N_7315,N_7258);
or U7685 (N_7685,N_7208,N_7097);
nand U7686 (N_7686,N_7233,N_7295);
nand U7687 (N_7687,N_7434,N_7150);
or U7688 (N_7688,N_7262,N_7463);
and U7689 (N_7689,N_7141,N_7178);
xnor U7690 (N_7690,N_7424,N_7243);
and U7691 (N_7691,N_7373,N_7207);
nor U7692 (N_7692,N_7488,N_7378);
and U7693 (N_7693,N_7191,N_7294);
nand U7694 (N_7694,N_7354,N_7442);
or U7695 (N_7695,N_7128,N_7327);
or U7696 (N_7696,N_7497,N_7091);
and U7697 (N_7697,N_7173,N_7176);
and U7698 (N_7698,N_7267,N_7385);
or U7699 (N_7699,N_7379,N_7495);
or U7700 (N_7700,N_7184,N_7213);
or U7701 (N_7701,N_7414,N_7119);
nor U7702 (N_7702,N_7461,N_7406);
and U7703 (N_7703,N_7081,N_7177);
and U7704 (N_7704,N_7192,N_7288);
nand U7705 (N_7705,N_7437,N_7083);
or U7706 (N_7706,N_7491,N_7123);
nand U7707 (N_7707,N_7204,N_7316);
nand U7708 (N_7708,N_7286,N_7397);
nand U7709 (N_7709,N_7298,N_7094);
and U7710 (N_7710,N_7114,N_7426);
nor U7711 (N_7711,N_7301,N_7175);
xnor U7712 (N_7712,N_7121,N_7077);
nor U7713 (N_7713,N_7413,N_7472);
nand U7714 (N_7714,N_7155,N_7018);
nor U7715 (N_7715,N_7070,N_7166);
or U7716 (N_7716,N_7169,N_7481);
xnor U7717 (N_7717,N_7035,N_7462);
nor U7718 (N_7718,N_7218,N_7357);
and U7719 (N_7719,N_7487,N_7014);
nand U7720 (N_7720,N_7253,N_7467);
or U7721 (N_7721,N_7271,N_7086);
nor U7722 (N_7722,N_7252,N_7224);
xor U7723 (N_7723,N_7493,N_7154);
xor U7724 (N_7724,N_7292,N_7165);
xnor U7725 (N_7725,N_7143,N_7494);
or U7726 (N_7726,N_7307,N_7356);
xnor U7727 (N_7727,N_7198,N_7239);
nand U7728 (N_7728,N_7484,N_7126);
or U7729 (N_7729,N_7268,N_7432);
or U7730 (N_7730,N_7133,N_7069);
and U7731 (N_7731,N_7458,N_7050);
or U7732 (N_7732,N_7202,N_7039);
xnor U7733 (N_7733,N_7326,N_7008);
and U7734 (N_7734,N_7075,N_7265);
nor U7735 (N_7735,N_7456,N_7103);
nor U7736 (N_7736,N_7244,N_7460);
xnor U7737 (N_7737,N_7340,N_7465);
and U7738 (N_7738,N_7190,N_7116);
or U7739 (N_7739,N_7033,N_7210);
nor U7740 (N_7740,N_7054,N_7389);
and U7741 (N_7741,N_7374,N_7377);
or U7742 (N_7742,N_7423,N_7453);
or U7743 (N_7743,N_7328,N_7360);
or U7744 (N_7744,N_7149,N_7278);
and U7745 (N_7745,N_7381,N_7034);
nand U7746 (N_7746,N_7027,N_7329);
xor U7747 (N_7747,N_7454,N_7254);
nand U7748 (N_7748,N_7241,N_7023);
xnor U7749 (N_7749,N_7164,N_7013);
nor U7750 (N_7750,N_7123,N_7010);
or U7751 (N_7751,N_7112,N_7127);
and U7752 (N_7752,N_7330,N_7355);
or U7753 (N_7753,N_7311,N_7429);
nor U7754 (N_7754,N_7038,N_7114);
and U7755 (N_7755,N_7372,N_7386);
nor U7756 (N_7756,N_7169,N_7452);
xor U7757 (N_7757,N_7309,N_7263);
nand U7758 (N_7758,N_7299,N_7493);
or U7759 (N_7759,N_7000,N_7387);
or U7760 (N_7760,N_7315,N_7262);
nand U7761 (N_7761,N_7430,N_7494);
nand U7762 (N_7762,N_7293,N_7389);
nor U7763 (N_7763,N_7433,N_7217);
nand U7764 (N_7764,N_7176,N_7072);
xnor U7765 (N_7765,N_7275,N_7139);
and U7766 (N_7766,N_7441,N_7412);
and U7767 (N_7767,N_7432,N_7394);
xnor U7768 (N_7768,N_7191,N_7000);
and U7769 (N_7769,N_7168,N_7428);
or U7770 (N_7770,N_7471,N_7254);
nand U7771 (N_7771,N_7039,N_7449);
nor U7772 (N_7772,N_7410,N_7372);
or U7773 (N_7773,N_7006,N_7156);
and U7774 (N_7774,N_7088,N_7154);
nor U7775 (N_7775,N_7411,N_7270);
or U7776 (N_7776,N_7008,N_7168);
xor U7777 (N_7777,N_7176,N_7264);
nor U7778 (N_7778,N_7282,N_7350);
or U7779 (N_7779,N_7217,N_7416);
nand U7780 (N_7780,N_7478,N_7189);
xor U7781 (N_7781,N_7052,N_7076);
or U7782 (N_7782,N_7057,N_7012);
nand U7783 (N_7783,N_7205,N_7179);
xor U7784 (N_7784,N_7125,N_7311);
nor U7785 (N_7785,N_7424,N_7092);
nor U7786 (N_7786,N_7436,N_7209);
and U7787 (N_7787,N_7089,N_7282);
xnor U7788 (N_7788,N_7366,N_7468);
nand U7789 (N_7789,N_7418,N_7141);
or U7790 (N_7790,N_7153,N_7338);
nor U7791 (N_7791,N_7497,N_7387);
nor U7792 (N_7792,N_7110,N_7042);
or U7793 (N_7793,N_7320,N_7046);
nand U7794 (N_7794,N_7054,N_7287);
nand U7795 (N_7795,N_7077,N_7357);
nand U7796 (N_7796,N_7034,N_7307);
or U7797 (N_7797,N_7449,N_7401);
or U7798 (N_7798,N_7347,N_7314);
xor U7799 (N_7799,N_7475,N_7369);
nand U7800 (N_7800,N_7369,N_7436);
nor U7801 (N_7801,N_7423,N_7420);
nor U7802 (N_7802,N_7089,N_7151);
nor U7803 (N_7803,N_7237,N_7002);
nand U7804 (N_7804,N_7027,N_7178);
and U7805 (N_7805,N_7261,N_7184);
or U7806 (N_7806,N_7054,N_7444);
nor U7807 (N_7807,N_7325,N_7056);
or U7808 (N_7808,N_7234,N_7116);
nor U7809 (N_7809,N_7456,N_7423);
xor U7810 (N_7810,N_7234,N_7433);
and U7811 (N_7811,N_7491,N_7120);
or U7812 (N_7812,N_7475,N_7160);
nand U7813 (N_7813,N_7081,N_7250);
nor U7814 (N_7814,N_7440,N_7111);
and U7815 (N_7815,N_7107,N_7156);
nand U7816 (N_7816,N_7437,N_7218);
and U7817 (N_7817,N_7238,N_7102);
and U7818 (N_7818,N_7115,N_7070);
nor U7819 (N_7819,N_7178,N_7374);
or U7820 (N_7820,N_7054,N_7388);
xnor U7821 (N_7821,N_7214,N_7168);
or U7822 (N_7822,N_7207,N_7475);
nor U7823 (N_7823,N_7145,N_7023);
xnor U7824 (N_7824,N_7087,N_7352);
xnor U7825 (N_7825,N_7033,N_7411);
nor U7826 (N_7826,N_7164,N_7476);
nand U7827 (N_7827,N_7296,N_7250);
nand U7828 (N_7828,N_7358,N_7124);
and U7829 (N_7829,N_7160,N_7434);
nand U7830 (N_7830,N_7399,N_7183);
nor U7831 (N_7831,N_7011,N_7174);
nand U7832 (N_7832,N_7186,N_7031);
and U7833 (N_7833,N_7248,N_7308);
or U7834 (N_7834,N_7378,N_7418);
xor U7835 (N_7835,N_7028,N_7435);
or U7836 (N_7836,N_7192,N_7281);
nand U7837 (N_7837,N_7483,N_7290);
and U7838 (N_7838,N_7384,N_7176);
nand U7839 (N_7839,N_7329,N_7490);
and U7840 (N_7840,N_7241,N_7152);
and U7841 (N_7841,N_7170,N_7154);
nor U7842 (N_7842,N_7043,N_7171);
nor U7843 (N_7843,N_7156,N_7015);
xnor U7844 (N_7844,N_7304,N_7011);
nand U7845 (N_7845,N_7108,N_7065);
nor U7846 (N_7846,N_7047,N_7143);
xor U7847 (N_7847,N_7017,N_7221);
nor U7848 (N_7848,N_7463,N_7287);
or U7849 (N_7849,N_7019,N_7378);
nand U7850 (N_7850,N_7022,N_7132);
nor U7851 (N_7851,N_7275,N_7160);
and U7852 (N_7852,N_7033,N_7103);
and U7853 (N_7853,N_7469,N_7278);
nand U7854 (N_7854,N_7318,N_7182);
nor U7855 (N_7855,N_7364,N_7396);
xnor U7856 (N_7856,N_7096,N_7203);
or U7857 (N_7857,N_7368,N_7173);
nand U7858 (N_7858,N_7286,N_7016);
nor U7859 (N_7859,N_7318,N_7217);
xnor U7860 (N_7860,N_7127,N_7156);
and U7861 (N_7861,N_7437,N_7481);
xnor U7862 (N_7862,N_7426,N_7020);
or U7863 (N_7863,N_7321,N_7481);
xor U7864 (N_7864,N_7372,N_7264);
xnor U7865 (N_7865,N_7114,N_7039);
xor U7866 (N_7866,N_7300,N_7150);
xnor U7867 (N_7867,N_7102,N_7163);
and U7868 (N_7868,N_7132,N_7294);
xor U7869 (N_7869,N_7121,N_7261);
nor U7870 (N_7870,N_7433,N_7316);
nor U7871 (N_7871,N_7153,N_7052);
or U7872 (N_7872,N_7360,N_7341);
and U7873 (N_7873,N_7106,N_7097);
or U7874 (N_7874,N_7113,N_7294);
and U7875 (N_7875,N_7408,N_7357);
or U7876 (N_7876,N_7091,N_7250);
nor U7877 (N_7877,N_7341,N_7279);
nor U7878 (N_7878,N_7414,N_7241);
nand U7879 (N_7879,N_7165,N_7344);
and U7880 (N_7880,N_7153,N_7114);
and U7881 (N_7881,N_7332,N_7190);
nand U7882 (N_7882,N_7170,N_7131);
nor U7883 (N_7883,N_7263,N_7290);
nor U7884 (N_7884,N_7068,N_7101);
xnor U7885 (N_7885,N_7289,N_7215);
xor U7886 (N_7886,N_7256,N_7408);
nor U7887 (N_7887,N_7020,N_7135);
nor U7888 (N_7888,N_7201,N_7268);
nand U7889 (N_7889,N_7239,N_7350);
and U7890 (N_7890,N_7030,N_7109);
nand U7891 (N_7891,N_7064,N_7083);
or U7892 (N_7892,N_7076,N_7459);
nand U7893 (N_7893,N_7104,N_7342);
or U7894 (N_7894,N_7162,N_7419);
or U7895 (N_7895,N_7385,N_7135);
and U7896 (N_7896,N_7369,N_7438);
nor U7897 (N_7897,N_7475,N_7081);
nor U7898 (N_7898,N_7134,N_7217);
or U7899 (N_7899,N_7050,N_7125);
and U7900 (N_7900,N_7166,N_7230);
nor U7901 (N_7901,N_7420,N_7038);
nand U7902 (N_7902,N_7023,N_7328);
nor U7903 (N_7903,N_7161,N_7379);
xor U7904 (N_7904,N_7058,N_7369);
or U7905 (N_7905,N_7048,N_7471);
nand U7906 (N_7906,N_7035,N_7211);
and U7907 (N_7907,N_7221,N_7408);
and U7908 (N_7908,N_7279,N_7375);
xor U7909 (N_7909,N_7300,N_7155);
nand U7910 (N_7910,N_7411,N_7103);
nor U7911 (N_7911,N_7296,N_7294);
xor U7912 (N_7912,N_7212,N_7397);
nand U7913 (N_7913,N_7461,N_7484);
and U7914 (N_7914,N_7381,N_7369);
nand U7915 (N_7915,N_7496,N_7410);
nor U7916 (N_7916,N_7058,N_7171);
nor U7917 (N_7917,N_7020,N_7408);
xnor U7918 (N_7918,N_7181,N_7332);
xnor U7919 (N_7919,N_7003,N_7362);
and U7920 (N_7920,N_7219,N_7162);
and U7921 (N_7921,N_7362,N_7433);
nand U7922 (N_7922,N_7190,N_7175);
nand U7923 (N_7923,N_7287,N_7022);
nand U7924 (N_7924,N_7153,N_7204);
nand U7925 (N_7925,N_7385,N_7160);
and U7926 (N_7926,N_7151,N_7385);
nor U7927 (N_7927,N_7289,N_7377);
xor U7928 (N_7928,N_7368,N_7217);
xor U7929 (N_7929,N_7061,N_7248);
and U7930 (N_7930,N_7268,N_7147);
xor U7931 (N_7931,N_7036,N_7174);
or U7932 (N_7932,N_7113,N_7101);
nor U7933 (N_7933,N_7306,N_7401);
nor U7934 (N_7934,N_7499,N_7229);
or U7935 (N_7935,N_7161,N_7242);
nor U7936 (N_7936,N_7166,N_7228);
nand U7937 (N_7937,N_7465,N_7297);
nand U7938 (N_7938,N_7203,N_7386);
nor U7939 (N_7939,N_7477,N_7256);
nor U7940 (N_7940,N_7440,N_7308);
nor U7941 (N_7941,N_7475,N_7446);
nand U7942 (N_7942,N_7186,N_7025);
nand U7943 (N_7943,N_7180,N_7109);
xor U7944 (N_7944,N_7142,N_7342);
xor U7945 (N_7945,N_7498,N_7358);
nor U7946 (N_7946,N_7306,N_7121);
or U7947 (N_7947,N_7403,N_7389);
nand U7948 (N_7948,N_7121,N_7447);
or U7949 (N_7949,N_7136,N_7295);
nand U7950 (N_7950,N_7396,N_7464);
nand U7951 (N_7951,N_7030,N_7222);
and U7952 (N_7952,N_7178,N_7158);
nand U7953 (N_7953,N_7254,N_7462);
nand U7954 (N_7954,N_7490,N_7186);
or U7955 (N_7955,N_7276,N_7448);
xnor U7956 (N_7956,N_7022,N_7021);
nand U7957 (N_7957,N_7448,N_7284);
and U7958 (N_7958,N_7423,N_7498);
xnor U7959 (N_7959,N_7408,N_7272);
nand U7960 (N_7960,N_7130,N_7424);
nand U7961 (N_7961,N_7352,N_7127);
or U7962 (N_7962,N_7305,N_7483);
nand U7963 (N_7963,N_7363,N_7114);
xnor U7964 (N_7964,N_7240,N_7261);
or U7965 (N_7965,N_7484,N_7011);
xor U7966 (N_7966,N_7370,N_7484);
nand U7967 (N_7967,N_7298,N_7333);
nor U7968 (N_7968,N_7220,N_7055);
and U7969 (N_7969,N_7458,N_7387);
and U7970 (N_7970,N_7148,N_7361);
and U7971 (N_7971,N_7074,N_7292);
nand U7972 (N_7972,N_7112,N_7369);
xnor U7973 (N_7973,N_7404,N_7192);
or U7974 (N_7974,N_7028,N_7404);
or U7975 (N_7975,N_7419,N_7100);
xor U7976 (N_7976,N_7402,N_7258);
and U7977 (N_7977,N_7419,N_7342);
or U7978 (N_7978,N_7223,N_7401);
nor U7979 (N_7979,N_7423,N_7298);
nor U7980 (N_7980,N_7162,N_7156);
and U7981 (N_7981,N_7145,N_7112);
and U7982 (N_7982,N_7438,N_7234);
xor U7983 (N_7983,N_7372,N_7295);
or U7984 (N_7984,N_7257,N_7287);
nor U7985 (N_7985,N_7221,N_7377);
nor U7986 (N_7986,N_7169,N_7287);
or U7987 (N_7987,N_7431,N_7150);
xor U7988 (N_7988,N_7360,N_7058);
nor U7989 (N_7989,N_7413,N_7149);
or U7990 (N_7990,N_7042,N_7268);
and U7991 (N_7991,N_7305,N_7296);
nor U7992 (N_7992,N_7199,N_7069);
nor U7993 (N_7993,N_7197,N_7375);
and U7994 (N_7994,N_7245,N_7225);
and U7995 (N_7995,N_7263,N_7443);
nand U7996 (N_7996,N_7382,N_7184);
or U7997 (N_7997,N_7075,N_7428);
nand U7998 (N_7998,N_7255,N_7054);
or U7999 (N_7999,N_7139,N_7162);
and U8000 (N_8000,N_7765,N_7976);
nor U8001 (N_8001,N_7927,N_7956);
xor U8002 (N_8002,N_7974,N_7999);
nand U8003 (N_8003,N_7758,N_7872);
and U8004 (N_8004,N_7560,N_7740);
nor U8005 (N_8005,N_7670,N_7785);
and U8006 (N_8006,N_7697,N_7716);
or U8007 (N_8007,N_7641,N_7917);
nor U8008 (N_8008,N_7985,N_7726);
or U8009 (N_8009,N_7720,N_7732);
or U8010 (N_8010,N_7950,N_7781);
nand U8011 (N_8011,N_7606,N_7522);
nor U8012 (N_8012,N_7508,N_7757);
nand U8013 (N_8013,N_7937,N_7736);
and U8014 (N_8014,N_7793,N_7884);
nor U8015 (N_8015,N_7624,N_7938);
and U8016 (N_8016,N_7898,N_7578);
nor U8017 (N_8017,N_7590,N_7609);
nor U8018 (N_8018,N_7975,N_7667);
and U8019 (N_8019,N_7799,N_7602);
xnor U8020 (N_8020,N_7782,N_7656);
xnor U8021 (N_8021,N_7674,N_7870);
nand U8022 (N_8022,N_7551,N_7998);
nor U8023 (N_8023,N_7693,N_7748);
and U8024 (N_8024,N_7626,N_7696);
nand U8025 (N_8025,N_7700,N_7822);
or U8026 (N_8026,N_7874,N_7661);
xnor U8027 (N_8027,N_7814,N_7509);
nand U8028 (N_8028,N_7623,N_7721);
nor U8029 (N_8029,N_7811,N_7797);
nand U8030 (N_8030,N_7891,N_7901);
or U8031 (N_8031,N_7692,N_7866);
and U8032 (N_8032,N_7902,N_7651);
and U8033 (N_8033,N_7830,N_7896);
xor U8034 (N_8034,N_7663,N_7689);
nand U8035 (N_8035,N_7614,N_7800);
or U8036 (N_8036,N_7550,N_7655);
xor U8037 (N_8037,N_7643,N_7636);
nand U8038 (N_8038,N_7649,N_7681);
and U8039 (N_8039,N_7573,N_7934);
xnor U8040 (N_8040,N_7885,N_7657);
and U8041 (N_8041,N_7719,N_7798);
or U8042 (N_8042,N_7841,N_7569);
and U8043 (N_8043,N_7665,N_7741);
and U8044 (N_8044,N_7727,N_7744);
nand U8045 (N_8045,N_7947,N_7943);
xor U8046 (N_8046,N_7805,N_7980);
nand U8047 (N_8047,N_7981,N_7581);
nor U8048 (N_8048,N_7959,N_7737);
xnor U8049 (N_8049,N_7989,N_7876);
nand U8050 (N_8050,N_7671,N_7599);
or U8051 (N_8051,N_7982,N_7645);
nand U8052 (N_8052,N_7541,N_7604);
and U8053 (N_8053,N_7933,N_7973);
and U8054 (N_8054,N_7936,N_7565);
nand U8055 (N_8055,N_7756,N_7892);
and U8056 (N_8056,N_7586,N_7640);
xnor U8057 (N_8057,N_7549,N_7789);
nor U8058 (N_8058,N_7829,N_7894);
and U8059 (N_8059,N_7559,N_7762);
nor U8060 (N_8060,N_7734,N_7960);
or U8061 (N_8061,N_7619,N_7555);
xnor U8062 (N_8062,N_7575,N_7646);
and U8063 (N_8063,N_7596,N_7571);
xor U8064 (N_8064,N_7775,N_7728);
xnor U8065 (N_8065,N_7988,N_7576);
and U8066 (N_8066,N_7572,N_7502);
nand U8067 (N_8067,N_7598,N_7929);
and U8068 (N_8068,N_7941,N_7831);
xor U8069 (N_8069,N_7882,N_7704);
xor U8070 (N_8070,N_7924,N_7895);
nand U8071 (N_8071,N_7582,N_7911);
nand U8072 (N_8072,N_7944,N_7577);
nand U8073 (N_8073,N_7629,N_7566);
and U8074 (N_8074,N_7877,N_7846);
nand U8075 (N_8075,N_7890,N_7879);
xnor U8076 (N_8076,N_7539,N_7628);
xnor U8077 (N_8077,N_7834,N_7856);
or U8078 (N_8078,N_7538,N_7567);
and U8079 (N_8079,N_7766,N_7966);
xor U8080 (N_8080,N_7540,N_7729);
or U8081 (N_8081,N_7817,N_7820);
and U8082 (N_8082,N_7978,N_7842);
xor U8083 (N_8083,N_7777,N_7913);
xnor U8084 (N_8084,N_7827,N_7850);
xor U8085 (N_8085,N_7583,N_7678);
nand U8086 (N_8086,N_7632,N_7587);
xor U8087 (N_8087,N_7588,N_7712);
xor U8088 (N_8088,N_7530,N_7591);
xnor U8089 (N_8089,N_7650,N_7796);
nor U8090 (N_8090,N_7897,N_7613);
nor U8091 (N_8091,N_7949,N_7642);
and U8092 (N_8092,N_7711,N_7516);
nor U8093 (N_8093,N_7562,N_7622);
nor U8094 (N_8094,N_7763,N_7969);
and U8095 (N_8095,N_7634,N_7881);
nor U8096 (N_8096,N_7992,N_7521);
nor U8097 (N_8097,N_7772,N_7750);
xnor U8098 (N_8098,N_7925,N_7564);
nand U8099 (N_8099,N_7620,N_7844);
nor U8100 (N_8100,N_7605,N_7506);
or U8101 (N_8101,N_7914,N_7589);
and U8102 (N_8102,N_7597,N_7867);
nor U8103 (N_8103,N_7504,N_7840);
or U8104 (N_8104,N_7812,N_7547);
nand U8105 (N_8105,N_7824,N_7951);
xor U8106 (N_8106,N_7679,N_7783);
or U8107 (N_8107,N_7742,N_7548);
xor U8108 (N_8108,N_7616,N_7687);
or U8109 (N_8109,N_7922,N_7733);
and U8110 (N_8110,N_7828,N_7791);
nor U8111 (N_8111,N_7826,N_7935);
and U8112 (N_8112,N_7669,N_7536);
nor U8113 (N_8113,N_7995,N_7909);
xnor U8114 (N_8114,N_7544,N_7875);
nor U8115 (N_8115,N_7520,N_7735);
nor U8116 (N_8116,N_7568,N_7675);
nor U8117 (N_8117,N_7691,N_7792);
and U8118 (N_8118,N_7784,N_7786);
nor U8119 (N_8119,N_7754,N_7601);
or U8120 (N_8120,N_7861,N_7921);
nand U8121 (N_8121,N_7857,N_7862);
and U8122 (N_8122,N_7958,N_7585);
xor U8123 (N_8123,N_7847,N_7858);
nand U8124 (N_8124,N_7694,N_7563);
and U8125 (N_8125,N_7610,N_7625);
xor U8126 (N_8126,N_7557,N_7570);
and U8127 (N_8127,N_7698,N_7715);
or U8128 (N_8128,N_7769,N_7702);
or U8129 (N_8129,N_7939,N_7940);
and U8130 (N_8130,N_7725,N_7916);
nand U8131 (N_8131,N_7545,N_7684);
nand U8132 (N_8132,N_7534,N_7767);
or U8133 (N_8133,N_7863,N_7528);
and U8134 (N_8134,N_7703,N_7963);
or U8135 (N_8135,N_7873,N_7752);
xnor U8136 (N_8136,N_7953,N_7535);
nand U8137 (N_8137,N_7617,N_7804);
and U8138 (N_8138,N_7864,N_7659);
and U8139 (N_8139,N_7851,N_7647);
xor U8140 (N_8140,N_7832,N_7531);
nand U8141 (N_8141,N_7753,N_7823);
or U8142 (N_8142,N_7816,N_7964);
nand U8143 (N_8143,N_7957,N_7580);
or U8144 (N_8144,N_7631,N_7554);
nor U8145 (N_8145,N_7903,N_7945);
and U8146 (N_8146,N_7600,N_7971);
xor U8147 (N_8147,N_7615,N_7654);
and U8148 (N_8148,N_7630,N_7759);
nor U8149 (N_8149,N_7690,N_7524);
or U8150 (N_8150,N_7854,N_7918);
xnor U8151 (N_8151,N_7833,N_7910);
nor U8152 (N_8152,N_7997,N_7806);
or U8153 (N_8153,N_7664,N_7923);
and U8154 (N_8154,N_7543,N_7984);
xnor U8155 (N_8155,N_7653,N_7778);
nor U8156 (N_8156,N_7836,N_7749);
or U8157 (N_8157,N_7714,N_7970);
and U8158 (N_8158,N_7608,N_7505);
or U8159 (N_8159,N_7707,N_7595);
nand U8160 (N_8160,N_7658,N_7787);
nand U8161 (N_8161,N_7865,N_7648);
xor U8162 (N_8162,N_7673,N_7774);
nand U8163 (N_8163,N_7611,N_7776);
nor U8164 (N_8164,N_7503,N_7660);
nand U8165 (N_8165,N_7760,N_7993);
xnor U8166 (N_8166,N_7771,N_7739);
or U8167 (N_8167,N_7819,N_7542);
xnor U8168 (N_8168,N_7848,N_7986);
or U8169 (N_8169,N_7904,N_7633);
nand U8170 (N_8170,N_7802,N_7529);
nor U8171 (N_8171,N_7790,N_7637);
xor U8172 (N_8172,N_7525,N_7869);
or U8173 (N_8173,N_7893,N_7676);
and U8174 (N_8174,N_7526,N_7501);
nor U8175 (N_8175,N_7906,N_7512);
nor U8176 (N_8176,N_7556,N_7558);
xor U8177 (N_8177,N_7932,N_7794);
nor U8178 (N_8178,N_7627,N_7618);
nor U8179 (N_8179,N_7731,N_7886);
and U8180 (N_8180,N_7513,N_7713);
nor U8181 (N_8181,N_7788,N_7983);
nand U8182 (N_8182,N_7518,N_7768);
nand U8183 (N_8183,N_7685,N_7803);
or U8184 (N_8184,N_7859,N_7967);
or U8185 (N_8185,N_7709,N_7579);
or U8186 (N_8186,N_7519,N_7880);
nand U8187 (N_8187,N_7818,N_7584);
nand U8188 (N_8188,N_7546,N_7722);
or U8189 (N_8189,N_7919,N_7990);
nand U8190 (N_8190,N_7889,N_7695);
xor U8191 (N_8191,N_7868,N_7593);
or U8192 (N_8192,N_7574,N_7773);
nor U8193 (N_8193,N_7533,N_7718);
xnor U8194 (N_8194,N_7607,N_7845);
nor U8195 (N_8195,N_7523,N_7668);
and U8196 (N_8196,N_7537,N_7652);
and U8197 (N_8197,N_7905,N_7835);
xor U8198 (N_8198,N_7977,N_7710);
nand U8199 (N_8199,N_7883,N_7514);
xor U8200 (N_8200,N_7592,N_7991);
and U8201 (N_8201,N_7942,N_7837);
nor U8202 (N_8202,N_7515,N_7532);
and U8203 (N_8203,N_7717,N_7764);
or U8204 (N_8204,N_7552,N_7644);
nand U8205 (N_8205,N_7915,N_7746);
or U8206 (N_8206,N_7666,N_7871);
xor U8207 (N_8207,N_7809,N_7930);
or U8208 (N_8208,N_7594,N_7510);
nor U8209 (N_8209,N_7808,N_7843);
or U8210 (N_8210,N_7855,N_7751);
or U8211 (N_8211,N_7928,N_7724);
and U8212 (N_8212,N_7852,N_7810);
xor U8213 (N_8213,N_7979,N_7888);
or U8214 (N_8214,N_7807,N_7994);
nor U8215 (N_8215,N_7839,N_7621);
nor U8216 (N_8216,N_7920,N_7706);
or U8217 (N_8217,N_7948,N_7511);
nand U8218 (N_8218,N_7779,N_7965);
nand U8219 (N_8219,N_7638,N_7500);
nor U8220 (N_8220,N_7815,N_7853);
and U8221 (N_8221,N_7747,N_7931);
nor U8222 (N_8222,N_7961,N_7908);
nor U8223 (N_8223,N_7683,N_7738);
and U8224 (N_8224,N_7705,N_7561);
nand U8225 (N_8225,N_7677,N_7780);
or U8226 (N_8226,N_7907,N_7795);
nor U8227 (N_8227,N_7761,N_7686);
nand U8228 (N_8228,N_7672,N_7743);
and U8229 (N_8229,N_7962,N_7887);
and U8230 (N_8230,N_7955,N_7825);
or U8231 (N_8231,N_7755,N_7987);
and U8232 (N_8232,N_7912,N_7723);
xnor U8233 (N_8233,N_7662,N_7701);
nor U8234 (N_8234,N_7745,N_7801);
and U8235 (N_8235,N_7770,N_7900);
or U8236 (N_8236,N_7708,N_7813);
nor U8237 (N_8237,N_7682,N_7639);
nor U8238 (N_8238,N_7849,N_7730);
nor U8239 (N_8239,N_7899,N_7527);
nor U8240 (N_8240,N_7972,N_7954);
and U8241 (N_8241,N_7926,N_7603);
nor U8242 (N_8242,N_7860,N_7635);
or U8243 (N_8243,N_7517,N_7821);
or U8244 (N_8244,N_7553,N_7507);
and U8245 (N_8245,N_7699,N_7838);
nor U8246 (N_8246,N_7946,N_7952);
and U8247 (N_8247,N_7680,N_7878);
or U8248 (N_8248,N_7968,N_7996);
nand U8249 (N_8249,N_7688,N_7612);
nor U8250 (N_8250,N_7760,N_7697);
nor U8251 (N_8251,N_7615,N_7501);
xor U8252 (N_8252,N_7535,N_7809);
or U8253 (N_8253,N_7825,N_7806);
nand U8254 (N_8254,N_7810,N_7617);
or U8255 (N_8255,N_7715,N_7895);
xnor U8256 (N_8256,N_7948,N_7566);
nor U8257 (N_8257,N_7929,N_7607);
nor U8258 (N_8258,N_7933,N_7597);
nor U8259 (N_8259,N_7674,N_7562);
nor U8260 (N_8260,N_7533,N_7678);
nand U8261 (N_8261,N_7775,N_7689);
and U8262 (N_8262,N_7569,N_7718);
xnor U8263 (N_8263,N_7736,N_7612);
nand U8264 (N_8264,N_7575,N_7818);
or U8265 (N_8265,N_7585,N_7952);
nor U8266 (N_8266,N_7969,N_7844);
or U8267 (N_8267,N_7604,N_7924);
or U8268 (N_8268,N_7709,N_7672);
nand U8269 (N_8269,N_7814,N_7739);
nor U8270 (N_8270,N_7699,N_7915);
or U8271 (N_8271,N_7811,N_7637);
nand U8272 (N_8272,N_7617,N_7548);
nor U8273 (N_8273,N_7907,N_7656);
and U8274 (N_8274,N_7622,N_7768);
nand U8275 (N_8275,N_7959,N_7661);
xor U8276 (N_8276,N_7514,N_7691);
nand U8277 (N_8277,N_7780,N_7638);
nor U8278 (N_8278,N_7883,N_7622);
or U8279 (N_8279,N_7565,N_7515);
xor U8280 (N_8280,N_7587,N_7685);
and U8281 (N_8281,N_7920,N_7664);
and U8282 (N_8282,N_7725,N_7547);
nand U8283 (N_8283,N_7752,N_7687);
or U8284 (N_8284,N_7640,N_7712);
or U8285 (N_8285,N_7803,N_7835);
and U8286 (N_8286,N_7567,N_7955);
nand U8287 (N_8287,N_7575,N_7712);
nand U8288 (N_8288,N_7669,N_7664);
nand U8289 (N_8289,N_7683,N_7771);
nand U8290 (N_8290,N_7716,N_7508);
xnor U8291 (N_8291,N_7645,N_7790);
nor U8292 (N_8292,N_7724,N_7886);
xor U8293 (N_8293,N_7944,N_7550);
xnor U8294 (N_8294,N_7887,N_7615);
xnor U8295 (N_8295,N_7544,N_7746);
and U8296 (N_8296,N_7610,N_7803);
xnor U8297 (N_8297,N_7595,N_7580);
xnor U8298 (N_8298,N_7776,N_7684);
nand U8299 (N_8299,N_7586,N_7597);
and U8300 (N_8300,N_7834,N_7631);
and U8301 (N_8301,N_7644,N_7787);
and U8302 (N_8302,N_7787,N_7669);
xnor U8303 (N_8303,N_7971,N_7827);
xnor U8304 (N_8304,N_7753,N_7889);
nor U8305 (N_8305,N_7611,N_7604);
or U8306 (N_8306,N_7949,N_7643);
xnor U8307 (N_8307,N_7957,N_7746);
xor U8308 (N_8308,N_7629,N_7529);
or U8309 (N_8309,N_7542,N_7982);
xnor U8310 (N_8310,N_7937,N_7548);
and U8311 (N_8311,N_7750,N_7812);
or U8312 (N_8312,N_7600,N_7979);
or U8313 (N_8313,N_7809,N_7996);
xnor U8314 (N_8314,N_7522,N_7740);
and U8315 (N_8315,N_7677,N_7771);
and U8316 (N_8316,N_7954,N_7945);
xor U8317 (N_8317,N_7727,N_7902);
and U8318 (N_8318,N_7908,N_7708);
or U8319 (N_8319,N_7910,N_7615);
and U8320 (N_8320,N_7643,N_7638);
nand U8321 (N_8321,N_7504,N_7857);
or U8322 (N_8322,N_7671,N_7998);
and U8323 (N_8323,N_7645,N_7654);
nor U8324 (N_8324,N_7833,N_7884);
nor U8325 (N_8325,N_7668,N_7616);
xnor U8326 (N_8326,N_7849,N_7760);
or U8327 (N_8327,N_7938,N_7967);
nand U8328 (N_8328,N_7785,N_7721);
xnor U8329 (N_8329,N_7744,N_7578);
and U8330 (N_8330,N_7584,N_7516);
nand U8331 (N_8331,N_7518,N_7967);
nand U8332 (N_8332,N_7527,N_7548);
xnor U8333 (N_8333,N_7877,N_7516);
nand U8334 (N_8334,N_7752,N_7615);
xnor U8335 (N_8335,N_7622,N_7919);
nor U8336 (N_8336,N_7764,N_7989);
and U8337 (N_8337,N_7546,N_7591);
xnor U8338 (N_8338,N_7854,N_7693);
nand U8339 (N_8339,N_7841,N_7614);
nand U8340 (N_8340,N_7613,N_7880);
or U8341 (N_8341,N_7939,N_7938);
or U8342 (N_8342,N_7645,N_7747);
nor U8343 (N_8343,N_7546,N_7723);
nor U8344 (N_8344,N_7823,N_7790);
and U8345 (N_8345,N_7719,N_7989);
nor U8346 (N_8346,N_7526,N_7683);
and U8347 (N_8347,N_7931,N_7934);
and U8348 (N_8348,N_7582,N_7875);
or U8349 (N_8349,N_7899,N_7575);
nor U8350 (N_8350,N_7817,N_7617);
nor U8351 (N_8351,N_7880,N_7909);
or U8352 (N_8352,N_7655,N_7769);
nand U8353 (N_8353,N_7910,N_7939);
xor U8354 (N_8354,N_7551,N_7580);
and U8355 (N_8355,N_7940,N_7749);
nor U8356 (N_8356,N_7609,N_7857);
or U8357 (N_8357,N_7953,N_7793);
nor U8358 (N_8358,N_7874,N_7662);
xnor U8359 (N_8359,N_7735,N_7610);
and U8360 (N_8360,N_7597,N_7842);
or U8361 (N_8361,N_7847,N_7810);
or U8362 (N_8362,N_7771,N_7642);
or U8363 (N_8363,N_7569,N_7595);
nand U8364 (N_8364,N_7794,N_7567);
nand U8365 (N_8365,N_7773,N_7638);
and U8366 (N_8366,N_7678,N_7654);
nor U8367 (N_8367,N_7956,N_7920);
or U8368 (N_8368,N_7597,N_7997);
or U8369 (N_8369,N_7828,N_7556);
or U8370 (N_8370,N_7753,N_7893);
or U8371 (N_8371,N_7896,N_7514);
nand U8372 (N_8372,N_7573,N_7815);
nand U8373 (N_8373,N_7814,N_7775);
xor U8374 (N_8374,N_7894,N_7850);
or U8375 (N_8375,N_7798,N_7735);
xnor U8376 (N_8376,N_7726,N_7986);
nand U8377 (N_8377,N_7804,N_7667);
and U8378 (N_8378,N_7543,N_7918);
nand U8379 (N_8379,N_7675,N_7572);
nand U8380 (N_8380,N_7817,N_7894);
xor U8381 (N_8381,N_7689,N_7537);
and U8382 (N_8382,N_7799,N_7701);
xnor U8383 (N_8383,N_7953,N_7760);
or U8384 (N_8384,N_7737,N_7597);
and U8385 (N_8385,N_7599,N_7902);
nor U8386 (N_8386,N_7715,N_7943);
xor U8387 (N_8387,N_7698,N_7602);
and U8388 (N_8388,N_7902,N_7628);
and U8389 (N_8389,N_7577,N_7795);
xor U8390 (N_8390,N_7816,N_7508);
xnor U8391 (N_8391,N_7792,N_7916);
xor U8392 (N_8392,N_7974,N_7551);
nand U8393 (N_8393,N_7820,N_7844);
xnor U8394 (N_8394,N_7905,N_7633);
xnor U8395 (N_8395,N_7926,N_7660);
xor U8396 (N_8396,N_7709,N_7606);
nand U8397 (N_8397,N_7697,N_7528);
nor U8398 (N_8398,N_7867,N_7607);
and U8399 (N_8399,N_7707,N_7887);
and U8400 (N_8400,N_7847,N_7609);
and U8401 (N_8401,N_7963,N_7590);
xnor U8402 (N_8402,N_7653,N_7926);
or U8403 (N_8403,N_7865,N_7937);
nand U8404 (N_8404,N_7537,N_7990);
xor U8405 (N_8405,N_7901,N_7641);
nor U8406 (N_8406,N_7947,N_7522);
nand U8407 (N_8407,N_7924,N_7540);
and U8408 (N_8408,N_7704,N_7684);
and U8409 (N_8409,N_7996,N_7931);
and U8410 (N_8410,N_7874,N_7785);
xnor U8411 (N_8411,N_7563,N_7796);
nand U8412 (N_8412,N_7820,N_7843);
xnor U8413 (N_8413,N_7759,N_7609);
xor U8414 (N_8414,N_7630,N_7879);
or U8415 (N_8415,N_7631,N_7921);
xnor U8416 (N_8416,N_7730,N_7740);
xor U8417 (N_8417,N_7717,N_7909);
nor U8418 (N_8418,N_7846,N_7816);
nand U8419 (N_8419,N_7689,N_7675);
nor U8420 (N_8420,N_7877,N_7628);
xnor U8421 (N_8421,N_7909,N_7746);
and U8422 (N_8422,N_7864,N_7716);
nor U8423 (N_8423,N_7752,N_7682);
nand U8424 (N_8424,N_7550,N_7688);
nand U8425 (N_8425,N_7933,N_7779);
nor U8426 (N_8426,N_7891,N_7992);
nand U8427 (N_8427,N_7543,N_7930);
nand U8428 (N_8428,N_7517,N_7809);
and U8429 (N_8429,N_7631,N_7980);
xor U8430 (N_8430,N_7790,N_7981);
and U8431 (N_8431,N_7913,N_7680);
or U8432 (N_8432,N_7500,N_7795);
or U8433 (N_8433,N_7742,N_7561);
nand U8434 (N_8434,N_7625,N_7571);
xor U8435 (N_8435,N_7636,N_7524);
nor U8436 (N_8436,N_7806,N_7949);
nand U8437 (N_8437,N_7916,N_7634);
nor U8438 (N_8438,N_7882,N_7820);
or U8439 (N_8439,N_7820,N_7578);
and U8440 (N_8440,N_7609,N_7741);
or U8441 (N_8441,N_7668,N_7507);
nand U8442 (N_8442,N_7825,N_7842);
xor U8443 (N_8443,N_7787,N_7963);
and U8444 (N_8444,N_7871,N_7866);
nand U8445 (N_8445,N_7638,N_7775);
and U8446 (N_8446,N_7939,N_7969);
nand U8447 (N_8447,N_7632,N_7919);
or U8448 (N_8448,N_7514,N_7853);
nor U8449 (N_8449,N_7831,N_7874);
nor U8450 (N_8450,N_7846,N_7720);
nor U8451 (N_8451,N_7835,N_7977);
xnor U8452 (N_8452,N_7563,N_7526);
nand U8453 (N_8453,N_7526,N_7610);
nand U8454 (N_8454,N_7957,N_7766);
nand U8455 (N_8455,N_7744,N_7673);
nand U8456 (N_8456,N_7909,N_7599);
xor U8457 (N_8457,N_7680,N_7844);
or U8458 (N_8458,N_7706,N_7572);
nor U8459 (N_8459,N_7779,N_7936);
nor U8460 (N_8460,N_7919,N_7991);
nand U8461 (N_8461,N_7725,N_7947);
or U8462 (N_8462,N_7831,N_7889);
nand U8463 (N_8463,N_7546,N_7635);
or U8464 (N_8464,N_7621,N_7954);
and U8465 (N_8465,N_7700,N_7772);
and U8466 (N_8466,N_7577,N_7836);
nor U8467 (N_8467,N_7601,N_7569);
nand U8468 (N_8468,N_7975,N_7618);
nand U8469 (N_8469,N_7836,N_7984);
nand U8470 (N_8470,N_7804,N_7607);
xor U8471 (N_8471,N_7720,N_7938);
or U8472 (N_8472,N_7840,N_7647);
nor U8473 (N_8473,N_7502,N_7862);
and U8474 (N_8474,N_7723,N_7929);
and U8475 (N_8475,N_7660,N_7580);
and U8476 (N_8476,N_7729,N_7925);
nand U8477 (N_8477,N_7659,N_7529);
xor U8478 (N_8478,N_7612,N_7724);
or U8479 (N_8479,N_7906,N_7661);
xor U8480 (N_8480,N_7546,N_7610);
or U8481 (N_8481,N_7711,N_7895);
nor U8482 (N_8482,N_7714,N_7533);
nor U8483 (N_8483,N_7993,N_7509);
or U8484 (N_8484,N_7807,N_7648);
and U8485 (N_8485,N_7517,N_7689);
nor U8486 (N_8486,N_7576,N_7676);
nor U8487 (N_8487,N_7916,N_7561);
nor U8488 (N_8488,N_7551,N_7814);
xor U8489 (N_8489,N_7554,N_7790);
or U8490 (N_8490,N_7538,N_7872);
and U8491 (N_8491,N_7579,N_7984);
nand U8492 (N_8492,N_7817,N_7997);
or U8493 (N_8493,N_7959,N_7876);
nor U8494 (N_8494,N_7832,N_7799);
and U8495 (N_8495,N_7585,N_7647);
nor U8496 (N_8496,N_7812,N_7965);
xor U8497 (N_8497,N_7811,N_7740);
xnor U8498 (N_8498,N_7627,N_7754);
and U8499 (N_8499,N_7604,N_7608);
xor U8500 (N_8500,N_8424,N_8417);
xnor U8501 (N_8501,N_8070,N_8157);
xnor U8502 (N_8502,N_8214,N_8174);
xnor U8503 (N_8503,N_8172,N_8378);
and U8504 (N_8504,N_8373,N_8176);
xor U8505 (N_8505,N_8251,N_8147);
and U8506 (N_8506,N_8493,N_8319);
and U8507 (N_8507,N_8278,N_8126);
and U8508 (N_8508,N_8369,N_8485);
nor U8509 (N_8509,N_8186,N_8374);
nand U8510 (N_8510,N_8124,N_8464);
or U8511 (N_8511,N_8137,N_8117);
nor U8512 (N_8512,N_8177,N_8104);
nor U8513 (N_8513,N_8330,N_8032);
nand U8514 (N_8514,N_8436,N_8021);
and U8515 (N_8515,N_8262,N_8487);
nor U8516 (N_8516,N_8290,N_8307);
or U8517 (N_8517,N_8063,N_8213);
xnor U8518 (N_8518,N_8030,N_8057);
and U8519 (N_8519,N_8444,N_8257);
xnor U8520 (N_8520,N_8324,N_8086);
xor U8521 (N_8521,N_8170,N_8250);
xnor U8522 (N_8522,N_8017,N_8089);
nor U8523 (N_8523,N_8038,N_8005);
or U8524 (N_8524,N_8349,N_8446);
or U8525 (N_8525,N_8354,N_8162);
nor U8526 (N_8526,N_8370,N_8434);
and U8527 (N_8527,N_8394,N_8052);
and U8528 (N_8528,N_8123,N_8026);
or U8529 (N_8529,N_8239,N_8060);
xor U8530 (N_8530,N_8050,N_8187);
nor U8531 (N_8531,N_8197,N_8087);
and U8532 (N_8532,N_8247,N_8184);
or U8533 (N_8533,N_8221,N_8199);
or U8534 (N_8534,N_8220,N_8058);
and U8535 (N_8535,N_8275,N_8405);
nor U8536 (N_8536,N_8027,N_8399);
nor U8537 (N_8537,N_8460,N_8108);
nor U8538 (N_8538,N_8410,N_8136);
nor U8539 (N_8539,N_8031,N_8191);
or U8540 (N_8540,N_8361,N_8272);
and U8541 (N_8541,N_8388,N_8094);
nand U8542 (N_8542,N_8376,N_8291);
xor U8543 (N_8543,N_8222,N_8238);
or U8544 (N_8544,N_8085,N_8280);
nor U8545 (N_8545,N_8461,N_8249);
xnor U8546 (N_8546,N_8044,N_8396);
and U8547 (N_8547,N_8178,N_8273);
xor U8548 (N_8548,N_8152,N_8336);
and U8549 (N_8549,N_8003,N_8457);
nor U8550 (N_8550,N_8043,N_8167);
nor U8551 (N_8551,N_8179,N_8345);
nand U8552 (N_8552,N_8252,N_8059);
nor U8553 (N_8553,N_8308,N_8053);
nor U8554 (N_8554,N_8259,N_8200);
xnor U8555 (N_8555,N_8289,N_8175);
nor U8556 (N_8556,N_8074,N_8453);
nor U8557 (N_8557,N_8007,N_8045);
nand U8558 (N_8558,N_8425,N_8389);
nor U8559 (N_8559,N_8452,N_8386);
nand U8560 (N_8560,N_8268,N_8287);
and U8561 (N_8561,N_8328,N_8406);
nor U8562 (N_8562,N_8042,N_8049);
or U8563 (N_8563,N_8107,N_8150);
and U8564 (N_8564,N_8196,N_8382);
and U8565 (N_8565,N_8366,N_8264);
nand U8566 (N_8566,N_8450,N_8277);
or U8567 (N_8567,N_8232,N_8304);
or U8568 (N_8568,N_8348,N_8484);
nand U8569 (N_8569,N_8056,N_8227);
or U8570 (N_8570,N_8471,N_8201);
or U8571 (N_8571,N_8371,N_8010);
or U8572 (N_8572,N_8437,N_8482);
or U8573 (N_8573,N_8113,N_8169);
nor U8574 (N_8574,N_8244,N_8332);
nand U8575 (N_8575,N_8022,N_8492);
nor U8576 (N_8576,N_8076,N_8047);
nor U8577 (N_8577,N_8171,N_8109);
xnor U8578 (N_8578,N_8216,N_8497);
nand U8579 (N_8579,N_8310,N_8215);
xnor U8580 (N_8580,N_8431,N_8456);
xor U8581 (N_8581,N_8339,N_8205);
nor U8582 (N_8582,N_8365,N_8305);
nor U8583 (N_8583,N_8148,N_8419);
or U8584 (N_8584,N_8357,N_8329);
xnor U8585 (N_8585,N_8080,N_8004);
nand U8586 (N_8586,N_8393,N_8037);
nand U8587 (N_8587,N_8292,N_8132);
nor U8588 (N_8588,N_8208,N_8270);
and U8589 (N_8589,N_8081,N_8019);
nand U8590 (N_8590,N_8013,N_8018);
or U8591 (N_8591,N_8055,N_8480);
xnor U8592 (N_8592,N_8188,N_8009);
xnor U8593 (N_8593,N_8276,N_8253);
nor U8594 (N_8594,N_8006,N_8435);
or U8595 (N_8595,N_8286,N_8432);
nand U8596 (N_8596,N_8494,N_8102);
xnor U8597 (N_8597,N_8149,N_8182);
nor U8598 (N_8598,N_8467,N_8428);
nor U8599 (N_8599,N_8195,N_8284);
nor U8600 (N_8600,N_8491,N_8210);
and U8601 (N_8601,N_8343,N_8161);
nor U8602 (N_8602,N_8311,N_8235);
xor U8603 (N_8603,N_8071,N_8130);
nand U8604 (N_8604,N_8029,N_8067);
or U8605 (N_8605,N_8254,N_8098);
nand U8606 (N_8606,N_8039,N_8267);
and U8607 (N_8607,N_8449,N_8285);
nand U8608 (N_8608,N_8119,N_8458);
nand U8609 (N_8609,N_8226,N_8346);
and U8610 (N_8610,N_8245,N_8411);
and U8611 (N_8611,N_8398,N_8111);
nand U8612 (N_8612,N_8092,N_8218);
and U8613 (N_8613,N_8317,N_8112);
or U8614 (N_8614,N_8133,N_8023);
and U8615 (N_8615,N_8282,N_8293);
xnor U8616 (N_8616,N_8443,N_8095);
or U8617 (N_8617,N_8001,N_8447);
nor U8618 (N_8618,N_8041,N_8016);
nor U8619 (N_8619,N_8015,N_8478);
and U8620 (N_8620,N_8141,N_8046);
nor U8621 (N_8621,N_8151,N_8440);
nor U8622 (N_8622,N_8402,N_8299);
xnor U8623 (N_8623,N_8156,N_8288);
nor U8624 (N_8624,N_8331,N_8142);
nor U8625 (N_8625,N_8298,N_8066);
and U8626 (N_8626,N_8413,N_8139);
nand U8627 (N_8627,N_8420,N_8103);
xnor U8628 (N_8628,N_8093,N_8229);
or U8629 (N_8629,N_8283,N_8498);
or U8630 (N_8630,N_8483,N_8140);
nand U8631 (N_8631,N_8163,N_8256);
or U8632 (N_8632,N_8155,N_8145);
nor U8633 (N_8633,N_8391,N_8203);
nand U8634 (N_8634,N_8068,N_8490);
and U8635 (N_8635,N_8474,N_8240);
and U8636 (N_8636,N_8372,N_8320);
nor U8637 (N_8637,N_8159,N_8091);
nor U8638 (N_8638,N_8212,N_8422);
nand U8639 (N_8639,N_8326,N_8408);
nand U8640 (N_8640,N_8033,N_8204);
or U8641 (N_8641,N_8316,N_8473);
nor U8642 (N_8642,N_8225,N_8384);
or U8643 (N_8643,N_8274,N_8279);
nor U8644 (N_8644,N_8427,N_8481);
and U8645 (N_8645,N_8000,N_8297);
nand U8646 (N_8646,N_8451,N_8322);
nand U8647 (N_8647,N_8164,N_8448);
nand U8648 (N_8648,N_8301,N_8407);
nand U8649 (N_8649,N_8358,N_8194);
and U8650 (N_8650,N_8255,N_8360);
nor U8651 (N_8651,N_8122,N_8106);
xnor U8652 (N_8652,N_8241,N_8048);
and U8653 (N_8653,N_8024,N_8488);
nor U8654 (N_8654,N_8198,N_8146);
or U8655 (N_8655,N_8219,N_8154);
xnor U8656 (N_8656,N_8295,N_8134);
nand U8657 (N_8657,N_8116,N_8064);
nor U8658 (N_8658,N_8160,N_8313);
and U8659 (N_8659,N_8395,N_8377);
nand U8660 (N_8660,N_8090,N_8468);
or U8661 (N_8661,N_8495,N_8125);
and U8662 (N_8662,N_8496,N_8028);
nor U8663 (N_8663,N_8403,N_8309);
nor U8664 (N_8664,N_8392,N_8025);
nor U8665 (N_8665,N_8323,N_8318);
nand U8666 (N_8666,N_8069,N_8340);
xor U8667 (N_8667,N_8368,N_8306);
xor U8668 (N_8668,N_8414,N_8034);
nand U8669 (N_8669,N_8135,N_8353);
nor U8670 (N_8670,N_8228,N_8248);
or U8671 (N_8671,N_8065,N_8101);
xnor U8672 (N_8672,N_8165,N_8083);
xnor U8673 (N_8673,N_8051,N_8131);
or U8674 (N_8674,N_8499,N_8477);
nor U8675 (N_8675,N_8231,N_8265);
nor U8676 (N_8676,N_8062,N_8404);
nor U8677 (N_8677,N_8439,N_8181);
or U8678 (N_8678,N_8421,N_8243);
nand U8679 (N_8679,N_8183,N_8223);
nor U8680 (N_8680,N_8294,N_8475);
nor U8681 (N_8681,N_8476,N_8350);
or U8682 (N_8682,N_8397,N_8012);
nor U8683 (N_8683,N_8347,N_8035);
xor U8684 (N_8684,N_8099,N_8296);
and U8685 (N_8685,N_8230,N_8158);
nor U8686 (N_8686,N_8362,N_8206);
or U8687 (N_8687,N_8462,N_8430);
and U8688 (N_8688,N_8415,N_8115);
nor U8689 (N_8689,N_8364,N_8084);
or U8690 (N_8690,N_8072,N_8466);
xor U8691 (N_8691,N_8390,N_8400);
and U8692 (N_8692,N_8401,N_8077);
nor U8693 (N_8693,N_8281,N_8011);
nand U8694 (N_8694,N_8110,N_8173);
nor U8695 (N_8695,N_8338,N_8105);
nand U8696 (N_8696,N_8100,N_8202);
and U8697 (N_8697,N_8379,N_8168);
nand U8698 (N_8698,N_8237,N_8075);
or U8699 (N_8699,N_8079,N_8192);
nand U8700 (N_8700,N_8314,N_8020);
nand U8701 (N_8701,N_8344,N_8143);
and U8702 (N_8702,N_8078,N_8337);
nor U8703 (N_8703,N_8454,N_8416);
nor U8704 (N_8704,N_8128,N_8097);
nor U8705 (N_8705,N_8441,N_8412);
and U8706 (N_8706,N_8138,N_8375);
xnor U8707 (N_8707,N_8014,N_8341);
xnor U8708 (N_8708,N_8207,N_8233);
or U8709 (N_8709,N_8383,N_8185);
xnor U8710 (N_8710,N_8302,N_8234);
or U8711 (N_8711,N_8470,N_8271);
nor U8712 (N_8712,N_8385,N_8263);
xnor U8713 (N_8713,N_8260,N_8442);
and U8714 (N_8714,N_8335,N_8486);
nor U8715 (N_8715,N_8190,N_8355);
xnor U8716 (N_8716,N_8088,N_8333);
nor U8717 (N_8717,N_8129,N_8166);
nor U8718 (N_8718,N_8315,N_8356);
or U8719 (N_8719,N_8367,N_8433);
nand U8720 (N_8720,N_8459,N_8445);
nor U8721 (N_8721,N_8351,N_8321);
xnor U8722 (N_8722,N_8472,N_8096);
nor U8723 (N_8723,N_8455,N_8325);
or U8724 (N_8724,N_8269,N_8438);
or U8725 (N_8725,N_8144,N_8418);
or U8726 (N_8726,N_8479,N_8342);
xnor U8727 (N_8727,N_8327,N_8380);
and U8728 (N_8728,N_8312,N_8469);
xnor U8729 (N_8729,N_8258,N_8303);
or U8730 (N_8730,N_8002,N_8381);
nand U8731 (N_8731,N_8352,N_8387);
nand U8732 (N_8732,N_8465,N_8429);
xor U8733 (N_8733,N_8236,N_8363);
nor U8734 (N_8734,N_8463,N_8121);
or U8735 (N_8735,N_8118,N_8266);
or U8736 (N_8736,N_8040,N_8334);
xor U8737 (N_8737,N_8114,N_8224);
nor U8738 (N_8738,N_8242,N_8082);
or U8739 (N_8739,N_8246,N_8409);
and U8740 (N_8740,N_8261,N_8359);
and U8741 (N_8741,N_8054,N_8423);
nand U8742 (N_8742,N_8127,N_8209);
nor U8743 (N_8743,N_8036,N_8153);
nor U8744 (N_8744,N_8189,N_8193);
or U8745 (N_8745,N_8217,N_8300);
xnor U8746 (N_8746,N_8211,N_8061);
nand U8747 (N_8747,N_8073,N_8180);
and U8748 (N_8748,N_8489,N_8426);
and U8749 (N_8749,N_8120,N_8008);
or U8750 (N_8750,N_8016,N_8389);
nand U8751 (N_8751,N_8263,N_8308);
and U8752 (N_8752,N_8391,N_8327);
xnor U8753 (N_8753,N_8468,N_8412);
and U8754 (N_8754,N_8230,N_8210);
and U8755 (N_8755,N_8150,N_8067);
or U8756 (N_8756,N_8424,N_8214);
nand U8757 (N_8757,N_8409,N_8330);
or U8758 (N_8758,N_8191,N_8060);
xnor U8759 (N_8759,N_8018,N_8352);
and U8760 (N_8760,N_8194,N_8389);
nand U8761 (N_8761,N_8169,N_8419);
and U8762 (N_8762,N_8335,N_8224);
or U8763 (N_8763,N_8454,N_8208);
and U8764 (N_8764,N_8414,N_8353);
xor U8765 (N_8765,N_8284,N_8119);
nor U8766 (N_8766,N_8130,N_8305);
and U8767 (N_8767,N_8067,N_8316);
nand U8768 (N_8768,N_8428,N_8448);
and U8769 (N_8769,N_8309,N_8363);
or U8770 (N_8770,N_8163,N_8149);
nand U8771 (N_8771,N_8164,N_8306);
xor U8772 (N_8772,N_8191,N_8489);
nor U8773 (N_8773,N_8079,N_8331);
or U8774 (N_8774,N_8461,N_8361);
nand U8775 (N_8775,N_8396,N_8196);
nand U8776 (N_8776,N_8101,N_8443);
nand U8777 (N_8777,N_8448,N_8017);
or U8778 (N_8778,N_8210,N_8301);
nand U8779 (N_8779,N_8246,N_8289);
nor U8780 (N_8780,N_8079,N_8087);
or U8781 (N_8781,N_8064,N_8148);
or U8782 (N_8782,N_8304,N_8243);
or U8783 (N_8783,N_8235,N_8377);
and U8784 (N_8784,N_8208,N_8423);
nor U8785 (N_8785,N_8164,N_8161);
xnor U8786 (N_8786,N_8258,N_8002);
and U8787 (N_8787,N_8035,N_8200);
or U8788 (N_8788,N_8434,N_8353);
xor U8789 (N_8789,N_8365,N_8413);
nand U8790 (N_8790,N_8450,N_8323);
xnor U8791 (N_8791,N_8148,N_8278);
and U8792 (N_8792,N_8313,N_8176);
xnor U8793 (N_8793,N_8047,N_8035);
nand U8794 (N_8794,N_8399,N_8431);
and U8795 (N_8795,N_8204,N_8103);
xor U8796 (N_8796,N_8087,N_8122);
and U8797 (N_8797,N_8491,N_8150);
xor U8798 (N_8798,N_8455,N_8156);
or U8799 (N_8799,N_8332,N_8009);
nand U8800 (N_8800,N_8435,N_8485);
nor U8801 (N_8801,N_8036,N_8155);
nand U8802 (N_8802,N_8309,N_8401);
nand U8803 (N_8803,N_8187,N_8069);
nor U8804 (N_8804,N_8227,N_8304);
nor U8805 (N_8805,N_8077,N_8413);
nand U8806 (N_8806,N_8377,N_8183);
nand U8807 (N_8807,N_8082,N_8397);
or U8808 (N_8808,N_8356,N_8481);
xnor U8809 (N_8809,N_8054,N_8178);
nor U8810 (N_8810,N_8436,N_8384);
xnor U8811 (N_8811,N_8277,N_8487);
or U8812 (N_8812,N_8100,N_8492);
xnor U8813 (N_8813,N_8325,N_8261);
and U8814 (N_8814,N_8004,N_8371);
and U8815 (N_8815,N_8066,N_8294);
xnor U8816 (N_8816,N_8085,N_8141);
xor U8817 (N_8817,N_8268,N_8219);
and U8818 (N_8818,N_8095,N_8102);
and U8819 (N_8819,N_8236,N_8149);
xor U8820 (N_8820,N_8069,N_8125);
and U8821 (N_8821,N_8169,N_8487);
xor U8822 (N_8822,N_8097,N_8422);
and U8823 (N_8823,N_8478,N_8323);
nor U8824 (N_8824,N_8434,N_8243);
nor U8825 (N_8825,N_8313,N_8283);
nand U8826 (N_8826,N_8178,N_8253);
or U8827 (N_8827,N_8361,N_8185);
nand U8828 (N_8828,N_8402,N_8215);
nand U8829 (N_8829,N_8212,N_8132);
nand U8830 (N_8830,N_8126,N_8178);
or U8831 (N_8831,N_8289,N_8158);
nor U8832 (N_8832,N_8043,N_8367);
or U8833 (N_8833,N_8363,N_8480);
and U8834 (N_8834,N_8035,N_8187);
nor U8835 (N_8835,N_8322,N_8112);
nor U8836 (N_8836,N_8427,N_8407);
and U8837 (N_8837,N_8229,N_8167);
nor U8838 (N_8838,N_8388,N_8343);
and U8839 (N_8839,N_8406,N_8306);
and U8840 (N_8840,N_8261,N_8267);
nand U8841 (N_8841,N_8336,N_8075);
or U8842 (N_8842,N_8165,N_8015);
xnor U8843 (N_8843,N_8281,N_8260);
nor U8844 (N_8844,N_8078,N_8144);
nor U8845 (N_8845,N_8388,N_8433);
xor U8846 (N_8846,N_8226,N_8151);
and U8847 (N_8847,N_8205,N_8071);
or U8848 (N_8848,N_8171,N_8277);
or U8849 (N_8849,N_8428,N_8468);
xor U8850 (N_8850,N_8483,N_8112);
nand U8851 (N_8851,N_8008,N_8031);
and U8852 (N_8852,N_8114,N_8380);
xor U8853 (N_8853,N_8001,N_8474);
and U8854 (N_8854,N_8202,N_8120);
and U8855 (N_8855,N_8124,N_8168);
nor U8856 (N_8856,N_8199,N_8122);
or U8857 (N_8857,N_8480,N_8403);
nor U8858 (N_8858,N_8415,N_8330);
nor U8859 (N_8859,N_8067,N_8092);
or U8860 (N_8860,N_8307,N_8039);
nand U8861 (N_8861,N_8284,N_8063);
nor U8862 (N_8862,N_8319,N_8440);
nand U8863 (N_8863,N_8300,N_8420);
nor U8864 (N_8864,N_8184,N_8035);
nor U8865 (N_8865,N_8484,N_8427);
xor U8866 (N_8866,N_8171,N_8135);
nor U8867 (N_8867,N_8343,N_8276);
nor U8868 (N_8868,N_8246,N_8112);
or U8869 (N_8869,N_8211,N_8377);
or U8870 (N_8870,N_8384,N_8288);
nor U8871 (N_8871,N_8183,N_8288);
or U8872 (N_8872,N_8413,N_8276);
and U8873 (N_8873,N_8347,N_8143);
nor U8874 (N_8874,N_8315,N_8246);
nand U8875 (N_8875,N_8432,N_8112);
and U8876 (N_8876,N_8339,N_8391);
nand U8877 (N_8877,N_8348,N_8100);
nor U8878 (N_8878,N_8416,N_8223);
nand U8879 (N_8879,N_8153,N_8154);
xnor U8880 (N_8880,N_8104,N_8480);
and U8881 (N_8881,N_8021,N_8212);
xor U8882 (N_8882,N_8408,N_8466);
nor U8883 (N_8883,N_8415,N_8137);
or U8884 (N_8884,N_8326,N_8443);
or U8885 (N_8885,N_8272,N_8153);
nor U8886 (N_8886,N_8139,N_8117);
xnor U8887 (N_8887,N_8018,N_8072);
nand U8888 (N_8888,N_8192,N_8102);
nand U8889 (N_8889,N_8163,N_8407);
xor U8890 (N_8890,N_8384,N_8286);
xor U8891 (N_8891,N_8198,N_8454);
xor U8892 (N_8892,N_8309,N_8367);
nor U8893 (N_8893,N_8476,N_8157);
nand U8894 (N_8894,N_8441,N_8046);
and U8895 (N_8895,N_8048,N_8004);
nor U8896 (N_8896,N_8160,N_8071);
or U8897 (N_8897,N_8364,N_8170);
nand U8898 (N_8898,N_8440,N_8235);
and U8899 (N_8899,N_8158,N_8262);
or U8900 (N_8900,N_8231,N_8210);
and U8901 (N_8901,N_8385,N_8267);
xor U8902 (N_8902,N_8008,N_8064);
or U8903 (N_8903,N_8236,N_8184);
xnor U8904 (N_8904,N_8203,N_8002);
or U8905 (N_8905,N_8347,N_8089);
nor U8906 (N_8906,N_8192,N_8139);
nand U8907 (N_8907,N_8101,N_8398);
or U8908 (N_8908,N_8248,N_8192);
nand U8909 (N_8909,N_8358,N_8064);
and U8910 (N_8910,N_8485,N_8214);
or U8911 (N_8911,N_8470,N_8152);
or U8912 (N_8912,N_8043,N_8033);
nand U8913 (N_8913,N_8242,N_8341);
xnor U8914 (N_8914,N_8173,N_8492);
and U8915 (N_8915,N_8364,N_8093);
nor U8916 (N_8916,N_8328,N_8028);
or U8917 (N_8917,N_8210,N_8371);
nand U8918 (N_8918,N_8365,N_8454);
nor U8919 (N_8919,N_8187,N_8170);
nand U8920 (N_8920,N_8375,N_8466);
xor U8921 (N_8921,N_8341,N_8169);
and U8922 (N_8922,N_8167,N_8390);
nor U8923 (N_8923,N_8402,N_8167);
nor U8924 (N_8924,N_8141,N_8369);
nand U8925 (N_8925,N_8273,N_8386);
nor U8926 (N_8926,N_8062,N_8489);
or U8927 (N_8927,N_8474,N_8254);
and U8928 (N_8928,N_8155,N_8331);
and U8929 (N_8929,N_8034,N_8092);
and U8930 (N_8930,N_8439,N_8185);
xnor U8931 (N_8931,N_8498,N_8073);
or U8932 (N_8932,N_8414,N_8124);
or U8933 (N_8933,N_8238,N_8192);
or U8934 (N_8934,N_8112,N_8491);
nand U8935 (N_8935,N_8422,N_8298);
nand U8936 (N_8936,N_8395,N_8056);
nor U8937 (N_8937,N_8301,N_8098);
nor U8938 (N_8938,N_8416,N_8435);
xor U8939 (N_8939,N_8209,N_8059);
xor U8940 (N_8940,N_8485,N_8310);
nand U8941 (N_8941,N_8333,N_8489);
xnor U8942 (N_8942,N_8272,N_8411);
nor U8943 (N_8943,N_8003,N_8127);
or U8944 (N_8944,N_8482,N_8229);
nand U8945 (N_8945,N_8436,N_8151);
and U8946 (N_8946,N_8386,N_8354);
nor U8947 (N_8947,N_8193,N_8348);
or U8948 (N_8948,N_8434,N_8160);
and U8949 (N_8949,N_8259,N_8195);
or U8950 (N_8950,N_8260,N_8354);
xor U8951 (N_8951,N_8214,N_8156);
nor U8952 (N_8952,N_8272,N_8364);
or U8953 (N_8953,N_8015,N_8169);
nor U8954 (N_8954,N_8255,N_8269);
or U8955 (N_8955,N_8156,N_8468);
nor U8956 (N_8956,N_8203,N_8207);
xor U8957 (N_8957,N_8426,N_8119);
nand U8958 (N_8958,N_8226,N_8054);
nor U8959 (N_8959,N_8260,N_8479);
xor U8960 (N_8960,N_8315,N_8344);
or U8961 (N_8961,N_8415,N_8336);
nor U8962 (N_8962,N_8130,N_8463);
and U8963 (N_8963,N_8260,N_8437);
xor U8964 (N_8964,N_8380,N_8237);
nor U8965 (N_8965,N_8108,N_8052);
nand U8966 (N_8966,N_8451,N_8094);
nand U8967 (N_8967,N_8167,N_8133);
nand U8968 (N_8968,N_8344,N_8462);
xnor U8969 (N_8969,N_8489,N_8009);
xor U8970 (N_8970,N_8493,N_8188);
nand U8971 (N_8971,N_8096,N_8279);
nand U8972 (N_8972,N_8349,N_8008);
or U8973 (N_8973,N_8273,N_8470);
and U8974 (N_8974,N_8017,N_8497);
and U8975 (N_8975,N_8349,N_8258);
or U8976 (N_8976,N_8079,N_8480);
nor U8977 (N_8977,N_8016,N_8353);
or U8978 (N_8978,N_8134,N_8294);
xnor U8979 (N_8979,N_8429,N_8419);
xnor U8980 (N_8980,N_8049,N_8002);
nand U8981 (N_8981,N_8391,N_8041);
nand U8982 (N_8982,N_8198,N_8475);
nand U8983 (N_8983,N_8071,N_8168);
and U8984 (N_8984,N_8484,N_8128);
or U8985 (N_8985,N_8091,N_8377);
or U8986 (N_8986,N_8100,N_8283);
or U8987 (N_8987,N_8469,N_8242);
nand U8988 (N_8988,N_8029,N_8008);
xor U8989 (N_8989,N_8076,N_8375);
nor U8990 (N_8990,N_8380,N_8249);
xnor U8991 (N_8991,N_8131,N_8219);
or U8992 (N_8992,N_8283,N_8404);
and U8993 (N_8993,N_8364,N_8457);
and U8994 (N_8994,N_8067,N_8392);
or U8995 (N_8995,N_8175,N_8072);
xor U8996 (N_8996,N_8263,N_8165);
xor U8997 (N_8997,N_8059,N_8474);
or U8998 (N_8998,N_8033,N_8329);
nand U8999 (N_8999,N_8027,N_8124);
nand U9000 (N_9000,N_8867,N_8973);
nand U9001 (N_9001,N_8727,N_8598);
or U9002 (N_9002,N_8741,N_8955);
nor U9003 (N_9003,N_8710,N_8987);
nor U9004 (N_9004,N_8768,N_8630);
xor U9005 (N_9005,N_8743,N_8798);
and U9006 (N_9006,N_8731,N_8652);
or U9007 (N_9007,N_8990,N_8542);
and U9008 (N_9008,N_8999,N_8528);
xor U9009 (N_9009,N_8986,N_8769);
nor U9010 (N_9010,N_8933,N_8570);
and U9011 (N_9011,N_8941,N_8690);
or U9012 (N_9012,N_8832,N_8762);
and U9013 (N_9013,N_8602,N_8868);
xor U9014 (N_9014,N_8548,N_8527);
xnor U9015 (N_9015,N_8526,N_8959);
nor U9016 (N_9016,N_8709,N_8782);
and U9017 (N_9017,N_8626,N_8500);
and U9018 (N_9018,N_8529,N_8827);
nand U9019 (N_9019,N_8755,N_8887);
nor U9020 (N_9020,N_8979,N_8681);
nand U9021 (N_9021,N_8616,N_8779);
and U9022 (N_9022,N_8932,N_8756);
and U9023 (N_9023,N_8549,N_8845);
nand U9024 (N_9024,N_8840,N_8924);
xor U9025 (N_9025,N_8670,N_8894);
xnor U9026 (N_9026,N_8774,N_8927);
nor U9027 (N_9027,N_8844,N_8574);
nand U9028 (N_9028,N_8884,N_8573);
nand U9029 (N_9029,N_8907,N_8882);
nand U9030 (N_9030,N_8917,N_8898);
nand U9031 (N_9031,N_8651,N_8722);
and U9032 (N_9032,N_8783,N_8878);
nor U9033 (N_9033,N_8596,N_8956);
xor U9034 (N_9034,N_8682,N_8708);
and U9035 (N_9035,N_8928,N_8974);
nand U9036 (N_9036,N_8629,N_8823);
or U9037 (N_9037,N_8846,N_8981);
and U9038 (N_9038,N_8833,N_8988);
or U9039 (N_9039,N_8648,N_8623);
or U9040 (N_9040,N_8749,N_8522);
or U9041 (N_9041,N_8516,N_8804);
nand U9042 (N_9042,N_8880,N_8584);
nor U9043 (N_9043,N_8506,N_8874);
xnor U9044 (N_9044,N_8938,N_8891);
or U9045 (N_9045,N_8655,N_8978);
and U9046 (N_9046,N_8712,N_8657);
and U9047 (N_9047,N_8591,N_8617);
or U9048 (N_9048,N_8696,N_8866);
nor U9049 (N_9049,N_8767,N_8537);
and U9050 (N_9050,N_8552,N_8571);
nor U9051 (N_9051,N_8951,N_8806);
xor U9052 (N_9052,N_8966,N_8847);
and U9053 (N_9053,N_8568,N_8675);
nor U9054 (N_9054,N_8634,N_8523);
and U9055 (N_9055,N_8638,N_8948);
xnor U9056 (N_9056,N_8699,N_8635);
xnor U9057 (N_9057,N_8647,N_8872);
nor U9058 (N_9058,N_8965,N_8740);
nand U9059 (N_9059,N_8569,N_8993);
and U9060 (N_9060,N_8751,N_8983);
and U9061 (N_9061,N_8923,N_8685);
xor U9062 (N_9062,N_8802,N_8621);
nor U9063 (N_9063,N_8539,N_8796);
xnor U9064 (N_9064,N_8788,N_8739);
nand U9065 (N_9065,N_8998,N_8953);
nor U9066 (N_9066,N_8614,N_8615);
nor U9067 (N_9067,N_8995,N_8888);
xnor U9068 (N_9068,N_8825,N_8915);
xnor U9069 (N_9069,N_8794,N_8579);
xnor U9070 (N_9070,N_8772,N_8989);
nor U9071 (N_9071,N_8719,N_8892);
and U9072 (N_9072,N_8771,N_8509);
nor U9073 (N_9073,N_8885,N_8581);
nor U9074 (N_9074,N_8831,N_8566);
or U9075 (N_9075,N_8814,N_8733);
or U9076 (N_9076,N_8922,N_8795);
xor U9077 (N_9077,N_8778,N_8534);
nor U9078 (N_9078,N_8883,N_8715);
nand U9079 (N_9079,N_8991,N_8780);
nand U9080 (N_9080,N_8590,N_8817);
nand U9081 (N_9081,N_8854,N_8513);
xnor U9082 (N_9082,N_8736,N_8962);
xor U9083 (N_9083,N_8656,N_8625);
xnor U9084 (N_9084,N_8575,N_8930);
nor U9085 (N_9085,N_8809,N_8863);
nor U9086 (N_9086,N_8687,N_8861);
xnor U9087 (N_9087,N_8912,N_8906);
nand U9088 (N_9088,N_8619,N_8641);
xor U9089 (N_9089,N_8692,N_8747);
xor U9090 (N_9090,N_8559,N_8632);
nor U9091 (N_9091,N_8934,N_8913);
and U9092 (N_9092,N_8673,N_8787);
and U9093 (N_9093,N_8726,N_8875);
nor U9094 (N_9094,N_8627,N_8577);
and U9095 (N_9095,N_8902,N_8903);
xor U9096 (N_9096,N_8609,N_8925);
and U9097 (N_9097,N_8698,N_8658);
nor U9098 (N_9098,N_8578,N_8889);
or U9099 (N_9099,N_8781,N_8611);
nor U9100 (N_9100,N_8791,N_8737);
or U9101 (N_9101,N_8760,N_8562);
nand U9102 (N_9102,N_8608,N_8518);
nand U9103 (N_9103,N_8856,N_8654);
or U9104 (N_9104,N_8536,N_8554);
nor U9105 (N_9105,N_8838,N_8954);
nand U9106 (N_9106,N_8950,N_8639);
nor U9107 (N_9107,N_8645,N_8807);
or U9108 (N_9108,N_8843,N_8969);
xnor U9109 (N_9109,N_8797,N_8680);
and U9110 (N_9110,N_8836,N_8700);
nor U9111 (N_9111,N_8663,N_8944);
and U9112 (N_9112,N_8541,N_8646);
or U9113 (N_9113,N_8612,N_8855);
and U9114 (N_9114,N_8734,N_8716);
or U9115 (N_9115,N_8775,N_8721);
or U9116 (N_9116,N_8752,N_8517);
and U9117 (N_9117,N_8770,N_8968);
nor U9118 (N_9118,N_8553,N_8653);
and U9119 (N_9119,N_8507,N_8811);
and U9120 (N_9120,N_8904,N_8929);
xor U9121 (N_9121,N_8703,N_8560);
and U9122 (N_9122,N_8865,N_8557);
or U9123 (N_9123,N_8600,N_8587);
nor U9124 (N_9124,N_8714,N_8588);
xnor U9125 (N_9125,N_8662,N_8786);
xor U9126 (N_9126,N_8693,N_8785);
and U9127 (N_9127,N_8815,N_8533);
and U9128 (N_9128,N_8538,N_8631);
nor U9129 (N_9129,N_8725,N_8812);
and U9130 (N_9130,N_8697,N_8940);
xor U9131 (N_9131,N_8567,N_8586);
and U9132 (N_9132,N_8821,N_8605);
and U9133 (N_9133,N_8871,N_8881);
nand U9134 (N_9134,N_8684,N_8593);
or U9135 (N_9135,N_8947,N_8618);
nor U9136 (N_9136,N_8558,N_8677);
xor U9137 (N_9137,N_8784,N_8637);
and U9138 (N_9138,N_8848,N_8563);
and U9139 (N_9139,N_8723,N_8551);
nand U9140 (N_9140,N_8985,N_8592);
or U9141 (N_9141,N_8572,N_8544);
nand U9142 (N_9142,N_8742,N_8624);
and U9143 (N_9143,N_8659,N_8744);
and U9144 (N_9144,N_8899,N_8705);
or U9145 (N_9145,N_8695,N_8642);
nor U9146 (N_9146,N_8818,N_8668);
or U9147 (N_9147,N_8543,N_8508);
or U9148 (N_9148,N_8839,N_8547);
or U9149 (N_9149,N_8620,N_8607);
and U9150 (N_9150,N_8688,N_8750);
and U9151 (N_9151,N_8644,N_8897);
nand U9152 (N_9152,N_8873,N_8852);
and U9153 (N_9153,N_8728,N_8819);
nand U9154 (N_9154,N_8519,N_8961);
nor U9155 (N_9155,N_8893,N_8801);
xnor U9156 (N_9156,N_8900,N_8958);
and U9157 (N_9157,N_8841,N_8765);
nor U9158 (N_9158,N_8870,N_8972);
nand U9159 (N_9159,N_8503,N_8975);
or U9160 (N_9160,N_8510,N_8957);
nor U9161 (N_9161,N_8540,N_8665);
and U9162 (N_9162,N_8674,N_8911);
nor U9163 (N_9163,N_8980,N_8816);
nand U9164 (N_9164,N_8920,N_8800);
nor U9165 (N_9165,N_8810,N_8691);
and U9166 (N_9166,N_8860,N_8758);
or U9167 (N_9167,N_8724,N_8515);
nand U9168 (N_9168,N_8976,N_8679);
and U9169 (N_9169,N_8859,N_8594);
xor U9170 (N_9170,N_8994,N_8753);
xnor U9171 (N_9171,N_8711,N_8945);
xor U9172 (N_9172,N_8820,N_8908);
nand U9173 (N_9173,N_8550,N_8745);
nand U9174 (N_9174,N_8876,N_8582);
nor U9175 (N_9175,N_8713,N_8761);
and U9176 (N_9176,N_8546,N_8501);
xnor U9177 (N_9177,N_8704,N_8813);
nor U9178 (N_9178,N_8921,N_8960);
nand U9179 (N_9179,N_8606,N_8792);
nor U9180 (N_9180,N_8901,N_8776);
nand U9181 (N_9181,N_8514,N_8970);
nor U9182 (N_9182,N_8849,N_8996);
and U9183 (N_9183,N_8597,N_8610);
nand U9184 (N_9184,N_8803,N_8520);
or U9185 (N_9185,N_8763,N_8826);
xnor U9186 (N_9186,N_8850,N_8585);
xnor U9187 (N_9187,N_8759,N_8525);
nand U9188 (N_9188,N_8909,N_8822);
nor U9189 (N_9189,N_8853,N_8748);
xnor U9190 (N_9190,N_8671,N_8946);
and U9191 (N_9191,N_8735,N_8511);
nor U9192 (N_9192,N_8936,N_8754);
nor U9193 (N_9193,N_8601,N_8524);
and U9194 (N_9194,N_8650,N_8676);
xor U9195 (N_9195,N_8678,N_8561);
or U9196 (N_9196,N_8512,N_8649);
xor U9197 (N_9197,N_8580,N_8706);
or U9198 (N_9198,N_8565,N_8857);
or U9199 (N_9199,N_8701,N_8757);
nor U9200 (N_9200,N_8683,N_8689);
nand U9201 (N_9201,N_8686,N_8837);
xor U9202 (N_9202,N_8746,N_8835);
nor U9203 (N_9203,N_8555,N_8952);
nand U9204 (N_9204,N_8877,N_8694);
xor U9205 (N_9205,N_8643,N_8521);
or U9206 (N_9206,N_8895,N_8707);
nand U9207 (N_9207,N_8977,N_8729);
nand U9208 (N_9208,N_8717,N_8842);
and U9209 (N_9209,N_8931,N_8599);
or U9210 (N_9210,N_8531,N_8982);
xor U9211 (N_9211,N_8622,N_8949);
or U9212 (N_9212,N_8914,N_8502);
nand U9213 (N_9213,N_8926,N_8943);
xor U9214 (N_9214,N_8666,N_8862);
and U9215 (N_9215,N_8777,N_8789);
xnor U9216 (N_9216,N_8919,N_8805);
and U9217 (N_9217,N_8613,N_8504);
and U9218 (N_9218,N_8738,N_8764);
and U9219 (N_9219,N_8971,N_8829);
or U9220 (N_9220,N_8702,N_8808);
nand U9221 (N_9221,N_8916,N_8633);
and U9222 (N_9222,N_8636,N_8718);
nand U9223 (N_9223,N_8997,N_8773);
xor U9224 (N_9224,N_8505,N_8660);
or U9225 (N_9225,N_8939,N_8640);
xnor U9226 (N_9226,N_8793,N_8790);
nor U9227 (N_9227,N_8890,N_8669);
or U9228 (N_9228,N_8963,N_8667);
and U9229 (N_9229,N_8964,N_8918);
nand U9230 (N_9230,N_8858,N_8589);
and U9231 (N_9231,N_8830,N_8564);
nand U9232 (N_9232,N_8879,N_8851);
nand U9233 (N_9233,N_8664,N_8672);
or U9234 (N_9234,N_8799,N_8992);
xnor U9235 (N_9235,N_8730,N_8967);
xor U9236 (N_9236,N_8910,N_8905);
and U9237 (N_9237,N_8545,N_8720);
nand U9238 (N_9238,N_8576,N_8896);
nand U9239 (N_9239,N_8604,N_8595);
or U9240 (N_9240,N_8824,N_8869);
xor U9241 (N_9241,N_8937,N_8535);
xnor U9242 (N_9242,N_8942,N_8532);
nand U9243 (N_9243,N_8661,N_8984);
or U9244 (N_9244,N_8886,N_8732);
nand U9245 (N_9245,N_8603,N_8583);
nand U9246 (N_9246,N_8530,N_8935);
xnor U9247 (N_9247,N_8556,N_8766);
nand U9248 (N_9248,N_8628,N_8834);
nand U9249 (N_9249,N_8864,N_8828);
or U9250 (N_9250,N_8826,N_8712);
and U9251 (N_9251,N_8689,N_8695);
or U9252 (N_9252,N_8703,N_8627);
nand U9253 (N_9253,N_8908,N_8990);
xnor U9254 (N_9254,N_8623,N_8602);
xor U9255 (N_9255,N_8596,N_8673);
and U9256 (N_9256,N_8701,N_8623);
xor U9257 (N_9257,N_8688,N_8797);
or U9258 (N_9258,N_8827,N_8605);
or U9259 (N_9259,N_8988,N_8832);
and U9260 (N_9260,N_8531,N_8583);
xnor U9261 (N_9261,N_8947,N_8979);
or U9262 (N_9262,N_8660,N_8618);
or U9263 (N_9263,N_8972,N_8602);
xor U9264 (N_9264,N_8531,N_8854);
nand U9265 (N_9265,N_8525,N_8505);
or U9266 (N_9266,N_8947,N_8609);
or U9267 (N_9267,N_8829,N_8826);
nand U9268 (N_9268,N_8648,N_8859);
and U9269 (N_9269,N_8667,N_8570);
nand U9270 (N_9270,N_8746,N_8547);
nor U9271 (N_9271,N_8687,N_8587);
and U9272 (N_9272,N_8762,N_8651);
xnor U9273 (N_9273,N_8679,N_8947);
nand U9274 (N_9274,N_8520,N_8743);
xnor U9275 (N_9275,N_8714,N_8848);
nor U9276 (N_9276,N_8831,N_8992);
and U9277 (N_9277,N_8727,N_8958);
or U9278 (N_9278,N_8527,N_8734);
nand U9279 (N_9279,N_8766,N_8569);
xor U9280 (N_9280,N_8678,N_8841);
nand U9281 (N_9281,N_8884,N_8562);
nand U9282 (N_9282,N_8770,N_8813);
or U9283 (N_9283,N_8804,N_8862);
nor U9284 (N_9284,N_8931,N_8846);
or U9285 (N_9285,N_8931,N_8810);
nand U9286 (N_9286,N_8943,N_8536);
xnor U9287 (N_9287,N_8547,N_8508);
nor U9288 (N_9288,N_8751,N_8742);
xnor U9289 (N_9289,N_8959,N_8872);
xnor U9290 (N_9290,N_8600,N_8773);
nand U9291 (N_9291,N_8795,N_8740);
nor U9292 (N_9292,N_8522,N_8664);
and U9293 (N_9293,N_8589,N_8616);
or U9294 (N_9294,N_8912,N_8635);
nor U9295 (N_9295,N_8911,N_8970);
nand U9296 (N_9296,N_8685,N_8941);
nand U9297 (N_9297,N_8793,N_8870);
xor U9298 (N_9298,N_8573,N_8549);
nand U9299 (N_9299,N_8608,N_8943);
nor U9300 (N_9300,N_8533,N_8942);
or U9301 (N_9301,N_8742,N_8719);
xnor U9302 (N_9302,N_8521,N_8553);
xnor U9303 (N_9303,N_8548,N_8920);
and U9304 (N_9304,N_8522,N_8945);
and U9305 (N_9305,N_8824,N_8668);
nand U9306 (N_9306,N_8951,N_8867);
xor U9307 (N_9307,N_8809,N_8946);
or U9308 (N_9308,N_8827,N_8934);
nand U9309 (N_9309,N_8640,N_8576);
or U9310 (N_9310,N_8530,N_8924);
xor U9311 (N_9311,N_8791,N_8685);
and U9312 (N_9312,N_8672,N_8621);
nor U9313 (N_9313,N_8720,N_8574);
or U9314 (N_9314,N_8678,N_8624);
or U9315 (N_9315,N_8682,N_8687);
xor U9316 (N_9316,N_8887,N_8500);
nand U9317 (N_9317,N_8750,N_8721);
xnor U9318 (N_9318,N_8611,N_8556);
nor U9319 (N_9319,N_8780,N_8737);
and U9320 (N_9320,N_8639,N_8787);
nand U9321 (N_9321,N_8912,N_8864);
nand U9322 (N_9322,N_8518,N_8936);
or U9323 (N_9323,N_8758,N_8688);
nand U9324 (N_9324,N_8512,N_8835);
nand U9325 (N_9325,N_8659,N_8589);
and U9326 (N_9326,N_8962,N_8761);
and U9327 (N_9327,N_8586,N_8678);
or U9328 (N_9328,N_8786,N_8775);
nor U9329 (N_9329,N_8816,N_8624);
nand U9330 (N_9330,N_8508,N_8721);
nor U9331 (N_9331,N_8613,N_8866);
xnor U9332 (N_9332,N_8584,N_8565);
and U9333 (N_9333,N_8808,N_8664);
and U9334 (N_9334,N_8901,N_8564);
xnor U9335 (N_9335,N_8707,N_8815);
nor U9336 (N_9336,N_8768,N_8543);
nand U9337 (N_9337,N_8692,N_8667);
nor U9338 (N_9338,N_8569,N_8969);
or U9339 (N_9339,N_8751,N_8845);
and U9340 (N_9340,N_8550,N_8535);
nand U9341 (N_9341,N_8715,N_8897);
nand U9342 (N_9342,N_8885,N_8701);
nand U9343 (N_9343,N_8753,N_8780);
and U9344 (N_9344,N_8783,N_8974);
or U9345 (N_9345,N_8862,N_8964);
nor U9346 (N_9346,N_8516,N_8527);
or U9347 (N_9347,N_8745,N_8721);
or U9348 (N_9348,N_8593,N_8962);
nor U9349 (N_9349,N_8714,N_8694);
xnor U9350 (N_9350,N_8622,N_8676);
nand U9351 (N_9351,N_8908,N_8826);
and U9352 (N_9352,N_8683,N_8880);
or U9353 (N_9353,N_8552,N_8508);
and U9354 (N_9354,N_8694,N_8800);
xor U9355 (N_9355,N_8608,N_8535);
xor U9356 (N_9356,N_8938,N_8861);
or U9357 (N_9357,N_8554,N_8798);
and U9358 (N_9358,N_8902,N_8927);
or U9359 (N_9359,N_8652,N_8683);
nand U9360 (N_9360,N_8894,N_8665);
nand U9361 (N_9361,N_8895,N_8613);
nand U9362 (N_9362,N_8874,N_8578);
xnor U9363 (N_9363,N_8854,N_8748);
and U9364 (N_9364,N_8794,N_8611);
nand U9365 (N_9365,N_8728,N_8892);
nor U9366 (N_9366,N_8817,N_8815);
or U9367 (N_9367,N_8540,N_8700);
nand U9368 (N_9368,N_8782,N_8539);
nor U9369 (N_9369,N_8831,N_8652);
xor U9370 (N_9370,N_8988,N_8625);
or U9371 (N_9371,N_8581,N_8510);
xor U9372 (N_9372,N_8801,N_8999);
xnor U9373 (N_9373,N_8701,N_8914);
nor U9374 (N_9374,N_8837,N_8793);
nand U9375 (N_9375,N_8582,N_8669);
or U9376 (N_9376,N_8550,N_8611);
xnor U9377 (N_9377,N_8503,N_8664);
or U9378 (N_9378,N_8856,N_8653);
nor U9379 (N_9379,N_8946,N_8806);
nand U9380 (N_9380,N_8639,N_8599);
or U9381 (N_9381,N_8573,N_8698);
or U9382 (N_9382,N_8806,N_8755);
xor U9383 (N_9383,N_8644,N_8865);
nand U9384 (N_9384,N_8671,N_8940);
xor U9385 (N_9385,N_8821,N_8773);
nand U9386 (N_9386,N_8824,N_8606);
xnor U9387 (N_9387,N_8789,N_8975);
or U9388 (N_9388,N_8576,N_8759);
or U9389 (N_9389,N_8572,N_8705);
nor U9390 (N_9390,N_8547,N_8612);
nor U9391 (N_9391,N_8695,N_8572);
nor U9392 (N_9392,N_8802,N_8837);
nor U9393 (N_9393,N_8680,N_8672);
or U9394 (N_9394,N_8697,N_8830);
xnor U9395 (N_9395,N_8860,N_8898);
and U9396 (N_9396,N_8956,N_8936);
nor U9397 (N_9397,N_8876,N_8695);
or U9398 (N_9398,N_8789,N_8821);
nand U9399 (N_9399,N_8914,N_8944);
xnor U9400 (N_9400,N_8685,N_8575);
and U9401 (N_9401,N_8721,N_8692);
nor U9402 (N_9402,N_8618,N_8858);
and U9403 (N_9403,N_8621,N_8631);
nand U9404 (N_9404,N_8774,N_8791);
or U9405 (N_9405,N_8784,N_8856);
nor U9406 (N_9406,N_8982,N_8656);
nand U9407 (N_9407,N_8611,N_8569);
nand U9408 (N_9408,N_8700,N_8766);
or U9409 (N_9409,N_8633,N_8868);
xnor U9410 (N_9410,N_8978,N_8554);
nand U9411 (N_9411,N_8958,N_8790);
nand U9412 (N_9412,N_8648,N_8923);
and U9413 (N_9413,N_8722,N_8501);
nand U9414 (N_9414,N_8758,N_8934);
and U9415 (N_9415,N_8935,N_8908);
or U9416 (N_9416,N_8537,N_8555);
or U9417 (N_9417,N_8591,N_8783);
nand U9418 (N_9418,N_8543,N_8748);
nand U9419 (N_9419,N_8955,N_8726);
and U9420 (N_9420,N_8633,N_8601);
and U9421 (N_9421,N_8539,N_8576);
nor U9422 (N_9422,N_8789,N_8749);
or U9423 (N_9423,N_8573,N_8934);
and U9424 (N_9424,N_8829,N_8812);
and U9425 (N_9425,N_8756,N_8958);
xnor U9426 (N_9426,N_8754,N_8649);
or U9427 (N_9427,N_8634,N_8711);
and U9428 (N_9428,N_8552,N_8720);
or U9429 (N_9429,N_8617,N_8515);
nand U9430 (N_9430,N_8793,N_8849);
xor U9431 (N_9431,N_8581,N_8751);
xnor U9432 (N_9432,N_8948,N_8854);
or U9433 (N_9433,N_8721,N_8619);
xnor U9434 (N_9434,N_8853,N_8554);
xor U9435 (N_9435,N_8644,N_8716);
and U9436 (N_9436,N_8509,N_8913);
and U9437 (N_9437,N_8588,N_8880);
xnor U9438 (N_9438,N_8503,N_8816);
and U9439 (N_9439,N_8961,N_8832);
or U9440 (N_9440,N_8589,N_8861);
xnor U9441 (N_9441,N_8695,N_8829);
or U9442 (N_9442,N_8598,N_8638);
or U9443 (N_9443,N_8643,N_8841);
or U9444 (N_9444,N_8652,N_8979);
nor U9445 (N_9445,N_8736,N_8624);
xnor U9446 (N_9446,N_8519,N_8550);
nor U9447 (N_9447,N_8719,N_8668);
and U9448 (N_9448,N_8770,N_8565);
nand U9449 (N_9449,N_8870,N_8733);
and U9450 (N_9450,N_8602,N_8800);
xor U9451 (N_9451,N_8609,N_8567);
nand U9452 (N_9452,N_8771,N_8693);
nor U9453 (N_9453,N_8896,N_8651);
and U9454 (N_9454,N_8755,N_8857);
nand U9455 (N_9455,N_8672,N_8698);
and U9456 (N_9456,N_8879,N_8801);
or U9457 (N_9457,N_8692,N_8794);
xnor U9458 (N_9458,N_8595,N_8886);
or U9459 (N_9459,N_8698,N_8594);
nor U9460 (N_9460,N_8968,N_8928);
and U9461 (N_9461,N_8869,N_8619);
or U9462 (N_9462,N_8553,N_8969);
nor U9463 (N_9463,N_8644,N_8860);
and U9464 (N_9464,N_8628,N_8586);
nand U9465 (N_9465,N_8691,N_8865);
xnor U9466 (N_9466,N_8795,N_8759);
nor U9467 (N_9467,N_8514,N_8908);
xor U9468 (N_9468,N_8795,N_8981);
nand U9469 (N_9469,N_8964,N_8851);
nor U9470 (N_9470,N_8766,N_8866);
or U9471 (N_9471,N_8738,N_8678);
nor U9472 (N_9472,N_8947,N_8702);
or U9473 (N_9473,N_8681,N_8573);
nand U9474 (N_9474,N_8600,N_8670);
nand U9475 (N_9475,N_8617,N_8602);
nand U9476 (N_9476,N_8842,N_8940);
and U9477 (N_9477,N_8574,N_8644);
or U9478 (N_9478,N_8609,N_8855);
xor U9479 (N_9479,N_8776,N_8801);
and U9480 (N_9480,N_8967,N_8900);
xnor U9481 (N_9481,N_8635,N_8951);
nor U9482 (N_9482,N_8640,N_8548);
or U9483 (N_9483,N_8627,N_8973);
and U9484 (N_9484,N_8682,N_8567);
or U9485 (N_9485,N_8814,N_8639);
nand U9486 (N_9486,N_8938,N_8959);
xnor U9487 (N_9487,N_8694,N_8726);
nand U9488 (N_9488,N_8588,N_8506);
nand U9489 (N_9489,N_8711,N_8760);
nand U9490 (N_9490,N_8727,N_8606);
or U9491 (N_9491,N_8728,N_8532);
nor U9492 (N_9492,N_8911,N_8919);
xnor U9493 (N_9493,N_8650,N_8635);
and U9494 (N_9494,N_8793,N_8736);
nor U9495 (N_9495,N_8563,N_8789);
or U9496 (N_9496,N_8823,N_8808);
nor U9497 (N_9497,N_8589,N_8658);
nor U9498 (N_9498,N_8612,N_8938);
or U9499 (N_9499,N_8959,N_8670);
or U9500 (N_9500,N_9085,N_9288);
xor U9501 (N_9501,N_9223,N_9389);
nand U9502 (N_9502,N_9180,N_9276);
xnor U9503 (N_9503,N_9478,N_9075);
nand U9504 (N_9504,N_9256,N_9307);
and U9505 (N_9505,N_9321,N_9299);
nand U9506 (N_9506,N_9116,N_9442);
and U9507 (N_9507,N_9434,N_9117);
nor U9508 (N_9508,N_9016,N_9291);
nand U9509 (N_9509,N_9397,N_9462);
and U9510 (N_9510,N_9029,N_9103);
and U9511 (N_9511,N_9018,N_9104);
or U9512 (N_9512,N_9199,N_9025);
and U9513 (N_9513,N_9471,N_9242);
or U9514 (N_9514,N_9494,N_9190);
xnor U9515 (N_9515,N_9187,N_9363);
xor U9516 (N_9516,N_9469,N_9449);
xor U9517 (N_9517,N_9273,N_9165);
nand U9518 (N_9518,N_9414,N_9129);
nor U9519 (N_9519,N_9219,N_9289);
or U9520 (N_9520,N_9404,N_9428);
nand U9521 (N_9521,N_9057,N_9480);
or U9522 (N_9522,N_9416,N_9341);
and U9523 (N_9523,N_9311,N_9235);
xnor U9524 (N_9524,N_9308,N_9079);
and U9525 (N_9525,N_9037,N_9171);
nand U9526 (N_9526,N_9267,N_9159);
nor U9527 (N_9527,N_9230,N_9246);
nor U9528 (N_9528,N_9422,N_9010);
nor U9529 (N_9529,N_9192,N_9244);
or U9530 (N_9530,N_9176,N_9233);
and U9531 (N_9531,N_9327,N_9460);
nand U9532 (N_9532,N_9204,N_9101);
nand U9533 (N_9533,N_9063,N_9384);
nand U9534 (N_9534,N_9381,N_9465);
and U9535 (N_9535,N_9275,N_9350);
or U9536 (N_9536,N_9214,N_9445);
xor U9537 (N_9537,N_9053,N_9263);
and U9538 (N_9538,N_9292,N_9438);
and U9539 (N_9539,N_9495,N_9412);
nand U9540 (N_9540,N_9481,N_9021);
xnor U9541 (N_9541,N_9312,N_9323);
or U9542 (N_9542,N_9425,N_9186);
or U9543 (N_9543,N_9486,N_9185);
nor U9544 (N_9544,N_9090,N_9277);
nor U9545 (N_9545,N_9177,N_9143);
nand U9546 (N_9546,N_9139,N_9482);
nor U9547 (N_9547,N_9406,N_9232);
and U9548 (N_9548,N_9487,N_9490);
or U9549 (N_9549,N_9330,N_9038);
or U9550 (N_9550,N_9319,N_9255);
nor U9551 (N_9551,N_9357,N_9393);
and U9552 (N_9552,N_9064,N_9137);
xor U9553 (N_9553,N_9202,N_9172);
or U9554 (N_9554,N_9118,N_9184);
and U9555 (N_9555,N_9448,N_9208);
nand U9556 (N_9556,N_9375,N_9499);
xor U9557 (N_9557,N_9151,N_9066);
or U9558 (N_9558,N_9338,N_9413);
or U9559 (N_9559,N_9033,N_9476);
xnor U9560 (N_9560,N_9050,N_9074);
xor U9561 (N_9561,N_9089,N_9377);
or U9562 (N_9562,N_9394,N_9450);
and U9563 (N_9563,N_9240,N_9367);
nor U9564 (N_9564,N_9484,N_9212);
nand U9565 (N_9565,N_9441,N_9360);
nand U9566 (N_9566,N_9453,N_9382);
nand U9567 (N_9567,N_9022,N_9132);
nand U9568 (N_9568,N_9354,N_9007);
or U9569 (N_9569,N_9415,N_9169);
nor U9570 (N_9570,N_9138,N_9142);
xnor U9571 (N_9571,N_9083,N_9313);
and U9572 (N_9572,N_9433,N_9152);
nor U9573 (N_9573,N_9432,N_9194);
and U9574 (N_9574,N_9229,N_9300);
or U9575 (N_9575,N_9126,N_9174);
nand U9576 (N_9576,N_9004,N_9168);
nand U9577 (N_9577,N_9003,N_9226);
nor U9578 (N_9578,N_9294,N_9253);
xnor U9579 (N_9579,N_9454,N_9306);
nor U9580 (N_9580,N_9156,N_9221);
nor U9581 (N_9581,N_9279,N_9410);
nor U9582 (N_9582,N_9069,N_9150);
nand U9583 (N_9583,N_9077,N_9154);
and U9584 (N_9584,N_9466,N_9366);
or U9585 (N_9585,N_9098,N_9297);
xnor U9586 (N_9586,N_9125,N_9228);
and U9587 (N_9587,N_9041,N_9322);
or U9588 (N_9588,N_9144,N_9222);
and U9589 (N_9589,N_9254,N_9456);
and U9590 (N_9590,N_9402,N_9318);
xnor U9591 (N_9591,N_9076,N_9483);
nand U9592 (N_9592,N_9237,N_9418);
nor U9593 (N_9593,N_9468,N_9260);
or U9594 (N_9594,N_9348,N_9131);
and U9595 (N_9595,N_9113,N_9369);
xor U9596 (N_9596,N_9030,N_9305);
nor U9597 (N_9597,N_9258,N_9200);
xnor U9598 (N_9598,N_9455,N_9164);
xnor U9599 (N_9599,N_9191,N_9044);
nand U9600 (N_9600,N_9281,N_9100);
nor U9601 (N_9601,N_9274,N_9148);
nand U9602 (N_9602,N_9224,N_9019);
xor U9603 (N_9603,N_9400,N_9310);
nor U9604 (N_9604,N_9387,N_9087);
and U9605 (N_9605,N_9470,N_9000);
xnor U9606 (N_9606,N_9439,N_9122);
or U9607 (N_9607,N_9488,N_9259);
and U9608 (N_9608,N_9067,N_9461);
xnor U9609 (N_9609,N_9315,N_9163);
or U9610 (N_9610,N_9032,N_9409);
nand U9611 (N_9611,N_9343,N_9197);
or U9612 (N_9612,N_9395,N_9464);
xnor U9613 (N_9613,N_9374,N_9006);
nor U9614 (N_9614,N_9026,N_9155);
nand U9615 (N_9615,N_9405,N_9140);
and U9616 (N_9616,N_9206,N_9326);
nand U9617 (N_9617,N_9396,N_9436);
and U9618 (N_9618,N_9265,N_9115);
or U9619 (N_9619,N_9463,N_9092);
or U9620 (N_9620,N_9111,N_9241);
nor U9621 (N_9621,N_9302,N_9344);
or U9622 (N_9622,N_9303,N_9437);
and U9623 (N_9623,N_9012,N_9009);
and U9624 (N_9624,N_9001,N_9179);
xor U9625 (N_9625,N_9061,N_9385);
or U9626 (N_9626,N_9271,N_9331);
xor U9627 (N_9627,N_9280,N_9342);
nand U9628 (N_9628,N_9036,N_9178);
or U9629 (N_9629,N_9304,N_9268);
or U9630 (N_9630,N_9065,N_9234);
and U9631 (N_9631,N_9093,N_9049);
or U9632 (N_9632,N_9136,N_9209);
xnor U9633 (N_9633,N_9062,N_9024);
and U9634 (N_9634,N_9457,N_9058);
and U9635 (N_9635,N_9210,N_9112);
or U9636 (N_9636,N_9262,N_9349);
nand U9637 (N_9637,N_9105,N_9380);
nor U9638 (N_9638,N_9351,N_9121);
nor U9639 (N_9639,N_9011,N_9120);
nor U9640 (N_9640,N_9046,N_9290);
nor U9641 (N_9641,N_9239,N_9278);
and U9642 (N_9642,N_9134,N_9035);
xnor U9643 (N_9643,N_9479,N_9145);
and U9644 (N_9644,N_9316,N_9443);
and U9645 (N_9645,N_9023,N_9325);
nor U9646 (N_9646,N_9459,N_9467);
or U9647 (N_9647,N_9207,N_9107);
xnor U9648 (N_9648,N_9293,N_9379);
and U9649 (N_9649,N_9153,N_9346);
or U9650 (N_9650,N_9213,N_9272);
or U9651 (N_9651,N_9017,N_9160);
nor U9652 (N_9652,N_9146,N_9411);
or U9653 (N_9653,N_9446,N_9236);
nand U9654 (N_9654,N_9158,N_9020);
xor U9655 (N_9655,N_9141,N_9489);
xnor U9656 (N_9656,N_9328,N_9368);
and U9657 (N_9657,N_9261,N_9485);
or U9658 (N_9658,N_9095,N_9408);
and U9659 (N_9659,N_9225,N_9162);
or U9660 (N_9660,N_9336,N_9361);
nand U9661 (N_9661,N_9073,N_9055);
nor U9662 (N_9662,N_9094,N_9472);
or U9663 (N_9663,N_9216,N_9014);
or U9664 (N_9664,N_9283,N_9048);
nor U9665 (N_9665,N_9353,N_9345);
nor U9666 (N_9666,N_9421,N_9435);
or U9667 (N_9667,N_9243,N_9175);
or U9668 (N_9668,N_9364,N_9334);
nand U9669 (N_9669,N_9447,N_9250);
xnor U9670 (N_9670,N_9183,N_9320);
xnor U9671 (N_9671,N_9043,N_9072);
or U9672 (N_9672,N_9173,N_9440);
nor U9673 (N_9673,N_9161,N_9227);
nand U9674 (N_9674,N_9188,N_9252);
nand U9675 (N_9675,N_9170,N_9193);
or U9676 (N_9676,N_9135,N_9071);
and U9677 (N_9677,N_9403,N_9287);
nand U9678 (N_9678,N_9427,N_9376);
and U9679 (N_9679,N_9042,N_9096);
or U9680 (N_9680,N_9295,N_9081);
nand U9681 (N_9681,N_9355,N_9264);
nor U9682 (N_9682,N_9220,N_9429);
and U9683 (N_9683,N_9123,N_9039);
and U9684 (N_9684,N_9157,N_9109);
and U9685 (N_9685,N_9247,N_9056);
nand U9686 (N_9686,N_9119,N_9045);
or U9687 (N_9687,N_9091,N_9149);
or U9688 (N_9688,N_9215,N_9370);
or U9689 (N_9689,N_9238,N_9231);
nor U9690 (N_9690,N_9047,N_9359);
or U9691 (N_9691,N_9086,N_9201);
and U9692 (N_9692,N_9329,N_9270);
xor U9693 (N_9693,N_9110,N_9352);
nand U9694 (N_9694,N_9059,N_9124);
nor U9695 (N_9695,N_9181,N_9373);
or U9696 (N_9696,N_9420,N_9417);
xor U9697 (N_9697,N_9040,N_9008);
and U9698 (N_9698,N_9251,N_9401);
nor U9699 (N_9699,N_9496,N_9282);
nand U9700 (N_9700,N_9477,N_9068);
and U9701 (N_9701,N_9078,N_9108);
nand U9702 (N_9702,N_9013,N_9099);
nor U9703 (N_9703,N_9390,N_9386);
or U9704 (N_9704,N_9080,N_9266);
or U9705 (N_9705,N_9362,N_9082);
and U9706 (N_9706,N_9196,N_9027);
and U9707 (N_9707,N_9473,N_9195);
and U9708 (N_9708,N_9424,N_9431);
nor U9709 (N_9709,N_9317,N_9070);
nand U9710 (N_9710,N_9167,N_9114);
nor U9711 (N_9711,N_9189,N_9452);
and U9712 (N_9712,N_9339,N_9015);
or U9713 (N_9713,N_9031,N_9298);
nand U9714 (N_9714,N_9493,N_9218);
nand U9715 (N_9715,N_9419,N_9084);
nor U9716 (N_9716,N_9309,N_9407);
or U9717 (N_9717,N_9314,N_9269);
xnor U9718 (N_9718,N_9444,N_9127);
or U9719 (N_9719,N_9166,N_9133);
nand U9720 (N_9720,N_9106,N_9128);
nor U9721 (N_9721,N_9399,N_9248);
and U9722 (N_9722,N_9391,N_9383);
nand U9723 (N_9723,N_9217,N_9388);
and U9724 (N_9724,N_9497,N_9324);
and U9725 (N_9725,N_9130,N_9052);
or U9726 (N_9726,N_9296,N_9356);
and U9727 (N_9727,N_9002,N_9451);
or U9728 (N_9728,N_9423,N_9205);
nor U9729 (N_9729,N_9284,N_9430);
or U9730 (N_9730,N_9335,N_9392);
nor U9731 (N_9731,N_9347,N_9028);
nand U9732 (N_9732,N_9337,N_9333);
xnor U9733 (N_9733,N_9398,N_9458);
nand U9734 (N_9734,N_9203,N_9475);
nand U9735 (N_9735,N_9257,N_9198);
nand U9736 (N_9736,N_9365,N_9426);
or U9737 (N_9737,N_9245,N_9211);
nand U9738 (N_9738,N_9285,N_9060);
and U9739 (N_9739,N_9340,N_9051);
and U9740 (N_9740,N_9301,N_9498);
nand U9741 (N_9741,N_9088,N_9286);
nand U9742 (N_9742,N_9378,N_9034);
nand U9743 (N_9743,N_9182,N_9005);
or U9744 (N_9744,N_9358,N_9097);
nand U9745 (N_9745,N_9054,N_9372);
and U9746 (N_9746,N_9492,N_9332);
and U9747 (N_9747,N_9371,N_9491);
and U9748 (N_9748,N_9102,N_9249);
and U9749 (N_9749,N_9474,N_9147);
nor U9750 (N_9750,N_9413,N_9155);
and U9751 (N_9751,N_9325,N_9289);
xnor U9752 (N_9752,N_9144,N_9101);
nor U9753 (N_9753,N_9426,N_9020);
xnor U9754 (N_9754,N_9406,N_9298);
and U9755 (N_9755,N_9406,N_9104);
nor U9756 (N_9756,N_9237,N_9479);
and U9757 (N_9757,N_9036,N_9255);
and U9758 (N_9758,N_9418,N_9195);
xor U9759 (N_9759,N_9315,N_9387);
nor U9760 (N_9760,N_9268,N_9031);
xor U9761 (N_9761,N_9158,N_9226);
xnor U9762 (N_9762,N_9413,N_9103);
xor U9763 (N_9763,N_9047,N_9074);
xor U9764 (N_9764,N_9070,N_9374);
or U9765 (N_9765,N_9429,N_9344);
xnor U9766 (N_9766,N_9246,N_9420);
and U9767 (N_9767,N_9004,N_9327);
nor U9768 (N_9768,N_9145,N_9316);
xnor U9769 (N_9769,N_9224,N_9450);
and U9770 (N_9770,N_9196,N_9358);
nand U9771 (N_9771,N_9383,N_9054);
or U9772 (N_9772,N_9329,N_9187);
nand U9773 (N_9773,N_9435,N_9372);
nor U9774 (N_9774,N_9286,N_9296);
xnor U9775 (N_9775,N_9412,N_9348);
xnor U9776 (N_9776,N_9207,N_9113);
and U9777 (N_9777,N_9357,N_9364);
xnor U9778 (N_9778,N_9113,N_9219);
or U9779 (N_9779,N_9050,N_9434);
nor U9780 (N_9780,N_9123,N_9446);
nand U9781 (N_9781,N_9484,N_9004);
or U9782 (N_9782,N_9438,N_9079);
nand U9783 (N_9783,N_9410,N_9223);
nor U9784 (N_9784,N_9449,N_9187);
nor U9785 (N_9785,N_9229,N_9128);
nor U9786 (N_9786,N_9332,N_9390);
nand U9787 (N_9787,N_9499,N_9455);
nor U9788 (N_9788,N_9148,N_9191);
and U9789 (N_9789,N_9178,N_9446);
xnor U9790 (N_9790,N_9409,N_9175);
and U9791 (N_9791,N_9400,N_9497);
nand U9792 (N_9792,N_9293,N_9328);
and U9793 (N_9793,N_9418,N_9322);
nor U9794 (N_9794,N_9276,N_9145);
or U9795 (N_9795,N_9319,N_9491);
nand U9796 (N_9796,N_9088,N_9384);
and U9797 (N_9797,N_9377,N_9476);
nand U9798 (N_9798,N_9396,N_9033);
nor U9799 (N_9799,N_9252,N_9376);
xor U9800 (N_9800,N_9408,N_9423);
xor U9801 (N_9801,N_9483,N_9429);
nor U9802 (N_9802,N_9065,N_9341);
nor U9803 (N_9803,N_9376,N_9332);
xnor U9804 (N_9804,N_9407,N_9083);
nor U9805 (N_9805,N_9003,N_9053);
and U9806 (N_9806,N_9029,N_9314);
and U9807 (N_9807,N_9477,N_9180);
and U9808 (N_9808,N_9036,N_9261);
or U9809 (N_9809,N_9393,N_9309);
or U9810 (N_9810,N_9236,N_9117);
nand U9811 (N_9811,N_9364,N_9346);
and U9812 (N_9812,N_9449,N_9068);
and U9813 (N_9813,N_9265,N_9393);
nand U9814 (N_9814,N_9347,N_9079);
or U9815 (N_9815,N_9449,N_9313);
nor U9816 (N_9816,N_9226,N_9177);
or U9817 (N_9817,N_9191,N_9472);
nand U9818 (N_9818,N_9361,N_9359);
and U9819 (N_9819,N_9387,N_9098);
and U9820 (N_9820,N_9367,N_9363);
nand U9821 (N_9821,N_9248,N_9352);
or U9822 (N_9822,N_9226,N_9001);
and U9823 (N_9823,N_9133,N_9245);
or U9824 (N_9824,N_9488,N_9433);
xor U9825 (N_9825,N_9328,N_9257);
nand U9826 (N_9826,N_9421,N_9121);
nand U9827 (N_9827,N_9463,N_9207);
nand U9828 (N_9828,N_9237,N_9244);
and U9829 (N_9829,N_9051,N_9014);
nor U9830 (N_9830,N_9052,N_9152);
xnor U9831 (N_9831,N_9283,N_9368);
nor U9832 (N_9832,N_9054,N_9258);
xnor U9833 (N_9833,N_9431,N_9063);
and U9834 (N_9834,N_9319,N_9089);
nor U9835 (N_9835,N_9346,N_9479);
or U9836 (N_9836,N_9284,N_9426);
nor U9837 (N_9837,N_9447,N_9012);
or U9838 (N_9838,N_9001,N_9326);
xor U9839 (N_9839,N_9111,N_9281);
nand U9840 (N_9840,N_9246,N_9121);
nand U9841 (N_9841,N_9243,N_9459);
nand U9842 (N_9842,N_9467,N_9478);
xor U9843 (N_9843,N_9360,N_9171);
or U9844 (N_9844,N_9034,N_9315);
xor U9845 (N_9845,N_9201,N_9108);
and U9846 (N_9846,N_9249,N_9143);
nor U9847 (N_9847,N_9233,N_9349);
and U9848 (N_9848,N_9192,N_9444);
nor U9849 (N_9849,N_9401,N_9263);
nor U9850 (N_9850,N_9071,N_9152);
nor U9851 (N_9851,N_9192,N_9451);
and U9852 (N_9852,N_9431,N_9456);
or U9853 (N_9853,N_9407,N_9080);
nor U9854 (N_9854,N_9071,N_9204);
nor U9855 (N_9855,N_9441,N_9306);
nand U9856 (N_9856,N_9104,N_9278);
xnor U9857 (N_9857,N_9190,N_9425);
nor U9858 (N_9858,N_9363,N_9062);
nand U9859 (N_9859,N_9057,N_9230);
or U9860 (N_9860,N_9089,N_9492);
and U9861 (N_9861,N_9311,N_9128);
or U9862 (N_9862,N_9236,N_9342);
nor U9863 (N_9863,N_9265,N_9100);
or U9864 (N_9864,N_9359,N_9211);
or U9865 (N_9865,N_9460,N_9004);
nand U9866 (N_9866,N_9201,N_9439);
or U9867 (N_9867,N_9252,N_9394);
or U9868 (N_9868,N_9277,N_9435);
nand U9869 (N_9869,N_9090,N_9477);
xnor U9870 (N_9870,N_9073,N_9348);
or U9871 (N_9871,N_9346,N_9081);
nor U9872 (N_9872,N_9269,N_9289);
nor U9873 (N_9873,N_9020,N_9215);
nor U9874 (N_9874,N_9213,N_9433);
and U9875 (N_9875,N_9227,N_9183);
xnor U9876 (N_9876,N_9175,N_9350);
nor U9877 (N_9877,N_9229,N_9201);
xnor U9878 (N_9878,N_9291,N_9168);
nor U9879 (N_9879,N_9305,N_9154);
or U9880 (N_9880,N_9275,N_9258);
and U9881 (N_9881,N_9265,N_9094);
nor U9882 (N_9882,N_9173,N_9351);
nand U9883 (N_9883,N_9037,N_9463);
nand U9884 (N_9884,N_9256,N_9188);
xor U9885 (N_9885,N_9297,N_9469);
nand U9886 (N_9886,N_9115,N_9329);
and U9887 (N_9887,N_9400,N_9088);
nor U9888 (N_9888,N_9364,N_9466);
and U9889 (N_9889,N_9313,N_9148);
or U9890 (N_9890,N_9396,N_9272);
xnor U9891 (N_9891,N_9141,N_9415);
and U9892 (N_9892,N_9414,N_9051);
or U9893 (N_9893,N_9164,N_9440);
or U9894 (N_9894,N_9377,N_9122);
xnor U9895 (N_9895,N_9168,N_9266);
or U9896 (N_9896,N_9258,N_9247);
xor U9897 (N_9897,N_9370,N_9051);
nand U9898 (N_9898,N_9334,N_9365);
or U9899 (N_9899,N_9378,N_9431);
nand U9900 (N_9900,N_9216,N_9494);
nor U9901 (N_9901,N_9334,N_9357);
nor U9902 (N_9902,N_9067,N_9102);
xor U9903 (N_9903,N_9349,N_9384);
nand U9904 (N_9904,N_9112,N_9342);
or U9905 (N_9905,N_9196,N_9167);
xor U9906 (N_9906,N_9212,N_9480);
xnor U9907 (N_9907,N_9046,N_9026);
nor U9908 (N_9908,N_9084,N_9246);
and U9909 (N_9909,N_9081,N_9041);
nor U9910 (N_9910,N_9211,N_9420);
xnor U9911 (N_9911,N_9225,N_9094);
nor U9912 (N_9912,N_9278,N_9309);
xor U9913 (N_9913,N_9378,N_9047);
nor U9914 (N_9914,N_9097,N_9247);
xor U9915 (N_9915,N_9102,N_9370);
nor U9916 (N_9916,N_9243,N_9204);
and U9917 (N_9917,N_9341,N_9313);
nand U9918 (N_9918,N_9178,N_9318);
nor U9919 (N_9919,N_9466,N_9349);
nor U9920 (N_9920,N_9139,N_9132);
xor U9921 (N_9921,N_9180,N_9362);
nand U9922 (N_9922,N_9093,N_9262);
nand U9923 (N_9923,N_9012,N_9116);
xnor U9924 (N_9924,N_9050,N_9136);
nand U9925 (N_9925,N_9073,N_9313);
xor U9926 (N_9926,N_9149,N_9156);
or U9927 (N_9927,N_9105,N_9106);
and U9928 (N_9928,N_9343,N_9114);
xnor U9929 (N_9929,N_9254,N_9150);
and U9930 (N_9930,N_9449,N_9380);
nor U9931 (N_9931,N_9462,N_9464);
nor U9932 (N_9932,N_9046,N_9277);
xnor U9933 (N_9933,N_9092,N_9064);
xor U9934 (N_9934,N_9039,N_9167);
xnor U9935 (N_9935,N_9134,N_9409);
or U9936 (N_9936,N_9364,N_9267);
xor U9937 (N_9937,N_9201,N_9473);
xnor U9938 (N_9938,N_9199,N_9495);
nor U9939 (N_9939,N_9021,N_9355);
xnor U9940 (N_9940,N_9186,N_9208);
or U9941 (N_9941,N_9099,N_9103);
and U9942 (N_9942,N_9454,N_9334);
nand U9943 (N_9943,N_9111,N_9348);
nand U9944 (N_9944,N_9272,N_9259);
and U9945 (N_9945,N_9295,N_9014);
nor U9946 (N_9946,N_9277,N_9248);
and U9947 (N_9947,N_9319,N_9340);
xnor U9948 (N_9948,N_9496,N_9427);
nor U9949 (N_9949,N_9150,N_9248);
nor U9950 (N_9950,N_9279,N_9255);
or U9951 (N_9951,N_9019,N_9073);
xor U9952 (N_9952,N_9262,N_9462);
or U9953 (N_9953,N_9396,N_9073);
or U9954 (N_9954,N_9380,N_9081);
or U9955 (N_9955,N_9247,N_9163);
nor U9956 (N_9956,N_9419,N_9227);
xnor U9957 (N_9957,N_9115,N_9228);
or U9958 (N_9958,N_9474,N_9239);
nor U9959 (N_9959,N_9016,N_9141);
nor U9960 (N_9960,N_9239,N_9472);
nand U9961 (N_9961,N_9158,N_9023);
nor U9962 (N_9962,N_9155,N_9372);
and U9963 (N_9963,N_9093,N_9261);
or U9964 (N_9964,N_9483,N_9197);
and U9965 (N_9965,N_9259,N_9435);
xnor U9966 (N_9966,N_9091,N_9379);
xnor U9967 (N_9967,N_9414,N_9052);
xnor U9968 (N_9968,N_9410,N_9458);
and U9969 (N_9969,N_9489,N_9495);
and U9970 (N_9970,N_9025,N_9008);
nor U9971 (N_9971,N_9255,N_9237);
or U9972 (N_9972,N_9406,N_9414);
or U9973 (N_9973,N_9213,N_9108);
nand U9974 (N_9974,N_9245,N_9046);
nand U9975 (N_9975,N_9290,N_9135);
and U9976 (N_9976,N_9485,N_9408);
xor U9977 (N_9977,N_9212,N_9025);
nor U9978 (N_9978,N_9442,N_9030);
xor U9979 (N_9979,N_9046,N_9339);
nor U9980 (N_9980,N_9377,N_9429);
and U9981 (N_9981,N_9275,N_9087);
or U9982 (N_9982,N_9022,N_9437);
xnor U9983 (N_9983,N_9476,N_9354);
and U9984 (N_9984,N_9007,N_9300);
and U9985 (N_9985,N_9112,N_9350);
and U9986 (N_9986,N_9275,N_9172);
or U9987 (N_9987,N_9021,N_9076);
or U9988 (N_9988,N_9282,N_9208);
nor U9989 (N_9989,N_9046,N_9256);
nor U9990 (N_9990,N_9071,N_9206);
nand U9991 (N_9991,N_9096,N_9268);
and U9992 (N_9992,N_9392,N_9346);
or U9993 (N_9993,N_9282,N_9006);
nand U9994 (N_9994,N_9154,N_9429);
and U9995 (N_9995,N_9297,N_9464);
nand U9996 (N_9996,N_9374,N_9496);
or U9997 (N_9997,N_9327,N_9140);
and U9998 (N_9998,N_9095,N_9124);
or U9999 (N_9999,N_9165,N_9464);
xnor U10000 (N_10000,N_9767,N_9905);
nor U10001 (N_10001,N_9506,N_9898);
or U10002 (N_10002,N_9927,N_9581);
nor U10003 (N_10003,N_9802,N_9566);
nand U10004 (N_10004,N_9979,N_9827);
and U10005 (N_10005,N_9607,N_9633);
nor U10006 (N_10006,N_9663,N_9504);
or U10007 (N_10007,N_9840,N_9712);
xnor U10008 (N_10008,N_9550,N_9542);
xor U10009 (N_10009,N_9588,N_9511);
or U10010 (N_10010,N_9935,N_9518);
and U10011 (N_10011,N_9931,N_9502);
or U10012 (N_10012,N_9619,N_9692);
nor U10013 (N_10013,N_9531,N_9590);
or U10014 (N_10014,N_9519,N_9780);
xor U10015 (N_10015,N_9822,N_9574);
xnor U10016 (N_10016,N_9717,N_9760);
or U10017 (N_10017,N_9592,N_9571);
and U10018 (N_10018,N_9996,N_9688);
nor U10019 (N_10019,N_9682,N_9989);
xor U10020 (N_10020,N_9917,N_9834);
nor U10021 (N_10021,N_9555,N_9553);
nor U10022 (N_10022,N_9899,N_9730);
and U10023 (N_10023,N_9573,N_9598);
nand U10024 (N_10024,N_9861,N_9686);
or U10025 (N_10025,N_9932,N_9572);
xnor U10026 (N_10026,N_9984,N_9784);
nand U10027 (N_10027,N_9738,N_9943);
and U10028 (N_10028,N_9835,N_9874);
xnor U10029 (N_10029,N_9746,N_9737);
nand U10030 (N_10030,N_9850,N_9774);
nor U10031 (N_10031,N_9761,N_9889);
or U10032 (N_10032,N_9911,N_9726);
nand U10033 (N_10033,N_9602,N_9657);
xor U10034 (N_10034,N_9525,N_9678);
nand U10035 (N_10035,N_9757,N_9806);
nor U10036 (N_10036,N_9941,N_9515);
or U10037 (N_10037,N_9665,N_9677);
nand U10038 (N_10038,N_9593,N_9788);
or U10039 (N_10039,N_9936,N_9548);
nor U10040 (N_10040,N_9981,N_9801);
xor U10041 (N_10041,N_9512,N_9980);
xnor U10042 (N_10042,N_9945,N_9513);
or U10043 (N_10043,N_9960,N_9683);
and U10044 (N_10044,N_9810,N_9994);
nor U10045 (N_10045,N_9972,N_9596);
and U10046 (N_10046,N_9918,N_9603);
nor U10047 (N_10047,N_9839,N_9636);
nor U10048 (N_10048,N_9564,N_9676);
or U10049 (N_10049,N_9896,N_9953);
xnor U10050 (N_10050,N_9570,N_9690);
and U10051 (N_10051,N_9854,N_9614);
or U10052 (N_10052,N_9700,N_9956);
or U10053 (N_10053,N_9949,N_9915);
xnor U10054 (N_10054,N_9904,N_9794);
and U10055 (N_10055,N_9939,N_9582);
nor U10056 (N_10056,N_9803,N_9567);
xnor U10057 (N_10057,N_9991,N_9797);
xnor U10058 (N_10058,N_9993,N_9514);
or U10059 (N_10059,N_9799,N_9894);
or U10060 (N_10060,N_9705,N_9733);
nor U10061 (N_10061,N_9618,N_9679);
nor U10062 (N_10062,N_9990,N_9948);
and U10063 (N_10063,N_9983,N_9819);
and U10064 (N_10064,N_9946,N_9569);
or U10065 (N_10065,N_9630,N_9615);
or U10066 (N_10066,N_9675,N_9786);
xnor U10067 (N_10067,N_9754,N_9658);
nand U10068 (N_10068,N_9897,N_9649);
nand U10069 (N_10069,N_9696,N_9589);
or U10070 (N_10070,N_9651,N_9547);
nor U10071 (N_10071,N_9597,N_9887);
xor U10072 (N_10072,N_9851,N_9743);
and U10073 (N_10073,N_9858,N_9622);
and U10074 (N_10074,N_9527,N_9882);
nor U10075 (N_10075,N_9620,N_9558);
xor U10076 (N_10076,N_9735,N_9976);
nand U10077 (N_10077,N_9758,N_9562);
xnor U10078 (N_10078,N_9585,N_9866);
or U10079 (N_10079,N_9540,N_9968);
nand U10080 (N_10080,N_9765,N_9561);
xor U10081 (N_10081,N_9845,N_9812);
xnor U10082 (N_10082,N_9950,N_9557);
nand U10083 (N_10083,N_9500,N_9975);
xnor U10084 (N_10084,N_9681,N_9734);
and U10085 (N_10085,N_9910,N_9568);
xor U10086 (N_10086,N_9709,N_9702);
nor U10087 (N_10087,N_9711,N_9701);
nand U10088 (N_10088,N_9727,N_9785);
and U10089 (N_10089,N_9503,N_9997);
nor U10090 (N_10090,N_9906,N_9901);
nand U10091 (N_10091,N_9719,N_9775);
xnor U10092 (N_10092,N_9923,N_9594);
xor U10093 (N_10093,N_9601,N_9672);
nor U10094 (N_10094,N_9963,N_9852);
and U10095 (N_10095,N_9565,N_9832);
xnor U10096 (N_10096,N_9947,N_9877);
nand U10097 (N_10097,N_9753,N_9778);
nor U10098 (N_10098,N_9862,N_9546);
or U10099 (N_10099,N_9773,N_9655);
and U10100 (N_10100,N_9684,N_9560);
xor U10101 (N_10101,N_9621,N_9584);
nand U10102 (N_10102,N_9699,N_9772);
nor U10103 (N_10103,N_9508,N_9982);
xnor U10104 (N_10104,N_9969,N_9604);
or U10105 (N_10105,N_9965,N_9795);
nor U10106 (N_10106,N_9608,N_9638);
xor U10107 (N_10107,N_9961,N_9731);
or U10108 (N_10108,N_9755,N_9591);
xor U10109 (N_10109,N_9954,N_9748);
or U10110 (N_10110,N_9776,N_9647);
nor U10111 (N_10111,N_9974,N_9576);
xnor U10112 (N_10112,N_9516,N_9792);
nand U10113 (N_10113,N_9800,N_9973);
nor U10114 (N_10114,N_9600,N_9713);
and U10115 (N_10115,N_9654,N_9742);
xnor U10116 (N_10116,N_9929,N_9707);
nor U10117 (N_10117,N_9507,N_9648);
or U10118 (N_10118,N_9818,N_9855);
nor U10119 (N_10119,N_9763,N_9859);
nand U10120 (N_10120,N_9706,N_9768);
nand U10121 (N_10121,N_9575,N_9787);
xor U10122 (N_10122,N_9611,N_9517);
and U10123 (N_10123,N_9632,N_9875);
nand U10124 (N_10124,N_9934,N_9728);
nor U10125 (N_10125,N_9885,N_9613);
or U10126 (N_10126,N_9667,N_9970);
or U10127 (N_10127,N_9830,N_9928);
nor U10128 (N_10128,N_9791,N_9641);
or U10129 (N_10129,N_9554,N_9781);
nand U10130 (N_10130,N_9739,N_9530);
and U10131 (N_10131,N_9745,N_9916);
nand U10132 (N_10132,N_9634,N_9646);
nor U10133 (N_10133,N_9868,N_9798);
and U10134 (N_10134,N_9964,N_9978);
nor U10135 (N_10135,N_9908,N_9749);
xnor U10136 (N_10136,N_9853,N_9955);
nand U10137 (N_10137,N_9520,N_9535);
and U10138 (N_10138,N_9999,N_9938);
and U10139 (N_10139,N_9987,N_9741);
nand U10140 (N_10140,N_9668,N_9942);
and U10141 (N_10141,N_9782,N_9586);
or U10142 (N_10142,N_9559,N_9544);
nand U10143 (N_10143,N_9771,N_9626);
nand U10144 (N_10144,N_9966,N_9878);
or U10145 (N_10145,N_9808,N_9766);
nor U10146 (N_10146,N_9959,N_9902);
nand U10147 (N_10147,N_9770,N_9642);
nor U10148 (N_10148,N_9521,N_9933);
xnor U10149 (N_10149,N_9724,N_9876);
and U10150 (N_10150,N_9789,N_9624);
or U10151 (N_10151,N_9809,N_9533);
and U10152 (N_10152,N_9595,N_9645);
xor U10153 (N_10153,N_9666,N_9714);
and U10154 (N_10154,N_9698,N_9725);
xor U10155 (N_10155,N_9631,N_9528);
and U10156 (N_10156,N_9612,N_9556);
or U10157 (N_10157,N_9879,N_9670);
and U10158 (N_10158,N_9545,N_9831);
or U10159 (N_10159,N_9524,N_9815);
nor U10160 (N_10160,N_9930,N_9659);
or U10161 (N_10161,N_9814,N_9995);
or U10162 (N_10162,N_9888,N_9577);
or U10163 (N_10163,N_9828,N_9580);
xnor U10164 (N_10164,N_9920,N_9844);
and U10165 (N_10165,N_9764,N_9625);
and U10166 (N_10166,N_9536,N_9762);
xnor U10167 (N_10167,N_9992,N_9922);
nand U10168 (N_10168,N_9985,N_9836);
xnor U10169 (N_10169,N_9541,N_9660);
nand U10170 (N_10170,N_9680,N_9671);
xnor U10171 (N_10171,N_9805,N_9986);
xnor U10172 (N_10172,N_9957,N_9715);
xnor U10173 (N_10173,N_9579,N_9509);
xor U10174 (N_10174,N_9813,N_9708);
or U10175 (N_10175,N_9744,N_9843);
nand U10176 (N_10176,N_9804,N_9796);
xnor U10177 (N_10177,N_9824,N_9951);
nor U10178 (N_10178,N_9759,N_9691);
and U10179 (N_10179,N_9944,N_9820);
or U10180 (N_10180,N_9609,N_9740);
xnor U10181 (N_10181,N_9895,N_9873);
and U10182 (N_10182,N_9842,N_9605);
or U10183 (N_10183,N_9529,N_9883);
nand U10184 (N_10184,N_9871,N_9998);
or U10185 (N_10185,N_9643,N_9661);
nor U10186 (N_10186,N_9913,N_9687);
nor U10187 (N_10187,N_9886,N_9937);
and U10188 (N_10188,N_9881,N_9685);
and U10189 (N_10189,N_9644,N_9736);
and U10190 (N_10190,N_9756,N_9870);
and U10191 (N_10191,N_9751,N_9669);
and U10192 (N_10192,N_9829,N_9848);
nor U10193 (N_10193,N_9697,N_9903);
nor U10194 (N_10194,N_9539,N_9940);
xnor U10195 (N_10195,N_9958,N_9718);
or U10196 (N_10196,N_9599,N_9857);
nand U10197 (N_10197,N_9720,N_9869);
nor U10198 (N_10198,N_9716,N_9526);
and U10199 (N_10199,N_9837,N_9732);
or U10200 (N_10200,N_9807,N_9721);
nor U10201 (N_10201,N_9900,N_9532);
and U10202 (N_10202,N_9865,N_9926);
xnor U10203 (N_10203,N_9750,N_9793);
nor U10204 (N_10204,N_9892,N_9921);
or U10205 (N_10205,N_9838,N_9616);
and U10206 (N_10206,N_9673,N_9747);
xor U10207 (N_10207,N_9628,N_9790);
xnor U10208 (N_10208,N_9823,N_9884);
nand U10209 (N_10209,N_9971,N_9637);
or U10210 (N_10210,N_9629,N_9872);
or U10211 (N_10211,N_9543,N_9695);
nand U10212 (N_10212,N_9549,N_9816);
nor U10213 (N_10213,N_9825,N_9640);
nor U10214 (N_10214,N_9962,N_9523);
or U10215 (N_10215,N_9639,N_9811);
or U10216 (N_10216,N_9891,N_9587);
xnor U10217 (N_10217,N_9967,N_9583);
or U10218 (N_10218,N_9729,N_9779);
nand U10219 (N_10219,N_9777,N_9893);
nor U10220 (N_10220,N_9914,N_9826);
or U10221 (N_10221,N_9849,N_9610);
nor U10222 (N_10222,N_9864,N_9909);
nor U10223 (N_10223,N_9925,N_9578);
nor U10224 (N_10224,N_9988,N_9769);
nand U10225 (N_10225,N_9912,N_9856);
or U10226 (N_10226,N_9635,N_9689);
nor U10227 (N_10227,N_9924,N_9723);
or U10228 (N_10228,N_9821,N_9551);
or U10229 (N_10229,N_9722,N_9847);
nand U10230 (N_10230,N_9652,N_9977);
or U10231 (N_10231,N_9606,N_9522);
and U10232 (N_10232,N_9505,N_9538);
nand U10233 (N_10233,N_9662,N_9694);
and U10234 (N_10234,N_9907,N_9674);
xnor U10235 (N_10235,N_9563,N_9693);
nor U10236 (N_10236,N_9919,N_9783);
or U10237 (N_10237,N_9703,N_9656);
or U10238 (N_10238,N_9890,N_9880);
nor U10239 (N_10239,N_9846,N_9817);
and U10240 (N_10240,N_9552,N_9841);
nor U10241 (N_10241,N_9510,N_9860);
or U10242 (N_10242,N_9627,N_9537);
nor U10243 (N_10243,N_9833,N_9617);
and U10244 (N_10244,N_9653,N_9952);
or U10245 (N_10245,N_9534,N_9867);
nand U10246 (N_10246,N_9704,N_9710);
and U10247 (N_10247,N_9623,N_9664);
nor U10248 (N_10248,N_9650,N_9752);
nor U10249 (N_10249,N_9501,N_9863);
and U10250 (N_10250,N_9516,N_9915);
xnor U10251 (N_10251,N_9642,N_9605);
and U10252 (N_10252,N_9799,N_9638);
nor U10253 (N_10253,N_9894,N_9707);
nand U10254 (N_10254,N_9600,N_9867);
xnor U10255 (N_10255,N_9816,N_9680);
or U10256 (N_10256,N_9810,N_9763);
nor U10257 (N_10257,N_9721,N_9970);
xnor U10258 (N_10258,N_9953,N_9598);
and U10259 (N_10259,N_9668,N_9723);
or U10260 (N_10260,N_9716,N_9899);
xnor U10261 (N_10261,N_9949,N_9982);
xnor U10262 (N_10262,N_9797,N_9660);
nand U10263 (N_10263,N_9956,N_9842);
nand U10264 (N_10264,N_9778,N_9806);
or U10265 (N_10265,N_9927,N_9521);
or U10266 (N_10266,N_9558,N_9598);
xnor U10267 (N_10267,N_9876,N_9536);
or U10268 (N_10268,N_9683,N_9577);
nand U10269 (N_10269,N_9991,N_9929);
nor U10270 (N_10270,N_9843,N_9830);
and U10271 (N_10271,N_9851,N_9618);
and U10272 (N_10272,N_9659,N_9933);
xnor U10273 (N_10273,N_9966,N_9872);
or U10274 (N_10274,N_9662,N_9921);
nor U10275 (N_10275,N_9896,N_9680);
or U10276 (N_10276,N_9974,N_9536);
nor U10277 (N_10277,N_9874,N_9763);
xnor U10278 (N_10278,N_9666,N_9841);
xnor U10279 (N_10279,N_9590,N_9611);
nand U10280 (N_10280,N_9941,N_9550);
nand U10281 (N_10281,N_9985,N_9637);
nor U10282 (N_10282,N_9638,N_9556);
or U10283 (N_10283,N_9951,N_9976);
nor U10284 (N_10284,N_9669,N_9719);
nor U10285 (N_10285,N_9813,N_9973);
nor U10286 (N_10286,N_9508,N_9530);
or U10287 (N_10287,N_9904,N_9959);
nor U10288 (N_10288,N_9508,N_9640);
and U10289 (N_10289,N_9504,N_9649);
or U10290 (N_10290,N_9988,N_9971);
or U10291 (N_10291,N_9993,N_9903);
nand U10292 (N_10292,N_9787,N_9723);
nand U10293 (N_10293,N_9735,N_9822);
or U10294 (N_10294,N_9678,N_9777);
or U10295 (N_10295,N_9849,N_9507);
xor U10296 (N_10296,N_9734,N_9706);
nand U10297 (N_10297,N_9977,N_9584);
and U10298 (N_10298,N_9609,N_9543);
nand U10299 (N_10299,N_9731,N_9529);
xnor U10300 (N_10300,N_9846,N_9621);
nand U10301 (N_10301,N_9505,N_9765);
or U10302 (N_10302,N_9853,N_9826);
nand U10303 (N_10303,N_9849,N_9504);
nand U10304 (N_10304,N_9776,N_9807);
and U10305 (N_10305,N_9976,N_9638);
nand U10306 (N_10306,N_9853,N_9666);
nand U10307 (N_10307,N_9815,N_9910);
nor U10308 (N_10308,N_9950,N_9926);
or U10309 (N_10309,N_9927,N_9619);
or U10310 (N_10310,N_9669,N_9960);
nor U10311 (N_10311,N_9675,N_9848);
xnor U10312 (N_10312,N_9974,N_9879);
xor U10313 (N_10313,N_9721,N_9615);
and U10314 (N_10314,N_9997,N_9908);
and U10315 (N_10315,N_9600,N_9800);
nand U10316 (N_10316,N_9716,N_9507);
or U10317 (N_10317,N_9909,N_9960);
nor U10318 (N_10318,N_9928,N_9724);
and U10319 (N_10319,N_9907,N_9643);
xnor U10320 (N_10320,N_9549,N_9809);
and U10321 (N_10321,N_9721,N_9923);
xnor U10322 (N_10322,N_9593,N_9750);
nor U10323 (N_10323,N_9740,N_9877);
xor U10324 (N_10324,N_9547,N_9701);
xor U10325 (N_10325,N_9552,N_9788);
or U10326 (N_10326,N_9708,N_9526);
and U10327 (N_10327,N_9961,N_9856);
xor U10328 (N_10328,N_9683,N_9938);
and U10329 (N_10329,N_9651,N_9536);
nor U10330 (N_10330,N_9599,N_9938);
xnor U10331 (N_10331,N_9957,N_9742);
nor U10332 (N_10332,N_9974,N_9901);
xnor U10333 (N_10333,N_9689,N_9535);
xor U10334 (N_10334,N_9834,N_9862);
nor U10335 (N_10335,N_9975,N_9572);
xnor U10336 (N_10336,N_9811,N_9582);
xnor U10337 (N_10337,N_9709,N_9975);
xor U10338 (N_10338,N_9975,N_9874);
and U10339 (N_10339,N_9726,N_9861);
xnor U10340 (N_10340,N_9624,N_9865);
nor U10341 (N_10341,N_9675,N_9719);
nor U10342 (N_10342,N_9887,N_9973);
and U10343 (N_10343,N_9575,N_9574);
xor U10344 (N_10344,N_9581,N_9654);
or U10345 (N_10345,N_9545,N_9818);
and U10346 (N_10346,N_9850,N_9531);
nor U10347 (N_10347,N_9542,N_9657);
xnor U10348 (N_10348,N_9774,N_9712);
nor U10349 (N_10349,N_9750,N_9761);
xnor U10350 (N_10350,N_9819,N_9765);
nor U10351 (N_10351,N_9731,N_9989);
and U10352 (N_10352,N_9786,N_9999);
or U10353 (N_10353,N_9701,N_9709);
and U10354 (N_10354,N_9558,N_9870);
and U10355 (N_10355,N_9518,N_9719);
or U10356 (N_10356,N_9508,N_9867);
nor U10357 (N_10357,N_9639,N_9834);
and U10358 (N_10358,N_9556,N_9928);
and U10359 (N_10359,N_9500,N_9827);
xnor U10360 (N_10360,N_9990,N_9935);
nor U10361 (N_10361,N_9550,N_9834);
and U10362 (N_10362,N_9990,N_9844);
and U10363 (N_10363,N_9748,N_9562);
or U10364 (N_10364,N_9631,N_9780);
or U10365 (N_10365,N_9928,N_9923);
nor U10366 (N_10366,N_9710,N_9974);
and U10367 (N_10367,N_9683,N_9832);
nor U10368 (N_10368,N_9807,N_9508);
xor U10369 (N_10369,N_9903,N_9686);
nand U10370 (N_10370,N_9692,N_9902);
xor U10371 (N_10371,N_9866,N_9677);
or U10372 (N_10372,N_9768,N_9761);
nand U10373 (N_10373,N_9631,N_9729);
nand U10374 (N_10374,N_9517,N_9865);
xor U10375 (N_10375,N_9647,N_9649);
or U10376 (N_10376,N_9756,N_9839);
or U10377 (N_10377,N_9900,N_9851);
and U10378 (N_10378,N_9594,N_9992);
nand U10379 (N_10379,N_9718,N_9552);
and U10380 (N_10380,N_9908,N_9611);
nor U10381 (N_10381,N_9547,N_9676);
nand U10382 (N_10382,N_9510,N_9802);
and U10383 (N_10383,N_9611,N_9975);
nor U10384 (N_10384,N_9558,N_9903);
xnor U10385 (N_10385,N_9618,N_9778);
nand U10386 (N_10386,N_9887,N_9844);
nor U10387 (N_10387,N_9767,N_9596);
xor U10388 (N_10388,N_9941,N_9759);
or U10389 (N_10389,N_9855,N_9822);
and U10390 (N_10390,N_9854,N_9790);
nor U10391 (N_10391,N_9788,N_9531);
or U10392 (N_10392,N_9867,N_9516);
or U10393 (N_10393,N_9552,N_9742);
and U10394 (N_10394,N_9738,N_9576);
nor U10395 (N_10395,N_9668,N_9837);
nor U10396 (N_10396,N_9749,N_9851);
or U10397 (N_10397,N_9908,N_9861);
xnor U10398 (N_10398,N_9769,N_9857);
nor U10399 (N_10399,N_9886,N_9673);
xnor U10400 (N_10400,N_9537,N_9641);
nand U10401 (N_10401,N_9718,N_9768);
or U10402 (N_10402,N_9651,N_9514);
and U10403 (N_10403,N_9824,N_9511);
nand U10404 (N_10404,N_9990,N_9795);
xnor U10405 (N_10405,N_9778,N_9719);
nor U10406 (N_10406,N_9979,N_9926);
or U10407 (N_10407,N_9972,N_9529);
and U10408 (N_10408,N_9554,N_9885);
and U10409 (N_10409,N_9788,N_9872);
and U10410 (N_10410,N_9694,N_9908);
xor U10411 (N_10411,N_9834,N_9676);
and U10412 (N_10412,N_9768,N_9545);
and U10413 (N_10413,N_9711,N_9770);
or U10414 (N_10414,N_9680,N_9881);
and U10415 (N_10415,N_9837,N_9722);
nor U10416 (N_10416,N_9805,N_9575);
nor U10417 (N_10417,N_9608,N_9814);
nand U10418 (N_10418,N_9635,N_9704);
nand U10419 (N_10419,N_9789,N_9785);
nor U10420 (N_10420,N_9756,N_9824);
xnor U10421 (N_10421,N_9535,N_9872);
or U10422 (N_10422,N_9644,N_9621);
and U10423 (N_10423,N_9901,N_9776);
and U10424 (N_10424,N_9545,N_9651);
xnor U10425 (N_10425,N_9776,N_9989);
nor U10426 (N_10426,N_9856,N_9703);
xnor U10427 (N_10427,N_9915,N_9722);
or U10428 (N_10428,N_9712,N_9683);
and U10429 (N_10429,N_9912,N_9970);
nor U10430 (N_10430,N_9786,N_9692);
and U10431 (N_10431,N_9815,N_9658);
and U10432 (N_10432,N_9548,N_9600);
nand U10433 (N_10433,N_9520,N_9511);
or U10434 (N_10434,N_9811,N_9677);
xor U10435 (N_10435,N_9507,N_9944);
nor U10436 (N_10436,N_9506,N_9836);
or U10437 (N_10437,N_9548,N_9509);
and U10438 (N_10438,N_9793,N_9659);
nor U10439 (N_10439,N_9611,N_9764);
nand U10440 (N_10440,N_9981,N_9525);
xnor U10441 (N_10441,N_9897,N_9629);
or U10442 (N_10442,N_9529,N_9780);
nor U10443 (N_10443,N_9955,N_9766);
and U10444 (N_10444,N_9566,N_9975);
nand U10445 (N_10445,N_9823,N_9982);
nor U10446 (N_10446,N_9993,N_9609);
xnor U10447 (N_10447,N_9748,N_9600);
nor U10448 (N_10448,N_9915,N_9654);
or U10449 (N_10449,N_9743,N_9760);
nand U10450 (N_10450,N_9699,N_9804);
xor U10451 (N_10451,N_9639,N_9816);
nor U10452 (N_10452,N_9675,N_9711);
xor U10453 (N_10453,N_9715,N_9629);
nor U10454 (N_10454,N_9799,N_9607);
nand U10455 (N_10455,N_9850,N_9890);
and U10456 (N_10456,N_9888,N_9644);
and U10457 (N_10457,N_9720,N_9641);
nand U10458 (N_10458,N_9736,N_9627);
xnor U10459 (N_10459,N_9843,N_9867);
nand U10460 (N_10460,N_9603,N_9884);
or U10461 (N_10461,N_9952,N_9573);
nand U10462 (N_10462,N_9811,N_9750);
and U10463 (N_10463,N_9557,N_9578);
or U10464 (N_10464,N_9973,N_9976);
and U10465 (N_10465,N_9845,N_9925);
nor U10466 (N_10466,N_9987,N_9830);
and U10467 (N_10467,N_9781,N_9716);
and U10468 (N_10468,N_9742,N_9735);
and U10469 (N_10469,N_9675,N_9659);
nand U10470 (N_10470,N_9621,N_9997);
nor U10471 (N_10471,N_9674,N_9934);
nor U10472 (N_10472,N_9916,N_9822);
xnor U10473 (N_10473,N_9941,N_9920);
and U10474 (N_10474,N_9752,N_9854);
nor U10475 (N_10475,N_9697,N_9651);
and U10476 (N_10476,N_9638,N_9796);
nor U10477 (N_10477,N_9897,N_9827);
nand U10478 (N_10478,N_9603,N_9695);
and U10479 (N_10479,N_9982,N_9680);
and U10480 (N_10480,N_9929,N_9744);
xor U10481 (N_10481,N_9669,N_9708);
xnor U10482 (N_10482,N_9555,N_9558);
and U10483 (N_10483,N_9819,N_9661);
or U10484 (N_10484,N_9774,N_9990);
nor U10485 (N_10485,N_9617,N_9524);
nor U10486 (N_10486,N_9958,N_9957);
nor U10487 (N_10487,N_9724,N_9912);
nand U10488 (N_10488,N_9970,N_9641);
xnor U10489 (N_10489,N_9877,N_9849);
nor U10490 (N_10490,N_9908,N_9682);
xor U10491 (N_10491,N_9558,N_9979);
nand U10492 (N_10492,N_9942,N_9610);
or U10493 (N_10493,N_9845,N_9612);
or U10494 (N_10494,N_9823,N_9562);
nand U10495 (N_10495,N_9786,N_9711);
or U10496 (N_10496,N_9832,N_9980);
and U10497 (N_10497,N_9867,N_9656);
nor U10498 (N_10498,N_9819,N_9868);
xnor U10499 (N_10499,N_9986,N_9943);
xor U10500 (N_10500,N_10319,N_10382);
or U10501 (N_10501,N_10356,N_10196);
or U10502 (N_10502,N_10467,N_10413);
and U10503 (N_10503,N_10214,N_10227);
and U10504 (N_10504,N_10412,N_10101);
nor U10505 (N_10505,N_10357,N_10417);
or U10506 (N_10506,N_10171,N_10405);
nand U10507 (N_10507,N_10085,N_10267);
xor U10508 (N_10508,N_10261,N_10194);
or U10509 (N_10509,N_10291,N_10240);
and U10510 (N_10510,N_10139,N_10201);
nor U10511 (N_10511,N_10480,N_10030);
or U10512 (N_10512,N_10179,N_10266);
or U10513 (N_10513,N_10048,N_10205);
or U10514 (N_10514,N_10178,N_10019);
nor U10515 (N_10515,N_10228,N_10292);
nand U10516 (N_10516,N_10286,N_10122);
xnor U10517 (N_10517,N_10089,N_10452);
nand U10518 (N_10518,N_10071,N_10077);
xor U10519 (N_10519,N_10470,N_10114);
xnor U10520 (N_10520,N_10409,N_10220);
xor U10521 (N_10521,N_10133,N_10198);
or U10522 (N_10522,N_10144,N_10116);
nor U10523 (N_10523,N_10431,N_10396);
nand U10524 (N_10524,N_10485,N_10410);
and U10525 (N_10525,N_10005,N_10164);
nor U10526 (N_10526,N_10065,N_10421);
and U10527 (N_10527,N_10060,N_10173);
or U10528 (N_10528,N_10394,N_10426);
or U10529 (N_10529,N_10035,N_10464);
or U10530 (N_10530,N_10370,N_10152);
nand U10531 (N_10531,N_10165,N_10104);
xnor U10532 (N_10532,N_10009,N_10036);
and U10533 (N_10533,N_10108,N_10314);
nor U10534 (N_10534,N_10224,N_10031);
nand U10535 (N_10535,N_10306,N_10444);
or U10536 (N_10536,N_10262,N_10100);
nor U10537 (N_10537,N_10202,N_10454);
or U10538 (N_10538,N_10492,N_10251);
and U10539 (N_10539,N_10182,N_10203);
and U10540 (N_10540,N_10424,N_10168);
nand U10541 (N_10541,N_10238,N_10024);
or U10542 (N_10542,N_10316,N_10148);
nor U10543 (N_10543,N_10127,N_10057);
and U10544 (N_10544,N_10347,N_10318);
or U10545 (N_10545,N_10377,N_10327);
or U10546 (N_10546,N_10226,N_10125);
nand U10547 (N_10547,N_10283,N_10337);
and U10548 (N_10548,N_10369,N_10481);
xnor U10549 (N_10549,N_10406,N_10279);
nor U10550 (N_10550,N_10325,N_10047);
nor U10551 (N_10551,N_10234,N_10372);
xnor U10552 (N_10552,N_10193,N_10263);
and U10553 (N_10553,N_10128,N_10425);
nor U10554 (N_10554,N_10358,N_10380);
nand U10555 (N_10555,N_10308,N_10155);
or U10556 (N_10556,N_10187,N_10335);
nor U10557 (N_10557,N_10004,N_10298);
nand U10558 (N_10558,N_10333,N_10320);
or U10559 (N_10559,N_10363,N_10430);
or U10560 (N_10560,N_10177,N_10373);
and U10561 (N_10561,N_10175,N_10222);
xnor U10562 (N_10562,N_10264,N_10072);
and U10563 (N_10563,N_10456,N_10008);
and U10564 (N_10564,N_10475,N_10123);
nand U10565 (N_10565,N_10053,N_10375);
nor U10566 (N_10566,N_10084,N_10029);
xor U10567 (N_10567,N_10058,N_10180);
or U10568 (N_10568,N_10388,N_10096);
nand U10569 (N_10569,N_10317,N_10403);
nand U10570 (N_10570,N_10346,N_10176);
and U10571 (N_10571,N_10290,N_10359);
nand U10572 (N_10572,N_10055,N_10387);
and U10573 (N_10573,N_10381,N_10239);
or U10574 (N_10574,N_10184,N_10093);
and U10575 (N_10575,N_10307,N_10069);
nor U10576 (N_10576,N_10212,N_10415);
nand U10577 (N_10577,N_10115,N_10254);
or U10578 (N_10578,N_10229,N_10206);
or U10579 (N_10579,N_10451,N_10132);
or U10580 (N_10580,N_10362,N_10259);
or U10581 (N_10581,N_10003,N_10199);
xor U10582 (N_10582,N_10231,N_10097);
nand U10583 (N_10583,N_10106,N_10256);
nor U10584 (N_10584,N_10404,N_10107);
nand U10585 (N_10585,N_10001,N_10443);
xor U10586 (N_10586,N_10477,N_10138);
nand U10587 (N_10587,N_10277,N_10192);
xor U10588 (N_10588,N_10195,N_10383);
or U10589 (N_10589,N_10275,N_10462);
or U10590 (N_10590,N_10401,N_10384);
and U10591 (N_10591,N_10488,N_10293);
or U10592 (N_10592,N_10305,N_10159);
nor U10593 (N_10593,N_10191,N_10343);
xor U10594 (N_10594,N_10252,N_10258);
or U10595 (N_10595,N_10341,N_10310);
xnor U10596 (N_10596,N_10437,N_10073);
or U10597 (N_10597,N_10109,N_10368);
or U10598 (N_10598,N_10336,N_10121);
nor U10599 (N_10599,N_10197,N_10010);
nor U10600 (N_10600,N_10459,N_10445);
or U10601 (N_10601,N_10338,N_10245);
or U10602 (N_10602,N_10329,N_10423);
nor U10603 (N_10603,N_10129,N_10389);
xnor U10604 (N_10604,N_10386,N_10011);
xnor U10605 (N_10605,N_10402,N_10130);
nor U10606 (N_10606,N_10257,N_10235);
xnor U10607 (N_10607,N_10304,N_10416);
or U10608 (N_10608,N_10294,N_10021);
nor U10609 (N_10609,N_10281,N_10427);
or U10610 (N_10610,N_10455,N_10006);
nor U10611 (N_10611,N_10350,N_10041);
nand U10612 (N_10612,N_10268,N_10418);
xor U10613 (N_10613,N_10040,N_10156);
xor U10614 (N_10614,N_10490,N_10142);
xnor U10615 (N_10615,N_10150,N_10349);
or U10616 (N_10616,N_10099,N_10473);
and U10617 (N_10617,N_10033,N_10140);
xnor U10618 (N_10618,N_10483,N_10478);
or U10619 (N_10619,N_10207,N_10117);
nand U10620 (N_10620,N_10113,N_10265);
and U10621 (N_10621,N_10393,N_10295);
or U10622 (N_10622,N_10246,N_10126);
xor U10623 (N_10623,N_10322,N_10045);
or U10624 (N_10624,N_10059,N_10225);
nand U10625 (N_10625,N_10050,N_10078);
xor U10626 (N_10626,N_10398,N_10284);
nor U10627 (N_10627,N_10061,N_10015);
and U10628 (N_10628,N_10174,N_10355);
xor U10629 (N_10629,N_10432,N_10374);
nor U10630 (N_10630,N_10280,N_10463);
nor U10631 (N_10631,N_10181,N_10494);
nor U10632 (N_10632,N_10124,N_10450);
or U10633 (N_10633,N_10497,N_10166);
nand U10634 (N_10634,N_10303,N_10052);
nand U10635 (N_10635,N_10399,N_10002);
xor U10636 (N_10636,N_10141,N_10103);
xnor U10637 (N_10637,N_10169,N_10371);
and U10638 (N_10638,N_10302,N_10479);
or U10639 (N_10639,N_10083,N_10422);
and U10640 (N_10640,N_10162,N_10330);
or U10641 (N_10641,N_10419,N_10120);
nor U10642 (N_10642,N_10081,N_10051);
nor U10643 (N_10643,N_10149,N_10056);
xnor U10644 (N_10644,N_10301,N_10157);
or U10645 (N_10645,N_10154,N_10495);
nor U10646 (N_10646,N_10408,N_10074);
or U10647 (N_10647,N_10365,N_10119);
nor U10648 (N_10648,N_10012,N_10210);
nor U10649 (N_10649,N_10461,N_10082);
nor U10650 (N_10650,N_10038,N_10020);
nand U10651 (N_10651,N_10208,N_10441);
xnor U10652 (N_10652,N_10062,N_10339);
nor U10653 (N_10653,N_10344,N_10269);
nand U10654 (N_10654,N_10489,N_10086);
and U10655 (N_10655,N_10498,N_10376);
or U10656 (N_10656,N_10049,N_10230);
nor U10657 (N_10657,N_10270,N_10324);
xor U10658 (N_10658,N_10447,N_10237);
and U10659 (N_10659,N_10025,N_10438);
and U10660 (N_10660,N_10364,N_10367);
nor U10661 (N_10661,N_10032,N_10278);
nor U10662 (N_10662,N_10158,N_10215);
nor U10663 (N_10663,N_10044,N_10209);
and U10664 (N_10664,N_10378,N_10146);
and U10665 (N_10665,N_10167,N_10385);
nand U10666 (N_10666,N_10249,N_10297);
xor U10667 (N_10667,N_10068,N_10448);
nand U10668 (N_10668,N_10242,N_10458);
nor U10669 (N_10669,N_10110,N_10190);
and U10670 (N_10670,N_10250,N_10326);
and U10671 (N_10671,N_10247,N_10486);
nand U10672 (N_10672,N_10241,N_10135);
nor U10673 (N_10673,N_10137,N_10037);
xnor U10674 (N_10674,N_10186,N_10145);
and U10675 (N_10675,N_10027,N_10070);
nand U10676 (N_10676,N_10172,N_10407);
and U10677 (N_10677,N_10469,N_10414);
or U10678 (N_10678,N_10018,N_10102);
xor U10679 (N_10679,N_10274,N_10026);
and U10680 (N_10680,N_10300,N_10457);
nor U10681 (N_10681,N_10439,N_10147);
xor U10682 (N_10682,N_10453,N_10233);
nor U10683 (N_10683,N_10088,N_10092);
nand U10684 (N_10684,N_10285,N_10446);
xnor U10685 (N_10685,N_10379,N_10465);
nand U10686 (N_10686,N_10312,N_10017);
xnor U10687 (N_10687,N_10309,N_10288);
xnor U10688 (N_10688,N_10323,N_10094);
xnor U10689 (N_10689,N_10034,N_10433);
and U10690 (N_10690,N_10223,N_10345);
or U10691 (N_10691,N_10066,N_10131);
and U10692 (N_10692,N_10232,N_10098);
or U10693 (N_10693,N_10436,N_10151);
xnor U10694 (N_10694,N_10442,N_10311);
nor U10695 (N_10695,N_10043,N_10468);
or U10696 (N_10696,N_10075,N_10022);
nor U10697 (N_10697,N_10315,N_10161);
xnor U10698 (N_10698,N_10218,N_10472);
and U10699 (N_10699,N_10067,N_10429);
nand U10700 (N_10700,N_10160,N_10491);
xnor U10701 (N_10701,N_10014,N_10090);
xnor U10702 (N_10702,N_10221,N_10360);
and U10703 (N_10703,N_10466,N_10200);
nand U10704 (N_10704,N_10342,N_10353);
nor U10705 (N_10705,N_10028,N_10007);
nor U10706 (N_10706,N_10428,N_10334);
and U10707 (N_10707,N_10328,N_10272);
or U10708 (N_10708,N_10105,N_10332);
or U10709 (N_10709,N_10042,N_10289);
or U10710 (N_10710,N_10248,N_10392);
or U10711 (N_10711,N_10016,N_10213);
nor U10712 (N_10712,N_10023,N_10493);
and U10713 (N_10713,N_10136,N_10087);
xnor U10714 (N_10714,N_10118,N_10366);
and U10715 (N_10715,N_10273,N_10091);
and U10716 (N_10716,N_10183,N_10313);
and U10717 (N_10717,N_10079,N_10204);
nand U10718 (N_10718,N_10276,N_10170);
xnor U10719 (N_10719,N_10143,N_10354);
and U10720 (N_10720,N_10244,N_10449);
nand U10721 (N_10721,N_10331,N_10063);
nor U10722 (N_10722,N_10189,N_10484);
nand U10723 (N_10723,N_10352,N_10395);
xor U10724 (N_10724,N_10271,N_10260);
or U10725 (N_10725,N_10080,N_10188);
nand U10726 (N_10726,N_10390,N_10216);
xor U10727 (N_10727,N_10219,N_10476);
and U10728 (N_10728,N_10471,N_10111);
xor U10729 (N_10729,N_10411,N_10361);
xor U10730 (N_10730,N_10013,N_10076);
nor U10731 (N_10731,N_10348,N_10420);
nor U10732 (N_10732,N_10435,N_10460);
nor U10733 (N_10733,N_10296,N_10112);
and U10734 (N_10734,N_10282,N_10217);
or U10735 (N_10735,N_10321,N_10440);
and U10736 (N_10736,N_10255,N_10287);
nor U10737 (N_10737,N_10474,N_10000);
and U10738 (N_10738,N_10397,N_10054);
nor U10739 (N_10739,N_10496,N_10351);
xnor U10740 (N_10740,N_10134,N_10064);
nand U10741 (N_10741,N_10434,N_10236);
nor U10742 (N_10742,N_10400,N_10163);
nand U10743 (N_10743,N_10299,N_10095);
nand U10744 (N_10744,N_10391,N_10153);
or U10745 (N_10745,N_10185,N_10482);
nor U10746 (N_10746,N_10253,N_10499);
or U10747 (N_10747,N_10211,N_10340);
or U10748 (N_10748,N_10046,N_10243);
or U10749 (N_10749,N_10039,N_10487);
nand U10750 (N_10750,N_10247,N_10371);
nor U10751 (N_10751,N_10387,N_10321);
nand U10752 (N_10752,N_10442,N_10294);
and U10753 (N_10753,N_10335,N_10398);
and U10754 (N_10754,N_10200,N_10436);
nor U10755 (N_10755,N_10340,N_10031);
xor U10756 (N_10756,N_10070,N_10471);
xnor U10757 (N_10757,N_10269,N_10395);
or U10758 (N_10758,N_10258,N_10173);
nand U10759 (N_10759,N_10428,N_10232);
nand U10760 (N_10760,N_10038,N_10149);
nor U10761 (N_10761,N_10389,N_10412);
xor U10762 (N_10762,N_10071,N_10496);
or U10763 (N_10763,N_10399,N_10454);
nor U10764 (N_10764,N_10391,N_10333);
xnor U10765 (N_10765,N_10149,N_10350);
nor U10766 (N_10766,N_10481,N_10056);
xnor U10767 (N_10767,N_10238,N_10284);
xor U10768 (N_10768,N_10242,N_10194);
xnor U10769 (N_10769,N_10356,N_10389);
nor U10770 (N_10770,N_10242,N_10259);
nand U10771 (N_10771,N_10171,N_10090);
or U10772 (N_10772,N_10390,N_10352);
nor U10773 (N_10773,N_10211,N_10016);
or U10774 (N_10774,N_10447,N_10066);
or U10775 (N_10775,N_10326,N_10447);
nand U10776 (N_10776,N_10404,N_10181);
xor U10777 (N_10777,N_10077,N_10210);
nand U10778 (N_10778,N_10343,N_10057);
nand U10779 (N_10779,N_10319,N_10263);
or U10780 (N_10780,N_10110,N_10070);
and U10781 (N_10781,N_10417,N_10372);
xnor U10782 (N_10782,N_10039,N_10412);
xnor U10783 (N_10783,N_10124,N_10461);
or U10784 (N_10784,N_10360,N_10127);
and U10785 (N_10785,N_10059,N_10181);
xor U10786 (N_10786,N_10437,N_10392);
nand U10787 (N_10787,N_10108,N_10036);
and U10788 (N_10788,N_10181,N_10453);
nand U10789 (N_10789,N_10463,N_10289);
and U10790 (N_10790,N_10300,N_10116);
and U10791 (N_10791,N_10345,N_10382);
and U10792 (N_10792,N_10070,N_10055);
nand U10793 (N_10793,N_10304,N_10017);
nor U10794 (N_10794,N_10441,N_10239);
nand U10795 (N_10795,N_10155,N_10257);
xor U10796 (N_10796,N_10090,N_10174);
or U10797 (N_10797,N_10396,N_10497);
or U10798 (N_10798,N_10381,N_10132);
or U10799 (N_10799,N_10435,N_10434);
nand U10800 (N_10800,N_10118,N_10386);
and U10801 (N_10801,N_10305,N_10027);
and U10802 (N_10802,N_10124,N_10055);
and U10803 (N_10803,N_10244,N_10404);
and U10804 (N_10804,N_10288,N_10277);
nor U10805 (N_10805,N_10263,N_10243);
nand U10806 (N_10806,N_10047,N_10233);
nor U10807 (N_10807,N_10268,N_10338);
xor U10808 (N_10808,N_10177,N_10372);
xnor U10809 (N_10809,N_10249,N_10301);
nor U10810 (N_10810,N_10140,N_10190);
or U10811 (N_10811,N_10090,N_10294);
nor U10812 (N_10812,N_10274,N_10262);
nand U10813 (N_10813,N_10193,N_10195);
xnor U10814 (N_10814,N_10304,N_10409);
and U10815 (N_10815,N_10371,N_10464);
nand U10816 (N_10816,N_10106,N_10229);
nand U10817 (N_10817,N_10399,N_10224);
nor U10818 (N_10818,N_10196,N_10099);
and U10819 (N_10819,N_10428,N_10092);
nor U10820 (N_10820,N_10373,N_10117);
xnor U10821 (N_10821,N_10034,N_10421);
nand U10822 (N_10822,N_10212,N_10375);
and U10823 (N_10823,N_10012,N_10126);
nor U10824 (N_10824,N_10200,N_10440);
and U10825 (N_10825,N_10126,N_10339);
and U10826 (N_10826,N_10371,N_10182);
nand U10827 (N_10827,N_10376,N_10412);
or U10828 (N_10828,N_10118,N_10026);
and U10829 (N_10829,N_10315,N_10426);
nand U10830 (N_10830,N_10049,N_10437);
nor U10831 (N_10831,N_10327,N_10454);
and U10832 (N_10832,N_10081,N_10361);
nor U10833 (N_10833,N_10493,N_10240);
nand U10834 (N_10834,N_10320,N_10341);
nand U10835 (N_10835,N_10404,N_10145);
and U10836 (N_10836,N_10495,N_10325);
nand U10837 (N_10837,N_10456,N_10269);
or U10838 (N_10838,N_10366,N_10384);
and U10839 (N_10839,N_10271,N_10462);
nand U10840 (N_10840,N_10321,N_10370);
xnor U10841 (N_10841,N_10231,N_10359);
or U10842 (N_10842,N_10247,N_10367);
and U10843 (N_10843,N_10333,N_10188);
xnor U10844 (N_10844,N_10178,N_10099);
or U10845 (N_10845,N_10219,N_10492);
and U10846 (N_10846,N_10236,N_10186);
xor U10847 (N_10847,N_10276,N_10205);
nor U10848 (N_10848,N_10358,N_10015);
xnor U10849 (N_10849,N_10107,N_10277);
xnor U10850 (N_10850,N_10103,N_10363);
and U10851 (N_10851,N_10201,N_10012);
and U10852 (N_10852,N_10141,N_10204);
nand U10853 (N_10853,N_10144,N_10292);
nand U10854 (N_10854,N_10459,N_10031);
nand U10855 (N_10855,N_10130,N_10284);
xnor U10856 (N_10856,N_10178,N_10041);
nor U10857 (N_10857,N_10101,N_10216);
xor U10858 (N_10858,N_10383,N_10460);
or U10859 (N_10859,N_10010,N_10168);
or U10860 (N_10860,N_10000,N_10467);
xnor U10861 (N_10861,N_10324,N_10290);
or U10862 (N_10862,N_10026,N_10102);
xor U10863 (N_10863,N_10242,N_10455);
and U10864 (N_10864,N_10031,N_10057);
xor U10865 (N_10865,N_10394,N_10436);
nor U10866 (N_10866,N_10128,N_10109);
nand U10867 (N_10867,N_10368,N_10152);
xnor U10868 (N_10868,N_10222,N_10440);
nand U10869 (N_10869,N_10315,N_10466);
nand U10870 (N_10870,N_10324,N_10130);
xor U10871 (N_10871,N_10300,N_10026);
nand U10872 (N_10872,N_10140,N_10341);
xor U10873 (N_10873,N_10370,N_10296);
nor U10874 (N_10874,N_10462,N_10126);
xnor U10875 (N_10875,N_10280,N_10295);
nor U10876 (N_10876,N_10419,N_10035);
xor U10877 (N_10877,N_10253,N_10083);
nand U10878 (N_10878,N_10226,N_10305);
nor U10879 (N_10879,N_10449,N_10101);
and U10880 (N_10880,N_10173,N_10191);
and U10881 (N_10881,N_10167,N_10242);
or U10882 (N_10882,N_10166,N_10343);
nor U10883 (N_10883,N_10006,N_10241);
and U10884 (N_10884,N_10294,N_10204);
and U10885 (N_10885,N_10369,N_10100);
and U10886 (N_10886,N_10408,N_10286);
nand U10887 (N_10887,N_10160,N_10316);
and U10888 (N_10888,N_10404,N_10123);
nand U10889 (N_10889,N_10375,N_10147);
or U10890 (N_10890,N_10319,N_10231);
or U10891 (N_10891,N_10355,N_10042);
or U10892 (N_10892,N_10037,N_10156);
and U10893 (N_10893,N_10370,N_10331);
or U10894 (N_10894,N_10443,N_10333);
and U10895 (N_10895,N_10072,N_10200);
or U10896 (N_10896,N_10315,N_10318);
or U10897 (N_10897,N_10055,N_10401);
xnor U10898 (N_10898,N_10455,N_10134);
nor U10899 (N_10899,N_10301,N_10402);
and U10900 (N_10900,N_10461,N_10088);
and U10901 (N_10901,N_10081,N_10046);
nor U10902 (N_10902,N_10421,N_10451);
nor U10903 (N_10903,N_10471,N_10159);
nor U10904 (N_10904,N_10115,N_10441);
nor U10905 (N_10905,N_10173,N_10268);
nor U10906 (N_10906,N_10179,N_10113);
or U10907 (N_10907,N_10436,N_10110);
or U10908 (N_10908,N_10488,N_10420);
xor U10909 (N_10909,N_10411,N_10137);
nor U10910 (N_10910,N_10275,N_10231);
xor U10911 (N_10911,N_10124,N_10405);
nor U10912 (N_10912,N_10112,N_10257);
xor U10913 (N_10913,N_10441,N_10440);
and U10914 (N_10914,N_10118,N_10294);
xor U10915 (N_10915,N_10128,N_10008);
or U10916 (N_10916,N_10431,N_10123);
nand U10917 (N_10917,N_10303,N_10009);
nor U10918 (N_10918,N_10069,N_10332);
nand U10919 (N_10919,N_10289,N_10382);
nor U10920 (N_10920,N_10313,N_10301);
nand U10921 (N_10921,N_10406,N_10313);
or U10922 (N_10922,N_10438,N_10054);
nor U10923 (N_10923,N_10332,N_10061);
xor U10924 (N_10924,N_10462,N_10185);
nand U10925 (N_10925,N_10095,N_10226);
and U10926 (N_10926,N_10461,N_10256);
or U10927 (N_10927,N_10342,N_10193);
xor U10928 (N_10928,N_10092,N_10200);
xnor U10929 (N_10929,N_10272,N_10485);
nor U10930 (N_10930,N_10435,N_10085);
and U10931 (N_10931,N_10039,N_10197);
nor U10932 (N_10932,N_10152,N_10466);
nand U10933 (N_10933,N_10497,N_10449);
nand U10934 (N_10934,N_10018,N_10038);
nand U10935 (N_10935,N_10313,N_10285);
nor U10936 (N_10936,N_10256,N_10436);
or U10937 (N_10937,N_10374,N_10270);
nor U10938 (N_10938,N_10146,N_10142);
nand U10939 (N_10939,N_10157,N_10484);
and U10940 (N_10940,N_10069,N_10127);
and U10941 (N_10941,N_10387,N_10044);
nor U10942 (N_10942,N_10076,N_10315);
xor U10943 (N_10943,N_10473,N_10169);
xor U10944 (N_10944,N_10446,N_10175);
and U10945 (N_10945,N_10123,N_10308);
xor U10946 (N_10946,N_10495,N_10229);
xnor U10947 (N_10947,N_10149,N_10411);
or U10948 (N_10948,N_10344,N_10082);
nand U10949 (N_10949,N_10370,N_10249);
and U10950 (N_10950,N_10289,N_10198);
nor U10951 (N_10951,N_10341,N_10369);
or U10952 (N_10952,N_10327,N_10332);
or U10953 (N_10953,N_10494,N_10497);
xnor U10954 (N_10954,N_10047,N_10478);
xor U10955 (N_10955,N_10347,N_10050);
nand U10956 (N_10956,N_10222,N_10416);
nand U10957 (N_10957,N_10037,N_10162);
and U10958 (N_10958,N_10433,N_10007);
xor U10959 (N_10959,N_10152,N_10028);
nand U10960 (N_10960,N_10124,N_10019);
xor U10961 (N_10961,N_10430,N_10160);
or U10962 (N_10962,N_10176,N_10180);
nand U10963 (N_10963,N_10468,N_10195);
xor U10964 (N_10964,N_10429,N_10390);
nor U10965 (N_10965,N_10422,N_10310);
or U10966 (N_10966,N_10335,N_10408);
nor U10967 (N_10967,N_10101,N_10149);
xor U10968 (N_10968,N_10124,N_10084);
nor U10969 (N_10969,N_10163,N_10294);
nor U10970 (N_10970,N_10083,N_10312);
or U10971 (N_10971,N_10327,N_10174);
and U10972 (N_10972,N_10219,N_10408);
and U10973 (N_10973,N_10265,N_10218);
and U10974 (N_10974,N_10496,N_10442);
or U10975 (N_10975,N_10353,N_10063);
and U10976 (N_10976,N_10212,N_10426);
or U10977 (N_10977,N_10411,N_10273);
nand U10978 (N_10978,N_10187,N_10247);
or U10979 (N_10979,N_10358,N_10176);
xnor U10980 (N_10980,N_10417,N_10325);
nand U10981 (N_10981,N_10298,N_10468);
and U10982 (N_10982,N_10329,N_10056);
or U10983 (N_10983,N_10013,N_10118);
or U10984 (N_10984,N_10382,N_10210);
and U10985 (N_10985,N_10460,N_10178);
or U10986 (N_10986,N_10025,N_10221);
xnor U10987 (N_10987,N_10184,N_10285);
nand U10988 (N_10988,N_10363,N_10202);
and U10989 (N_10989,N_10363,N_10445);
nor U10990 (N_10990,N_10494,N_10127);
nor U10991 (N_10991,N_10234,N_10021);
nor U10992 (N_10992,N_10199,N_10452);
nand U10993 (N_10993,N_10388,N_10077);
nand U10994 (N_10994,N_10451,N_10211);
xnor U10995 (N_10995,N_10137,N_10127);
nand U10996 (N_10996,N_10022,N_10416);
nor U10997 (N_10997,N_10448,N_10095);
and U10998 (N_10998,N_10246,N_10369);
or U10999 (N_10999,N_10134,N_10465);
or U11000 (N_11000,N_10807,N_10835);
nand U11001 (N_11001,N_10707,N_10511);
nor U11002 (N_11002,N_10672,N_10990);
nand U11003 (N_11003,N_10921,N_10586);
or U11004 (N_11004,N_10768,N_10713);
and U11005 (N_11005,N_10681,N_10683);
nand U11006 (N_11006,N_10877,N_10565);
and U11007 (N_11007,N_10640,N_10972);
nor U11008 (N_11008,N_10793,N_10609);
xnor U11009 (N_11009,N_10744,N_10880);
nor U11010 (N_11010,N_10992,N_10950);
and U11011 (N_11011,N_10561,N_10675);
nand U11012 (N_11012,N_10906,N_10529);
xor U11013 (N_11013,N_10890,N_10520);
nand U11014 (N_11014,N_10548,N_10542);
nor U11015 (N_11015,N_10616,N_10706);
nor U11016 (N_11016,N_10957,N_10948);
xnor U11017 (N_11017,N_10704,N_10836);
xnor U11018 (N_11018,N_10708,N_10770);
nor U11019 (N_11019,N_10766,N_10999);
and U11020 (N_11020,N_10997,N_10513);
and U11021 (N_11021,N_10832,N_10850);
or U11022 (N_11022,N_10522,N_10691);
and U11023 (N_11023,N_10748,N_10965);
and U11024 (N_11024,N_10996,N_10699);
or U11025 (N_11025,N_10914,N_10525);
nand U11026 (N_11026,N_10620,N_10858);
xor U11027 (N_11027,N_10781,N_10827);
xor U11028 (N_11028,N_10570,N_10834);
nand U11029 (N_11029,N_10651,N_10593);
xor U11030 (N_11030,N_10682,N_10897);
nand U11031 (N_11031,N_10749,N_10650);
xor U11032 (N_11032,N_10902,N_10842);
nor U11033 (N_11033,N_10567,N_10856);
and U11034 (N_11034,N_10879,N_10639);
nor U11035 (N_11035,N_10979,N_10645);
or U11036 (N_11036,N_10841,N_10790);
or U11037 (N_11037,N_10503,N_10732);
nand U11038 (N_11038,N_10539,N_10769);
and U11039 (N_11039,N_10760,N_10846);
nor U11040 (N_11040,N_10578,N_10753);
xor U11041 (N_11041,N_10989,N_10915);
xor U11042 (N_11042,N_10688,N_10961);
nand U11043 (N_11043,N_10805,N_10727);
or U11044 (N_11044,N_10978,N_10730);
and U11045 (N_11045,N_10696,N_10637);
nand U11046 (N_11046,N_10538,N_10819);
xnor U11047 (N_11047,N_10767,N_10589);
nand U11048 (N_11048,N_10919,N_10636);
nand U11049 (N_11049,N_10502,N_10632);
xor U11050 (N_11050,N_10554,N_10563);
and U11051 (N_11051,N_10527,N_10679);
nand U11052 (N_11052,N_10888,N_10864);
nor U11053 (N_11053,N_10943,N_10772);
and U11054 (N_11054,N_10701,N_10544);
nor U11055 (N_11055,N_10558,N_10778);
nor U11056 (N_11056,N_10981,N_10971);
nand U11057 (N_11057,N_10531,N_10606);
nor U11058 (N_11058,N_10714,N_10505);
nand U11059 (N_11059,N_10519,N_10952);
or U11060 (N_11060,N_10956,N_10630);
and U11061 (N_11061,N_10776,N_10725);
and U11062 (N_11062,N_10722,N_10745);
xnor U11063 (N_11063,N_10625,N_10739);
xnor U11064 (N_11064,N_10799,N_10986);
nor U11065 (N_11065,N_10809,N_10677);
nor U11066 (N_11066,N_10559,N_10951);
and U11067 (N_11067,N_10723,N_10654);
or U11068 (N_11068,N_10711,N_10810);
nand U11069 (N_11069,N_10551,N_10811);
or U11070 (N_11070,N_10692,N_10761);
xor U11071 (N_11071,N_10506,N_10912);
nor U11072 (N_11072,N_10823,N_10881);
nand U11073 (N_11073,N_10817,N_10631);
xnor U11074 (N_11074,N_10607,N_10905);
xnor U11075 (N_11075,N_10621,N_10964);
and U11076 (N_11076,N_10967,N_10755);
nand U11077 (N_11077,N_10818,N_10710);
or U11078 (N_11078,N_10878,N_10695);
and U11079 (N_11079,N_10762,N_10741);
nor U11080 (N_11080,N_10633,N_10541);
nand U11081 (N_11081,N_10641,N_10794);
or U11082 (N_11082,N_10900,N_10629);
and U11083 (N_11083,N_10798,N_10945);
nor U11084 (N_11084,N_10994,N_10825);
nor U11085 (N_11085,N_10754,N_10715);
or U11086 (N_11086,N_10930,N_10617);
or U11087 (N_11087,N_10597,N_10931);
and U11088 (N_11088,N_10815,N_10546);
xor U11089 (N_11089,N_10975,N_10535);
xor U11090 (N_11090,N_10742,N_10602);
or U11091 (N_11091,N_10892,N_10816);
or U11092 (N_11092,N_10826,N_10765);
or U11093 (N_11093,N_10608,N_10598);
and U11094 (N_11094,N_10954,N_10847);
xor U11095 (N_11095,N_10938,N_10782);
nand U11096 (N_11096,N_10916,N_10581);
nor U11097 (N_11097,N_10624,N_10791);
or U11098 (N_11098,N_10737,N_10733);
nand U11099 (N_11099,N_10557,N_10909);
and U11100 (N_11100,N_10628,N_10980);
xnor U11101 (N_11101,N_10547,N_10569);
and U11102 (N_11102,N_10500,N_10573);
and U11103 (N_11103,N_10987,N_10974);
or U11104 (N_11104,N_10564,N_10984);
and U11105 (N_11105,N_10869,N_10876);
or U11106 (N_11106,N_10545,N_10526);
and U11107 (N_11107,N_10703,N_10797);
nor U11108 (N_11108,N_10649,N_10949);
xor U11109 (N_11109,N_10893,N_10851);
or U11110 (N_11110,N_10911,N_10611);
nor U11111 (N_11111,N_10627,N_10947);
xor U11112 (N_11112,N_10686,N_10687);
nand U11113 (N_11113,N_10813,N_10728);
or U11114 (N_11114,N_10595,N_10668);
nor U11115 (N_11115,N_10838,N_10849);
xnor U11116 (N_11116,N_10599,N_10872);
and U11117 (N_11117,N_10623,N_10953);
and U11118 (N_11118,N_10924,N_10576);
nor U11119 (N_11119,N_10689,N_10575);
xor U11120 (N_11120,N_10925,N_10516);
nor U11121 (N_11121,N_10923,N_10820);
nand U11122 (N_11122,N_10837,N_10963);
xnor U11123 (N_11123,N_10792,N_10812);
xor U11124 (N_11124,N_10870,N_10536);
or U11125 (N_11125,N_10543,N_10592);
nand U11126 (N_11126,N_10577,N_10552);
or U11127 (N_11127,N_10635,N_10933);
or U11128 (N_11128,N_10663,N_10763);
or U11129 (N_11129,N_10644,N_10610);
xnor U11130 (N_11130,N_10709,N_10553);
nand U11131 (N_11131,N_10862,N_10787);
and U11132 (N_11132,N_10712,N_10659);
nor U11133 (N_11133,N_10795,N_10619);
nand U11134 (N_11134,N_10676,N_10868);
and U11135 (N_11135,N_10752,N_10588);
and U11136 (N_11136,N_10904,N_10803);
and U11137 (N_11137,N_10901,N_10674);
and U11138 (N_11138,N_10508,N_10603);
xnor U11139 (N_11139,N_10800,N_10998);
nand U11140 (N_11140,N_10895,N_10775);
or U11141 (N_11141,N_10671,N_10518);
nand U11142 (N_11142,N_10774,N_10653);
nand U11143 (N_11143,N_10991,N_10562);
nand U11144 (N_11144,N_10796,N_10962);
and U11145 (N_11145,N_10764,N_10885);
or U11146 (N_11146,N_10751,N_10560);
nor U11147 (N_11147,N_10604,N_10666);
and U11148 (N_11148,N_10955,N_10647);
xnor U11149 (N_11149,N_10910,N_10936);
nor U11150 (N_11150,N_10521,N_10731);
and U11151 (N_11151,N_10969,N_10937);
or U11152 (N_11152,N_10697,N_10995);
xnor U11153 (N_11153,N_10882,N_10808);
and U11154 (N_11154,N_10786,N_10966);
xnor U11155 (N_11155,N_10960,N_10549);
nor U11156 (N_11156,N_10783,N_10638);
nand U11157 (N_11157,N_10678,N_10585);
or U11158 (N_11158,N_10747,N_10612);
xor U11159 (N_11159,N_10555,N_10779);
and U11160 (N_11160,N_10828,N_10759);
nand U11161 (N_11161,N_10524,N_10985);
nand U11162 (N_11162,N_10514,N_10515);
nand U11163 (N_11163,N_10643,N_10928);
nor U11164 (N_11164,N_10814,N_10777);
xnor U11165 (N_11165,N_10926,N_10771);
and U11166 (N_11166,N_10568,N_10702);
nor U11167 (N_11167,N_10939,N_10579);
nand U11168 (N_11168,N_10883,N_10587);
and U11169 (N_11169,N_10591,N_10746);
or U11170 (N_11170,N_10773,N_10942);
or U11171 (N_11171,N_10845,N_10684);
xor U11172 (N_11172,N_10556,N_10865);
and U11173 (N_11173,N_10920,N_10572);
nor U11174 (N_11174,N_10824,N_10866);
nand U11175 (N_11175,N_10664,N_10660);
and U11176 (N_11176,N_10922,N_10750);
or U11177 (N_11177,N_10907,N_10615);
nand U11178 (N_11178,N_10642,N_10863);
or U11179 (N_11179,N_10669,N_10861);
nand U11180 (N_11180,N_10622,N_10894);
or U11181 (N_11181,N_10871,N_10917);
xnor U11182 (N_11182,N_10721,N_10873);
nand U11183 (N_11183,N_10512,N_10594);
or U11184 (N_11184,N_10736,N_10517);
nand U11185 (N_11185,N_10789,N_10970);
nor U11186 (N_11186,N_10973,N_10932);
xor U11187 (N_11187,N_10889,N_10719);
xor U11188 (N_11188,N_10618,N_10694);
nand U11189 (N_11189,N_10605,N_10648);
and U11190 (N_11190,N_10662,N_10927);
and U11191 (N_11191,N_10685,N_10988);
nor U11192 (N_11192,N_10854,N_10537);
or U11193 (N_11193,N_10528,N_10839);
xor U11194 (N_11194,N_10740,N_10801);
or U11195 (N_11195,N_10670,N_10959);
xnor U11196 (N_11196,N_10540,N_10584);
or U11197 (N_11197,N_10756,N_10652);
nor U11198 (N_11198,N_10887,N_10896);
nor U11199 (N_11199,N_10855,N_10698);
xnor U11200 (N_11200,N_10946,N_10501);
nor U11201 (N_11201,N_10658,N_10859);
nor U11202 (N_11202,N_10891,N_10982);
nand U11203 (N_11203,N_10886,N_10843);
nand U11204 (N_11204,N_10550,N_10918);
nor U11205 (N_11205,N_10574,N_10780);
or U11206 (N_11206,N_10852,N_10833);
xnor U11207 (N_11207,N_10530,N_10729);
nor U11208 (N_11208,N_10976,N_10596);
xor U11209 (N_11209,N_10724,N_10690);
and U11210 (N_11210,N_10507,N_10743);
nor U11211 (N_11211,N_10844,N_10788);
nand U11212 (N_11212,N_10655,N_10720);
nand U11213 (N_11213,N_10898,N_10580);
xor U11214 (N_11214,N_10532,N_10738);
or U11215 (N_11215,N_10735,N_10700);
nand U11216 (N_11216,N_10661,N_10582);
nand U11217 (N_11217,N_10614,N_10734);
or U11218 (N_11218,N_10533,N_10830);
and U11219 (N_11219,N_10983,N_10993);
nand U11220 (N_11220,N_10831,N_10935);
nand U11221 (N_11221,N_10853,N_10634);
nor U11222 (N_11222,N_10875,N_10718);
or U11223 (N_11223,N_10903,N_10656);
nor U11224 (N_11224,N_10958,N_10758);
or U11225 (N_11225,N_10802,N_10757);
or U11226 (N_11226,N_10867,N_10899);
nand U11227 (N_11227,N_10829,N_10667);
nor U11228 (N_11228,N_10680,N_10857);
nor U11229 (N_11229,N_10600,N_10583);
and U11230 (N_11230,N_10726,N_10860);
or U11231 (N_11231,N_10566,N_10848);
or U11232 (N_11232,N_10534,N_10613);
and U11233 (N_11233,N_10693,N_10504);
xor U11234 (N_11234,N_10806,N_10509);
nand U11235 (N_11235,N_10944,N_10804);
or U11236 (N_11236,N_10822,N_10523);
and U11237 (N_11237,N_10940,N_10705);
nand U11238 (N_11238,N_10941,N_10716);
or U11239 (N_11239,N_10785,N_10665);
and U11240 (N_11240,N_10934,N_10884);
xnor U11241 (N_11241,N_10874,N_10590);
xnor U11242 (N_11242,N_10510,N_10913);
nand U11243 (N_11243,N_10908,N_10626);
or U11244 (N_11244,N_10821,N_10673);
nand U11245 (N_11245,N_10977,N_10784);
or U11246 (N_11246,N_10571,N_10646);
xnor U11247 (N_11247,N_10929,N_10717);
nor U11248 (N_11248,N_10601,N_10657);
or U11249 (N_11249,N_10968,N_10840);
nor U11250 (N_11250,N_10613,N_10706);
or U11251 (N_11251,N_10564,N_10584);
nand U11252 (N_11252,N_10595,N_10671);
nand U11253 (N_11253,N_10586,N_10763);
and U11254 (N_11254,N_10504,N_10963);
nor U11255 (N_11255,N_10704,N_10879);
nand U11256 (N_11256,N_10988,N_10555);
and U11257 (N_11257,N_10677,N_10609);
and U11258 (N_11258,N_10636,N_10789);
xnor U11259 (N_11259,N_10988,N_10801);
nor U11260 (N_11260,N_10570,N_10611);
and U11261 (N_11261,N_10706,N_10546);
or U11262 (N_11262,N_10527,N_10522);
nor U11263 (N_11263,N_10864,N_10775);
and U11264 (N_11264,N_10680,N_10759);
nand U11265 (N_11265,N_10842,N_10742);
or U11266 (N_11266,N_10821,N_10920);
or U11267 (N_11267,N_10907,N_10510);
xnor U11268 (N_11268,N_10686,N_10964);
nor U11269 (N_11269,N_10781,N_10565);
nand U11270 (N_11270,N_10649,N_10819);
xor U11271 (N_11271,N_10691,N_10679);
or U11272 (N_11272,N_10685,N_10633);
nand U11273 (N_11273,N_10827,N_10761);
nand U11274 (N_11274,N_10985,N_10775);
nor U11275 (N_11275,N_10644,N_10963);
nand U11276 (N_11276,N_10588,N_10781);
or U11277 (N_11277,N_10654,N_10865);
nor U11278 (N_11278,N_10977,N_10547);
or U11279 (N_11279,N_10794,N_10966);
and U11280 (N_11280,N_10679,N_10712);
nand U11281 (N_11281,N_10917,N_10852);
xnor U11282 (N_11282,N_10735,N_10542);
and U11283 (N_11283,N_10743,N_10803);
and U11284 (N_11284,N_10698,N_10535);
or U11285 (N_11285,N_10912,N_10571);
or U11286 (N_11286,N_10677,N_10668);
nor U11287 (N_11287,N_10635,N_10504);
and U11288 (N_11288,N_10905,N_10921);
nor U11289 (N_11289,N_10716,N_10533);
and U11290 (N_11290,N_10823,N_10856);
xor U11291 (N_11291,N_10773,N_10724);
xnor U11292 (N_11292,N_10709,N_10946);
nand U11293 (N_11293,N_10508,N_10895);
and U11294 (N_11294,N_10943,N_10756);
and U11295 (N_11295,N_10753,N_10712);
xnor U11296 (N_11296,N_10809,N_10851);
xnor U11297 (N_11297,N_10809,N_10738);
and U11298 (N_11298,N_10710,N_10954);
nand U11299 (N_11299,N_10853,N_10585);
and U11300 (N_11300,N_10779,N_10717);
nand U11301 (N_11301,N_10968,N_10722);
or U11302 (N_11302,N_10882,N_10531);
xor U11303 (N_11303,N_10550,N_10646);
or U11304 (N_11304,N_10766,N_10971);
xor U11305 (N_11305,N_10859,N_10957);
nor U11306 (N_11306,N_10636,N_10586);
nand U11307 (N_11307,N_10952,N_10888);
or U11308 (N_11308,N_10618,N_10523);
or U11309 (N_11309,N_10921,N_10648);
nor U11310 (N_11310,N_10912,N_10896);
nor U11311 (N_11311,N_10568,N_10698);
and U11312 (N_11312,N_10565,N_10736);
or U11313 (N_11313,N_10705,N_10668);
and U11314 (N_11314,N_10992,N_10622);
and U11315 (N_11315,N_10770,N_10760);
or U11316 (N_11316,N_10902,N_10639);
and U11317 (N_11317,N_10921,N_10854);
xnor U11318 (N_11318,N_10704,N_10976);
xor U11319 (N_11319,N_10996,N_10979);
xor U11320 (N_11320,N_10991,N_10591);
or U11321 (N_11321,N_10550,N_10795);
or U11322 (N_11322,N_10580,N_10894);
or U11323 (N_11323,N_10832,N_10559);
nor U11324 (N_11324,N_10868,N_10829);
and U11325 (N_11325,N_10697,N_10595);
nand U11326 (N_11326,N_10900,N_10506);
xor U11327 (N_11327,N_10678,N_10970);
xnor U11328 (N_11328,N_10712,N_10674);
nand U11329 (N_11329,N_10894,N_10742);
nor U11330 (N_11330,N_10972,N_10869);
or U11331 (N_11331,N_10728,N_10782);
nand U11332 (N_11332,N_10671,N_10701);
xor U11333 (N_11333,N_10630,N_10519);
or U11334 (N_11334,N_10532,N_10761);
nor U11335 (N_11335,N_10939,N_10531);
or U11336 (N_11336,N_10841,N_10947);
or U11337 (N_11337,N_10736,N_10797);
or U11338 (N_11338,N_10606,N_10683);
nand U11339 (N_11339,N_10880,N_10858);
xnor U11340 (N_11340,N_10727,N_10506);
nor U11341 (N_11341,N_10538,N_10683);
xnor U11342 (N_11342,N_10722,N_10875);
nand U11343 (N_11343,N_10567,N_10981);
nor U11344 (N_11344,N_10853,N_10532);
and U11345 (N_11345,N_10747,N_10891);
xor U11346 (N_11346,N_10761,N_10758);
nor U11347 (N_11347,N_10539,N_10816);
nor U11348 (N_11348,N_10754,N_10763);
nor U11349 (N_11349,N_10769,N_10559);
xnor U11350 (N_11350,N_10603,N_10741);
nand U11351 (N_11351,N_10748,N_10652);
or U11352 (N_11352,N_10825,N_10676);
nand U11353 (N_11353,N_10801,N_10619);
and U11354 (N_11354,N_10752,N_10823);
or U11355 (N_11355,N_10846,N_10944);
nor U11356 (N_11356,N_10526,N_10696);
nor U11357 (N_11357,N_10634,N_10872);
and U11358 (N_11358,N_10605,N_10927);
and U11359 (N_11359,N_10506,N_10954);
nand U11360 (N_11360,N_10587,N_10997);
and U11361 (N_11361,N_10715,N_10531);
nand U11362 (N_11362,N_10874,N_10976);
or U11363 (N_11363,N_10519,N_10824);
nor U11364 (N_11364,N_10642,N_10726);
or U11365 (N_11365,N_10599,N_10656);
or U11366 (N_11366,N_10977,N_10961);
and U11367 (N_11367,N_10581,N_10623);
and U11368 (N_11368,N_10898,N_10540);
xnor U11369 (N_11369,N_10561,N_10895);
or U11370 (N_11370,N_10599,N_10865);
xnor U11371 (N_11371,N_10677,N_10576);
or U11372 (N_11372,N_10983,N_10902);
xnor U11373 (N_11373,N_10919,N_10503);
nand U11374 (N_11374,N_10813,N_10601);
nor U11375 (N_11375,N_10611,N_10663);
nand U11376 (N_11376,N_10621,N_10521);
nand U11377 (N_11377,N_10650,N_10864);
xnor U11378 (N_11378,N_10921,N_10692);
and U11379 (N_11379,N_10830,N_10948);
xor U11380 (N_11380,N_10578,N_10811);
nand U11381 (N_11381,N_10943,N_10790);
nor U11382 (N_11382,N_10620,N_10592);
and U11383 (N_11383,N_10825,N_10869);
and U11384 (N_11384,N_10726,N_10778);
or U11385 (N_11385,N_10828,N_10883);
and U11386 (N_11386,N_10833,N_10732);
xor U11387 (N_11387,N_10714,N_10544);
or U11388 (N_11388,N_10761,N_10958);
xor U11389 (N_11389,N_10789,N_10511);
and U11390 (N_11390,N_10915,N_10500);
nor U11391 (N_11391,N_10788,N_10588);
or U11392 (N_11392,N_10719,N_10784);
or U11393 (N_11393,N_10973,N_10612);
xor U11394 (N_11394,N_10836,N_10712);
xnor U11395 (N_11395,N_10512,N_10712);
and U11396 (N_11396,N_10786,N_10597);
xnor U11397 (N_11397,N_10524,N_10554);
nand U11398 (N_11398,N_10655,N_10911);
xnor U11399 (N_11399,N_10838,N_10518);
or U11400 (N_11400,N_10858,N_10564);
xor U11401 (N_11401,N_10831,N_10897);
nor U11402 (N_11402,N_10817,N_10762);
nand U11403 (N_11403,N_10689,N_10750);
xnor U11404 (N_11404,N_10531,N_10661);
or U11405 (N_11405,N_10693,N_10552);
or U11406 (N_11406,N_10939,N_10912);
and U11407 (N_11407,N_10967,N_10916);
and U11408 (N_11408,N_10642,N_10672);
nor U11409 (N_11409,N_10692,N_10951);
nor U11410 (N_11410,N_10681,N_10758);
nand U11411 (N_11411,N_10570,N_10898);
and U11412 (N_11412,N_10662,N_10524);
nor U11413 (N_11413,N_10732,N_10607);
nor U11414 (N_11414,N_10842,N_10528);
or U11415 (N_11415,N_10603,N_10841);
or U11416 (N_11416,N_10606,N_10803);
xnor U11417 (N_11417,N_10949,N_10833);
nand U11418 (N_11418,N_10697,N_10646);
xnor U11419 (N_11419,N_10852,N_10976);
or U11420 (N_11420,N_10867,N_10949);
nor U11421 (N_11421,N_10920,N_10921);
or U11422 (N_11422,N_10528,N_10996);
xor U11423 (N_11423,N_10960,N_10849);
xor U11424 (N_11424,N_10944,N_10863);
nand U11425 (N_11425,N_10731,N_10922);
nor U11426 (N_11426,N_10601,N_10830);
nand U11427 (N_11427,N_10886,N_10521);
xnor U11428 (N_11428,N_10584,N_10510);
or U11429 (N_11429,N_10746,N_10983);
xnor U11430 (N_11430,N_10720,N_10922);
nor U11431 (N_11431,N_10995,N_10638);
xor U11432 (N_11432,N_10546,N_10664);
or U11433 (N_11433,N_10607,N_10638);
xor U11434 (N_11434,N_10971,N_10923);
or U11435 (N_11435,N_10841,N_10748);
nand U11436 (N_11436,N_10780,N_10993);
nand U11437 (N_11437,N_10813,N_10750);
nand U11438 (N_11438,N_10895,N_10877);
or U11439 (N_11439,N_10935,N_10759);
xnor U11440 (N_11440,N_10822,N_10929);
or U11441 (N_11441,N_10721,N_10982);
nand U11442 (N_11442,N_10674,N_10886);
nand U11443 (N_11443,N_10982,N_10557);
nand U11444 (N_11444,N_10916,N_10955);
nand U11445 (N_11445,N_10503,N_10544);
xnor U11446 (N_11446,N_10748,N_10883);
nor U11447 (N_11447,N_10860,N_10777);
xor U11448 (N_11448,N_10601,N_10687);
nor U11449 (N_11449,N_10718,N_10551);
nor U11450 (N_11450,N_10570,N_10534);
or U11451 (N_11451,N_10521,N_10878);
nand U11452 (N_11452,N_10678,N_10501);
and U11453 (N_11453,N_10585,N_10819);
xnor U11454 (N_11454,N_10713,N_10588);
nor U11455 (N_11455,N_10986,N_10937);
nor U11456 (N_11456,N_10961,N_10755);
nor U11457 (N_11457,N_10868,N_10982);
nor U11458 (N_11458,N_10840,N_10678);
nand U11459 (N_11459,N_10889,N_10936);
or U11460 (N_11460,N_10521,N_10722);
nor U11461 (N_11461,N_10991,N_10973);
or U11462 (N_11462,N_10927,N_10744);
nand U11463 (N_11463,N_10591,N_10502);
xnor U11464 (N_11464,N_10942,N_10546);
xnor U11465 (N_11465,N_10669,N_10985);
xor U11466 (N_11466,N_10806,N_10792);
xor U11467 (N_11467,N_10745,N_10683);
and U11468 (N_11468,N_10785,N_10693);
xnor U11469 (N_11469,N_10952,N_10807);
nor U11470 (N_11470,N_10514,N_10598);
nand U11471 (N_11471,N_10728,N_10677);
nand U11472 (N_11472,N_10552,N_10960);
and U11473 (N_11473,N_10617,N_10656);
nor U11474 (N_11474,N_10830,N_10743);
xor U11475 (N_11475,N_10859,N_10521);
nor U11476 (N_11476,N_10535,N_10867);
nand U11477 (N_11477,N_10963,N_10696);
nor U11478 (N_11478,N_10691,N_10888);
nand U11479 (N_11479,N_10966,N_10501);
or U11480 (N_11480,N_10646,N_10755);
and U11481 (N_11481,N_10682,N_10910);
or U11482 (N_11482,N_10504,N_10550);
and U11483 (N_11483,N_10568,N_10750);
nand U11484 (N_11484,N_10587,N_10875);
nand U11485 (N_11485,N_10545,N_10604);
xor U11486 (N_11486,N_10534,N_10728);
or U11487 (N_11487,N_10596,N_10690);
xnor U11488 (N_11488,N_10906,N_10977);
or U11489 (N_11489,N_10909,N_10715);
and U11490 (N_11490,N_10727,N_10653);
nand U11491 (N_11491,N_10830,N_10581);
and U11492 (N_11492,N_10696,N_10625);
nor U11493 (N_11493,N_10634,N_10665);
nor U11494 (N_11494,N_10662,N_10709);
nor U11495 (N_11495,N_10503,N_10821);
and U11496 (N_11496,N_10706,N_10544);
and U11497 (N_11497,N_10581,N_10502);
and U11498 (N_11498,N_10706,N_10537);
or U11499 (N_11499,N_10906,N_10690);
nand U11500 (N_11500,N_11459,N_11319);
nor U11501 (N_11501,N_11178,N_11120);
xnor U11502 (N_11502,N_11285,N_11113);
nand U11503 (N_11503,N_11355,N_11040);
xnor U11504 (N_11504,N_11123,N_11324);
or U11505 (N_11505,N_11346,N_11337);
and U11506 (N_11506,N_11339,N_11226);
and U11507 (N_11507,N_11354,N_11102);
and U11508 (N_11508,N_11410,N_11073);
or U11509 (N_11509,N_11338,N_11399);
xor U11510 (N_11510,N_11079,N_11024);
nand U11511 (N_11511,N_11303,N_11100);
nor U11512 (N_11512,N_11035,N_11363);
nor U11513 (N_11513,N_11219,N_11058);
and U11514 (N_11514,N_11137,N_11236);
or U11515 (N_11515,N_11315,N_11187);
or U11516 (N_11516,N_11037,N_11259);
xor U11517 (N_11517,N_11179,N_11275);
or U11518 (N_11518,N_11046,N_11320);
nand U11519 (N_11519,N_11062,N_11468);
and U11520 (N_11520,N_11281,N_11034);
xnor U11521 (N_11521,N_11496,N_11116);
nor U11522 (N_11522,N_11237,N_11483);
nor U11523 (N_11523,N_11371,N_11186);
or U11524 (N_11524,N_11292,N_11366);
or U11525 (N_11525,N_11183,N_11191);
or U11526 (N_11526,N_11299,N_11432);
and U11527 (N_11527,N_11009,N_11499);
xnor U11528 (N_11528,N_11447,N_11429);
xnor U11529 (N_11529,N_11039,N_11398);
nor U11530 (N_11530,N_11203,N_11061);
xnor U11531 (N_11531,N_11312,N_11038);
xnor U11532 (N_11532,N_11165,N_11420);
xor U11533 (N_11533,N_11193,N_11241);
nand U11534 (N_11534,N_11243,N_11151);
xnor U11535 (N_11535,N_11020,N_11416);
xnor U11536 (N_11536,N_11052,N_11387);
nand U11537 (N_11537,N_11247,N_11492);
or U11538 (N_11538,N_11016,N_11351);
xor U11539 (N_11539,N_11345,N_11010);
xnor U11540 (N_11540,N_11407,N_11457);
and U11541 (N_11541,N_11172,N_11385);
and U11542 (N_11542,N_11198,N_11087);
and U11543 (N_11543,N_11199,N_11152);
nand U11544 (N_11544,N_11284,N_11099);
or U11545 (N_11545,N_11174,N_11002);
xnor U11546 (N_11546,N_11445,N_11290);
nor U11547 (N_11547,N_11450,N_11173);
nor U11548 (N_11548,N_11094,N_11091);
xor U11549 (N_11549,N_11357,N_11467);
xor U11550 (N_11550,N_11111,N_11273);
or U11551 (N_11551,N_11049,N_11030);
and U11552 (N_11552,N_11015,N_11159);
and U11553 (N_11553,N_11149,N_11456);
nor U11554 (N_11554,N_11434,N_11437);
nor U11555 (N_11555,N_11489,N_11001);
xnor U11556 (N_11556,N_11068,N_11287);
and U11557 (N_11557,N_11309,N_11274);
or U11558 (N_11558,N_11025,N_11378);
nor U11559 (N_11559,N_11029,N_11271);
and U11560 (N_11560,N_11466,N_11369);
nand U11561 (N_11561,N_11098,N_11426);
xor U11562 (N_11562,N_11164,N_11096);
nor U11563 (N_11563,N_11056,N_11263);
nand U11564 (N_11564,N_11406,N_11107);
and U11565 (N_11565,N_11300,N_11074);
nand U11566 (N_11566,N_11086,N_11332);
xor U11567 (N_11567,N_11258,N_11490);
nand U11568 (N_11568,N_11197,N_11019);
nor U11569 (N_11569,N_11280,N_11234);
nand U11570 (N_11570,N_11409,N_11394);
and U11571 (N_11571,N_11310,N_11491);
nand U11572 (N_11572,N_11372,N_11211);
xor U11573 (N_11573,N_11497,N_11452);
nand U11574 (N_11574,N_11155,N_11063);
nor U11575 (N_11575,N_11214,N_11449);
or U11576 (N_11576,N_11064,N_11383);
nand U11577 (N_11577,N_11270,N_11440);
nand U11578 (N_11578,N_11117,N_11423);
nor U11579 (N_11579,N_11140,N_11231);
or U11580 (N_11580,N_11185,N_11485);
or U11581 (N_11581,N_11408,N_11377);
or U11582 (N_11582,N_11458,N_11112);
xor U11583 (N_11583,N_11255,N_11139);
nor U11584 (N_11584,N_11433,N_11042);
or U11585 (N_11585,N_11359,N_11031);
and U11586 (N_11586,N_11043,N_11430);
nor U11587 (N_11587,N_11122,N_11133);
xor U11588 (N_11588,N_11352,N_11368);
nand U11589 (N_11589,N_11184,N_11257);
xnor U11590 (N_11590,N_11367,N_11207);
or U11591 (N_11591,N_11028,N_11256);
nor U11592 (N_11592,N_11375,N_11204);
nor U11593 (N_11593,N_11435,N_11305);
nand U11594 (N_11594,N_11047,N_11069);
xor U11595 (N_11595,N_11143,N_11004);
and U11596 (N_11596,N_11252,N_11484);
nor U11597 (N_11597,N_11109,N_11134);
nor U11598 (N_11598,N_11106,N_11041);
and U11599 (N_11599,N_11018,N_11446);
and U11600 (N_11600,N_11402,N_11253);
nand U11601 (N_11601,N_11147,N_11262);
and U11602 (N_11602,N_11481,N_11053);
and U11603 (N_11603,N_11036,N_11021);
and U11604 (N_11604,N_11431,N_11311);
nand U11605 (N_11605,N_11180,N_11386);
xor U11606 (N_11606,N_11390,N_11048);
xnor U11607 (N_11607,N_11264,N_11059);
and U11608 (N_11608,N_11453,N_11417);
and U11609 (N_11609,N_11331,N_11230);
and U11610 (N_11610,N_11293,N_11384);
nand U11611 (N_11611,N_11182,N_11395);
nor U11612 (N_11612,N_11477,N_11168);
and U11613 (N_11613,N_11391,N_11150);
xor U11614 (N_11614,N_11279,N_11007);
or U11615 (N_11615,N_11250,N_11475);
and U11616 (N_11616,N_11327,N_11200);
nand U11617 (N_11617,N_11192,N_11014);
nor U11618 (N_11618,N_11356,N_11013);
nor U11619 (N_11619,N_11488,N_11469);
nor U11620 (N_11620,N_11220,N_11050);
nand U11621 (N_11621,N_11487,N_11415);
or U11622 (N_11622,N_11413,N_11289);
and U11623 (N_11623,N_11254,N_11454);
xnor U11624 (N_11624,N_11295,N_11333);
nor U11625 (N_11625,N_11428,N_11397);
nor U11626 (N_11626,N_11114,N_11006);
or U11627 (N_11627,N_11474,N_11439);
nand U11628 (N_11628,N_11210,N_11067);
nand U11629 (N_11629,N_11343,N_11077);
nor U11630 (N_11630,N_11422,N_11451);
xnor U11631 (N_11631,N_11153,N_11405);
and U11632 (N_11632,N_11205,N_11498);
and U11633 (N_11633,N_11260,N_11022);
or U11634 (N_11634,N_11216,N_11379);
and U11635 (N_11635,N_11162,N_11127);
nand U11636 (N_11636,N_11023,N_11085);
xnor U11637 (N_11637,N_11361,N_11065);
and U11638 (N_11638,N_11131,N_11365);
xnor U11639 (N_11639,N_11225,N_11393);
nor U11640 (N_11640,N_11125,N_11121);
nor U11641 (N_11641,N_11334,N_11081);
and U11642 (N_11642,N_11245,N_11227);
nor U11643 (N_11643,N_11232,N_11321);
or U11644 (N_11644,N_11160,N_11328);
nor U11645 (N_11645,N_11078,N_11201);
nand U11646 (N_11646,N_11146,N_11104);
and U11647 (N_11647,N_11224,N_11071);
xnor U11648 (N_11648,N_11082,N_11438);
nor U11649 (N_11649,N_11269,N_11436);
xor U11650 (N_11650,N_11494,N_11132);
and U11651 (N_11651,N_11266,N_11248);
or U11652 (N_11652,N_11129,N_11011);
nor U11653 (N_11653,N_11403,N_11218);
and U11654 (N_11654,N_11412,N_11421);
xnor U11655 (N_11655,N_11308,N_11176);
nor U11656 (N_11656,N_11288,N_11476);
or U11657 (N_11657,N_11340,N_11144);
nor U11658 (N_11658,N_11166,N_11240);
xor U11659 (N_11659,N_11026,N_11388);
or U11660 (N_11660,N_11441,N_11291);
nor U11661 (N_11661,N_11326,N_11418);
and U11662 (N_11662,N_11228,N_11088);
nor U11663 (N_11663,N_11017,N_11080);
or U11664 (N_11664,N_11246,N_11470);
and U11665 (N_11665,N_11206,N_11465);
and U11666 (N_11666,N_11154,N_11108);
nor U11667 (N_11667,N_11265,N_11350);
and U11668 (N_11668,N_11054,N_11089);
or U11669 (N_11669,N_11462,N_11463);
and U11670 (N_11670,N_11084,N_11304);
or U11671 (N_11671,N_11464,N_11196);
xor U11672 (N_11672,N_11000,N_11145);
nand U11673 (N_11673,N_11296,N_11419);
xnor U11674 (N_11674,N_11381,N_11115);
nor U11675 (N_11675,N_11349,N_11344);
or U11676 (N_11676,N_11090,N_11307);
or U11677 (N_11677,N_11472,N_11194);
xor U11678 (N_11678,N_11083,N_11126);
and U11679 (N_11679,N_11444,N_11480);
or U11680 (N_11680,N_11124,N_11072);
and U11681 (N_11681,N_11471,N_11323);
nand U11682 (N_11682,N_11181,N_11342);
nor U11683 (N_11683,N_11493,N_11302);
nor U11684 (N_11684,N_11076,N_11233);
or U11685 (N_11685,N_11142,N_11482);
xor U11686 (N_11686,N_11128,N_11156);
xnor U11687 (N_11687,N_11443,N_11136);
or U11688 (N_11688,N_11217,N_11335);
or U11689 (N_11689,N_11396,N_11374);
nand U11690 (N_11690,N_11360,N_11175);
xnor U11691 (N_11691,N_11358,N_11347);
xor U11692 (N_11692,N_11404,N_11425);
nor U11693 (N_11693,N_11244,N_11301);
xnor U11694 (N_11694,N_11325,N_11313);
or U11695 (N_11695,N_11277,N_11130);
or U11696 (N_11696,N_11373,N_11392);
nor U11697 (N_11697,N_11070,N_11093);
nand U11698 (N_11698,N_11188,N_11495);
and U11699 (N_11699,N_11268,N_11479);
nor U11700 (N_11700,N_11400,N_11318);
and U11701 (N_11701,N_11370,N_11148);
and U11702 (N_11702,N_11330,N_11283);
xor U11703 (N_11703,N_11157,N_11336);
nand U11704 (N_11704,N_11382,N_11348);
nor U11705 (N_11705,N_11251,N_11389);
xor U11706 (N_11706,N_11306,N_11005);
nand U11707 (N_11707,N_11066,N_11092);
or U11708 (N_11708,N_11473,N_11135);
or U11709 (N_11709,N_11032,N_11012);
nand U11710 (N_11710,N_11118,N_11212);
xor U11711 (N_11711,N_11163,N_11261);
xor U11712 (N_11712,N_11195,N_11235);
nand U11713 (N_11713,N_11239,N_11341);
or U11714 (N_11714,N_11242,N_11353);
nand U11715 (N_11715,N_11272,N_11055);
or U11716 (N_11716,N_11401,N_11297);
and U11717 (N_11717,N_11223,N_11362);
or U11718 (N_11718,N_11329,N_11141);
and U11719 (N_11719,N_11190,N_11103);
nand U11720 (N_11720,N_11110,N_11044);
or U11721 (N_11721,N_11169,N_11167);
xor U11722 (N_11722,N_11486,N_11286);
and U11723 (N_11723,N_11278,N_11177);
xnor U11724 (N_11724,N_11189,N_11171);
nor U11725 (N_11725,N_11060,N_11411);
and U11726 (N_11726,N_11097,N_11282);
xor U11727 (N_11727,N_11003,N_11222);
nor U11728 (N_11728,N_11161,N_11276);
nor U11729 (N_11729,N_11364,N_11322);
nor U11730 (N_11730,N_11105,N_11033);
nor U11731 (N_11731,N_11461,N_11427);
nand U11732 (N_11732,N_11249,N_11138);
nand U11733 (N_11733,N_11314,N_11158);
or U11734 (N_11734,N_11095,N_11448);
or U11735 (N_11735,N_11119,N_11478);
nor U11736 (N_11736,N_11294,N_11442);
and U11737 (N_11737,N_11424,N_11238);
nor U11738 (N_11738,N_11317,N_11213);
and U11739 (N_11739,N_11229,N_11209);
xnor U11740 (N_11740,N_11208,N_11455);
xor U11741 (N_11741,N_11460,N_11215);
nor U11742 (N_11742,N_11298,N_11414);
and U11743 (N_11743,N_11057,N_11376);
and U11744 (N_11744,N_11267,N_11075);
and U11745 (N_11745,N_11008,N_11380);
and U11746 (N_11746,N_11101,N_11316);
and U11747 (N_11747,N_11051,N_11045);
nand U11748 (N_11748,N_11202,N_11221);
or U11749 (N_11749,N_11027,N_11170);
xor U11750 (N_11750,N_11381,N_11101);
or U11751 (N_11751,N_11001,N_11011);
nand U11752 (N_11752,N_11207,N_11260);
and U11753 (N_11753,N_11133,N_11257);
nor U11754 (N_11754,N_11121,N_11413);
nand U11755 (N_11755,N_11071,N_11150);
nand U11756 (N_11756,N_11405,N_11308);
and U11757 (N_11757,N_11004,N_11495);
xor U11758 (N_11758,N_11176,N_11059);
nor U11759 (N_11759,N_11492,N_11397);
nor U11760 (N_11760,N_11167,N_11362);
xor U11761 (N_11761,N_11487,N_11474);
and U11762 (N_11762,N_11055,N_11325);
nand U11763 (N_11763,N_11156,N_11456);
and U11764 (N_11764,N_11461,N_11288);
nor U11765 (N_11765,N_11250,N_11469);
and U11766 (N_11766,N_11175,N_11017);
or U11767 (N_11767,N_11149,N_11089);
nand U11768 (N_11768,N_11041,N_11191);
xor U11769 (N_11769,N_11053,N_11113);
or U11770 (N_11770,N_11006,N_11212);
nand U11771 (N_11771,N_11123,N_11162);
nor U11772 (N_11772,N_11121,N_11054);
nor U11773 (N_11773,N_11373,N_11305);
or U11774 (N_11774,N_11008,N_11131);
or U11775 (N_11775,N_11242,N_11215);
nor U11776 (N_11776,N_11361,N_11261);
nor U11777 (N_11777,N_11048,N_11143);
and U11778 (N_11778,N_11056,N_11275);
nor U11779 (N_11779,N_11117,N_11316);
xnor U11780 (N_11780,N_11146,N_11071);
and U11781 (N_11781,N_11137,N_11348);
xnor U11782 (N_11782,N_11262,N_11337);
nand U11783 (N_11783,N_11047,N_11366);
xor U11784 (N_11784,N_11206,N_11284);
nor U11785 (N_11785,N_11394,N_11396);
xnor U11786 (N_11786,N_11060,N_11195);
xnor U11787 (N_11787,N_11297,N_11058);
nand U11788 (N_11788,N_11327,N_11216);
nand U11789 (N_11789,N_11353,N_11438);
and U11790 (N_11790,N_11378,N_11107);
xnor U11791 (N_11791,N_11303,N_11008);
nor U11792 (N_11792,N_11018,N_11421);
and U11793 (N_11793,N_11123,N_11423);
nand U11794 (N_11794,N_11091,N_11420);
nor U11795 (N_11795,N_11131,N_11465);
xor U11796 (N_11796,N_11370,N_11047);
or U11797 (N_11797,N_11131,N_11066);
nor U11798 (N_11798,N_11471,N_11086);
or U11799 (N_11799,N_11417,N_11189);
nand U11800 (N_11800,N_11084,N_11419);
nor U11801 (N_11801,N_11400,N_11244);
nor U11802 (N_11802,N_11103,N_11258);
and U11803 (N_11803,N_11231,N_11273);
or U11804 (N_11804,N_11274,N_11260);
xnor U11805 (N_11805,N_11236,N_11419);
xor U11806 (N_11806,N_11429,N_11419);
and U11807 (N_11807,N_11239,N_11107);
xor U11808 (N_11808,N_11050,N_11090);
and U11809 (N_11809,N_11410,N_11086);
or U11810 (N_11810,N_11415,N_11100);
nor U11811 (N_11811,N_11382,N_11494);
or U11812 (N_11812,N_11333,N_11220);
xnor U11813 (N_11813,N_11444,N_11212);
xnor U11814 (N_11814,N_11104,N_11253);
nor U11815 (N_11815,N_11274,N_11063);
and U11816 (N_11816,N_11451,N_11266);
and U11817 (N_11817,N_11318,N_11179);
nor U11818 (N_11818,N_11399,N_11450);
and U11819 (N_11819,N_11398,N_11479);
and U11820 (N_11820,N_11462,N_11050);
xnor U11821 (N_11821,N_11033,N_11073);
nor U11822 (N_11822,N_11149,N_11491);
nand U11823 (N_11823,N_11406,N_11218);
xor U11824 (N_11824,N_11203,N_11314);
or U11825 (N_11825,N_11172,N_11387);
or U11826 (N_11826,N_11486,N_11269);
xor U11827 (N_11827,N_11218,N_11134);
nand U11828 (N_11828,N_11266,N_11388);
nand U11829 (N_11829,N_11033,N_11288);
or U11830 (N_11830,N_11372,N_11157);
or U11831 (N_11831,N_11142,N_11484);
and U11832 (N_11832,N_11285,N_11180);
nor U11833 (N_11833,N_11042,N_11201);
and U11834 (N_11834,N_11391,N_11190);
xnor U11835 (N_11835,N_11155,N_11381);
nand U11836 (N_11836,N_11256,N_11113);
or U11837 (N_11837,N_11116,N_11155);
or U11838 (N_11838,N_11140,N_11314);
and U11839 (N_11839,N_11063,N_11082);
nand U11840 (N_11840,N_11149,N_11358);
or U11841 (N_11841,N_11071,N_11302);
and U11842 (N_11842,N_11096,N_11495);
or U11843 (N_11843,N_11348,N_11054);
xnor U11844 (N_11844,N_11416,N_11140);
nand U11845 (N_11845,N_11372,N_11482);
nand U11846 (N_11846,N_11227,N_11173);
and U11847 (N_11847,N_11310,N_11245);
xor U11848 (N_11848,N_11429,N_11437);
and U11849 (N_11849,N_11021,N_11462);
and U11850 (N_11850,N_11136,N_11391);
or U11851 (N_11851,N_11024,N_11154);
and U11852 (N_11852,N_11180,N_11379);
or U11853 (N_11853,N_11273,N_11137);
nor U11854 (N_11854,N_11274,N_11050);
and U11855 (N_11855,N_11283,N_11124);
xor U11856 (N_11856,N_11075,N_11484);
or U11857 (N_11857,N_11282,N_11091);
nor U11858 (N_11858,N_11054,N_11419);
nor U11859 (N_11859,N_11264,N_11397);
nor U11860 (N_11860,N_11359,N_11323);
nand U11861 (N_11861,N_11199,N_11128);
nor U11862 (N_11862,N_11194,N_11142);
or U11863 (N_11863,N_11256,N_11016);
and U11864 (N_11864,N_11138,N_11010);
and U11865 (N_11865,N_11334,N_11390);
and U11866 (N_11866,N_11019,N_11154);
or U11867 (N_11867,N_11333,N_11065);
or U11868 (N_11868,N_11408,N_11230);
or U11869 (N_11869,N_11359,N_11186);
nand U11870 (N_11870,N_11298,N_11345);
and U11871 (N_11871,N_11237,N_11477);
or U11872 (N_11872,N_11178,N_11044);
nand U11873 (N_11873,N_11363,N_11337);
xor U11874 (N_11874,N_11235,N_11220);
xnor U11875 (N_11875,N_11487,N_11105);
xor U11876 (N_11876,N_11242,N_11168);
nor U11877 (N_11877,N_11427,N_11130);
xor U11878 (N_11878,N_11009,N_11104);
nand U11879 (N_11879,N_11043,N_11499);
xor U11880 (N_11880,N_11373,N_11163);
or U11881 (N_11881,N_11013,N_11242);
or U11882 (N_11882,N_11111,N_11456);
xor U11883 (N_11883,N_11074,N_11340);
xor U11884 (N_11884,N_11118,N_11241);
nor U11885 (N_11885,N_11392,N_11437);
and U11886 (N_11886,N_11156,N_11091);
xor U11887 (N_11887,N_11228,N_11358);
or U11888 (N_11888,N_11183,N_11094);
nand U11889 (N_11889,N_11320,N_11286);
and U11890 (N_11890,N_11456,N_11041);
and U11891 (N_11891,N_11465,N_11188);
and U11892 (N_11892,N_11269,N_11390);
and U11893 (N_11893,N_11209,N_11085);
or U11894 (N_11894,N_11109,N_11349);
and U11895 (N_11895,N_11381,N_11044);
xnor U11896 (N_11896,N_11293,N_11415);
nor U11897 (N_11897,N_11368,N_11351);
or U11898 (N_11898,N_11095,N_11457);
nand U11899 (N_11899,N_11169,N_11361);
xnor U11900 (N_11900,N_11118,N_11073);
xor U11901 (N_11901,N_11443,N_11277);
xor U11902 (N_11902,N_11385,N_11323);
xor U11903 (N_11903,N_11049,N_11052);
xor U11904 (N_11904,N_11481,N_11412);
nand U11905 (N_11905,N_11007,N_11124);
nor U11906 (N_11906,N_11450,N_11497);
and U11907 (N_11907,N_11086,N_11061);
nor U11908 (N_11908,N_11475,N_11467);
xor U11909 (N_11909,N_11421,N_11060);
nand U11910 (N_11910,N_11000,N_11321);
xor U11911 (N_11911,N_11051,N_11121);
xnor U11912 (N_11912,N_11219,N_11398);
nor U11913 (N_11913,N_11449,N_11377);
nor U11914 (N_11914,N_11476,N_11442);
or U11915 (N_11915,N_11365,N_11050);
or U11916 (N_11916,N_11427,N_11389);
xor U11917 (N_11917,N_11214,N_11366);
or U11918 (N_11918,N_11034,N_11158);
xor U11919 (N_11919,N_11070,N_11204);
xnor U11920 (N_11920,N_11410,N_11368);
and U11921 (N_11921,N_11130,N_11374);
and U11922 (N_11922,N_11163,N_11181);
or U11923 (N_11923,N_11128,N_11277);
nand U11924 (N_11924,N_11382,N_11007);
xor U11925 (N_11925,N_11314,N_11063);
xnor U11926 (N_11926,N_11470,N_11000);
nor U11927 (N_11927,N_11020,N_11287);
nor U11928 (N_11928,N_11494,N_11376);
and U11929 (N_11929,N_11045,N_11429);
and U11930 (N_11930,N_11094,N_11459);
and U11931 (N_11931,N_11433,N_11304);
xor U11932 (N_11932,N_11118,N_11247);
and U11933 (N_11933,N_11362,N_11405);
nand U11934 (N_11934,N_11190,N_11267);
nand U11935 (N_11935,N_11283,N_11274);
nand U11936 (N_11936,N_11036,N_11099);
xnor U11937 (N_11937,N_11491,N_11215);
xnor U11938 (N_11938,N_11159,N_11140);
nor U11939 (N_11939,N_11318,N_11301);
xnor U11940 (N_11940,N_11281,N_11137);
or U11941 (N_11941,N_11397,N_11192);
nor U11942 (N_11942,N_11178,N_11497);
nand U11943 (N_11943,N_11312,N_11066);
and U11944 (N_11944,N_11333,N_11436);
and U11945 (N_11945,N_11280,N_11458);
or U11946 (N_11946,N_11258,N_11325);
nand U11947 (N_11947,N_11195,N_11464);
nand U11948 (N_11948,N_11047,N_11075);
and U11949 (N_11949,N_11180,N_11134);
and U11950 (N_11950,N_11482,N_11411);
nand U11951 (N_11951,N_11283,N_11355);
nand U11952 (N_11952,N_11193,N_11332);
xnor U11953 (N_11953,N_11104,N_11285);
nand U11954 (N_11954,N_11373,N_11301);
or U11955 (N_11955,N_11499,N_11196);
nand U11956 (N_11956,N_11410,N_11288);
and U11957 (N_11957,N_11064,N_11078);
nor U11958 (N_11958,N_11221,N_11369);
nand U11959 (N_11959,N_11048,N_11331);
xor U11960 (N_11960,N_11247,N_11119);
and U11961 (N_11961,N_11332,N_11275);
and U11962 (N_11962,N_11463,N_11132);
or U11963 (N_11963,N_11140,N_11410);
and U11964 (N_11964,N_11307,N_11248);
and U11965 (N_11965,N_11203,N_11175);
or U11966 (N_11966,N_11024,N_11322);
nor U11967 (N_11967,N_11194,N_11180);
nor U11968 (N_11968,N_11159,N_11270);
or U11969 (N_11969,N_11141,N_11084);
and U11970 (N_11970,N_11298,N_11055);
nand U11971 (N_11971,N_11206,N_11442);
nor U11972 (N_11972,N_11261,N_11064);
nand U11973 (N_11973,N_11267,N_11425);
nand U11974 (N_11974,N_11402,N_11178);
and U11975 (N_11975,N_11145,N_11351);
nor U11976 (N_11976,N_11497,N_11132);
xnor U11977 (N_11977,N_11293,N_11490);
xnor U11978 (N_11978,N_11487,N_11276);
nor U11979 (N_11979,N_11146,N_11407);
and U11980 (N_11980,N_11131,N_11256);
xor U11981 (N_11981,N_11494,N_11000);
nand U11982 (N_11982,N_11073,N_11284);
and U11983 (N_11983,N_11358,N_11452);
and U11984 (N_11984,N_11403,N_11294);
nor U11985 (N_11985,N_11231,N_11023);
xor U11986 (N_11986,N_11460,N_11380);
and U11987 (N_11987,N_11247,N_11200);
xor U11988 (N_11988,N_11330,N_11457);
nor U11989 (N_11989,N_11139,N_11158);
nand U11990 (N_11990,N_11148,N_11265);
nand U11991 (N_11991,N_11273,N_11031);
or U11992 (N_11992,N_11310,N_11119);
and U11993 (N_11993,N_11409,N_11247);
nor U11994 (N_11994,N_11249,N_11231);
and U11995 (N_11995,N_11485,N_11477);
and U11996 (N_11996,N_11018,N_11169);
and U11997 (N_11997,N_11192,N_11323);
or U11998 (N_11998,N_11413,N_11319);
nor U11999 (N_11999,N_11225,N_11283);
xnor U12000 (N_12000,N_11951,N_11549);
nor U12001 (N_12001,N_11758,N_11527);
nand U12002 (N_12002,N_11807,N_11547);
nor U12003 (N_12003,N_11653,N_11755);
nor U12004 (N_12004,N_11710,N_11628);
nor U12005 (N_12005,N_11737,N_11812);
or U12006 (N_12006,N_11963,N_11696);
and U12007 (N_12007,N_11808,N_11919);
xnor U12008 (N_12008,N_11679,N_11955);
nor U12009 (N_12009,N_11872,N_11792);
and U12010 (N_12010,N_11716,N_11833);
or U12011 (N_12011,N_11917,N_11687);
nand U12012 (N_12012,N_11868,N_11957);
nand U12013 (N_12013,N_11797,N_11846);
nor U12014 (N_12014,N_11504,N_11865);
xnor U12015 (N_12015,N_11941,N_11916);
or U12016 (N_12016,N_11510,N_11829);
xor U12017 (N_12017,N_11715,N_11802);
xnor U12018 (N_12018,N_11811,N_11814);
and U12019 (N_12019,N_11761,N_11592);
and U12020 (N_12020,N_11892,N_11555);
or U12021 (N_12021,N_11961,N_11795);
and U12022 (N_12022,N_11933,N_11560);
and U12023 (N_12023,N_11521,N_11890);
and U12024 (N_12024,N_11852,N_11987);
xor U12025 (N_12025,N_11581,N_11967);
nor U12026 (N_12026,N_11702,N_11713);
nand U12027 (N_12027,N_11924,N_11898);
nor U12028 (N_12028,N_11636,N_11566);
nor U12029 (N_12029,N_11650,N_11821);
or U12030 (N_12030,N_11945,N_11763);
nor U12031 (N_12031,N_11670,N_11950);
and U12032 (N_12032,N_11753,N_11966);
xor U12033 (N_12033,N_11762,N_11507);
xor U12034 (N_12034,N_11837,N_11879);
xnor U12035 (N_12035,N_11845,N_11648);
nor U12036 (N_12036,N_11714,N_11739);
nor U12037 (N_12037,N_11783,N_11569);
nand U12038 (N_12038,N_11567,N_11532);
nor U12039 (N_12039,N_11907,N_11631);
nand U12040 (N_12040,N_11883,N_11861);
nor U12041 (N_12041,N_11529,N_11973);
xnor U12042 (N_12042,N_11623,N_11757);
nand U12043 (N_12043,N_11667,N_11836);
or U12044 (N_12044,N_11749,N_11645);
nor U12045 (N_12045,N_11576,N_11748);
or U12046 (N_12046,N_11859,N_11780);
xnor U12047 (N_12047,N_11642,N_11588);
nand U12048 (N_12048,N_11777,N_11663);
nand U12049 (N_12049,N_11585,N_11751);
or U12050 (N_12050,N_11920,N_11596);
nand U12051 (N_12051,N_11732,N_11662);
nand U12052 (N_12052,N_11771,N_11727);
xnor U12053 (N_12053,N_11734,N_11880);
nand U12054 (N_12054,N_11864,N_11982);
and U12055 (N_12055,N_11705,N_11711);
or U12056 (N_12056,N_11994,N_11834);
or U12057 (N_12057,N_11838,N_11577);
and U12058 (N_12058,N_11980,N_11743);
or U12059 (N_12059,N_11523,N_11528);
and U12060 (N_12060,N_11793,N_11736);
nor U12061 (N_12061,N_11826,N_11765);
nand U12062 (N_12062,N_11733,N_11799);
or U12063 (N_12063,N_11551,N_11774);
nand U12064 (N_12064,N_11925,N_11535);
or U12065 (N_12065,N_11773,N_11768);
and U12066 (N_12066,N_11553,N_11508);
and U12067 (N_12067,N_11522,N_11526);
or U12068 (N_12068,N_11629,N_11786);
nand U12069 (N_12069,N_11656,N_11894);
and U12070 (N_12070,N_11700,N_11790);
nor U12071 (N_12071,N_11904,N_11842);
xnor U12072 (N_12072,N_11544,N_11726);
or U12073 (N_12073,N_11841,N_11899);
nor U12074 (N_12074,N_11889,N_11661);
or U12075 (N_12075,N_11689,N_11927);
nor U12076 (N_12076,N_11888,N_11591);
or U12077 (N_12077,N_11813,N_11738);
or U12078 (N_12078,N_11954,N_11693);
xor U12079 (N_12079,N_11608,N_11796);
nand U12080 (N_12080,N_11819,N_11997);
xor U12081 (N_12081,N_11960,N_11568);
nor U12082 (N_12082,N_11622,N_11692);
xor U12083 (N_12083,N_11514,N_11956);
or U12084 (N_12084,N_11723,N_11896);
or U12085 (N_12085,N_11630,N_11988);
nor U12086 (N_12086,N_11534,N_11855);
nand U12087 (N_12087,N_11962,N_11570);
or U12088 (N_12088,N_11647,N_11969);
or U12089 (N_12089,N_11984,N_11775);
nor U12090 (N_12090,N_11926,N_11564);
xnor U12091 (N_12091,N_11978,N_11610);
nor U12092 (N_12092,N_11600,N_11515);
or U12093 (N_12093,N_11539,N_11981);
nor U12094 (N_12094,N_11789,N_11694);
or U12095 (N_12095,N_11858,N_11586);
or U12096 (N_12096,N_11860,N_11906);
or U12097 (N_12097,N_11706,N_11977);
nand U12098 (N_12098,N_11989,N_11659);
xnor U12099 (N_12099,N_11707,N_11519);
xnor U12100 (N_12100,N_11634,N_11557);
xor U12101 (N_12101,N_11719,N_11953);
and U12102 (N_12102,N_11506,N_11875);
and U12103 (N_12103,N_11903,N_11582);
or U12104 (N_12104,N_11923,N_11513);
xnor U12105 (N_12105,N_11905,N_11857);
nand U12106 (N_12106,N_11938,N_11708);
and U12107 (N_12107,N_11990,N_11633);
and U12108 (N_12108,N_11823,N_11545);
xnor U12109 (N_12109,N_11729,N_11558);
nand U12110 (N_12110,N_11878,N_11972);
and U12111 (N_12111,N_11505,N_11844);
xor U12112 (N_12112,N_11541,N_11998);
xnor U12113 (N_12113,N_11788,N_11822);
xor U12114 (N_12114,N_11922,N_11603);
nor U12115 (N_12115,N_11787,N_11500);
nand U12116 (N_12116,N_11512,N_11556);
xnor U12117 (N_12117,N_11816,N_11542);
or U12118 (N_12118,N_11983,N_11625);
nor U12119 (N_12119,N_11717,N_11578);
nand U12120 (N_12120,N_11760,N_11530);
or U12121 (N_12121,N_11818,N_11800);
and U12122 (N_12122,N_11843,N_11537);
or U12123 (N_12123,N_11611,N_11911);
and U12124 (N_12124,N_11887,N_11518);
or U12125 (N_12125,N_11895,N_11583);
and U12126 (N_12126,N_11691,N_11617);
and U12127 (N_12127,N_11563,N_11803);
and U12128 (N_12128,N_11703,N_11654);
nand U12129 (N_12129,N_11604,N_11935);
nor U12130 (N_12130,N_11971,N_11877);
and U12131 (N_12131,N_11674,N_11804);
or U12132 (N_12132,N_11606,N_11718);
and U12133 (N_12133,N_11921,N_11632);
or U12134 (N_12134,N_11735,N_11698);
nor U12135 (N_12135,N_11502,N_11697);
nand U12136 (N_12136,N_11533,N_11942);
nor U12137 (N_12137,N_11828,N_11572);
nand U12138 (N_12138,N_11665,N_11912);
and U12139 (N_12139,N_11785,N_11641);
nor U12140 (N_12140,N_11574,N_11620);
and U12141 (N_12141,N_11619,N_11722);
and U12142 (N_12142,N_11839,N_11747);
or U12143 (N_12143,N_11658,N_11680);
xnor U12144 (N_12144,N_11575,N_11866);
nor U12145 (N_12145,N_11959,N_11893);
xnor U12146 (N_12146,N_11550,N_11546);
xnor U12147 (N_12147,N_11638,N_11985);
and U12148 (N_12148,N_11835,N_11543);
and U12149 (N_12149,N_11536,N_11509);
nor U12150 (N_12150,N_11902,N_11832);
or U12151 (N_12151,N_11759,N_11613);
nor U12152 (N_12152,N_11934,N_11970);
nor U12153 (N_12153,N_11939,N_11750);
nor U12154 (N_12154,N_11810,N_11516);
nand U12155 (N_12155,N_11996,N_11913);
nor U12156 (N_12156,N_11684,N_11851);
nor U12157 (N_12157,N_11579,N_11931);
or U12158 (N_12158,N_11695,N_11740);
xor U12159 (N_12159,N_11699,N_11720);
or U12160 (N_12160,N_11979,N_11815);
and U12161 (N_12161,N_11643,N_11914);
and U12162 (N_12162,N_11652,N_11741);
nor U12163 (N_12163,N_11686,N_11856);
or U12164 (N_12164,N_11964,N_11712);
and U12165 (N_12165,N_11637,N_11940);
nor U12166 (N_12166,N_11615,N_11986);
nand U12167 (N_12167,N_11772,N_11624);
nor U12168 (N_12168,N_11791,N_11639);
or U12169 (N_12169,N_11874,N_11809);
xnor U12170 (N_12170,N_11976,N_11820);
xnor U12171 (N_12171,N_11936,N_11669);
or U12172 (N_12172,N_11850,N_11649);
and U12173 (N_12173,N_11730,N_11602);
nand U12174 (N_12174,N_11779,N_11869);
nand U12175 (N_12175,N_11531,N_11766);
or U12176 (N_12176,N_11830,N_11690);
and U12177 (N_12177,N_11618,N_11672);
nor U12178 (N_12178,N_11794,N_11995);
nand U12179 (N_12179,N_11863,N_11752);
nor U12180 (N_12180,N_11881,N_11784);
xor U12181 (N_12181,N_11937,N_11520);
nor U12182 (N_12182,N_11848,N_11552);
and U12183 (N_12183,N_11511,N_11798);
nor U12184 (N_12184,N_11817,N_11503);
or U12185 (N_12185,N_11781,N_11559);
nor U12186 (N_12186,N_11805,N_11947);
nand U12187 (N_12187,N_11580,N_11876);
and U12188 (N_12188,N_11548,N_11946);
nand U12189 (N_12189,N_11900,N_11673);
xor U12190 (N_12190,N_11824,N_11958);
and U12191 (N_12191,N_11664,N_11616);
nand U12192 (N_12192,N_11948,N_11677);
nand U12193 (N_12193,N_11932,N_11873);
xor U12194 (N_12194,N_11671,N_11721);
nor U12195 (N_12195,N_11965,N_11968);
or U12196 (N_12196,N_11646,N_11746);
nor U12197 (N_12197,N_11884,N_11992);
nor U12198 (N_12198,N_11908,N_11778);
xor U12199 (N_12199,N_11909,N_11867);
and U12200 (N_12200,N_11949,N_11597);
or U12201 (N_12201,N_11593,N_11882);
and U12202 (N_12202,N_11517,N_11745);
and U12203 (N_12203,N_11525,N_11840);
and U12204 (N_12204,N_11704,N_11993);
xnor U12205 (N_12205,N_11767,N_11827);
nand U12206 (N_12206,N_11655,N_11657);
or U12207 (N_12207,N_11501,N_11621);
xor U12208 (N_12208,N_11554,N_11930);
xor U12209 (N_12209,N_11886,N_11540);
nor U12210 (N_12210,N_11871,N_11589);
nand U12211 (N_12211,N_11682,N_11609);
nand U12212 (N_12212,N_11991,N_11668);
or U12213 (N_12213,N_11782,N_11952);
or U12214 (N_12214,N_11599,N_11731);
nand U12215 (N_12215,N_11885,N_11929);
or U12216 (N_12216,N_11862,N_11915);
xor U12217 (N_12217,N_11605,N_11897);
and U12218 (N_12218,N_11614,N_11565);
nand U12219 (N_12219,N_11849,N_11644);
nand U12220 (N_12220,N_11831,N_11601);
or U12221 (N_12221,N_11944,N_11561);
xor U12222 (N_12222,N_11584,N_11776);
nand U12223 (N_12223,N_11678,N_11675);
xnor U12224 (N_12224,N_11769,N_11891);
nor U12225 (N_12225,N_11901,N_11627);
nand U12226 (N_12226,N_11688,N_11573);
and U12227 (N_12227,N_11854,N_11651);
nand U12228 (N_12228,N_11742,N_11562);
and U12229 (N_12229,N_11756,N_11928);
and U12230 (N_12230,N_11612,N_11975);
or U12231 (N_12231,N_11744,N_11870);
and U12232 (N_12232,N_11770,N_11595);
or U12233 (N_12233,N_11594,N_11709);
or U12234 (N_12234,N_11635,N_11999);
and U12235 (N_12235,N_11701,N_11681);
nand U12236 (N_12236,N_11725,N_11538);
nor U12237 (N_12237,N_11666,N_11728);
xor U12238 (N_12238,N_11943,N_11626);
nand U12239 (N_12239,N_11853,N_11764);
nor U12240 (N_12240,N_11587,N_11754);
nand U12241 (N_12241,N_11683,N_11974);
nand U12242 (N_12242,N_11847,N_11660);
nor U12243 (N_12243,N_11524,N_11685);
and U12244 (N_12244,N_11676,N_11806);
and U12245 (N_12245,N_11590,N_11724);
or U12246 (N_12246,N_11801,N_11825);
and U12247 (N_12247,N_11918,N_11640);
nand U12248 (N_12248,N_11910,N_11607);
nor U12249 (N_12249,N_11598,N_11571);
nand U12250 (N_12250,N_11808,N_11984);
or U12251 (N_12251,N_11580,N_11913);
nor U12252 (N_12252,N_11574,N_11878);
and U12253 (N_12253,N_11775,N_11689);
or U12254 (N_12254,N_11914,N_11997);
xnor U12255 (N_12255,N_11854,N_11767);
nor U12256 (N_12256,N_11838,N_11872);
xnor U12257 (N_12257,N_11750,N_11793);
nand U12258 (N_12258,N_11680,N_11638);
and U12259 (N_12259,N_11584,N_11697);
and U12260 (N_12260,N_11790,N_11847);
and U12261 (N_12261,N_11603,N_11718);
nand U12262 (N_12262,N_11771,N_11976);
nor U12263 (N_12263,N_11995,N_11846);
nand U12264 (N_12264,N_11971,N_11535);
or U12265 (N_12265,N_11832,N_11912);
nor U12266 (N_12266,N_11552,N_11761);
nor U12267 (N_12267,N_11630,N_11546);
nand U12268 (N_12268,N_11553,N_11875);
or U12269 (N_12269,N_11679,N_11961);
nor U12270 (N_12270,N_11794,N_11627);
nor U12271 (N_12271,N_11958,N_11975);
and U12272 (N_12272,N_11721,N_11584);
and U12273 (N_12273,N_11609,N_11543);
nand U12274 (N_12274,N_11677,N_11859);
and U12275 (N_12275,N_11865,N_11660);
xor U12276 (N_12276,N_11619,N_11506);
nor U12277 (N_12277,N_11555,N_11685);
or U12278 (N_12278,N_11852,N_11680);
nor U12279 (N_12279,N_11989,N_11766);
or U12280 (N_12280,N_11933,N_11731);
nand U12281 (N_12281,N_11943,N_11953);
nand U12282 (N_12282,N_11921,N_11812);
nor U12283 (N_12283,N_11662,N_11783);
or U12284 (N_12284,N_11804,N_11976);
or U12285 (N_12285,N_11618,N_11632);
and U12286 (N_12286,N_11542,N_11973);
or U12287 (N_12287,N_11640,N_11905);
nand U12288 (N_12288,N_11806,N_11757);
nand U12289 (N_12289,N_11669,N_11580);
nand U12290 (N_12290,N_11637,N_11782);
and U12291 (N_12291,N_11712,N_11542);
nand U12292 (N_12292,N_11905,N_11500);
nor U12293 (N_12293,N_11761,N_11528);
nor U12294 (N_12294,N_11932,N_11517);
and U12295 (N_12295,N_11995,N_11984);
or U12296 (N_12296,N_11707,N_11634);
nor U12297 (N_12297,N_11702,N_11949);
nor U12298 (N_12298,N_11516,N_11729);
or U12299 (N_12299,N_11589,N_11965);
xnor U12300 (N_12300,N_11889,N_11893);
or U12301 (N_12301,N_11818,N_11748);
nor U12302 (N_12302,N_11693,N_11948);
or U12303 (N_12303,N_11956,N_11926);
nand U12304 (N_12304,N_11715,N_11550);
and U12305 (N_12305,N_11828,N_11650);
and U12306 (N_12306,N_11572,N_11771);
xor U12307 (N_12307,N_11654,N_11691);
and U12308 (N_12308,N_11533,N_11654);
and U12309 (N_12309,N_11705,N_11535);
or U12310 (N_12310,N_11952,N_11850);
or U12311 (N_12311,N_11715,N_11778);
nor U12312 (N_12312,N_11547,N_11718);
nor U12313 (N_12313,N_11879,N_11501);
nand U12314 (N_12314,N_11970,N_11614);
nor U12315 (N_12315,N_11593,N_11570);
xor U12316 (N_12316,N_11532,N_11658);
and U12317 (N_12317,N_11631,N_11818);
nand U12318 (N_12318,N_11675,N_11862);
xor U12319 (N_12319,N_11526,N_11985);
or U12320 (N_12320,N_11717,N_11740);
nor U12321 (N_12321,N_11651,N_11764);
nor U12322 (N_12322,N_11546,N_11645);
nor U12323 (N_12323,N_11842,N_11629);
nor U12324 (N_12324,N_11991,N_11586);
nand U12325 (N_12325,N_11612,N_11621);
nor U12326 (N_12326,N_11860,N_11707);
xor U12327 (N_12327,N_11808,N_11816);
or U12328 (N_12328,N_11633,N_11586);
xnor U12329 (N_12329,N_11545,N_11804);
nor U12330 (N_12330,N_11597,N_11718);
nor U12331 (N_12331,N_11823,N_11640);
or U12332 (N_12332,N_11924,N_11819);
xor U12333 (N_12333,N_11890,N_11949);
and U12334 (N_12334,N_11854,N_11716);
and U12335 (N_12335,N_11861,N_11871);
and U12336 (N_12336,N_11858,N_11961);
and U12337 (N_12337,N_11518,N_11903);
or U12338 (N_12338,N_11937,N_11948);
nor U12339 (N_12339,N_11736,N_11879);
xnor U12340 (N_12340,N_11695,N_11633);
xnor U12341 (N_12341,N_11958,N_11943);
or U12342 (N_12342,N_11705,N_11679);
nand U12343 (N_12343,N_11821,N_11625);
nor U12344 (N_12344,N_11708,N_11842);
and U12345 (N_12345,N_11700,N_11932);
nor U12346 (N_12346,N_11883,N_11813);
nor U12347 (N_12347,N_11708,N_11779);
and U12348 (N_12348,N_11691,N_11511);
xnor U12349 (N_12349,N_11577,N_11702);
and U12350 (N_12350,N_11663,N_11781);
or U12351 (N_12351,N_11650,N_11544);
nor U12352 (N_12352,N_11539,N_11590);
xnor U12353 (N_12353,N_11691,N_11712);
and U12354 (N_12354,N_11676,N_11881);
nor U12355 (N_12355,N_11503,N_11840);
xnor U12356 (N_12356,N_11563,N_11740);
nand U12357 (N_12357,N_11826,N_11663);
nand U12358 (N_12358,N_11693,N_11830);
xor U12359 (N_12359,N_11698,N_11815);
nor U12360 (N_12360,N_11599,N_11761);
xor U12361 (N_12361,N_11872,N_11935);
nor U12362 (N_12362,N_11584,N_11560);
nor U12363 (N_12363,N_11535,N_11632);
nor U12364 (N_12364,N_11744,N_11807);
xnor U12365 (N_12365,N_11782,N_11745);
xor U12366 (N_12366,N_11627,N_11874);
or U12367 (N_12367,N_11951,N_11511);
nor U12368 (N_12368,N_11885,N_11735);
nand U12369 (N_12369,N_11963,N_11991);
nor U12370 (N_12370,N_11568,N_11599);
or U12371 (N_12371,N_11809,N_11545);
nor U12372 (N_12372,N_11940,N_11620);
nand U12373 (N_12373,N_11647,N_11984);
nand U12374 (N_12374,N_11819,N_11689);
nor U12375 (N_12375,N_11662,N_11849);
nor U12376 (N_12376,N_11501,N_11945);
nand U12377 (N_12377,N_11947,N_11869);
xnor U12378 (N_12378,N_11844,N_11922);
and U12379 (N_12379,N_11737,N_11855);
or U12380 (N_12380,N_11625,N_11799);
nor U12381 (N_12381,N_11600,N_11586);
nor U12382 (N_12382,N_11545,N_11753);
xor U12383 (N_12383,N_11607,N_11696);
and U12384 (N_12384,N_11773,N_11891);
and U12385 (N_12385,N_11507,N_11755);
or U12386 (N_12386,N_11600,N_11730);
and U12387 (N_12387,N_11896,N_11948);
nand U12388 (N_12388,N_11935,N_11564);
xor U12389 (N_12389,N_11570,N_11744);
nor U12390 (N_12390,N_11675,N_11543);
and U12391 (N_12391,N_11756,N_11949);
nand U12392 (N_12392,N_11750,N_11506);
or U12393 (N_12393,N_11657,N_11667);
nor U12394 (N_12394,N_11639,N_11562);
and U12395 (N_12395,N_11621,N_11685);
or U12396 (N_12396,N_11578,N_11649);
nor U12397 (N_12397,N_11888,N_11812);
and U12398 (N_12398,N_11766,N_11887);
xnor U12399 (N_12399,N_11879,N_11982);
and U12400 (N_12400,N_11767,N_11832);
nand U12401 (N_12401,N_11938,N_11574);
nor U12402 (N_12402,N_11753,N_11810);
nand U12403 (N_12403,N_11590,N_11809);
nor U12404 (N_12404,N_11932,N_11977);
or U12405 (N_12405,N_11857,N_11841);
and U12406 (N_12406,N_11787,N_11723);
nand U12407 (N_12407,N_11507,N_11615);
and U12408 (N_12408,N_11631,N_11618);
nand U12409 (N_12409,N_11850,N_11788);
or U12410 (N_12410,N_11841,N_11571);
nand U12411 (N_12411,N_11808,N_11648);
nor U12412 (N_12412,N_11528,N_11667);
and U12413 (N_12413,N_11814,N_11973);
and U12414 (N_12414,N_11534,N_11758);
xnor U12415 (N_12415,N_11643,N_11569);
nand U12416 (N_12416,N_11872,N_11937);
or U12417 (N_12417,N_11719,N_11579);
xor U12418 (N_12418,N_11891,N_11803);
nor U12419 (N_12419,N_11537,N_11849);
xor U12420 (N_12420,N_11577,N_11544);
xor U12421 (N_12421,N_11944,N_11886);
and U12422 (N_12422,N_11900,N_11530);
and U12423 (N_12423,N_11980,N_11588);
or U12424 (N_12424,N_11535,N_11541);
and U12425 (N_12425,N_11640,N_11993);
xor U12426 (N_12426,N_11680,N_11822);
nor U12427 (N_12427,N_11752,N_11837);
nand U12428 (N_12428,N_11652,N_11928);
and U12429 (N_12429,N_11521,N_11598);
nand U12430 (N_12430,N_11827,N_11699);
nor U12431 (N_12431,N_11842,N_11501);
nand U12432 (N_12432,N_11947,N_11566);
nand U12433 (N_12433,N_11670,N_11805);
nand U12434 (N_12434,N_11554,N_11694);
nand U12435 (N_12435,N_11927,N_11813);
xnor U12436 (N_12436,N_11695,N_11978);
nor U12437 (N_12437,N_11894,N_11936);
or U12438 (N_12438,N_11978,N_11859);
or U12439 (N_12439,N_11656,N_11869);
or U12440 (N_12440,N_11729,N_11941);
xnor U12441 (N_12441,N_11851,N_11508);
xnor U12442 (N_12442,N_11685,N_11744);
nand U12443 (N_12443,N_11556,N_11513);
xnor U12444 (N_12444,N_11953,N_11765);
and U12445 (N_12445,N_11922,N_11642);
nor U12446 (N_12446,N_11842,N_11766);
xor U12447 (N_12447,N_11602,N_11804);
or U12448 (N_12448,N_11718,N_11948);
or U12449 (N_12449,N_11878,N_11862);
nor U12450 (N_12450,N_11854,N_11880);
and U12451 (N_12451,N_11596,N_11504);
or U12452 (N_12452,N_11543,N_11562);
nand U12453 (N_12453,N_11716,N_11914);
nand U12454 (N_12454,N_11946,N_11687);
nor U12455 (N_12455,N_11514,N_11926);
nor U12456 (N_12456,N_11790,N_11932);
nor U12457 (N_12457,N_11674,N_11735);
and U12458 (N_12458,N_11617,N_11758);
and U12459 (N_12459,N_11721,N_11800);
nor U12460 (N_12460,N_11919,N_11816);
or U12461 (N_12461,N_11553,N_11971);
or U12462 (N_12462,N_11779,N_11680);
xor U12463 (N_12463,N_11793,N_11672);
nand U12464 (N_12464,N_11863,N_11585);
or U12465 (N_12465,N_11904,N_11710);
nand U12466 (N_12466,N_11715,N_11812);
nor U12467 (N_12467,N_11910,N_11583);
or U12468 (N_12468,N_11504,N_11672);
nor U12469 (N_12469,N_11676,N_11897);
and U12470 (N_12470,N_11899,N_11837);
nand U12471 (N_12471,N_11500,N_11929);
and U12472 (N_12472,N_11700,N_11639);
nor U12473 (N_12473,N_11826,N_11539);
nor U12474 (N_12474,N_11746,N_11959);
nand U12475 (N_12475,N_11518,N_11610);
nor U12476 (N_12476,N_11837,N_11617);
nand U12477 (N_12477,N_11980,N_11715);
nand U12478 (N_12478,N_11944,N_11814);
or U12479 (N_12479,N_11855,N_11649);
xnor U12480 (N_12480,N_11651,N_11644);
nor U12481 (N_12481,N_11747,N_11865);
nand U12482 (N_12482,N_11983,N_11659);
nand U12483 (N_12483,N_11785,N_11751);
or U12484 (N_12484,N_11943,N_11720);
xor U12485 (N_12485,N_11672,N_11908);
xor U12486 (N_12486,N_11678,N_11562);
or U12487 (N_12487,N_11719,N_11844);
nor U12488 (N_12488,N_11970,N_11894);
nand U12489 (N_12489,N_11635,N_11543);
xor U12490 (N_12490,N_11550,N_11669);
nand U12491 (N_12491,N_11969,N_11575);
nand U12492 (N_12492,N_11599,N_11777);
and U12493 (N_12493,N_11868,N_11840);
or U12494 (N_12494,N_11757,N_11824);
or U12495 (N_12495,N_11683,N_11827);
nand U12496 (N_12496,N_11782,N_11552);
nand U12497 (N_12497,N_11774,N_11659);
and U12498 (N_12498,N_11814,N_11504);
xnor U12499 (N_12499,N_11784,N_11709);
xor U12500 (N_12500,N_12089,N_12231);
or U12501 (N_12501,N_12107,N_12250);
and U12502 (N_12502,N_12312,N_12292);
xnor U12503 (N_12503,N_12417,N_12409);
nand U12504 (N_12504,N_12192,N_12196);
nand U12505 (N_12505,N_12449,N_12149);
nor U12506 (N_12506,N_12368,N_12461);
or U12507 (N_12507,N_12220,N_12392);
xnor U12508 (N_12508,N_12337,N_12363);
and U12509 (N_12509,N_12353,N_12229);
and U12510 (N_12510,N_12094,N_12162);
nor U12511 (N_12511,N_12009,N_12328);
nand U12512 (N_12512,N_12139,N_12140);
nand U12513 (N_12513,N_12418,N_12232);
nand U12514 (N_12514,N_12460,N_12233);
and U12515 (N_12515,N_12433,N_12013);
xor U12516 (N_12516,N_12097,N_12186);
nand U12517 (N_12517,N_12100,N_12058);
or U12518 (N_12518,N_12123,N_12226);
and U12519 (N_12519,N_12334,N_12432);
nand U12520 (N_12520,N_12429,N_12281);
or U12521 (N_12521,N_12258,N_12434);
nand U12522 (N_12522,N_12470,N_12238);
nand U12523 (N_12523,N_12468,N_12003);
and U12524 (N_12524,N_12038,N_12126);
xor U12525 (N_12525,N_12357,N_12419);
or U12526 (N_12526,N_12266,N_12129);
nor U12527 (N_12527,N_12069,N_12227);
nor U12528 (N_12528,N_12318,N_12336);
xnor U12529 (N_12529,N_12093,N_12424);
nand U12530 (N_12530,N_12218,N_12222);
xor U12531 (N_12531,N_12067,N_12396);
or U12532 (N_12532,N_12382,N_12488);
xnor U12533 (N_12533,N_12316,N_12447);
or U12534 (N_12534,N_12381,N_12207);
or U12535 (N_12535,N_12402,N_12020);
and U12536 (N_12536,N_12413,N_12237);
nand U12537 (N_12537,N_12469,N_12050);
xor U12538 (N_12538,N_12480,N_12303);
nand U12539 (N_12539,N_12319,N_12389);
and U12540 (N_12540,N_12298,N_12344);
nand U12541 (N_12541,N_12407,N_12133);
nand U12542 (N_12542,N_12053,N_12311);
nor U12543 (N_12543,N_12172,N_12484);
or U12544 (N_12544,N_12446,N_12057);
nor U12545 (N_12545,N_12113,N_12411);
nor U12546 (N_12546,N_12309,N_12314);
xnor U12547 (N_12547,N_12205,N_12261);
nand U12548 (N_12548,N_12387,N_12153);
nand U12549 (N_12549,N_12335,N_12265);
nor U12550 (N_12550,N_12170,N_12457);
and U12551 (N_12551,N_12166,N_12048);
or U12552 (N_12552,N_12324,N_12206);
and U12553 (N_12553,N_12304,N_12277);
xnor U12554 (N_12554,N_12280,N_12428);
and U12555 (N_12555,N_12364,N_12359);
or U12556 (N_12556,N_12412,N_12084);
nor U12557 (N_12557,N_12142,N_12037);
or U12558 (N_12558,N_12085,N_12014);
nor U12559 (N_12559,N_12184,N_12251);
nand U12560 (N_12560,N_12492,N_12150);
and U12561 (N_12561,N_12090,N_12061);
nor U12562 (N_12562,N_12071,N_12269);
nor U12563 (N_12563,N_12175,N_12098);
or U12564 (N_12564,N_12493,N_12242);
xor U12565 (N_12565,N_12030,N_12305);
xnor U12566 (N_12566,N_12439,N_12465);
xor U12567 (N_12567,N_12235,N_12438);
xor U12568 (N_12568,N_12494,N_12390);
nand U12569 (N_12569,N_12183,N_12145);
or U12570 (N_12570,N_12330,N_12224);
and U12571 (N_12571,N_12295,N_12036);
xor U12572 (N_12572,N_12462,N_12474);
nor U12573 (N_12573,N_12477,N_12262);
and U12574 (N_12574,N_12210,N_12383);
nand U12575 (N_12575,N_12105,N_12119);
or U12576 (N_12576,N_12391,N_12486);
nor U12577 (N_12577,N_12329,N_12195);
nor U12578 (N_12578,N_12120,N_12137);
nor U12579 (N_12579,N_12035,N_12406);
nand U12580 (N_12580,N_12127,N_12108);
xor U12581 (N_12581,N_12293,N_12342);
nand U12582 (N_12582,N_12082,N_12083);
nor U12583 (N_12583,N_12249,N_12467);
and U12584 (N_12584,N_12495,N_12187);
and U12585 (N_12585,N_12369,N_12333);
xnor U12586 (N_12586,N_12349,N_12306);
or U12587 (N_12587,N_12112,N_12482);
or U12588 (N_12588,N_12033,N_12178);
nor U12589 (N_12589,N_12109,N_12209);
nor U12590 (N_12590,N_12146,N_12135);
nand U12591 (N_12591,N_12259,N_12095);
nand U12592 (N_12592,N_12204,N_12450);
nor U12593 (N_12593,N_12271,N_12288);
nand U12594 (N_12594,N_12346,N_12499);
nand U12595 (N_12595,N_12156,N_12475);
xor U12596 (N_12596,N_12198,N_12267);
nand U12597 (N_12597,N_12386,N_12323);
or U12598 (N_12598,N_12018,N_12039);
and U12599 (N_12599,N_12115,N_12217);
nor U12600 (N_12600,N_12138,N_12077);
nor U12601 (N_12601,N_12017,N_12032);
and U12602 (N_12602,N_12375,N_12315);
and U12603 (N_12603,N_12004,N_12169);
and U12604 (N_12604,N_12310,N_12110);
or U12605 (N_12605,N_12173,N_12455);
or U12606 (N_12606,N_12430,N_12221);
nor U12607 (N_12607,N_12471,N_12044);
and U12608 (N_12608,N_12283,N_12078);
nor U12609 (N_12609,N_12106,N_12352);
and U12610 (N_12610,N_12415,N_12163);
and U12611 (N_12611,N_12144,N_12385);
xnor U12612 (N_12612,N_12174,N_12476);
nor U12613 (N_12613,N_12131,N_12074);
and U12614 (N_12614,N_12241,N_12022);
xnor U12615 (N_12615,N_12219,N_12079);
nand U12616 (N_12616,N_12479,N_12168);
nor U12617 (N_12617,N_12028,N_12076);
nor U12618 (N_12618,N_12422,N_12148);
nor U12619 (N_12619,N_12073,N_12308);
or U12620 (N_12620,N_12473,N_12070);
and U12621 (N_12621,N_12245,N_12463);
or U12622 (N_12622,N_12301,N_12092);
nand U12623 (N_12623,N_12208,N_12299);
nand U12624 (N_12624,N_12377,N_12254);
or U12625 (N_12625,N_12102,N_12435);
and U12626 (N_12626,N_12374,N_12286);
nor U12627 (N_12627,N_12361,N_12257);
nand U12628 (N_12628,N_12440,N_12203);
or U12629 (N_12629,N_12481,N_12290);
and U12630 (N_12630,N_12317,N_12404);
xnor U12631 (N_12631,N_12045,N_12001);
nor U12632 (N_12632,N_12136,N_12080);
or U12633 (N_12633,N_12040,N_12398);
nor U12634 (N_12634,N_12459,N_12051);
nand U12635 (N_12635,N_12284,N_12046);
or U12636 (N_12636,N_12025,N_12021);
xnor U12637 (N_12637,N_12274,N_12380);
or U12638 (N_12638,N_12152,N_12285);
or U12639 (N_12639,N_12483,N_12397);
or U12640 (N_12640,N_12452,N_12190);
and U12641 (N_12641,N_12176,N_12427);
or U12642 (N_12642,N_12270,N_12276);
nand U12643 (N_12643,N_12244,N_12448);
and U12644 (N_12644,N_12068,N_12322);
and U12645 (N_12645,N_12236,N_12031);
or U12646 (N_12646,N_12049,N_12372);
nand U12647 (N_12647,N_12185,N_12130);
nand U12648 (N_12648,N_12200,N_12015);
and U12649 (N_12649,N_12487,N_12075);
nand U12650 (N_12650,N_12279,N_12060);
and U12651 (N_12651,N_12191,N_12012);
and U12652 (N_12652,N_12088,N_12117);
and U12653 (N_12653,N_12275,N_12408);
xor U12654 (N_12654,N_12348,N_12215);
and U12655 (N_12655,N_12072,N_12326);
nand U12656 (N_12656,N_12000,N_12472);
and U12657 (N_12657,N_12291,N_12167);
or U12658 (N_12658,N_12201,N_12054);
nor U12659 (N_12659,N_12064,N_12410);
xnor U12660 (N_12660,N_12273,N_12423);
nand U12661 (N_12661,N_12216,N_12300);
nor U12662 (N_12662,N_12052,N_12345);
nand U12663 (N_12663,N_12122,N_12320);
nor U12664 (N_12664,N_12491,N_12395);
nand U12665 (N_12665,N_12151,N_12338);
or U12666 (N_12666,N_12260,N_12376);
or U12667 (N_12667,N_12347,N_12096);
xor U12668 (N_12668,N_12453,N_12490);
and U12669 (N_12669,N_12181,N_12425);
nand U12670 (N_12670,N_12008,N_12340);
nor U12671 (N_12671,N_12059,N_12087);
or U12672 (N_12672,N_12128,N_12091);
and U12673 (N_12673,N_12247,N_12321);
xor U12674 (N_12674,N_12379,N_12199);
nor U12675 (N_12675,N_12367,N_12023);
or U12676 (N_12676,N_12124,N_12441);
or U12677 (N_12677,N_12444,N_12354);
nor U12678 (N_12678,N_12339,N_12263);
and U12679 (N_12679,N_12225,N_12062);
and U12680 (N_12680,N_12116,N_12211);
nor U12681 (N_12681,N_12055,N_12327);
and U12682 (N_12682,N_12043,N_12213);
xor U12683 (N_12683,N_12026,N_12005);
nand U12684 (N_12684,N_12313,N_12405);
nor U12685 (N_12685,N_12464,N_12498);
xnor U12686 (N_12686,N_12373,N_12081);
nand U12687 (N_12687,N_12370,N_12442);
nor U12688 (N_12688,N_12268,N_12193);
xnor U12689 (N_12689,N_12234,N_12399);
nor U12690 (N_12690,N_12302,N_12240);
nand U12691 (N_12691,N_12401,N_12437);
nand U12692 (N_12692,N_12256,N_12016);
xor U12693 (N_12693,N_12350,N_12065);
or U12694 (N_12694,N_12388,N_12164);
or U12695 (N_12695,N_12223,N_12165);
nand U12696 (N_12696,N_12157,N_12027);
and U12697 (N_12697,N_12378,N_12443);
and U12698 (N_12698,N_12414,N_12159);
nand U12699 (N_12699,N_12458,N_12066);
nor U12700 (N_12700,N_12239,N_12099);
nor U12701 (N_12701,N_12197,N_12485);
and U12702 (N_12702,N_12114,N_12202);
xor U12703 (N_12703,N_12147,N_12325);
xor U12704 (N_12704,N_12047,N_12182);
nand U12705 (N_12705,N_12264,N_12154);
nand U12706 (N_12706,N_12171,N_12282);
or U12707 (N_12707,N_12189,N_12118);
and U12708 (N_12708,N_12466,N_12394);
xor U12709 (N_12709,N_12436,N_12421);
or U12710 (N_12710,N_12177,N_12497);
xnor U12711 (N_12711,N_12143,N_12362);
nand U12712 (N_12712,N_12111,N_12253);
xor U12713 (N_12713,N_12356,N_12451);
nand U12714 (N_12714,N_12358,N_12002);
and U12715 (N_12715,N_12307,N_12416);
nand U12716 (N_12716,N_12214,N_12180);
nor U12717 (N_12717,N_12029,N_12041);
xnor U12718 (N_12718,N_12331,N_12296);
nand U12719 (N_12719,N_12341,N_12034);
or U12720 (N_12720,N_12431,N_12355);
or U12721 (N_12721,N_12006,N_12252);
nand U12722 (N_12722,N_12212,N_12024);
and U12723 (N_12723,N_12141,N_12393);
nor U12724 (N_12724,N_12351,N_12243);
nor U12725 (N_12725,N_12426,N_12297);
nor U12726 (N_12726,N_12161,N_12019);
xnor U12727 (N_12727,N_12332,N_12121);
or U12728 (N_12728,N_12011,N_12366);
nor U12729 (N_12729,N_12160,N_12400);
and U12730 (N_12730,N_12155,N_12158);
or U12731 (N_12731,N_12228,N_12125);
xnor U12732 (N_12732,N_12179,N_12194);
nor U12733 (N_12733,N_12056,N_12343);
nor U12734 (N_12734,N_12132,N_12042);
or U12735 (N_12735,N_12489,N_12384);
nor U12736 (N_12736,N_12360,N_12101);
or U12737 (N_12737,N_12188,N_12230);
xnor U12738 (N_12738,N_12294,N_12010);
and U12739 (N_12739,N_12086,N_12278);
and U12740 (N_12740,N_12365,N_12496);
or U12741 (N_12741,N_12272,N_12255);
or U12742 (N_12742,N_12403,N_12063);
nand U12743 (N_12743,N_12287,N_12248);
and U12744 (N_12744,N_12454,N_12103);
nand U12745 (N_12745,N_12007,N_12104);
or U12746 (N_12746,N_12420,N_12445);
xnor U12747 (N_12747,N_12371,N_12134);
nand U12748 (N_12748,N_12456,N_12478);
and U12749 (N_12749,N_12246,N_12289);
nand U12750 (N_12750,N_12117,N_12308);
xor U12751 (N_12751,N_12260,N_12320);
xor U12752 (N_12752,N_12415,N_12272);
nand U12753 (N_12753,N_12418,N_12137);
or U12754 (N_12754,N_12044,N_12061);
and U12755 (N_12755,N_12258,N_12356);
and U12756 (N_12756,N_12090,N_12327);
nand U12757 (N_12757,N_12061,N_12299);
nor U12758 (N_12758,N_12035,N_12486);
xor U12759 (N_12759,N_12309,N_12353);
or U12760 (N_12760,N_12362,N_12412);
and U12761 (N_12761,N_12325,N_12005);
and U12762 (N_12762,N_12455,N_12112);
xor U12763 (N_12763,N_12291,N_12158);
xor U12764 (N_12764,N_12259,N_12129);
nor U12765 (N_12765,N_12392,N_12196);
and U12766 (N_12766,N_12311,N_12484);
nand U12767 (N_12767,N_12387,N_12359);
nor U12768 (N_12768,N_12272,N_12151);
or U12769 (N_12769,N_12108,N_12073);
xor U12770 (N_12770,N_12326,N_12156);
nor U12771 (N_12771,N_12086,N_12003);
xor U12772 (N_12772,N_12137,N_12074);
nand U12773 (N_12773,N_12183,N_12181);
xnor U12774 (N_12774,N_12073,N_12357);
nand U12775 (N_12775,N_12195,N_12447);
nand U12776 (N_12776,N_12258,N_12029);
nand U12777 (N_12777,N_12029,N_12489);
nand U12778 (N_12778,N_12393,N_12423);
and U12779 (N_12779,N_12182,N_12317);
or U12780 (N_12780,N_12124,N_12425);
or U12781 (N_12781,N_12249,N_12321);
or U12782 (N_12782,N_12482,N_12305);
or U12783 (N_12783,N_12287,N_12212);
nor U12784 (N_12784,N_12091,N_12338);
xnor U12785 (N_12785,N_12130,N_12445);
xnor U12786 (N_12786,N_12337,N_12351);
nor U12787 (N_12787,N_12050,N_12339);
nor U12788 (N_12788,N_12017,N_12126);
or U12789 (N_12789,N_12251,N_12476);
nor U12790 (N_12790,N_12461,N_12456);
and U12791 (N_12791,N_12396,N_12227);
nand U12792 (N_12792,N_12299,N_12183);
xor U12793 (N_12793,N_12293,N_12308);
or U12794 (N_12794,N_12054,N_12349);
nor U12795 (N_12795,N_12002,N_12396);
nand U12796 (N_12796,N_12486,N_12197);
nand U12797 (N_12797,N_12367,N_12469);
nor U12798 (N_12798,N_12004,N_12022);
nand U12799 (N_12799,N_12335,N_12488);
and U12800 (N_12800,N_12170,N_12079);
nor U12801 (N_12801,N_12016,N_12375);
xor U12802 (N_12802,N_12222,N_12299);
and U12803 (N_12803,N_12289,N_12330);
xnor U12804 (N_12804,N_12403,N_12052);
and U12805 (N_12805,N_12170,N_12357);
and U12806 (N_12806,N_12126,N_12157);
and U12807 (N_12807,N_12416,N_12081);
and U12808 (N_12808,N_12379,N_12218);
nand U12809 (N_12809,N_12044,N_12144);
and U12810 (N_12810,N_12029,N_12482);
and U12811 (N_12811,N_12108,N_12293);
and U12812 (N_12812,N_12331,N_12461);
or U12813 (N_12813,N_12307,N_12420);
nand U12814 (N_12814,N_12373,N_12073);
nand U12815 (N_12815,N_12456,N_12066);
nor U12816 (N_12816,N_12313,N_12026);
and U12817 (N_12817,N_12164,N_12031);
or U12818 (N_12818,N_12046,N_12109);
nor U12819 (N_12819,N_12008,N_12201);
and U12820 (N_12820,N_12057,N_12285);
nand U12821 (N_12821,N_12257,N_12171);
nand U12822 (N_12822,N_12007,N_12469);
nand U12823 (N_12823,N_12450,N_12148);
nor U12824 (N_12824,N_12231,N_12225);
nor U12825 (N_12825,N_12152,N_12318);
xor U12826 (N_12826,N_12465,N_12147);
xnor U12827 (N_12827,N_12181,N_12067);
xnor U12828 (N_12828,N_12223,N_12286);
nor U12829 (N_12829,N_12208,N_12377);
or U12830 (N_12830,N_12495,N_12329);
nor U12831 (N_12831,N_12295,N_12085);
or U12832 (N_12832,N_12142,N_12241);
nand U12833 (N_12833,N_12071,N_12465);
and U12834 (N_12834,N_12078,N_12271);
and U12835 (N_12835,N_12075,N_12447);
or U12836 (N_12836,N_12264,N_12199);
and U12837 (N_12837,N_12448,N_12125);
xnor U12838 (N_12838,N_12299,N_12471);
nor U12839 (N_12839,N_12366,N_12259);
nand U12840 (N_12840,N_12363,N_12109);
or U12841 (N_12841,N_12162,N_12237);
xor U12842 (N_12842,N_12239,N_12432);
xor U12843 (N_12843,N_12113,N_12174);
xnor U12844 (N_12844,N_12429,N_12313);
and U12845 (N_12845,N_12453,N_12268);
xnor U12846 (N_12846,N_12119,N_12301);
nand U12847 (N_12847,N_12239,N_12286);
nand U12848 (N_12848,N_12352,N_12318);
nor U12849 (N_12849,N_12363,N_12490);
xnor U12850 (N_12850,N_12034,N_12021);
nor U12851 (N_12851,N_12488,N_12288);
nor U12852 (N_12852,N_12344,N_12495);
nand U12853 (N_12853,N_12365,N_12107);
or U12854 (N_12854,N_12139,N_12377);
nor U12855 (N_12855,N_12490,N_12102);
nor U12856 (N_12856,N_12098,N_12451);
and U12857 (N_12857,N_12125,N_12202);
or U12858 (N_12858,N_12038,N_12470);
nor U12859 (N_12859,N_12031,N_12232);
nand U12860 (N_12860,N_12250,N_12017);
nor U12861 (N_12861,N_12164,N_12342);
and U12862 (N_12862,N_12144,N_12158);
or U12863 (N_12863,N_12259,N_12455);
nand U12864 (N_12864,N_12438,N_12161);
and U12865 (N_12865,N_12134,N_12173);
nand U12866 (N_12866,N_12264,N_12176);
or U12867 (N_12867,N_12028,N_12346);
or U12868 (N_12868,N_12274,N_12172);
and U12869 (N_12869,N_12414,N_12274);
or U12870 (N_12870,N_12005,N_12362);
xor U12871 (N_12871,N_12182,N_12044);
or U12872 (N_12872,N_12296,N_12067);
and U12873 (N_12873,N_12083,N_12393);
or U12874 (N_12874,N_12266,N_12130);
and U12875 (N_12875,N_12216,N_12351);
or U12876 (N_12876,N_12448,N_12122);
and U12877 (N_12877,N_12085,N_12156);
nor U12878 (N_12878,N_12493,N_12350);
and U12879 (N_12879,N_12375,N_12065);
and U12880 (N_12880,N_12358,N_12156);
xor U12881 (N_12881,N_12466,N_12002);
or U12882 (N_12882,N_12133,N_12143);
or U12883 (N_12883,N_12403,N_12332);
xor U12884 (N_12884,N_12036,N_12004);
nand U12885 (N_12885,N_12214,N_12406);
or U12886 (N_12886,N_12248,N_12394);
nand U12887 (N_12887,N_12087,N_12321);
nand U12888 (N_12888,N_12478,N_12496);
or U12889 (N_12889,N_12456,N_12395);
or U12890 (N_12890,N_12499,N_12116);
and U12891 (N_12891,N_12454,N_12243);
xor U12892 (N_12892,N_12445,N_12282);
nand U12893 (N_12893,N_12076,N_12398);
nand U12894 (N_12894,N_12042,N_12074);
nor U12895 (N_12895,N_12242,N_12118);
and U12896 (N_12896,N_12144,N_12244);
or U12897 (N_12897,N_12062,N_12243);
nand U12898 (N_12898,N_12141,N_12073);
and U12899 (N_12899,N_12369,N_12091);
xnor U12900 (N_12900,N_12326,N_12219);
or U12901 (N_12901,N_12285,N_12401);
nand U12902 (N_12902,N_12299,N_12013);
nand U12903 (N_12903,N_12274,N_12116);
nand U12904 (N_12904,N_12363,N_12390);
nor U12905 (N_12905,N_12461,N_12228);
xor U12906 (N_12906,N_12380,N_12095);
nand U12907 (N_12907,N_12161,N_12454);
or U12908 (N_12908,N_12091,N_12026);
and U12909 (N_12909,N_12163,N_12401);
xor U12910 (N_12910,N_12264,N_12146);
nor U12911 (N_12911,N_12026,N_12143);
and U12912 (N_12912,N_12035,N_12409);
nor U12913 (N_12913,N_12171,N_12152);
xor U12914 (N_12914,N_12200,N_12036);
or U12915 (N_12915,N_12005,N_12495);
and U12916 (N_12916,N_12111,N_12154);
or U12917 (N_12917,N_12230,N_12434);
xor U12918 (N_12918,N_12206,N_12195);
nand U12919 (N_12919,N_12325,N_12070);
and U12920 (N_12920,N_12290,N_12309);
and U12921 (N_12921,N_12314,N_12019);
xnor U12922 (N_12922,N_12109,N_12250);
and U12923 (N_12923,N_12436,N_12307);
xor U12924 (N_12924,N_12021,N_12110);
nand U12925 (N_12925,N_12213,N_12144);
nor U12926 (N_12926,N_12175,N_12210);
nor U12927 (N_12927,N_12220,N_12279);
xnor U12928 (N_12928,N_12175,N_12455);
nor U12929 (N_12929,N_12333,N_12070);
or U12930 (N_12930,N_12431,N_12120);
nand U12931 (N_12931,N_12391,N_12301);
or U12932 (N_12932,N_12297,N_12198);
nand U12933 (N_12933,N_12014,N_12069);
nor U12934 (N_12934,N_12203,N_12000);
or U12935 (N_12935,N_12101,N_12485);
or U12936 (N_12936,N_12239,N_12024);
or U12937 (N_12937,N_12181,N_12272);
nand U12938 (N_12938,N_12325,N_12132);
nand U12939 (N_12939,N_12348,N_12499);
or U12940 (N_12940,N_12006,N_12441);
xnor U12941 (N_12941,N_12163,N_12493);
and U12942 (N_12942,N_12370,N_12419);
xnor U12943 (N_12943,N_12072,N_12486);
nor U12944 (N_12944,N_12346,N_12029);
xnor U12945 (N_12945,N_12369,N_12334);
nor U12946 (N_12946,N_12463,N_12012);
nor U12947 (N_12947,N_12048,N_12401);
nor U12948 (N_12948,N_12235,N_12244);
and U12949 (N_12949,N_12387,N_12270);
nor U12950 (N_12950,N_12045,N_12016);
and U12951 (N_12951,N_12301,N_12319);
nand U12952 (N_12952,N_12102,N_12491);
nor U12953 (N_12953,N_12260,N_12317);
nand U12954 (N_12954,N_12050,N_12467);
nor U12955 (N_12955,N_12095,N_12174);
or U12956 (N_12956,N_12167,N_12408);
and U12957 (N_12957,N_12445,N_12328);
nand U12958 (N_12958,N_12284,N_12200);
nand U12959 (N_12959,N_12357,N_12456);
nor U12960 (N_12960,N_12026,N_12331);
or U12961 (N_12961,N_12230,N_12353);
and U12962 (N_12962,N_12018,N_12195);
nand U12963 (N_12963,N_12429,N_12222);
and U12964 (N_12964,N_12452,N_12458);
and U12965 (N_12965,N_12152,N_12468);
nor U12966 (N_12966,N_12478,N_12472);
nor U12967 (N_12967,N_12075,N_12066);
nor U12968 (N_12968,N_12373,N_12212);
xnor U12969 (N_12969,N_12187,N_12055);
and U12970 (N_12970,N_12124,N_12404);
xor U12971 (N_12971,N_12064,N_12151);
nand U12972 (N_12972,N_12493,N_12051);
xor U12973 (N_12973,N_12209,N_12389);
nand U12974 (N_12974,N_12167,N_12047);
and U12975 (N_12975,N_12140,N_12064);
and U12976 (N_12976,N_12134,N_12108);
and U12977 (N_12977,N_12038,N_12186);
nor U12978 (N_12978,N_12106,N_12361);
nand U12979 (N_12979,N_12149,N_12356);
nand U12980 (N_12980,N_12294,N_12082);
or U12981 (N_12981,N_12089,N_12208);
xnor U12982 (N_12982,N_12093,N_12374);
nor U12983 (N_12983,N_12313,N_12349);
nand U12984 (N_12984,N_12113,N_12156);
and U12985 (N_12985,N_12054,N_12260);
xnor U12986 (N_12986,N_12205,N_12350);
nor U12987 (N_12987,N_12201,N_12270);
nor U12988 (N_12988,N_12252,N_12402);
or U12989 (N_12989,N_12304,N_12475);
xor U12990 (N_12990,N_12225,N_12050);
xor U12991 (N_12991,N_12211,N_12271);
nand U12992 (N_12992,N_12466,N_12025);
and U12993 (N_12993,N_12083,N_12377);
or U12994 (N_12994,N_12075,N_12476);
nor U12995 (N_12995,N_12451,N_12304);
nor U12996 (N_12996,N_12287,N_12356);
nor U12997 (N_12997,N_12153,N_12115);
or U12998 (N_12998,N_12437,N_12026);
xor U12999 (N_12999,N_12030,N_12332);
and U13000 (N_13000,N_12811,N_12698);
xor U13001 (N_13001,N_12541,N_12790);
nor U13002 (N_13002,N_12722,N_12599);
nand U13003 (N_13003,N_12704,N_12894);
nor U13004 (N_13004,N_12775,N_12995);
or U13005 (N_13005,N_12523,N_12844);
xor U13006 (N_13006,N_12840,N_12761);
xor U13007 (N_13007,N_12782,N_12501);
or U13008 (N_13008,N_12584,N_12688);
and U13009 (N_13009,N_12615,N_12621);
or U13010 (N_13010,N_12574,N_12636);
nand U13011 (N_13011,N_12838,N_12510);
nor U13012 (N_13012,N_12757,N_12724);
xor U13013 (N_13013,N_12581,N_12971);
or U13014 (N_13014,N_12723,N_12793);
and U13015 (N_13015,N_12705,N_12877);
nor U13016 (N_13016,N_12856,N_12717);
xnor U13017 (N_13017,N_12559,N_12889);
nor U13018 (N_13018,N_12719,N_12817);
nand U13019 (N_13019,N_12921,N_12766);
and U13020 (N_13020,N_12853,N_12693);
xor U13021 (N_13021,N_12792,N_12617);
nand U13022 (N_13022,N_12742,N_12940);
and U13023 (N_13023,N_12732,N_12842);
nor U13024 (N_13024,N_12804,N_12537);
nand U13025 (N_13025,N_12843,N_12708);
nand U13026 (N_13026,N_12999,N_12568);
nor U13027 (N_13027,N_12866,N_12947);
or U13028 (N_13028,N_12819,N_12828);
xor U13029 (N_13029,N_12968,N_12992);
or U13030 (N_13030,N_12699,N_12593);
or U13031 (N_13031,N_12925,N_12653);
nand U13032 (N_13032,N_12884,N_12578);
xor U13033 (N_13033,N_12718,N_12952);
nor U13034 (N_13034,N_12878,N_12847);
or U13035 (N_13035,N_12656,N_12594);
xnor U13036 (N_13036,N_12809,N_12700);
nand U13037 (N_13037,N_12545,N_12676);
nor U13038 (N_13038,N_12648,N_12920);
and U13039 (N_13039,N_12778,N_12610);
xnor U13040 (N_13040,N_12726,N_12575);
or U13041 (N_13041,N_12706,N_12748);
nand U13042 (N_13042,N_12794,N_12964);
and U13043 (N_13043,N_12773,N_12528);
nor U13044 (N_13044,N_12978,N_12601);
nor U13045 (N_13045,N_12507,N_12784);
nor U13046 (N_13046,N_12588,N_12598);
nand U13047 (N_13047,N_12763,N_12808);
nand U13048 (N_13048,N_12609,N_12570);
and U13049 (N_13049,N_12977,N_12513);
nand U13050 (N_13050,N_12918,N_12987);
and U13051 (N_13051,N_12668,N_12572);
nor U13052 (N_13052,N_12777,N_12550);
or U13053 (N_13053,N_12924,N_12512);
and U13054 (N_13054,N_12919,N_12839);
nor U13055 (N_13055,N_12679,N_12872);
and U13056 (N_13056,N_12511,N_12701);
or U13057 (N_13057,N_12882,N_12988);
xnor U13058 (N_13058,N_12639,N_12611);
xnor U13059 (N_13059,N_12579,N_12576);
or U13060 (N_13060,N_12674,N_12739);
and U13061 (N_13061,N_12604,N_12551);
nor U13062 (N_13062,N_12681,N_12755);
and U13063 (N_13063,N_12595,N_12797);
or U13064 (N_13064,N_12682,N_12616);
xnor U13065 (N_13065,N_12963,N_12986);
xnor U13066 (N_13066,N_12506,N_12941);
xor U13067 (N_13067,N_12519,N_12862);
or U13068 (N_13068,N_12665,N_12531);
or U13069 (N_13069,N_12933,N_12630);
nand U13070 (N_13070,N_12509,N_12565);
nand U13071 (N_13071,N_12851,N_12927);
or U13072 (N_13072,N_12503,N_12926);
nand U13073 (N_13073,N_12996,N_12715);
nand U13074 (N_13074,N_12950,N_12951);
xnor U13075 (N_13075,N_12898,N_12622);
xor U13076 (N_13076,N_12547,N_12953);
and U13077 (N_13077,N_12721,N_12967);
xnor U13078 (N_13078,N_12984,N_12803);
nand U13079 (N_13079,N_12944,N_12955);
nand U13080 (N_13080,N_12922,N_12534);
xor U13081 (N_13081,N_12786,N_12983);
xnor U13082 (N_13082,N_12532,N_12695);
nand U13083 (N_13083,N_12857,N_12900);
xor U13084 (N_13084,N_12629,N_12657);
nand U13085 (N_13085,N_12798,N_12860);
xnor U13086 (N_13086,N_12897,N_12613);
or U13087 (N_13087,N_12634,N_12644);
and U13088 (N_13088,N_12652,N_12678);
nand U13089 (N_13089,N_12692,N_12991);
and U13090 (N_13090,N_12890,N_12834);
xnor U13091 (N_13091,N_12765,N_12555);
nor U13092 (N_13092,N_12727,N_12590);
xnor U13093 (N_13093,N_12910,N_12603);
nor U13094 (N_13094,N_12896,N_12875);
nor U13095 (N_13095,N_12549,N_12571);
or U13096 (N_13096,N_12768,N_12820);
and U13097 (N_13097,N_12743,N_12702);
or U13098 (N_13098,N_12923,N_12799);
or U13099 (N_13099,N_12666,N_12689);
nor U13100 (N_13100,N_12597,N_12907);
and U13101 (N_13101,N_12769,N_12660);
nor U13102 (N_13102,N_12902,N_12813);
nand U13103 (N_13103,N_12887,N_12841);
and U13104 (N_13104,N_12573,N_12558);
nand U13105 (N_13105,N_12873,N_12779);
and U13106 (N_13106,N_12974,N_12904);
nor U13107 (N_13107,N_12788,N_12626);
nand U13108 (N_13108,N_12680,N_12731);
nand U13109 (N_13109,N_12650,N_12942);
and U13110 (N_13110,N_12567,N_12937);
xnor U13111 (N_13111,N_12911,N_12795);
nand U13112 (N_13112,N_12754,N_12980);
nand U13113 (N_13113,N_12893,N_12961);
and U13114 (N_13114,N_12749,N_12837);
nand U13115 (N_13115,N_12871,N_12807);
xnor U13116 (N_13116,N_12711,N_12520);
nand U13117 (N_13117,N_12753,N_12526);
xor U13118 (N_13118,N_12989,N_12916);
nor U13119 (N_13119,N_12734,N_12865);
nand U13120 (N_13120,N_12957,N_12525);
nor U13121 (N_13121,N_12787,N_12728);
or U13122 (N_13122,N_12976,N_12858);
nor U13123 (N_13123,N_12552,N_12934);
nor U13124 (N_13124,N_12654,N_12970);
nor U13125 (N_13125,N_12959,N_12670);
nand U13126 (N_13126,N_12855,N_12880);
nor U13127 (N_13127,N_12850,N_12929);
xor U13128 (N_13128,N_12605,N_12876);
or U13129 (N_13129,N_12810,N_12677);
xnor U13130 (N_13130,N_12548,N_12789);
nor U13131 (N_13131,N_12835,N_12538);
xnor U13132 (N_13132,N_12883,N_12874);
or U13133 (N_13133,N_12939,N_12938);
nand U13134 (N_13134,N_12539,N_12891);
or U13135 (N_13135,N_12901,N_12580);
or U13136 (N_13136,N_12824,N_12675);
and U13137 (N_13137,N_12852,N_12535);
nor U13138 (N_13138,N_12710,N_12752);
nor U13139 (N_13139,N_12564,N_12741);
nor U13140 (N_13140,N_12931,N_12515);
nand U13141 (N_13141,N_12829,N_12909);
nand U13142 (N_13142,N_12914,N_12521);
or U13143 (N_13143,N_12767,N_12600);
xnor U13144 (N_13144,N_12928,N_12776);
xor U13145 (N_13145,N_12885,N_12899);
nor U13146 (N_13146,N_12703,N_12661);
nor U13147 (N_13147,N_12720,N_12879);
xor U13148 (N_13148,N_12832,N_12903);
and U13149 (N_13149,N_12659,N_12563);
nand U13150 (N_13150,N_12806,N_12972);
or U13151 (N_13151,N_12518,N_12713);
nor U13152 (N_13152,N_12994,N_12774);
or U13153 (N_13153,N_12958,N_12982);
nor U13154 (N_13154,N_12587,N_12729);
nor U13155 (N_13155,N_12631,N_12770);
and U13156 (N_13156,N_12536,N_12936);
nor U13157 (N_13157,N_12687,N_12672);
or U13158 (N_13158,N_12979,N_12759);
nand U13159 (N_13159,N_12906,N_12540);
xnor U13160 (N_13160,N_12791,N_12709);
nor U13161 (N_13161,N_12821,N_12527);
or U13162 (N_13162,N_12740,N_12869);
xnor U13163 (N_13163,N_12608,N_12888);
and U13164 (N_13164,N_12606,N_12602);
or U13165 (N_13165,N_12745,N_12805);
xnor U13166 (N_13166,N_12589,N_12764);
nand U13167 (N_13167,N_12750,N_12746);
nand U13168 (N_13168,N_12867,N_12658);
xnor U13169 (N_13169,N_12854,N_12756);
xor U13170 (N_13170,N_12935,N_12635);
nor U13171 (N_13171,N_12685,N_12990);
nor U13172 (N_13172,N_12975,N_12554);
or U13173 (N_13173,N_12530,N_12533);
nand U13174 (N_13174,N_12744,N_12823);
or U13175 (N_13175,N_12641,N_12667);
nand U13176 (N_13176,N_12502,N_12671);
xor U13177 (N_13177,N_12772,N_12825);
or U13178 (N_13178,N_12771,N_12544);
xor U13179 (N_13179,N_12915,N_12633);
and U13180 (N_13180,N_12997,N_12892);
nand U13181 (N_13181,N_12998,N_12973);
xnor U13182 (N_13182,N_12627,N_12624);
and U13183 (N_13183,N_12663,N_12673);
and U13184 (N_13184,N_12725,N_12881);
or U13185 (N_13185,N_12669,N_12816);
xnor U13186 (N_13186,N_12505,N_12945);
and U13187 (N_13187,N_12831,N_12524);
nand U13188 (N_13188,N_12625,N_12762);
nand U13189 (N_13189,N_12785,N_12886);
or U13190 (N_13190,N_12569,N_12684);
or U13191 (N_13191,N_12504,N_12690);
and U13192 (N_13192,N_12845,N_12949);
nand U13193 (N_13193,N_12751,N_12801);
nor U13194 (N_13194,N_12802,N_12815);
nor U13195 (N_13195,N_12560,N_12758);
or U13196 (N_13196,N_12960,N_12956);
nand U13197 (N_13197,N_12546,N_12591);
and U13198 (N_13198,N_12696,N_12566);
and U13199 (N_13199,N_12508,N_12848);
and U13200 (N_13200,N_12895,N_12814);
nand U13201 (N_13201,N_12716,N_12943);
nor U13202 (N_13202,N_12614,N_12868);
xor U13203 (N_13203,N_12542,N_12529);
xnor U13204 (N_13204,N_12637,N_12730);
and U13205 (N_13205,N_12628,N_12596);
nor U13206 (N_13206,N_12500,N_12683);
nor U13207 (N_13207,N_12664,N_12646);
xnor U13208 (N_13208,N_12686,N_12781);
and U13209 (N_13209,N_12905,N_12800);
nand U13210 (N_13210,N_12583,N_12736);
nand U13211 (N_13211,N_12582,N_12516);
xor U13212 (N_13212,N_12522,N_12612);
and U13213 (N_13213,N_12812,N_12735);
or U13214 (N_13214,N_12561,N_12623);
or U13215 (N_13215,N_12738,N_12863);
xnor U13216 (N_13216,N_12836,N_12864);
or U13217 (N_13217,N_12783,N_12946);
nand U13218 (N_13218,N_12649,N_12643);
and U13219 (N_13219,N_12556,N_12917);
and U13220 (N_13220,N_12859,N_12826);
nor U13221 (N_13221,N_12932,N_12849);
or U13222 (N_13222,N_12543,N_12655);
nand U13223 (N_13223,N_12993,N_12760);
nand U13224 (N_13224,N_12714,N_12619);
xnor U13225 (N_13225,N_12737,N_12981);
nor U13226 (N_13226,N_12733,N_12912);
xnor U13227 (N_13227,N_12620,N_12930);
xnor U13228 (N_13228,N_12638,N_12592);
nand U13229 (N_13229,N_12780,N_12577);
nand U13230 (N_13230,N_12707,N_12846);
and U13231 (N_13231,N_12965,N_12969);
or U13232 (N_13232,N_12647,N_12712);
or U13233 (N_13233,N_12645,N_12557);
or U13234 (N_13234,N_12697,N_12747);
or U13235 (N_13235,N_12818,N_12632);
xor U13236 (N_13236,N_12913,N_12517);
or U13237 (N_13237,N_12830,N_12585);
nand U13238 (N_13238,N_12861,N_12796);
nand U13239 (N_13239,N_12870,N_12985);
and U13240 (N_13240,N_12694,N_12948);
or U13241 (N_13241,N_12691,N_12827);
or U13242 (N_13242,N_12822,N_12966);
nand U13243 (N_13243,N_12640,N_12962);
xnor U13244 (N_13244,N_12833,N_12586);
or U13245 (N_13245,N_12562,N_12651);
or U13246 (N_13246,N_12642,N_12954);
nand U13247 (N_13247,N_12662,N_12607);
nor U13248 (N_13248,N_12514,N_12618);
nand U13249 (N_13249,N_12908,N_12553);
xnor U13250 (N_13250,N_12810,N_12506);
and U13251 (N_13251,N_12816,N_12599);
nor U13252 (N_13252,N_12505,N_12894);
or U13253 (N_13253,N_12641,N_12900);
or U13254 (N_13254,N_12606,N_12632);
xnor U13255 (N_13255,N_12948,N_12941);
nor U13256 (N_13256,N_12825,N_12826);
nand U13257 (N_13257,N_12950,N_12676);
xor U13258 (N_13258,N_12618,N_12538);
nand U13259 (N_13259,N_12904,N_12943);
or U13260 (N_13260,N_12647,N_12912);
nor U13261 (N_13261,N_12615,N_12859);
nor U13262 (N_13262,N_12518,N_12698);
or U13263 (N_13263,N_12595,N_12707);
and U13264 (N_13264,N_12780,N_12552);
nor U13265 (N_13265,N_12618,N_12908);
nor U13266 (N_13266,N_12683,N_12622);
or U13267 (N_13267,N_12722,N_12623);
nor U13268 (N_13268,N_12783,N_12916);
or U13269 (N_13269,N_12936,N_12775);
nor U13270 (N_13270,N_12804,N_12632);
xor U13271 (N_13271,N_12534,N_12686);
nor U13272 (N_13272,N_12663,N_12711);
xnor U13273 (N_13273,N_12992,N_12730);
nor U13274 (N_13274,N_12702,N_12720);
xor U13275 (N_13275,N_12906,N_12609);
or U13276 (N_13276,N_12642,N_12940);
xor U13277 (N_13277,N_12722,N_12636);
or U13278 (N_13278,N_12761,N_12990);
xor U13279 (N_13279,N_12863,N_12710);
nor U13280 (N_13280,N_12815,N_12925);
and U13281 (N_13281,N_12912,N_12899);
nor U13282 (N_13282,N_12690,N_12758);
and U13283 (N_13283,N_12562,N_12534);
nor U13284 (N_13284,N_12702,N_12690);
or U13285 (N_13285,N_12501,N_12592);
and U13286 (N_13286,N_12569,N_12688);
nand U13287 (N_13287,N_12854,N_12820);
nor U13288 (N_13288,N_12971,N_12770);
nor U13289 (N_13289,N_12563,N_12786);
and U13290 (N_13290,N_12995,N_12703);
nor U13291 (N_13291,N_12603,N_12832);
and U13292 (N_13292,N_12774,N_12735);
and U13293 (N_13293,N_12541,N_12889);
or U13294 (N_13294,N_12815,N_12949);
nor U13295 (N_13295,N_12814,N_12634);
or U13296 (N_13296,N_12784,N_12880);
nor U13297 (N_13297,N_12866,N_12889);
and U13298 (N_13298,N_12870,N_12820);
and U13299 (N_13299,N_12694,N_12700);
nand U13300 (N_13300,N_12843,N_12886);
nand U13301 (N_13301,N_12821,N_12573);
and U13302 (N_13302,N_12594,N_12603);
xnor U13303 (N_13303,N_12827,N_12531);
and U13304 (N_13304,N_12909,N_12643);
or U13305 (N_13305,N_12819,N_12974);
nor U13306 (N_13306,N_12752,N_12804);
or U13307 (N_13307,N_12532,N_12964);
nand U13308 (N_13308,N_12877,N_12737);
nand U13309 (N_13309,N_12827,N_12977);
or U13310 (N_13310,N_12722,N_12961);
and U13311 (N_13311,N_12832,N_12934);
xnor U13312 (N_13312,N_12994,N_12602);
and U13313 (N_13313,N_12759,N_12599);
or U13314 (N_13314,N_12857,N_12856);
xor U13315 (N_13315,N_12768,N_12574);
xor U13316 (N_13316,N_12799,N_12520);
nor U13317 (N_13317,N_12842,N_12558);
and U13318 (N_13318,N_12503,N_12922);
and U13319 (N_13319,N_12981,N_12670);
and U13320 (N_13320,N_12693,N_12690);
nor U13321 (N_13321,N_12627,N_12522);
xor U13322 (N_13322,N_12977,N_12735);
and U13323 (N_13323,N_12654,N_12765);
xor U13324 (N_13324,N_12939,N_12583);
xnor U13325 (N_13325,N_12925,N_12761);
xor U13326 (N_13326,N_12681,N_12673);
nor U13327 (N_13327,N_12626,N_12650);
xnor U13328 (N_13328,N_12819,N_12853);
or U13329 (N_13329,N_12605,N_12805);
or U13330 (N_13330,N_12537,N_12933);
nand U13331 (N_13331,N_12944,N_12842);
and U13332 (N_13332,N_12897,N_12909);
xor U13333 (N_13333,N_12545,N_12641);
nor U13334 (N_13334,N_12842,N_12542);
nand U13335 (N_13335,N_12990,N_12806);
nand U13336 (N_13336,N_12734,N_12949);
xor U13337 (N_13337,N_12961,N_12864);
or U13338 (N_13338,N_12808,N_12606);
nand U13339 (N_13339,N_12870,N_12553);
or U13340 (N_13340,N_12939,N_12800);
nor U13341 (N_13341,N_12671,N_12959);
nor U13342 (N_13342,N_12889,N_12844);
xnor U13343 (N_13343,N_12843,N_12616);
or U13344 (N_13344,N_12618,N_12836);
xor U13345 (N_13345,N_12878,N_12771);
xor U13346 (N_13346,N_12574,N_12709);
xor U13347 (N_13347,N_12598,N_12850);
nor U13348 (N_13348,N_12787,N_12581);
nor U13349 (N_13349,N_12740,N_12734);
nor U13350 (N_13350,N_12744,N_12850);
and U13351 (N_13351,N_12591,N_12504);
and U13352 (N_13352,N_12646,N_12922);
xnor U13353 (N_13353,N_12884,N_12583);
or U13354 (N_13354,N_12655,N_12860);
nor U13355 (N_13355,N_12732,N_12753);
nand U13356 (N_13356,N_12918,N_12593);
and U13357 (N_13357,N_12667,N_12871);
xor U13358 (N_13358,N_12928,N_12565);
and U13359 (N_13359,N_12798,N_12777);
xnor U13360 (N_13360,N_12835,N_12511);
and U13361 (N_13361,N_12850,N_12944);
nand U13362 (N_13362,N_12939,N_12788);
nor U13363 (N_13363,N_12855,N_12805);
and U13364 (N_13364,N_12936,N_12571);
or U13365 (N_13365,N_12510,N_12994);
nor U13366 (N_13366,N_12561,N_12586);
nand U13367 (N_13367,N_12546,N_12868);
nand U13368 (N_13368,N_12528,N_12913);
nand U13369 (N_13369,N_12818,N_12777);
nor U13370 (N_13370,N_12660,N_12882);
nor U13371 (N_13371,N_12601,N_12754);
nand U13372 (N_13372,N_12989,N_12883);
and U13373 (N_13373,N_12779,N_12858);
and U13374 (N_13374,N_12937,N_12833);
nor U13375 (N_13375,N_12772,N_12980);
nor U13376 (N_13376,N_12566,N_12791);
nor U13377 (N_13377,N_12524,N_12691);
and U13378 (N_13378,N_12779,N_12764);
xnor U13379 (N_13379,N_12625,N_12600);
and U13380 (N_13380,N_12746,N_12567);
nand U13381 (N_13381,N_12819,N_12947);
and U13382 (N_13382,N_12871,N_12705);
xnor U13383 (N_13383,N_12867,N_12576);
nor U13384 (N_13384,N_12853,N_12991);
and U13385 (N_13385,N_12880,N_12762);
nand U13386 (N_13386,N_12949,N_12990);
or U13387 (N_13387,N_12576,N_12833);
xor U13388 (N_13388,N_12617,N_12599);
or U13389 (N_13389,N_12863,N_12764);
nand U13390 (N_13390,N_12722,N_12957);
and U13391 (N_13391,N_12546,N_12840);
nand U13392 (N_13392,N_12814,N_12581);
xor U13393 (N_13393,N_12526,N_12632);
and U13394 (N_13394,N_12789,N_12654);
or U13395 (N_13395,N_12811,N_12824);
and U13396 (N_13396,N_12712,N_12813);
and U13397 (N_13397,N_12905,N_12505);
nor U13398 (N_13398,N_12939,N_12985);
or U13399 (N_13399,N_12851,N_12594);
and U13400 (N_13400,N_12950,N_12766);
xnor U13401 (N_13401,N_12500,N_12966);
xor U13402 (N_13402,N_12769,N_12636);
and U13403 (N_13403,N_12709,N_12666);
and U13404 (N_13404,N_12706,N_12761);
nand U13405 (N_13405,N_12590,N_12670);
xor U13406 (N_13406,N_12876,N_12927);
xor U13407 (N_13407,N_12817,N_12740);
or U13408 (N_13408,N_12624,N_12987);
nand U13409 (N_13409,N_12862,N_12834);
nor U13410 (N_13410,N_12531,N_12880);
nor U13411 (N_13411,N_12747,N_12549);
nor U13412 (N_13412,N_12943,N_12987);
xnor U13413 (N_13413,N_12573,N_12517);
and U13414 (N_13414,N_12836,N_12631);
nand U13415 (N_13415,N_12832,N_12987);
and U13416 (N_13416,N_12766,N_12991);
and U13417 (N_13417,N_12690,N_12622);
and U13418 (N_13418,N_12587,N_12994);
nor U13419 (N_13419,N_12954,N_12786);
nand U13420 (N_13420,N_12844,N_12587);
nand U13421 (N_13421,N_12996,N_12683);
nor U13422 (N_13422,N_12896,N_12644);
and U13423 (N_13423,N_12671,N_12966);
or U13424 (N_13424,N_12703,N_12563);
nand U13425 (N_13425,N_12632,N_12679);
or U13426 (N_13426,N_12866,N_12978);
or U13427 (N_13427,N_12689,N_12729);
and U13428 (N_13428,N_12728,N_12774);
nor U13429 (N_13429,N_12752,N_12501);
nand U13430 (N_13430,N_12554,N_12854);
nand U13431 (N_13431,N_12635,N_12934);
and U13432 (N_13432,N_12812,N_12730);
nand U13433 (N_13433,N_12815,N_12957);
or U13434 (N_13434,N_12627,N_12745);
and U13435 (N_13435,N_12566,N_12663);
xor U13436 (N_13436,N_12815,N_12845);
and U13437 (N_13437,N_12911,N_12893);
nand U13438 (N_13438,N_12958,N_12567);
nand U13439 (N_13439,N_12526,N_12767);
nor U13440 (N_13440,N_12923,N_12621);
nand U13441 (N_13441,N_12918,N_12522);
nor U13442 (N_13442,N_12817,N_12819);
nand U13443 (N_13443,N_12857,N_12573);
nor U13444 (N_13444,N_12826,N_12762);
nand U13445 (N_13445,N_12736,N_12861);
or U13446 (N_13446,N_12674,N_12638);
or U13447 (N_13447,N_12632,N_12901);
nand U13448 (N_13448,N_12645,N_12550);
and U13449 (N_13449,N_12931,N_12563);
or U13450 (N_13450,N_12711,N_12995);
nor U13451 (N_13451,N_12752,N_12868);
nor U13452 (N_13452,N_12616,N_12838);
nor U13453 (N_13453,N_12970,N_12724);
nor U13454 (N_13454,N_12876,N_12926);
nand U13455 (N_13455,N_12581,N_12954);
nor U13456 (N_13456,N_12602,N_12935);
xor U13457 (N_13457,N_12883,N_12721);
nor U13458 (N_13458,N_12882,N_12518);
or U13459 (N_13459,N_12840,N_12564);
nor U13460 (N_13460,N_12644,N_12633);
or U13461 (N_13461,N_12997,N_12907);
nor U13462 (N_13462,N_12758,N_12660);
and U13463 (N_13463,N_12783,N_12922);
nor U13464 (N_13464,N_12508,N_12675);
and U13465 (N_13465,N_12531,N_12762);
nor U13466 (N_13466,N_12853,N_12870);
or U13467 (N_13467,N_12820,N_12801);
nand U13468 (N_13468,N_12884,N_12518);
and U13469 (N_13469,N_12830,N_12846);
nand U13470 (N_13470,N_12583,N_12650);
and U13471 (N_13471,N_12649,N_12535);
nor U13472 (N_13472,N_12635,N_12741);
xor U13473 (N_13473,N_12792,N_12763);
nand U13474 (N_13474,N_12655,N_12994);
xor U13475 (N_13475,N_12891,N_12708);
xor U13476 (N_13476,N_12675,N_12933);
nor U13477 (N_13477,N_12757,N_12704);
nor U13478 (N_13478,N_12724,N_12904);
xor U13479 (N_13479,N_12946,N_12731);
nand U13480 (N_13480,N_12651,N_12631);
nor U13481 (N_13481,N_12554,N_12871);
xnor U13482 (N_13482,N_12988,N_12937);
or U13483 (N_13483,N_12814,N_12929);
or U13484 (N_13484,N_12573,N_12562);
xor U13485 (N_13485,N_12899,N_12735);
nor U13486 (N_13486,N_12820,N_12552);
and U13487 (N_13487,N_12697,N_12788);
nor U13488 (N_13488,N_12774,N_12755);
xor U13489 (N_13489,N_12564,N_12552);
or U13490 (N_13490,N_12719,N_12858);
xnor U13491 (N_13491,N_12546,N_12612);
or U13492 (N_13492,N_12716,N_12961);
xor U13493 (N_13493,N_12540,N_12691);
nor U13494 (N_13494,N_12587,N_12596);
nand U13495 (N_13495,N_12956,N_12764);
or U13496 (N_13496,N_12928,N_12719);
and U13497 (N_13497,N_12679,N_12576);
or U13498 (N_13498,N_12557,N_12709);
nor U13499 (N_13499,N_12645,N_12587);
nand U13500 (N_13500,N_13013,N_13067);
nor U13501 (N_13501,N_13053,N_13133);
nor U13502 (N_13502,N_13342,N_13038);
or U13503 (N_13503,N_13220,N_13070);
and U13504 (N_13504,N_13226,N_13290);
nor U13505 (N_13505,N_13228,N_13493);
nor U13506 (N_13506,N_13004,N_13196);
and U13507 (N_13507,N_13237,N_13003);
xnor U13508 (N_13508,N_13163,N_13080);
nand U13509 (N_13509,N_13169,N_13295);
or U13510 (N_13510,N_13094,N_13093);
xnor U13511 (N_13511,N_13275,N_13023);
and U13512 (N_13512,N_13106,N_13077);
nand U13513 (N_13513,N_13308,N_13151);
or U13514 (N_13514,N_13118,N_13112);
nor U13515 (N_13515,N_13294,N_13395);
xnor U13516 (N_13516,N_13417,N_13071);
and U13517 (N_13517,N_13389,N_13204);
nor U13518 (N_13518,N_13249,N_13393);
or U13519 (N_13519,N_13218,N_13364);
and U13520 (N_13520,N_13154,N_13422);
and U13521 (N_13521,N_13471,N_13054);
and U13522 (N_13522,N_13260,N_13254);
and U13523 (N_13523,N_13059,N_13410);
or U13524 (N_13524,N_13245,N_13207);
and U13525 (N_13525,N_13480,N_13376);
nor U13526 (N_13526,N_13205,N_13247);
xor U13527 (N_13527,N_13402,N_13005);
and U13528 (N_13528,N_13333,N_13000);
nor U13529 (N_13529,N_13336,N_13128);
nand U13530 (N_13530,N_13432,N_13406);
nor U13531 (N_13531,N_13208,N_13174);
xnor U13532 (N_13532,N_13160,N_13031);
and U13533 (N_13533,N_13474,N_13442);
xor U13534 (N_13534,N_13449,N_13124);
nand U13535 (N_13535,N_13391,N_13462);
and U13536 (N_13536,N_13338,N_13274);
nand U13537 (N_13537,N_13001,N_13048);
nor U13538 (N_13538,N_13026,N_13036);
and U13539 (N_13539,N_13147,N_13414);
nor U13540 (N_13540,N_13490,N_13426);
nand U13541 (N_13541,N_13136,N_13496);
or U13542 (N_13542,N_13195,N_13337);
or U13543 (N_13543,N_13375,N_13020);
nand U13544 (N_13544,N_13351,N_13134);
nand U13545 (N_13545,N_13327,N_13286);
or U13546 (N_13546,N_13314,N_13132);
nor U13547 (N_13547,N_13448,N_13084);
or U13548 (N_13548,N_13390,N_13252);
nand U13549 (N_13549,N_13244,N_13498);
and U13550 (N_13550,N_13323,N_13350);
nand U13551 (N_13551,N_13344,N_13266);
and U13552 (N_13552,N_13325,N_13100);
or U13553 (N_13553,N_13170,N_13074);
nor U13554 (N_13554,N_13461,N_13387);
and U13555 (N_13555,N_13045,N_13483);
or U13556 (N_13556,N_13158,N_13135);
nand U13557 (N_13557,N_13475,N_13201);
xor U13558 (N_13558,N_13453,N_13185);
or U13559 (N_13559,N_13159,N_13024);
and U13560 (N_13560,N_13485,N_13078);
or U13561 (N_13561,N_13428,N_13111);
nor U13562 (N_13562,N_13289,N_13386);
and U13563 (N_13563,N_13371,N_13146);
and U13564 (N_13564,N_13262,N_13246);
and U13565 (N_13565,N_13097,N_13303);
nor U13566 (N_13566,N_13029,N_13380);
nor U13567 (N_13567,N_13401,N_13231);
or U13568 (N_13568,N_13049,N_13122);
nand U13569 (N_13569,N_13041,N_13460);
xnor U13570 (N_13570,N_13438,N_13319);
nand U13571 (N_13571,N_13152,N_13330);
nand U13572 (N_13572,N_13110,N_13119);
and U13573 (N_13573,N_13037,N_13372);
nand U13574 (N_13574,N_13370,N_13312);
nor U13575 (N_13575,N_13358,N_13014);
nor U13576 (N_13576,N_13162,N_13463);
or U13577 (N_13577,N_13413,N_13412);
and U13578 (N_13578,N_13011,N_13306);
nor U13579 (N_13579,N_13469,N_13473);
or U13580 (N_13580,N_13348,N_13369);
xor U13581 (N_13581,N_13360,N_13114);
nand U13582 (N_13582,N_13176,N_13304);
or U13583 (N_13583,N_13141,N_13271);
nand U13584 (N_13584,N_13148,N_13221);
and U13585 (N_13585,N_13316,N_13399);
and U13586 (N_13586,N_13057,N_13092);
or U13587 (N_13587,N_13302,N_13009);
and U13588 (N_13588,N_13063,N_13108);
nand U13589 (N_13589,N_13157,N_13285);
xor U13590 (N_13590,N_13378,N_13145);
and U13591 (N_13591,N_13040,N_13030);
nand U13592 (N_13592,N_13035,N_13476);
or U13593 (N_13593,N_13181,N_13310);
nor U13594 (N_13594,N_13039,N_13165);
nor U13595 (N_13595,N_13392,N_13318);
or U13596 (N_13596,N_13086,N_13434);
or U13597 (N_13597,N_13255,N_13409);
nand U13598 (N_13598,N_13486,N_13206);
or U13599 (N_13599,N_13243,N_13065);
nor U13600 (N_13600,N_13349,N_13222);
and U13601 (N_13601,N_13352,N_13288);
nand U13602 (N_13602,N_13489,N_13497);
and U13603 (N_13603,N_13293,N_13335);
or U13604 (N_13604,N_13028,N_13427);
or U13605 (N_13605,N_13436,N_13332);
nand U13606 (N_13606,N_13385,N_13216);
or U13607 (N_13607,N_13361,N_13305);
or U13608 (N_13608,N_13367,N_13235);
and U13609 (N_13609,N_13217,N_13354);
nand U13610 (N_13610,N_13472,N_13033);
and U13611 (N_13611,N_13464,N_13055);
and U13612 (N_13612,N_13066,N_13006);
or U13613 (N_13613,N_13405,N_13015);
or U13614 (N_13614,N_13443,N_13214);
and U13615 (N_13615,N_13396,N_13281);
nor U13616 (N_13616,N_13018,N_13400);
nor U13617 (N_13617,N_13149,N_13355);
or U13618 (N_13618,N_13088,N_13334);
nand U13619 (N_13619,N_13492,N_13189);
or U13620 (N_13620,N_13034,N_13224);
nor U13621 (N_13621,N_13435,N_13459);
or U13622 (N_13622,N_13073,N_13347);
xnor U13623 (N_13623,N_13016,N_13309);
and U13624 (N_13624,N_13050,N_13415);
or U13625 (N_13625,N_13099,N_13025);
nor U13626 (N_13626,N_13282,N_13076);
nand U13627 (N_13627,N_13043,N_13383);
or U13628 (N_13628,N_13107,N_13424);
nor U13629 (N_13629,N_13127,N_13215);
nand U13630 (N_13630,N_13184,N_13081);
and U13631 (N_13631,N_13256,N_13212);
and U13632 (N_13632,N_13441,N_13002);
and U13633 (N_13633,N_13156,N_13253);
xor U13634 (N_13634,N_13328,N_13115);
or U13635 (N_13635,N_13175,N_13276);
and U13636 (N_13636,N_13230,N_13191);
xor U13637 (N_13637,N_13467,N_13056);
nand U13638 (N_13638,N_13340,N_13433);
xor U13639 (N_13639,N_13403,N_13283);
nand U13640 (N_13640,N_13368,N_13484);
xnor U13641 (N_13641,N_13447,N_13192);
xnor U13642 (N_13642,N_13418,N_13116);
nand U13643 (N_13643,N_13095,N_13455);
nor U13644 (N_13644,N_13047,N_13173);
nand U13645 (N_13645,N_13103,N_13085);
nor U13646 (N_13646,N_13126,N_13227);
or U13647 (N_13647,N_13280,N_13121);
nor U13648 (N_13648,N_13143,N_13346);
nor U13649 (N_13649,N_13250,N_13384);
nand U13650 (N_13650,N_13365,N_13104);
nand U13651 (N_13651,N_13322,N_13313);
xor U13652 (N_13652,N_13123,N_13278);
or U13653 (N_13653,N_13270,N_13379);
or U13654 (N_13654,N_13420,N_13202);
and U13655 (N_13655,N_13416,N_13439);
nand U13656 (N_13656,N_13017,N_13144);
nand U13657 (N_13657,N_13190,N_13263);
and U13658 (N_13658,N_13488,N_13357);
nand U13659 (N_13659,N_13272,N_13423);
nand U13660 (N_13660,N_13284,N_13219);
nand U13661 (N_13661,N_13445,N_13478);
xnor U13662 (N_13662,N_13153,N_13321);
nor U13663 (N_13663,N_13150,N_13339);
and U13664 (N_13664,N_13075,N_13200);
and U13665 (N_13665,N_13072,N_13491);
xnor U13666 (N_13666,N_13166,N_13362);
nand U13667 (N_13667,N_13331,N_13404);
and U13668 (N_13668,N_13203,N_13248);
and U13669 (N_13669,N_13481,N_13373);
nand U13670 (N_13670,N_13456,N_13477);
nand U13671 (N_13671,N_13240,N_13320);
nand U13672 (N_13672,N_13421,N_13277);
nand U13673 (N_13673,N_13010,N_13171);
nand U13674 (N_13674,N_13105,N_13466);
xor U13675 (N_13675,N_13164,N_13209);
nand U13676 (N_13676,N_13044,N_13259);
xnor U13677 (N_13677,N_13382,N_13140);
nand U13678 (N_13678,N_13225,N_13082);
nand U13679 (N_13679,N_13251,N_13155);
nor U13680 (N_13680,N_13142,N_13326);
nand U13681 (N_13681,N_13180,N_13457);
nor U13682 (N_13682,N_13012,N_13161);
xnor U13683 (N_13683,N_13234,N_13408);
xnor U13684 (N_13684,N_13213,N_13300);
nand U13685 (N_13685,N_13064,N_13374);
xnor U13686 (N_13686,N_13411,N_13345);
or U13687 (N_13687,N_13487,N_13307);
xor U13688 (N_13688,N_13046,N_13032);
and U13689 (N_13689,N_13087,N_13098);
nor U13690 (N_13690,N_13458,N_13397);
and U13691 (N_13691,N_13052,N_13019);
and U13692 (N_13692,N_13186,N_13102);
nor U13693 (N_13693,N_13091,N_13356);
xnor U13694 (N_13694,N_13168,N_13198);
or U13695 (N_13695,N_13109,N_13363);
and U13696 (N_13696,N_13296,N_13257);
nor U13697 (N_13697,N_13398,N_13437);
xnor U13698 (N_13698,N_13187,N_13177);
nor U13699 (N_13699,N_13299,N_13193);
xnor U13700 (N_13700,N_13482,N_13499);
nand U13701 (N_13701,N_13468,N_13341);
nand U13702 (N_13702,N_13494,N_13236);
nor U13703 (N_13703,N_13229,N_13291);
nand U13704 (N_13704,N_13470,N_13172);
or U13705 (N_13705,N_13096,N_13021);
nor U13706 (N_13706,N_13261,N_13465);
and U13707 (N_13707,N_13139,N_13241);
nand U13708 (N_13708,N_13265,N_13239);
and U13709 (N_13709,N_13419,N_13431);
nand U13710 (N_13710,N_13407,N_13027);
nor U13711 (N_13711,N_13324,N_13125);
xnor U13712 (N_13712,N_13317,N_13232);
nand U13713 (N_13713,N_13450,N_13131);
nand U13714 (N_13714,N_13130,N_13233);
nor U13715 (N_13715,N_13329,N_13129);
nor U13716 (N_13716,N_13183,N_13287);
and U13717 (N_13717,N_13366,N_13451);
xor U13718 (N_13718,N_13138,N_13258);
or U13719 (N_13719,N_13452,N_13429);
xnor U13720 (N_13720,N_13051,N_13188);
nand U13721 (N_13721,N_13042,N_13068);
xnor U13722 (N_13722,N_13079,N_13060);
or U13723 (N_13723,N_13430,N_13425);
nor U13724 (N_13724,N_13101,N_13061);
and U13725 (N_13725,N_13394,N_13223);
nand U13726 (N_13726,N_13022,N_13120);
nor U13727 (N_13727,N_13359,N_13279);
nand U13728 (N_13728,N_13264,N_13495);
nand U13729 (N_13729,N_13090,N_13007);
xor U13730 (N_13730,N_13454,N_13211);
xnor U13731 (N_13731,N_13311,N_13167);
nor U13732 (N_13732,N_13377,N_13089);
and U13733 (N_13733,N_13298,N_13199);
nand U13734 (N_13734,N_13210,N_13446);
and U13735 (N_13735,N_13297,N_13479);
nand U13736 (N_13736,N_13242,N_13269);
nor U13737 (N_13737,N_13117,N_13137);
nand U13738 (N_13738,N_13062,N_13058);
nor U13739 (N_13739,N_13273,N_13083);
nor U13740 (N_13740,N_13381,N_13179);
xnor U13741 (N_13741,N_13353,N_13292);
nand U13742 (N_13742,N_13069,N_13178);
nor U13743 (N_13743,N_13008,N_13315);
or U13744 (N_13744,N_13197,N_13440);
or U13745 (N_13745,N_13194,N_13268);
and U13746 (N_13746,N_13267,N_13301);
or U13747 (N_13747,N_13182,N_13343);
nor U13748 (N_13748,N_13238,N_13388);
and U13749 (N_13749,N_13444,N_13113);
or U13750 (N_13750,N_13029,N_13165);
xor U13751 (N_13751,N_13433,N_13187);
and U13752 (N_13752,N_13109,N_13071);
nor U13753 (N_13753,N_13454,N_13193);
nand U13754 (N_13754,N_13363,N_13210);
nor U13755 (N_13755,N_13075,N_13179);
xor U13756 (N_13756,N_13027,N_13389);
and U13757 (N_13757,N_13119,N_13194);
and U13758 (N_13758,N_13479,N_13219);
nand U13759 (N_13759,N_13150,N_13022);
and U13760 (N_13760,N_13473,N_13351);
nor U13761 (N_13761,N_13473,N_13025);
or U13762 (N_13762,N_13339,N_13343);
and U13763 (N_13763,N_13135,N_13366);
and U13764 (N_13764,N_13136,N_13273);
xnor U13765 (N_13765,N_13434,N_13046);
nor U13766 (N_13766,N_13417,N_13047);
nand U13767 (N_13767,N_13381,N_13076);
nand U13768 (N_13768,N_13310,N_13464);
or U13769 (N_13769,N_13440,N_13005);
and U13770 (N_13770,N_13164,N_13034);
xnor U13771 (N_13771,N_13123,N_13370);
nor U13772 (N_13772,N_13167,N_13381);
and U13773 (N_13773,N_13498,N_13424);
or U13774 (N_13774,N_13077,N_13075);
and U13775 (N_13775,N_13044,N_13194);
xor U13776 (N_13776,N_13204,N_13297);
nand U13777 (N_13777,N_13270,N_13431);
and U13778 (N_13778,N_13045,N_13332);
nor U13779 (N_13779,N_13361,N_13172);
xor U13780 (N_13780,N_13130,N_13204);
nor U13781 (N_13781,N_13185,N_13419);
nor U13782 (N_13782,N_13380,N_13247);
or U13783 (N_13783,N_13054,N_13134);
nand U13784 (N_13784,N_13003,N_13078);
nand U13785 (N_13785,N_13403,N_13358);
nand U13786 (N_13786,N_13065,N_13318);
nor U13787 (N_13787,N_13408,N_13089);
or U13788 (N_13788,N_13497,N_13164);
xnor U13789 (N_13789,N_13469,N_13234);
nand U13790 (N_13790,N_13133,N_13153);
xor U13791 (N_13791,N_13228,N_13029);
nor U13792 (N_13792,N_13464,N_13057);
nor U13793 (N_13793,N_13490,N_13196);
and U13794 (N_13794,N_13229,N_13037);
xor U13795 (N_13795,N_13426,N_13085);
nor U13796 (N_13796,N_13422,N_13104);
and U13797 (N_13797,N_13053,N_13143);
or U13798 (N_13798,N_13027,N_13141);
nand U13799 (N_13799,N_13460,N_13458);
or U13800 (N_13800,N_13348,N_13010);
nand U13801 (N_13801,N_13011,N_13125);
and U13802 (N_13802,N_13259,N_13466);
nand U13803 (N_13803,N_13026,N_13322);
and U13804 (N_13804,N_13430,N_13142);
and U13805 (N_13805,N_13177,N_13259);
or U13806 (N_13806,N_13129,N_13205);
or U13807 (N_13807,N_13119,N_13379);
nand U13808 (N_13808,N_13081,N_13430);
and U13809 (N_13809,N_13210,N_13250);
nor U13810 (N_13810,N_13005,N_13241);
nor U13811 (N_13811,N_13065,N_13499);
or U13812 (N_13812,N_13123,N_13075);
xnor U13813 (N_13813,N_13374,N_13204);
nor U13814 (N_13814,N_13497,N_13333);
nor U13815 (N_13815,N_13139,N_13426);
xor U13816 (N_13816,N_13138,N_13487);
nand U13817 (N_13817,N_13341,N_13457);
and U13818 (N_13818,N_13003,N_13471);
and U13819 (N_13819,N_13002,N_13293);
nand U13820 (N_13820,N_13498,N_13469);
nor U13821 (N_13821,N_13455,N_13461);
nor U13822 (N_13822,N_13244,N_13050);
or U13823 (N_13823,N_13472,N_13156);
nand U13824 (N_13824,N_13015,N_13032);
xor U13825 (N_13825,N_13234,N_13410);
xnor U13826 (N_13826,N_13127,N_13279);
or U13827 (N_13827,N_13415,N_13087);
nor U13828 (N_13828,N_13053,N_13445);
nor U13829 (N_13829,N_13478,N_13118);
nand U13830 (N_13830,N_13447,N_13152);
or U13831 (N_13831,N_13336,N_13151);
and U13832 (N_13832,N_13341,N_13494);
xor U13833 (N_13833,N_13110,N_13351);
xor U13834 (N_13834,N_13132,N_13177);
or U13835 (N_13835,N_13438,N_13360);
xor U13836 (N_13836,N_13487,N_13474);
or U13837 (N_13837,N_13042,N_13065);
nand U13838 (N_13838,N_13184,N_13452);
and U13839 (N_13839,N_13053,N_13061);
nand U13840 (N_13840,N_13214,N_13172);
nor U13841 (N_13841,N_13449,N_13275);
nand U13842 (N_13842,N_13328,N_13161);
nor U13843 (N_13843,N_13140,N_13308);
nand U13844 (N_13844,N_13138,N_13060);
xor U13845 (N_13845,N_13137,N_13403);
or U13846 (N_13846,N_13430,N_13015);
nor U13847 (N_13847,N_13251,N_13372);
nand U13848 (N_13848,N_13113,N_13244);
and U13849 (N_13849,N_13140,N_13236);
nand U13850 (N_13850,N_13271,N_13047);
xnor U13851 (N_13851,N_13059,N_13075);
and U13852 (N_13852,N_13499,N_13204);
nor U13853 (N_13853,N_13339,N_13022);
and U13854 (N_13854,N_13309,N_13494);
or U13855 (N_13855,N_13064,N_13469);
nand U13856 (N_13856,N_13201,N_13283);
xor U13857 (N_13857,N_13496,N_13085);
and U13858 (N_13858,N_13468,N_13060);
or U13859 (N_13859,N_13002,N_13469);
nand U13860 (N_13860,N_13284,N_13326);
or U13861 (N_13861,N_13351,N_13101);
nor U13862 (N_13862,N_13192,N_13346);
xnor U13863 (N_13863,N_13396,N_13158);
nand U13864 (N_13864,N_13241,N_13118);
nor U13865 (N_13865,N_13028,N_13254);
nand U13866 (N_13866,N_13401,N_13140);
and U13867 (N_13867,N_13048,N_13011);
and U13868 (N_13868,N_13189,N_13105);
xnor U13869 (N_13869,N_13184,N_13219);
or U13870 (N_13870,N_13408,N_13196);
and U13871 (N_13871,N_13262,N_13112);
xnor U13872 (N_13872,N_13288,N_13472);
xnor U13873 (N_13873,N_13126,N_13499);
or U13874 (N_13874,N_13103,N_13215);
or U13875 (N_13875,N_13042,N_13418);
or U13876 (N_13876,N_13273,N_13044);
xnor U13877 (N_13877,N_13131,N_13262);
nor U13878 (N_13878,N_13444,N_13336);
and U13879 (N_13879,N_13455,N_13010);
xor U13880 (N_13880,N_13333,N_13308);
or U13881 (N_13881,N_13261,N_13122);
or U13882 (N_13882,N_13072,N_13283);
and U13883 (N_13883,N_13115,N_13437);
nor U13884 (N_13884,N_13114,N_13299);
and U13885 (N_13885,N_13480,N_13342);
or U13886 (N_13886,N_13234,N_13039);
nand U13887 (N_13887,N_13399,N_13493);
nand U13888 (N_13888,N_13286,N_13228);
nand U13889 (N_13889,N_13043,N_13165);
xor U13890 (N_13890,N_13198,N_13033);
xor U13891 (N_13891,N_13342,N_13456);
nor U13892 (N_13892,N_13432,N_13255);
nand U13893 (N_13893,N_13343,N_13374);
and U13894 (N_13894,N_13430,N_13180);
or U13895 (N_13895,N_13467,N_13431);
xor U13896 (N_13896,N_13162,N_13287);
or U13897 (N_13897,N_13316,N_13459);
nand U13898 (N_13898,N_13010,N_13404);
nand U13899 (N_13899,N_13119,N_13311);
xor U13900 (N_13900,N_13093,N_13296);
or U13901 (N_13901,N_13102,N_13189);
or U13902 (N_13902,N_13127,N_13154);
and U13903 (N_13903,N_13328,N_13304);
and U13904 (N_13904,N_13126,N_13421);
and U13905 (N_13905,N_13025,N_13372);
or U13906 (N_13906,N_13226,N_13484);
and U13907 (N_13907,N_13013,N_13158);
or U13908 (N_13908,N_13476,N_13038);
xnor U13909 (N_13909,N_13162,N_13200);
nand U13910 (N_13910,N_13021,N_13115);
xor U13911 (N_13911,N_13152,N_13233);
or U13912 (N_13912,N_13204,N_13057);
nor U13913 (N_13913,N_13339,N_13138);
and U13914 (N_13914,N_13273,N_13238);
nand U13915 (N_13915,N_13489,N_13124);
nand U13916 (N_13916,N_13235,N_13074);
nand U13917 (N_13917,N_13103,N_13222);
xor U13918 (N_13918,N_13240,N_13036);
nand U13919 (N_13919,N_13409,N_13375);
nor U13920 (N_13920,N_13154,N_13348);
and U13921 (N_13921,N_13180,N_13318);
nand U13922 (N_13922,N_13324,N_13040);
or U13923 (N_13923,N_13024,N_13124);
nand U13924 (N_13924,N_13277,N_13107);
or U13925 (N_13925,N_13124,N_13358);
and U13926 (N_13926,N_13432,N_13005);
nand U13927 (N_13927,N_13180,N_13345);
xor U13928 (N_13928,N_13019,N_13214);
or U13929 (N_13929,N_13376,N_13155);
and U13930 (N_13930,N_13415,N_13496);
xnor U13931 (N_13931,N_13438,N_13373);
nor U13932 (N_13932,N_13374,N_13462);
xnor U13933 (N_13933,N_13063,N_13389);
and U13934 (N_13934,N_13204,N_13164);
xnor U13935 (N_13935,N_13332,N_13386);
xnor U13936 (N_13936,N_13184,N_13198);
and U13937 (N_13937,N_13389,N_13381);
and U13938 (N_13938,N_13230,N_13270);
or U13939 (N_13939,N_13416,N_13261);
xor U13940 (N_13940,N_13123,N_13219);
nor U13941 (N_13941,N_13067,N_13350);
xor U13942 (N_13942,N_13488,N_13126);
nor U13943 (N_13943,N_13094,N_13295);
and U13944 (N_13944,N_13367,N_13003);
nand U13945 (N_13945,N_13483,N_13114);
or U13946 (N_13946,N_13201,N_13422);
nor U13947 (N_13947,N_13085,N_13355);
and U13948 (N_13948,N_13467,N_13408);
nor U13949 (N_13949,N_13336,N_13465);
or U13950 (N_13950,N_13183,N_13190);
nand U13951 (N_13951,N_13204,N_13244);
or U13952 (N_13952,N_13017,N_13264);
xnor U13953 (N_13953,N_13156,N_13479);
and U13954 (N_13954,N_13165,N_13111);
nor U13955 (N_13955,N_13444,N_13496);
xnor U13956 (N_13956,N_13155,N_13255);
or U13957 (N_13957,N_13258,N_13030);
xor U13958 (N_13958,N_13135,N_13222);
and U13959 (N_13959,N_13493,N_13381);
or U13960 (N_13960,N_13071,N_13486);
nand U13961 (N_13961,N_13459,N_13302);
nand U13962 (N_13962,N_13276,N_13345);
or U13963 (N_13963,N_13200,N_13253);
or U13964 (N_13964,N_13061,N_13383);
nand U13965 (N_13965,N_13076,N_13111);
nor U13966 (N_13966,N_13341,N_13476);
nor U13967 (N_13967,N_13004,N_13078);
nand U13968 (N_13968,N_13101,N_13492);
and U13969 (N_13969,N_13461,N_13477);
nor U13970 (N_13970,N_13028,N_13341);
and U13971 (N_13971,N_13487,N_13362);
nor U13972 (N_13972,N_13024,N_13190);
and U13973 (N_13973,N_13421,N_13332);
xnor U13974 (N_13974,N_13043,N_13451);
xnor U13975 (N_13975,N_13038,N_13195);
xor U13976 (N_13976,N_13163,N_13121);
and U13977 (N_13977,N_13097,N_13124);
nor U13978 (N_13978,N_13270,N_13387);
or U13979 (N_13979,N_13321,N_13063);
or U13980 (N_13980,N_13202,N_13472);
nand U13981 (N_13981,N_13429,N_13321);
nor U13982 (N_13982,N_13479,N_13255);
nand U13983 (N_13983,N_13416,N_13185);
or U13984 (N_13984,N_13150,N_13430);
and U13985 (N_13985,N_13101,N_13188);
nand U13986 (N_13986,N_13265,N_13152);
nor U13987 (N_13987,N_13195,N_13164);
nand U13988 (N_13988,N_13111,N_13023);
or U13989 (N_13989,N_13241,N_13230);
or U13990 (N_13990,N_13369,N_13026);
nand U13991 (N_13991,N_13408,N_13299);
and U13992 (N_13992,N_13200,N_13371);
or U13993 (N_13993,N_13254,N_13430);
or U13994 (N_13994,N_13116,N_13218);
xnor U13995 (N_13995,N_13333,N_13206);
nor U13996 (N_13996,N_13303,N_13410);
nand U13997 (N_13997,N_13444,N_13072);
nor U13998 (N_13998,N_13369,N_13279);
xor U13999 (N_13999,N_13339,N_13194);
or U14000 (N_14000,N_13616,N_13892);
or U14001 (N_14001,N_13973,N_13523);
xor U14002 (N_14002,N_13826,N_13526);
xnor U14003 (N_14003,N_13505,N_13681);
nand U14004 (N_14004,N_13545,N_13918);
xor U14005 (N_14005,N_13580,N_13860);
xor U14006 (N_14006,N_13634,N_13613);
xor U14007 (N_14007,N_13666,N_13902);
or U14008 (N_14008,N_13956,N_13875);
nand U14009 (N_14009,N_13767,N_13774);
nor U14010 (N_14010,N_13736,N_13727);
xor U14011 (N_14011,N_13869,N_13661);
nor U14012 (N_14012,N_13744,N_13565);
nor U14013 (N_14013,N_13962,N_13808);
nor U14014 (N_14014,N_13998,N_13608);
xnor U14015 (N_14015,N_13656,N_13582);
and U14016 (N_14016,N_13759,N_13995);
nand U14017 (N_14017,N_13805,N_13802);
xnor U14018 (N_14018,N_13702,N_13695);
or U14019 (N_14019,N_13894,N_13690);
nor U14020 (N_14020,N_13692,N_13859);
nand U14021 (N_14021,N_13618,N_13972);
and U14022 (N_14022,N_13612,N_13974);
nand U14023 (N_14023,N_13701,N_13551);
and U14024 (N_14024,N_13778,N_13528);
and U14025 (N_14025,N_13696,N_13668);
and U14026 (N_14026,N_13984,N_13575);
and U14027 (N_14027,N_13753,N_13558);
or U14028 (N_14028,N_13627,N_13828);
and U14029 (N_14029,N_13733,N_13831);
nor U14030 (N_14030,N_13748,N_13585);
or U14031 (N_14031,N_13760,N_13939);
xnor U14032 (N_14032,N_13851,N_13581);
or U14033 (N_14033,N_13694,N_13586);
or U14034 (N_14034,N_13504,N_13691);
and U14035 (N_14035,N_13795,N_13550);
or U14036 (N_14036,N_13710,N_13509);
nor U14037 (N_14037,N_13963,N_13740);
or U14038 (N_14038,N_13532,N_13573);
and U14039 (N_14039,N_13643,N_13849);
and U14040 (N_14040,N_13810,N_13923);
or U14041 (N_14041,N_13556,N_13951);
xnor U14042 (N_14042,N_13986,N_13823);
nand U14043 (N_14043,N_13960,N_13857);
xor U14044 (N_14044,N_13780,N_13850);
or U14045 (N_14045,N_13728,N_13641);
or U14046 (N_14046,N_13978,N_13819);
xor U14047 (N_14047,N_13766,N_13721);
xnor U14048 (N_14048,N_13913,N_13830);
and U14049 (N_14049,N_13846,N_13662);
nand U14050 (N_14050,N_13834,N_13822);
xor U14051 (N_14051,N_13703,N_13909);
and U14052 (N_14052,N_13757,N_13655);
xnor U14053 (N_14053,N_13679,N_13779);
nor U14054 (N_14054,N_13711,N_13862);
nand U14055 (N_14055,N_13506,N_13966);
or U14056 (N_14056,N_13976,N_13597);
nand U14057 (N_14057,N_13867,N_13631);
xor U14058 (N_14058,N_13591,N_13642);
nand U14059 (N_14059,N_13958,N_13595);
or U14060 (N_14060,N_13969,N_13572);
and U14061 (N_14061,N_13599,N_13633);
or U14062 (N_14062,N_13650,N_13559);
or U14063 (N_14063,N_13997,N_13699);
or U14064 (N_14064,N_13855,N_13989);
nor U14065 (N_14065,N_13878,N_13932);
or U14066 (N_14066,N_13950,N_13929);
nor U14067 (N_14067,N_13578,N_13538);
nor U14068 (N_14068,N_13947,N_13835);
and U14069 (N_14069,N_13773,N_13571);
nor U14070 (N_14070,N_13786,N_13790);
and U14071 (N_14071,N_13503,N_13924);
nand U14072 (N_14072,N_13907,N_13563);
nor U14073 (N_14073,N_13874,N_13953);
or U14074 (N_14074,N_13747,N_13734);
nor U14075 (N_14075,N_13754,N_13732);
or U14076 (N_14076,N_13886,N_13665);
and U14077 (N_14077,N_13873,N_13501);
nand U14078 (N_14078,N_13521,N_13516);
nand U14079 (N_14079,N_13657,N_13787);
nor U14080 (N_14080,N_13741,N_13916);
and U14081 (N_14081,N_13856,N_13629);
nor U14082 (N_14082,N_13970,N_13900);
xnor U14083 (N_14083,N_13583,N_13917);
nand U14084 (N_14084,N_13776,N_13912);
and U14085 (N_14085,N_13698,N_13725);
nand U14086 (N_14086,N_13716,N_13833);
nor U14087 (N_14087,N_13513,N_13925);
or U14088 (N_14088,N_13649,N_13872);
and U14089 (N_14089,N_13793,N_13530);
xor U14090 (N_14090,N_13821,N_13884);
nand U14091 (N_14091,N_13659,N_13731);
nand U14092 (N_14092,N_13714,N_13677);
and U14093 (N_14093,N_13965,N_13600);
nor U14094 (N_14094,N_13535,N_13804);
nand U14095 (N_14095,N_13593,N_13844);
nor U14096 (N_14096,N_13782,N_13824);
or U14097 (N_14097,N_13686,N_13680);
nand U14098 (N_14098,N_13983,N_13682);
nand U14099 (N_14099,N_13982,N_13660);
nand U14100 (N_14100,N_13549,N_13635);
and U14101 (N_14101,N_13652,N_13626);
nand U14102 (N_14102,N_13930,N_13993);
xor U14103 (N_14103,N_13933,N_13981);
nand U14104 (N_14104,N_13937,N_13683);
or U14105 (N_14105,N_13697,N_13945);
xnor U14106 (N_14106,N_13737,N_13743);
or U14107 (N_14107,N_13858,N_13817);
xor U14108 (N_14108,N_13547,N_13534);
xor U14109 (N_14109,N_13529,N_13533);
or U14110 (N_14110,N_13606,N_13898);
nand U14111 (N_14111,N_13895,N_13531);
nand U14112 (N_14112,N_13796,N_13584);
nand U14113 (N_14113,N_13864,N_13605);
xnor U14114 (N_14114,N_13887,N_13685);
nand U14115 (N_14115,N_13771,N_13765);
or U14116 (N_14116,N_13836,N_13646);
nand U14117 (N_14117,N_13919,N_13619);
and U14118 (N_14118,N_13783,N_13624);
nand U14119 (N_14119,N_13815,N_13706);
nor U14120 (N_14120,N_13746,N_13617);
nand U14121 (N_14121,N_13952,N_13964);
nor U14122 (N_14122,N_13684,N_13664);
and U14123 (N_14123,N_13994,N_13752);
xor U14124 (N_14124,N_13724,N_13514);
and U14125 (N_14125,N_13921,N_13901);
nor U14126 (N_14126,N_13904,N_13673);
and U14127 (N_14127,N_13968,N_13825);
or U14128 (N_14128,N_13812,N_13502);
nand U14129 (N_14129,N_13798,N_13590);
nand U14130 (N_14130,N_13676,N_13893);
nor U14131 (N_14131,N_13770,N_13853);
and U14132 (N_14132,N_13996,N_13906);
nor U14133 (N_14133,N_13675,N_13512);
or U14134 (N_14134,N_13990,N_13881);
nand U14135 (N_14135,N_13543,N_13651);
nor U14136 (N_14136,N_13941,N_13999);
nor U14137 (N_14137,N_13623,N_13839);
or U14138 (N_14138,N_13566,N_13899);
xnor U14139 (N_14139,N_13596,N_13720);
nor U14140 (N_14140,N_13557,N_13561);
and U14141 (N_14141,N_13840,N_13868);
and U14142 (N_14142,N_13519,N_13761);
nor U14143 (N_14143,N_13722,N_13576);
and U14144 (N_14144,N_13838,N_13877);
xor U14145 (N_14145,N_13940,N_13520);
nor U14146 (N_14146,N_13789,N_13546);
nor U14147 (N_14147,N_13946,N_13942);
nand U14148 (N_14148,N_13614,N_13562);
nand U14149 (N_14149,N_13570,N_13926);
nor U14150 (N_14150,N_13890,N_13671);
nor U14151 (N_14151,N_13517,N_13645);
or U14152 (N_14152,N_13791,N_13943);
nand U14153 (N_14153,N_13669,N_13922);
or U14154 (N_14154,N_13587,N_13977);
nor U14155 (N_14155,N_13837,N_13522);
xor U14156 (N_14156,N_13717,N_13814);
xor U14157 (N_14157,N_13980,N_13750);
xor U14158 (N_14158,N_13979,N_13644);
xnor U14159 (N_14159,N_13949,N_13525);
or U14160 (N_14160,N_13708,N_13865);
and U14161 (N_14161,N_13967,N_13621);
and U14162 (N_14162,N_13553,N_13735);
xnor U14163 (N_14163,N_13674,N_13755);
xor U14164 (N_14164,N_13935,N_13807);
or U14165 (N_14165,N_13764,N_13891);
or U14166 (N_14166,N_13961,N_13672);
xnor U14167 (N_14167,N_13800,N_13920);
xnor U14168 (N_14168,N_13985,N_13647);
xnor U14169 (N_14169,N_13832,N_13507);
or U14170 (N_14170,N_13866,N_13914);
and U14171 (N_14171,N_13630,N_13663);
xor U14172 (N_14172,N_13537,N_13511);
xor U14173 (N_14173,N_13738,N_13542);
xnor U14174 (N_14174,N_13745,N_13987);
and U14175 (N_14175,N_13622,N_13871);
nor U14176 (N_14176,N_13667,N_13615);
nand U14177 (N_14177,N_13718,N_13688);
xnor U14178 (N_14178,N_13607,N_13510);
or U14179 (N_14179,N_13848,N_13620);
nand U14180 (N_14180,N_13876,N_13775);
and U14181 (N_14181,N_13948,N_13792);
and U14182 (N_14182,N_13577,N_13628);
or U14183 (N_14183,N_13555,N_13648);
or U14184 (N_14184,N_13713,N_13707);
nand U14185 (N_14185,N_13784,N_13625);
or U14186 (N_14186,N_13632,N_13957);
xnor U14187 (N_14187,N_13944,N_13845);
xor U14188 (N_14188,N_13678,N_13730);
nand U14189 (N_14189,N_13579,N_13910);
xnor U14190 (N_14190,N_13729,N_13589);
nand U14191 (N_14191,N_13689,N_13539);
nand U14192 (N_14192,N_13809,N_13975);
and U14193 (N_14193,N_13726,N_13544);
or U14194 (N_14194,N_13540,N_13653);
xnor U14195 (N_14195,N_13554,N_13803);
nor U14196 (N_14196,N_13794,N_13971);
nand U14197 (N_14197,N_13654,N_13888);
or U14198 (N_14198,N_13785,N_13936);
nor U14199 (N_14199,N_13954,N_13749);
nand U14200 (N_14200,N_13594,N_13799);
or U14201 (N_14201,N_13806,N_13638);
or U14202 (N_14202,N_13788,N_13991);
nor U14203 (N_14203,N_13700,N_13604);
xnor U14204 (N_14204,N_13811,N_13777);
and U14205 (N_14205,N_13911,N_13854);
xnor U14206 (N_14206,N_13598,N_13928);
nand U14207 (N_14207,N_13541,N_13897);
and U14208 (N_14208,N_13863,N_13903);
and U14209 (N_14209,N_13885,N_13843);
and U14210 (N_14210,N_13801,N_13818);
or U14211 (N_14211,N_13568,N_13762);
and U14212 (N_14212,N_13781,N_13719);
or U14213 (N_14213,N_13518,N_13959);
or U14214 (N_14214,N_13847,N_13829);
and U14215 (N_14215,N_13955,N_13603);
nand U14216 (N_14216,N_13569,N_13601);
or U14217 (N_14217,N_13889,N_13915);
nand U14218 (N_14218,N_13592,N_13739);
nand U14219 (N_14219,N_13564,N_13609);
and U14220 (N_14220,N_13709,N_13879);
nor U14221 (N_14221,N_13934,N_13905);
xnor U14222 (N_14222,N_13693,N_13552);
or U14223 (N_14223,N_13880,N_13797);
nor U14224 (N_14224,N_13670,N_13756);
nor U14225 (N_14225,N_13882,N_13640);
or U14226 (N_14226,N_13567,N_13896);
and U14227 (N_14227,N_13938,N_13758);
xnor U14228 (N_14228,N_13813,N_13524);
or U14229 (N_14229,N_13527,N_13560);
or U14230 (N_14230,N_13723,N_13841);
xor U14231 (N_14231,N_13742,N_13763);
xnor U14232 (N_14232,N_13769,N_13820);
xor U14233 (N_14233,N_13610,N_13772);
nor U14234 (N_14234,N_13715,N_13636);
nand U14235 (N_14235,N_13637,N_13658);
nor U14236 (N_14236,N_13548,N_13816);
xnor U14237 (N_14237,N_13992,N_13602);
or U14238 (N_14238,N_13588,N_13500);
nor U14239 (N_14239,N_13639,N_13508);
and U14240 (N_14240,N_13768,N_13883);
xor U14241 (N_14241,N_13515,N_13931);
nor U14242 (N_14242,N_13852,N_13712);
or U14243 (N_14243,N_13827,N_13687);
nor U14244 (N_14244,N_13842,N_13927);
xor U14245 (N_14245,N_13704,N_13908);
nor U14246 (N_14246,N_13751,N_13705);
and U14247 (N_14247,N_13861,N_13870);
and U14248 (N_14248,N_13574,N_13611);
and U14249 (N_14249,N_13536,N_13988);
or U14250 (N_14250,N_13899,N_13891);
xor U14251 (N_14251,N_13714,N_13587);
nor U14252 (N_14252,N_13849,N_13798);
nor U14253 (N_14253,N_13723,N_13789);
xnor U14254 (N_14254,N_13503,N_13905);
or U14255 (N_14255,N_13529,N_13858);
xor U14256 (N_14256,N_13941,N_13791);
or U14257 (N_14257,N_13804,N_13644);
or U14258 (N_14258,N_13556,N_13670);
and U14259 (N_14259,N_13878,N_13723);
nor U14260 (N_14260,N_13712,N_13813);
or U14261 (N_14261,N_13983,N_13910);
nand U14262 (N_14262,N_13556,N_13980);
nand U14263 (N_14263,N_13869,N_13749);
and U14264 (N_14264,N_13995,N_13692);
and U14265 (N_14265,N_13801,N_13573);
or U14266 (N_14266,N_13501,N_13655);
xnor U14267 (N_14267,N_13914,N_13759);
nor U14268 (N_14268,N_13718,N_13924);
nand U14269 (N_14269,N_13672,N_13741);
and U14270 (N_14270,N_13806,N_13991);
nor U14271 (N_14271,N_13930,N_13752);
or U14272 (N_14272,N_13664,N_13748);
and U14273 (N_14273,N_13981,N_13924);
nand U14274 (N_14274,N_13736,N_13672);
nand U14275 (N_14275,N_13978,N_13797);
nand U14276 (N_14276,N_13860,N_13969);
nor U14277 (N_14277,N_13551,N_13901);
nor U14278 (N_14278,N_13528,N_13700);
nand U14279 (N_14279,N_13712,N_13690);
nor U14280 (N_14280,N_13751,N_13682);
or U14281 (N_14281,N_13623,N_13868);
nand U14282 (N_14282,N_13988,N_13960);
nor U14283 (N_14283,N_13984,N_13573);
and U14284 (N_14284,N_13979,N_13713);
or U14285 (N_14285,N_13840,N_13998);
xnor U14286 (N_14286,N_13846,N_13504);
or U14287 (N_14287,N_13817,N_13952);
xor U14288 (N_14288,N_13671,N_13896);
and U14289 (N_14289,N_13845,N_13599);
and U14290 (N_14290,N_13770,N_13561);
nor U14291 (N_14291,N_13920,N_13822);
or U14292 (N_14292,N_13986,N_13687);
or U14293 (N_14293,N_13504,N_13532);
nor U14294 (N_14294,N_13991,N_13616);
xor U14295 (N_14295,N_13919,N_13681);
xor U14296 (N_14296,N_13597,N_13878);
or U14297 (N_14297,N_13942,N_13524);
and U14298 (N_14298,N_13888,N_13942);
xor U14299 (N_14299,N_13852,N_13718);
or U14300 (N_14300,N_13829,N_13792);
nand U14301 (N_14301,N_13687,N_13857);
or U14302 (N_14302,N_13613,N_13791);
and U14303 (N_14303,N_13548,N_13715);
nand U14304 (N_14304,N_13660,N_13945);
or U14305 (N_14305,N_13921,N_13757);
xnor U14306 (N_14306,N_13940,N_13723);
nand U14307 (N_14307,N_13800,N_13673);
nor U14308 (N_14308,N_13571,N_13613);
nor U14309 (N_14309,N_13605,N_13885);
xnor U14310 (N_14310,N_13976,N_13672);
xnor U14311 (N_14311,N_13779,N_13686);
nor U14312 (N_14312,N_13638,N_13633);
nor U14313 (N_14313,N_13714,N_13874);
or U14314 (N_14314,N_13806,N_13681);
and U14315 (N_14315,N_13830,N_13664);
nand U14316 (N_14316,N_13654,N_13733);
xor U14317 (N_14317,N_13730,N_13997);
nand U14318 (N_14318,N_13867,N_13780);
and U14319 (N_14319,N_13820,N_13527);
nand U14320 (N_14320,N_13880,N_13910);
and U14321 (N_14321,N_13657,N_13746);
and U14322 (N_14322,N_13607,N_13897);
xnor U14323 (N_14323,N_13712,N_13907);
nand U14324 (N_14324,N_13966,N_13732);
xor U14325 (N_14325,N_13875,N_13542);
nor U14326 (N_14326,N_13578,N_13884);
xor U14327 (N_14327,N_13572,N_13852);
nand U14328 (N_14328,N_13509,N_13618);
nand U14329 (N_14329,N_13542,N_13906);
and U14330 (N_14330,N_13628,N_13632);
and U14331 (N_14331,N_13601,N_13696);
or U14332 (N_14332,N_13614,N_13639);
xnor U14333 (N_14333,N_13607,N_13538);
nand U14334 (N_14334,N_13629,N_13808);
nor U14335 (N_14335,N_13706,N_13505);
nand U14336 (N_14336,N_13550,N_13910);
nor U14337 (N_14337,N_13651,N_13798);
nor U14338 (N_14338,N_13557,N_13635);
or U14339 (N_14339,N_13712,N_13877);
nand U14340 (N_14340,N_13529,N_13847);
and U14341 (N_14341,N_13854,N_13692);
nor U14342 (N_14342,N_13943,N_13774);
xnor U14343 (N_14343,N_13579,N_13665);
or U14344 (N_14344,N_13559,N_13864);
nor U14345 (N_14345,N_13509,N_13915);
nor U14346 (N_14346,N_13708,N_13696);
and U14347 (N_14347,N_13814,N_13567);
and U14348 (N_14348,N_13970,N_13565);
nor U14349 (N_14349,N_13881,N_13934);
nor U14350 (N_14350,N_13594,N_13575);
xor U14351 (N_14351,N_13921,N_13910);
and U14352 (N_14352,N_13849,N_13819);
xnor U14353 (N_14353,N_13749,N_13502);
xnor U14354 (N_14354,N_13933,N_13926);
and U14355 (N_14355,N_13761,N_13889);
nor U14356 (N_14356,N_13775,N_13615);
nor U14357 (N_14357,N_13817,N_13717);
nor U14358 (N_14358,N_13983,N_13728);
nor U14359 (N_14359,N_13526,N_13705);
and U14360 (N_14360,N_13535,N_13642);
nor U14361 (N_14361,N_13720,N_13731);
or U14362 (N_14362,N_13918,N_13832);
or U14363 (N_14363,N_13768,N_13726);
nor U14364 (N_14364,N_13672,N_13808);
or U14365 (N_14365,N_13945,N_13745);
xor U14366 (N_14366,N_13628,N_13933);
or U14367 (N_14367,N_13563,N_13654);
or U14368 (N_14368,N_13840,N_13768);
xnor U14369 (N_14369,N_13620,N_13789);
nand U14370 (N_14370,N_13731,N_13859);
and U14371 (N_14371,N_13520,N_13601);
xnor U14372 (N_14372,N_13863,N_13857);
nor U14373 (N_14373,N_13718,N_13616);
xnor U14374 (N_14374,N_13836,N_13808);
or U14375 (N_14375,N_13643,N_13972);
nor U14376 (N_14376,N_13862,N_13574);
nand U14377 (N_14377,N_13826,N_13577);
nor U14378 (N_14378,N_13948,N_13510);
nand U14379 (N_14379,N_13776,N_13680);
and U14380 (N_14380,N_13798,N_13605);
or U14381 (N_14381,N_13899,N_13573);
and U14382 (N_14382,N_13925,N_13743);
xnor U14383 (N_14383,N_13910,N_13947);
nor U14384 (N_14384,N_13885,N_13529);
nor U14385 (N_14385,N_13848,N_13867);
and U14386 (N_14386,N_13761,N_13881);
and U14387 (N_14387,N_13640,N_13734);
and U14388 (N_14388,N_13735,N_13760);
xor U14389 (N_14389,N_13710,N_13750);
nand U14390 (N_14390,N_13886,N_13947);
nor U14391 (N_14391,N_13845,N_13832);
and U14392 (N_14392,N_13811,N_13509);
nor U14393 (N_14393,N_13927,N_13719);
nor U14394 (N_14394,N_13636,N_13952);
or U14395 (N_14395,N_13527,N_13985);
nand U14396 (N_14396,N_13769,N_13828);
and U14397 (N_14397,N_13605,N_13575);
and U14398 (N_14398,N_13720,N_13868);
nor U14399 (N_14399,N_13873,N_13686);
and U14400 (N_14400,N_13973,N_13694);
or U14401 (N_14401,N_13780,N_13866);
xnor U14402 (N_14402,N_13860,N_13914);
and U14403 (N_14403,N_13830,N_13815);
xor U14404 (N_14404,N_13751,N_13927);
nand U14405 (N_14405,N_13814,N_13793);
nor U14406 (N_14406,N_13551,N_13544);
or U14407 (N_14407,N_13941,N_13546);
xnor U14408 (N_14408,N_13735,N_13931);
nand U14409 (N_14409,N_13733,N_13861);
xor U14410 (N_14410,N_13975,N_13856);
nor U14411 (N_14411,N_13519,N_13789);
or U14412 (N_14412,N_13678,N_13863);
or U14413 (N_14413,N_13514,N_13909);
or U14414 (N_14414,N_13914,N_13853);
or U14415 (N_14415,N_13884,N_13955);
and U14416 (N_14416,N_13598,N_13581);
xnor U14417 (N_14417,N_13553,N_13801);
nor U14418 (N_14418,N_13646,N_13673);
or U14419 (N_14419,N_13969,N_13597);
xor U14420 (N_14420,N_13683,N_13560);
xnor U14421 (N_14421,N_13711,N_13819);
and U14422 (N_14422,N_13668,N_13809);
and U14423 (N_14423,N_13902,N_13843);
nand U14424 (N_14424,N_13940,N_13828);
and U14425 (N_14425,N_13562,N_13827);
nand U14426 (N_14426,N_13833,N_13579);
or U14427 (N_14427,N_13715,N_13880);
nand U14428 (N_14428,N_13594,N_13628);
xor U14429 (N_14429,N_13511,N_13551);
or U14430 (N_14430,N_13750,N_13717);
and U14431 (N_14431,N_13561,N_13729);
xnor U14432 (N_14432,N_13672,N_13798);
nor U14433 (N_14433,N_13686,N_13519);
or U14434 (N_14434,N_13939,N_13786);
nand U14435 (N_14435,N_13992,N_13659);
nand U14436 (N_14436,N_13713,N_13606);
xnor U14437 (N_14437,N_13906,N_13561);
xor U14438 (N_14438,N_13664,N_13864);
or U14439 (N_14439,N_13769,N_13669);
nor U14440 (N_14440,N_13905,N_13661);
and U14441 (N_14441,N_13604,N_13870);
and U14442 (N_14442,N_13826,N_13698);
nand U14443 (N_14443,N_13986,N_13612);
nor U14444 (N_14444,N_13831,N_13968);
nand U14445 (N_14445,N_13819,N_13837);
xnor U14446 (N_14446,N_13501,N_13742);
xnor U14447 (N_14447,N_13854,N_13574);
xor U14448 (N_14448,N_13675,N_13783);
nand U14449 (N_14449,N_13805,N_13587);
xnor U14450 (N_14450,N_13906,N_13695);
or U14451 (N_14451,N_13625,N_13514);
nor U14452 (N_14452,N_13965,N_13786);
nor U14453 (N_14453,N_13749,N_13999);
and U14454 (N_14454,N_13836,N_13713);
or U14455 (N_14455,N_13564,N_13614);
nor U14456 (N_14456,N_13900,N_13833);
and U14457 (N_14457,N_13910,N_13636);
xnor U14458 (N_14458,N_13901,N_13876);
xor U14459 (N_14459,N_13541,N_13804);
and U14460 (N_14460,N_13903,N_13827);
nand U14461 (N_14461,N_13521,N_13590);
or U14462 (N_14462,N_13649,N_13857);
nand U14463 (N_14463,N_13552,N_13744);
or U14464 (N_14464,N_13983,N_13530);
and U14465 (N_14465,N_13644,N_13506);
nand U14466 (N_14466,N_13836,N_13560);
nand U14467 (N_14467,N_13903,N_13528);
nor U14468 (N_14468,N_13629,N_13978);
and U14469 (N_14469,N_13509,N_13866);
nand U14470 (N_14470,N_13803,N_13595);
and U14471 (N_14471,N_13665,N_13870);
or U14472 (N_14472,N_13617,N_13504);
or U14473 (N_14473,N_13885,N_13572);
xor U14474 (N_14474,N_13803,N_13876);
nor U14475 (N_14475,N_13817,N_13799);
and U14476 (N_14476,N_13909,N_13720);
nor U14477 (N_14477,N_13549,N_13809);
nor U14478 (N_14478,N_13779,N_13518);
nand U14479 (N_14479,N_13992,N_13563);
or U14480 (N_14480,N_13810,N_13946);
nor U14481 (N_14481,N_13944,N_13858);
xnor U14482 (N_14482,N_13778,N_13816);
xnor U14483 (N_14483,N_13540,N_13888);
nor U14484 (N_14484,N_13978,N_13805);
xnor U14485 (N_14485,N_13723,N_13786);
nor U14486 (N_14486,N_13649,N_13557);
xnor U14487 (N_14487,N_13835,N_13846);
and U14488 (N_14488,N_13891,N_13679);
and U14489 (N_14489,N_13670,N_13517);
and U14490 (N_14490,N_13835,N_13721);
and U14491 (N_14491,N_13856,N_13976);
or U14492 (N_14492,N_13999,N_13864);
or U14493 (N_14493,N_13646,N_13787);
nand U14494 (N_14494,N_13704,N_13864);
or U14495 (N_14495,N_13748,N_13998);
nor U14496 (N_14496,N_13700,N_13914);
or U14497 (N_14497,N_13551,N_13648);
or U14498 (N_14498,N_13800,N_13980);
or U14499 (N_14499,N_13662,N_13657);
nand U14500 (N_14500,N_14383,N_14046);
xor U14501 (N_14501,N_14055,N_14420);
and U14502 (N_14502,N_14240,N_14411);
nand U14503 (N_14503,N_14419,N_14007);
nand U14504 (N_14504,N_14180,N_14436);
nand U14505 (N_14505,N_14076,N_14344);
and U14506 (N_14506,N_14345,N_14427);
nand U14507 (N_14507,N_14356,N_14156);
nand U14508 (N_14508,N_14278,N_14161);
or U14509 (N_14509,N_14190,N_14230);
nand U14510 (N_14510,N_14021,N_14438);
and U14511 (N_14511,N_14402,N_14410);
or U14512 (N_14512,N_14065,N_14255);
nand U14513 (N_14513,N_14243,N_14381);
and U14514 (N_14514,N_14086,N_14472);
nand U14515 (N_14515,N_14331,N_14448);
or U14516 (N_14516,N_14437,N_14263);
xnor U14517 (N_14517,N_14042,N_14132);
nand U14518 (N_14518,N_14440,N_14075);
nand U14519 (N_14519,N_14292,N_14314);
nor U14520 (N_14520,N_14144,N_14178);
nor U14521 (N_14521,N_14157,N_14128);
nand U14522 (N_14522,N_14492,N_14400);
xnor U14523 (N_14523,N_14030,N_14455);
nand U14524 (N_14524,N_14407,N_14103);
nor U14525 (N_14525,N_14223,N_14095);
and U14526 (N_14526,N_14034,N_14272);
and U14527 (N_14527,N_14110,N_14188);
nand U14528 (N_14528,N_14265,N_14122);
nor U14529 (N_14529,N_14094,N_14304);
nand U14530 (N_14530,N_14166,N_14215);
xor U14531 (N_14531,N_14357,N_14346);
nor U14532 (N_14532,N_14010,N_14111);
xor U14533 (N_14533,N_14158,N_14481);
xnor U14534 (N_14534,N_14241,N_14298);
and U14535 (N_14535,N_14315,N_14456);
or U14536 (N_14536,N_14429,N_14432);
nand U14537 (N_14537,N_14426,N_14499);
xnor U14538 (N_14538,N_14062,N_14171);
nand U14539 (N_14539,N_14350,N_14395);
and U14540 (N_14540,N_14490,N_14313);
nand U14541 (N_14541,N_14183,N_14300);
xnor U14542 (N_14542,N_14373,N_14480);
or U14543 (N_14543,N_14248,N_14113);
xor U14544 (N_14544,N_14452,N_14382);
and U14545 (N_14545,N_14323,N_14229);
or U14546 (N_14546,N_14134,N_14201);
nand U14547 (N_14547,N_14127,N_14195);
nand U14548 (N_14548,N_14031,N_14074);
or U14549 (N_14549,N_14377,N_14434);
nor U14550 (N_14550,N_14376,N_14302);
nand U14551 (N_14551,N_14468,N_14431);
nor U14552 (N_14552,N_14477,N_14203);
and U14553 (N_14553,N_14092,N_14471);
or U14554 (N_14554,N_14288,N_14151);
nand U14555 (N_14555,N_14285,N_14486);
nor U14556 (N_14556,N_14496,N_14206);
and U14557 (N_14557,N_14261,N_14406);
xnor U14558 (N_14558,N_14101,N_14318);
xnor U14559 (N_14559,N_14153,N_14238);
or U14560 (N_14560,N_14341,N_14069);
and U14561 (N_14561,N_14102,N_14038);
xnor U14562 (N_14562,N_14309,N_14317);
and U14563 (N_14563,N_14231,N_14367);
xnor U14564 (N_14564,N_14469,N_14028);
nand U14565 (N_14565,N_14416,N_14286);
or U14566 (N_14566,N_14123,N_14289);
nor U14567 (N_14567,N_14093,N_14295);
nor U14568 (N_14568,N_14077,N_14476);
or U14569 (N_14569,N_14320,N_14004);
or U14570 (N_14570,N_14297,N_14482);
or U14571 (N_14571,N_14015,N_14254);
and U14572 (N_14572,N_14061,N_14269);
or U14573 (N_14573,N_14162,N_14022);
or U14574 (N_14574,N_14019,N_14365);
nand U14575 (N_14575,N_14170,N_14305);
nand U14576 (N_14576,N_14167,N_14234);
or U14577 (N_14577,N_14488,N_14441);
xor U14578 (N_14578,N_14002,N_14033);
nand U14579 (N_14579,N_14404,N_14497);
and U14580 (N_14580,N_14032,N_14273);
xor U14581 (N_14581,N_14287,N_14369);
and U14582 (N_14582,N_14090,N_14168);
xor U14583 (N_14583,N_14275,N_14258);
or U14584 (N_14584,N_14053,N_14221);
nand U14585 (N_14585,N_14237,N_14364);
or U14586 (N_14586,N_14324,N_14462);
nor U14587 (N_14587,N_14185,N_14140);
or U14588 (N_14588,N_14164,N_14239);
and U14589 (N_14589,N_14461,N_14425);
and U14590 (N_14590,N_14299,N_14199);
or U14591 (N_14591,N_14413,N_14036);
and U14592 (N_14592,N_14041,N_14334);
and U14593 (N_14593,N_14349,N_14016);
xor U14594 (N_14594,N_14387,N_14091);
xor U14595 (N_14595,N_14388,N_14296);
nor U14596 (N_14596,N_14421,N_14085);
nand U14597 (N_14597,N_14202,N_14179);
or U14598 (N_14598,N_14114,N_14301);
nand U14599 (N_14599,N_14329,N_14154);
or U14600 (N_14600,N_14050,N_14130);
and U14601 (N_14601,N_14423,N_14037);
xnor U14602 (N_14602,N_14379,N_14175);
or U14603 (N_14603,N_14143,N_14232);
and U14604 (N_14604,N_14131,N_14217);
or U14605 (N_14605,N_14256,N_14267);
nand U14606 (N_14606,N_14212,N_14150);
or U14607 (N_14607,N_14332,N_14218);
and U14608 (N_14608,N_14129,N_14118);
xor U14609 (N_14609,N_14244,N_14057);
or U14610 (N_14610,N_14017,N_14359);
or U14611 (N_14611,N_14398,N_14080);
nand U14612 (N_14612,N_14498,N_14040);
nand U14613 (N_14613,N_14116,N_14347);
and U14614 (N_14614,N_14271,N_14354);
xor U14615 (N_14615,N_14181,N_14165);
nor U14616 (N_14616,N_14460,N_14391);
nor U14617 (N_14617,N_14049,N_14099);
nand U14618 (N_14618,N_14368,N_14467);
xnor U14619 (N_14619,N_14393,N_14339);
or U14620 (N_14620,N_14282,N_14348);
and U14621 (N_14621,N_14063,N_14182);
and U14622 (N_14622,N_14196,N_14495);
nand U14623 (N_14623,N_14408,N_14245);
or U14624 (N_14624,N_14446,N_14112);
and U14625 (N_14625,N_14013,N_14279);
or U14626 (N_14626,N_14281,N_14358);
nor U14627 (N_14627,N_14378,N_14204);
xor U14628 (N_14628,N_14264,N_14430);
nor U14629 (N_14629,N_14355,N_14072);
nor U14630 (N_14630,N_14253,N_14280);
and U14631 (N_14631,N_14048,N_14216);
and U14632 (N_14632,N_14043,N_14336);
nand U14633 (N_14633,N_14390,N_14169);
and U14634 (N_14634,N_14056,N_14361);
nor U14635 (N_14635,N_14330,N_14186);
or U14636 (N_14636,N_14087,N_14039);
or U14637 (N_14637,N_14159,N_14242);
or U14638 (N_14638,N_14249,N_14465);
xnor U14639 (N_14639,N_14194,N_14070);
xor U14640 (N_14640,N_14403,N_14173);
and U14641 (N_14641,N_14384,N_14463);
nand U14642 (N_14642,N_14454,N_14145);
or U14643 (N_14643,N_14208,N_14172);
nor U14644 (N_14644,N_14052,N_14119);
nor U14645 (N_14645,N_14415,N_14225);
xor U14646 (N_14646,N_14227,N_14306);
nor U14647 (N_14647,N_14290,N_14401);
and U14648 (N_14648,N_14311,N_14228);
xnor U14649 (N_14649,N_14222,N_14360);
nand U14650 (N_14650,N_14374,N_14328);
nand U14651 (N_14651,N_14060,N_14139);
xnor U14652 (N_14652,N_14018,N_14136);
nand U14653 (N_14653,N_14108,N_14088);
nand U14654 (N_14654,N_14197,N_14485);
nand U14655 (N_14655,N_14489,N_14176);
nor U14656 (N_14656,N_14450,N_14079);
xnor U14657 (N_14657,N_14316,N_14433);
and U14658 (N_14658,N_14193,N_14326);
nor U14659 (N_14659,N_14200,N_14372);
xnor U14660 (N_14660,N_14274,N_14475);
xnor U14661 (N_14661,N_14445,N_14294);
xor U14662 (N_14662,N_14214,N_14370);
and U14663 (N_14663,N_14447,N_14308);
xor U14664 (N_14664,N_14337,N_14259);
nor U14665 (N_14665,N_14246,N_14351);
and U14666 (N_14666,N_14064,N_14014);
xor U14667 (N_14667,N_14147,N_14135);
nor U14668 (N_14668,N_14459,N_14138);
and U14669 (N_14669,N_14386,N_14284);
xnor U14670 (N_14670,N_14152,N_14453);
nor U14671 (N_14671,N_14209,N_14029);
nor U14672 (N_14672,N_14213,N_14011);
and U14673 (N_14673,N_14458,N_14124);
xor U14674 (N_14674,N_14192,N_14005);
nor U14675 (N_14675,N_14268,N_14220);
nor U14676 (N_14676,N_14117,N_14198);
nand U14677 (N_14677,N_14457,N_14397);
xnor U14678 (N_14678,N_14045,N_14371);
and U14679 (N_14679,N_14003,N_14035);
nand U14680 (N_14680,N_14148,N_14078);
and U14681 (N_14681,N_14047,N_14474);
nor U14682 (N_14682,N_14149,N_14352);
nand U14683 (N_14683,N_14435,N_14283);
nand U14684 (N_14684,N_14473,N_14266);
nand U14685 (N_14685,N_14020,N_14366);
nor U14686 (N_14686,N_14073,N_14001);
nand U14687 (N_14687,N_14068,N_14325);
and U14688 (N_14688,N_14252,N_14027);
or U14689 (N_14689,N_14418,N_14262);
or U14690 (N_14690,N_14487,N_14233);
nor U14691 (N_14691,N_14363,N_14008);
nor U14692 (N_14692,N_14470,N_14338);
xor U14693 (N_14693,N_14051,N_14303);
nor U14694 (N_14694,N_14026,N_14177);
nor U14695 (N_14695,N_14478,N_14120);
and U14696 (N_14696,N_14493,N_14219);
xor U14697 (N_14697,N_14115,N_14082);
xnor U14698 (N_14698,N_14412,N_14483);
nor U14699 (N_14699,N_14058,N_14009);
xnor U14700 (N_14700,N_14098,N_14321);
and U14701 (N_14701,N_14236,N_14442);
nand U14702 (N_14702,N_14141,N_14044);
nand U14703 (N_14703,N_14121,N_14422);
and U14704 (N_14704,N_14466,N_14399);
nand U14705 (N_14705,N_14409,N_14067);
and U14706 (N_14706,N_14054,N_14362);
nor U14707 (N_14707,N_14333,N_14327);
nor U14708 (N_14708,N_14443,N_14439);
xor U14709 (N_14709,N_14012,N_14109);
or U14710 (N_14710,N_14071,N_14089);
and U14711 (N_14711,N_14444,N_14137);
nor U14712 (N_14712,N_14210,N_14097);
and U14713 (N_14713,N_14006,N_14396);
xnor U14714 (N_14714,N_14226,N_14310);
or U14715 (N_14715,N_14424,N_14312);
and U14716 (N_14716,N_14024,N_14133);
or U14717 (N_14717,N_14293,N_14307);
xnor U14718 (N_14718,N_14322,N_14277);
xor U14719 (N_14719,N_14146,N_14000);
and U14720 (N_14720,N_14251,N_14142);
nand U14721 (N_14721,N_14319,N_14428);
or U14722 (N_14722,N_14491,N_14449);
or U14723 (N_14723,N_14389,N_14335);
nor U14724 (N_14724,N_14081,N_14375);
or U14725 (N_14725,N_14184,N_14479);
nor U14726 (N_14726,N_14096,N_14189);
and U14727 (N_14727,N_14163,N_14207);
or U14728 (N_14728,N_14224,N_14494);
and U14729 (N_14729,N_14023,N_14107);
nor U14730 (N_14730,N_14270,N_14250);
nand U14731 (N_14731,N_14191,N_14340);
nand U14732 (N_14732,N_14291,N_14394);
xor U14733 (N_14733,N_14126,N_14025);
nand U14734 (N_14734,N_14417,N_14380);
nand U14735 (N_14735,N_14160,N_14187);
and U14736 (N_14736,N_14342,N_14392);
or U14737 (N_14737,N_14100,N_14257);
and U14738 (N_14738,N_14084,N_14260);
or U14739 (N_14739,N_14414,N_14235);
nand U14740 (N_14740,N_14106,N_14105);
and U14741 (N_14741,N_14211,N_14276);
nor U14742 (N_14742,N_14405,N_14464);
nand U14743 (N_14743,N_14484,N_14125);
or U14744 (N_14744,N_14451,N_14066);
xor U14745 (N_14745,N_14247,N_14083);
and U14746 (N_14746,N_14059,N_14343);
nor U14747 (N_14747,N_14353,N_14155);
xnor U14748 (N_14748,N_14205,N_14104);
nand U14749 (N_14749,N_14174,N_14385);
xnor U14750 (N_14750,N_14212,N_14354);
nand U14751 (N_14751,N_14285,N_14012);
nand U14752 (N_14752,N_14047,N_14428);
nand U14753 (N_14753,N_14040,N_14379);
nand U14754 (N_14754,N_14391,N_14411);
nor U14755 (N_14755,N_14224,N_14052);
or U14756 (N_14756,N_14187,N_14024);
nand U14757 (N_14757,N_14324,N_14173);
and U14758 (N_14758,N_14472,N_14312);
nand U14759 (N_14759,N_14108,N_14005);
nand U14760 (N_14760,N_14440,N_14153);
and U14761 (N_14761,N_14233,N_14117);
nor U14762 (N_14762,N_14182,N_14215);
or U14763 (N_14763,N_14393,N_14026);
or U14764 (N_14764,N_14088,N_14045);
nor U14765 (N_14765,N_14353,N_14074);
or U14766 (N_14766,N_14058,N_14394);
or U14767 (N_14767,N_14183,N_14216);
nand U14768 (N_14768,N_14497,N_14475);
or U14769 (N_14769,N_14077,N_14264);
and U14770 (N_14770,N_14100,N_14443);
or U14771 (N_14771,N_14249,N_14357);
or U14772 (N_14772,N_14453,N_14169);
nor U14773 (N_14773,N_14401,N_14218);
nor U14774 (N_14774,N_14334,N_14435);
and U14775 (N_14775,N_14439,N_14490);
nor U14776 (N_14776,N_14347,N_14257);
or U14777 (N_14777,N_14178,N_14237);
or U14778 (N_14778,N_14113,N_14021);
or U14779 (N_14779,N_14027,N_14297);
and U14780 (N_14780,N_14307,N_14130);
nor U14781 (N_14781,N_14471,N_14099);
xor U14782 (N_14782,N_14360,N_14263);
or U14783 (N_14783,N_14442,N_14301);
and U14784 (N_14784,N_14286,N_14187);
or U14785 (N_14785,N_14437,N_14136);
nor U14786 (N_14786,N_14419,N_14342);
nand U14787 (N_14787,N_14210,N_14429);
and U14788 (N_14788,N_14372,N_14146);
xnor U14789 (N_14789,N_14385,N_14263);
and U14790 (N_14790,N_14001,N_14150);
or U14791 (N_14791,N_14092,N_14076);
nor U14792 (N_14792,N_14184,N_14363);
or U14793 (N_14793,N_14236,N_14418);
nand U14794 (N_14794,N_14119,N_14397);
nor U14795 (N_14795,N_14379,N_14250);
and U14796 (N_14796,N_14413,N_14196);
xnor U14797 (N_14797,N_14150,N_14409);
nand U14798 (N_14798,N_14274,N_14489);
or U14799 (N_14799,N_14303,N_14206);
and U14800 (N_14800,N_14018,N_14317);
nand U14801 (N_14801,N_14285,N_14133);
and U14802 (N_14802,N_14152,N_14094);
xor U14803 (N_14803,N_14015,N_14104);
xor U14804 (N_14804,N_14321,N_14424);
xnor U14805 (N_14805,N_14142,N_14455);
nor U14806 (N_14806,N_14267,N_14320);
nor U14807 (N_14807,N_14302,N_14320);
xnor U14808 (N_14808,N_14482,N_14115);
nand U14809 (N_14809,N_14449,N_14158);
or U14810 (N_14810,N_14333,N_14332);
or U14811 (N_14811,N_14430,N_14439);
or U14812 (N_14812,N_14409,N_14002);
or U14813 (N_14813,N_14212,N_14074);
and U14814 (N_14814,N_14256,N_14070);
xnor U14815 (N_14815,N_14037,N_14005);
nor U14816 (N_14816,N_14284,N_14206);
or U14817 (N_14817,N_14093,N_14455);
xor U14818 (N_14818,N_14385,N_14002);
xor U14819 (N_14819,N_14246,N_14449);
xor U14820 (N_14820,N_14269,N_14127);
nand U14821 (N_14821,N_14261,N_14227);
nand U14822 (N_14822,N_14262,N_14294);
and U14823 (N_14823,N_14396,N_14180);
or U14824 (N_14824,N_14000,N_14353);
and U14825 (N_14825,N_14443,N_14352);
or U14826 (N_14826,N_14256,N_14193);
xnor U14827 (N_14827,N_14353,N_14306);
nor U14828 (N_14828,N_14268,N_14190);
xor U14829 (N_14829,N_14044,N_14397);
nand U14830 (N_14830,N_14411,N_14104);
nor U14831 (N_14831,N_14458,N_14154);
nand U14832 (N_14832,N_14497,N_14012);
xor U14833 (N_14833,N_14320,N_14094);
nor U14834 (N_14834,N_14402,N_14123);
and U14835 (N_14835,N_14441,N_14231);
and U14836 (N_14836,N_14252,N_14228);
or U14837 (N_14837,N_14188,N_14495);
and U14838 (N_14838,N_14232,N_14112);
nor U14839 (N_14839,N_14323,N_14439);
and U14840 (N_14840,N_14428,N_14322);
nand U14841 (N_14841,N_14393,N_14478);
and U14842 (N_14842,N_14320,N_14120);
nand U14843 (N_14843,N_14050,N_14376);
or U14844 (N_14844,N_14308,N_14278);
xnor U14845 (N_14845,N_14466,N_14167);
and U14846 (N_14846,N_14249,N_14121);
xor U14847 (N_14847,N_14063,N_14443);
or U14848 (N_14848,N_14315,N_14140);
or U14849 (N_14849,N_14364,N_14415);
or U14850 (N_14850,N_14224,N_14092);
nand U14851 (N_14851,N_14414,N_14384);
nor U14852 (N_14852,N_14481,N_14126);
nor U14853 (N_14853,N_14497,N_14329);
and U14854 (N_14854,N_14088,N_14071);
nand U14855 (N_14855,N_14098,N_14018);
and U14856 (N_14856,N_14405,N_14096);
or U14857 (N_14857,N_14123,N_14455);
nand U14858 (N_14858,N_14126,N_14385);
or U14859 (N_14859,N_14209,N_14232);
xnor U14860 (N_14860,N_14264,N_14057);
or U14861 (N_14861,N_14167,N_14250);
and U14862 (N_14862,N_14423,N_14007);
or U14863 (N_14863,N_14406,N_14401);
and U14864 (N_14864,N_14198,N_14099);
xnor U14865 (N_14865,N_14372,N_14178);
nand U14866 (N_14866,N_14455,N_14495);
and U14867 (N_14867,N_14008,N_14404);
nor U14868 (N_14868,N_14481,N_14427);
and U14869 (N_14869,N_14428,N_14191);
nand U14870 (N_14870,N_14428,N_14230);
nand U14871 (N_14871,N_14322,N_14127);
nand U14872 (N_14872,N_14474,N_14091);
and U14873 (N_14873,N_14045,N_14489);
and U14874 (N_14874,N_14334,N_14368);
xnor U14875 (N_14875,N_14461,N_14446);
or U14876 (N_14876,N_14069,N_14403);
xnor U14877 (N_14877,N_14210,N_14137);
xor U14878 (N_14878,N_14284,N_14058);
nor U14879 (N_14879,N_14344,N_14445);
nand U14880 (N_14880,N_14495,N_14296);
and U14881 (N_14881,N_14140,N_14423);
nand U14882 (N_14882,N_14275,N_14396);
or U14883 (N_14883,N_14179,N_14391);
nor U14884 (N_14884,N_14337,N_14013);
nor U14885 (N_14885,N_14361,N_14087);
and U14886 (N_14886,N_14273,N_14126);
nor U14887 (N_14887,N_14363,N_14051);
or U14888 (N_14888,N_14079,N_14422);
nor U14889 (N_14889,N_14288,N_14367);
nand U14890 (N_14890,N_14273,N_14485);
nor U14891 (N_14891,N_14460,N_14443);
xor U14892 (N_14892,N_14467,N_14261);
nor U14893 (N_14893,N_14012,N_14078);
nand U14894 (N_14894,N_14032,N_14241);
nand U14895 (N_14895,N_14133,N_14213);
and U14896 (N_14896,N_14030,N_14116);
nor U14897 (N_14897,N_14305,N_14064);
and U14898 (N_14898,N_14013,N_14153);
nor U14899 (N_14899,N_14096,N_14267);
nor U14900 (N_14900,N_14412,N_14039);
xor U14901 (N_14901,N_14249,N_14093);
or U14902 (N_14902,N_14003,N_14145);
xnor U14903 (N_14903,N_14076,N_14228);
xor U14904 (N_14904,N_14118,N_14321);
xor U14905 (N_14905,N_14421,N_14341);
or U14906 (N_14906,N_14253,N_14261);
xnor U14907 (N_14907,N_14404,N_14426);
nor U14908 (N_14908,N_14325,N_14087);
nand U14909 (N_14909,N_14361,N_14342);
or U14910 (N_14910,N_14145,N_14032);
or U14911 (N_14911,N_14008,N_14036);
nand U14912 (N_14912,N_14350,N_14180);
xor U14913 (N_14913,N_14489,N_14117);
or U14914 (N_14914,N_14222,N_14299);
nor U14915 (N_14915,N_14483,N_14067);
xnor U14916 (N_14916,N_14210,N_14231);
nand U14917 (N_14917,N_14199,N_14495);
and U14918 (N_14918,N_14189,N_14454);
nand U14919 (N_14919,N_14064,N_14081);
or U14920 (N_14920,N_14297,N_14009);
and U14921 (N_14921,N_14412,N_14473);
or U14922 (N_14922,N_14093,N_14470);
or U14923 (N_14923,N_14043,N_14161);
or U14924 (N_14924,N_14302,N_14307);
nand U14925 (N_14925,N_14334,N_14247);
nand U14926 (N_14926,N_14039,N_14071);
nand U14927 (N_14927,N_14321,N_14081);
or U14928 (N_14928,N_14483,N_14162);
nand U14929 (N_14929,N_14144,N_14279);
nor U14930 (N_14930,N_14112,N_14196);
nand U14931 (N_14931,N_14091,N_14284);
xnor U14932 (N_14932,N_14401,N_14350);
xor U14933 (N_14933,N_14264,N_14384);
or U14934 (N_14934,N_14165,N_14024);
nand U14935 (N_14935,N_14308,N_14390);
nor U14936 (N_14936,N_14497,N_14308);
nand U14937 (N_14937,N_14338,N_14397);
and U14938 (N_14938,N_14361,N_14121);
nand U14939 (N_14939,N_14101,N_14274);
xnor U14940 (N_14940,N_14424,N_14143);
nor U14941 (N_14941,N_14025,N_14052);
xor U14942 (N_14942,N_14349,N_14051);
xnor U14943 (N_14943,N_14275,N_14095);
nand U14944 (N_14944,N_14365,N_14026);
and U14945 (N_14945,N_14376,N_14098);
nand U14946 (N_14946,N_14301,N_14263);
xnor U14947 (N_14947,N_14387,N_14453);
nor U14948 (N_14948,N_14015,N_14058);
and U14949 (N_14949,N_14394,N_14156);
nand U14950 (N_14950,N_14330,N_14301);
and U14951 (N_14951,N_14062,N_14221);
nor U14952 (N_14952,N_14314,N_14214);
and U14953 (N_14953,N_14270,N_14093);
xnor U14954 (N_14954,N_14263,N_14123);
nor U14955 (N_14955,N_14448,N_14369);
and U14956 (N_14956,N_14375,N_14487);
nor U14957 (N_14957,N_14003,N_14174);
and U14958 (N_14958,N_14400,N_14056);
nand U14959 (N_14959,N_14082,N_14179);
nand U14960 (N_14960,N_14207,N_14208);
or U14961 (N_14961,N_14191,N_14020);
xnor U14962 (N_14962,N_14335,N_14270);
xor U14963 (N_14963,N_14245,N_14353);
and U14964 (N_14964,N_14249,N_14355);
xor U14965 (N_14965,N_14359,N_14433);
nor U14966 (N_14966,N_14224,N_14397);
xnor U14967 (N_14967,N_14113,N_14345);
nand U14968 (N_14968,N_14003,N_14109);
nand U14969 (N_14969,N_14076,N_14244);
and U14970 (N_14970,N_14416,N_14437);
nand U14971 (N_14971,N_14415,N_14403);
nand U14972 (N_14972,N_14235,N_14384);
nand U14973 (N_14973,N_14187,N_14240);
nand U14974 (N_14974,N_14436,N_14191);
nor U14975 (N_14975,N_14304,N_14068);
xnor U14976 (N_14976,N_14320,N_14342);
xnor U14977 (N_14977,N_14253,N_14115);
and U14978 (N_14978,N_14483,N_14382);
nor U14979 (N_14979,N_14156,N_14206);
or U14980 (N_14980,N_14015,N_14493);
nor U14981 (N_14981,N_14147,N_14385);
nor U14982 (N_14982,N_14163,N_14350);
nor U14983 (N_14983,N_14310,N_14316);
xnor U14984 (N_14984,N_14335,N_14319);
xor U14985 (N_14985,N_14096,N_14094);
or U14986 (N_14986,N_14113,N_14177);
nor U14987 (N_14987,N_14102,N_14180);
nand U14988 (N_14988,N_14103,N_14093);
xnor U14989 (N_14989,N_14209,N_14169);
nand U14990 (N_14990,N_14301,N_14274);
nor U14991 (N_14991,N_14483,N_14424);
nand U14992 (N_14992,N_14212,N_14376);
and U14993 (N_14993,N_14292,N_14173);
nand U14994 (N_14994,N_14318,N_14140);
nor U14995 (N_14995,N_14344,N_14351);
nand U14996 (N_14996,N_14359,N_14129);
and U14997 (N_14997,N_14447,N_14249);
or U14998 (N_14998,N_14488,N_14289);
or U14999 (N_14999,N_14013,N_14227);
xnor U15000 (N_15000,N_14906,N_14923);
or U15001 (N_15001,N_14978,N_14514);
xnor U15002 (N_15002,N_14811,N_14714);
nand U15003 (N_15003,N_14567,N_14931);
xnor U15004 (N_15004,N_14946,N_14684);
xor U15005 (N_15005,N_14842,N_14607);
nand U15006 (N_15006,N_14747,N_14565);
xnor U15007 (N_15007,N_14970,N_14879);
and U15008 (N_15008,N_14589,N_14550);
xnor U15009 (N_15009,N_14717,N_14955);
or U15010 (N_15010,N_14629,N_14905);
nand U15011 (N_15011,N_14705,N_14785);
nand U15012 (N_15012,N_14506,N_14536);
nand U15013 (N_15013,N_14969,N_14912);
nand U15014 (N_15014,N_14973,N_14758);
or U15015 (N_15015,N_14624,N_14633);
xor U15016 (N_15016,N_14543,N_14981);
nand U15017 (N_15017,N_14726,N_14526);
nor U15018 (N_15018,N_14582,N_14601);
nand U15019 (N_15019,N_14767,N_14549);
or U15020 (N_15020,N_14694,N_14659);
or U15021 (N_15021,N_14616,N_14824);
and U15022 (N_15022,N_14655,N_14852);
xnor U15023 (N_15023,N_14826,N_14977);
or U15024 (N_15024,N_14766,N_14701);
nand U15025 (N_15025,N_14871,N_14832);
or U15026 (N_15026,N_14604,N_14803);
nand U15027 (N_15027,N_14802,N_14516);
nor U15028 (N_15028,N_14552,N_14672);
nor U15029 (N_15029,N_14736,N_14935);
nand U15030 (N_15030,N_14892,N_14542);
xor U15031 (N_15031,N_14816,N_14927);
xnor U15032 (N_15032,N_14806,N_14630);
or U15033 (N_15033,N_14541,N_14699);
nor U15034 (N_15034,N_14687,N_14738);
or U15035 (N_15035,N_14798,N_14891);
xor U15036 (N_15036,N_14670,N_14743);
nand U15037 (N_15037,N_14606,N_14553);
or U15038 (N_15038,N_14942,N_14580);
xor U15039 (N_15039,N_14535,N_14681);
nand U15040 (N_15040,N_14799,N_14716);
xor U15041 (N_15041,N_14651,N_14609);
nor U15042 (N_15042,N_14932,N_14576);
nand U15043 (N_15043,N_14709,N_14858);
nand U15044 (N_15044,N_14857,N_14791);
nand U15045 (N_15045,N_14765,N_14654);
xnor U15046 (N_15046,N_14628,N_14943);
nand U15047 (N_15047,N_14810,N_14723);
and U15048 (N_15048,N_14784,N_14501);
and U15049 (N_15049,N_14938,N_14611);
xnor U15050 (N_15050,N_14827,N_14841);
and U15051 (N_15051,N_14886,N_14727);
nor U15052 (N_15052,N_14789,N_14911);
xor U15053 (N_15053,N_14612,N_14779);
nor U15054 (N_15054,N_14641,N_14704);
nand U15055 (N_15055,N_14960,N_14749);
or U15056 (N_15056,N_14586,N_14594);
xor U15057 (N_15057,N_14903,N_14639);
xor U15058 (N_15058,N_14623,N_14631);
xor U15059 (N_15059,N_14603,N_14861);
or U15060 (N_15060,N_14668,N_14908);
or U15061 (N_15061,N_14508,N_14708);
nor U15062 (N_15062,N_14794,N_14698);
nand U15063 (N_15063,N_14518,N_14614);
nand U15064 (N_15064,N_14529,N_14730);
nand U15065 (N_15065,N_14850,N_14894);
nor U15066 (N_15066,N_14561,N_14712);
xnor U15067 (N_15067,N_14882,N_14729);
nor U15068 (N_15068,N_14953,N_14926);
nor U15069 (N_15069,N_14674,N_14590);
xnor U15070 (N_15070,N_14657,N_14801);
nand U15071 (N_15071,N_14875,N_14665);
nor U15072 (N_15072,N_14869,N_14962);
xor U15073 (N_15073,N_14588,N_14817);
nand U15074 (N_15074,N_14989,N_14741);
nor U15075 (N_15075,N_14997,N_14814);
nor U15076 (N_15076,N_14732,N_14994);
or U15077 (N_15077,N_14921,N_14573);
and U15078 (N_15078,N_14618,N_14913);
xnor U15079 (N_15079,N_14829,N_14900);
xnor U15080 (N_15080,N_14683,N_14673);
and U15081 (N_15081,N_14933,N_14854);
nor U15082 (N_15082,N_14823,N_14809);
xor U15083 (N_15083,N_14548,N_14534);
and U15084 (N_15084,N_14795,N_14838);
xnor U15085 (N_15085,N_14507,N_14787);
and U15086 (N_15086,N_14597,N_14556);
nor U15087 (N_15087,N_14728,N_14721);
nor U15088 (N_15088,N_14980,N_14577);
or U15089 (N_15089,N_14939,N_14539);
and U15090 (N_15090,N_14936,N_14568);
nand U15091 (N_15091,N_14948,N_14650);
nor U15092 (N_15092,N_14735,N_14914);
nor U15093 (N_15093,N_14972,N_14924);
or U15094 (N_15094,N_14984,N_14621);
or U15095 (N_15095,N_14961,N_14528);
nor U15096 (N_15096,N_14523,N_14515);
nand U15097 (N_15097,N_14706,N_14746);
nand U15098 (N_15098,N_14837,N_14775);
nor U15099 (N_15099,N_14988,N_14693);
nor U15100 (N_15100,N_14663,N_14517);
xor U15101 (N_15101,N_14627,N_14622);
and U15102 (N_15102,N_14648,N_14888);
nand U15103 (N_15103,N_14700,N_14733);
nand U15104 (N_15104,N_14971,N_14881);
nand U15105 (N_15105,N_14761,N_14596);
nor U15106 (N_15106,N_14557,N_14546);
xnor U15107 (N_15107,N_14719,N_14975);
or U15108 (N_15108,N_14757,N_14748);
nor U15109 (N_15109,N_14739,N_14711);
or U15110 (N_15110,N_14918,N_14608);
and U15111 (N_15111,N_14679,N_14848);
and U15112 (N_15112,N_14992,N_14579);
and U15113 (N_15113,N_14909,N_14521);
and U15114 (N_15114,N_14689,N_14774);
xnor U15115 (N_15115,N_14602,N_14640);
or U15116 (N_15116,N_14660,N_14676);
and U15117 (N_15117,N_14707,N_14522);
xnor U15118 (N_15118,N_14725,N_14941);
or U15119 (N_15119,N_14896,N_14585);
or U15120 (N_15120,N_14985,N_14859);
nor U15121 (N_15121,N_14635,N_14560);
nor U15122 (N_15122,N_14950,N_14759);
nor U15123 (N_15123,N_14677,N_14866);
and U15124 (N_15124,N_14904,N_14537);
xor U15125 (N_15125,N_14937,N_14664);
and U15126 (N_15126,N_14790,N_14887);
or U15127 (N_15127,N_14952,N_14916);
xnor U15128 (N_15128,N_14667,N_14554);
xor U15129 (N_15129,N_14696,N_14867);
nand U15130 (N_15130,N_14532,N_14976);
and U15131 (N_15131,N_14883,N_14974);
nand U15132 (N_15132,N_14922,N_14995);
or U15133 (N_15133,N_14524,N_14617);
and U15134 (N_15134,N_14525,N_14744);
or U15135 (N_15135,N_14605,N_14919);
xor U15136 (N_15136,N_14862,N_14813);
nor U15137 (N_15137,N_14865,N_14527);
nor U15138 (N_15138,N_14956,N_14772);
nor U15139 (N_15139,N_14845,N_14807);
xor U15140 (N_15140,N_14658,N_14770);
nor U15141 (N_15141,N_14511,N_14610);
and U15142 (N_15142,N_14745,N_14513);
xnor U15143 (N_15143,N_14649,N_14901);
and U15144 (N_15144,N_14703,N_14695);
or U15145 (N_15145,N_14752,N_14893);
or U15146 (N_15146,N_14968,N_14958);
nand U15147 (N_15147,N_14724,N_14600);
and U15148 (N_15148,N_14671,N_14688);
or U15149 (N_15149,N_14804,N_14575);
xnor U15150 (N_15150,N_14737,N_14678);
and U15151 (N_15151,N_14998,N_14959);
xnor U15152 (N_15152,N_14940,N_14788);
nand U15153 (N_15153,N_14873,N_14574);
nand U15154 (N_15154,N_14599,N_14662);
xor U15155 (N_15155,N_14797,N_14880);
xnor U15156 (N_15156,N_14945,N_14500);
or U15157 (N_15157,N_14868,N_14592);
nor U15158 (N_15158,N_14764,N_14957);
xor U15159 (N_15159,N_14856,N_14889);
or U15160 (N_15160,N_14661,N_14853);
and U15161 (N_15161,N_14877,N_14686);
nor U15162 (N_15162,N_14780,N_14769);
and U15163 (N_15163,N_14503,N_14634);
nor U15164 (N_15164,N_14645,N_14828);
nor U15165 (N_15165,N_14815,N_14545);
nor U15166 (N_15166,N_14834,N_14983);
and U15167 (N_15167,N_14991,N_14825);
nand U15168 (N_15168,N_14812,N_14999);
or U15169 (N_15169,N_14502,N_14768);
and U15170 (N_15170,N_14840,N_14690);
and U15171 (N_15171,N_14808,N_14895);
xnor U15172 (N_15172,N_14835,N_14591);
xnor U15173 (N_15173,N_14636,N_14849);
xor U15174 (N_15174,N_14564,N_14777);
or U15175 (N_15175,N_14642,N_14509);
nand U15176 (N_15176,N_14965,N_14734);
or U15177 (N_15177,N_14530,N_14833);
xor U15178 (N_15178,N_14864,N_14771);
or U15179 (N_15179,N_14710,N_14884);
nand U15180 (N_15180,N_14519,N_14680);
nand U15181 (N_15181,N_14750,N_14756);
or U15182 (N_15182,N_14782,N_14839);
or U15183 (N_15183,N_14843,N_14967);
or U15184 (N_15184,N_14644,N_14776);
nor U15185 (N_15185,N_14966,N_14578);
or U15186 (N_15186,N_14544,N_14954);
and U15187 (N_15187,N_14510,N_14647);
or U15188 (N_15188,N_14572,N_14653);
and U15189 (N_15189,N_14563,N_14818);
or U15190 (N_15190,N_14547,N_14692);
nand U15191 (N_15191,N_14819,N_14929);
nand U15192 (N_15192,N_14702,N_14566);
xor U15193 (N_15193,N_14620,N_14637);
or U15194 (N_15194,N_14713,N_14718);
nor U15195 (N_15195,N_14643,N_14876);
and U15196 (N_15196,N_14949,N_14855);
xor U15197 (N_15197,N_14619,N_14551);
xor U15198 (N_15198,N_14951,N_14754);
xor U15199 (N_15199,N_14751,N_14652);
and U15200 (N_15200,N_14505,N_14656);
and U15201 (N_15201,N_14715,N_14786);
or U15202 (N_15202,N_14885,N_14846);
nand U15203 (N_15203,N_14982,N_14831);
or U15204 (N_15204,N_14822,N_14793);
nand U15205 (N_15205,N_14538,N_14615);
nor U15206 (N_15206,N_14874,N_14763);
or U15207 (N_15207,N_14836,N_14666);
or U15208 (N_15208,N_14979,N_14598);
xor U15209 (N_15209,N_14504,N_14934);
and U15210 (N_15210,N_14964,N_14646);
nor U15211 (N_15211,N_14531,N_14915);
or U15212 (N_15212,N_14632,N_14902);
and U15213 (N_15213,N_14821,N_14928);
xor U15214 (N_15214,N_14990,N_14820);
xnor U15215 (N_15215,N_14675,N_14587);
nor U15216 (N_15216,N_14760,N_14593);
and U15217 (N_15217,N_14872,N_14762);
or U15218 (N_15218,N_14753,N_14720);
nand U15219 (N_15219,N_14559,N_14860);
or U15220 (N_15220,N_14947,N_14558);
nand U15221 (N_15221,N_14783,N_14930);
or U15222 (N_15222,N_14844,N_14569);
xnor U15223 (N_15223,N_14773,N_14555);
or U15224 (N_15224,N_14682,N_14562);
nor U15225 (N_15225,N_14691,N_14925);
xor U15226 (N_15226,N_14863,N_14996);
xnor U15227 (N_15227,N_14890,N_14697);
nand U15228 (N_15228,N_14626,N_14781);
or U15229 (N_15229,N_14987,N_14778);
xor U15230 (N_15230,N_14595,N_14685);
and U15231 (N_15231,N_14847,N_14805);
nand U15232 (N_15232,N_14920,N_14993);
and U15233 (N_15233,N_14898,N_14899);
and U15234 (N_15234,N_14512,N_14613);
nor U15235 (N_15235,N_14520,N_14570);
and U15236 (N_15236,N_14800,N_14870);
nand U15237 (N_15237,N_14583,N_14584);
or U15238 (N_15238,N_14669,N_14796);
and U15239 (N_15239,N_14878,N_14540);
xnor U15240 (N_15240,N_14963,N_14910);
nand U15241 (N_15241,N_14625,N_14907);
xor U15242 (N_15242,N_14571,N_14638);
or U15243 (N_15243,N_14742,N_14917);
xnor U15244 (N_15244,N_14897,N_14755);
or U15245 (N_15245,N_14944,N_14581);
and U15246 (N_15246,N_14722,N_14851);
xor U15247 (N_15247,N_14830,N_14533);
nand U15248 (N_15248,N_14740,N_14792);
nor U15249 (N_15249,N_14986,N_14731);
and U15250 (N_15250,N_14811,N_14546);
nor U15251 (N_15251,N_14844,N_14706);
and U15252 (N_15252,N_14613,N_14807);
nor U15253 (N_15253,N_14735,N_14838);
and U15254 (N_15254,N_14720,N_14692);
nand U15255 (N_15255,N_14677,N_14924);
or U15256 (N_15256,N_14799,N_14632);
nor U15257 (N_15257,N_14829,N_14706);
and U15258 (N_15258,N_14969,N_14753);
nand U15259 (N_15259,N_14987,N_14802);
and U15260 (N_15260,N_14733,N_14757);
and U15261 (N_15261,N_14941,N_14532);
nand U15262 (N_15262,N_14807,N_14589);
nor U15263 (N_15263,N_14886,N_14661);
nor U15264 (N_15264,N_14880,N_14513);
xor U15265 (N_15265,N_14875,N_14698);
and U15266 (N_15266,N_14632,N_14937);
xnor U15267 (N_15267,N_14881,N_14532);
or U15268 (N_15268,N_14755,N_14740);
nor U15269 (N_15269,N_14830,N_14761);
xor U15270 (N_15270,N_14841,N_14904);
and U15271 (N_15271,N_14526,N_14838);
and U15272 (N_15272,N_14864,N_14706);
or U15273 (N_15273,N_14655,N_14904);
or U15274 (N_15274,N_14816,N_14824);
nand U15275 (N_15275,N_14516,N_14613);
nor U15276 (N_15276,N_14974,N_14653);
and U15277 (N_15277,N_14602,N_14925);
or U15278 (N_15278,N_14870,N_14914);
nand U15279 (N_15279,N_14903,N_14732);
nand U15280 (N_15280,N_14869,N_14651);
nand U15281 (N_15281,N_14950,N_14571);
nand U15282 (N_15282,N_14807,N_14741);
nand U15283 (N_15283,N_14746,N_14705);
xnor U15284 (N_15284,N_14677,N_14590);
nor U15285 (N_15285,N_14678,N_14536);
xor U15286 (N_15286,N_14758,N_14613);
nand U15287 (N_15287,N_14587,N_14738);
or U15288 (N_15288,N_14511,N_14813);
nor U15289 (N_15289,N_14664,N_14849);
xor U15290 (N_15290,N_14756,N_14916);
nand U15291 (N_15291,N_14566,N_14627);
nand U15292 (N_15292,N_14592,N_14700);
or U15293 (N_15293,N_14742,N_14861);
xnor U15294 (N_15294,N_14750,N_14837);
or U15295 (N_15295,N_14597,N_14842);
xor U15296 (N_15296,N_14812,N_14903);
nor U15297 (N_15297,N_14995,N_14953);
xor U15298 (N_15298,N_14970,N_14642);
nor U15299 (N_15299,N_14701,N_14583);
or U15300 (N_15300,N_14755,N_14843);
xor U15301 (N_15301,N_14919,N_14548);
or U15302 (N_15302,N_14553,N_14615);
nor U15303 (N_15303,N_14959,N_14662);
nor U15304 (N_15304,N_14624,N_14610);
or U15305 (N_15305,N_14928,N_14843);
xor U15306 (N_15306,N_14548,N_14658);
or U15307 (N_15307,N_14611,N_14626);
or U15308 (N_15308,N_14911,N_14921);
nor U15309 (N_15309,N_14941,N_14533);
xor U15310 (N_15310,N_14856,N_14716);
nand U15311 (N_15311,N_14771,N_14986);
and U15312 (N_15312,N_14639,N_14982);
nand U15313 (N_15313,N_14705,N_14621);
nor U15314 (N_15314,N_14925,N_14965);
xnor U15315 (N_15315,N_14580,N_14820);
or U15316 (N_15316,N_14637,N_14573);
nand U15317 (N_15317,N_14876,N_14502);
nor U15318 (N_15318,N_14878,N_14775);
xor U15319 (N_15319,N_14742,N_14758);
and U15320 (N_15320,N_14858,N_14844);
or U15321 (N_15321,N_14729,N_14580);
and U15322 (N_15322,N_14633,N_14955);
xnor U15323 (N_15323,N_14840,N_14925);
xnor U15324 (N_15324,N_14582,N_14757);
or U15325 (N_15325,N_14889,N_14567);
nand U15326 (N_15326,N_14579,N_14854);
nand U15327 (N_15327,N_14811,N_14577);
or U15328 (N_15328,N_14898,N_14689);
nand U15329 (N_15329,N_14640,N_14908);
nor U15330 (N_15330,N_14665,N_14991);
or U15331 (N_15331,N_14764,N_14834);
xor U15332 (N_15332,N_14560,N_14866);
nand U15333 (N_15333,N_14555,N_14828);
or U15334 (N_15334,N_14783,N_14763);
xor U15335 (N_15335,N_14673,N_14685);
nand U15336 (N_15336,N_14581,N_14868);
nor U15337 (N_15337,N_14798,N_14625);
and U15338 (N_15338,N_14816,N_14768);
or U15339 (N_15339,N_14787,N_14545);
and U15340 (N_15340,N_14511,N_14795);
xnor U15341 (N_15341,N_14827,N_14870);
and U15342 (N_15342,N_14977,N_14594);
nor U15343 (N_15343,N_14945,N_14561);
nand U15344 (N_15344,N_14939,N_14531);
xnor U15345 (N_15345,N_14792,N_14958);
xnor U15346 (N_15346,N_14533,N_14719);
or U15347 (N_15347,N_14670,N_14855);
xnor U15348 (N_15348,N_14809,N_14926);
and U15349 (N_15349,N_14674,N_14596);
and U15350 (N_15350,N_14834,N_14618);
nor U15351 (N_15351,N_14501,N_14939);
nand U15352 (N_15352,N_14516,N_14897);
nor U15353 (N_15353,N_14921,N_14558);
nand U15354 (N_15354,N_14934,N_14580);
or U15355 (N_15355,N_14887,N_14985);
nor U15356 (N_15356,N_14548,N_14645);
or U15357 (N_15357,N_14607,N_14733);
xor U15358 (N_15358,N_14532,N_14929);
nor U15359 (N_15359,N_14528,N_14903);
nand U15360 (N_15360,N_14566,N_14902);
and U15361 (N_15361,N_14619,N_14889);
nand U15362 (N_15362,N_14924,N_14583);
nor U15363 (N_15363,N_14590,N_14574);
nand U15364 (N_15364,N_14502,N_14748);
and U15365 (N_15365,N_14575,N_14981);
nand U15366 (N_15366,N_14591,N_14882);
xnor U15367 (N_15367,N_14984,N_14961);
or U15368 (N_15368,N_14560,N_14789);
and U15369 (N_15369,N_14734,N_14698);
nand U15370 (N_15370,N_14622,N_14956);
nand U15371 (N_15371,N_14957,N_14537);
or U15372 (N_15372,N_14766,N_14634);
or U15373 (N_15373,N_14839,N_14985);
and U15374 (N_15374,N_14715,N_14760);
and U15375 (N_15375,N_14734,N_14966);
nor U15376 (N_15376,N_14531,N_14760);
xor U15377 (N_15377,N_14846,N_14811);
and U15378 (N_15378,N_14560,N_14510);
or U15379 (N_15379,N_14938,N_14925);
nor U15380 (N_15380,N_14501,N_14680);
xnor U15381 (N_15381,N_14519,N_14708);
or U15382 (N_15382,N_14922,N_14557);
nand U15383 (N_15383,N_14542,N_14849);
nand U15384 (N_15384,N_14676,N_14904);
nand U15385 (N_15385,N_14642,N_14811);
xnor U15386 (N_15386,N_14674,N_14642);
or U15387 (N_15387,N_14846,N_14629);
nand U15388 (N_15388,N_14787,N_14804);
nand U15389 (N_15389,N_14615,N_14832);
and U15390 (N_15390,N_14571,N_14628);
nand U15391 (N_15391,N_14719,N_14657);
xor U15392 (N_15392,N_14501,N_14653);
nand U15393 (N_15393,N_14668,N_14822);
or U15394 (N_15394,N_14991,N_14909);
nor U15395 (N_15395,N_14825,N_14530);
nand U15396 (N_15396,N_14925,N_14974);
nor U15397 (N_15397,N_14909,N_14518);
nor U15398 (N_15398,N_14867,N_14778);
or U15399 (N_15399,N_14815,N_14680);
nor U15400 (N_15400,N_14908,N_14861);
or U15401 (N_15401,N_14876,N_14577);
nand U15402 (N_15402,N_14890,N_14918);
or U15403 (N_15403,N_14676,N_14914);
or U15404 (N_15404,N_14685,N_14703);
or U15405 (N_15405,N_14967,N_14820);
nor U15406 (N_15406,N_14740,N_14534);
xnor U15407 (N_15407,N_14612,N_14915);
xor U15408 (N_15408,N_14836,N_14669);
or U15409 (N_15409,N_14772,N_14588);
nor U15410 (N_15410,N_14849,N_14659);
or U15411 (N_15411,N_14749,N_14620);
xor U15412 (N_15412,N_14796,N_14981);
nand U15413 (N_15413,N_14596,N_14625);
xor U15414 (N_15414,N_14939,N_14766);
nand U15415 (N_15415,N_14533,N_14997);
or U15416 (N_15416,N_14986,N_14881);
xnor U15417 (N_15417,N_14545,N_14821);
and U15418 (N_15418,N_14850,N_14969);
nor U15419 (N_15419,N_14522,N_14978);
and U15420 (N_15420,N_14949,N_14764);
or U15421 (N_15421,N_14828,N_14992);
xnor U15422 (N_15422,N_14609,N_14758);
nand U15423 (N_15423,N_14556,N_14654);
nand U15424 (N_15424,N_14744,N_14860);
or U15425 (N_15425,N_14770,N_14728);
or U15426 (N_15426,N_14649,N_14928);
and U15427 (N_15427,N_14995,N_14568);
xor U15428 (N_15428,N_14999,N_14909);
and U15429 (N_15429,N_14885,N_14851);
nand U15430 (N_15430,N_14700,N_14781);
xnor U15431 (N_15431,N_14518,N_14699);
xnor U15432 (N_15432,N_14801,N_14872);
and U15433 (N_15433,N_14685,N_14770);
xnor U15434 (N_15434,N_14740,N_14832);
or U15435 (N_15435,N_14786,N_14881);
xnor U15436 (N_15436,N_14764,N_14758);
nand U15437 (N_15437,N_14806,N_14670);
xnor U15438 (N_15438,N_14990,N_14824);
or U15439 (N_15439,N_14924,N_14884);
or U15440 (N_15440,N_14948,N_14737);
nor U15441 (N_15441,N_14867,N_14507);
nand U15442 (N_15442,N_14816,N_14851);
and U15443 (N_15443,N_14964,N_14801);
nand U15444 (N_15444,N_14532,N_14671);
nor U15445 (N_15445,N_14628,N_14738);
or U15446 (N_15446,N_14591,N_14842);
nor U15447 (N_15447,N_14934,N_14961);
nor U15448 (N_15448,N_14537,N_14642);
nor U15449 (N_15449,N_14501,N_14729);
nor U15450 (N_15450,N_14849,N_14719);
nand U15451 (N_15451,N_14578,N_14632);
xor U15452 (N_15452,N_14829,N_14744);
or U15453 (N_15453,N_14556,N_14530);
nor U15454 (N_15454,N_14951,N_14822);
or U15455 (N_15455,N_14879,N_14739);
xor U15456 (N_15456,N_14797,N_14865);
nand U15457 (N_15457,N_14891,N_14810);
xnor U15458 (N_15458,N_14744,N_14617);
xnor U15459 (N_15459,N_14802,N_14999);
nand U15460 (N_15460,N_14643,N_14652);
or U15461 (N_15461,N_14848,N_14723);
xor U15462 (N_15462,N_14642,N_14666);
xor U15463 (N_15463,N_14895,N_14985);
xnor U15464 (N_15464,N_14530,N_14505);
nand U15465 (N_15465,N_14583,N_14982);
xor U15466 (N_15466,N_14535,N_14855);
or U15467 (N_15467,N_14643,N_14731);
xnor U15468 (N_15468,N_14851,N_14877);
xnor U15469 (N_15469,N_14993,N_14841);
nor U15470 (N_15470,N_14547,N_14693);
and U15471 (N_15471,N_14967,N_14881);
and U15472 (N_15472,N_14858,N_14695);
nor U15473 (N_15473,N_14865,N_14892);
nand U15474 (N_15474,N_14853,N_14829);
or U15475 (N_15475,N_14942,N_14908);
nand U15476 (N_15476,N_14714,N_14609);
xor U15477 (N_15477,N_14882,N_14814);
and U15478 (N_15478,N_14711,N_14559);
nand U15479 (N_15479,N_14718,N_14649);
and U15480 (N_15480,N_14694,N_14622);
and U15481 (N_15481,N_14634,N_14902);
nor U15482 (N_15482,N_14595,N_14720);
nand U15483 (N_15483,N_14636,N_14956);
and U15484 (N_15484,N_14981,N_14553);
nand U15485 (N_15485,N_14805,N_14658);
and U15486 (N_15486,N_14910,N_14926);
or U15487 (N_15487,N_14683,N_14615);
xor U15488 (N_15488,N_14970,N_14660);
nor U15489 (N_15489,N_14603,N_14684);
nor U15490 (N_15490,N_14645,N_14975);
and U15491 (N_15491,N_14865,N_14742);
nand U15492 (N_15492,N_14714,N_14820);
nor U15493 (N_15493,N_14678,N_14685);
nor U15494 (N_15494,N_14950,N_14638);
nor U15495 (N_15495,N_14598,N_14778);
xor U15496 (N_15496,N_14933,N_14944);
nand U15497 (N_15497,N_14828,N_14532);
nor U15498 (N_15498,N_14572,N_14595);
and U15499 (N_15499,N_14664,N_14544);
nor U15500 (N_15500,N_15300,N_15048);
nand U15501 (N_15501,N_15331,N_15071);
or U15502 (N_15502,N_15204,N_15181);
and U15503 (N_15503,N_15091,N_15141);
nor U15504 (N_15504,N_15168,N_15039);
and U15505 (N_15505,N_15394,N_15382);
nand U15506 (N_15506,N_15279,N_15421);
nor U15507 (N_15507,N_15208,N_15156);
and U15508 (N_15508,N_15325,N_15232);
nor U15509 (N_15509,N_15079,N_15165);
nand U15510 (N_15510,N_15121,N_15342);
nor U15511 (N_15511,N_15040,N_15195);
nand U15512 (N_15512,N_15174,N_15410);
and U15513 (N_15513,N_15041,N_15182);
nor U15514 (N_15514,N_15096,N_15332);
nor U15515 (N_15515,N_15015,N_15225);
nand U15516 (N_15516,N_15160,N_15109);
and U15517 (N_15517,N_15294,N_15367);
or U15518 (N_15518,N_15173,N_15350);
xnor U15519 (N_15519,N_15044,N_15050);
nand U15520 (N_15520,N_15283,N_15073);
nand U15521 (N_15521,N_15319,N_15357);
xor U15522 (N_15522,N_15134,N_15488);
nor U15523 (N_15523,N_15406,N_15102);
and U15524 (N_15524,N_15428,N_15179);
xnor U15525 (N_15525,N_15224,N_15155);
xor U15526 (N_15526,N_15199,N_15218);
or U15527 (N_15527,N_15494,N_15444);
nand U15528 (N_15528,N_15497,N_15143);
or U15529 (N_15529,N_15403,N_15392);
or U15530 (N_15530,N_15068,N_15329);
or U15531 (N_15531,N_15347,N_15483);
xnor U15532 (N_15532,N_15315,N_15476);
nor U15533 (N_15533,N_15405,N_15256);
xor U15534 (N_15534,N_15021,N_15250);
xor U15535 (N_15535,N_15498,N_15390);
xor U15536 (N_15536,N_15280,N_15380);
nor U15537 (N_15537,N_15378,N_15239);
nor U15538 (N_15538,N_15043,N_15164);
or U15539 (N_15539,N_15138,N_15070);
nor U15540 (N_15540,N_15275,N_15062);
xnor U15541 (N_15541,N_15177,N_15284);
xnor U15542 (N_15542,N_15020,N_15397);
or U15543 (N_15543,N_15217,N_15274);
xnor U15544 (N_15544,N_15118,N_15482);
or U15545 (N_15545,N_15242,N_15408);
and U15546 (N_15546,N_15167,N_15411);
nand U15547 (N_15547,N_15265,N_15277);
and U15548 (N_15548,N_15231,N_15078);
xor U15549 (N_15549,N_15148,N_15478);
or U15550 (N_15550,N_15477,N_15158);
nand U15551 (N_15551,N_15320,N_15180);
nand U15552 (N_15552,N_15067,N_15309);
xnor U15553 (N_15553,N_15082,N_15339);
nand U15554 (N_15554,N_15462,N_15424);
and U15555 (N_15555,N_15171,N_15415);
xor U15556 (N_15556,N_15293,N_15370);
and U15557 (N_15557,N_15024,N_15456);
nor U15558 (N_15558,N_15058,N_15324);
nor U15559 (N_15559,N_15057,N_15150);
nand U15560 (N_15560,N_15356,N_15417);
and U15561 (N_15561,N_15384,N_15372);
nor U15562 (N_15562,N_15166,N_15090);
and U15563 (N_15563,N_15425,N_15402);
or U15564 (N_15564,N_15423,N_15323);
and U15565 (N_15565,N_15053,N_15375);
nor U15566 (N_15566,N_15414,N_15278);
nand U15567 (N_15567,N_15445,N_15122);
xor U15568 (N_15568,N_15396,N_15254);
or U15569 (N_15569,N_15258,N_15426);
and U15570 (N_15570,N_15340,N_15151);
xnor U15571 (N_15571,N_15216,N_15175);
nor U15572 (N_15572,N_15318,N_15213);
nand U15573 (N_15573,N_15328,N_15139);
or U15574 (N_15574,N_15471,N_15271);
or U15575 (N_15575,N_15412,N_15066);
or U15576 (N_15576,N_15076,N_15446);
nand U15577 (N_15577,N_15114,N_15314);
or U15578 (N_15578,N_15334,N_15341);
xnor U15579 (N_15579,N_15391,N_15023);
nor U15580 (N_15580,N_15363,N_15313);
nand U15581 (N_15581,N_15119,N_15100);
and U15582 (N_15582,N_15248,N_15144);
or U15583 (N_15583,N_15310,N_15107);
and U15584 (N_15584,N_15029,N_15115);
and U15585 (N_15585,N_15321,N_15436);
nand U15586 (N_15586,N_15223,N_15205);
or U15587 (N_15587,N_15172,N_15192);
nand U15588 (N_15588,N_15170,N_15188);
nor U15589 (N_15589,N_15452,N_15000);
or U15590 (N_15590,N_15008,N_15465);
nand U15591 (N_15591,N_15002,N_15296);
and U15592 (N_15592,N_15336,N_15433);
xnor U15593 (N_15593,N_15450,N_15330);
xor U15594 (N_15594,N_15492,N_15381);
nand U15595 (N_15595,N_15466,N_15418);
nor U15596 (N_15596,N_15472,N_15260);
nand U15597 (N_15597,N_15147,N_15491);
nand U15598 (N_15598,N_15128,N_15055);
nor U15599 (N_15599,N_15369,N_15261);
or U15600 (N_15600,N_15352,N_15443);
or U15601 (N_15601,N_15276,N_15273);
nor U15602 (N_15602,N_15022,N_15012);
nand U15603 (N_15603,N_15312,N_15110);
xnor U15604 (N_15604,N_15094,N_15063);
xnor U15605 (N_15605,N_15010,N_15441);
or U15606 (N_15606,N_15270,N_15133);
xnor U15607 (N_15607,N_15186,N_15049);
nand U15608 (N_15608,N_15458,N_15159);
or U15609 (N_15609,N_15437,N_15474);
nand U15610 (N_15610,N_15243,N_15292);
nor U15611 (N_15611,N_15487,N_15489);
and U15612 (N_15612,N_15153,N_15108);
nor U15613 (N_15613,N_15095,N_15101);
nor U15614 (N_15614,N_15374,N_15286);
and U15615 (N_15615,N_15289,N_15311);
nand U15616 (N_15616,N_15282,N_15061);
or U15617 (N_15617,N_15221,N_15305);
nor U15618 (N_15618,N_15210,N_15016);
or U15619 (N_15619,N_15035,N_15442);
or U15620 (N_15620,N_15364,N_15197);
and U15621 (N_15621,N_15353,N_15187);
nor U15622 (N_15622,N_15077,N_15361);
nor U15623 (N_15623,N_15299,N_15255);
xor U15624 (N_15624,N_15327,N_15463);
nand U15625 (N_15625,N_15263,N_15371);
or U15626 (N_15626,N_15127,N_15257);
nand U15627 (N_15627,N_15304,N_15354);
nand U15628 (N_15628,N_15413,N_15338);
nor U15629 (N_15629,N_15129,N_15237);
or U15630 (N_15630,N_15163,N_15196);
xor U15631 (N_15631,N_15026,N_15429);
xnor U15632 (N_15632,N_15475,N_15081);
nand U15633 (N_15633,N_15287,N_15084);
nand U15634 (N_15634,N_15348,N_15295);
or U15635 (N_15635,N_15496,N_15430);
nor U15636 (N_15636,N_15075,N_15365);
and U15637 (N_15637,N_15395,N_15266);
xor U15638 (N_15638,N_15461,N_15161);
nand U15639 (N_15639,N_15473,N_15269);
xor U15640 (N_15640,N_15033,N_15203);
nand U15641 (N_15641,N_15307,N_15220);
nand U15642 (N_15642,N_15056,N_15290);
or U15643 (N_15643,N_15301,N_15051);
or U15644 (N_15644,N_15302,N_15099);
and U15645 (N_15645,N_15235,N_15316);
or U15646 (N_15646,N_15025,N_15240);
nand U15647 (N_15647,N_15132,N_15422);
or U15648 (N_15648,N_15125,N_15288);
xor U15649 (N_15649,N_15136,N_15401);
xor U15650 (N_15650,N_15103,N_15470);
xnor U15651 (N_15651,N_15386,N_15383);
nand U15652 (N_15652,N_15014,N_15137);
or U15653 (N_15653,N_15226,N_15400);
nand U15654 (N_15654,N_15135,N_15211);
nand U15655 (N_15655,N_15459,N_15416);
nand U15656 (N_15656,N_15233,N_15467);
and U15657 (N_15657,N_15080,N_15484);
nand U15658 (N_15658,N_15335,N_15183);
or U15659 (N_15659,N_15398,N_15004);
nor U15660 (N_15660,N_15435,N_15030);
nand U15661 (N_15661,N_15317,N_15162);
xor U15662 (N_15662,N_15018,N_15252);
nor U15663 (N_15663,N_15454,N_15176);
or U15664 (N_15664,N_15326,N_15126);
and U15665 (N_15665,N_15149,N_15045);
and U15666 (N_15666,N_15031,N_15069);
and U15667 (N_15667,N_15448,N_15447);
nor U15668 (N_15668,N_15373,N_15086);
nand U15669 (N_15669,N_15479,N_15007);
xnor U15670 (N_15670,N_15368,N_15038);
and U15671 (N_15671,N_15111,N_15229);
nand U15672 (N_15672,N_15457,N_15189);
or U15673 (N_15673,N_15106,N_15333);
and U15674 (N_15674,N_15419,N_15194);
nor U15675 (N_15675,N_15431,N_15389);
and U15676 (N_15676,N_15366,N_15200);
nor U15677 (N_15677,N_15469,N_15493);
xor U15678 (N_15678,N_15253,N_15009);
xnor U15679 (N_15679,N_15427,N_15268);
and U15680 (N_15680,N_15184,N_15191);
and U15681 (N_15681,N_15360,N_15404);
nand U15682 (N_15682,N_15207,N_15298);
xor U15683 (N_15683,N_15098,N_15434);
and U15684 (N_15684,N_15351,N_15169);
nor U15685 (N_15685,N_15495,N_15297);
or U15686 (N_15686,N_15306,N_15214);
or U15687 (N_15687,N_15190,N_15215);
nand U15688 (N_15688,N_15006,N_15085);
nor U15689 (N_15689,N_15142,N_15227);
xor U15690 (N_15690,N_15027,N_15453);
or U15691 (N_15691,N_15272,N_15193);
and U15692 (N_15692,N_15499,N_15245);
nor U15693 (N_15693,N_15054,N_15005);
xor U15694 (N_15694,N_15480,N_15490);
nor U15695 (N_15695,N_15449,N_15262);
nor U15696 (N_15696,N_15346,N_15322);
nor U15697 (N_15697,N_15120,N_15198);
nor U15698 (N_15698,N_15097,N_15281);
and U15699 (N_15699,N_15124,N_15238);
nor U15700 (N_15700,N_15247,N_15451);
nor U15701 (N_15701,N_15407,N_15152);
xnor U15702 (N_15702,N_15432,N_15013);
and U15703 (N_15703,N_15481,N_15251);
or U15704 (N_15704,N_15130,N_15157);
nor U15705 (N_15705,N_15345,N_15093);
and U15706 (N_15706,N_15105,N_15065);
and U15707 (N_15707,N_15145,N_15178);
or U15708 (N_15708,N_15264,N_15379);
or U15709 (N_15709,N_15438,N_15037);
xor U15710 (N_15710,N_15249,N_15117);
or U15711 (N_15711,N_15267,N_15439);
and U15712 (N_15712,N_15291,N_15042);
and U15713 (N_15713,N_15359,N_15337);
nor U15714 (N_15714,N_15034,N_15385);
nand U15715 (N_15715,N_15185,N_15440);
nand U15716 (N_15716,N_15486,N_15485);
or U15717 (N_15717,N_15028,N_15092);
nand U15718 (N_15718,N_15420,N_15001);
and U15719 (N_15719,N_15064,N_15123);
or U15720 (N_15720,N_15244,N_15344);
nor U15721 (N_15721,N_15003,N_15259);
and U15722 (N_15722,N_15388,N_15399);
or U15723 (N_15723,N_15377,N_15140);
xnor U15724 (N_15724,N_15241,N_15468);
and U15725 (N_15725,N_15032,N_15230);
or U15726 (N_15726,N_15036,N_15464);
nand U15727 (N_15727,N_15131,N_15052);
nor U15728 (N_15728,N_15046,N_15376);
and U15729 (N_15729,N_15074,N_15455);
nor U15730 (N_15730,N_15246,N_15212);
xor U15731 (N_15731,N_15355,N_15219);
nor U15732 (N_15732,N_15222,N_15011);
or U15733 (N_15733,N_15236,N_15393);
xor U15734 (N_15734,N_15059,N_15209);
nand U15735 (N_15735,N_15308,N_15234);
or U15736 (N_15736,N_15017,N_15113);
nor U15737 (N_15737,N_15460,N_15362);
nand U15738 (N_15738,N_15087,N_15206);
xnor U15739 (N_15739,N_15116,N_15088);
xor U15740 (N_15740,N_15112,N_15358);
xnor U15741 (N_15741,N_15343,N_15202);
nand U15742 (N_15742,N_15047,N_15089);
or U15743 (N_15743,N_15285,N_15154);
and U15744 (N_15744,N_15303,N_15146);
nor U15745 (N_15745,N_15228,N_15201);
nor U15746 (N_15746,N_15072,N_15387);
nor U15747 (N_15747,N_15019,N_15104);
xor U15748 (N_15748,N_15083,N_15060);
xor U15749 (N_15749,N_15349,N_15409);
or U15750 (N_15750,N_15474,N_15401);
nor U15751 (N_15751,N_15402,N_15404);
nor U15752 (N_15752,N_15412,N_15135);
nor U15753 (N_15753,N_15174,N_15079);
nand U15754 (N_15754,N_15063,N_15162);
nand U15755 (N_15755,N_15197,N_15106);
nand U15756 (N_15756,N_15442,N_15096);
and U15757 (N_15757,N_15360,N_15295);
nor U15758 (N_15758,N_15235,N_15399);
or U15759 (N_15759,N_15406,N_15369);
nand U15760 (N_15760,N_15102,N_15329);
and U15761 (N_15761,N_15417,N_15199);
nor U15762 (N_15762,N_15251,N_15055);
nor U15763 (N_15763,N_15082,N_15030);
nand U15764 (N_15764,N_15271,N_15101);
or U15765 (N_15765,N_15258,N_15378);
xnor U15766 (N_15766,N_15255,N_15332);
nand U15767 (N_15767,N_15376,N_15084);
nor U15768 (N_15768,N_15312,N_15126);
nand U15769 (N_15769,N_15389,N_15135);
and U15770 (N_15770,N_15419,N_15355);
nor U15771 (N_15771,N_15446,N_15180);
and U15772 (N_15772,N_15194,N_15246);
nand U15773 (N_15773,N_15175,N_15429);
nor U15774 (N_15774,N_15091,N_15144);
nand U15775 (N_15775,N_15106,N_15023);
and U15776 (N_15776,N_15283,N_15368);
xnor U15777 (N_15777,N_15349,N_15463);
nor U15778 (N_15778,N_15115,N_15007);
nor U15779 (N_15779,N_15138,N_15249);
or U15780 (N_15780,N_15314,N_15162);
xor U15781 (N_15781,N_15244,N_15037);
nand U15782 (N_15782,N_15359,N_15001);
and U15783 (N_15783,N_15412,N_15464);
nor U15784 (N_15784,N_15393,N_15213);
nand U15785 (N_15785,N_15079,N_15447);
nand U15786 (N_15786,N_15465,N_15437);
or U15787 (N_15787,N_15269,N_15228);
or U15788 (N_15788,N_15194,N_15156);
and U15789 (N_15789,N_15335,N_15316);
and U15790 (N_15790,N_15179,N_15334);
and U15791 (N_15791,N_15173,N_15052);
nor U15792 (N_15792,N_15298,N_15339);
or U15793 (N_15793,N_15473,N_15325);
nor U15794 (N_15794,N_15298,N_15497);
xnor U15795 (N_15795,N_15222,N_15432);
xor U15796 (N_15796,N_15482,N_15027);
or U15797 (N_15797,N_15264,N_15173);
and U15798 (N_15798,N_15419,N_15372);
nor U15799 (N_15799,N_15471,N_15280);
and U15800 (N_15800,N_15112,N_15479);
nor U15801 (N_15801,N_15015,N_15132);
or U15802 (N_15802,N_15169,N_15153);
and U15803 (N_15803,N_15439,N_15441);
xnor U15804 (N_15804,N_15087,N_15413);
nor U15805 (N_15805,N_15195,N_15192);
nand U15806 (N_15806,N_15364,N_15315);
nor U15807 (N_15807,N_15140,N_15130);
or U15808 (N_15808,N_15200,N_15348);
or U15809 (N_15809,N_15404,N_15262);
nor U15810 (N_15810,N_15289,N_15216);
nor U15811 (N_15811,N_15426,N_15279);
nand U15812 (N_15812,N_15033,N_15078);
or U15813 (N_15813,N_15294,N_15378);
xnor U15814 (N_15814,N_15264,N_15309);
or U15815 (N_15815,N_15237,N_15219);
xor U15816 (N_15816,N_15147,N_15337);
xnor U15817 (N_15817,N_15275,N_15372);
nor U15818 (N_15818,N_15236,N_15418);
and U15819 (N_15819,N_15272,N_15265);
or U15820 (N_15820,N_15069,N_15327);
xnor U15821 (N_15821,N_15085,N_15181);
xor U15822 (N_15822,N_15454,N_15416);
or U15823 (N_15823,N_15169,N_15154);
nor U15824 (N_15824,N_15124,N_15367);
nand U15825 (N_15825,N_15095,N_15073);
and U15826 (N_15826,N_15493,N_15342);
nand U15827 (N_15827,N_15031,N_15315);
nand U15828 (N_15828,N_15175,N_15081);
or U15829 (N_15829,N_15129,N_15053);
or U15830 (N_15830,N_15092,N_15013);
nor U15831 (N_15831,N_15376,N_15005);
nor U15832 (N_15832,N_15441,N_15046);
and U15833 (N_15833,N_15322,N_15366);
or U15834 (N_15834,N_15464,N_15163);
and U15835 (N_15835,N_15462,N_15161);
nor U15836 (N_15836,N_15137,N_15022);
and U15837 (N_15837,N_15106,N_15107);
nor U15838 (N_15838,N_15008,N_15341);
xor U15839 (N_15839,N_15056,N_15139);
nand U15840 (N_15840,N_15410,N_15070);
nor U15841 (N_15841,N_15455,N_15464);
or U15842 (N_15842,N_15194,N_15055);
nand U15843 (N_15843,N_15046,N_15108);
and U15844 (N_15844,N_15346,N_15380);
or U15845 (N_15845,N_15181,N_15413);
xnor U15846 (N_15846,N_15428,N_15267);
nor U15847 (N_15847,N_15290,N_15233);
xnor U15848 (N_15848,N_15407,N_15473);
and U15849 (N_15849,N_15298,N_15099);
or U15850 (N_15850,N_15090,N_15199);
and U15851 (N_15851,N_15364,N_15493);
nand U15852 (N_15852,N_15446,N_15424);
nor U15853 (N_15853,N_15441,N_15321);
nand U15854 (N_15854,N_15040,N_15208);
nand U15855 (N_15855,N_15428,N_15349);
xnor U15856 (N_15856,N_15294,N_15406);
and U15857 (N_15857,N_15239,N_15098);
and U15858 (N_15858,N_15303,N_15188);
xor U15859 (N_15859,N_15495,N_15333);
nand U15860 (N_15860,N_15388,N_15305);
nor U15861 (N_15861,N_15375,N_15333);
xor U15862 (N_15862,N_15290,N_15405);
xor U15863 (N_15863,N_15294,N_15025);
or U15864 (N_15864,N_15034,N_15117);
and U15865 (N_15865,N_15475,N_15049);
and U15866 (N_15866,N_15117,N_15312);
xor U15867 (N_15867,N_15071,N_15481);
and U15868 (N_15868,N_15088,N_15387);
and U15869 (N_15869,N_15337,N_15111);
xor U15870 (N_15870,N_15040,N_15376);
nor U15871 (N_15871,N_15064,N_15002);
and U15872 (N_15872,N_15435,N_15144);
and U15873 (N_15873,N_15411,N_15292);
nand U15874 (N_15874,N_15287,N_15390);
nor U15875 (N_15875,N_15484,N_15023);
xnor U15876 (N_15876,N_15226,N_15477);
nor U15877 (N_15877,N_15037,N_15273);
nor U15878 (N_15878,N_15111,N_15259);
or U15879 (N_15879,N_15241,N_15049);
nor U15880 (N_15880,N_15085,N_15339);
or U15881 (N_15881,N_15433,N_15287);
nor U15882 (N_15882,N_15107,N_15218);
and U15883 (N_15883,N_15123,N_15047);
or U15884 (N_15884,N_15200,N_15012);
xnor U15885 (N_15885,N_15063,N_15051);
nand U15886 (N_15886,N_15131,N_15311);
and U15887 (N_15887,N_15443,N_15156);
xor U15888 (N_15888,N_15333,N_15243);
nor U15889 (N_15889,N_15008,N_15183);
nand U15890 (N_15890,N_15272,N_15360);
and U15891 (N_15891,N_15492,N_15478);
nand U15892 (N_15892,N_15453,N_15288);
nand U15893 (N_15893,N_15412,N_15046);
nand U15894 (N_15894,N_15468,N_15014);
xor U15895 (N_15895,N_15229,N_15465);
or U15896 (N_15896,N_15358,N_15340);
nand U15897 (N_15897,N_15259,N_15460);
nand U15898 (N_15898,N_15324,N_15121);
and U15899 (N_15899,N_15195,N_15244);
nand U15900 (N_15900,N_15235,N_15439);
nor U15901 (N_15901,N_15201,N_15104);
and U15902 (N_15902,N_15021,N_15278);
nand U15903 (N_15903,N_15177,N_15030);
or U15904 (N_15904,N_15039,N_15383);
nor U15905 (N_15905,N_15073,N_15364);
nor U15906 (N_15906,N_15122,N_15377);
nand U15907 (N_15907,N_15250,N_15355);
xor U15908 (N_15908,N_15271,N_15492);
or U15909 (N_15909,N_15140,N_15438);
or U15910 (N_15910,N_15499,N_15046);
nand U15911 (N_15911,N_15444,N_15145);
xnor U15912 (N_15912,N_15432,N_15150);
nand U15913 (N_15913,N_15049,N_15419);
or U15914 (N_15914,N_15465,N_15342);
nand U15915 (N_15915,N_15032,N_15411);
nor U15916 (N_15916,N_15394,N_15203);
or U15917 (N_15917,N_15017,N_15248);
nand U15918 (N_15918,N_15006,N_15001);
nor U15919 (N_15919,N_15005,N_15102);
or U15920 (N_15920,N_15116,N_15358);
nor U15921 (N_15921,N_15421,N_15230);
or U15922 (N_15922,N_15019,N_15444);
or U15923 (N_15923,N_15402,N_15069);
nor U15924 (N_15924,N_15102,N_15253);
and U15925 (N_15925,N_15061,N_15375);
nor U15926 (N_15926,N_15174,N_15425);
nand U15927 (N_15927,N_15176,N_15422);
nor U15928 (N_15928,N_15090,N_15213);
nand U15929 (N_15929,N_15123,N_15390);
or U15930 (N_15930,N_15285,N_15249);
nor U15931 (N_15931,N_15037,N_15020);
and U15932 (N_15932,N_15185,N_15264);
nand U15933 (N_15933,N_15236,N_15096);
and U15934 (N_15934,N_15118,N_15093);
and U15935 (N_15935,N_15335,N_15058);
and U15936 (N_15936,N_15363,N_15281);
xnor U15937 (N_15937,N_15475,N_15392);
or U15938 (N_15938,N_15009,N_15384);
xor U15939 (N_15939,N_15122,N_15162);
and U15940 (N_15940,N_15358,N_15177);
nand U15941 (N_15941,N_15235,N_15390);
nor U15942 (N_15942,N_15360,N_15270);
and U15943 (N_15943,N_15176,N_15213);
and U15944 (N_15944,N_15352,N_15156);
or U15945 (N_15945,N_15036,N_15420);
and U15946 (N_15946,N_15301,N_15457);
nor U15947 (N_15947,N_15090,N_15243);
xnor U15948 (N_15948,N_15396,N_15056);
nor U15949 (N_15949,N_15220,N_15115);
xnor U15950 (N_15950,N_15146,N_15375);
nor U15951 (N_15951,N_15493,N_15183);
xnor U15952 (N_15952,N_15190,N_15270);
and U15953 (N_15953,N_15319,N_15218);
and U15954 (N_15954,N_15417,N_15431);
or U15955 (N_15955,N_15051,N_15171);
and U15956 (N_15956,N_15138,N_15440);
nand U15957 (N_15957,N_15092,N_15280);
or U15958 (N_15958,N_15323,N_15165);
or U15959 (N_15959,N_15173,N_15422);
nor U15960 (N_15960,N_15045,N_15150);
or U15961 (N_15961,N_15284,N_15258);
and U15962 (N_15962,N_15242,N_15464);
or U15963 (N_15963,N_15194,N_15006);
or U15964 (N_15964,N_15066,N_15230);
nor U15965 (N_15965,N_15484,N_15482);
nor U15966 (N_15966,N_15179,N_15321);
nor U15967 (N_15967,N_15039,N_15059);
nand U15968 (N_15968,N_15293,N_15294);
or U15969 (N_15969,N_15404,N_15004);
and U15970 (N_15970,N_15133,N_15303);
xor U15971 (N_15971,N_15497,N_15175);
nor U15972 (N_15972,N_15177,N_15386);
nor U15973 (N_15973,N_15071,N_15276);
and U15974 (N_15974,N_15050,N_15400);
xor U15975 (N_15975,N_15076,N_15091);
and U15976 (N_15976,N_15300,N_15320);
or U15977 (N_15977,N_15026,N_15377);
xnor U15978 (N_15978,N_15398,N_15110);
nor U15979 (N_15979,N_15149,N_15331);
and U15980 (N_15980,N_15407,N_15383);
or U15981 (N_15981,N_15247,N_15123);
and U15982 (N_15982,N_15320,N_15238);
or U15983 (N_15983,N_15229,N_15479);
nor U15984 (N_15984,N_15214,N_15198);
or U15985 (N_15985,N_15291,N_15427);
nand U15986 (N_15986,N_15204,N_15134);
and U15987 (N_15987,N_15436,N_15076);
and U15988 (N_15988,N_15157,N_15446);
nor U15989 (N_15989,N_15239,N_15321);
xor U15990 (N_15990,N_15344,N_15094);
or U15991 (N_15991,N_15195,N_15329);
nor U15992 (N_15992,N_15461,N_15201);
or U15993 (N_15993,N_15368,N_15124);
xnor U15994 (N_15994,N_15128,N_15171);
or U15995 (N_15995,N_15344,N_15365);
and U15996 (N_15996,N_15115,N_15411);
or U15997 (N_15997,N_15379,N_15253);
and U15998 (N_15998,N_15002,N_15033);
or U15999 (N_15999,N_15368,N_15178);
nor U16000 (N_16000,N_15969,N_15551);
nor U16001 (N_16001,N_15596,N_15783);
nor U16002 (N_16002,N_15982,N_15930);
or U16003 (N_16003,N_15534,N_15537);
or U16004 (N_16004,N_15713,N_15543);
nand U16005 (N_16005,N_15999,N_15791);
nand U16006 (N_16006,N_15950,N_15861);
nor U16007 (N_16007,N_15769,N_15943);
and U16008 (N_16008,N_15604,N_15709);
nor U16009 (N_16009,N_15504,N_15587);
xor U16010 (N_16010,N_15839,N_15581);
and U16011 (N_16011,N_15585,N_15641);
or U16012 (N_16012,N_15571,N_15984);
and U16013 (N_16013,N_15664,N_15561);
nor U16014 (N_16014,N_15921,N_15723);
nand U16015 (N_16015,N_15647,N_15883);
nor U16016 (N_16016,N_15817,N_15759);
nand U16017 (N_16017,N_15846,N_15805);
xor U16018 (N_16018,N_15795,N_15570);
and U16019 (N_16019,N_15563,N_15755);
or U16020 (N_16020,N_15955,N_15710);
xor U16021 (N_16021,N_15716,N_15597);
nand U16022 (N_16022,N_15699,N_15559);
or U16023 (N_16023,N_15836,N_15888);
nand U16024 (N_16024,N_15612,N_15514);
nor U16025 (N_16025,N_15764,N_15960);
nand U16026 (N_16026,N_15756,N_15794);
nand U16027 (N_16027,N_15936,N_15761);
xnor U16028 (N_16028,N_15981,N_15864);
or U16029 (N_16029,N_15757,N_15568);
xnor U16030 (N_16030,N_15607,N_15816);
and U16031 (N_16031,N_15944,N_15935);
nor U16032 (N_16032,N_15517,N_15815);
nor U16033 (N_16033,N_15626,N_15547);
and U16034 (N_16034,N_15698,N_15535);
xor U16035 (N_16035,N_15859,N_15851);
or U16036 (N_16036,N_15747,N_15745);
nand U16037 (N_16037,N_15988,N_15826);
xor U16038 (N_16038,N_15727,N_15951);
nand U16039 (N_16039,N_15733,N_15925);
xnor U16040 (N_16040,N_15601,N_15555);
nand U16041 (N_16041,N_15825,N_15767);
nand U16042 (N_16042,N_15998,N_15651);
or U16043 (N_16043,N_15676,N_15506);
xnor U16044 (N_16044,N_15758,N_15661);
or U16045 (N_16045,N_15746,N_15763);
nor U16046 (N_16046,N_15541,N_15917);
xor U16047 (N_16047,N_15558,N_15688);
nand U16048 (N_16048,N_15516,N_15907);
or U16049 (N_16049,N_15569,N_15693);
and U16050 (N_16050,N_15913,N_15734);
or U16051 (N_16051,N_15616,N_15515);
nand U16052 (N_16052,N_15949,N_15670);
nor U16053 (N_16053,N_15659,N_15971);
and U16054 (N_16054,N_15726,N_15995);
and U16055 (N_16055,N_15731,N_15831);
xor U16056 (N_16056,N_15674,N_15735);
xor U16057 (N_16057,N_15991,N_15625);
and U16058 (N_16058,N_15793,N_15802);
xor U16059 (N_16059,N_15738,N_15784);
xnor U16060 (N_16060,N_15961,N_15885);
nor U16061 (N_16061,N_15752,N_15941);
nand U16062 (N_16062,N_15806,N_15507);
and U16063 (N_16063,N_15821,N_15583);
xnor U16064 (N_16064,N_15781,N_15617);
nor U16065 (N_16065,N_15695,N_15832);
xor U16066 (N_16066,N_15939,N_15989);
and U16067 (N_16067,N_15584,N_15855);
or U16068 (N_16068,N_15655,N_15512);
and U16069 (N_16069,N_15849,N_15744);
and U16070 (N_16070,N_15690,N_15996);
xnor U16071 (N_16071,N_15639,N_15990);
and U16072 (N_16072,N_15798,N_15954);
nand U16073 (N_16073,N_15813,N_15714);
nor U16074 (N_16074,N_15788,N_15508);
nand U16075 (N_16075,N_15994,N_15980);
and U16076 (N_16076,N_15653,N_15526);
nand U16077 (N_16077,N_15818,N_15657);
nand U16078 (N_16078,N_15860,N_15611);
or U16079 (N_16079,N_15751,N_15997);
nand U16080 (N_16080,N_15685,N_15856);
xor U16081 (N_16081,N_15683,N_15536);
or U16082 (N_16082,N_15684,N_15705);
or U16083 (N_16083,N_15932,N_15622);
nand U16084 (N_16084,N_15775,N_15533);
xnor U16085 (N_16085,N_15841,N_15681);
and U16086 (N_16086,N_15545,N_15829);
or U16087 (N_16087,N_15708,N_15992);
xor U16088 (N_16088,N_15500,N_15503);
and U16089 (N_16089,N_15636,N_15728);
nor U16090 (N_16090,N_15777,N_15801);
or U16091 (N_16091,N_15696,N_15530);
nand U16092 (N_16092,N_15787,N_15579);
nand U16093 (N_16093,N_15656,N_15598);
xor U16094 (N_16094,N_15863,N_15706);
nor U16095 (N_16095,N_15874,N_15901);
nor U16096 (N_16096,N_15799,N_15770);
nor U16097 (N_16097,N_15965,N_15934);
xor U16098 (N_16098,N_15729,N_15593);
or U16099 (N_16099,N_15672,N_15887);
and U16100 (N_16100,N_15986,N_15987);
nand U16101 (N_16101,N_15910,N_15619);
nand U16102 (N_16102,N_15892,N_15968);
and U16103 (N_16103,N_15704,N_15848);
nor U16104 (N_16104,N_15635,N_15608);
nor U16105 (N_16105,N_15527,N_15976);
and U16106 (N_16106,N_15665,N_15948);
nand U16107 (N_16107,N_15889,N_15890);
nor U16108 (N_16108,N_15947,N_15592);
nor U16109 (N_16109,N_15937,N_15700);
nor U16110 (N_16110,N_15771,N_15689);
nand U16111 (N_16111,N_15804,N_15953);
xnor U16112 (N_16112,N_15623,N_15786);
and U16113 (N_16113,N_15509,N_15800);
nand U16114 (N_16114,N_15737,N_15675);
and U16115 (N_16115,N_15966,N_15580);
or U16116 (N_16116,N_15754,N_15518);
or U16117 (N_16117,N_15796,N_15712);
and U16118 (N_16118,N_15896,N_15511);
nor U16119 (N_16119,N_15605,N_15797);
and U16120 (N_16120,N_15834,N_15642);
or U16121 (N_16121,N_15573,N_15828);
xnor U16122 (N_16122,N_15915,N_15865);
nor U16123 (N_16123,N_15557,N_15654);
xnor U16124 (N_16124,N_15790,N_15808);
xnor U16125 (N_16125,N_15906,N_15835);
nand U16126 (N_16126,N_15614,N_15565);
or U16127 (N_16127,N_15590,N_15602);
xnor U16128 (N_16128,N_15720,N_15524);
nor U16129 (N_16129,N_15967,N_15721);
xnor U16130 (N_16130,N_15959,N_15697);
nor U16131 (N_16131,N_15594,N_15680);
and U16132 (N_16132,N_15567,N_15538);
and U16133 (N_16133,N_15868,N_15750);
nand U16134 (N_16134,N_15753,N_15926);
or U16135 (N_16135,N_15633,N_15898);
and U16136 (N_16136,N_15975,N_15631);
or U16137 (N_16137,N_15502,N_15717);
nor U16138 (N_16138,N_15927,N_15958);
xnor U16139 (N_16139,N_15844,N_15707);
or U16140 (N_16140,N_15814,N_15933);
or U16141 (N_16141,N_15867,N_15615);
nand U16142 (N_16142,N_15785,N_15586);
nor U16143 (N_16143,N_15748,N_15918);
nand U16144 (N_16144,N_15609,N_15519);
and U16145 (N_16145,N_15810,N_15629);
xnor U16146 (N_16146,N_15760,N_15811);
nor U16147 (N_16147,N_15591,N_15682);
nor U16148 (N_16148,N_15701,N_15776);
and U16149 (N_16149,N_15722,N_15973);
nand U16150 (N_16150,N_15956,N_15854);
nor U16151 (N_16151,N_15852,N_15599);
nor U16152 (N_16152,N_15879,N_15556);
nor U16153 (N_16153,N_15673,N_15575);
nor U16154 (N_16154,N_15692,N_15725);
nor U16155 (N_16155,N_15938,N_15550);
xnor U16156 (N_16156,N_15691,N_15539);
nand U16157 (N_16157,N_15897,N_15895);
or U16158 (N_16158,N_15711,N_15866);
and U16159 (N_16159,N_15902,N_15830);
or U16160 (N_16160,N_15899,N_15715);
nand U16161 (N_16161,N_15658,N_15627);
nor U16162 (N_16162,N_15838,N_15827);
xnor U16163 (N_16163,N_15595,N_15566);
xor U16164 (N_16164,N_15732,N_15552);
and U16165 (N_16165,N_15606,N_15946);
xor U16166 (N_16166,N_15924,N_15544);
xnor U16167 (N_16167,N_15807,N_15853);
or U16168 (N_16168,N_15650,N_15893);
or U16169 (N_16169,N_15553,N_15529);
or U16170 (N_16170,N_15677,N_15979);
or U16171 (N_16171,N_15873,N_15719);
or U16172 (N_16172,N_15678,N_15875);
or U16173 (N_16173,N_15978,N_15513);
nor U16174 (N_16174,N_15974,N_15876);
or U16175 (N_16175,N_15572,N_15962);
nand U16176 (N_16176,N_15869,N_15576);
and U16177 (N_16177,N_15923,N_15880);
nand U16178 (N_16178,N_15600,N_15778);
nand U16179 (N_16179,N_15643,N_15803);
xnor U16180 (N_16180,N_15621,N_15909);
and U16181 (N_16181,N_15894,N_15779);
nand U16182 (N_16182,N_15850,N_15522);
xnor U16183 (N_16183,N_15702,N_15662);
and U16184 (N_16184,N_15645,N_15667);
nor U16185 (N_16185,N_15970,N_15822);
or U16186 (N_16186,N_15877,N_15789);
and U16187 (N_16187,N_15884,N_15718);
xnor U16188 (N_16188,N_15542,N_15774);
and U16189 (N_16189,N_15520,N_15574);
xor U16190 (N_16190,N_15847,N_15582);
nor U16191 (N_16191,N_15531,N_15765);
xor U16192 (N_16192,N_15963,N_15687);
or U16193 (N_16193,N_15510,N_15549);
nor U16194 (N_16194,N_15964,N_15928);
or U16195 (N_16195,N_15843,N_15858);
and U16196 (N_16196,N_15773,N_15686);
xnor U16197 (N_16197,N_15837,N_15546);
and U16198 (N_16198,N_15819,N_15501);
nor U16199 (N_16199,N_15620,N_15812);
nor U16200 (N_16200,N_15916,N_15630);
or U16201 (N_16201,N_15548,N_15741);
and U16202 (N_16202,N_15603,N_15782);
or U16203 (N_16203,N_15945,N_15912);
or U16204 (N_16204,N_15624,N_15862);
and U16205 (N_16205,N_15532,N_15618);
and U16206 (N_16206,N_15881,N_15983);
nand U16207 (N_16207,N_15820,N_15554);
and U16208 (N_16208,N_15649,N_15957);
nand U16209 (N_16209,N_15823,N_15766);
and U16210 (N_16210,N_15588,N_15919);
nand U16211 (N_16211,N_15900,N_15564);
nor U16212 (N_16212,N_15740,N_15628);
xnor U16213 (N_16213,N_15809,N_15668);
xor U16214 (N_16214,N_15914,N_15613);
nand U16215 (N_16215,N_15644,N_15922);
xnor U16216 (N_16216,N_15666,N_15882);
or U16217 (N_16217,N_15905,N_15505);
xor U16218 (N_16218,N_15857,N_15952);
or U16219 (N_16219,N_15525,N_15993);
nor U16220 (N_16220,N_15872,N_15640);
nor U16221 (N_16221,N_15660,N_15736);
nor U16222 (N_16222,N_15942,N_15560);
and U16223 (N_16223,N_15878,N_15792);
nand U16224 (N_16224,N_15772,N_15703);
and U16225 (N_16225,N_15562,N_15833);
nor U16226 (N_16226,N_15637,N_15931);
xor U16227 (N_16227,N_15679,N_15652);
and U16228 (N_16228,N_15972,N_15929);
xnor U16229 (N_16229,N_15648,N_15768);
nand U16230 (N_16230,N_15908,N_15743);
and U16231 (N_16231,N_15646,N_15870);
nand U16232 (N_16232,N_15578,N_15871);
and U16233 (N_16233,N_15824,N_15920);
or U16234 (N_16234,N_15891,N_15528);
xnor U16235 (N_16235,N_15638,N_15886);
nand U16236 (N_16236,N_15840,N_15739);
or U16237 (N_16237,N_15730,N_15749);
and U16238 (N_16238,N_15742,N_15523);
and U16239 (N_16239,N_15589,N_15663);
and U16240 (N_16240,N_15780,N_15694);
or U16241 (N_16241,N_15904,N_15632);
or U16242 (N_16242,N_15634,N_15610);
and U16243 (N_16243,N_15842,N_15577);
or U16244 (N_16244,N_15762,N_15911);
or U16245 (N_16245,N_15903,N_15940);
xor U16246 (N_16246,N_15724,N_15985);
nor U16247 (N_16247,N_15977,N_15845);
and U16248 (N_16248,N_15521,N_15669);
nand U16249 (N_16249,N_15671,N_15540);
xor U16250 (N_16250,N_15760,N_15698);
or U16251 (N_16251,N_15701,N_15709);
and U16252 (N_16252,N_15935,N_15762);
nand U16253 (N_16253,N_15622,N_15631);
and U16254 (N_16254,N_15931,N_15849);
or U16255 (N_16255,N_15678,N_15689);
nor U16256 (N_16256,N_15583,N_15736);
nand U16257 (N_16257,N_15549,N_15835);
nor U16258 (N_16258,N_15721,N_15957);
nor U16259 (N_16259,N_15921,N_15608);
xnor U16260 (N_16260,N_15902,N_15743);
and U16261 (N_16261,N_15582,N_15871);
or U16262 (N_16262,N_15891,N_15710);
xor U16263 (N_16263,N_15601,N_15901);
or U16264 (N_16264,N_15914,N_15810);
nand U16265 (N_16265,N_15501,N_15695);
xor U16266 (N_16266,N_15954,N_15782);
or U16267 (N_16267,N_15645,N_15590);
nand U16268 (N_16268,N_15881,N_15696);
nor U16269 (N_16269,N_15949,N_15918);
nand U16270 (N_16270,N_15530,N_15682);
or U16271 (N_16271,N_15914,N_15698);
nand U16272 (N_16272,N_15504,N_15987);
nor U16273 (N_16273,N_15741,N_15575);
and U16274 (N_16274,N_15645,N_15654);
xor U16275 (N_16275,N_15962,N_15687);
nand U16276 (N_16276,N_15587,N_15778);
and U16277 (N_16277,N_15608,N_15831);
xnor U16278 (N_16278,N_15623,N_15961);
nor U16279 (N_16279,N_15787,N_15626);
xnor U16280 (N_16280,N_15785,N_15530);
and U16281 (N_16281,N_15594,N_15738);
or U16282 (N_16282,N_15503,N_15665);
nand U16283 (N_16283,N_15894,N_15569);
nand U16284 (N_16284,N_15748,N_15775);
and U16285 (N_16285,N_15642,N_15813);
xor U16286 (N_16286,N_15605,N_15526);
nor U16287 (N_16287,N_15834,N_15929);
nand U16288 (N_16288,N_15655,N_15621);
and U16289 (N_16289,N_15869,N_15527);
nor U16290 (N_16290,N_15700,N_15541);
or U16291 (N_16291,N_15935,N_15719);
and U16292 (N_16292,N_15850,N_15992);
or U16293 (N_16293,N_15861,N_15771);
or U16294 (N_16294,N_15877,N_15670);
or U16295 (N_16295,N_15769,N_15507);
and U16296 (N_16296,N_15620,N_15993);
and U16297 (N_16297,N_15597,N_15797);
or U16298 (N_16298,N_15872,N_15675);
and U16299 (N_16299,N_15931,N_15838);
and U16300 (N_16300,N_15667,N_15957);
and U16301 (N_16301,N_15918,N_15637);
or U16302 (N_16302,N_15916,N_15573);
nor U16303 (N_16303,N_15762,N_15958);
or U16304 (N_16304,N_15677,N_15664);
nor U16305 (N_16305,N_15796,N_15819);
and U16306 (N_16306,N_15625,N_15739);
and U16307 (N_16307,N_15647,N_15785);
nor U16308 (N_16308,N_15955,N_15910);
xor U16309 (N_16309,N_15958,N_15541);
nand U16310 (N_16310,N_15577,N_15708);
xnor U16311 (N_16311,N_15738,N_15960);
nor U16312 (N_16312,N_15839,N_15933);
or U16313 (N_16313,N_15788,N_15917);
nand U16314 (N_16314,N_15654,N_15964);
nor U16315 (N_16315,N_15732,N_15544);
nor U16316 (N_16316,N_15712,N_15644);
or U16317 (N_16317,N_15537,N_15878);
and U16318 (N_16318,N_15943,N_15966);
or U16319 (N_16319,N_15650,N_15685);
nand U16320 (N_16320,N_15688,N_15819);
or U16321 (N_16321,N_15919,N_15594);
or U16322 (N_16322,N_15536,N_15626);
and U16323 (N_16323,N_15925,N_15929);
or U16324 (N_16324,N_15843,N_15673);
and U16325 (N_16325,N_15653,N_15856);
and U16326 (N_16326,N_15845,N_15729);
xnor U16327 (N_16327,N_15568,N_15817);
nor U16328 (N_16328,N_15795,N_15920);
and U16329 (N_16329,N_15883,N_15902);
and U16330 (N_16330,N_15684,N_15949);
and U16331 (N_16331,N_15901,N_15730);
or U16332 (N_16332,N_15535,N_15669);
and U16333 (N_16333,N_15603,N_15920);
nor U16334 (N_16334,N_15842,N_15917);
or U16335 (N_16335,N_15750,N_15814);
nor U16336 (N_16336,N_15540,N_15607);
nor U16337 (N_16337,N_15600,N_15654);
xnor U16338 (N_16338,N_15932,N_15776);
xnor U16339 (N_16339,N_15773,N_15951);
and U16340 (N_16340,N_15900,N_15607);
and U16341 (N_16341,N_15834,N_15728);
nor U16342 (N_16342,N_15771,N_15508);
and U16343 (N_16343,N_15834,N_15811);
or U16344 (N_16344,N_15934,N_15584);
xnor U16345 (N_16345,N_15917,N_15717);
and U16346 (N_16346,N_15969,N_15998);
nor U16347 (N_16347,N_15818,N_15762);
or U16348 (N_16348,N_15600,N_15522);
or U16349 (N_16349,N_15895,N_15790);
nand U16350 (N_16350,N_15950,N_15573);
nand U16351 (N_16351,N_15828,N_15981);
xnor U16352 (N_16352,N_15709,N_15567);
or U16353 (N_16353,N_15919,N_15693);
xnor U16354 (N_16354,N_15838,N_15536);
and U16355 (N_16355,N_15996,N_15903);
and U16356 (N_16356,N_15734,N_15888);
nor U16357 (N_16357,N_15650,N_15665);
nand U16358 (N_16358,N_15871,N_15654);
or U16359 (N_16359,N_15948,N_15557);
nand U16360 (N_16360,N_15617,N_15867);
xnor U16361 (N_16361,N_15605,N_15592);
xor U16362 (N_16362,N_15701,N_15789);
and U16363 (N_16363,N_15503,N_15891);
xnor U16364 (N_16364,N_15945,N_15981);
or U16365 (N_16365,N_15797,N_15600);
xnor U16366 (N_16366,N_15644,N_15844);
nor U16367 (N_16367,N_15523,N_15547);
or U16368 (N_16368,N_15958,N_15887);
nand U16369 (N_16369,N_15556,N_15783);
nor U16370 (N_16370,N_15941,N_15698);
xnor U16371 (N_16371,N_15701,N_15860);
and U16372 (N_16372,N_15798,N_15665);
nor U16373 (N_16373,N_15584,N_15547);
or U16374 (N_16374,N_15994,N_15703);
and U16375 (N_16375,N_15806,N_15687);
nor U16376 (N_16376,N_15657,N_15627);
xnor U16377 (N_16377,N_15688,N_15892);
nor U16378 (N_16378,N_15958,N_15609);
nand U16379 (N_16379,N_15778,N_15596);
nor U16380 (N_16380,N_15511,N_15965);
xor U16381 (N_16381,N_15606,N_15889);
xor U16382 (N_16382,N_15946,N_15962);
and U16383 (N_16383,N_15724,N_15833);
xor U16384 (N_16384,N_15892,N_15859);
xnor U16385 (N_16385,N_15592,N_15749);
nand U16386 (N_16386,N_15801,N_15733);
nor U16387 (N_16387,N_15852,N_15660);
xnor U16388 (N_16388,N_15742,N_15984);
xor U16389 (N_16389,N_15815,N_15662);
nor U16390 (N_16390,N_15916,N_15624);
nand U16391 (N_16391,N_15865,N_15749);
or U16392 (N_16392,N_15942,N_15867);
nand U16393 (N_16393,N_15802,N_15911);
xnor U16394 (N_16394,N_15714,N_15705);
and U16395 (N_16395,N_15879,N_15598);
or U16396 (N_16396,N_15518,N_15841);
and U16397 (N_16397,N_15644,N_15770);
nand U16398 (N_16398,N_15968,N_15948);
and U16399 (N_16399,N_15594,N_15560);
nand U16400 (N_16400,N_15520,N_15740);
nor U16401 (N_16401,N_15556,N_15705);
and U16402 (N_16402,N_15657,N_15752);
xnor U16403 (N_16403,N_15885,N_15628);
nor U16404 (N_16404,N_15750,N_15747);
nor U16405 (N_16405,N_15663,N_15768);
or U16406 (N_16406,N_15825,N_15736);
xnor U16407 (N_16407,N_15533,N_15754);
nor U16408 (N_16408,N_15722,N_15792);
nand U16409 (N_16409,N_15562,N_15507);
xor U16410 (N_16410,N_15967,N_15514);
nor U16411 (N_16411,N_15931,N_15740);
nor U16412 (N_16412,N_15817,N_15618);
xor U16413 (N_16413,N_15799,N_15709);
nand U16414 (N_16414,N_15830,N_15645);
xor U16415 (N_16415,N_15593,N_15987);
xor U16416 (N_16416,N_15883,N_15776);
and U16417 (N_16417,N_15903,N_15922);
nor U16418 (N_16418,N_15811,N_15979);
or U16419 (N_16419,N_15709,N_15736);
xor U16420 (N_16420,N_15916,N_15589);
xnor U16421 (N_16421,N_15931,N_15990);
or U16422 (N_16422,N_15968,N_15652);
and U16423 (N_16423,N_15877,N_15513);
xnor U16424 (N_16424,N_15975,N_15869);
or U16425 (N_16425,N_15899,N_15620);
or U16426 (N_16426,N_15917,N_15525);
nor U16427 (N_16427,N_15535,N_15764);
nor U16428 (N_16428,N_15768,N_15971);
xor U16429 (N_16429,N_15895,N_15941);
and U16430 (N_16430,N_15500,N_15651);
and U16431 (N_16431,N_15851,N_15863);
and U16432 (N_16432,N_15995,N_15978);
or U16433 (N_16433,N_15954,N_15810);
nand U16434 (N_16434,N_15659,N_15535);
and U16435 (N_16435,N_15565,N_15523);
nand U16436 (N_16436,N_15701,N_15788);
nand U16437 (N_16437,N_15916,N_15893);
xnor U16438 (N_16438,N_15943,N_15801);
or U16439 (N_16439,N_15559,N_15757);
xnor U16440 (N_16440,N_15809,N_15644);
and U16441 (N_16441,N_15760,N_15931);
xnor U16442 (N_16442,N_15930,N_15537);
xor U16443 (N_16443,N_15699,N_15673);
or U16444 (N_16444,N_15556,N_15665);
xnor U16445 (N_16445,N_15760,N_15739);
xnor U16446 (N_16446,N_15678,N_15606);
and U16447 (N_16447,N_15592,N_15815);
nand U16448 (N_16448,N_15662,N_15549);
nor U16449 (N_16449,N_15876,N_15677);
nand U16450 (N_16450,N_15995,N_15611);
xor U16451 (N_16451,N_15521,N_15737);
and U16452 (N_16452,N_15951,N_15947);
xnor U16453 (N_16453,N_15867,N_15669);
or U16454 (N_16454,N_15845,N_15582);
nand U16455 (N_16455,N_15509,N_15874);
nor U16456 (N_16456,N_15614,N_15871);
or U16457 (N_16457,N_15707,N_15895);
nand U16458 (N_16458,N_15741,N_15642);
nor U16459 (N_16459,N_15810,N_15509);
or U16460 (N_16460,N_15582,N_15904);
xnor U16461 (N_16461,N_15574,N_15617);
nor U16462 (N_16462,N_15535,N_15645);
and U16463 (N_16463,N_15511,N_15715);
or U16464 (N_16464,N_15751,N_15695);
and U16465 (N_16465,N_15651,N_15563);
and U16466 (N_16466,N_15805,N_15568);
and U16467 (N_16467,N_15777,N_15620);
nor U16468 (N_16468,N_15633,N_15924);
xor U16469 (N_16469,N_15956,N_15545);
nand U16470 (N_16470,N_15589,N_15668);
nand U16471 (N_16471,N_15695,N_15800);
xnor U16472 (N_16472,N_15501,N_15861);
nor U16473 (N_16473,N_15758,N_15586);
and U16474 (N_16474,N_15788,N_15506);
nor U16475 (N_16475,N_15751,N_15834);
nor U16476 (N_16476,N_15702,N_15809);
nand U16477 (N_16477,N_15599,N_15885);
nand U16478 (N_16478,N_15785,N_15659);
nor U16479 (N_16479,N_15890,N_15993);
or U16480 (N_16480,N_15631,N_15908);
nand U16481 (N_16481,N_15606,N_15809);
nor U16482 (N_16482,N_15963,N_15822);
nand U16483 (N_16483,N_15988,N_15790);
nand U16484 (N_16484,N_15678,N_15568);
and U16485 (N_16485,N_15545,N_15714);
and U16486 (N_16486,N_15822,N_15865);
nand U16487 (N_16487,N_15602,N_15839);
nand U16488 (N_16488,N_15955,N_15582);
or U16489 (N_16489,N_15864,N_15770);
xnor U16490 (N_16490,N_15650,N_15620);
and U16491 (N_16491,N_15908,N_15770);
nand U16492 (N_16492,N_15682,N_15769);
and U16493 (N_16493,N_15889,N_15501);
and U16494 (N_16494,N_15528,N_15811);
or U16495 (N_16495,N_15861,N_15587);
xnor U16496 (N_16496,N_15696,N_15506);
and U16497 (N_16497,N_15527,N_15921);
xnor U16498 (N_16498,N_15842,N_15621);
and U16499 (N_16499,N_15775,N_15984);
or U16500 (N_16500,N_16363,N_16123);
nor U16501 (N_16501,N_16168,N_16378);
and U16502 (N_16502,N_16241,N_16099);
nand U16503 (N_16503,N_16266,N_16333);
and U16504 (N_16504,N_16461,N_16190);
xor U16505 (N_16505,N_16237,N_16196);
and U16506 (N_16506,N_16351,N_16205);
xnor U16507 (N_16507,N_16213,N_16398);
nor U16508 (N_16508,N_16222,N_16456);
or U16509 (N_16509,N_16267,N_16125);
nor U16510 (N_16510,N_16150,N_16498);
nor U16511 (N_16511,N_16252,N_16119);
or U16512 (N_16512,N_16175,N_16288);
nor U16513 (N_16513,N_16298,N_16373);
xor U16514 (N_16514,N_16256,N_16491);
nor U16515 (N_16515,N_16407,N_16146);
nor U16516 (N_16516,N_16318,N_16199);
nand U16517 (N_16517,N_16272,N_16321);
and U16518 (N_16518,N_16035,N_16376);
nor U16519 (N_16519,N_16496,N_16102);
or U16520 (N_16520,N_16105,N_16019);
and U16521 (N_16521,N_16460,N_16081);
and U16522 (N_16522,N_16417,N_16446);
nor U16523 (N_16523,N_16142,N_16157);
nand U16524 (N_16524,N_16499,N_16039);
nand U16525 (N_16525,N_16480,N_16313);
xor U16526 (N_16526,N_16463,N_16184);
and U16527 (N_16527,N_16476,N_16438);
nor U16528 (N_16528,N_16051,N_16330);
and U16529 (N_16529,N_16218,N_16185);
or U16530 (N_16530,N_16067,N_16250);
nor U16531 (N_16531,N_16022,N_16061);
nor U16532 (N_16532,N_16354,N_16308);
nor U16533 (N_16533,N_16377,N_16064);
nor U16534 (N_16534,N_16270,N_16197);
xor U16535 (N_16535,N_16207,N_16134);
or U16536 (N_16536,N_16301,N_16093);
and U16537 (N_16537,N_16012,N_16046);
xnor U16538 (N_16538,N_16443,N_16489);
and U16539 (N_16539,N_16231,N_16486);
and U16540 (N_16540,N_16140,N_16158);
and U16541 (N_16541,N_16278,N_16088);
nor U16542 (N_16542,N_16441,N_16089);
nor U16543 (N_16543,N_16478,N_16467);
nand U16544 (N_16544,N_16450,N_16208);
nand U16545 (N_16545,N_16018,N_16139);
or U16546 (N_16546,N_16405,N_16385);
xor U16547 (N_16547,N_16317,N_16495);
nor U16548 (N_16548,N_16397,N_16442);
or U16549 (N_16549,N_16282,N_16118);
and U16550 (N_16550,N_16364,N_16217);
nor U16551 (N_16551,N_16116,N_16429);
nor U16552 (N_16552,N_16257,N_16269);
nor U16553 (N_16553,N_16437,N_16179);
nor U16554 (N_16554,N_16078,N_16017);
or U16555 (N_16555,N_16328,N_16249);
or U16556 (N_16556,N_16043,N_16127);
xnor U16557 (N_16557,N_16126,N_16128);
or U16558 (N_16558,N_16007,N_16242);
nand U16559 (N_16559,N_16220,N_16409);
nor U16560 (N_16560,N_16041,N_16448);
nor U16561 (N_16561,N_16106,N_16014);
nor U16562 (N_16562,N_16396,N_16477);
nor U16563 (N_16563,N_16097,N_16466);
or U16564 (N_16564,N_16284,N_16003);
xnor U16565 (N_16565,N_16245,N_16246);
nand U16566 (N_16566,N_16255,N_16136);
and U16567 (N_16567,N_16493,N_16206);
nand U16568 (N_16568,N_16183,N_16280);
xnor U16569 (N_16569,N_16411,N_16037);
nand U16570 (N_16570,N_16482,N_16268);
or U16571 (N_16571,N_16144,N_16188);
xnor U16572 (N_16572,N_16165,N_16164);
xor U16573 (N_16573,N_16030,N_16204);
nor U16574 (N_16574,N_16389,N_16294);
nand U16575 (N_16575,N_16350,N_16178);
xnor U16576 (N_16576,N_16391,N_16264);
xnor U16577 (N_16577,N_16054,N_16044);
nor U16578 (N_16578,N_16420,N_16015);
and U16579 (N_16579,N_16327,N_16345);
nand U16580 (N_16580,N_16173,N_16349);
xnor U16581 (N_16581,N_16445,N_16388);
and U16582 (N_16582,N_16110,N_16332);
or U16583 (N_16583,N_16274,N_16152);
and U16584 (N_16584,N_16113,N_16342);
or U16585 (N_16585,N_16029,N_16481);
xor U16586 (N_16586,N_16135,N_16132);
nand U16587 (N_16587,N_16107,N_16419);
or U16588 (N_16588,N_16426,N_16219);
nor U16589 (N_16589,N_16209,N_16200);
xor U16590 (N_16590,N_16372,N_16352);
xor U16591 (N_16591,N_16357,N_16449);
and U16592 (N_16592,N_16234,N_16343);
nor U16593 (N_16593,N_16186,N_16227);
nand U16594 (N_16594,N_16457,N_16251);
nor U16595 (N_16595,N_16225,N_16083);
or U16596 (N_16596,N_16131,N_16247);
nor U16597 (N_16597,N_16076,N_16386);
and U16598 (N_16598,N_16198,N_16296);
nand U16599 (N_16599,N_16005,N_16117);
nand U16600 (N_16600,N_16211,N_16101);
or U16601 (N_16601,N_16040,N_16244);
nand U16602 (N_16602,N_16277,N_16096);
nor U16603 (N_16603,N_16236,N_16038);
xor U16604 (N_16604,N_16303,N_16452);
nor U16605 (N_16605,N_16195,N_16375);
xnor U16606 (N_16606,N_16341,N_16399);
nand U16607 (N_16607,N_16235,N_16468);
nor U16608 (N_16608,N_16302,N_16002);
or U16609 (N_16609,N_16162,N_16060);
xnor U16610 (N_16610,N_16337,N_16260);
nor U16611 (N_16611,N_16436,N_16229);
nor U16612 (N_16612,N_16291,N_16428);
nor U16613 (N_16613,N_16307,N_16155);
or U16614 (N_16614,N_16406,N_16403);
nand U16615 (N_16615,N_16070,N_16009);
xor U16616 (N_16616,N_16472,N_16034);
nor U16617 (N_16617,N_16304,N_16336);
or U16618 (N_16618,N_16122,N_16124);
or U16619 (N_16619,N_16138,N_16394);
xnor U16620 (N_16620,N_16418,N_16057);
xor U16621 (N_16621,N_16379,N_16412);
or U16622 (N_16622,N_16362,N_16079);
or U16623 (N_16623,N_16114,N_16320);
xnor U16624 (N_16624,N_16404,N_16483);
xnor U16625 (N_16625,N_16447,N_16090);
nor U16626 (N_16626,N_16355,N_16292);
nand U16627 (N_16627,N_16154,N_16026);
or U16628 (N_16628,N_16028,N_16177);
nor U16629 (N_16629,N_16176,N_16435);
and U16630 (N_16630,N_16020,N_16230);
nor U16631 (N_16631,N_16484,N_16427);
nor U16632 (N_16632,N_16383,N_16141);
nand U16633 (N_16633,N_16212,N_16103);
nand U16634 (N_16634,N_16221,N_16316);
or U16635 (N_16635,N_16410,N_16042);
and U16636 (N_16636,N_16238,N_16193);
xor U16637 (N_16637,N_16371,N_16422);
xor U16638 (N_16638,N_16370,N_16374);
or U16639 (N_16639,N_16361,N_16494);
and U16640 (N_16640,N_16414,N_16344);
and U16641 (N_16641,N_16254,N_16423);
or U16642 (N_16642,N_16432,N_16348);
and U16643 (N_16643,N_16109,N_16071);
xor U16644 (N_16644,N_16228,N_16047);
nor U16645 (N_16645,N_16239,N_16130);
xnor U16646 (N_16646,N_16080,N_16055);
nand U16647 (N_16647,N_16334,N_16329);
or U16648 (N_16648,N_16339,N_16380);
or U16649 (N_16649,N_16074,N_16408);
xnor U16650 (N_16650,N_16210,N_16492);
xor U16651 (N_16651,N_16315,N_16147);
nor U16652 (N_16652,N_16112,N_16335);
and U16653 (N_16653,N_16312,N_16149);
nor U16654 (N_16654,N_16058,N_16360);
nand U16655 (N_16655,N_16223,N_16233);
xnor U16656 (N_16656,N_16133,N_16273);
xnor U16657 (N_16657,N_16077,N_16368);
or U16658 (N_16658,N_16395,N_16050);
nor U16659 (N_16659,N_16027,N_16243);
nand U16660 (N_16660,N_16433,N_16401);
xnor U16661 (N_16661,N_16263,N_16082);
and U16662 (N_16662,N_16279,N_16137);
xor U16663 (N_16663,N_16453,N_16487);
nand U16664 (N_16664,N_16194,N_16300);
nor U16665 (N_16665,N_16434,N_16240);
nor U16666 (N_16666,N_16000,N_16319);
and U16667 (N_16667,N_16470,N_16170);
and U16668 (N_16668,N_16166,N_16095);
nor U16669 (N_16669,N_16474,N_16032);
and U16670 (N_16670,N_16023,N_16224);
or U16671 (N_16671,N_16290,N_16087);
nor U16672 (N_16672,N_16276,N_16285);
nor U16673 (N_16673,N_16072,N_16145);
or U16674 (N_16674,N_16171,N_16275);
xnor U16675 (N_16675,N_16458,N_16293);
and U16676 (N_16676,N_16013,N_16172);
nor U16677 (N_16677,N_16010,N_16143);
xnor U16678 (N_16678,N_16473,N_16084);
nand U16679 (N_16679,N_16092,N_16465);
and U16680 (N_16680,N_16326,N_16073);
nand U16681 (N_16681,N_16309,N_16008);
nand U16682 (N_16682,N_16108,N_16393);
and U16683 (N_16683,N_16098,N_16094);
nand U16684 (N_16684,N_16356,N_16085);
nor U16685 (N_16685,N_16366,N_16086);
or U16686 (N_16686,N_16187,N_16066);
or U16687 (N_16687,N_16048,N_16359);
or U16688 (N_16688,N_16031,N_16049);
or U16689 (N_16689,N_16384,N_16462);
or U16690 (N_16690,N_16163,N_16036);
xor U16691 (N_16691,N_16283,N_16402);
or U16692 (N_16692,N_16331,N_16439);
and U16693 (N_16693,N_16232,N_16305);
xor U16694 (N_16694,N_16056,N_16338);
nand U16695 (N_16695,N_16181,N_16271);
xor U16696 (N_16696,N_16253,N_16011);
or U16697 (N_16697,N_16400,N_16129);
nor U16698 (N_16698,N_16148,N_16004);
nand U16699 (N_16699,N_16424,N_16115);
or U16700 (N_16700,N_16295,N_16286);
nand U16701 (N_16701,N_16214,N_16068);
and U16702 (N_16702,N_16469,N_16001);
or U16703 (N_16703,N_16347,N_16262);
nor U16704 (N_16704,N_16287,N_16192);
and U16705 (N_16705,N_16455,N_16201);
xnor U16706 (N_16706,N_16100,N_16180);
nor U16707 (N_16707,N_16421,N_16024);
nand U16708 (N_16708,N_16297,N_16261);
or U16709 (N_16709,N_16159,N_16353);
or U16710 (N_16710,N_16160,N_16053);
nor U16711 (N_16711,N_16306,N_16111);
and U16712 (N_16712,N_16340,N_16413);
or U16713 (N_16713,N_16226,N_16063);
nand U16714 (N_16714,N_16069,N_16161);
nand U16715 (N_16715,N_16153,N_16265);
or U16716 (N_16716,N_16025,N_16324);
and U16717 (N_16717,N_16033,N_16387);
xor U16718 (N_16718,N_16454,N_16346);
xor U16719 (N_16719,N_16451,N_16202);
xnor U16720 (N_16720,N_16120,N_16156);
nand U16721 (N_16721,N_16390,N_16416);
and U16722 (N_16722,N_16075,N_16016);
or U16723 (N_16723,N_16497,N_16358);
xnor U16724 (N_16724,N_16258,N_16065);
nor U16725 (N_16725,N_16440,N_16392);
xnor U16726 (N_16726,N_16062,N_16299);
and U16727 (N_16727,N_16325,N_16006);
and U16728 (N_16728,N_16174,N_16382);
and U16729 (N_16729,N_16169,N_16151);
and U16730 (N_16730,N_16430,N_16464);
nand U16731 (N_16731,N_16314,N_16059);
nand U16732 (N_16732,N_16365,N_16121);
and U16733 (N_16733,N_16322,N_16381);
and U16734 (N_16734,N_16052,N_16471);
nor U16735 (N_16735,N_16475,N_16488);
and U16736 (N_16736,N_16104,N_16369);
xnor U16737 (N_16737,N_16415,N_16216);
nand U16738 (N_16738,N_16021,N_16323);
nor U16739 (N_16739,N_16459,N_16281);
nor U16740 (N_16740,N_16311,N_16091);
and U16741 (N_16741,N_16248,N_16425);
nand U16742 (N_16742,N_16310,N_16215);
nand U16743 (N_16743,N_16490,N_16182);
nor U16744 (N_16744,N_16289,N_16367);
xnor U16745 (N_16745,N_16203,N_16045);
and U16746 (N_16746,N_16167,N_16191);
xnor U16747 (N_16747,N_16479,N_16259);
xor U16748 (N_16748,N_16189,N_16444);
xnor U16749 (N_16749,N_16485,N_16431);
and U16750 (N_16750,N_16455,N_16209);
xnor U16751 (N_16751,N_16283,N_16443);
or U16752 (N_16752,N_16013,N_16102);
or U16753 (N_16753,N_16104,N_16479);
nor U16754 (N_16754,N_16269,N_16238);
or U16755 (N_16755,N_16399,N_16439);
or U16756 (N_16756,N_16155,N_16408);
or U16757 (N_16757,N_16314,N_16471);
or U16758 (N_16758,N_16145,N_16370);
and U16759 (N_16759,N_16495,N_16245);
and U16760 (N_16760,N_16063,N_16003);
nor U16761 (N_16761,N_16470,N_16331);
nor U16762 (N_16762,N_16447,N_16169);
nand U16763 (N_16763,N_16021,N_16455);
or U16764 (N_16764,N_16493,N_16360);
or U16765 (N_16765,N_16380,N_16143);
and U16766 (N_16766,N_16130,N_16063);
or U16767 (N_16767,N_16129,N_16134);
xor U16768 (N_16768,N_16461,N_16176);
nor U16769 (N_16769,N_16218,N_16236);
nor U16770 (N_16770,N_16007,N_16021);
xnor U16771 (N_16771,N_16243,N_16026);
and U16772 (N_16772,N_16435,N_16051);
nand U16773 (N_16773,N_16333,N_16463);
or U16774 (N_16774,N_16061,N_16191);
xnor U16775 (N_16775,N_16412,N_16432);
and U16776 (N_16776,N_16341,N_16255);
xor U16777 (N_16777,N_16379,N_16464);
or U16778 (N_16778,N_16456,N_16013);
xor U16779 (N_16779,N_16400,N_16152);
or U16780 (N_16780,N_16401,N_16089);
xnor U16781 (N_16781,N_16222,N_16150);
and U16782 (N_16782,N_16174,N_16067);
nor U16783 (N_16783,N_16358,N_16217);
or U16784 (N_16784,N_16062,N_16287);
nor U16785 (N_16785,N_16270,N_16352);
or U16786 (N_16786,N_16487,N_16184);
or U16787 (N_16787,N_16244,N_16310);
nor U16788 (N_16788,N_16485,N_16464);
and U16789 (N_16789,N_16152,N_16328);
nand U16790 (N_16790,N_16226,N_16086);
and U16791 (N_16791,N_16145,N_16352);
and U16792 (N_16792,N_16077,N_16356);
or U16793 (N_16793,N_16326,N_16332);
nor U16794 (N_16794,N_16433,N_16327);
nand U16795 (N_16795,N_16217,N_16093);
and U16796 (N_16796,N_16267,N_16239);
and U16797 (N_16797,N_16218,N_16086);
and U16798 (N_16798,N_16059,N_16124);
nor U16799 (N_16799,N_16282,N_16374);
xnor U16800 (N_16800,N_16052,N_16483);
or U16801 (N_16801,N_16357,N_16433);
nand U16802 (N_16802,N_16021,N_16297);
and U16803 (N_16803,N_16288,N_16478);
xnor U16804 (N_16804,N_16077,N_16450);
nand U16805 (N_16805,N_16404,N_16297);
nor U16806 (N_16806,N_16195,N_16399);
or U16807 (N_16807,N_16099,N_16100);
nor U16808 (N_16808,N_16164,N_16247);
nor U16809 (N_16809,N_16487,N_16062);
nand U16810 (N_16810,N_16135,N_16252);
xor U16811 (N_16811,N_16430,N_16248);
and U16812 (N_16812,N_16073,N_16350);
nor U16813 (N_16813,N_16430,N_16145);
nand U16814 (N_16814,N_16165,N_16190);
xnor U16815 (N_16815,N_16179,N_16463);
or U16816 (N_16816,N_16231,N_16393);
nor U16817 (N_16817,N_16346,N_16085);
or U16818 (N_16818,N_16050,N_16407);
nand U16819 (N_16819,N_16316,N_16016);
xnor U16820 (N_16820,N_16158,N_16479);
nor U16821 (N_16821,N_16102,N_16299);
nand U16822 (N_16822,N_16432,N_16439);
nor U16823 (N_16823,N_16382,N_16474);
xnor U16824 (N_16824,N_16273,N_16091);
nor U16825 (N_16825,N_16045,N_16206);
or U16826 (N_16826,N_16122,N_16044);
nand U16827 (N_16827,N_16446,N_16448);
or U16828 (N_16828,N_16221,N_16023);
or U16829 (N_16829,N_16491,N_16372);
nand U16830 (N_16830,N_16305,N_16364);
and U16831 (N_16831,N_16465,N_16159);
nor U16832 (N_16832,N_16130,N_16143);
xnor U16833 (N_16833,N_16400,N_16411);
nand U16834 (N_16834,N_16196,N_16340);
nor U16835 (N_16835,N_16435,N_16402);
nand U16836 (N_16836,N_16323,N_16248);
xor U16837 (N_16837,N_16422,N_16272);
nor U16838 (N_16838,N_16198,N_16101);
or U16839 (N_16839,N_16290,N_16098);
or U16840 (N_16840,N_16082,N_16070);
xnor U16841 (N_16841,N_16301,N_16141);
nor U16842 (N_16842,N_16184,N_16190);
or U16843 (N_16843,N_16086,N_16250);
nand U16844 (N_16844,N_16068,N_16453);
xor U16845 (N_16845,N_16316,N_16333);
xor U16846 (N_16846,N_16458,N_16312);
and U16847 (N_16847,N_16030,N_16485);
nor U16848 (N_16848,N_16053,N_16280);
nand U16849 (N_16849,N_16255,N_16092);
and U16850 (N_16850,N_16480,N_16440);
or U16851 (N_16851,N_16166,N_16062);
nor U16852 (N_16852,N_16385,N_16270);
or U16853 (N_16853,N_16089,N_16480);
and U16854 (N_16854,N_16019,N_16028);
nand U16855 (N_16855,N_16182,N_16346);
or U16856 (N_16856,N_16387,N_16447);
nor U16857 (N_16857,N_16207,N_16384);
or U16858 (N_16858,N_16131,N_16473);
xor U16859 (N_16859,N_16016,N_16211);
xnor U16860 (N_16860,N_16100,N_16032);
nor U16861 (N_16861,N_16268,N_16252);
or U16862 (N_16862,N_16044,N_16289);
or U16863 (N_16863,N_16320,N_16143);
nand U16864 (N_16864,N_16074,N_16348);
xor U16865 (N_16865,N_16393,N_16308);
nor U16866 (N_16866,N_16265,N_16172);
nor U16867 (N_16867,N_16133,N_16380);
xnor U16868 (N_16868,N_16436,N_16180);
and U16869 (N_16869,N_16247,N_16188);
nand U16870 (N_16870,N_16462,N_16010);
nand U16871 (N_16871,N_16454,N_16266);
or U16872 (N_16872,N_16341,N_16425);
or U16873 (N_16873,N_16274,N_16384);
nand U16874 (N_16874,N_16224,N_16114);
and U16875 (N_16875,N_16010,N_16047);
nor U16876 (N_16876,N_16360,N_16351);
and U16877 (N_16877,N_16373,N_16284);
xor U16878 (N_16878,N_16011,N_16378);
and U16879 (N_16879,N_16049,N_16373);
nand U16880 (N_16880,N_16449,N_16298);
xor U16881 (N_16881,N_16219,N_16290);
and U16882 (N_16882,N_16450,N_16363);
nor U16883 (N_16883,N_16494,N_16451);
nor U16884 (N_16884,N_16208,N_16226);
and U16885 (N_16885,N_16196,N_16309);
nor U16886 (N_16886,N_16269,N_16186);
xor U16887 (N_16887,N_16153,N_16405);
nor U16888 (N_16888,N_16330,N_16380);
xor U16889 (N_16889,N_16478,N_16417);
xnor U16890 (N_16890,N_16306,N_16371);
and U16891 (N_16891,N_16364,N_16441);
xor U16892 (N_16892,N_16326,N_16022);
xnor U16893 (N_16893,N_16081,N_16326);
and U16894 (N_16894,N_16418,N_16101);
nor U16895 (N_16895,N_16238,N_16060);
or U16896 (N_16896,N_16053,N_16066);
nand U16897 (N_16897,N_16223,N_16456);
nand U16898 (N_16898,N_16059,N_16397);
nor U16899 (N_16899,N_16202,N_16059);
nand U16900 (N_16900,N_16488,N_16171);
nor U16901 (N_16901,N_16189,N_16256);
or U16902 (N_16902,N_16418,N_16002);
nand U16903 (N_16903,N_16266,N_16126);
nand U16904 (N_16904,N_16399,N_16334);
nand U16905 (N_16905,N_16231,N_16467);
or U16906 (N_16906,N_16382,N_16067);
xnor U16907 (N_16907,N_16064,N_16003);
xnor U16908 (N_16908,N_16432,N_16075);
and U16909 (N_16909,N_16309,N_16206);
or U16910 (N_16910,N_16277,N_16453);
nand U16911 (N_16911,N_16178,N_16117);
xnor U16912 (N_16912,N_16438,N_16116);
nor U16913 (N_16913,N_16035,N_16353);
and U16914 (N_16914,N_16389,N_16289);
xor U16915 (N_16915,N_16324,N_16131);
xor U16916 (N_16916,N_16447,N_16137);
and U16917 (N_16917,N_16399,N_16031);
or U16918 (N_16918,N_16335,N_16218);
xor U16919 (N_16919,N_16035,N_16286);
xor U16920 (N_16920,N_16202,N_16242);
nor U16921 (N_16921,N_16048,N_16357);
nor U16922 (N_16922,N_16197,N_16194);
xnor U16923 (N_16923,N_16015,N_16281);
and U16924 (N_16924,N_16437,N_16497);
or U16925 (N_16925,N_16132,N_16078);
nand U16926 (N_16926,N_16285,N_16175);
nor U16927 (N_16927,N_16135,N_16036);
nand U16928 (N_16928,N_16489,N_16233);
or U16929 (N_16929,N_16304,N_16088);
and U16930 (N_16930,N_16475,N_16378);
nand U16931 (N_16931,N_16219,N_16369);
nor U16932 (N_16932,N_16016,N_16047);
or U16933 (N_16933,N_16192,N_16478);
xnor U16934 (N_16934,N_16245,N_16066);
nand U16935 (N_16935,N_16431,N_16291);
xnor U16936 (N_16936,N_16299,N_16491);
and U16937 (N_16937,N_16192,N_16123);
nand U16938 (N_16938,N_16258,N_16262);
and U16939 (N_16939,N_16357,N_16035);
xor U16940 (N_16940,N_16131,N_16426);
or U16941 (N_16941,N_16483,N_16371);
or U16942 (N_16942,N_16066,N_16013);
xor U16943 (N_16943,N_16292,N_16412);
nand U16944 (N_16944,N_16275,N_16357);
nor U16945 (N_16945,N_16324,N_16192);
xor U16946 (N_16946,N_16217,N_16012);
nand U16947 (N_16947,N_16346,N_16172);
or U16948 (N_16948,N_16465,N_16399);
or U16949 (N_16949,N_16297,N_16181);
nand U16950 (N_16950,N_16415,N_16099);
and U16951 (N_16951,N_16122,N_16414);
nor U16952 (N_16952,N_16137,N_16060);
and U16953 (N_16953,N_16214,N_16030);
or U16954 (N_16954,N_16391,N_16482);
or U16955 (N_16955,N_16118,N_16148);
nor U16956 (N_16956,N_16271,N_16412);
nand U16957 (N_16957,N_16247,N_16379);
nor U16958 (N_16958,N_16320,N_16423);
xnor U16959 (N_16959,N_16216,N_16278);
and U16960 (N_16960,N_16076,N_16096);
or U16961 (N_16961,N_16109,N_16389);
xnor U16962 (N_16962,N_16391,N_16252);
nor U16963 (N_16963,N_16302,N_16214);
nor U16964 (N_16964,N_16413,N_16125);
nand U16965 (N_16965,N_16363,N_16037);
nor U16966 (N_16966,N_16487,N_16415);
xnor U16967 (N_16967,N_16482,N_16346);
nor U16968 (N_16968,N_16305,N_16167);
xnor U16969 (N_16969,N_16251,N_16278);
xnor U16970 (N_16970,N_16491,N_16282);
nand U16971 (N_16971,N_16462,N_16017);
xor U16972 (N_16972,N_16497,N_16251);
and U16973 (N_16973,N_16365,N_16024);
nand U16974 (N_16974,N_16332,N_16469);
or U16975 (N_16975,N_16019,N_16149);
or U16976 (N_16976,N_16133,N_16004);
nand U16977 (N_16977,N_16406,N_16371);
nand U16978 (N_16978,N_16175,N_16282);
xnor U16979 (N_16979,N_16143,N_16276);
and U16980 (N_16980,N_16115,N_16179);
and U16981 (N_16981,N_16282,N_16268);
xor U16982 (N_16982,N_16013,N_16393);
or U16983 (N_16983,N_16003,N_16362);
nor U16984 (N_16984,N_16214,N_16358);
and U16985 (N_16985,N_16158,N_16181);
xnor U16986 (N_16986,N_16158,N_16125);
nor U16987 (N_16987,N_16308,N_16086);
nor U16988 (N_16988,N_16367,N_16196);
or U16989 (N_16989,N_16273,N_16274);
nor U16990 (N_16990,N_16237,N_16197);
nand U16991 (N_16991,N_16256,N_16460);
or U16992 (N_16992,N_16442,N_16418);
nor U16993 (N_16993,N_16310,N_16063);
nand U16994 (N_16994,N_16344,N_16431);
and U16995 (N_16995,N_16121,N_16122);
nor U16996 (N_16996,N_16308,N_16101);
and U16997 (N_16997,N_16497,N_16427);
and U16998 (N_16998,N_16401,N_16338);
nor U16999 (N_16999,N_16168,N_16390);
nor U17000 (N_17000,N_16972,N_16635);
and U17001 (N_17001,N_16747,N_16612);
or U17002 (N_17002,N_16620,N_16576);
and U17003 (N_17003,N_16994,N_16896);
and U17004 (N_17004,N_16753,N_16586);
nor U17005 (N_17005,N_16939,N_16502);
xor U17006 (N_17006,N_16998,N_16530);
or U17007 (N_17007,N_16901,N_16834);
xor U17008 (N_17008,N_16552,N_16568);
nor U17009 (N_17009,N_16599,N_16903);
and U17010 (N_17010,N_16566,N_16942);
nor U17011 (N_17011,N_16973,N_16557);
nand U17012 (N_17012,N_16583,N_16917);
nor U17013 (N_17013,N_16625,N_16543);
or U17014 (N_17014,N_16914,N_16816);
xnor U17015 (N_17015,N_16936,N_16899);
or U17016 (N_17016,N_16758,N_16760);
nor U17017 (N_17017,N_16825,N_16590);
xor U17018 (N_17018,N_16797,N_16793);
and U17019 (N_17019,N_16822,N_16680);
and U17020 (N_17020,N_16713,N_16648);
or U17021 (N_17021,N_16556,N_16892);
or U17022 (N_17022,N_16943,N_16869);
nand U17023 (N_17023,N_16545,N_16640);
or U17024 (N_17024,N_16655,N_16656);
and U17025 (N_17025,N_16961,N_16958);
nand U17026 (N_17026,N_16909,N_16670);
nand U17027 (N_17027,N_16720,N_16513);
xnor U17028 (N_17028,N_16875,N_16742);
nor U17029 (N_17029,N_16796,N_16995);
and U17030 (N_17030,N_16887,N_16633);
xor U17031 (N_17031,N_16947,N_16759);
nor U17032 (N_17032,N_16578,N_16592);
or U17033 (N_17033,N_16630,N_16567);
nand U17034 (N_17034,N_16750,N_16559);
or U17035 (N_17035,N_16831,N_16639);
xor U17036 (N_17036,N_16649,N_16919);
and U17037 (N_17037,N_16980,N_16621);
nor U17038 (N_17038,N_16951,N_16724);
or U17039 (N_17039,N_16996,N_16575);
or U17040 (N_17040,N_16697,N_16693);
nor U17041 (N_17041,N_16833,N_16626);
xnor U17042 (N_17042,N_16631,N_16835);
and U17043 (N_17043,N_16827,N_16546);
and U17044 (N_17044,N_16595,N_16930);
or U17045 (N_17045,N_16520,N_16946);
and U17046 (N_17046,N_16969,N_16673);
and U17047 (N_17047,N_16940,N_16739);
or U17048 (N_17048,N_16527,N_16982);
xnor U17049 (N_17049,N_16554,N_16840);
and U17050 (N_17050,N_16651,N_16810);
and U17051 (N_17051,N_16800,N_16910);
xor U17052 (N_17052,N_16855,N_16676);
nor U17053 (N_17053,N_16574,N_16868);
xor U17054 (N_17054,N_16560,N_16859);
xnor U17055 (N_17055,N_16820,N_16732);
or U17056 (N_17056,N_16518,N_16853);
nand U17057 (N_17057,N_16591,N_16521);
and U17058 (N_17058,N_16778,N_16911);
nand U17059 (N_17059,N_16999,N_16522);
xor U17060 (N_17060,N_16788,N_16532);
nor U17061 (N_17061,N_16811,N_16614);
and U17062 (N_17062,N_16769,N_16873);
nor U17063 (N_17063,N_16849,N_16658);
and U17064 (N_17064,N_16741,N_16846);
nor U17065 (N_17065,N_16832,N_16815);
or U17066 (N_17066,N_16550,N_16765);
nor U17067 (N_17067,N_16891,N_16989);
nand U17068 (N_17068,N_16681,N_16852);
xor U17069 (N_17069,N_16971,N_16689);
or U17070 (N_17070,N_16781,N_16701);
xnor U17071 (N_17071,N_16871,N_16627);
xnor U17072 (N_17072,N_16606,N_16885);
or U17073 (N_17073,N_16642,N_16959);
xor U17074 (N_17074,N_16782,N_16510);
or U17075 (N_17075,N_16728,N_16636);
xor U17076 (N_17076,N_16812,N_16506);
or U17077 (N_17077,N_16691,N_16861);
xnor U17078 (N_17078,N_16838,N_16955);
xor U17079 (N_17079,N_16582,N_16533);
nor U17080 (N_17080,N_16704,N_16682);
nand U17081 (N_17081,N_16945,N_16604);
and U17082 (N_17082,N_16824,N_16783);
and U17083 (N_17083,N_16924,N_16524);
nand U17084 (N_17084,N_16927,N_16949);
nor U17085 (N_17085,N_16798,N_16751);
or U17086 (N_17086,N_16746,N_16572);
and U17087 (N_17087,N_16744,N_16601);
nand U17088 (N_17088,N_16699,N_16990);
xor U17089 (N_17089,N_16770,N_16664);
or U17090 (N_17090,N_16893,N_16826);
xor U17091 (N_17091,N_16652,N_16843);
nor U17092 (N_17092,N_16929,N_16860);
nor U17093 (N_17093,N_16986,N_16774);
nand U17094 (N_17094,N_16613,N_16677);
xor U17095 (N_17095,N_16886,N_16987);
nand U17096 (N_17096,N_16856,N_16779);
nand U17097 (N_17097,N_16617,N_16503);
or U17098 (N_17098,N_16702,N_16684);
nor U17099 (N_17099,N_16611,N_16794);
and U17100 (N_17100,N_16596,N_16512);
and U17101 (N_17101,N_16628,N_16666);
and U17102 (N_17102,N_16675,N_16763);
nand U17103 (N_17103,N_16694,N_16555);
nor U17104 (N_17104,N_16637,N_16509);
nand U17105 (N_17105,N_16967,N_16938);
xor U17106 (N_17106,N_16952,N_16890);
nor U17107 (N_17107,N_16823,N_16773);
xor U17108 (N_17108,N_16711,N_16933);
and U17109 (N_17109,N_16979,N_16937);
or U17110 (N_17110,N_16602,N_16618);
xnor U17111 (N_17111,N_16957,N_16950);
nand U17112 (N_17112,N_16733,N_16997);
or U17113 (N_17113,N_16535,N_16841);
xor U17114 (N_17114,N_16641,N_16553);
and U17115 (N_17115,N_16603,N_16531);
xor U17116 (N_17116,N_16516,N_16716);
or U17117 (N_17117,N_16809,N_16818);
nand U17118 (N_17118,N_16683,N_16696);
nand U17119 (N_17119,N_16692,N_16771);
nand U17120 (N_17120,N_16705,N_16507);
nor U17121 (N_17121,N_16948,N_16668);
nand U17122 (N_17122,N_16643,N_16548);
and U17123 (N_17123,N_16784,N_16964);
xnor U17124 (N_17124,N_16821,N_16610);
or U17125 (N_17125,N_16888,N_16738);
and U17126 (N_17126,N_16991,N_16593);
nor U17127 (N_17127,N_16736,N_16844);
nor U17128 (N_17128,N_16864,N_16953);
xnor U17129 (N_17129,N_16845,N_16926);
and U17130 (N_17130,N_16906,N_16881);
nor U17131 (N_17131,N_16672,N_16928);
xor U17132 (N_17132,N_16857,N_16992);
nor U17133 (N_17133,N_16983,N_16544);
nor U17134 (N_17134,N_16504,N_16828);
nand U17135 (N_17135,N_16536,N_16565);
nand U17136 (N_17136,N_16904,N_16632);
and U17137 (N_17137,N_16538,N_16570);
nand U17138 (N_17138,N_16540,N_16839);
or U17139 (N_17139,N_16922,N_16710);
nor U17140 (N_17140,N_16975,N_16665);
xor U17141 (N_17141,N_16638,N_16960);
or U17142 (N_17142,N_16976,N_16663);
xnor U17143 (N_17143,N_16646,N_16659);
xnor U17144 (N_17144,N_16785,N_16525);
or U17145 (N_17145,N_16848,N_16594);
nor U17146 (N_17146,N_16740,N_16584);
or U17147 (N_17147,N_16805,N_16787);
nand U17148 (N_17148,N_16863,N_16837);
nor U17149 (N_17149,N_16882,N_16842);
nor U17150 (N_17150,N_16645,N_16598);
nor U17151 (N_17151,N_16597,N_16970);
xor U17152 (N_17152,N_16789,N_16768);
nor U17153 (N_17153,N_16915,N_16709);
or U17154 (N_17154,N_16907,N_16752);
xnor U17155 (N_17155,N_16718,N_16714);
nand U17156 (N_17156,N_16647,N_16687);
xor U17157 (N_17157,N_16977,N_16808);
or U17158 (N_17158,N_16847,N_16726);
and U17159 (N_17159,N_16619,N_16529);
xor U17160 (N_17160,N_16748,N_16993);
xor U17161 (N_17161,N_16854,N_16913);
or U17162 (N_17162,N_16622,N_16708);
or U17163 (N_17163,N_16690,N_16581);
and U17164 (N_17164,N_16962,N_16674);
or U17165 (N_17165,N_16577,N_16703);
or U17166 (N_17166,N_16608,N_16902);
or U17167 (N_17167,N_16877,N_16660);
nor U17168 (N_17168,N_16561,N_16934);
or U17169 (N_17169,N_16981,N_16700);
and U17170 (N_17170,N_16829,N_16539);
and U17171 (N_17171,N_16984,N_16884);
and U17172 (N_17172,N_16925,N_16722);
nand U17173 (N_17173,N_16735,N_16935);
nor U17174 (N_17174,N_16657,N_16978);
xnor U17175 (N_17175,N_16806,N_16894);
xor U17176 (N_17176,N_16897,N_16900);
and U17177 (N_17177,N_16776,N_16571);
nor U17178 (N_17178,N_16721,N_16616);
and U17179 (N_17179,N_16623,N_16505);
and U17180 (N_17180,N_16819,N_16688);
and U17181 (N_17181,N_16764,N_16923);
and U17182 (N_17182,N_16790,N_16745);
and U17183 (N_17183,N_16558,N_16653);
and U17184 (N_17184,N_16932,N_16795);
xnor U17185 (N_17185,N_16500,N_16755);
nor U17186 (N_17186,N_16523,N_16879);
nand U17187 (N_17187,N_16654,N_16850);
nand U17188 (N_17188,N_16876,N_16916);
nand U17189 (N_17189,N_16836,N_16729);
nand U17190 (N_17190,N_16830,N_16944);
xor U17191 (N_17191,N_16920,N_16537);
nor U17192 (N_17192,N_16685,N_16956);
or U17193 (N_17193,N_16813,N_16579);
nand U17194 (N_17194,N_16707,N_16589);
nand U17195 (N_17195,N_16580,N_16526);
nor U17196 (N_17196,N_16667,N_16965);
nor U17197 (N_17197,N_16588,N_16501);
and U17198 (N_17198,N_16547,N_16511);
xor U17199 (N_17199,N_16791,N_16817);
and U17200 (N_17200,N_16731,N_16851);
nand U17201 (N_17201,N_16880,N_16931);
nor U17202 (N_17202,N_16889,N_16609);
nor U17203 (N_17203,N_16629,N_16650);
nand U17204 (N_17204,N_16534,N_16968);
and U17205 (N_17205,N_16767,N_16662);
and U17206 (N_17206,N_16905,N_16802);
or U17207 (N_17207,N_16883,N_16743);
and U17208 (N_17208,N_16585,N_16727);
xnor U17209 (N_17209,N_16562,N_16814);
and U17210 (N_17210,N_16941,N_16730);
and U17211 (N_17211,N_16870,N_16587);
xnor U17212 (N_17212,N_16807,N_16573);
or U17213 (N_17213,N_16723,N_16563);
nand U17214 (N_17214,N_16803,N_16754);
nand U17215 (N_17215,N_16719,N_16706);
or U17216 (N_17216,N_16514,N_16963);
nor U17217 (N_17217,N_16799,N_16717);
nand U17218 (N_17218,N_16908,N_16974);
nand U17219 (N_17219,N_16715,N_16615);
xor U17220 (N_17220,N_16569,N_16761);
xnor U17221 (N_17221,N_16508,N_16686);
xor U17222 (N_17222,N_16872,N_16867);
nand U17223 (N_17223,N_16985,N_16866);
and U17224 (N_17224,N_16762,N_16862);
xor U17225 (N_17225,N_16634,N_16772);
and U17226 (N_17226,N_16749,N_16541);
or U17227 (N_17227,N_16600,N_16712);
nand U17228 (N_17228,N_16766,N_16542);
nand U17229 (N_17229,N_16858,N_16780);
nor U17230 (N_17230,N_16517,N_16644);
and U17231 (N_17231,N_16605,N_16988);
nor U17232 (N_17232,N_16912,N_16698);
and U17233 (N_17233,N_16624,N_16695);
nand U17234 (N_17234,N_16756,N_16878);
nand U17235 (N_17235,N_16669,N_16757);
or U17236 (N_17236,N_16725,N_16804);
xor U17237 (N_17237,N_16564,N_16865);
nor U17238 (N_17238,N_16519,N_16918);
nand U17239 (N_17239,N_16777,N_16898);
nand U17240 (N_17240,N_16679,N_16528);
and U17241 (N_17241,N_16874,N_16954);
and U17242 (N_17242,N_16734,N_16671);
nor U17243 (N_17243,N_16966,N_16678);
xnor U17244 (N_17244,N_16551,N_16786);
nor U17245 (N_17245,N_16921,N_16661);
nor U17246 (N_17246,N_16895,N_16801);
nor U17247 (N_17247,N_16737,N_16775);
and U17248 (N_17248,N_16792,N_16515);
or U17249 (N_17249,N_16549,N_16607);
nand U17250 (N_17250,N_16940,N_16612);
nand U17251 (N_17251,N_16824,N_16996);
or U17252 (N_17252,N_16616,N_16689);
nand U17253 (N_17253,N_16602,N_16697);
nor U17254 (N_17254,N_16925,N_16817);
or U17255 (N_17255,N_16682,N_16864);
nor U17256 (N_17256,N_16504,N_16509);
nor U17257 (N_17257,N_16744,N_16874);
nand U17258 (N_17258,N_16958,N_16980);
nor U17259 (N_17259,N_16798,N_16940);
xor U17260 (N_17260,N_16831,N_16882);
xnor U17261 (N_17261,N_16557,N_16925);
xnor U17262 (N_17262,N_16763,N_16700);
or U17263 (N_17263,N_16582,N_16792);
nand U17264 (N_17264,N_16744,N_16938);
and U17265 (N_17265,N_16822,N_16718);
xnor U17266 (N_17266,N_16895,N_16766);
or U17267 (N_17267,N_16736,N_16878);
nand U17268 (N_17268,N_16766,N_16528);
or U17269 (N_17269,N_16592,N_16768);
nand U17270 (N_17270,N_16876,N_16697);
xnor U17271 (N_17271,N_16845,N_16847);
nand U17272 (N_17272,N_16636,N_16552);
nand U17273 (N_17273,N_16859,N_16773);
and U17274 (N_17274,N_16957,N_16951);
and U17275 (N_17275,N_16563,N_16916);
nor U17276 (N_17276,N_16765,N_16746);
nand U17277 (N_17277,N_16756,N_16560);
or U17278 (N_17278,N_16663,N_16813);
nor U17279 (N_17279,N_16674,N_16861);
xor U17280 (N_17280,N_16637,N_16706);
and U17281 (N_17281,N_16925,N_16769);
nor U17282 (N_17282,N_16625,N_16929);
nand U17283 (N_17283,N_16504,N_16740);
and U17284 (N_17284,N_16897,N_16940);
or U17285 (N_17285,N_16654,N_16591);
or U17286 (N_17286,N_16719,N_16677);
and U17287 (N_17287,N_16587,N_16781);
xnor U17288 (N_17288,N_16707,N_16799);
xnor U17289 (N_17289,N_16793,N_16788);
or U17290 (N_17290,N_16903,N_16790);
nor U17291 (N_17291,N_16624,N_16963);
and U17292 (N_17292,N_16949,N_16776);
nor U17293 (N_17293,N_16856,N_16928);
and U17294 (N_17294,N_16614,N_16503);
xnor U17295 (N_17295,N_16718,N_16563);
and U17296 (N_17296,N_16863,N_16711);
nand U17297 (N_17297,N_16822,N_16559);
nor U17298 (N_17298,N_16823,N_16850);
nand U17299 (N_17299,N_16506,N_16986);
xor U17300 (N_17300,N_16774,N_16753);
nand U17301 (N_17301,N_16896,N_16883);
nand U17302 (N_17302,N_16940,N_16729);
or U17303 (N_17303,N_16648,N_16996);
and U17304 (N_17304,N_16649,N_16758);
or U17305 (N_17305,N_16810,N_16694);
and U17306 (N_17306,N_16602,N_16976);
or U17307 (N_17307,N_16981,N_16592);
and U17308 (N_17308,N_16924,N_16666);
or U17309 (N_17309,N_16633,N_16551);
nor U17310 (N_17310,N_16668,N_16653);
and U17311 (N_17311,N_16668,N_16684);
or U17312 (N_17312,N_16502,N_16696);
and U17313 (N_17313,N_16965,N_16572);
xnor U17314 (N_17314,N_16726,N_16971);
and U17315 (N_17315,N_16515,N_16890);
or U17316 (N_17316,N_16909,N_16644);
and U17317 (N_17317,N_16731,N_16852);
xnor U17318 (N_17318,N_16595,N_16695);
xor U17319 (N_17319,N_16691,N_16675);
nor U17320 (N_17320,N_16589,N_16961);
nand U17321 (N_17321,N_16679,N_16601);
and U17322 (N_17322,N_16707,N_16621);
nand U17323 (N_17323,N_16895,N_16901);
and U17324 (N_17324,N_16577,N_16529);
xor U17325 (N_17325,N_16951,N_16520);
nor U17326 (N_17326,N_16644,N_16940);
xor U17327 (N_17327,N_16600,N_16532);
or U17328 (N_17328,N_16911,N_16843);
nor U17329 (N_17329,N_16975,N_16607);
and U17330 (N_17330,N_16809,N_16869);
nand U17331 (N_17331,N_16885,N_16707);
xnor U17332 (N_17332,N_16661,N_16892);
and U17333 (N_17333,N_16604,N_16977);
and U17334 (N_17334,N_16894,N_16606);
nand U17335 (N_17335,N_16835,N_16770);
nor U17336 (N_17336,N_16880,N_16970);
xnor U17337 (N_17337,N_16531,N_16726);
xnor U17338 (N_17338,N_16539,N_16584);
nand U17339 (N_17339,N_16930,N_16547);
nand U17340 (N_17340,N_16500,N_16925);
xor U17341 (N_17341,N_16594,N_16931);
and U17342 (N_17342,N_16712,N_16791);
nand U17343 (N_17343,N_16808,N_16773);
nand U17344 (N_17344,N_16823,N_16752);
and U17345 (N_17345,N_16695,N_16849);
and U17346 (N_17346,N_16915,N_16962);
or U17347 (N_17347,N_16519,N_16864);
and U17348 (N_17348,N_16593,N_16871);
or U17349 (N_17349,N_16591,N_16833);
xor U17350 (N_17350,N_16575,N_16603);
nor U17351 (N_17351,N_16714,N_16697);
nor U17352 (N_17352,N_16674,N_16867);
and U17353 (N_17353,N_16951,N_16778);
nor U17354 (N_17354,N_16981,N_16699);
nor U17355 (N_17355,N_16656,N_16661);
or U17356 (N_17356,N_16921,N_16822);
nand U17357 (N_17357,N_16925,N_16551);
nand U17358 (N_17358,N_16841,N_16563);
or U17359 (N_17359,N_16885,N_16991);
or U17360 (N_17360,N_16643,N_16768);
nor U17361 (N_17361,N_16906,N_16915);
nor U17362 (N_17362,N_16529,N_16763);
xor U17363 (N_17363,N_16567,N_16676);
nand U17364 (N_17364,N_16901,N_16832);
nand U17365 (N_17365,N_16690,N_16687);
nor U17366 (N_17366,N_16732,N_16990);
xnor U17367 (N_17367,N_16796,N_16915);
and U17368 (N_17368,N_16905,N_16714);
or U17369 (N_17369,N_16537,N_16963);
nand U17370 (N_17370,N_16928,N_16764);
xor U17371 (N_17371,N_16670,N_16680);
or U17372 (N_17372,N_16783,N_16815);
and U17373 (N_17373,N_16916,N_16724);
xnor U17374 (N_17374,N_16991,N_16612);
nor U17375 (N_17375,N_16961,N_16842);
nand U17376 (N_17376,N_16602,N_16656);
and U17377 (N_17377,N_16681,N_16577);
xor U17378 (N_17378,N_16611,N_16754);
or U17379 (N_17379,N_16861,N_16781);
or U17380 (N_17380,N_16991,N_16674);
and U17381 (N_17381,N_16795,N_16555);
nor U17382 (N_17382,N_16795,N_16561);
xnor U17383 (N_17383,N_16999,N_16821);
nor U17384 (N_17384,N_16945,N_16958);
nand U17385 (N_17385,N_16944,N_16573);
nand U17386 (N_17386,N_16586,N_16758);
nor U17387 (N_17387,N_16698,N_16768);
nor U17388 (N_17388,N_16983,N_16529);
xnor U17389 (N_17389,N_16920,N_16612);
or U17390 (N_17390,N_16730,N_16731);
xor U17391 (N_17391,N_16784,N_16688);
nor U17392 (N_17392,N_16779,N_16626);
nor U17393 (N_17393,N_16998,N_16758);
nand U17394 (N_17394,N_16938,N_16949);
nand U17395 (N_17395,N_16817,N_16524);
xor U17396 (N_17396,N_16553,N_16846);
and U17397 (N_17397,N_16946,N_16916);
or U17398 (N_17398,N_16892,N_16890);
nor U17399 (N_17399,N_16936,N_16793);
xor U17400 (N_17400,N_16656,N_16688);
nor U17401 (N_17401,N_16639,N_16961);
nor U17402 (N_17402,N_16598,N_16623);
and U17403 (N_17403,N_16849,N_16833);
nand U17404 (N_17404,N_16960,N_16762);
or U17405 (N_17405,N_16672,N_16894);
nand U17406 (N_17406,N_16967,N_16668);
or U17407 (N_17407,N_16683,N_16750);
nand U17408 (N_17408,N_16880,N_16500);
or U17409 (N_17409,N_16680,N_16903);
nor U17410 (N_17410,N_16814,N_16763);
xor U17411 (N_17411,N_16729,N_16726);
xor U17412 (N_17412,N_16788,N_16770);
xor U17413 (N_17413,N_16863,N_16654);
nand U17414 (N_17414,N_16746,N_16699);
xnor U17415 (N_17415,N_16820,N_16652);
nand U17416 (N_17416,N_16926,N_16978);
nand U17417 (N_17417,N_16774,N_16865);
nor U17418 (N_17418,N_16604,N_16554);
or U17419 (N_17419,N_16821,N_16514);
nor U17420 (N_17420,N_16678,N_16794);
and U17421 (N_17421,N_16989,N_16773);
and U17422 (N_17422,N_16680,N_16725);
xnor U17423 (N_17423,N_16915,N_16775);
or U17424 (N_17424,N_16886,N_16671);
nand U17425 (N_17425,N_16680,N_16840);
and U17426 (N_17426,N_16671,N_16733);
and U17427 (N_17427,N_16735,N_16545);
nor U17428 (N_17428,N_16945,N_16541);
nor U17429 (N_17429,N_16715,N_16548);
xor U17430 (N_17430,N_16733,N_16969);
and U17431 (N_17431,N_16787,N_16963);
or U17432 (N_17432,N_16724,N_16878);
xnor U17433 (N_17433,N_16934,N_16985);
and U17434 (N_17434,N_16806,N_16760);
and U17435 (N_17435,N_16582,N_16679);
or U17436 (N_17436,N_16881,N_16789);
and U17437 (N_17437,N_16817,N_16802);
nor U17438 (N_17438,N_16781,N_16726);
and U17439 (N_17439,N_16922,N_16927);
or U17440 (N_17440,N_16798,N_16807);
and U17441 (N_17441,N_16582,N_16794);
or U17442 (N_17442,N_16642,N_16540);
nand U17443 (N_17443,N_16764,N_16983);
nand U17444 (N_17444,N_16591,N_16829);
nand U17445 (N_17445,N_16870,N_16524);
nor U17446 (N_17446,N_16822,N_16672);
or U17447 (N_17447,N_16896,N_16625);
nand U17448 (N_17448,N_16655,N_16819);
nand U17449 (N_17449,N_16603,N_16795);
xnor U17450 (N_17450,N_16799,N_16665);
and U17451 (N_17451,N_16571,N_16786);
or U17452 (N_17452,N_16940,N_16971);
nor U17453 (N_17453,N_16897,N_16808);
xnor U17454 (N_17454,N_16957,N_16706);
xor U17455 (N_17455,N_16606,N_16846);
nand U17456 (N_17456,N_16654,N_16707);
or U17457 (N_17457,N_16764,N_16575);
or U17458 (N_17458,N_16607,N_16588);
nor U17459 (N_17459,N_16506,N_16531);
or U17460 (N_17460,N_16564,N_16639);
nand U17461 (N_17461,N_16670,N_16544);
xor U17462 (N_17462,N_16917,N_16829);
and U17463 (N_17463,N_16764,N_16657);
xnor U17464 (N_17464,N_16589,N_16653);
nand U17465 (N_17465,N_16574,N_16505);
xor U17466 (N_17466,N_16583,N_16688);
nor U17467 (N_17467,N_16839,N_16529);
nor U17468 (N_17468,N_16549,N_16963);
nand U17469 (N_17469,N_16902,N_16690);
and U17470 (N_17470,N_16928,N_16951);
or U17471 (N_17471,N_16946,N_16815);
nor U17472 (N_17472,N_16761,N_16966);
and U17473 (N_17473,N_16801,N_16949);
nand U17474 (N_17474,N_16643,N_16786);
nand U17475 (N_17475,N_16602,N_16971);
and U17476 (N_17476,N_16794,N_16997);
nor U17477 (N_17477,N_16589,N_16698);
xnor U17478 (N_17478,N_16995,N_16562);
and U17479 (N_17479,N_16899,N_16877);
nor U17480 (N_17480,N_16698,N_16717);
xnor U17481 (N_17481,N_16774,N_16567);
and U17482 (N_17482,N_16549,N_16746);
nand U17483 (N_17483,N_16841,N_16559);
and U17484 (N_17484,N_16666,N_16993);
nand U17485 (N_17485,N_16772,N_16665);
and U17486 (N_17486,N_16951,N_16642);
xor U17487 (N_17487,N_16605,N_16832);
nand U17488 (N_17488,N_16949,N_16538);
and U17489 (N_17489,N_16523,N_16581);
nand U17490 (N_17490,N_16712,N_16547);
nand U17491 (N_17491,N_16626,N_16879);
nor U17492 (N_17492,N_16778,N_16570);
nor U17493 (N_17493,N_16563,N_16741);
nor U17494 (N_17494,N_16937,N_16588);
or U17495 (N_17495,N_16969,N_16757);
nor U17496 (N_17496,N_16573,N_16644);
and U17497 (N_17497,N_16543,N_16706);
and U17498 (N_17498,N_16705,N_16864);
nand U17499 (N_17499,N_16604,N_16886);
xor U17500 (N_17500,N_17441,N_17200);
or U17501 (N_17501,N_17078,N_17053);
or U17502 (N_17502,N_17120,N_17329);
nor U17503 (N_17503,N_17280,N_17307);
xor U17504 (N_17504,N_17143,N_17133);
xnor U17505 (N_17505,N_17251,N_17389);
nor U17506 (N_17506,N_17434,N_17195);
and U17507 (N_17507,N_17080,N_17141);
and U17508 (N_17508,N_17085,N_17221);
or U17509 (N_17509,N_17289,N_17225);
xor U17510 (N_17510,N_17153,N_17127);
nor U17511 (N_17511,N_17247,N_17360);
or U17512 (N_17512,N_17048,N_17325);
nor U17513 (N_17513,N_17458,N_17284);
xor U17514 (N_17514,N_17437,N_17430);
or U17515 (N_17515,N_17366,N_17173);
nor U17516 (N_17516,N_17497,N_17056);
nand U17517 (N_17517,N_17040,N_17345);
or U17518 (N_17518,N_17298,N_17005);
or U17519 (N_17519,N_17213,N_17115);
xor U17520 (N_17520,N_17044,N_17445);
and U17521 (N_17521,N_17217,N_17494);
and U17522 (N_17522,N_17318,N_17302);
xnor U17523 (N_17523,N_17015,N_17493);
xor U17524 (N_17524,N_17238,N_17268);
nor U17525 (N_17525,N_17065,N_17347);
and U17526 (N_17526,N_17062,N_17265);
and U17527 (N_17527,N_17147,N_17435);
or U17528 (N_17528,N_17266,N_17034);
nor U17529 (N_17529,N_17379,N_17261);
or U17530 (N_17530,N_17113,N_17449);
nor U17531 (N_17531,N_17296,N_17183);
xor U17532 (N_17532,N_17042,N_17267);
nor U17533 (N_17533,N_17477,N_17020);
or U17534 (N_17534,N_17124,N_17371);
nor U17535 (N_17535,N_17125,N_17241);
xnor U17536 (N_17536,N_17287,N_17237);
nand U17537 (N_17537,N_17285,N_17220);
or U17538 (N_17538,N_17337,N_17310);
nor U17539 (N_17539,N_17073,N_17013);
xnor U17540 (N_17540,N_17414,N_17180);
and U17541 (N_17541,N_17372,N_17172);
nor U17542 (N_17542,N_17390,N_17304);
nor U17543 (N_17543,N_17242,N_17384);
or U17544 (N_17544,N_17194,N_17232);
nor U17545 (N_17545,N_17017,N_17111);
xor U17546 (N_17546,N_17160,N_17109);
nand U17547 (N_17547,N_17166,N_17264);
nand U17548 (N_17548,N_17161,N_17159);
nand U17549 (N_17549,N_17218,N_17203);
nor U17550 (N_17550,N_17002,N_17433);
xnor U17551 (N_17551,N_17416,N_17359);
or U17552 (N_17552,N_17239,N_17275);
nor U17553 (N_17553,N_17076,N_17401);
nand U17554 (N_17554,N_17156,N_17398);
xnor U17555 (N_17555,N_17228,N_17474);
nand U17556 (N_17556,N_17061,N_17370);
nor U17557 (N_17557,N_17152,N_17394);
nand U17558 (N_17558,N_17096,N_17427);
nor U17559 (N_17559,N_17052,N_17186);
nor U17560 (N_17560,N_17019,N_17462);
nand U17561 (N_17561,N_17098,N_17381);
xnor U17562 (N_17562,N_17240,N_17171);
nand U17563 (N_17563,N_17103,N_17229);
xor U17564 (N_17564,N_17272,N_17444);
xnor U17565 (N_17565,N_17431,N_17460);
nor U17566 (N_17566,N_17352,N_17206);
nor U17567 (N_17567,N_17039,N_17349);
nor U17568 (N_17568,N_17475,N_17350);
xor U17569 (N_17569,N_17047,N_17255);
and U17570 (N_17570,N_17059,N_17361);
and U17571 (N_17571,N_17105,N_17404);
nand U17572 (N_17572,N_17138,N_17313);
and U17573 (N_17573,N_17421,N_17029);
or U17574 (N_17574,N_17465,N_17169);
xnor U17575 (N_17575,N_17295,N_17305);
nor U17576 (N_17576,N_17190,N_17234);
nand U17577 (N_17577,N_17248,N_17198);
or U17578 (N_17578,N_17151,N_17091);
nand U17579 (N_17579,N_17193,N_17342);
and U17580 (N_17580,N_17426,N_17452);
nor U17581 (N_17581,N_17354,N_17069);
nand U17582 (N_17582,N_17294,N_17094);
or U17583 (N_17583,N_17009,N_17252);
or U17584 (N_17584,N_17417,N_17231);
xnor U17585 (N_17585,N_17301,N_17227);
or U17586 (N_17586,N_17425,N_17388);
or U17587 (N_17587,N_17300,N_17283);
and U17588 (N_17588,N_17461,N_17451);
xor U17589 (N_17589,N_17333,N_17413);
nand U17590 (N_17590,N_17204,N_17386);
xnor U17591 (N_17591,N_17101,N_17216);
nand U17592 (N_17592,N_17438,N_17378);
and U17593 (N_17593,N_17000,N_17025);
nor U17594 (N_17594,N_17468,N_17167);
nand U17595 (N_17595,N_17402,N_17050);
and U17596 (N_17596,N_17224,N_17214);
nor U17597 (N_17597,N_17212,N_17112);
and U17598 (N_17598,N_17117,N_17336);
and U17599 (N_17599,N_17079,N_17100);
or U17600 (N_17600,N_17170,N_17409);
and U17601 (N_17601,N_17095,N_17419);
nor U17602 (N_17602,N_17396,N_17145);
and U17603 (N_17603,N_17055,N_17373);
xnor U17604 (N_17604,N_17415,N_17297);
and U17605 (N_17605,N_17278,N_17230);
nand U17606 (N_17606,N_17358,N_17154);
nor U17607 (N_17607,N_17142,N_17012);
nor U17608 (N_17608,N_17243,N_17448);
xor U17609 (N_17609,N_17439,N_17330);
nor U17610 (N_17610,N_17008,N_17057);
nor U17611 (N_17611,N_17024,N_17033);
nor U17612 (N_17612,N_17406,N_17092);
and U17613 (N_17613,N_17312,N_17383);
xor U17614 (N_17614,N_17067,N_17498);
xnor U17615 (N_17615,N_17339,N_17487);
nand U17616 (N_17616,N_17410,N_17060);
or U17617 (N_17617,N_17321,N_17282);
nand U17618 (N_17618,N_17269,N_17471);
or U17619 (N_17619,N_17028,N_17355);
nand U17620 (N_17620,N_17082,N_17382);
and U17621 (N_17621,N_17496,N_17089);
or U17622 (N_17622,N_17162,N_17420);
xor U17623 (N_17623,N_17031,N_17139);
and U17624 (N_17624,N_17215,N_17326);
xor U17625 (N_17625,N_17070,N_17236);
nor U17626 (N_17626,N_17107,N_17185);
and U17627 (N_17627,N_17357,N_17293);
nor U17628 (N_17628,N_17341,N_17041);
or U17629 (N_17629,N_17314,N_17130);
and U17630 (N_17630,N_17155,N_17385);
nor U17631 (N_17631,N_17469,N_17126);
nand U17632 (N_17632,N_17208,N_17322);
and U17633 (N_17633,N_17118,N_17442);
or U17634 (N_17634,N_17363,N_17397);
xor U17635 (N_17635,N_17472,N_17188);
or U17636 (N_17636,N_17158,N_17483);
xnor U17637 (N_17637,N_17090,N_17174);
or U17638 (N_17638,N_17099,N_17270);
xor U17639 (N_17639,N_17340,N_17026);
nor U17640 (N_17640,N_17271,N_17018);
and U17641 (N_17641,N_17315,N_17233);
or U17642 (N_17642,N_17068,N_17257);
and U17643 (N_17643,N_17088,N_17184);
nand U17644 (N_17644,N_17351,N_17299);
and U17645 (N_17645,N_17467,N_17146);
and U17646 (N_17646,N_17258,N_17244);
nor U17647 (N_17647,N_17205,N_17331);
nand U17648 (N_17648,N_17481,N_17087);
and U17649 (N_17649,N_17136,N_17260);
and U17650 (N_17650,N_17286,N_17077);
and U17651 (N_17651,N_17476,N_17209);
xor U17652 (N_17652,N_17405,N_17473);
nand U17653 (N_17653,N_17377,N_17292);
nand U17654 (N_17654,N_17392,N_17317);
and U17655 (N_17655,N_17010,N_17182);
and U17656 (N_17656,N_17132,N_17051);
or U17657 (N_17657,N_17479,N_17121);
xor U17658 (N_17658,N_17177,N_17346);
and U17659 (N_17659,N_17466,N_17485);
nor U17660 (N_17660,N_17192,N_17181);
nand U17661 (N_17661,N_17246,N_17344);
nand U17662 (N_17662,N_17165,N_17369);
or U17663 (N_17663,N_17334,N_17066);
nand U17664 (N_17664,N_17211,N_17011);
and U17665 (N_17665,N_17074,N_17245);
nor U17666 (N_17666,N_17353,N_17491);
and U17667 (N_17667,N_17075,N_17478);
or U17668 (N_17668,N_17395,N_17168);
and U17669 (N_17669,N_17253,N_17399);
and U17670 (N_17670,N_17480,N_17016);
xor U17671 (N_17671,N_17316,N_17064);
nor U17672 (N_17672,N_17273,N_17023);
nor U17673 (N_17673,N_17490,N_17083);
and U17674 (N_17674,N_17484,N_17362);
xor U17675 (N_17675,N_17309,N_17290);
nand U17676 (N_17676,N_17412,N_17021);
nor U17677 (N_17677,N_17400,N_17263);
nand U17678 (N_17678,N_17097,N_17187);
or U17679 (N_17679,N_17328,N_17488);
or U17680 (N_17680,N_17164,N_17422);
and U17681 (N_17681,N_17320,N_17004);
nand U17682 (N_17682,N_17119,N_17223);
and U17683 (N_17683,N_17207,N_17411);
nor U17684 (N_17684,N_17447,N_17222);
nor U17685 (N_17685,N_17093,N_17086);
nor U17686 (N_17686,N_17407,N_17281);
or U17687 (N_17687,N_17175,N_17429);
and U17688 (N_17688,N_17499,N_17274);
nor U17689 (N_17689,N_17279,N_17495);
nor U17690 (N_17690,N_17219,N_17201);
and U17691 (N_17691,N_17288,N_17324);
or U17692 (N_17692,N_17250,N_17408);
and U17693 (N_17693,N_17176,N_17393);
nand U17694 (N_17694,N_17356,N_17122);
nor U17695 (N_17695,N_17235,N_17327);
or U17696 (N_17696,N_17335,N_17432);
and U17697 (N_17697,N_17276,N_17338);
nor U17698 (N_17698,N_17376,N_17129);
and U17699 (N_17699,N_17464,N_17054);
or U17700 (N_17700,N_17492,N_17178);
and U17701 (N_17701,N_17084,N_17403);
and U17702 (N_17702,N_17311,N_17368);
nor U17703 (N_17703,N_17179,N_17197);
xor U17704 (N_17704,N_17001,N_17259);
nor U17705 (N_17705,N_17038,N_17043);
and U17706 (N_17706,N_17482,N_17443);
or U17707 (N_17707,N_17332,N_17470);
nor U17708 (N_17708,N_17063,N_17037);
and U17709 (N_17709,N_17030,N_17249);
nor U17710 (N_17710,N_17367,N_17446);
nand U17711 (N_17711,N_17457,N_17058);
or U17712 (N_17712,N_17149,N_17418);
or U17713 (N_17713,N_17391,N_17108);
xor U17714 (N_17714,N_17003,N_17226);
nand U17715 (N_17715,N_17104,N_17277);
nor U17716 (N_17716,N_17036,N_17455);
and U17717 (N_17717,N_17453,N_17110);
xor U17718 (N_17718,N_17428,N_17374);
nand U17719 (N_17719,N_17072,N_17007);
xor U17720 (N_17720,N_17319,N_17014);
nor U17721 (N_17721,N_17148,N_17456);
nand U17722 (N_17722,N_17116,N_17202);
xor U17723 (N_17723,N_17256,N_17199);
or U17724 (N_17724,N_17364,N_17150);
nor U17725 (N_17725,N_17323,N_17144);
and U17726 (N_17726,N_17045,N_17348);
and U17727 (N_17727,N_17106,N_17459);
nor U17728 (N_17728,N_17308,N_17046);
nor U17729 (N_17729,N_17423,N_17343);
and U17730 (N_17730,N_17436,N_17306);
nand U17731 (N_17731,N_17387,N_17006);
or U17732 (N_17732,N_17440,N_17157);
nor U17733 (N_17733,N_17254,N_17140);
nor U17734 (N_17734,N_17081,N_17071);
and U17735 (N_17735,N_17365,N_17123);
xor U17736 (N_17736,N_17375,N_17196);
nand U17737 (N_17737,N_17131,N_17049);
and U17738 (N_17738,N_17262,N_17137);
or U17739 (N_17739,N_17114,N_17450);
xor U17740 (N_17740,N_17022,N_17424);
and U17741 (N_17741,N_17128,N_17191);
nor U17742 (N_17742,N_17027,N_17035);
nand U17743 (N_17743,N_17163,N_17135);
xnor U17744 (N_17744,N_17489,N_17189);
and U17745 (N_17745,N_17291,N_17210);
nand U17746 (N_17746,N_17454,N_17032);
nor U17747 (N_17747,N_17134,N_17102);
and U17748 (N_17748,N_17303,N_17463);
or U17749 (N_17749,N_17486,N_17380);
nor U17750 (N_17750,N_17453,N_17122);
nor U17751 (N_17751,N_17450,N_17470);
nand U17752 (N_17752,N_17257,N_17122);
xor U17753 (N_17753,N_17418,N_17266);
or U17754 (N_17754,N_17329,N_17424);
xor U17755 (N_17755,N_17287,N_17366);
nor U17756 (N_17756,N_17368,N_17483);
nand U17757 (N_17757,N_17393,N_17350);
xor U17758 (N_17758,N_17305,N_17167);
or U17759 (N_17759,N_17442,N_17070);
xnor U17760 (N_17760,N_17244,N_17387);
xor U17761 (N_17761,N_17277,N_17412);
and U17762 (N_17762,N_17276,N_17178);
and U17763 (N_17763,N_17114,N_17045);
or U17764 (N_17764,N_17229,N_17387);
xor U17765 (N_17765,N_17435,N_17408);
nand U17766 (N_17766,N_17170,N_17489);
nor U17767 (N_17767,N_17070,N_17448);
and U17768 (N_17768,N_17360,N_17483);
nand U17769 (N_17769,N_17077,N_17358);
nor U17770 (N_17770,N_17480,N_17213);
or U17771 (N_17771,N_17330,N_17268);
nor U17772 (N_17772,N_17342,N_17432);
nand U17773 (N_17773,N_17193,N_17486);
nand U17774 (N_17774,N_17193,N_17441);
nor U17775 (N_17775,N_17161,N_17403);
and U17776 (N_17776,N_17036,N_17495);
or U17777 (N_17777,N_17050,N_17288);
and U17778 (N_17778,N_17394,N_17081);
xnor U17779 (N_17779,N_17060,N_17193);
nand U17780 (N_17780,N_17313,N_17260);
and U17781 (N_17781,N_17176,N_17129);
or U17782 (N_17782,N_17470,N_17376);
nor U17783 (N_17783,N_17278,N_17296);
nand U17784 (N_17784,N_17244,N_17100);
nor U17785 (N_17785,N_17246,N_17217);
or U17786 (N_17786,N_17290,N_17043);
and U17787 (N_17787,N_17316,N_17271);
or U17788 (N_17788,N_17008,N_17277);
nor U17789 (N_17789,N_17221,N_17186);
nand U17790 (N_17790,N_17355,N_17020);
nor U17791 (N_17791,N_17121,N_17372);
or U17792 (N_17792,N_17146,N_17102);
xnor U17793 (N_17793,N_17443,N_17077);
xnor U17794 (N_17794,N_17466,N_17221);
or U17795 (N_17795,N_17347,N_17117);
or U17796 (N_17796,N_17433,N_17499);
nor U17797 (N_17797,N_17409,N_17289);
nor U17798 (N_17798,N_17023,N_17217);
xnor U17799 (N_17799,N_17002,N_17090);
or U17800 (N_17800,N_17108,N_17100);
or U17801 (N_17801,N_17296,N_17010);
nand U17802 (N_17802,N_17363,N_17444);
and U17803 (N_17803,N_17390,N_17452);
nor U17804 (N_17804,N_17204,N_17097);
nand U17805 (N_17805,N_17293,N_17042);
nor U17806 (N_17806,N_17287,N_17343);
or U17807 (N_17807,N_17264,N_17455);
and U17808 (N_17808,N_17350,N_17435);
xor U17809 (N_17809,N_17177,N_17450);
nor U17810 (N_17810,N_17326,N_17245);
xor U17811 (N_17811,N_17124,N_17367);
xor U17812 (N_17812,N_17450,N_17378);
or U17813 (N_17813,N_17064,N_17353);
xor U17814 (N_17814,N_17213,N_17310);
xor U17815 (N_17815,N_17245,N_17008);
nor U17816 (N_17816,N_17246,N_17375);
nor U17817 (N_17817,N_17361,N_17284);
or U17818 (N_17818,N_17004,N_17181);
and U17819 (N_17819,N_17049,N_17133);
xor U17820 (N_17820,N_17306,N_17478);
or U17821 (N_17821,N_17428,N_17309);
nand U17822 (N_17822,N_17105,N_17251);
xor U17823 (N_17823,N_17139,N_17037);
xor U17824 (N_17824,N_17376,N_17449);
or U17825 (N_17825,N_17417,N_17395);
and U17826 (N_17826,N_17071,N_17293);
or U17827 (N_17827,N_17383,N_17373);
or U17828 (N_17828,N_17059,N_17360);
nand U17829 (N_17829,N_17452,N_17321);
nand U17830 (N_17830,N_17464,N_17106);
nor U17831 (N_17831,N_17355,N_17463);
xnor U17832 (N_17832,N_17345,N_17020);
nand U17833 (N_17833,N_17009,N_17114);
or U17834 (N_17834,N_17417,N_17412);
nand U17835 (N_17835,N_17272,N_17458);
xor U17836 (N_17836,N_17000,N_17103);
nand U17837 (N_17837,N_17108,N_17296);
nor U17838 (N_17838,N_17363,N_17225);
nor U17839 (N_17839,N_17436,N_17300);
nand U17840 (N_17840,N_17244,N_17369);
xnor U17841 (N_17841,N_17200,N_17015);
xnor U17842 (N_17842,N_17053,N_17073);
xnor U17843 (N_17843,N_17041,N_17091);
xor U17844 (N_17844,N_17149,N_17439);
and U17845 (N_17845,N_17312,N_17375);
nor U17846 (N_17846,N_17496,N_17052);
nand U17847 (N_17847,N_17348,N_17066);
and U17848 (N_17848,N_17420,N_17254);
nor U17849 (N_17849,N_17303,N_17006);
nor U17850 (N_17850,N_17428,N_17008);
nor U17851 (N_17851,N_17025,N_17183);
nor U17852 (N_17852,N_17087,N_17211);
nand U17853 (N_17853,N_17286,N_17232);
and U17854 (N_17854,N_17118,N_17068);
and U17855 (N_17855,N_17312,N_17438);
or U17856 (N_17856,N_17087,N_17059);
or U17857 (N_17857,N_17456,N_17340);
or U17858 (N_17858,N_17485,N_17233);
nand U17859 (N_17859,N_17330,N_17337);
nand U17860 (N_17860,N_17097,N_17312);
nand U17861 (N_17861,N_17020,N_17229);
nand U17862 (N_17862,N_17127,N_17417);
nand U17863 (N_17863,N_17030,N_17379);
and U17864 (N_17864,N_17131,N_17327);
and U17865 (N_17865,N_17456,N_17403);
xnor U17866 (N_17866,N_17336,N_17273);
nand U17867 (N_17867,N_17017,N_17012);
xor U17868 (N_17868,N_17202,N_17320);
nor U17869 (N_17869,N_17253,N_17405);
xnor U17870 (N_17870,N_17395,N_17266);
nor U17871 (N_17871,N_17250,N_17460);
or U17872 (N_17872,N_17258,N_17289);
and U17873 (N_17873,N_17407,N_17191);
nand U17874 (N_17874,N_17248,N_17074);
or U17875 (N_17875,N_17112,N_17228);
nor U17876 (N_17876,N_17475,N_17247);
nor U17877 (N_17877,N_17155,N_17086);
nor U17878 (N_17878,N_17491,N_17220);
and U17879 (N_17879,N_17454,N_17496);
or U17880 (N_17880,N_17224,N_17083);
or U17881 (N_17881,N_17013,N_17158);
nor U17882 (N_17882,N_17154,N_17431);
and U17883 (N_17883,N_17405,N_17059);
xor U17884 (N_17884,N_17103,N_17045);
nor U17885 (N_17885,N_17411,N_17394);
or U17886 (N_17886,N_17324,N_17315);
xnor U17887 (N_17887,N_17487,N_17238);
and U17888 (N_17888,N_17471,N_17255);
nand U17889 (N_17889,N_17067,N_17306);
and U17890 (N_17890,N_17010,N_17319);
xnor U17891 (N_17891,N_17432,N_17497);
nand U17892 (N_17892,N_17018,N_17408);
and U17893 (N_17893,N_17245,N_17449);
nor U17894 (N_17894,N_17132,N_17321);
xor U17895 (N_17895,N_17448,N_17145);
nor U17896 (N_17896,N_17342,N_17125);
nor U17897 (N_17897,N_17221,N_17123);
or U17898 (N_17898,N_17447,N_17489);
or U17899 (N_17899,N_17202,N_17355);
nand U17900 (N_17900,N_17176,N_17405);
nor U17901 (N_17901,N_17364,N_17213);
nand U17902 (N_17902,N_17072,N_17456);
xor U17903 (N_17903,N_17225,N_17136);
or U17904 (N_17904,N_17097,N_17209);
xor U17905 (N_17905,N_17173,N_17484);
xnor U17906 (N_17906,N_17463,N_17296);
xor U17907 (N_17907,N_17034,N_17362);
xor U17908 (N_17908,N_17368,N_17127);
and U17909 (N_17909,N_17497,N_17212);
xor U17910 (N_17910,N_17383,N_17234);
nor U17911 (N_17911,N_17327,N_17005);
nand U17912 (N_17912,N_17343,N_17055);
xnor U17913 (N_17913,N_17357,N_17276);
xnor U17914 (N_17914,N_17079,N_17456);
xnor U17915 (N_17915,N_17489,N_17316);
nand U17916 (N_17916,N_17314,N_17117);
and U17917 (N_17917,N_17069,N_17084);
nor U17918 (N_17918,N_17067,N_17229);
or U17919 (N_17919,N_17480,N_17382);
xor U17920 (N_17920,N_17402,N_17376);
or U17921 (N_17921,N_17113,N_17224);
or U17922 (N_17922,N_17465,N_17385);
nor U17923 (N_17923,N_17382,N_17436);
and U17924 (N_17924,N_17111,N_17439);
or U17925 (N_17925,N_17181,N_17159);
nand U17926 (N_17926,N_17132,N_17111);
nand U17927 (N_17927,N_17134,N_17488);
xnor U17928 (N_17928,N_17420,N_17020);
nor U17929 (N_17929,N_17208,N_17202);
nor U17930 (N_17930,N_17498,N_17089);
xor U17931 (N_17931,N_17262,N_17357);
nand U17932 (N_17932,N_17193,N_17450);
xnor U17933 (N_17933,N_17478,N_17322);
nor U17934 (N_17934,N_17096,N_17131);
or U17935 (N_17935,N_17385,N_17218);
nand U17936 (N_17936,N_17288,N_17140);
xnor U17937 (N_17937,N_17211,N_17380);
or U17938 (N_17938,N_17428,N_17499);
and U17939 (N_17939,N_17378,N_17225);
or U17940 (N_17940,N_17319,N_17440);
and U17941 (N_17941,N_17134,N_17059);
and U17942 (N_17942,N_17191,N_17486);
nor U17943 (N_17943,N_17455,N_17386);
or U17944 (N_17944,N_17140,N_17335);
nor U17945 (N_17945,N_17370,N_17271);
or U17946 (N_17946,N_17102,N_17480);
xor U17947 (N_17947,N_17237,N_17044);
nand U17948 (N_17948,N_17384,N_17481);
xnor U17949 (N_17949,N_17190,N_17032);
nor U17950 (N_17950,N_17330,N_17467);
and U17951 (N_17951,N_17062,N_17427);
nor U17952 (N_17952,N_17112,N_17345);
and U17953 (N_17953,N_17071,N_17235);
or U17954 (N_17954,N_17234,N_17054);
xnor U17955 (N_17955,N_17330,N_17233);
nand U17956 (N_17956,N_17287,N_17126);
nand U17957 (N_17957,N_17358,N_17458);
or U17958 (N_17958,N_17253,N_17364);
nor U17959 (N_17959,N_17397,N_17043);
nand U17960 (N_17960,N_17122,N_17120);
nand U17961 (N_17961,N_17455,N_17272);
nor U17962 (N_17962,N_17457,N_17132);
nand U17963 (N_17963,N_17069,N_17433);
nand U17964 (N_17964,N_17035,N_17186);
xnor U17965 (N_17965,N_17397,N_17443);
or U17966 (N_17966,N_17080,N_17120);
xnor U17967 (N_17967,N_17004,N_17187);
xnor U17968 (N_17968,N_17238,N_17342);
nand U17969 (N_17969,N_17088,N_17209);
nor U17970 (N_17970,N_17416,N_17165);
xor U17971 (N_17971,N_17228,N_17372);
nand U17972 (N_17972,N_17169,N_17223);
nor U17973 (N_17973,N_17406,N_17416);
xnor U17974 (N_17974,N_17154,N_17257);
nor U17975 (N_17975,N_17489,N_17399);
xor U17976 (N_17976,N_17401,N_17074);
and U17977 (N_17977,N_17477,N_17213);
xor U17978 (N_17978,N_17286,N_17328);
nand U17979 (N_17979,N_17121,N_17120);
nor U17980 (N_17980,N_17027,N_17375);
xnor U17981 (N_17981,N_17203,N_17329);
nor U17982 (N_17982,N_17057,N_17291);
xor U17983 (N_17983,N_17051,N_17355);
nand U17984 (N_17984,N_17279,N_17352);
or U17985 (N_17985,N_17144,N_17334);
and U17986 (N_17986,N_17249,N_17345);
nor U17987 (N_17987,N_17096,N_17102);
nand U17988 (N_17988,N_17244,N_17190);
nor U17989 (N_17989,N_17298,N_17022);
nand U17990 (N_17990,N_17377,N_17096);
nor U17991 (N_17991,N_17267,N_17402);
and U17992 (N_17992,N_17221,N_17418);
or U17993 (N_17993,N_17184,N_17065);
xor U17994 (N_17994,N_17055,N_17266);
xor U17995 (N_17995,N_17248,N_17095);
nand U17996 (N_17996,N_17079,N_17254);
nor U17997 (N_17997,N_17198,N_17312);
xor U17998 (N_17998,N_17438,N_17365);
xor U17999 (N_17999,N_17007,N_17436);
nor U18000 (N_18000,N_17783,N_17761);
nor U18001 (N_18001,N_17938,N_17904);
or U18002 (N_18002,N_17713,N_17670);
nand U18003 (N_18003,N_17678,N_17986);
nor U18004 (N_18004,N_17797,N_17805);
nor U18005 (N_18005,N_17943,N_17529);
nand U18006 (N_18006,N_17710,N_17769);
or U18007 (N_18007,N_17849,N_17756);
xnor U18008 (N_18008,N_17758,N_17975);
or U18009 (N_18009,N_17693,N_17755);
nand U18010 (N_18010,N_17559,N_17626);
and U18011 (N_18011,N_17926,N_17861);
nand U18012 (N_18012,N_17820,N_17663);
xor U18013 (N_18013,N_17882,N_17563);
nand U18014 (N_18014,N_17645,N_17969);
nand U18015 (N_18015,N_17729,N_17657);
or U18016 (N_18016,N_17618,N_17779);
nor U18017 (N_18017,N_17537,N_17964);
and U18018 (N_18018,N_17891,N_17649);
and U18019 (N_18019,N_17680,N_17522);
nor U18020 (N_18020,N_17633,N_17936);
nand U18021 (N_18021,N_17990,N_17772);
or U18022 (N_18022,N_17617,N_17946);
or U18023 (N_18023,N_17698,N_17658);
and U18024 (N_18024,N_17875,N_17933);
or U18025 (N_18025,N_17997,N_17564);
or U18026 (N_18026,N_17767,N_17907);
and U18027 (N_18027,N_17738,N_17793);
nor U18028 (N_18028,N_17505,N_17570);
xor U18029 (N_18029,N_17578,N_17801);
nor U18030 (N_18030,N_17668,N_17571);
or U18031 (N_18031,N_17838,N_17593);
or U18032 (N_18032,N_17836,N_17749);
and U18033 (N_18033,N_17695,N_17546);
xor U18034 (N_18034,N_17700,N_17606);
nor U18035 (N_18035,N_17665,N_17798);
and U18036 (N_18036,N_17818,N_17995);
or U18037 (N_18037,N_17650,N_17583);
and U18038 (N_18038,N_17994,N_17746);
nand U18039 (N_18039,N_17551,N_17955);
nor U18040 (N_18040,N_17978,N_17586);
or U18041 (N_18041,N_17776,N_17603);
nor U18042 (N_18042,N_17972,N_17962);
or U18043 (N_18043,N_17701,N_17900);
nor U18044 (N_18044,N_17810,N_17591);
and U18045 (N_18045,N_17582,N_17515);
nand U18046 (N_18046,N_17817,N_17886);
nor U18047 (N_18047,N_17655,N_17902);
nor U18048 (N_18048,N_17619,N_17653);
xnor U18049 (N_18049,N_17961,N_17862);
or U18050 (N_18050,N_17858,N_17737);
and U18051 (N_18051,N_17624,N_17974);
and U18052 (N_18052,N_17516,N_17641);
or U18053 (N_18053,N_17952,N_17535);
xor U18054 (N_18054,N_17868,N_17834);
and U18055 (N_18055,N_17945,N_17677);
nor U18056 (N_18056,N_17527,N_17682);
nor U18057 (N_18057,N_17764,N_17830);
nor U18058 (N_18058,N_17799,N_17828);
nand U18059 (N_18059,N_17599,N_17745);
xor U18060 (N_18060,N_17659,N_17689);
or U18061 (N_18061,N_17719,N_17681);
xor U18062 (N_18062,N_17574,N_17855);
and U18063 (N_18063,N_17601,N_17837);
or U18064 (N_18064,N_17747,N_17743);
or U18065 (N_18065,N_17925,N_17850);
xor U18066 (N_18066,N_17898,N_17876);
and U18067 (N_18067,N_17811,N_17757);
and U18068 (N_18068,N_17560,N_17735);
nand U18069 (N_18069,N_17565,N_17513);
nand U18070 (N_18070,N_17924,N_17860);
and U18071 (N_18071,N_17621,N_17730);
xnor U18072 (N_18072,N_17647,N_17935);
nand U18073 (N_18073,N_17821,N_17542);
xor U18074 (N_18074,N_17960,N_17775);
nand U18075 (N_18075,N_17726,N_17800);
nand U18076 (N_18076,N_17781,N_17620);
nor U18077 (N_18077,N_17789,N_17813);
nor U18078 (N_18078,N_17552,N_17991);
xor U18079 (N_18079,N_17521,N_17625);
or U18080 (N_18080,N_17632,N_17976);
xnor U18081 (N_18081,N_17556,N_17637);
nand U18082 (N_18082,N_17672,N_17917);
nand U18083 (N_18083,N_17751,N_17567);
or U18084 (N_18084,N_17534,N_17733);
nor U18085 (N_18085,N_17533,N_17629);
nand U18086 (N_18086,N_17768,N_17806);
and U18087 (N_18087,N_17883,N_17598);
nor U18088 (N_18088,N_17888,N_17708);
and U18089 (N_18089,N_17644,N_17506);
nor U18090 (N_18090,N_17538,N_17980);
and U18091 (N_18091,N_17832,N_17794);
xor U18092 (N_18092,N_17615,N_17690);
and U18093 (N_18093,N_17909,N_17592);
nor U18094 (N_18094,N_17833,N_17628);
xnor U18095 (N_18095,N_17877,N_17854);
xnor U18096 (N_18096,N_17796,N_17989);
nand U18097 (N_18097,N_17892,N_17717);
xnor U18098 (N_18098,N_17687,N_17580);
or U18099 (N_18099,N_17740,N_17895);
xnor U18100 (N_18100,N_17750,N_17587);
or U18101 (N_18101,N_17508,N_17627);
and U18102 (N_18102,N_17760,N_17992);
xnor U18103 (N_18103,N_17863,N_17514);
and U18104 (N_18104,N_17608,N_17654);
nand U18105 (N_18105,N_17770,N_17503);
or U18106 (N_18106,N_17727,N_17584);
or U18107 (N_18107,N_17525,N_17967);
nand U18108 (N_18108,N_17963,N_17981);
and U18109 (N_18109,N_17763,N_17539);
and U18110 (N_18110,N_17970,N_17667);
nand U18111 (N_18111,N_17511,N_17993);
nand U18112 (N_18112,N_17613,N_17576);
or U18113 (N_18113,N_17694,N_17893);
or U18114 (N_18114,N_17896,N_17906);
and U18115 (N_18115,N_17787,N_17673);
nor U18116 (N_18116,N_17814,N_17662);
or U18117 (N_18117,N_17928,N_17867);
nand U18118 (N_18118,N_17942,N_17716);
nor U18119 (N_18119,N_17922,N_17872);
nor U18120 (N_18120,N_17610,N_17754);
and U18121 (N_18121,N_17709,N_17819);
or U18122 (N_18122,N_17742,N_17822);
xnor U18123 (N_18123,N_17519,N_17611);
and U18124 (N_18124,N_17845,N_17616);
nor U18125 (N_18125,N_17941,N_17815);
and U18126 (N_18126,N_17785,N_17696);
or U18127 (N_18127,N_17953,N_17864);
nor U18128 (N_18128,N_17884,N_17512);
and U18129 (N_18129,N_17510,N_17968);
nor U18130 (N_18130,N_17622,N_17531);
xor U18131 (N_18131,N_17550,N_17699);
and U18132 (N_18132,N_17866,N_17859);
nor U18133 (N_18133,N_17736,N_17724);
xor U18134 (N_18134,N_17762,N_17500);
and U18135 (N_18135,N_17752,N_17734);
xnor U18136 (N_18136,N_17966,N_17596);
and U18137 (N_18137,N_17977,N_17804);
nor U18138 (N_18138,N_17623,N_17913);
nor U18139 (N_18139,N_17612,N_17518);
xor U18140 (N_18140,N_17841,N_17930);
nor U18141 (N_18141,N_17791,N_17949);
xor U18142 (N_18142,N_17722,N_17605);
nand U18143 (N_18143,N_17651,N_17532);
nor U18144 (N_18144,N_17914,N_17524);
and U18145 (N_18145,N_17642,N_17741);
nor U18146 (N_18146,N_17530,N_17685);
and U18147 (N_18147,N_17725,N_17575);
nand U18148 (N_18148,N_17509,N_17697);
and U18149 (N_18149,N_17865,N_17544);
nor U18150 (N_18150,N_17950,N_17979);
nand U18151 (N_18151,N_17923,N_17912);
or U18152 (N_18152,N_17573,N_17631);
or U18153 (N_18153,N_17840,N_17501);
nor U18154 (N_18154,N_17703,N_17869);
xnor U18155 (N_18155,N_17604,N_17517);
or U18156 (N_18156,N_17848,N_17857);
nor U18157 (N_18157,N_17705,N_17988);
and U18158 (N_18158,N_17825,N_17777);
and U18159 (N_18159,N_17894,N_17744);
nand U18160 (N_18160,N_17874,N_17853);
and U18161 (N_18161,N_17948,N_17634);
nor U18162 (N_18162,N_17640,N_17784);
nand U18163 (N_18163,N_17648,N_17939);
nor U18164 (N_18164,N_17577,N_17720);
nand U18165 (N_18165,N_17790,N_17971);
xor U18166 (N_18166,N_17905,N_17998);
nor U18167 (N_18167,N_17569,N_17664);
xor U18168 (N_18168,N_17932,N_17636);
nand U18169 (N_18169,N_17915,N_17526);
nor U18170 (N_18170,N_17780,N_17973);
xnor U18171 (N_18171,N_17607,N_17951);
nor U18172 (N_18172,N_17773,N_17985);
nand U18173 (N_18173,N_17721,N_17782);
and U18174 (N_18174,N_17839,N_17712);
nand U18175 (N_18175,N_17844,N_17590);
or U18176 (N_18176,N_17630,N_17929);
and U18177 (N_18177,N_17666,N_17808);
nand U18178 (N_18178,N_17683,N_17554);
or U18179 (N_18179,N_17520,N_17829);
nand U18180 (N_18180,N_17809,N_17944);
nor U18181 (N_18181,N_17771,N_17954);
nand U18182 (N_18182,N_17553,N_17879);
nand U18183 (N_18183,N_17684,N_17919);
nand U18184 (N_18184,N_17675,N_17502);
nand U18185 (N_18185,N_17878,N_17691);
nor U18186 (N_18186,N_17831,N_17851);
nor U18187 (N_18187,N_17549,N_17558);
xor U18188 (N_18188,N_17600,N_17885);
xnor U18189 (N_18189,N_17507,N_17807);
nor U18190 (N_18190,N_17897,N_17816);
xnor U18191 (N_18191,N_17660,N_17823);
or U18192 (N_18192,N_17581,N_17786);
nor U18193 (N_18193,N_17908,N_17589);
nor U18194 (N_18194,N_17568,N_17723);
nor U18195 (N_18195,N_17983,N_17802);
and U18196 (N_18196,N_17852,N_17555);
and U18197 (N_18197,N_17910,N_17842);
nor U18198 (N_18198,N_17788,N_17999);
or U18199 (N_18199,N_17557,N_17987);
nand U18200 (N_18200,N_17901,N_17566);
or U18201 (N_18201,N_17847,N_17585);
xnor U18202 (N_18202,N_17702,N_17728);
nand U18203 (N_18203,N_17889,N_17595);
and U18204 (N_18204,N_17543,N_17614);
and U18205 (N_18205,N_17843,N_17541);
nor U18206 (N_18206,N_17548,N_17957);
xnor U18207 (N_18207,N_17937,N_17940);
xnor U18208 (N_18208,N_17870,N_17956);
and U18209 (N_18209,N_17661,N_17827);
nor U18210 (N_18210,N_17759,N_17921);
or U18211 (N_18211,N_17679,N_17602);
and U18212 (N_18212,N_17982,N_17887);
nor U18213 (N_18213,N_17748,N_17674);
and U18214 (N_18214,N_17873,N_17871);
nand U18215 (N_18215,N_17545,N_17714);
or U18216 (N_18216,N_17732,N_17856);
and U18217 (N_18217,N_17911,N_17890);
nor U18218 (N_18218,N_17916,N_17669);
xnor U18219 (N_18219,N_17635,N_17765);
nor U18220 (N_18220,N_17918,N_17766);
nor U18221 (N_18221,N_17947,N_17934);
and U18222 (N_18222,N_17753,N_17597);
or U18223 (N_18223,N_17639,N_17504);
and U18224 (N_18224,N_17706,N_17778);
and U18225 (N_18225,N_17881,N_17927);
xnor U18226 (N_18226,N_17686,N_17646);
and U18227 (N_18227,N_17931,N_17652);
nor U18228 (N_18228,N_17899,N_17718);
nand U18229 (N_18229,N_17536,N_17846);
and U18230 (N_18230,N_17656,N_17588);
xnor U18231 (N_18231,N_17774,N_17711);
xnor U18232 (N_18232,N_17824,N_17903);
or U18233 (N_18233,N_17920,N_17638);
nor U18234 (N_18234,N_17739,N_17561);
and U18235 (N_18235,N_17688,N_17547);
nand U18236 (N_18236,N_17643,N_17958);
and U18237 (N_18237,N_17523,N_17579);
or U18238 (N_18238,N_17812,N_17540);
and U18239 (N_18239,N_17594,N_17965);
nand U18240 (N_18240,N_17671,N_17562);
and U18241 (N_18241,N_17959,N_17795);
nand U18242 (N_18242,N_17792,N_17826);
or U18243 (N_18243,N_17880,N_17692);
and U18244 (N_18244,N_17715,N_17803);
nor U18245 (N_18245,N_17609,N_17528);
or U18246 (N_18246,N_17835,N_17676);
or U18247 (N_18247,N_17984,N_17996);
xnor U18248 (N_18248,N_17572,N_17707);
or U18249 (N_18249,N_17731,N_17704);
or U18250 (N_18250,N_17959,N_17758);
xnor U18251 (N_18251,N_17970,N_17895);
or U18252 (N_18252,N_17721,N_17673);
nor U18253 (N_18253,N_17977,N_17935);
nor U18254 (N_18254,N_17661,N_17843);
or U18255 (N_18255,N_17714,N_17562);
and U18256 (N_18256,N_17964,N_17759);
and U18257 (N_18257,N_17692,N_17794);
nor U18258 (N_18258,N_17810,N_17614);
nor U18259 (N_18259,N_17927,N_17563);
or U18260 (N_18260,N_17640,N_17923);
xnor U18261 (N_18261,N_17879,N_17603);
and U18262 (N_18262,N_17943,N_17836);
and U18263 (N_18263,N_17786,N_17783);
nand U18264 (N_18264,N_17701,N_17803);
nand U18265 (N_18265,N_17699,N_17651);
and U18266 (N_18266,N_17513,N_17582);
nor U18267 (N_18267,N_17521,N_17687);
or U18268 (N_18268,N_17916,N_17943);
and U18269 (N_18269,N_17577,N_17556);
nand U18270 (N_18270,N_17767,N_17734);
nand U18271 (N_18271,N_17933,N_17625);
or U18272 (N_18272,N_17955,N_17557);
and U18273 (N_18273,N_17916,N_17869);
nor U18274 (N_18274,N_17539,N_17726);
nand U18275 (N_18275,N_17636,N_17561);
nor U18276 (N_18276,N_17645,N_17944);
and U18277 (N_18277,N_17948,N_17814);
or U18278 (N_18278,N_17937,N_17973);
nand U18279 (N_18279,N_17843,N_17567);
nand U18280 (N_18280,N_17650,N_17752);
nor U18281 (N_18281,N_17692,N_17984);
and U18282 (N_18282,N_17861,N_17743);
xnor U18283 (N_18283,N_17568,N_17698);
or U18284 (N_18284,N_17822,N_17550);
or U18285 (N_18285,N_17957,N_17752);
or U18286 (N_18286,N_17727,N_17962);
and U18287 (N_18287,N_17664,N_17648);
and U18288 (N_18288,N_17730,N_17519);
nand U18289 (N_18289,N_17785,N_17959);
nor U18290 (N_18290,N_17689,N_17838);
xor U18291 (N_18291,N_17763,N_17551);
xnor U18292 (N_18292,N_17787,N_17966);
or U18293 (N_18293,N_17834,N_17782);
xor U18294 (N_18294,N_17999,N_17910);
xor U18295 (N_18295,N_17977,N_17766);
nor U18296 (N_18296,N_17675,N_17706);
xnor U18297 (N_18297,N_17617,N_17520);
and U18298 (N_18298,N_17566,N_17737);
nor U18299 (N_18299,N_17847,N_17717);
nor U18300 (N_18300,N_17977,N_17758);
xnor U18301 (N_18301,N_17929,N_17562);
nand U18302 (N_18302,N_17789,N_17757);
nand U18303 (N_18303,N_17998,N_17906);
and U18304 (N_18304,N_17808,N_17800);
nand U18305 (N_18305,N_17524,N_17521);
xnor U18306 (N_18306,N_17766,N_17937);
nor U18307 (N_18307,N_17613,N_17964);
or U18308 (N_18308,N_17589,N_17657);
or U18309 (N_18309,N_17941,N_17995);
and U18310 (N_18310,N_17585,N_17857);
and U18311 (N_18311,N_17956,N_17985);
nand U18312 (N_18312,N_17686,N_17639);
or U18313 (N_18313,N_17727,N_17772);
or U18314 (N_18314,N_17834,N_17867);
nor U18315 (N_18315,N_17625,N_17528);
and U18316 (N_18316,N_17572,N_17849);
or U18317 (N_18317,N_17718,N_17613);
and U18318 (N_18318,N_17543,N_17620);
or U18319 (N_18319,N_17944,N_17982);
or U18320 (N_18320,N_17530,N_17803);
nor U18321 (N_18321,N_17603,N_17548);
or U18322 (N_18322,N_17890,N_17944);
and U18323 (N_18323,N_17710,N_17771);
xor U18324 (N_18324,N_17966,N_17551);
xnor U18325 (N_18325,N_17860,N_17787);
nor U18326 (N_18326,N_17760,N_17631);
and U18327 (N_18327,N_17916,N_17918);
nand U18328 (N_18328,N_17607,N_17975);
or U18329 (N_18329,N_17729,N_17923);
or U18330 (N_18330,N_17887,N_17893);
or U18331 (N_18331,N_17899,N_17794);
xor U18332 (N_18332,N_17718,N_17749);
xnor U18333 (N_18333,N_17701,N_17711);
xor U18334 (N_18334,N_17650,N_17569);
and U18335 (N_18335,N_17977,N_17822);
or U18336 (N_18336,N_17611,N_17806);
nand U18337 (N_18337,N_17663,N_17515);
xnor U18338 (N_18338,N_17757,N_17608);
and U18339 (N_18339,N_17595,N_17583);
and U18340 (N_18340,N_17849,N_17662);
nor U18341 (N_18341,N_17567,N_17692);
nor U18342 (N_18342,N_17666,N_17563);
xor U18343 (N_18343,N_17737,N_17514);
xnor U18344 (N_18344,N_17511,N_17539);
nor U18345 (N_18345,N_17844,N_17801);
nor U18346 (N_18346,N_17735,N_17621);
xor U18347 (N_18347,N_17883,N_17619);
and U18348 (N_18348,N_17979,N_17732);
and U18349 (N_18349,N_17746,N_17770);
nand U18350 (N_18350,N_17551,N_17788);
or U18351 (N_18351,N_17874,N_17817);
nand U18352 (N_18352,N_17524,N_17923);
nor U18353 (N_18353,N_17898,N_17544);
xnor U18354 (N_18354,N_17566,N_17718);
nand U18355 (N_18355,N_17770,N_17923);
nand U18356 (N_18356,N_17626,N_17812);
and U18357 (N_18357,N_17918,N_17985);
nor U18358 (N_18358,N_17675,N_17652);
xnor U18359 (N_18359,N_17754,N_17526);
nor U18360 (N_18360,N_17975,N_17591);
nor U18361 (N_18361,N_17684,N_17990);
xnor U18362 (N_18362,N_17886,N_17974);
or U18363 (N_18363,N_17964,N_17910);
and U18364 (N_18364,N_17594,N_17679);
nor U18365 (N_18365,N_17749,N_17666);
or U18366 (N_18366,N_17787,N_17969);
or U18367 (N_18367,N_17884,N_17661);
nor U18368 (N_18368,N_17918,N_17967);
or U18369 (N_18369,N_17859,N_17748);
nand U18370 (N_18370,N_17822,N_17891);
and U18371 (N_18371,N_17632,N_17834);
nor U18372 (N_18372,N_17707,N_17841);
nand U18373 (N_18373,N_17982,N_17593);
or U18374 (N_18374,N_17846,N_17900);
or U18375 (N_18375,N_17665,N_17871);
nor U18376 (N_18376,N_17721,N_17706);
xnor U18377 (N_18377,N_17719,N_17549);
or U18378 (N_18378,N_17748,N_17586);
nand U18379 (N_18379,N_17715,N_17675);
and U18380 (N_18380,N_17521,N_17757);
or U18381 (N_18381,N_17636,N_17953);
nand U18382 (N_18382,N_17512,N_17632);
xnor U18383 (N_18383,N_17972,N_17582);
nand U18384 (N_18384,N_17958,N_17942);
or U18385 (N_18385,N_17891,N_17721);
nand U18386 (N_18386,N_17748,N_17523);
nor U18387 (N_18387,N_17704,N_17895);
and U18388 (N_18388,N_17889,N_17734);
nand U18389 (N_18389,N_17507,N_17749);
and U18390 (N_18390,N_17641,N_17634);
xnor U18391 (N_18391,N_17536,N_17706);
nand U18392 (N_18392,N_17918,N_17883);
or U18393 (N_18393,N_17774,N_17723);
xnor U18394 (N_18394,N_17578,N_17807);
xor U18395 (N_18395,N_17591,N_17862);
and U18396 (N_18396,N_17670,N_17627);
xnor U18397 (N_18397,N_17710,N_17847);
nand U18398 (N_18398,N_17594,N_17834);
xnor U18399 (N_18399,N_17848,N_17831);
nor U18400 (N_18400,N_17556,N_17954);
and U18401 (N_18401,N_17599,N_17849);
or U18402 (N_18402,N_17903,N_17934);
and U18403 (N_18403,N_17822,N_17938);
nand U18404 (N_18404,N_17889,N_17876);
or U18405 (N_18405,N_17723,N_17959);
nor U18406 (N_18406,N_17811,N_17891);
nor U18407 (N_18407,N_17995,N_17635);
xor U18408 (N_18408,N_17578,N_17645);
nor U18409 (N_18409,N_17598,N_17936);
or U18410 (N_18410,N_17711,N_17740);
nor U18411 (N_18411,N_17832,N_17828);
nand U18412 (N_18412,N_17802,N_17921);
nand U18413 (N_18413,N_17551,N_17544);
xor U18414 (N_18414,N_17963,N_17745);
xnor U18415 (N_18415,N_17907,N_17510);
nand U18416 (N_18416,N_17655,N_17728);
nand U18417 (N_18417,N_17730,N_17767);
or U18418 (N_18418,N_17782,N_17980);
and U18419 (N_18419,N_17871,N_17638);
xor U18420 (N_18420,N_17734,N_17692);
and U18421 (N_18421,N_17980,N_17759);
xnor U18422 (N_18422,N_17622,N_17772);
xor U18423 (N_18423,N_17742,N_17692);
and U18424 (N_18424,N_17830,N_17616);
nand U18425 (N_18425,N_17813,N_17636);
nor U18426 (N_18426,N_17775,N_17984);
nor U18427 (N_18427,N_17501,N_17833);
nor U18428 (N_18428,N_17828,N_17729);
nand U18429 (N_18429,N_17520,N_17985);
and U18430 (N_18430,N_17799,N_17539);
and U18431 (N_18431,N_17716,N_17803);
nor U18432 (N_18432,N_17718,N_17748);
xnor U18433 (N_18433,N_17703,N_17814);
xnor U18434 (N_18434,N_17889,N_17758);
or U18435 (N_18435,N_17659,N_17946);
and U18436 (N_18436,N_17662,N_17583);
xor U18437 (N_18437,N_17604,N_17730);
nand U18438 (N_18438,N_17502,N_17878);
xor U18439 (N_18439,N_17544,N_17634);
or U18440 (N_18440,N_17615,N_17978);
nand U18441 (N_18441,N_17886,N_17862);
or U18442 (N_18442,N_17539,N_17959);
and U18443 (N_18443,N_17598,N_17792);
or U18444 (N_18444,N_17928,N_17670);
xnor U18445 (N_18445,N_17996,N_17744);
and U18446 (N_18446,N_17664,N_17502);
or U18447 (N_18447,N_17533,N_17531);
and U18448 (N_18448,N_17827,N_17561);
nor U18449 (N_18449,N_17559,N_17502);
xor U18450 (N_18450,N_17758,N_17654);
nor U18451 (N_18451,N_17739,N_17749);
and U18452 (N_18452,N_17506,N_17933);
nand U18453 (N_18453,N_17618,N_17631);
or U18454 (N_18454,N_17723,N_17694);
and U18455 (N_18455,N_17779,N_17567);
xnor U18456 (N_18456,N_17712,N_17754);
nand U18457 (N_18457,N_17880,N_17848);
nor U18458 (N_18458,N_17857,N_17934);
nand U18459 (N_18459,N_17929,N_17769);
xnor U18460 (N_18460,N_17648,N_17925);
xnor U18461 (N_18461,N_17765,N_17723);
xnor U18462 (N_18462,N_17623,N_17673);
xnor U18463 (N_18463,N_17596,N_17606);
or U18464 (N_18464,N_17882,N_17619);
or U18465 (N_18465,N_17902,N_17799);
nand U18466 (N_18466,N_17600,N_17717);
xnor U18467 (N_18467,N_17705,N_17899);
and U18468 (N_18468,N_17747,N_17893);
or U18469 (N_18469,N_17780,N_17850);
xnor U18470 (N_18470,N_17902,N_17663);
or U18471 (N_18471,N_17814,N_17663);
or U18472 (N_18472,N_17893,N_17643);
nor U18473 (N_18473,N_17508,N_17926);
and U18474 (N_18474,N_17512,N_17661);
xnor U18475 (N_18475,N_17501,N_17536);
nand U18476 (N_18476,N_17882,N_17746);
or U18477 (N_18477,N_17794,N_17710);
xnor U18478 (N_18478,N_17501,N_17997);
nand U18479 (N_18479,N_17915,N_17658);
nor U18480 (N_18480,N_17609,N_17503);
or U18481 (N_18481,N_17973,N_17699);
or U18482 (N_18482,N_17503,N_17818);
or U18483 (N_18483,N_17757,N_17669);
and U18484 (N_18484,N_17599,N_17762);
and U18485 (N_18485,N_17930,N_17585);
xnor U18486 (N_18486,N_17730,N_17940);
and U18487 (N_18487,N_17952,N_17659);
nor U18488 (N_18488,N_17657,N_17855);
and U18489 (N_18489,N_17712,N_17895);
nand U18490 (N_18490,N_17859,N_17729);
nand U18491 (N_18491,N_17981,N_17939);
and U18492 (N_18492,N_17763,N_17608);
and U18493 (N_18493,N_17909,N_17727);
nand U18494 (N_18494,N_17590,N_17617);
nor U18495 (N_18495,N_17831,N_17647);
nor U18496 (N_18496,N_17642,N_17768);
and U18497 (N_18497,N_17951,N_17844);
xor U18498 (N_18498,N_17788,N_17808);
nor U18499 (N_18499,N_17788,N_17943);
nor U18500 (N_18500,N_18265,N_18223);
xor U18501 (N_18501,N_18288,N_18139);
nor U18502 (N_18502,N_18434,N_18266);
nand U18503 (N_18503,N_18394,N_18301);
xnor U18504 (N_18504,N_18171,N_18407);
or U18505 (N_18505,N_18308,N_18114);
or U18506 (N_18506,N_18340,N_18268);
nor U18507 (N_18507,N_18249,N_18406);
or U18508 (N_18508,N_18314,N_18059);
xor U18509 (N_18509,N_18413,N_18399);
xor U18510 (N_18510,N_18057,N_18339);
xnor U18511 (N_18511,N_18447,N_18263);
or U18512 (N_18512,N_18219,N_18190);
or U18513 (N_18513,N_18296,N_18346);
nand U18514 (N_18514,N_18078,N_18076);
nand U18515 (N_18515,N_18095,N_18155);
nand U18516 (N_18516,N_18361,N_18238);
nor U18517 (N_18517,N_18082,N_18294);
nor U18518 (N_18518,N_18018,N_18123);
or U18519 (N_18519,N_18388,N_18277);
and U18520 (N_18520,N_18485,N_18320);
xnor U18521 (N_18521,N_18408,N_18316);
nand U18522 (N_18522,N_18211,N_18183);
nand U18523 (N_18523,N_18271,N_18205);
nor U18524 (N_18524,N_18455,N_18027);
or U18525 (N_18525,N_18172,N_18003);
xor U18526 (N_18526,N_18317,N_18257);
nor U18527 (N_18527,N_18306,N_18477);
xor U18528 (N_18528,N_18479,N_18453);
or U18529 (N_18529,N_18198,N_18181);
nor U18530 (N_18530,N_18307,N_18116);
xor U18531 (N_18531,N_18375,N_18086);
or U18532 (N_18532,N_18430,N_18411);
and U18533 (N_18533,N_18440,N_18212);
xor U18534 (N_18534,N_18300,N_18298);
xnor U18535 (N_18535,N_18305,N_18460);
xnor U18536 (N_18536,N_18157,N_18169);
and U18537 (N_18537,N_18262,N_18229);
xor U18538 (N_18538,N_18044,N_18033);
or U18539 (N_18539,N_18063,N_18355);
or U18540 (N_18540,N_18309,N_18255);
and U18541 (N_18541,N_18213,N_18174);
xnor U18542 (N_18542,N_18292,N_18295);
and U18543 (N_18543,N_18079,N_18242);
nand U18544 (N_18544,N_18337,N_18387);
nor U18545 (N_18545,N_18378,N_18352);
nand U18546 (N_18546,N_18410,N_18454);
xnor U18547 (N_18547,N_18001,N_18083);
and U18548 (N_18548,N_18280,N_18336);
nand U18549 (N_18549,N_18208,N_18045);
and U18550 (N_18550,N_18445,N_18243);
or U18551 (N_18551,N_18210,N_18469);
xnor U18552 (N_18552,N_18285,N_18152);
xor U18553 (N_18553,N_18014,N_18096);
nand U18554 (N_18554,N_18207,N_18233);
or U18555 (N_18555,N_18290,N_18438);
and U18556 (N_18556,N_18144,N_18374);
nand U18557 (N_18557,N_18250,N_18237);
and U18558 (N_18558,N_18256,N_18429);
nand U18559 (N_18559,N_18269,N_18209);
nor U18560 (N_18560,N_18131,N_18273);
or U18561 (N_18561,N_18017,N_18103);
or U18562 (N_18562,N_18185,N_18244);
and U18563 (N_18563,N_18481,N_18088);
nor U18564 (N_18564,N_18357,N_18492);
xnor U18565 (N_18565,N_18145,N_18193);
and U18566 (N_18566,N_18239,N_18068);
nor U18567 (N_18567,N_18401,N_18071);
and U18568 (N_18568,N_18197,N_18302);
xor U18569 (N_18569,N_18052,N_18030);
nand U18570 (N_18570,N_18004,N_18313);
or U18571 (N_18571,N_18154,N_18436);
xor U18572 (N_18572,N_18498,N_18478);
xor U18573 (N_18573,N_18435,N_18090);
nor U18574 (N_18574,N_18377,N_18202);
and U18575 (N_18575,N_18457,N_18019);
or U18576 (N_18576,N_18113,N_18168);
nand U18577 (N_18577,N_18091,N_18372);
xor U18578 (N_18578,N_18136,N_18102);
nand U18579 (N_18579,N_18291,N_18234);
or U18580 (N_18580,N_18162,N_18267);
and U18581 (N_18581,N_18039,N_18452);
and U18582 (N_18582,N_18332,N_18140);
nor U18583 (N_18583,N_18343,N_18137);
and U18584 (N_18584,N_18367,N_18448);
xnor U18585 (N_18585,N_18393,N_18041);
xnor U18586 (N_18586,N_18177,N_18159);
nand U18587 (N_18587,N_18437,N_18247);
or U18588 (N_18588,N_18354,N_18390);
xnor U18589 (N_18589,N_18272,N_18466);
or U18590 (N_18590,N_18134,N_18442);
and U18591 (N_18591,N_18489,N_18077);
xnor U18592 (N_18592,N_18024,N_18356);
nand U18593 (N_18593,N_18335,N_18391);
nor U18594 (N_18594,N_18165,N_18389);
xor U18595 (N_18595,N_18328,N_18104);
xnor U18596 (N_18596,N_18164,N_18400);
or U18597 (N_18597,N_18409,N_18423);
xor U18598 (N_18598,N_18194,N_18147);
nand U18599 (N_18599,N_18376,N_18206);
and U18600 (N_18600,N_18381,N_18125);
and U18601 (N_18601,N_18473,N_18425);
xnor U18602 (N_18602,N_18111,N_18022);
xor U18603 (N_18603,N_18451,N_18065);
nand U18604 (N_18604,N_18135,N_18220);
and U18605 (N_18605,N_18258,N_18098);
xnor U18606 (N_18606,N_18215,N_18032);
xor U18607 (N_18607,N_18318,N_18126);
or U18608 (N_18608,N_18491,N_18184);
nor U18609 (N_18609,N_18276,N_18153);
nor U18610 (N_18610,N_18405,N_18297);
or U18611 (N_18611,N_18061,N_18311);
or U18612 (N_18612,N_18118,N_18497);
nor U18613 (N_18613,N_18225,N_18040);
and U18614 (N_18614,N_18443,N_18365);
and U18615 (N_18615,N_18251,N_18120);
or U18616 (N_18616,N_18055,N_18218);
nor U18617 (N_18617,N_18427,N_18494);
nor U18618 (N_18618,N_18087,N_18151);
nand U18619 (N_18619,N_18379,N_18331);
and U18620 (N_18620,N_18402,N_18025);
nand U18621 (N_18621,N_18037,N_18161);
or U18622 (N_18622,N_18128,N_18217);
nor U18623 (N_18623,N_18304,N_18428);
xnor U18624 (N_18624,N_18006,N_18124);
and U18625 (N_18625,N_18049,N_18461);
or U18626 (N_18626,N_18094,N_18468);
nand U18627 (N_18627,N_18338,N_18299);
nor U18628 (N_18628,N_18146,N_18048);
nor U18629 (N_18629,N_18488,N_18278);
xor U18630 (N_18630,N_18380,N_18284);
nand U18631 (N_18631,N_18382,N_18475);
and U18632 (N_18632,N_18010,N_18282);
nand U18633 (N_18633,N_18064,N_18450);
nor U18634 (N_18634,N_18397,N_18456);
nor U18635 (N_18635,N_18034,N_18241);
nor U18636 (N_18636,N_18362,N_18201);
nand U18637 (N_18637,N_18166,N_18035);
xnor U18638 (N_18638,N_18439,N_18227);
or U18639 (N_18639,N_18093,N_18395);
xnor U18640 (N_18640,N_18424,N_18031);
nand U18641 (N_18641,N_18175,N_18329);
xnor U18642 (N_18642,N_18149,N_18472);
and U18643 (N_18643,N_18353,N_18046);
or U18644 (N_18644,N_18349,N_18259);
xnor U18645 (N_18645,N_18279,N_18493);
nor U18646 (N_18646,N_18023,N_18188);
xor U18647 (N_18647,N_18287,N_18245);
and U18648 (N_18648,N_18345,N_18412);
nor U18649 (N_18649,N_18176,N_18254);
nor U18650 (N_18650,N_18444,N_18156);
and U18651 (N_18651,N_18417,N_18129);
and U18652 (N_18652,N_18016,N_18471);
nand U18653 (N_18653,N_18101,N_18084);
and U18654 (N_18654,N_18404,N_18289);
nor U18655 (N_18655,N_18270,N_18248);
or U18656 (N_18656,N_18363,N_18109);
xor U18657 (N_18657,N_18216,N_18369);
nor U18658 (N_18658,N_18420,N_18403);
nand U18659 (N_18659,N_18150,N_18105);
and U18660 (N_18660,N_18459,N_18026);
and U18661 (N_18661,N_18414,N_18119);
and U18662 (N_18662,N_18054,N_18187);
nand U18663 (N_18663,N_18275,N_18051);
and U18664 (N_18664,N_18013,N_18462);
xnor U18665 (N_18665,N_18143,N_18253);
and U18666 (N_18666,N_18323,N_18231);
or U18667 (N_18667,N_18224,N_18232);
and U18668 (N_18668,N_18246,N_18110);
xnor U18669 (N_18669,N_18195,N_18221);
nand U18670 (N_18670,N_18074,N_18163);
and U18671 (N_18671,N_18419,N_18008);
and U18672 (N_18672,N_18326,N_18100);
nand U18673 (N_18673,N_18431,N_18333);
nor U18674 (N_18674,N_18396,N_18484);
or U18675 (N_18675,N_18069,N_18073);
or U18676 (N_18676,N_18312,N_18107);
nor U18677 (N_18677,N_18458,N_18056);
xnor U18678 (N_18678,N_18315,N_18228);
or U18679 (N_18679,N_18321,N_18133);
nand U18680 (N_18680,N_18366,N_18483);
and U18681 (N_18681,N_18348,N_18286);
xnor U18682 (N_18682,N_18204,N_18189);
nand U18683 (N_18683,N_18368,N_18415);
or U18684 (N_18684,N_18421,N_18132);
or U18685 (N_18685,N_18303,N_18260);
xnor U18686 (N_18686,N_18236,N_18050);
nand U18687 (N_18687,N_18020,N_18196);
or U18688 (N_18688,N_18112,N_18433);
nor U18689 (N_18689,N_18342,N_18099);
and U18690 (N_18690,N_18179,N_18138);
nor U18691 (N_18691,N_18170,N_18191);
xor U18692 (N_18692,N_18474,N_18000);
and U18693 (N_18693,N_18180,N_18097);
or U18694 (N_18694,N_18386,N_18038);
xor U18695 (N_18695,N_18344,N_18067);
or U18696 (N_18696,N_18127,N_18130);
nand U18697 (N_18697,N_18058,N_18036);
nor U18698 (N_18698,N_18160,N_18085);
or U18699 (N_18699,N_18293,N_18106);
or U18700 (N_18700,N_18360,N_18005);
xnor U18701 (N_18701,N_18080,N_18226);
xnor U18702 (N_18702,N_18072,N_18370);
or U18703 (N_18703,N_18482,N_18319);
nand U18704 (N_18704,N_18141,N_18476);
and U18705 (N_18705,N_18384,N_18383);
nor U18706 (N_18706,N_18015,N_18062);
or U18707 (N_18707,N_18350,N_18214);
or U18708 (N_18708,N_18261,N_18392);
or U18709 (N_18709,N_18398,N_18324);
nor U18710 (N_18710,N_18449,N_18446);
nand U18711 (N_18711,N_18199,N_18499);
xor U18712 (N_18712,N_18089,N_18182);
nand U18713 (N_18713,N_18115,N_18117);
nand U18714 (N_18714,N_18042,N_18178);
xnor U18715 (N_18715,N_18167,N_18465);
xnor U18716 (N_18716,N_18330,N_18230);
nor U18717 (N_18717,N_18148,N_18463);
xor U18718 (N_18718,N_18371,N_18490);
or U18719 (N_18719,N_18487,N_18347);
and U18720 (N_18720,N_18235,N_18060);
nor U18721 (N_18721,N_18364,N_18467);
nand U18722 (N_18722,N_18108,N_18047);
nor U18723 (N_18723,N_18358,N_18200);
and U18724 (N_18724,N_18173,N_18252);
nor U18725 (N_18725,N_18310,N_18441);
or U18726 (N_18726,N_18418,N_18327);
xor U18727 (N_18727,N_18496,N_18009);
nor U18728 (N_18728,N_18341,N_18203);
and U18729 (N_18729,N_18385,N_18142);
nor U18730 (N_18730,N_18186,N_18066);
xnor U18731 (N_18731,N_18495,N_18432);
xnor U18732 (N_18732,N_18158,N_18426);
or U18733 (N_18733,N_18264,N_18002);
or U18734 (N_18734,N_18021,N_18351);
nor U18735 (N_18735,N_18029,N_18070);
nand U18736 (N_18736,N_18192,N_18416);
and U18737 (N_18737,N_18422,N_18464);
nor U18738 (N_18738,N_18012,N_18281);
nand U18739 (N_18739,N_18373,N_18322);
nand U18740 (N_18740,N_18480,N_18011);
nand U18741 (N_18741,N_18359,N_18053);
and U18742 (N_18742,N_18007,N_18122);
or U18743 (N_18743,N_18334,N_18274);
nor U18744 (N_18744,N_18092,N_18043);
nand U18745 (N_18745,N_18028,N_18486);
nand U18746 (N_18746,N_18121,N_18240);
nor U18747 (N_18747,N_18075,N_18470);
nor U18748 (N_18748,N_18283,N_18222);
nand U18749 (N_18749,N_18081,N_18325);
nand U18750 (N_18750,N_18442,N_18315);
nand U18751 (N_18751,N_18433,N_18239);
xor U18752 (N_18752,N_18354,N_18224);
nand U18753 (N_18753,N_18061,N_18330);
nor U18754 (N_18754,N_18114,N_18415);
or U18755 (N_18755,N_18152,N_18323);
nor U18756 (N_18756,N_18132,N_18346);
and U18757 (N_18757,N_18426,N_18342);
or U18758 (N_18758,N_18419,N_18473);
xnor U18759 (N_18759,N_18236,N_18000);
nor U18760 (N_18760,N_18267,N_18195);
or U18761 (N_18761,N_18200,N_18058);
nor U18762 (N_18762,N_18010,N_18352);
xnor U18763 (N_18763,N_18180,N_18473);
nand U18764 (N_18764,N_18396,N_18336);
nor U18765 (N_18765,N_18464,N_18065);
and U18766 (N_18766,N_18187,N_18042);
and U18767 (N_18767,N_18166,N_18496);
nand U18768 (N_18768,N_18067,N_18096);
nor U18769 (N_18769,N_18155,N_18415);
nand U18770 (N_18770,N_18474,N_18149);
and U18771 (N_18771,N_18070,N_18183);
nand U18772 (N_18772,N_18030,N_18218);
nor U18773 (N_18773,N_18099,N_18374);
nor U18774 (N_18774,N_18413,N_18194);
and U18775 (N_18775,N_18251,N_18025);
or U18776 (N_18776,N_18203,N_18408);
and U18777 (N_18777,N_18179,N_18210);
and U18778 (N_18778,N_18194,N_18123);
xor U18779 (N_18779,N_18252,N_18021);
and U18780 (N_18780,N_18380,N_18212);
xnor U18781 (N_18781,N_18462,N_18036);
xnor U18782 (N_18782,N_18312,N_18118);
or U18783 (N_18783,N_18416,N_18003);
and U18784 (N_18784,N_18457,N_18178);
and U18785 (N_18785,N_18410,N_18484);
and U18786 (N_18786,N_18283,N_18321);
and U18787 (N_18787,N_18196,N_18398);
and U18788 (N_18788,N_18263,N_18494);
and U18789 (N_18789,N_18470,N_18137);
xnor U18790 (N_18790,N_18472,N_18137);
nand U18791 (N_18791,N_18043,N_18179);
or U18792 (N_18792,N_18078,N_18015);
nor U18793 (N_18793,N_18266,N_18173);
or U18794 (N_18794,N_18198,N_18171);
xor U18795 (N_18795,N_18087,N_18365);
xnor U18796 (N_18796,N_18296,N_18078);
nor U18797 (N_18797,N_18005,N_18041);
nand U18798 (N_18798,N_18055,N_18174);
xnor U18799 (N_18799,N_18473,N_18024);
and U18800 (N_18800,N_18469,N_18326);
xor U18801 (N_18801,N_18232,N_18025);
nor U18802 (N_18802,N_18223,N_18390);
nand U18803 (N_18803,N_18110,N_18464);
nor U18804 (N_18804,N_18016,N_18126);
or U18805 (N_18805,N_18498,N_18442);
xor U18806 (N_18806,N_18289,N_18234);
and U18807 (N_18807,N_18063,N_18357);
xnor U18808 (N_18808,N_18006,N_18180);
xnor U18809 (N_18809,N_18409,N_18297);
nor U18810 (N_18810,N_18363,N_18441);
nor U18811 (N_18811,N_18211,N_18458);
nor U18812 (N_18812,N_18301,N_18131);
or U18813 (N_18813,N_18367,N_18157);
nor U18814 (N_18814,N_18021,N_18470);
or U18815 (N_18815,N_18119,N_18134);
nor U18816 (N_18816,N_18001,N_18455);
nor U18817 (N_18817,N_18390,N_18496);
and U18818 (N_18818,N_18081,N_18342);
nand U18819 (N_18819,N_18029,N_18078);
nor U18820 (N_18820,N_18261,N_18004);
nor U18821 (N_18821,N_18003,N_18118);
or U18822 (N_18822,N_18403,N_18461);
nor U18823 (N_18823,N_18330,N_18371);
xor U18824 (N_18824,N_18437,N_18088);
or U18825 (N_18825,N_18109,N_18226);
nand U18826 (N_18826,N_18305,N_18359);
nand U18827 (N_18827,N_18020,N_18499);
nand U18828 (N_18828,N_18084,N_18485);
or U18829 (N_18829,N_18051,N_18401);
or U18830 (N_18830,N_18155,N_18310);
xnor U18831 (N_18831,N_18143,N_18309);
and U18832 (N_18832,N_18498,N_18161);
xor U18833 (N_18833,N_18001,N_18032);
and U18834 (N_18834,N_18027,N_18369);
nand U18835 (N_18835,N_18201,N_18456);
xnor U18836 (N_18836,N_18001,N_18332);
nand U18837 (N_18837,N_18330,N_18235);
or U18838 (N_18838,N_18389,N_18444);
xnor U18839 (N_18839,N_18104,N_18087);
or U18840 (N_18840,N_18284,N_18424);
nor U18841 (N_18841,N_18378,N_18270);
nand U18842 (N_18842,N_18404,N_18217);
or U18843 (N_18843,N_18487,N_18299);
nand U18844 (N_18844,N_18349,N_18268);
or U18845 (N_18845,N_18120,N_18190);
xnor U18846 (N_18846,N_18176,N_18497);
nand U18847 (N_18847,N_18091,N_18106);
and U18848 (N_18848,N_18465,N_18303);
xnor U18849 (N_18849,N_18046,N_18217);
or U18850 (N_18850,N_18347,N_18361);
xor U18851 (N_18851,N_18342,N_18451);
and U18852 (N_18852,N_18120,N_18062);
or U18853 (N_18853,N_18405,N_18421);
or U18854 (N_18854,N_18273,N_18067);
nor U18855 (N_18855,N_18040,N_18267);
nor U18856 (N_18856,N_18035,N_18423);
nand U18857 (N_18857,N_18180,N_18125);
or U18858 (N_18858,N_18191,N_18130);
or U18859 (N_18859,N_18038,N_18456);
and U18860 (N_18860,N_18290,N_18384);
or U18861 (N_18861,N_18023,N_18129);
xnor U18862 (N_18862,N_18464,N_18458);
nor U18863 (N_18863,N_18071,N_18091);
nand U18864 (N_18864,N_18046,N_18056);
nor U18865 (N_18865,N_18069,N_18262);
nand U18866 (N_18866,N_18279,N_18007);
nor U18867 (N_18867,N_18224,N_18459);
nand U18868 (N_18868,N_18444,N_18303);
nand U18869 (N_18869,N_18103,N_18247);
and U18870 (N_18870,N_18282,N_18151);
nand U18871 (N_18871,N_18253,N_18250);
nor U18872 (N_18872,N_18477,N_18277);
and U18873 (N_18873,N_18381,N_18428);
xor U18874 (N_18874,N_18160,N_18246);
nor U18875 (N_18875,N_18135,N_18168);
or U18876 (N_18876,N_18219,N_18263);
nor U18877 (N_18877,N_18453,N_18324);
and U18878 (N_18878,N_18452,N_18431);
nor U18879 (N_18879,N_18381,N_18007);
and U18880 (N_18880,N_18232,N_18311);
nor U18881 (N_18881,N_18159,N_18196);
nand U18882 (N_18882,N_18498,N_18430);
xnor U18883 (N_18883,N_18297,N_18106);
and U18884 (N_18884,N_18081,N_18272);
nor U18885 (N_18885,N_18024,N_18160);
xnor U18886 (N_18886,N_18095,N_18179);
or U18887 (N_18887,N_18305,N_18289);
nor U18888 (N_18888,N_18088,N_18350);
and U18889 (N_18889,N_18491,N_18139);
xnor U18890 (N_18890,N_18068,N_18098);
nor U18891 (N_18891,N_18332,N_18374);
nor U18892 (N_18892,N_18296,N_18487);
nand U18893 (N_18893,N_18252,N_18387);
xor U18894 (N_18894,N_18077,N_18487);
nor U18895 (N_18895,N_18422,N_18107);
or U18896 (N_18896,N_18128,N_18154);
or U18897 (N_18897,N_18120,N_18339);
or U18898 (N_18898,N_18208,N_18294);
xnor U18899 (N_18899,N_18138,N_18326);
and U18900 (N_18900,N_18373,N_18424);
xnor U18901 (N_18901,N_18368,N_18126);
and U18902 (N_18902,N_18304,N_18311);
xnor U18903 (N_18903,N_18430,N_18246);
and U18904 (N_18904,N_18233,N_18121);
xor U18905 (N_18905,N_18076,N_18391);
nor U18906 (N_18906,N_18384,N_18366);
xor U18907 (N_18907,N_18032,N_18007);
nand U18908 (N_18908,N_18004,N_18021);
or U18909 (N_18909,N_18436,N_18101);
or U18910 (N_18910,N_18374,N_18183);
nor U18911 (N_18911,N_18044,N_18007);
nand U18912 (N_18912,N_18114,N_18148);
nor U18913 (N_18913,N_18144,N_18266);
and U18914 (N_18914,N_18342,N_18109);
xor U18915 (N_18915,N_18202,N_18077);
nand U18916 (N_18916,N_18206,N_18381);
xor U18917 (N_18917,N_18003,N_18224);
and U18918 (N_18918,N_18235,N_18025);
or U18919 (N_18919,N_18082,N_18430);
xor U18920 (N_18920,N_18321,N_18427);
nor U18921 (N_18921,N_18185,N_18409);
nor U18922 (N_18922,N_18411,N_18036);
and U18923 (N_18923,N_18334,N_18394);
and U18924 (N_18924,N_18459,N_18210);
nor U18925 (N_18925,N_18225,N_18367);
nand U18926 (N_18926,N_18454,N_18386);
or U18927 (N_18927,N_18015,N_18012);
or U18928 (N_18928,N_18450,N_18141);
nor U18929 (N_18929,N_18264,N_18416);
and U18930 (N_18930,N_18371,N_18179);
or U18931 (N_18931,N_18381,N_18217);
nand U18932 (N_18932,N_18339,N_18353);
or U18933 (N_18933,N_18022,N_18396);
and U18934 (N_18934,N_18285,N_18058);
or U18935 (N_18935,N_18498,N_18116);
nor U18936 (N_18936,N_18346,N_18456);
nand U18937 (N_18937,N_18237,N_18071);
nor U18938 (N_18938,N_18256,N_18023);
or U18939 (N_18939,N_18363,N_18028);
and U18940 (N_18940,N_18061,N_18046);
nor U18941 (N_18941,N_18258,N_18084);
xor U18942 (N_18942,N_18186,N_18159);
and U18943 (N_18943,N_18463,N_18287);
or U18944 (N_18944,N_18276,N_18335);
nand U18945 (N_18945,N_18068,N_18148);
xnor U18946 (N_18946,N_18497,N_18405);
nor U18947 (N_18947,N_18312,N_18052);
or U18948 (N_18948,N_18087,N_18359);
nor U18949 (N_18949,N_18352,N_18274);
or U18950 (N_18950,N_18457,N_18173);
xor U18951 (N_18951,N_18101,N_18374);
or U18952 (N_18952,N_18128,N_18468);
nor U18953 (N_18953,N_18385,N_18068);
nor U18954 (N_18954,N_18205,N_18156);
nand U18955 (N_18955,N_18162,N_18399);
xnor U18956 (N_18956,N_18437,N_18192);
and U18957 (N_18957,N_18340,N_18025);
or U18958 (N_18958,N_18067,N_18289);
xnor U18959 (N_18959,N_18426,N_18210);
nor U18960 (N_18960,N_18283,N_18037);
or U18961 (N_18961,N_18226,N_18105);
xnor U18962 (N_18962,N_18107,N_18292);
or U18963 (N_18963,N_18380,N_18318);
nand U18964 (N_18964,N_18390,N_18113);
nor U18965 (N_18965,N_18072,N_18055);
or U18966 (N_18966,N_18322,N_18126);
xnor U18967 (N_18967,N_18386,N_18096);
and U18968 (N_18968,N_18488,N_18481);
or U18969 (N_18969,N_18392,N_18264);
or U18970 (N_18970,N_18168,N_18008);
nand U18971 (N_18971,N_18397,N_18046);
and U18972 (N_18972,N_18293,N_18214);
or U18973 (N_18973,N_18337,N_18409);
and U18974 (N_18974,N_18016,N_18342);
nand U18975 (N_18975,N_18111,N_18495);
and U18976 (N_18976,N_18060,N_18069);
xnor U18977 (N_18977,N_18325,N_18035);
nand U18978 (N_18978,N_18121,N_18355);
xor U18979 (N_18979,N_18188,N_18211);
nand U18980 (N_18980,N_18464,N_18221);
and U18981 (N_18981,N_18255,N_18231);
or U18982 (N_18982,N_18051,N_18145);
xor U18983 (N_18983,N_18303,N_18033);
xor U18984 (N_18984,N_18177,N_18058);
nor U18985 (N_18985,N_18229,N_18274);
xnor U18986 (N_18986,N_18054,N_18062);
nor U18987 (N_18987,N_18003,N_18200);
and U18988 (N_18988,N_18329,N_18481);
xor U18989 (N_18989,N_18496,N_18003);
nand U18990 (N_18990,N_18147,N_18325);
xnor U18991 (N_18991,N_18354,N_18360);
or U18992 (N_18992,N_18186,N_18241);
nor U18993 (N_18993,N_18395,N_18469);
or U18994 (N_18994,N_18385,N_18196);
or U18995 (N_18995,N_18400,N_18044);
xor U18996 (N_18996,N_18329,N_18338);
nand U18997 (N_18997,N_18401,N_18337);
nor U18998 (N_18998,N_18206,N_18093);
nand U18999 (N_18999,N_18408,N_18286);
nor U19000 (N_19000,N_18974,N_18788);
or U19001 (N_19001,N_18809,N_18530);
and U19002 (N_19002,N_18818,N_18537);
and U19003 (N_19003,N_18825,N_18538);
or U19004 (N_19004,N_18900,N_18649);
nor U19005 (N_19005,N_18815,N_18601);
nor U19006 (N_19006,N_18557,N_18946);
nand U19007 (N_19007,N_18830,N_18618);
or U19008 (N_19008,N_18858,N_18515);
xor U19009 (N_19009,N_18510,N_18984);
nor U19010 (N_19010,N_18912,N_18624);
nor U19011 (N_19011,N_18636,N_18550);
xnor U19012 (N_19012,N_18954,N_18747);
and U19013 (N_19013,N_18727,N_18643);
or U19014 (N_19014,N_18591,N_18993);
nor U19015 (N_19015,N_18603,N_18542);
and U19016 (N_19016,N_18936,N_18867);
xnor U19017 (N_19017,N_18876,N_18926);
xnor U19018 (N_19018,N_18855,N_18857);
xnor U19019 (N_19019,N_18764,N_18999);
and U19020 (N_19020,N_18918,N_18774);
and U19021 (N_19021,N_18890,N_18715);
xnor U19022 (N_19022,N_18713,N_18901);
and U19023 (N_19023,N_18579,N_18821);
nand U19024 (N_19024,N_18506,N_18932);
xor U19025 (N_19025,N_18997,N_18634);
or U19026 (N_19026,N_18808,N_18767);
xor U19027 (N_19027,N_18752,N_18578);
nor U19028 (N_19028,N_18728,N_18760);
and U19029 (N_19029,N_18834,N_18735);
nor U19030 (N_19030,N_18742,N_18968);
and U19031 (N_19031,N_18991,N_18902);
nor U19032 (N_19032,N_18642,N_18672);
nand U19033 (N_19033,N_18629,N_18560);
nand U19034 (N_19034,N_18721,N_18934);
nand U19035 (N_19035,N_18921,N_18535);
and U19036 (N_19036,N_18706,N_18920);
nor U19037 (N_19037,N_18688,N_18869);
xnor U19038 (N_19038,N_18667,N_18776);
nand U19039 (N_19039,N_18651,N_18754);
nand U19040 (N_19040,N_18574,N_18518);
xnor U19041 (N_19041,N_18609,N_18543);
or U19042 (N_19042,N_18803,N_18816);
nor U19043 (N_19043,N_18546,N_18948);
nand U19044 (N_19044,N_18689,N_18547);
xnor U19045 (N_19045,N_18782,N_18888);
or U19046 (N_19046,N_18973,N_18568);
and U19047 (N_19047,N_18566,N_18509);
nand U19048 (N_19048,N_18870,N_18795);
nor U19049 (N_19049,N_18873,N_18982);
or U19050 (N_19050,N_18909,N_18573);
or U19051 (N_19051,N_18940,N_18503);
nand U19052 (N_19052,N_18963,N_18887);
or U19053 (N_19053,N_18925,N_18520);
nor U19054 (N_19054,N_18981,N_18919);
and U19055 (N_19055,N_18726,N_18511);
nand U19056 (N_19056,N_18790,N_18734);
or U19057 (N_19057,N_18617,N_18710);
nor U19058 (N_19058,N_18598,N_18614);
nor U19059 (N_19059,N_18894,N_18584);
or U19060 (N_19060,N_18580,N_18517);
nor U19061 (N_19061,N_18720,N_18625);
xor U19062 (N_19062,N_18635,N_18645);
xnor U19063 (N_19063,N_18526,N_18971);
or U19064 (N_19064,N_18949,N_18756);
nand U19065 (N_19065,N_18836,N_18928);
nor U19066 (N_19066,N_18620,N_18794);
nand U19067 (N_19067,N_18929,N_18978);
nor U19068 (N_19068,N_18707,N_18632);
xor U19069 (N_19069,N_18570,N_18783);
and U19070 (N_19070,N_18831,N_18504);
nand U19071 (N_19071,N_18804,N_18581);
xnor U19072 (N_19072,N_18759,N_18676);
nor U19073 (N_19073,N_18505,N_18915);
xor U19074 (N_19074,N_18866,N_18730);
xor U19075 (N_19075,N_18668,N_18988);
xnor U19076 (N_19076,N_18844,N_18813);
and U19077 (N_19077,N_18679,N_18883);
or U19078 (N_19078,N_18576,N_18608);
xnor U19079 (N_19079,N_18619,N_18874);
nor U19080 (N_19080,N_18702,N_18739);
xor U19081 (N_19081,N_18701,N_18910);
or U19082 (N_19082,N_18663,N_18746);
or U19083 (N_19083,N_18621,N_18588);
or U19084 (N_19084,N_18558,N_18716);
xor U19085 (N_19085,N_18605,N_18514);
nand U19086 (N_19086,N_18757,N_18881);
or U19087 (N_19087,N_18811,N_18638);
nand U19088 (N_19088,N_18744,N_18650);
and U19089 (N_19089,N_18678,N_18951);
nor U19090 (N_19090,N_18889,N_18938);
xor U19091 (N_19091,N_18563,N_18849);
nand U19092 (N_19092,N_18556,N_18812);
and U19093 (N_19093,N_18906,N_18914);
nor U19094 (N_19094,N_18630,N_18554);
nor U19095 (N_19095,N_18930,N_18741);
and U19096 (N_19096,N_18805,N_18819);
nand U19097 (N_19097,N_18523,N_18541);
nor U19098 (N_19098,N_18913,N_18772);
nand U19099 (N_19099,N_18718,N_18972);
nor U19100 (N_19100,N_18512,N_18690);
nor U19101 (N_19101,N_18736,N_18685);
nor U19102 (N_19102,N_18989,N_18841);
nor U19103 (N_19103,N_18545,N_18648);
and U19104 (N_19104,N_18878,N_18674);
nand U19105 (N_19105,N_18564,N_18691);
and U19106 (N_19106,N_18501,N_18923);
nand U19107 (N_19107,N_18755,N_18846);
xnor U19108 (N_19108,N_18937,N_18641);
and U19109 (N_19109,N_18778,N_18786);
and U19110 (N_19110,N_18848,N_18687);
nand U19111 (N_19111,N_18959,N_18749);
or U19112 (N_19112,N_18665,N_18839);
and U19113 (N_19113,N_18548,N_18737);
nand U19114 (N_19114,N_18986,N_18507);
or U19115 (N_19115,N_18670,N_18571);
nor U19116 (N_19116,N_18994,N_18750);
nand U19117 (N_19117,N_18891,N_18696);
or U19118 (N_19118,N_18657,N_18555);
nor U19119 (N_19119,N_18673,N_18582);
nand U19120 (N_19120,N_18704,N_18644);
xnor U19121 (N_19121,N_18861,N_18882);
and U19122 (N_19122,N_18899,N_18765);
nand U19123 (N_19123,N_18964,N_18904);
xnor U19124 (N_19124,N_18800,N_18723);
nor U19125 (N_19125,N_18793,N_18682);
and U19126 (N_19126,N_18758,N_18561);
nand U19127 (N_19127,N_18748,N_18513);
xnor U19128 (N_19128,N_18733,N_18500);
xnor U19129 (N_19129,N_18985,N_18864);
and U19130 (N_19130,N_18699,N_18751);
nand U19131 (N_19131,N_18753,N_18787);
xor U19132 (N_19132,N_18549,N_18528);
and U19133 (N_19133,N_18851,N_18669);
nor U19134 (N_19134,N_18616,N_18895);
xnor U19135 (N_19135,N_18875,N_18762);
and U19136 (N_19136,N_18828,N_18911);
nor U19137 (N_19137,N_18955,N_18935);
nand U19138 (N_19138,N_18536,N_18656);
or U19139 (N_19139,N_18658,N_18990);
and U19140 (N_19140,N_18802,N_18586);
and U19141 (N_19141,N_18987,N_18960);
nor U19142 (N_19142,N_18627,N_18666);
nor U19143 (N_19143,N_18975,N_18664);
nand U19144 (N_19144,N_18976,N_18810);
xnor U19145 (N_19145,N_18850,N_18797);
and U19146 (N_19146,N_18695,N_18612);
xnor U19147 (N_19147,N_18943,N_18950);
xnor U19148 (N_19148,N_18969,N_18933);
nor U19149 (N_19149,N_18847,N_18686);
xnor U19150 (N_19150,N_18525,N_18768);
xor U19151 (N_19151,N_18607,N_18725);
or U19152 (N_19152,N_18789,N_18908);
xor U19153 (N_19153,N_18771,N_18958);
and U19154 (N_19154,N_18952,N_18660);
or U19155 (N_19155,N_18917,N_18653);
and U19156 (N_19156,N_18508,N_18709);
nand U19157 (N_19157,N_18631,N_18903);
and U19158 (N_19158,N_18927,N_18626);
and U19159 (N_19159,N_18872,N_18845);
nand U19160 (N_19160,N_18569,N_18532);
or U19161 (N_19161,N_18521,N_18965);
nand U19162 (N_19162,N_18662,N_18559);
nand U19163 (N_19163,N_18613,N_18792);
nand U19164 (N_19164,N_18639,N_18977);
xnor U19165 (N_19165,N_18594,N_18731);
and U19166 (N_19166,N_18675,N_18529);
nand U19167 (N_19167,N_18995,N_18807);
xnor U19168 (N_19168,N_18829,N_18945);
or U19169 (N_19169,N_18898,N_18743);
xnor U19170 (N_19170,N_18646,N_18777);
nor U19171 (N_19171,N_18962,N_18738);
nor U19172 (N_19172,N_18708,N_18732);
and U19173 (N_19173,N_18833,N_18589);
or U19174 (N_19174,N_18996,N_18865);
nand U19175 (N_19175,N_18860,N_18775);
nand U19176 (N_19176,N_18814,N_18597);
or U19177 (N_19177,N_18843,N_18681);
nor U19178 (N_19178,N_18717,N_18637);
xor U19179 (N_19179,N_18961,N_18966);
and U19180 (N_19180,N_18583,N_18533);
nor U19181 (N_19181,N_18868,N_18892);
nor U19182 (N_19182,N_18827,N_18593);
or U19183 (N_19183,N_18823,N_18553);
xor U19184 (N_19184,N_18980,N_18859);
xnor U19185 (N_19185,N_18697,N_18552);
and U19186 (N_19186,N_18628,N_18798);
nor U19187 (N_19187,N_18692,N_18893);
xnor U19188 (N_19188,N_18539,N_18516);
nor U19189 (N_19189,N_18998,N_18842);
or U19190 (N_19190,N_18779,N_18801);
and U19191 (N_19191,N_18595,N_18886);
nand U19192 (N_19192,N_18837,N_18585);
or U19193 (N_19193,N_18785,N_18654);
nor U19194 (N_19194,N_18773,N_18745);
or U19195 (N_19195,N_18540,N_18820);
nor U19196 (N_19196,N_18769,N_18680);
and U19197 (N_19197,N_18712,N_18729);
nand U19198 (N_19198,N_18652,N_18791);
and U19199 (N_19199,N_18916,N_18572);
or U19200 (N_19200,N_18711,N_18602);
nand U19201 (N_19201,N_18544,N_18615);
xnor U19202 (N_19202,N_18822,N_18806);
and U19203 (N_19203,N_18611,N_18905);
nand U19204 (N_19204,N_18897,N_18562);
nor U19205 (N_19205,N_18939,N_18885);
and U19206 (N_19206,N_18575,N_18524);
xnor U19207 (N_19207,N_18671,N_18796);
xor U19208 (N_19208,N_18719,N_18655);
xnor U19209 (N_19209,N_18519,N_18684);
and U19210 (N_19210,N_18931,N_18714);
nor U19211 (N_19211,N_18817,N_18884);
nor U19212 (N_19212,N_18502,N_18979);
xnor U19213 (N_19213,N_18677,N_18592);
nor U19214 (N_19214,N_18838,N_18703);
nand U19215 (N_19215,N_18832,N_18871);
or U19216 (N_19216,N_18683,N_18659);
and U19217 (N_19217,N_18862,N_18610);
and U19218 (N_19218,N_18770,N_18606);
xor U19219 (N_19219,N_18761,N_18600);
and U19220 (N_19220,N_18922,N_18599);
and U19221 (N_19221,N_18693,N_18835);
or U19222 (N_19222,N_18880,N_18863);
nor U19223 (N_19223,N_18970,N_18766);
and U19224 (N_19224,N_18947,N_18824);
or U19225 (N_19225,N_18907,N_18854);
nand U19226 (N_19226,N_18698,N_18879);
xnor U19227 (N_19227,N_18577,N_18781);
and U19228 (N_19228,N_18622,N_18700);
or U19229 (N_19229,N_18694,N_18780);
xnor U19230 (N_19230,N_18992,N_18740);
and U19231 (N_19231,N_18942,N_18522);
or U19232 (N_19232,N_18840,N_18590);
xnor U19233 (N_19233,N_18705,N_18640);
and U19234 (N_19234,N_18944,N_18567);
xnor U19235 (N_19235,N_18956,N_18647);
xnor U19236 (N_19236,N_18527,N_18941);
nor U19237 (N_19237,N_18877,N_18784);
or U19238 (N_19238,N_18633,N_18763);
xnor U19239 (N_19239,N_18953,N_18551);
and U19240 (N_19240,N_18604,N_18896);
and U19241 (N_19241,N_18853,N_18799);
xor U19242 (N_19242,N_18983,N_18856);
xnor U19243 (N_19243,N_18957,N_18661);
and U19244 (N_19244,N_18826,N_18596);
nor U19245 (N_19245,N_18852,N_18967);
nand U19246 (N_19246,N_18722,N_18587);
xor U19247 (N_19247,N_18924,N_18565);
and U19248 (N_19248,N_18534,N_18531);
or U19249 (N_19249,N_18623,N_18724);
xor U19250 (N_19250,N_18637,N_18716);
or U19251 (N_19251,N_18684,N_18663);
nor U19252 (N_19252,N_18917,N_18856);
and U19253 (N_19253,N_18839,N_18941);
and U19254 (N_19254,N_18640,N_18950);
nand U19255 (N_19255,N_18751,N_18642);
or U19256 (N_19256,N_18543,N_18843);
nor U19257 (N_19257,N_18637,N_18625);
nand U19258 (N_19258,N_18716,N_18675);
nand U19259 (N_19259,N_18719,N_18630);
or U19260 (N_19260,N_18504,N_18512);
nor U19261 (N_19261,N_18577,N_18950);
nor U19262 (N_19262,N_18537,N_18556);
nand U19263 (N_19263,N_18880,N_18747);
nand U19264 (N_19264,N_18893,N_18712);
nand U19265 (N_19265,N_18977,N_18868);
nor U19266 (N_19266,N_18940,N_18864);
nand U19267 (N_19267,N_18795,N_18591);
xor U19268 (N_19268,N_18878,N_18857);
nand U19269 (N_19269,N_18579,N_18855);
xnor U19270 (N_19270,N_18689,N_18631);
nand U19271 (N_19271,N_18669,N_18821);
xnor U19272 (N_19272,N_18600,N_18644);
or U19273 (N_19273,N_18584,N_18644);
nor U19274 (N_19274,N_18955,N_18695);
nor U19275 (N_19275,N_18586,N_18834);
and U19276 (N_19276,N_18874,N_18567);
nand U19277 (N_19277,N_18522,N_18763);
and U19278 (N_19278,N_18836,N_18856);
and U19279 (N_19279,N_18567,N_18790);
xnor U19280 (N_19280,N_18993,N_18724);
nand U19281 (N_19281,N_18753,N_18711);
and U19282 (N_19282,N_18997,N_18580);
and U19283 (N_19283,N_18665,N_18522);
xor U19284 (N_19284,N_18611,N_18938);
nor U19285 (N_19285,N_18501,N_18643);
and U19286 (N_19286,N_18831,N_18950);
nand U19287 (N_19287,N_18870,N_18960);
or U19288 (N_19288,N_18955,N_18580);
nand U19289 (N_19289,N_18958,N_18624);
xor U19290 (N_19290,N_18508,N_18561);
or U19291 (N_19291,N_18633,N_18893);
nand U19292 (N_19292,N_18694,N_18851);
and U19293 (N_19293,N_18688,N_18669);
and U19294 (N_19294,N_18682,N_18992);
xor U19295 (N_19295,N_18601,N_18582);
nand U19296 (N_19296,N_18874,N_18528);
or U19297 (N_19297,N_18734,N_18732);
xnor U19298 (N_19298,N_18947,N_18560);
nand U19299 (N_19299,N_18893,N_18971);
nand U19300 (N_19300,N_18790,N_18908);
and U19301 (N_19301,N_18774,N_18975);
nor U19302 (N_19302,N_18887,N_18836);
nor U19303 (N_19303,N_18963,N_18582);
and U19304 (N_19304,N_18522,N_18946);
xnor U19305 (N_19305,N_18885,N_18956);
nor U19306 (N_19306,N_18929,N_18641);
xor U19307 (N_19307,N_18832,N_18973);
and U19308 (N_19308,N_18570,N_18828);
xnor U19309 (N_19309,N_18859,N_18685);
or U19310 (N_19310,N_18758,N_18975);
xnor U19311 (N_19311,N_18947,N_18981);
and U19312 (N_19312,N_18730,N_18778);
xor U19313 (N_19313,N_18872,N_18535);
and U19314 (N_19314,N_18695,N_18771);
nand U19315 (N_19315,N_18793,N_18713);
or U19316 (N_19316,N_18822,N_18676);
nor U19317 (N_19317,N_18867,N_18695);
and U19318 (N_19318,N_18822,N_18680);
nand U19319 (N_19319,N_18941,N_18985);
and U19320 (N_19320,N_18835,N_18786);
and U19321 (N_19321,N_18968,N_18779);
and U19322 (N_19322,N_18922,N_18937);
and U19323 (N_19323,N_18624,N_18771);
nand U19324 (N_19324,N_18674,N_18805);
nor U19325 (N_19325,N_18652,N_18757);
nand U19326 (N_19326,N_18518,N_18780);
nor U19327 (N_19327,N_18838,N_18875);
nand U19328 (N_19328,N_18681,N_18724);
or U19329 (N_19329,N_18861,N_18919);
nand U19330 (N_19330,N_18834,N_18580);
nand U19331 (N_19331,N_18994,N_18533);
and U19332 (N_19332,N_18955,N_18813);
nand U19333 (N_19333,N_18602,N_18534);
nor U19334 (N_19334,N_18552,N_18627);
nand U19335 (N_19335,N_18594,N_18814);
nor U19336 (N_19336,N_18701,N_18717);
xnor U19337 (N_19337,N_18903,N_18645);
nand U19338 (N_19338,N_18567,N_18658);
and U19339 (N_19339,N_18934,N_18981);
nor U19340 (N_19340,N_18686,N_18589);
or U19341 (N_19341,N_18956,N_18986);
and U19342 (N_19342,N_18836,N_18844);
nor U19343 (N_19343,N_18713,N_18728);
and U19344 (N_19344,N_18734,N_18960);
or U19345 (N_19345,N_18547,N_18626);
nor U19346 (N_19346,N_18680,N_18669);
and U19347 (N_19347,N_18581,N_18662);
and U19348 (N_19348,N_18717,N_18743);
and U19349 (N_19349,N_18597,N_18909);
xnor U19350 (N_19350,N_18617,N_18934);
or U19351 (N_19351,N_18565,N_18824);
nor U19352 (N_19352,N_18509,N_18525);
and U19353 (N_19353,N_18583,N_18886);
nand U19354 (N_19354,N_18768,N_18539);
xor U19355 (N_19355,N_18952,N_18942);
or U19356 (N_19356,N_18986,N_18607);
nand U19357 (N_19357,N_18992,N_18941);
xnor U19358 (N_19358,N_18940,N_18845);
xor U19359 (N_19359,N_18746,N_18892);
nor U19360 (N_19360,N_18849,N_18550);
nand U19361 (N_19361,N_18848,N_18885);
nand U19362 (N_19362,N_18661,N_18942);
nand U19363 (N_19363,N_18587,N_18879);
xor U19364 (N_19364,N_18622,N_18543);
or U19365 (N_19365,N_18891,N_18907);
nor U19366 (N_19366,N_18835,N_18942);
xor U19367 (N_19367,N_18926,N_18712);
or U19368 (N_19368,N_18710,N_18587);
or U19369 (N_19369,N_18667,N_18900);
nand U19370 (N_19370,N_18865,N_18629);
or U19371 (N_19371,N_18667,N_18963);
xor U19372 (N_19372,N_18562,N_18812);
nor U19373 (N_19373,N_18863,N_18823);
or U19374 (N_19374,N_18516,N_18877);
nor U19375 (N_19375,N_18556,N_18608);
xnor U19376 (N_19376,N_18954,N_18525);
nor U19377 (N_19377,N_18987,N_18858);
and U19378 (N_19378,N_18599,N_18852);
nand U19379 (N_19379,N_18729,N_18551);
xnor U19380 (N_19380,N_18578,N_18598);
xor U19381 (N_19381,N_18949,N_18973);
nand U19382 (N_19382,N_18639,N_18521);
or U19383 (N_19383,N_18526,N_18766);
and U19384 (N_19384,N_18747,N_18843);
and U19385 (N_19385,N_18880,N_18679);
and U19386 (N_19386,N_18787,N_18953);
xnor U19387 (N_19387,N_18860,N_18645);
xor U19388 (N_19388,N_18832,N_18884);
or U19389 (N_19389,N_18665,N_18761);
or U19390 (N_19390,N_18873,N_18767);
nor U19391 (N_19391,N_18959,N_18900);
or U19392 (N_19392,N_18994,N_18839);
or U19393 (N_19393,N_18805,N_18758);
and U19394 (N_19394,N_18599,N_18877);
xor U19395 (N_19395,N_18776,N_18739);
or U19396 (N_19396,N_18512,N_18892);
and U19397 (N_19397,N_18639,N_18713);
and U19398 (N_19398,N_18764,N_18731);
and U19399 (N_19399,N_18685,N_18799);
nor U19400 (N_19400,N_18584,N_18556);
nand U19401 (N_19401,N_18631,N_18541);
or U19402 (N_19402,N_18914,N_18885);
xnor U19403 (N_19403,N_18544,N_18849);
and U19404 (N_19404,N_18781,N_18596);
and U19405 (N_19405,N_18867,N_18759);
nand U19406 (N_19406,N_18524,N_18705);
nand U19407 (N_19407,N_18573,N_18908);
and U19408 (N_19408,N_18697,N_18733);
or U19409 (N_19409,N_18926,N_18627);
or U19410 (N_19410,N_18952,N_18737);
xor U19411 (N_19411,N_18850,N_18626);
nand U19412 (N_19412,N_18832,N_18777);
nor U19413 (N_19413,N_18896,N_18876);
and U19414 (N_19414,N_18811,N_18870);
or U19415 (N_19415,N_18782,N_18623);
nand U19416 (N_19416,N_18767,N_18811);
xnor U19417 (N_19417,N_18813,N_18554);
or U19418 (N_19418,N_18929,N_18864);
nand U19419 (N_19419,N_18746,N_18602);
and U19420 (N_19420,N_18842,N_18740);
or U19421 (N_19421,N_18574,N_18572);
nor U19422 (N_19422,N_18691,N_18912);
and U19423 (N_19423,N_18946,N_18997);
nand U19424 (N_19424,N_18759,N_18725);
nand U19425 (N_19425,N_18842,N_18560);
and U19426 (N_19426,N_18698,N_18988);
or U19427 (N_19427,N_18927,N_18899);
nor U19428 (N_19428,N_18909,N_18754);
or U19429 (N_19429,N_18901,N_18770);
nand U19430 (N_19430,N_18780,N_18795);
or U19431 (N_19431,N_18886,N_18877);
nor U19432 (N_19432,N_18670,N_18877);
nor U19433 (N_19433,N_18552,N_18875);
nand U19434 (N_19434,N_18806,N_18913);
nor U19435 (N_19435,N_18759,N_18655);
xnor U19436 (N_19436,N_18513,N_18671);
nor U19437 (N_19437,N_18964,N_18803);
or U19438 (N_19438,N_18979,N_18601);
nand U19439 (N_19439,N_18701,N_18994);
or U19440 (N_19440,N_18722,N_18941);
or U19441 (N_19441,N_18792,N_18813);
or U19442 (N_19442,N_18902,N_18816);
xor U19443 (N_19443,N_18648,N_18657);
or U19444 (N_19444,N_18700,N_18893);
nand U19445 (N_19445,N_18653,N_18615);
xnor U19446 (N_19446,N_18547,N_18735);
nor U19447 (N_19447,N_18962,N_18814);
nand U19448 (N_19448,N_18658,N_18717);
or U19449 (N_19449,N_18747,N_18983);
and U19450 (N_19450,N_18510,N_18835);
nor U19451 (N_19451,N_18983,N_18806);
or U19452 (N_19452,N_18607,N_18914);
nand U19453 (N_19453,N_18730,N_18507);
and U19454 (N_19454,N_18829,N_18750);
xnor U19455 (N_19455,N_18863,N_18924);
xnor U19456 (N_19456,N_18506,N_18557);
nand U19457 (N_19457,N_18899,N_18723);
nand U19458 (N_19458,N_18700,N_18776);
or U19459 (N_19459,N_18711,N_18956);
and U19460 (N_19460,N_18732,N_18790);
and U19461 (N_19461,N_18937,N_18705);
nor U19462 (N_19462,N_18628,N_18939);
nor U19463 (N_19463,N_18898,N_18581);
or U19464 (N_19464,N_18886,N_18526);
xnor U19465 (N_19465,N_18686,N_18841);
and U19466 (N_19466,N_18663,N_18788);
and U19467 (N_19467,N_18562,N_18944);
xnor U19468 (N_19468,N_18840,N_18924);
or U19469 (N_19469,N_18537,N_18708);
and U19470 (N_19470,N_18680,N_18784);
and U19471 (N_19471,N_18533,N_18778);
and U19472 (N_19472,N_18734,N_18916);
nand U19473 (N_19473,N_18511,N_18940);
and U19474 (N_19474,N_18977,N_18702);
or U19475 (N_19475,N_18533,N_18813);
nor U19476 (N_19476,N_18684,N_18799);
or U19477 (N_19477,N_18650,N_18787);
or U19478 (N_19478,N_18687,N_18980);
nor U19479 (N_19479,N_18670,N_18964);
or U19480 (N_19480,N_18901,N_18571);
or U19481 (N_19481,N_18572,N_18796);
nand U19482 (N_19482,N_18764,N_18902);
or U19483 (N_19483,N_18616,N_18742);
nand U19484 (N_19484,N_18912,N_18758);
xnor U19485 (N_19485,N_18580,N_18549);
nor U19486 (N_19486,N_18624,N_18557);
xnor U19487 (N_19487,N_18769,N_18738);
and U19488 (N_19488,N_18841,N_18679);
xnor U19489 (N_19489,N_18610,N_18789);
and U19490 (N_19490,N_18795,N_18813);
nor U19491 (N_19491,N_18648,N_18720);
nand U19492 (N_19492,N_18744,N_18787);
or U19493 (N_19493,N_18868,N_18620);
xor U19494 (N_19494,N_18883,N_18637);
and U19495 (N_19495,N_18661,N_18785);
nand U19496 (N_19496,N_18846,N_18532);
xor U19497 (N_19497,N_18902,N_18945);
nand U19498 (N_19498,N_18631,N_18529);
and U19499 (N_19499,N_18919,N_18693);
xnor U19500 (N_19500,N_19054,N_19281);
nand U19501 (N_19501,N_19062,N_19142);
nand U19502 (N_19502,N_19388,N_19446);
nor U19503 (N_19503,N_19223,N_19111);
nor U19504 (N_19504,N_19473,N_19452);
nand U19505 (N_19505,N_19072,N_19418);
nand U19506 (N_19506,N_19409,N_19063);
nand U19507 (N_19507,N_19386,N_19244);
nor U19508 (N_19508,N_19147,N_19265);
or U19509 (N_19509,N_19382,N_19058);
xor U19510 (N_19510,N_19442,N_19331);
xor U19511 (N_19511,N_19474,N_19314);
and U19512 (N_19512,N_19343,N_19148);
nor U19513 (N_19513,N_19172,N_19396);
xor U19514 (N_19514,N_19346,N_19470);
or U19515 (N_19515,N_19425,N_19469);
and U19516 (N_19516,N_19431,N_19341);
nand U19517 (N_19517,N_19157,N_19415);
and U19518 (N_19518,N_19158,N_19435);
and U19519 (N_19519,N_19352,N_19486);
or U19520 (N_19520,N_19332,N_19195);
and U19521 (N_19521,N_19347,N_19086);
nand U19522 (N_19522,N_19159,N_19309);
xor U19523 (N_19523,N_19115,N_19497);
xnor U19524 (N_19524,N_19356,N_19334);
nor U19525 (N_19525,N_19216,N_19394);
xor U19526 (N_19526,N_19238,N_19459);
and U19527 (N_19527,N_19079,N_19137);
xor U19528 (N_19528,N_19291,N_19248);
xor U19529 (N_19529,N_19263,N_19283);
nand U19530 (N_19530,N_19108,N_19024);
nand U19531 (N_19531,N_19190,N_19253);
xor U19532 (N_19532,N_19096,N_19162);
nand U19533 (N_19533,N_19071,N_19034);
nand U19534 (N_19534,N_19488,N_19041);
and U19535 (N_19535,N_19095,N_19479);
nor U19536 (N_19536,N_19363,N_19462);
and U19537 (N_19537,N_19203,N_19304);
xor U19538 (N_19538,N_19427,N_19299);
nor U19539 (N_19539,N_19392,N_19270);
xnor U19540 (N_19540,N_19303,N_19466);
nor U19541 (N_19541,N_19116,N_19053);
xnor U19542 (N_19542,N_19428,N_19027);
nor U19543 (N_19543,N_19235,N_19323);
and U19544 (N_19544,N_19328,N_19298);
xor U19545 (N_19545,N_19353,N_19191);
xnor U19546 (N_19546,N_19450,N_19165);
nand U19547 (N_19547,N_19198,N_19308);
xor U19548 (N_19548,N_19066,N_19060);
and U19549 (N_19549,N_19440,N_19239);
nand U19550 (N_19550,N_19374,N_19245);
or U19551 (N_19551,N_19210,N_19133);
xor U19552 (N_19552,N_19493,N_19068);
nand U19553 (N_19553,N_19187,N_19141);
xor U19554 (N_19554,N_19109,N_19406);
xnor U19555 (N_19555,N_19230,N_19075);
and U19556 (N_19556,N_19483,N_19098);
nand U19557 (N_19557,N_19206,N_19188);
nand U19558 (N_19558,N_19391,N_19246);
nand U19559 (N_19559,N_19177,N_19232);
and U19560 (N_19560,N_19321,N_19498);
nor U19561 (N_19561,N_19224,N_19448);
and U19562 (N_19562,N_19390,N_19010);
or U19563 (N_19563,N_19173,N_19164);
or U19564 (N_19564,N_19377,N_19082);
and U19565 (N_19565,N_19128,N_19181);
nand U19566 (N_19566,N_19324,N_19194);
nand U19567 (N_19567,N_19043,N_19376);
or U19568 (N_19568,N_19375,N_19453);
nand U19569 (N_19569,N_19430,N_19080);
or U19570 (N_19570,N_19261,N_19478);
and U19571 (N_19571,N_19397,N_19026);
nor U19572 (N_19572,N_19022,N_19379);
xor U19573 (N_19573,N_19495,N_19124);
or U19574 (N_19574,N_19273,N_19135);
and U19575 (N_19575,N_19077,N_19000);
nor U19576 (N_19576,N_19204,N_19278);
nand U19577 (N_19577,N_19121,N_19342);
nor U19578 (N_19578,N_19107,N_19170);
xor U19579 (N_19579,N_19357,N_19254);
and U19580 (N_19580,N_19084,N_19345);
or U19581 (N_19581,N_19127,N_19130);
and U19582 (N_19582,N_19477,N_19014);
and U19583 (N_19583,N_19404,N_19085);
xor U19584 (N_19584,N_19426,N_19290);
nor U19585 (N_19585,N_19344,N_19046);
nor U19586 (N_19586,N_19259,N_19174);
xor U19587 (N_19587,N_19134,N_19018);
nand U19588 (N_19588,N_19280,N_19484);
xor U19589 (N_19589,N_19132,N_19241);
nor U19590 (N_19590,N_19136,N_19306);
and U19591 (N_19591,N_19381,N_19364);
xor U19592 (N_19592,N_19411,N_19403);
xor U19593 (N_19593,N_19153,N_19393);
or U19594 (N_19594,N_19015,N_19312);
xor U19595 (N_19595,N_19358,N_19091);
xnor U19596 (N_19596,N_19202,N_19185);
or U19597 (N_19597,N_19481,N_19025);
or U19598 (N_19598,N_19419,N_19468);
nor U19599 (N_19599,N_19178,N_19400);
nand U19600 (N_19600,N_19326,N_19255);
xor U19601 (N_19601,N_19316,N_19422);
or U19602 (N_19602,N_19208,N_19252);
nor U19603 (N_19603,N_19247,N_19414);
nor U19604 (N_19604,N_19189,N_19256);
nor U19605 (N_19605,N_19274,N_19036);
xor U19606 (N_19606,N_19269,N_19186);
nand U19607 (N_19607,N_19337,N_19047);
nand U19608 (N_19608,N_19350,N_19480);
nor U19609 (N_19609,N_19219,N_19013);
or U19610 (N_19610,N_19131,N_19327);
and U19611 (N_19611,N_19045,N_19033);
or U19612 (N_19612,N_19297,N_19351);
nor U19613 (N_19613,N_19160,N_19197);
or U19614 (N_19614,N_19372,N_19221);
or U19615 (N_19615,N_19104,N_19310);
xor U19616 (N_19616,N_19285,N_19008);
nand U19617 (N_19617,N_19476,N_19007);
nand U19618 (N_19618,N_19020,N_19105);
nor U19619 (N_19619,N_19083,N_19152);
and U19620 (N_19620,N_19482,N_19338);
xnor U19621 (N_19621,N_19052,N_19184);
nand U19622 (N_19622,N_19092,N_19125);
nor U19623 (N_19623,N_19038,N_19284);
nand U19624 (N_19624,N_19268,N_19492);
or U19625 (N_19625,N_19236,N_19264);
nor U19626 (N_19626,N_19183,N_19067);
or U19627 (N_19627,N_19023,N_19362);
and U19628 (N_19628,N_19485,N_19444);
nor U19629 (N_19629,N_19120,N_19271);
xnor U19630 (N_19630,N_19056,N_19163);
xnor U19631 (N_19631,N_19074,N_19401);
or U19632 (N_19632,N_19410,N_19301);
nor U19633 (N_19633,N_19361,N_19367);
nor U19634 (N_19634,N_19103,N_19461);
xor U19635 (N_19635,N_19168,N_19349);
nand U19636 (N_19636,N_19467,N_19017);
or U19637 (N_19637,N_19171,N_19055);
or U19638 (N_19638,N_19156,N_19296);
nand U19639 (N_19639,N_19455,N_19436);
or U19640 (N_19640,N_19383,N_19424);
nand U19641 (N_19641,N_19429,N_19368);
xor U19642 (N_19642,N_19201,N_19472);
and U19643 (N_19643,N_19030,N_19395);
nand U19644 (N_19644,N_19398,N_19293);
and U19645 (N_19645,N_19145,N_19340);
xnor U19646 (N_19646,N_19001,N_19262);
or U19647 (N_19647,N_19294,N_19012);
or U19648 (N_19648,N_19100,N_19218);
nor U19649 (N_19649,N_19009,N_19258);
or U19650 (N_19650,N_19200,N_19069);
or U19651 (N_19651,N_19335,N_19222);
xor U19652 (N_19652,N_19339,N_19405);
xor U19653 (N_19653,N_19319,N_19408);
nand U19654 (N_19654,N_19412,N_19196);
nand U19655 (N_19655,N_19011,N_19438);
or U19656 (N_19656,N_19275,N_19300);
nand U19657 (N_19657,N_19463,N_19114);
nor U19658 (N_19658,N_19214,N_19193);
nor U19659 (N_19659,N_19433,N_19005);
xnor U19660 (N_19660,N_19051,N_19048);
or U19661 (N_19661,N_19276,N_19102);
or U19662 (N_19662,N_19458,N_19078);
nor U19663 (N_19663,N_19279,N_19369);
and U19664 (N_19664,N_19464,N_19322);
nor U19665 (N_19665,N_19305,N_19049);
and U19666 (N_19666,N_19267,N_19035);
nor U19667 (N_19667,N_19019,N_19028);
nand U19668 (N_19668,N_19112,N_19389);
nand U19669 (N_19669,N_19217,N_19138);
nor U19670 (N_19670,N_19061,N_19402);
nor U19671 (N_19671,N_19315,N_19122);
or U19672 (N_19672,N_19064,N_19150);
or U19673 (N_19673,N_19329,N_19059);
xnor U19674 (N_19674,N_19113,N_19228);
xor U19675 (N_19675,N_19155,N_19295);
or U19676 (N_19676,N_19454,N_19151);
nand U19677 (N_19677,N_19289,N_19231);
nor U19678 (N_19678,N_19336,N_19129);
nor U19679 (N_19679,N_19447,N_19387);
nor U19680 (N_19680,N_19226,N_19443);
and U19681 (N_19681,N_19094,N_19118);
and U19682 (N_19682,N_19257,N_19211);
nor U19683 (N_19683,N_19161,N_19292);
nor U19684 (N_19684,N_19209,N_19097);
nor U19685 (N_19685,N_19207,N_19101);
or U19686 (N_19686,N_19050,N_19359);
nand U19687 (N_19687,N_19365,N_19491);
xnor U19688 (N_19688,N_19039,N_19237);
nor U19689 (N_19689,N_19149,N_19076);
or U19690 (N_19690,N_19166,N_19499);
xor U19691 (N_19691,N_19456,N_19154);
nor U19692 (N_19692,N_19234,N_19099);
and U19693 (N_19693,N_19354,N_19313);
xnor U19694 (N_19694,N_19044,N_19260);
nor U19695 (N_19695,N_19250,N_19437);
and U19696 (N_19696,N_19385,N_19169);
xnor U19697 (N_19697,N_19251,N_19006);
and U19698 (N_19698,N_19494,N_19272);
nor U19699 (N_19699,N_19441,N_19370);
and U19700 (N_19700,N_19212,N_19366);
nand U19701 (N_19701,N_19199,N_19355);
xnor U19702 (N_19702,N_19016,N_19266);
xor U19703 (N_19703,N_19021,N_19240);
nand U19704 (N_19704,N_19144,N_19317);
nand U19705 (N_19705,N_19065,N_19325);
or U19706 (N_19706,N_19249,N_19457);
and U19707 (N_19707,N_19090,N_19176);
xnor U19708 (N_19708,N_19282,N_19004);
xnor U19709 (N_19709,N_19003,N_19089);
nor U19710 (N_19710,N_19373,N_19378);
nand U19711 (N_19711,N_19220,N_19073);
xnor U19712 (N_19712,N_19243,N_19432);
nand U19713 (N_19713,N_19348,N_19330);
nor U19714 (N_19714,N_19070,N_19286);
or U19715 (N_19715,N_19421,N_19487);
nand U19716 (N_19716,N_19123,N_19182);
nand U19717 (N_19717,N_19287,N_19119);
nand U19718 (N_19718,N_19140,N_19180);
and U19719 (N_19719,N_19399,N_19233);
nand U19720 (N_19720,N_19380,N_19360);
nand U19721 (N_19721,N_19496,N_19037);
nor U19722 (N_19722,N_19139,N_19179);
xor U19723 (N_19723,N_19445,N_19227);
xor U19724 (N_19724,N_19439,N_19471);
and U19725 (N_19725,N_19192,N_19057);
nor U19726 (N_19726,N_19318,N_19417);
nand U19727 (N_19727,N_19423,N_19081);
nor U19728 (N_19728,N_19146,N_19032);
nand U19729 (N_19729,N_19489,N_19167);
nor U19730 (N_19730,N_19093,N_19320);
nand U19731 (N_19731,N_19213,N_19475);
xor U19732 (N_19732,N_19040,N_19088);
nand U19733 (N_19733,N_19333,N_19384);
nand U19734 (N_19734,N_19302,N_19413);
xor U19735 (N_19735,N_19215,N_19002);
nor U19736 (N_19736,N_19407,N_19110);
and U19737 (N_19737,N_19288,N_19242);
xnor U19738 (N_19738,N_19225,N_19205);
nor U19739 (N_19739,N_19117,N_19106);
nand U19740 (N_19740,N_19175,N_19449);
nand U19741 (N_19741,N_19451,N_19042);
nor U19742 (N_19742,N_19087,N_19434);
nor U19743 (N_19743,N_19416,N_19420);
nor U19744 (N_19744,N_19371,N_19229);
nor U19745 (N_19745,N_19031,N_19307);
nor U19746 (N_19746,N_19277,N_19029);
nand U19747 (N_19747,N_19311,N_19143);
nand U19748 (N_19748,N_19490,N_19465);
or U19749 (N_19749,N_19460,N_19126);
nand U19750 (N_19750,N_19172,N_19145);
or U19751 (N_19751,N_19103,N_19011);
and U19752 (N_19752,N_19305,N_19082);
and U19753 (N_19753,N_19421,N_19001);
nand U19754 (N_19754,N_19413,N_19179);
and U19755 (N_19755,N_19454,N_19319);
xor U19756 (N_19756,N_19188,N_19149);
or U19757 (N_19757,N_19488,N_19315);
nor U19758 (N_19758,N_19457,N_19013);
or U19759 (N_19759,N_19343,N_19284);
nor U19760 (N_19760,N_19157,N_19083);
nor U19761 (N_19761,N_19052,N_19163);
xnor U19762 (N_19762,N_19349,N_19029);
nor U19763 (N_19763,N_19015,N_19327);
nor U19764 (N_19764,N_19182,N_19142);
nor U19765 (N_19765,N_19315,N_19485);
and U19766 (N_19766,N_19021,N_19494);
nor U19767 (N_19767,N_19046,N_19298);
or U19768 (N_19768,N_19103,N_19230);
and U19769 (N_19769,N_19337,N_19286);
nand U19770 (N_19770,N_19307,N_19080);
or U19771 (N_19771,N_19416,N_19498);
nand U19772 (N_19772,N_19311,N_19052);
nor U19773 (N_19773,N_19087,N_19321);
or U19774 (N_19774,N_19158,N_19305);
xor U19775 (N_19775,N_19305,N_19072);
xor U19776 (N_19776,N_19323,N_19177);
and U19777 (N_19777,N_19038,N_19106);
or U19778 (N_19778,N_19419,N_19277);
and U19779 (N_19779,N_19322,N_19415);
and U19780 (N_19780,N_19064,N_19398);
nand U19781 (N_19781,N_19284,N_19370);
nand U19782 (N_19782,N_19217,N_19013);
nor U19783 (N_19783,N_19046,N_19285);
nor U19784 (N_19784,N_19284,N_19378);
nand U19785 (N_19785,N_19018,N_19237);
nor U19786 (N_19786,N_19154,N_19336);
nor U19787 (N_19787,N_19066,N_19127);
and U19788 (N_19788,N_19436,N_19217);
nand U19789 (N_19789,N_19162,N_19395);
or U19790 (N_19790,N_19231,N_19359);
and U19791 (N_19791,N_19427,N_19320);
nand U19792 (N_19792,N_19008,N_19142);
or U19793 (N_19793,N_19488,N_19042);
or U19794 (N_19794,N_19407,N_19469);
nand U19795 (N_19795,N_19170,N_19287);
xnor U19796 (N_19796,N_19284,N_19099);
xor U19797 (N_19797,N_19100,N_19490);
nor U19798 (N_19798,N_19077,N_19468);
nor U19799 (N_19799,N_19273,N_19008);
xnor U19800 (N_19800,N_19009,N_19120);
and U19801 (N_19801,N_19471,N_19493);
xnor U19802 (N_19802,N_19456,N_19359);
and U19803 (N_19803,N_19151,N_19270);
and U19804 (N_19804,N_19241,N_19365);
nor U19805 (N_19805,N_19213,N_19369);
nor U19806 (N_19806,N_19250,N_19228);
nand U19807 (N_19807,N_19336,N_19237);
nor U19808 (N_19808,N_19138,N_19442);
nor U19809 (N_19809,N_19220,N_19391);
nor U19810 (N_19810,N_19214,N_19026);
nor U19811 (N_19811,N_19115,N_19264);
and U19812 (N_19812,N_19244,N_19085);
nor U19813 (N_19813,N_19072,N_19106);
xnor U19814 (N_19814,N_19303,N_19170);
or U19815 (N_19815,N_19471,N_19291);
nor U19816 (N_19816,N_19024,N_19303);
and U19817 (N_19817,N_19470,N_19182);
nor U19818 (N_19818,N_19214,N_19204);
and U19819 (N_19819,N_19252,N_19480);
xor U19820 (N_19820,N_19017,N_19171);
xor U19821 (N_19821,N_19025,N_19057);
xor U19822 (N_19822,N_19135,N_19390);
xor U19823 (N_19823,N_19102,N_19459);
nor U19824 (N_19824,N_19047,N_19473);
or U19825 (N_19825,N_19061,N_19050);
or U19826 (N_19826,N_19219,N_19229);
nor U19827 (N_19827,N_19101,N_19088);
xor U19828 (N_19828,N_19035,N_19469);
nor U19829 (N_19829,N_19307,N_19238);
or U19830 (N_19830,N_19352,N_19068);
or U19831 (N_19831,N_19300,N_19129);
and U19832 (N_19832,N_19372,N_19062);
and U19833 (N_19833,N_19076,N_19402);
or U19834 (N_19834,N_19008,N_19478);
or U19835 (N_19835,N_19063,N_19387);
and U19836 (N_19836,N_19395,N_19449);
nor U19837 (N_19837,N_19332,N_19049);
nor U19838 (N_19838,N_19474,N_19014);
or U19839 (N_19839,N_19286,N_19291);
and U19840 (N_19840,N_19050,N_19328);
and U19841 (N_19841,N_19220,N_19237);
and U19842 (N_19842,N_19225,N_19385);
or U19843 (N_19843,N_19443,N_19126);
or U19844 (N_19844,N_19051,N_19296);
nand U19845 (N_19845,N_19333,N_19406);
nor U19846 (N_19846,N_19361,N_19276);
or U19847 (N_19847,N_19006,N_19094);
nand U19848 (N_19848,N_19342,N_19048);
nor U19849 (N_19849,N_19461,N_19173);
nand U19850 (N_19850,N_19133,N_19156);
nor U19851 (N_19851,N_19023,N_19430);
or U19852 (N_19852,N_19176,N_19453);
and U19853 (N_19853,N_19216,N_19007);
nand U19854 (N_19854,N_19487,N_19116);
and U19855 (N_19855,N_19354,N_19257);
or U19856 (N_19856,N_19085,N_19126);
nand U19857 (N_19857,N_19422,N_19139);
and U19858 (N_19858,N_19065,N_19237);
nor U19859 (N_19859,N_19123,N_19382);
xor U19860 (N_19860,N_19419,N_19016);
nor U19861 (N_19861,N_19366,N_19237);
and U19862 (N_19862,N_19218,N_19019);
or U19863 (N_19863,N_19351,N_19080);
nand U19864 (N_19864,N_19085,N_19033);
or U19865 (N_19865,N_19282,N_19465);
nor U19866 (N_19866,N_19248,N_19438);
xor U19867 (N_19867,N_19444,N_19354);
and U19868 (N_19868,N_19474,N_19313);
and U19869 (N_19869,N_19217,N_19177);
or U19870 (N_19870,N_19458,N_19358);
nand U19871 (N_19871,N_19348,N_19468);
or U19872 (N_19872,N_19476,N_19411);
xor U19873 (N_19873,N_19344,N_19125);
nor U19874 (N_19874,N_19110,N_19272);
or U19875 (N_19875,N_19342,N_19228);
xor U19876 (N_19876,N_19059,N_19421);
nor U19877 (N_19877,N_19386,N_19054);
nand U19878 (N_19878,N_19144,N_19268);
nand U19879 (N_19879,N_19108,N_19206);
xnor U19880 (N_19880,N_19250,N_19402);
xnor U19881 (N_19881,N_19092,N_19196);
nand U19882 (N_19882,N_19006,N_19096);
nand U19883 (N_19883,N_19149,N_19073);
nand U19884 (N_19884,N_19068,N_19326);
and U19885 (N_19885,N_19008,N_19335);
nor U19886 (N_19886,N_19401,N_19253);
xnor U19887 (N_19887,N_19040,N_19079);
nand U19888 (N_19888,N_19268,N_19401);
nand U19889 (N_19889,N_19091,N_19483);
and U19890 (N_19890,N_19284,N_19418);
xor U19891 (N_19891,N_19210,N_19493);
nor U19892 (N_19892,N_19449,N_19259);
and U19893 (N_19893,N_19132,N_19428);
or U19894 (N_19894,N_19405,N_19143);
nor U19895 (N_19895,N_19329,N_19052);
xnor U19896 (N_19896,N_19024,N_19411);
or U19897 (N_19897,N_19091,N_19176);
and U19898 (N_19898,N_19451,N_19262);
or U19899 (N_19899,N_19426,N_19464);
nor U19900 (N_19900,N_19171,N_19219);
nand U19901 (N_19901,N_19012,N_19482);
and U19902 (N_19902,N_19493,N_19422);
or U19903 (N_19903,N_19234,N_19323);
nor U19904 (N_19904,N_19411,N_19099);
and U19905 (N_19905,N_19285,N_19373);
nor U19906 (N_19906,N_19149,N_19479);
xor U19907 (N_19907,N_19352,N_19450);
or U19908 (N_19908,N_19181,N_19225);
or U19909 (N_19909,N_19074,N_19002);
and U19910 (N_19910,N_19199,N_19063);
or U19911 (N_19911,N_19074,N_19300);
nor U19912 (N_19912,N_19067,N_19350);
or U19913 (N_19913,N_19359,N_19436);
nor U19914 (N_19914,N_19136,N_19464);
xor U19915 (N_19915,N_19343,N_19330);
nor U19916 (N_19916,N_19485,N_19237);
xor U19917 (N_19917,N_19098,N_19203);
nand U19918 (N_19918,N_19083,N_19331);
and U19919 (N_19919,N_19454,N_19448);
xnor U19920 (N_19920,N_19052,N_19300);
nor U19921 (N_19921,N_19036,N_19013);
nor U19922 (N_19922,N_19071,N_19210);
nor U19923 (N_19923,N_19105,N_19352);
nor U19924 (N_19924,N_19019,N_19317);
and U19925 (N_19925,N_19271,N_19269);
and U19926 (N_19926,N_19113,N_19477);
xor U19927 (N_19927,N_19467,N_19057);
nand U19928 (N_19928,N_19297,N_19265);
nor U19929 (N_19929,N_19249,N_19499);
nor U19930 (N_19930,N_19050,N_19357);
or U19931 (N_19931,N_19380,N_19453);
xnor U19932 (N_19932,N_19037,N_19208);
or U19933 (N_19933,N_19022,N_19417);
xor U19934 (N_19934,N_19315,N_19083);
or U19935 (N_19935,N_19313,N_19067);
nand U19936 (N_19936,N_19468,N_19190);
or U19937 (N_19937,N_19391,N_19372);
and U19938 (N_19938,N_19461,N_19140);
and U19939 (N_19939,N_19474,N_19232);
nand U19940 (N_19940,N_19428,N_19449);
nand U19941 (N_19941,N_19118,N_19002);
xor U19942 (N_19942,N_19190,N_19221);
or U19943 (N_19943,N_19350,N_19472);
nand U19944 (N_19944,N_19005,N_19095);
nor U19945 (N_19945,N_19287,N_19250);
or U19946 (N_19946,N_19374,N_19066);
and U19947 (N_19947,N_19022,N_19215);
xor U19948 (N_19948,N_19281,N_19383);
nand U19949 (N_19949,N_19057,N_19062);
and U19950 (N_19950,N_19348,N_19398);
and U19951 (N_19951,N_19428,N_19137);
nand U19952 (N_19952,N_19454,N_19150);
and U19953 (N_19953,N_19296,N_19275);
nor U19954 (N_19954,N_19224,N_19368);
or U19955 (N_19955,N_19406,N_19046);
nor U19956 (N_19956,N_19026,N_19470);
nand U19957 (N_19957,N_19050,N_19000);
and U19958 (N_19958,N_19082,N_19448);
nor U19959 (N_19959,N_19403,N_19355);
nor U19960 (N_19960,N_19103,N_19343);
and U19961 (N_19961,N_19381,N_19397);
or U19962 (N_19962,N_19298,N_19087);
or U19963 (N_19963,N_19299,N_19459);
nand U19964 (N_19964,N_19314,N_19010);
and U19965 (N_19965,N_19182,N_19255);
nand U19966 (N_19966,N_19139,N_19255);
nor U19967 (N_19967,N_19355,N_19446);
nor U19968 (N_19968,N_19046,N_19401);
and U19969 (N_19969,N_19023,N_19304);
nand U19970 (N_19970,N_19415,N_19087);
nor U19971 (N_19971,N_19364,N_19229);
nand U19972 (N_19972,N_19493,N_19201);
nor U19973 (N_19973,N_19468,N_19016);
nand U19974 (N_19974,N_19257,N_19075);
or U19975 (N_19975,N_19380,N_19226);
nor U19976 (N_19976,N_19465,N_19201);
nor U19977 (N_19977,N_19104,N_19385);
xor U19978 (N_19978,N_19359,N_19089);
xnor U19979 (N_19979,N_19499,N_19182);
xor U19980 (N_19980,N_19280,N_19313);
xor U19981 (N_19981,N_19219,N_19446);
xnor U19982 (N_19982,N_19284,N_19265);
or U19983 (N_19983,N_19098,N_19324);
nor U19984 (N_19984,N_19289,N_19428);
nor U19985 (N_19985,N_19459,N_19070);
xnor U19986 (N_19986,N_19113,N_19339);
and U19987 (N_19987,N_19325,N_19404);
nor U19988 (N_19988,N_19359,N_19461);
and U19989 (N_19989,N_19061,N_19493);
nand U19990 (N_19990,N_19055,N_19321);
nand U19991 (N_19991,N_19042,N_19208);
or U19992 (N_19992,N_19196,N_19044);
xnor U19993 (N_19993,N_19237,N_19474);
and U19994 (N_19994,N_19074,N_19116);
xor U19995 (N_19995,N_19059,N_19000);
xnor U19996 (N_19996,N_19338,N_19419);
nor U19997 (N_19997,N_19494,N_19364);
and U19998 (N_19998,N_19482,N_19249);
and U19999 (N_19999,N_19138,N_19159);
or U20000 (N_20000,N_19516,N_19761);
nand U20001 (N_20001,N_19510,N_19779);
or U20002 (N_20002,N_19864,N_19949);
or U20003 (N_20003,N_19693,N_19591);
and U20004 (N_20004,N_19702,N_19902);
and U20005 (N_20005,N_19858,N_19912);
or U20006 (N_20006,N_19571,N_19915);
or U20007 (N_20007,N_19964,N_19894);
nor U20008 (N_20008,N_19877,N_19951);
nor U20009 (N_20009,N_19579,N_19670);
and U20010 (N_20010,N_19808,N_19852);
nor U20011 (N_20011,N_19961,N_19703);
nor U20012 (N_20012,N_19757,N_19501);
and U20013 (N_20013,N_19946,N_19514);
or U20014 (N_20014,N_19942,N_19764);
or U20015 (N_20015,N_19650,N_19513);
nand U20016 (N_20016,N_19874,N_19537);
and U20017 (N_20017,N_19704,N_19809);
xor U20018 (N_20018,N_19847,N_19802);
or U20019 (N_20019,N_19661,N_19713);
nor U20020 (N_20020,N_19633,N_19724);
or U20021 (N_20021,N_19508,N_19963);
nand U20022 (N_20022,N_19672,N_19971);
nand U20023 (N_20023,N_19876,N_19934);
and U20024 (N_20024,N_19935,N_19891);
xor U20025 (N_20025,N_19739,N_19583);
xnor U20026 (N_20026,N_19622,N_19683);
nand U20027 (N_20027,N_19899,N_19829);
and U20028 (N_20028,N_19780,N_19958);
or U20029 (N_20029,N_19924,N_19986);
xor U20030 (N_20030,N_19792,N_19542);
or U20031 (N_20031,N_19828,N_19791);
and U20032 (N_20032,N_19860,N_19502);
xor U20033 (N_20033,N_19675,N_19766);
xor U20034 (N_20034,N_19612,N_19561);
and U20035 (N_20035,N_19782,N_19937);
nor U20036 (N_20036,N_19669,N_19699);
xnor U20037 (N_20037,N_19646,N_19656);
nor U20038 (N_20038,N_19707,N_19639);
and U20039 (N_20039,N_19846,N_19574);
and U20040 (N_20040,N_19658,N_19567);
and U20041 (N_20041,N_19705,N_19851);
nand U20042 (N_20042,N_19726,N_19817);
or U20043 (N_20043,N_19805,N_19523);
or U20044 (N_20044,N_19565,N_19831);
or U20045 (N_20045,N_19970,N_19833);
or U20046 (N_20046,N_19668,N_19957);
nand U20047 (N_20047,N_19888,N_19590);
xor U20048 (N_20048,N_19746,N_19740);
and U20049 (N_20049,N_19834,N_19840);
and U20050 (N_20050,N_19914,N_19556);
nand U20051 (N_20051,N_19988,N_19641);
nand U20052 (N_20052,N_19992,N_19652);
or U20053 (N_20053,N_19917,N_19967);
or U20054 (N_20054,N_19528,N_19532);
nand U20055 (N_20055,N_19547,N_19798);
nand U20056 (N_20056,N_19816,N_19619);
or U20057 (N_20057,N_19947,N_19944);
or U20058 (N_20058,N_19870,N_19637);
xnor U20059 (N_20059,N_19889,N_19842);
xor U20060 (N_20060,N_19687,N_19714);
nand U20061 (N_20061,N_19885,N_19535);
nand U20062 (N_20062,N_19898,N_19807);
and U20063 (N_20063,N_19578,N_19850);
xor U20064 (N_20064,N_19555,N_19674);
or U20065 (N_20065,N_19625,N_19742);
xnor U20066 (N_20066,N_19526,N_19938);
xor U20067 (N_20067,N_19901,N_19673);
nor U20068 (N_20068,N_19697,N_19984);
nor U20069 (N_20069,N_19760,N_19500);
xor U20070 (N_20070,N_19908,N_19995);
and U20071 (N_20071,N_19589,N_19618);
and U20072 (N_20072,N_19727,N_19977);
nor U20073 (N_20073,N_19839,N_19982);
and U20074 (N_20074,N_19796,N_19954);
and U20075 (N_20075,N_19651,N_19887);
and U20076 (N_20076,N_19654,N_19920);
nor U20077 (N_20077,N_19631,N_19715);
nor U20078 (N_20078,N_19932,N_19595);
or U20079 (N_20079,N_19962,N_19538);
xnor U20080 (N_20080,N_19710,N_19677);
and U20081 (N_20081,N_19621,N_19793);
xor U20082 (N_20082,N_19611,N_19666);
nand U20083 (N_20083,N_19781,N_19557);
xnor U20084 (N_20084,N_19733,N_19925);
and U20085 (N_20085,N_19506,N_19563);
xnor U20086 (N_20086,N_19832,N_19552);
nor U20087 (N_20087,N_19533,N_19968);
xnor U20088 (N_20088,N_19709,N_19730);
xor U20089 (N_20089,N_19620,N_19728);
or U20090 (N_20090,N_19572,N_19911);
and U20091 (N_20091,N_19985,N_19734);
xor U20092 (N_20092,N_19863,N_19799);
nor U20093 (N_20093,N_19873,N_19721);
nor U20094 (N_20094,N_19955,N_19684);
nor U20095 (N_20095,N_19856,N_19754);
and U20096 (N_20096,N_19784,N_19830);
nand U20097 (N_20097,N_19504,N_19753);
or U20098 (N_20098,N_19745,N_19723);
xnor U20099 (N_20099,N_19685,N_19866);
nor U20100 (N_20100,N_19940,N_19653);
nand U20101 (N_20101,N_19550,N_19539);
or U20102 (N_20102,N_19731,N_19806);
or U20103 (N_20103,N_19789,N_19628);
or U20104 (N_20104,N_19606,N_19797);
nand U20105 (N_20105,N_19872,N_19862);
or U20106 (N_20106,N_19783,N_19900);
xor U20107 (N_20107,N_19662,N_19857);
and U20108 (N_20108,N_19698,N_19773);
xor U20109 (N_20109,N_19608,N_19998);
and U20110 (N_20110,N_19975,N_19741);
nand U20111 (N_20111,N_19577,N_19680);
nor U20112 (N_20112,N_19979,N_19544);
or U20113 (N_20113,N_19960,N_19747);
nor U20114 (N_20114,N_19815,N_19930);
or U20115 (N_20115,N_19649,N_19838);
xnor U20116 (N_20116,N_19616,N_19729);
or U20117 (N_20117,N_19913,N_19923);
xor U20118 (N_20118,N_19562,N_19800);
xor U20119 (N_20119,N_19517,N_19593);
or U20120 (N_20120,N_19823,N_19795);
and U20121 (N_20121,N_19640,N_19818);
nor U20122 (N_20122,N_19682,N_19529);
nor U20123 (N_20123,N_19569,N_19647);
nor U20124 (N_20124,N_19859,N_19629);
xnor U20125 (N_20125,N_19893,N_19660);
xnor U20126 (N_20126,N_19849,N_19814);
or U20127 (N_20127,N_19587,N_19719);
or U20128 (N_20128,N_19566,N_19627);
and U20129 (N_20129,N_19610,N_19844);
xnor U20130 (N_20130,N_19762,N_19676);
xor U20131 (N_20131,N_19599,N_19999);
or U20132 (N_20132,N_19597,N_19879);
nand U20133 (N_20133,N_19884,N_19548);
and U20134 (N_20134,N_19813,N_19867);
xnor U20135 (N_20135,N_19663,N_19965);
xor U20136 (N_20136,N_19630,N_19522);
nand U20137 (N_20137,N_19880,N_19895);
nand U20138 (N_20138,N_19643,N_19575);
xor U20139 (N_20139,N_19671,N_19748);
or U20140 (N_20140,N_19777,N_19755);
or U20141 (N_20141,N_19507,N_19648);
and U20142 (N_20142,N_19695,N_19580);
nand U20143 (N_20143,N_19617,N_19804);
nand U20144 (N_20144,N_19765,N_19665);
and U20145 (N_20145,N_19869,N_19758);
nand U20146 (N_20146,N_19751,N_19546);
nor U20147 (N_20147,N_19551,N_19716);
or U20148 (N_20148,N_19701,N_19657);
nor U20149 (N_20149,N_19875,N_19512);
nor U20150 (N_20150,N_19598,N_19503);
and U20151 (N_20151,N_19564,N_19768);
xnor U20152 (N_20152,N_19763,N_19978);
or U20153 (N_20153,N_19868,N_19545);
nor U20154 (N_20154,N_19664,N_19624);
nand U20155 (N_20155,N_19638,N_19910);
nand U20156 (N_20156,N_19694,N_19626);
nor U20157 (N_20157,N_19634,N_19835);
or U20158 (N_20158,N_19774,N_19511);
and U20159 (N_20159,N_19553,N_19738);
nand U20160 (N_20160,N_19520,N_19576);
or U20161 (N_20161,N_19827,N_19836);
nor U20162 (N_20162,N_19882,N_19689);
and U20163 (N_20163,N_19903,N_19854);
and U20164 (N_20164,N_19688,N_19994);
or U20165 (N_20165,N_19604,N_19991);
xor U20166 (N_20166,N_19615,N_19600);
or U20167 (N_20167,N_19794,N_19905);
or U20168 (N_20168,N_19776,N_19655);
and U20169 (N_20169,N_19558,N_19744);
nand U20170 (N_20170,N_19559,N_19959);
nor U20171 (N_20171,N_19700,N_19973);
xnor U20172 (N_20172,N_19525,N_19554);
xnor U20173 (N_20173,N_19890,N_19841);
and U20174 (N_20174,N_19936,N_19881);
nand U20175 (N_20175,N_19770,N_19976);
nand U20176 (N_20176,N_19993,N_19931);
and U20177 (N_20177,N_19956,N_19843);
and U20178 (N_20178,N_19752,N_19560);
nor U20179 (N_20179,N_19926,N_19603);
xnor U20180 (N_20180,N_19922,N_19886);
or U20181 (N_20181,N_19540,N_19586);
nor U20182 (N_20182,N_19582,N_19918);
nand U20183 (N_20183,N_19594,N_19848);
xnor U20184 (N_20184,N_19896,N_19969);
xor U20185 (N_20185,N_19644,N_19585);
nor U20186 (N_20186,N_19596,N_19790);
or U20187 (N_20187,N_19801,N_19845);
xor U20188 (N_20188,N_19518,N_19711);
nor U20189 (N_20189,N_19588,N_19735);
nand U20190 (N_20190,N_19524,N_19929);
nand U20191 (N_20191,N_19549,N_19614);
xor U20192 (N_20192,N_19855,N_19897);
and U20193 (N_20193,N_19570,N_19659);
or U20194 (N_20194,N_19717,N_19950);
and U20195 (N_20195,N_19605,N_19691);
xnor U20196 (N_20196,N_19636,N_19759);
xor U20197 (N_20197,N_19945,N_19667);
and U20198 (N_20198,N_19632,N_19990);
or U20199 (N_20199,N_19645,N_19778);
nand U20200 (N_20200,N_19941,N_19749);
xnor U20201 (N_20201,N_19916,N_19906);
and U20202 (N_20202,N_19706,N_19812);
and U20203 (N_20203,N_19811,N_19708);
nand U20204 (N_20204,N_19865,N_19718);
nand U20205 (N_20205,N_19581,N_19681);
xor U20206 (N_20206,N_19825,N_19788);
or U20207 (N_20207,N_19786,N_19983);
or U20208 (N_20208,N_19939,N_19821);
nor U20209 (N_20209,N_19953,N_19530);
nand U20210 (N_20210,N_19592,N_19623);
nand U20211 (N_20211,N_19527,N_19536);
and U20212 (N_20212,N_19837,N_19987);
and U20213 (N_20213,N_19927,N_19981);
nor U20214 (N_20214,N_19787,N_19803);
nand U20215 (N_20215,N_19732,N_19519);
nor U20216 (N_20216,N_19521,N_19686);
and U20217 (N_20217,N_19607,N_19505);
nand U20218 (N_20218,N_19743,N_19573);
nand U20219 (N_20219,N_19725,N_19678);
nand U20220 (N_20220,N_19819,N_19609);
nor U20221 (N_20221,N_19853,N_19907);
and U20222 (N_20222,N_19822,N_19642);
xor U20223 (N_20223,N_19692,N_19531);
xor U20224 (N_20224,N_19568,N_19767);
and U20225 (N_20225,N_19712,N_19769);
and U20226 (N_20226,N_19584,N_19772);
or U20227 (N_20227,N_19972,N_19826);
and U20228 (N_20228,N_19824,N_19919);
xnor U20229 (N_20229,N_19974,N_19966);
and U20230 (N_20230,N_19737,N_19720);
and U20231 (N_20231,N_19679,N_19602);
or U20232 (N_20232,N_19980,N_19921);
or U20233 (N_20233,N_19613,N_19750);
nand U20234 (N_20234,N_19785,N_19515);
nand U20235 (N_20235,N_19722,N_19601);
nor U20236 (N_20236,N_19952,N_19928);
xor U20237 (N_20237,N_19820,N_19541);
and U20238 (N_20238,N_19904,N_19534);
or U20239 (N_20239,N_19635,N_19543);
and U20240 (N_20240,N_19861,N_19997);
or U20241 (N_20241,N_19883,N_19933);
nand U20242 (N_20242,N_19871,N_19810);
nor U20243 (N_20243,N_19690,N_19878);
xnor U20244 (N_20244,N_19909,N_19736);
xnor U20245 (N_20245,N_19892,N_19775);
nand U20246 (N_20246,N_19989,N_19771);
and U20247 (N_20247,N_19996,N_19509);
xor U20248 (N_20248,N_19943,N_19696);
nor U20249 (N_20249,N_19756,N_19948);
xnor U20250 (N_20250,N_19913,N_19588);
and U20251 (N_20251,N_19964,N_19880);
or U20252 (N_20252,N_19500,N_19561);
or U20253 (N_20253,N_19642,N_19549);
or U20254 (N_20254,N_19998,N_19816);
or U20255 (N_20255,N_19814,N_19562);
or U20256 (N_20256,N_19827,N_19568);
nand U20257 (N_20257,N_19904,N_19780);
and U20258 (N_20258,N_19623,N_19953);
nor U20259 (N_20259,N_19991,N_19949);
nor U20260 (N_20260,N_19769,N_19839);
xnor U20261 (N_20261,N_19612,N_19554);
nand U20262 (N_20262,N_19778,N_19851);
or U20263 (N_20263,N_19586,N_19545);
nor U20264 (N_20264,N_19551,N_19628);
nor U20265 (N_20265,N_19832,N_19687);
nor U20266 (N_20266,N_19690,N_19640);
or U20267 (N_20267,N_19552,N_19612);
nor U20268 (N_20268,N_19808,N_19732);
and U20269 (N_20269,N_19724,N_19516);
nand U20270 (N_20270,N_19741,N_19953);
or U20271 (N_20271,N_19966,N_19629);
xor U20272 (N_20272,N_19777,N_19876);
nand U20273 (N_20273,N_19821,N_19504);
xor U20274 (N_20274,N_19656,N_19541);
xor U20275 (N_20275,N_19559,N_19951);
nor U20276 (N_20276,N_19993,N_19733);
or U20277 (N_20277,N_19968,N_19540);
or U20278 (N_20278,N_19580,N_19659);
and U20279 (N_20279,N_19557,N_19766);
nand U20280 (N_20280,N_19558,N_19832);
and U20281 (N_20281,N_19616,N_19815);
nor U20282 (N_20282,N_19935,N_19572);
nand U20283 (N_20283,N_19866,N_19628);
and U20284 (N_20284,N_19994,N_19560);
and U20285 (N_20285,N_19513,N_19561);
xnor U20286 (N_20286,N_19631,N_19784);
xnor U20287 (N_20287,N_19686,N_19653);
xnor U20288 (N_20288,N_19542,N_19563);
and U20289 (N_20289,N_19938,N_19943);
or U20290 (N_20290,N_19837,N_19818);
nor U20291 (N_20291,N_19599,N_19571);
xor U20292 (N_20292,N_19907,N_19806);
nor U20293 (N_20293,N_19773,N_19587);
nand U20294 (N_20294,N_19639,N_19531);
or U20295 (N_20295,N_19729,N_19964);
and U20296 (N_20296,N_19941,N_19904);
and U20297 (N_20297,N_19871,N_19812);
nand U20298 (N_20298,N_19899,N_19555);
and U20299 (N_20299,N_19927,N_19588);
nor U20300 (N_20300,N_19955,N_19602);
nor U20301 (N_20301,N_19606,N_19666);
nand U20302 (N_20302,N_19581,N_19570);
nor U20303 (N_20303,N_19570,N_19542);
and U20304 (N_20304,N_19640,N_19856);
or U20305 (N_20305,N_19559,N_19622);
or U20306 (N_20306,N_19875,N_19792);
and U20307 (N_20307,N_19644,N_19676);
and U20308 (N_20308,N_19660,N_19574);
xor U20309 (N_20309,N_19533,N_19796);
nand U20310 (N_20310,N_19511,N_19988);
or U20311 (N_20311,N_19577,N_19853);
or U20312 (N_20312,N_19667,N_19901);
xor U20313 (N_20313,N_19606,N_19680);
and U20314 (N_20314,N_19746,N_19794);
nor U20315 (N_20315,N_19778,N_19681);
or U20316 (N_20316,N_19505,N_19914);
nand U20317 (N_20317,N_19773,N_19764);
xor U20318 (N_20318,N_19619,N_19918);
xnor U20319 (N_20319,N_19763,N_19737);
nor U20320 (N_20320,N_19929,N_19787);
xnor U20321 (N_20321,N_19971,N_19815);
nor U20322 (N_20322,N_19860,N_19723);
nand U20323 (N_20323,N_19772,N_19939);
nand U20324 (N_20324,N_19595,N_19567);
and U20325 (N_20325,N_19834,N_19690);
xnor U20326 (N_20326,N_19652,N_19948);
nand U20327 (N_20327,N_19826,N_19676);
and U20328 (N_20328,N_19847,N_19668);
xor U20329 (N_20329,N_19568,N_19691);
or U20330 (N_20330,N_19875,N_19947);
and U20331 (N_20331,N_19783,N_19778);
or U20332 (N_20332,N_19845,N_19862);
and U20333 (N_20333,N_19631,N_19716);
or U20334 (N_20334,N_19515,N_19772);
nor U20335 (N_20335,N_19527,N_19622);
and U20336 (N_20336,N_19572,N_19791);
nor U20337 (N_20337,N_19953,N_19876);
or U20338 (N_20338,N_19969,N_19900);
nor U20339 (N_20339,N_19962,N_19640);
or U20340 (N_20340,N_19828,N_19549);
xor U20341 (N_20341,N_19547,N_19802);
and U20342 (N_20342,N_19783,N_19524);
nand U20343 (N_20343,N_19918,N_19615);
nand U20344 (N_20344,N_19970,N_19844);
or U20345 (N_20345,N_19706,N_19735);
nor U20346 (N_20346,N_19886,N_19894);
nor U20347 (N_20347,N_19583,N_19824);
or U20348 (N_20348,N_19683,N_19872);
and U20349 (N_20349,N_19628,N_19629);
or U20350 (N_20350,N_19711,N_19664);
or U20351 (N_20351,N_19580,N_19577);
xnor U20352 (N_20352,N_19857,N_19674);
xor U20353 (N_20353,N_19609,N_19758);
xnor U20354 (N_20354,N_19861,N_19871);
and U20355 (N_20355,N_19964,N_19802);
nor U20356 (N_20356,N_19525,N_19678);
xnor U20357 (N_20357,N_19904,N_19751);
xor U20358 (N_20358,N_19652,N_19955);
nand U20359 (N_20359,N_19934,N_19767);
xnor U20360 (N_20360,N_19796,N_19817);
xor U20361 (N_20361,N_19872,N_19911);
or U20362 (N_20362,N_19603,N_19877);
nand U20363 (N_20363,N_19759,N_19703);
xor U20364 (N_20364,N_19886,N_19974);
nor U20365 (N_20365,N_19525,N_19805);
nor U20366 (N_20366,N_19531,N_19693);
xor U20367 (N_20367,N_19824,N_19762);
nand U20368 (N_20368,N_19915,N_19596);
and U20369 (N_20369,N_19997,N_19708);
nand U20370 (N_20370,N_19987,N_19725);
nand U20371 (N_20371,N_19597,N_19926);
xor U20372 (N_20372,N_19524,N_19869);
nor U20373 (N_20373,N_19514,N_19756);
nand U20374 (N_20374,N_19528,N_19973);
xor U20375 (N_20375,N_19868,N_19626);
or U20376 (N_20376,N_19765,N_19934);
nor U20377 (N_20377,N_19668,N_19956);
xnor U20378 (N_20378,N_19904,N_19662);
nand U20379 (N_20379,N_19993,N_19736);
and U20380 (N_20380,N_19961,N_19545);
nor U20381 (N_20381,N_19606,N_19652);
and U20382 (N_20382,N_19877,N_19533);
nand U20383 (N_20383,N_19696,N_19784);
or U20384 (N_20384,N_19832,N_19659);
nand U20385 (N_20385,N_19805,N_19593);
xnor U20386 (N_20386,N_19862,N_19851);
or U20387 (N_20387,N_19560,N_19936);
xor U20388 (N_20388,N_19567,N_19569);
nor U20389 (N_20389,N_19975,N_19811);
and U20390 (N_20390,N_19589,N_19703);
nand U20391 (N_20391,N_19533,N_19805);
xnor U20392 (N_20392,N_19958,N_19586);
or U20393 (N_20393,N_19505,N_19657);
or U20394 (N_20394,N_19504,N_19932);
or U20395 (N_20395,N_19878,N_19703);
xor U20396 (N_20396,N_19550,N_19501);
xor U20397 (N_20397,N_19873,N_19772);
xor U20398 (N_20398,N_19911,N_19737);
or U20399 (N_20399,N_19629,N_19553);
nand U20400 (N_20400,N_19500,N_19787);
xnor U20401 (N_20401,N_19973,N_19588);
nor U20402 (N_20402,N_19592,N_19672);
and U20403 (N_20403,N_19513,N_19783);
nand U20404 (N_20404,N_19979,N_19534);
nand U20405 (N_20405,N_19789,N_19816);
nor U20406 (N_20406,N_19970,N_19874);
xnor U20407 (N_20407,N_19779,N_19537);
xor U20408 (N_20408,N_19534,N_19631);
nor U20409 (N_20409,N_19543,N_19986);
nand U20410 (N_20410,N_19755,N_19740);
xor U20411 (N_20411,N_19727,N_19978);
nand U20412 (N_20412,N_19510,N_19813);
nor U20413 (N_20413,N_19691,N_19833);
nor U20414 (N_20414,N_19996,N_19773);
nor U20415 (N_20415,N_19840,N_19796);
xor U20416 (N_20416,N_19570,N_19671);
or U20417 (N_20417,N_19581,N_19578);
and U20418 (N_20418,N_19533,N_19572);
and U20419 (N_20419,N_19600,N_19701);
and U20420 (N_20420,N_19605,N_19539);
nand U20421 (N_20421,N_19981,N_19546);
and U20422 (N_20422,N_19631,N_19665);
nor U20423 (N_20423,N_19509,N_19936);
or U20424 (N_20424,N_19892,N_19601);
nand U20425 (N_20425,N_19890,N_19886);
xnor U20426 (N_20426,N_19997,N_19782);
nand U20427 (N_20427,N_19781,N_19892);
or U20428 (N_20428,N_19689,N_19886);
nand U20429 (N_20429,N_19710,N_19788);
nor U20430 (N_20430,N_19876,N_19828);
xor U20431 (N_20431,N_19522,N_19603);
nor U20432 (N_20432,N_19749,N_19508);
or U20433 (N_20433,N_19661,N_19571);
nand U20434 (N_20434,N_19952,N_19667);
xor U20435 (N_20435,N_19834,N_19981);
or U20436 (N_20436,N_19986,N_19678);
or U20437 (N_20437,N_19637,N_19779);
nand U20438 (N_20438,N_19575,N_19831);
and U20439 (N_20439,N_19611,N_19890);
nor U20440 (N_20440,N_19644,N_19911);
xnor U20441 (N_20441,N_19666,N_19653);
or U20442 (N_20442,N_19923,N_19549);
nand U20443 (N_20443,N_19558,N_19919);
or U20444 (N_20444,N_19832,N_19819);
nand U20445 (N_20445,N_19946,N_19885);
nor U20446 (N_20446,N_19564,N_19547);
nand U20447 (N_20447,N_19539,N_19597);
xnor U20448 (N_20448,N_19888,N_19773);
xor U20449 (N_20449,N_19645,N_19590);
and U20450 (N_20450,N_19574,N_19860);
or U20451 (N_20451,N_19930,N_19819);
nand U20452 (N_20452,N_19637,N_19621);
xnor U20453 (N_20453,N_19850,N_19786);
nand U20454 (N_20454,N_19597,N_19723);
nand U20455 (N_20455,N_19983,N_19773);
nand U20456 (N_20456,N_19654,N_19800);
and U20457 (N_20457,N_19695,N_19677);
or U20458 (N_20458,N_19575,N_19806);
nand U20459 (N_20459,N_19786,N_19680);
and U20460 (N_20460,N_19973,N_19542);
xnor U20461 (N_20461,N_19622,N_19742);
or U20462 (N_20462,N_19702,N_19510);
or U20463 (N_20463,N_19638,N_19982);
or U20464 (N_20464,N_19949,N_19769);
nor U20465 (N_20465,N_19507,N_19855);
or U20466 (N_20466,N_19948,N_19959);
nand U20467 (N_20467,N_19923,N_19837);
and U20468 (N_20468,N_19561,N_19988);
xnor U20469 (N_20469,N_19787,N_19995);
or U20470 (N_20470,N_19662,N_19716);
xor U20471 (N_20471,N_19728,N_19944);
or U20472 (N_20472,N_19803,N_19778);
xnor U20473 (N_20473,N_19642,N_19969);
nor U20474 (N_20474,N_19675,N_19971);
xnor U20475 (N_20475,N_19569,N_19511);
or U20476 (N_20476,N_19773,N_19627);
or U20477 (N_20477,N_19888,N_19952);
nand U20478 (N_20478,N_19805,N_19730);
and U20479 (N_20479,N_19610,N_19887);
or U20480 (N_20480,N_19866,N_19870);
or U20481 (N_20481,N_19820,N_19793);
nor U20482 (N_20482,N_19752,N_19711);
nor U20483 (N_20483,N_19975,N_19778);
nor U20484 (N_20484,N_19573,N_19640);
nor U20485 (N_20485,N_19904,N_19624);
and U20486 (N_20486,N_19953,N_19561);
nor U20487 (N_20487,N_19940,N_19622);
and U20488 (N_20488,N_19533,N_19782);
or U20489 (N_20489,N_19924,N_19915);
xor U20490 (N_20490,N_19676,N_19884);
and U20491 (N_20491,N_19524,N_19601);
or U20492 (N_20492,N_19779,N_19927);
nor U20493 (N_20493,N_19669,N_19798);
xnor U20494 (N_20494,N_19717,N_19622);
nand U20495 (N_20495,N_19543,N_19533);
nand U20496 (N_20496,N_19647,N_19749);
and U20497 (N_20497,N_19998,N_19682);
nand U20498 (N_20498,N_19700,N_19611);
or U20499 (N_20499,N_19799,N_19540);
xor U20500 (N_20500,N_20429,N_20323);
xnor U20501 (N_20501,N_20225,N_20215);
nor U20502 (N_20502,N_20014,N_20007);
nor U20503 (N_20503,N_20259,N_20171);
nor U20504 (N_20504,N_20421,N_20335);
nor U20505 (N_20505,N_20164,N_20015);
xnor U20506 (N_20506,N_20208,N_20357);
nor U20507 (N_20507,N_20165,N_20248);
nand U20508 (N_20508,N_20040,N_20163);
nor U20509 (N_20509,N_20145,N_20337);
xor U20510 (N_20510,N_20127,N_20422);
and U20511 (N_20511,N_20081,N_20334);
and U20512 (N_20512,N_20201,N_20031);
and U20513 (N_20513,N_20440,N_20012);
nor U20514 (N_20514,N_20463,N_20155);
and U20515 (N_20515,N_20350,N_20411);
nor U20516 (N_20516,N_20394,N_20432);
or U20517 (N_20517,N_20090,N_20453);
xnor U20518 (N_20518,N_20373,N_20021);
xor U20519 (N_20519,N_20181,N_20405);
xor U20520 (N_20520,N_20486,N_20467);
and U20521 (N_20521,N_20317,N_20172);
nand U20522 (N_20522,N_20389,N_20434);
nor U20523 (N_20523,N_20410,N_20112);
or U20524 (N_20524,N_20044,N_20094);
nor U20525 (N_20525,N_20151,N_20079);
or U20526 (N_20526,N_20420,N_20193);
or U20527 (N_20527,N_20371,N_20472);
nand U20528 (N_20528,N_20068,N_20384);
or U20529 (N_20529,N_20365,N_20297);
xor U20530 (N_20530,N_20345,N_20366);
nand U20531 (N_20531,N_20180,N_20426);
xor U20532 (N_20532,N_20053,N_20298);
nand U20533 (N_20533,N_20244,N_20257);
nand U20534 (N_20534,N_20025,N_20439);
or U20535 (N_20535,N_20119,N_20062);
nand U20536 (N_20536,N_20316,N_20454);
nor U20537 (N_20537,N_20184,N_20234);
and U20538 (N_20538,N_20362,N_20498);
and U20539 (N_20539,N_20205,N_20149);
xor U20540 (N_20540,N_20416,N_20437);
xor U20541 (N_20541,N_20199,N_20159);
xor U20542 (N_20542,N_20280,N_20261);
xor U20543 (N_20543,N_20085,N_20256);
xnor U20544 (N_20544,N_20448,N_20377);
nor U20545 (N_20545,N_20153,N_20202);
nand U20546 (N_20546,N_20427,N_20478);
or U20547 (N_20547,N_20188,N_20032);
nand U20548 (N_20548,N_20104,N_20333);
xnor U20549 (N_20549,N_20482,N_20459);
and U20550 (N_20550,N_20003,N_20358);
xor U20551 (N_20551,N_20018,N_20457);
xnor U20552 (N_20552,N_20057,N_20056);
xnor U20553 (N_20553,N_20131,N_20237);
and U20554 (N_20554,N_20026,N_20230);
nand U20555 (N_20555,N_20361,N_20226);
or U20556 (N_20556,N_20247,N_20446);
nand U20557 (N_20557,N_20239,N_20279);
xor U20558 (N_20558,N_20344,N_20236);
nor U20559 (N_20559,N_20400,N_20102);
nor U20560 (N_20560,N_20418,N_20255);
or U20561 (N_20561,N_20229,N_20108);
xnor U20562 (N_20562,N_20238,N_20273);
nand U20563 (N_20563,N_20197,N_20060);
xor U20564 (N_20564,N_20260,N_20277);
xor U20565 (N_20565,N_20047,N_20319);
xor U20566 (N_20566,N_20253,N_20294);
nand U20567 (N_20567,N_20049,N_20072);
nor U20568 (N_20568,N_20243,N_20495);
nand U20569 (N_20569,N_20251,N_20222);
nor U20570 (N_20570,N_20218,N_20302);
xor U20571 (N_20571,N_20262,N_20336);
xnor U20572 (N_20572,N_20070,N_20211);
or U20573 (N_20573,N_20156,N_20084);
and U20574 (N_20574,N_20168,N_20479);
xnor U20575 (N_20575,N_20200,N_20122);
or U20576 (N_20576,N_20158,N_20374);
nor U20577 (N_20577,N_20150,N_20438);
xor U20578 (N_20578,N_20488,N_20010);
or U20579 (N_20579,N_20324,N_20378);
nand U20580 (N_20580,N_20338,N_20162);
nand U20581 (N_20581,N_20073,N_20235);
or U20582 (N_20582,N_20456,N_20497);
or U20583 (N_20583,N_20398,N_20091);
or U20584 (N_20584,N_20332,N_20415);
nor U20585 (N_20585,N_20231,N_20413);
or U20586 (N_20586,N_20223,N_20143);
xor U20587 (N_20587,N_20441,N_20008);
xor U20588 (N_20588,N_20340,N_20460);
or U20589 (N_20589,N_20083,N_20187);
xnor U20590 (N_20590,N_20175,N_20227);
nand U20591 (N_20591,N_20423,N_20349);
nand U20592 (N_20592,N_20354,N_20372);
nor U20593 (N_20593,N_20216,N_20138);
and U20594 (N_20594,N_20481,N_20086);
and U20595 (N_20595,N_20381,N_20061);
or U20596 (N_20596,N_20249,N_20196);
xnor U20597 (N_20597,N_20469,N_20359);
nand U20598 (N_20598,N_20191,N_20036);
nand U20599 (N_20599,N_20137,N_20265);
and U20600 (N_20600,N_20161,N_20152);
or U20601 (N_20601,N_20281,N_20355);
or U20602 (N_20602,N_20451,N_20414);
xnor U20603 (N_20603,N_20470,N_20407);
or U20604 (N_20604,N_20046,N_20055);
nand U20605 (N_20605,N_20089,N_20269);
and U20606 (N_20606,N_20190,N_20473);
or U20607 (N_20607,N_20114,N_20206);
nor U20608 (N_20608,N_20106,N_20326);
nor U20609 (N_20609,N_20033,N_20417);
or U20610 (N_20610,N_20096,N_20097);
nor U20611 (N_20611,N_20054,N_20169);
nand U20612 (N_20612,N_20397,N_20487);
nand U20613 (N_20613,N_20154,N_20458);
nor U20614 (N_20614,N_20077,N_20483);
or U20615 (N_20615,N_20020,N_20071);
nand U20616 (N_20616,N_20477,N_20314);
and U20617 (N_20617,N_20004,N_20117);
or U20618 (N_20618,N_20499,N_20351);
and U20619 (N_20619,N_20066,N_20490);
and U20620 (N_20620,N_20376,N_20116);
or U20621 (N_20621,N_20093,N_20179);
and U20622 (N_20622,N_20368,N_20311);
nand U20623 (N_20623,N_20348,N_20042);
nand U20624 (N_20624,N_20301,N_20295);
nor U20625 (N_20625,N_20075,N_20041);
and U20626 (N_20626,N_20424,N_20011);
nand U20627 (N_20627,N_20139,N_20270);
nand U20628 (N_20628,N_20339,N_20303);
nand U20629 (N_20629,N_20217,N_20288);
nand U20630 (N_20630,N_20052,N_20494);
or U20631 (N_20631,N_20329,N_20035);
or U20632 (N_20632,N_20493,N_20148);
xor U20633 (N_20633,N_20118,N_20289);
xor U20634 (N_20634,N_20363,N_20409);
and U20635 (N_20635,N_20121,N_20375);
and U20636 (N_20636,N_20321,N_20310);
nor U20637 (N_20637,N_20465,N_20210);
nor U20638 (N_20638,N_20419,N_20198);
and U20639 (N_20639,N_20177,N_20461);
nand U20640 (N_20640,N_20275,N_20385);
nand U20641 (N_20641,N_20396,N_20123);
nand U20642 (N_20642,N_20105,N_20278);
xor U20643 (N_20643,N_20356,N_20360);
or U20644 (N_20644,N_20485,N_20233);
or U20645 (N_20645,N_20330,N_20209);
nor U20646 (N_20646,N_20252,N_20034);
nor U20647 (N_20647,N_20095,N_20263);
and U20648 (N_20648,N_20299,N_20325);
xnor U20649 (N_20649,N_20287,N_20284);
or U20650 (N_20650,N_20489,N_20100);
or U20651 (N_20651,N_20078,N_20176);
xnor U20652 (N_20652,N_20291,N_20293);
nand U20653 (N_20653,N_20195,N_20370);
and U20654 (N_20654,N_20144,N_20080);
xor U20655 (N_20655,N_20125,N_20327);
or U20656 (N_20656,N_20082,N_20173);
xor U20657 (N_20657,N_20272,N_20103);
nor U20658 (N_20658,N_20386,N_20312);
nor U20659 (N_20659,N_20444,N_20039);
or U20660 (N_20660,N_20267,N_20067);
nor U20661 (N_20661,N_20285,N_20124);
xnor U20662 (N_20662,N_20115,N_20341);
nor U20663 (N_20663,N_20449,N_20099);
and U20664 (N_20664,N_20076,N_20491);
or U20665 (N_20665,N_20250,N_20213);
and U20666 (N_20666,N_20274,N_20264);
nand U20667 (N_20667,N_20445,N_20282);
and U20668 (N_20668,N_20002,N_20296);
xnor U20669 (N_20669,N_20132,N_20388);
nand U20670 (N_20670,N_20464,N_20430);
or U20671 (N_20671,N_20048,N_20313);
xnor U20672 (N_20672,N_20024,N_20369);
nand U20673 (N_20673,N_20246,N_20059);
nand U20674 (N_20674,N_20455,N_20194);
nand U20675 (N_20675,N_20142,N_20006);
xor U20676 (N_20676,N_20387,N_20343);
nand U20677 (N_20677,N_20245,N_20027);
nor U20678 (N_20678,N_20391,N_20276);
xor U20679 (N_20679,N_20307,N_20401);
nor U20680 (N_20680,N_20065,N_20480);
nor U20681 (N_20681,N_20186,N_20240);
xnor U20682 (N_20682,N_20379,N_20170);
and U20683 (N_20683,N_20111,N_20029);
nand U20684 (N_20684,N_20346,N_20043);
and U20685 (N_20685,N_20492,N_20128);
nand U20686 (N_20686,N_20166,N_20050);
xor U20687 (N_20687,N_20005,N_20308);
xnor U20688 (N_20688,N_20074,N_20242);
and U20689 (N_20689,N_20028,N_20178);
nand U20690 (N_20690,N_20212,N_20134);
xor U20691 (N_20691,N_20309,N_20126);
or U20692 (N_20692,N_20390,N_20203);
xnor U20693 (N_20693,N_20271,N_20147);
xor U20694 (N_20694,N_20022,N_20266);
xnor U20695 (N_20695,N_20192,N_20305);
nand U20696 (N_20696,N_20185,N_20157);
or U20697 (N_20697,N_20331,N_20364);
nand U20698 (N_20698,N_20136,N_20098);
or U20699 (N_20699,N_20189,N_20110);
nor U20700 (N_20700,N_20038,N_20462);
or U20701 (N_20701,N_20380,N_20241);
and U20702 (N_20702,N_20107,N_20290);
and U20703 (N_20703,N_20322,N_20353);
xor U20704 (N_20704,N_20254,N_20442);
nand U20705 (N_20705,N_20292,N_20051);
and U20706 (N_20706,N_20219,N_20129);
and U20707 (N_20707,N_20431,N_20088);
xnor U20708 (N_20708,N_20069,N_20183);
or U20709 (N_20709,N_20433,N_20130);
xor U20710 (N_20710,N_20220,N_20063);
or U20711 (N_20711,N_20224,N_20045);
and U20712 (N_20712,N_20399,N_20412);
xnor U20713 (N_20713,N_20174,N_20017);
nor U20714 (N_20714,N_20320,N_20087);
or U20715 (N_20715,N_20286,N_20113);
xor U20716 (N_20716,N_20133,N_20392);
xor U20717 (N_20717,N_20304,N_20484);
nand U20718 (N_20718,N_20109,N_20383);
and U20719 (N_20719,N_20300,N_20443);
xnor U20720 (N_20720,N_20395,N_20393);
or U20721 (N_20721,N_20135,N_20475);
or U20722 (N_20722,N_20476,N_20141);
or U20723 (N_20723,N_20000,N_20435);
nand U20724 (N_20724,N_20232,N_20101);
and U20725 (N_20725,N_20182,N_20450);
nor U20726 (N_20726,N_20001,N_20013);
nand U20727 (N_20727,N_20228,N_20471);
nor U20728 (N_20728,N_20167,N_20452);
and U20729 (N_20729,N_20120,N_20204);
nor U20730 (N_20730,N_20221,N_20160);
and U20731 (N_20731,N_20318,N_20092);
nand U20732 (N_20732,N_20064,N_20406);
nand U20733 (N_20733,N_20474,N_20019);
xnor U20734 (N_20734,N_20447,N_20023);
and U20735 (N_20735,N_20352,N_20258);
xor U20736 (N_20736,N_20408,N_20367);
or U20737 (N_20737,N_20436,N_20402);
nor U20738 (N_20738,N_20214,N_20283);
and U20739 (N_20739,N_20328,N_20425);
or U20740 (N_20740,N_20140,N_20347);
xor U20741 (N_20741,N_20030,N_20428);
and U20742 (N_20742,N_20496,N_20342);
nor U20743 (N_20743,N_20466,N_20037);
xnor U20744 (N_20744,N_20009,N_20468);
and U20745 (N_20745,N_20382,N_20207);
nand U20746 (N_20746,N_20268,N_20404);
and U20747 (N_20747,N_20058,N_20146);
xnor U20748 (N_20748,N_20306,N_20016);
xor U20749 (N_20749,N_20403,N_20315);
and U20750 (N_20750,N_20380,N_20369);
or U20751 (N_20751,N_20267,N_20068);
xor U20752 (N_20752,N_20457,N_20093);
nand U20753 (N_20753,N_20290,N_20018);
nor U20754 (N_20754,N_20469,N_20053);
nor U20755 (N_20755,N_20185,N_20003);
nand U20756 (N_20756,N_20422,N_20088);
nand U20757 (N_20757,N_20076,N_20170);
and U20758 (N_20758,N_20362,N_20198);
xor U20759 (N_20759,N_20297,N_20011);
nand U20760 (N_20760,N_20016,N_20142);
nand U20761 (N_20761,N_20394,N_20383);
nor U20762 (N_20762,N_20175,N_20153);
or U20763 (N_20763,N_20339,N_20156);
or U20764 (N_20764,N_20054,N_20066);
or U20765 (N_20765,N_20410,N_20227);
and U20766 (N_20766,N_20249,N_20185);
xnor U20767 (N_20767,N_20409,N_20349);
xnor U20768 (N_20768,N_20221,N_20319);
and U20769 (N_20769,N_20029,N_20319);
nor U20770 (N_20770,N_20493,N_20086);
or U20771 (N_20771,N_20346,N_20050);
xor U20772 (N_20772,N_20129,N_20307);
nor U20773 (N_20773,N_20350,N_20210);
nor U20774 (N_20774,N_20449,N_20351);
xor U20775 (N_20775,N_20317,N_20254);
nor U20776 (N_20776,N_20386,N_20364);
nand U20777 (N_20777,N_20076,N_20023);
xnor U20778 (N_20778,N_20005,N_20335);
or U20779 (N_20779,N_20093,N_20084);
nand U20780 (N_20780,N_20489,N_20356);
nor U20781 (N_20781,N_20004,N_20277);
xnor U20782 (N_20782,N_20076,N_20240);
xor U20783 (N_20783,N_20347,N_20165);
xor U20784 (N_20784,N_20303,N_20266);
or U20785 (N_20785,N_20279,N_20385);
or U20786 (N_20786,N_20374,N_20146);
nand U20787 (N_20787,N_20407,N_20185);
or U20788 (N_20788,N_20140,N_20100);
nor U20789 (N_20789,N_20177,N_20008);
nor U20790 (N_20790,N_20146,N_20479);
nand U20791 (N_20791,N_20318,N_20304);
xnor U20792 (N_20792,N_20234,N_20207);
or U20793 (N_20793,N_20075,N_20280);
nor U20794 (N_20794,N_20300,N_20391);
and U20795 (N_20795,N_20070,N_20400);
nand U20796 (N_20796,N_20055,N_20377);
and U20797 (N_20797,N_20309,N_20474);
xor U20798 (N_20798,N_20442,N_20489);
nor U20799 (N_20799,N_20270,N_20193);
nor U20800 (N_20800,N_20444,N_20287);
and U20801 (N_20801,N_20362,N_20220);
xor U20802 (N_20802,N_20059,N_20422);
or U20803 (N_20803,N_20050,N_20273);
and U20804 (N_20804,N_20241,N_20235);
xnor U20805 (N_20805,N_20162,N_20045);
or U20806 (N_20806,N_20402,N_20327);
nor U20807 (N_20807,N_20013,N_20439);
nor U20808 (N_20808,N_20375,N_20411);
xnor U20809 (N_20809,N_20258,N_20075);
nand U20810 (N_20810,N_20189,N_20137);
or U20811 (N_20811,N_20146,N_20441);
nand U20812 (N_20812,N_20380,N_20345);
and U20813 (N_20813,N_20157,N_20230);
nand U20814 (N_20814,N_20321,N_20171);
or U20815 (N_20815,N_20248,N_20161);
nor U20816 (N_20816,N_20143,N_20400);
nand U20817 (N_20817,N_20336,N_20404);
or U20818 (N_20818,N_20126,N_20009);
nor U20819 (N_20819,N_20091,N_20201);
or U20820 (N_20820,N_20235,N_20103);
nor U20821 (N_20821,N_20474,N_20202);
or U20822 (N_20822,N_20153,N_20178);
nand U20823 (N_20823,N_20137,N_20038);
and U20824 (N_20824,N_20172,N_20252);
or U20825 (N_20825,N_20178,N_20270);
or U20826 (N_20826,N_20151,N_20009);
nand U20827 (N_20827,N_20249,N_20092);
or U20828 (N_20828,N_20081,N_20271);
nor U20829 (N_20829,N_20096,N_20413);
nor U20830 (N_20830,N_20304,N_20092);
nand U20831 (N_20831,N_20163,N_20338);
nand U20832 (N_20832,N_20145,N_20291);
xor U20833 (N_20833,N_20149,N_20403);
and U20834 (N_20834,N_20135,N_20233);
xor U20835 (N_20835,N_20075,N_20334);
nand U20836 (N_20836,N_20405,N_20148);
nor U20837 (N_20837,N_20349,N_20294);
nand U20838 (N_20838,N_20332,N_20206);
nand U20839 (N_20839,N_20385,N_20207);
or U20840 (N_20840,N_20297,N_20454);
and U20841 (N_20841,N_20076,N_20288);
nand U20842 (N_20842,N_20397,N_20414);
or U20843 (N_20843,N_20283,N_20322);
nand U20844 (N_20844,N_20246,N_20456);
or U20845 (N_20845,N_20073,N_20173);
xor U20846 (N_20846,N_20424,N_20277);
and U20847 (N_20847,N_20484,N_20327);
nor U20848 (N_20848,N_20311,N_20113);
and U20849 (N_20849,N_20391,N_20133);
and U20850 (N_20850,N_20070,N_20042);
or U20851 (N_20851,N_20253,N_20434);
nand U20852 (N_20852,N_20361,N_20115);
xor U20853 (N_20853,N_20498,N_20152);
or U20854 (N_20854,N_20459,N_20038);
or U20855 (N_20855,N_20002,N_20023);
nor U20856 (N_20856,N_20065,N_20162);
and U20857 (N_20857,N_20341,N_20057);
nand U20858 (N_20858,N_20413,N_20479);
nor U20859 (N_20859,N_20405,N_20128);
and U20860 (N_20860,N_20341,N_20130);
nand U20861 (N_20861,N_20147,N_20062);
xor U20862 (N_20862,N_20317,N_20138);
nor U20863 (N_20863,N_20451,N_20039);
nand U20864 (N_20864,N_20091,N_20262);
or U20865 (N_20865,N_20116,N_20037);
and U20866 (N_20866,N_20019,N_20240);
or U20867 (N_20867,N_20226,N_20183);
and U20868 (N_20868,N_20201,N_20448);
or U20869 (N_20869,N_20337,N_20405);
or U20870 (N_20870,N_20107,N_20499);
nand U20871 (N_20871,N_20179,N_20448);
nand U20872 (N_20872,N_20281,N_20133);
xnor U20873 (N_20873,N_20498,N_20409);
or U20874 (N_20874,N_20107,N_20198);
and U20875 (N_20875,N_20149,N_20386);
nor U20876 (N_20876,N_20086,N_20438);
nand U20877 (N_20877,N_20426,N_20362);
xor U20878 (N_20878,N_20179,N_20043);
xor U20879 (N_20879,N_20204,N_20412);
nand U20880 (N_20880,N_20003,N_20133);
xor U20881 (N_20881,N_20479,N_20328);
or U20882 (N_20882,N_20369,N_20165);
or U20883 (N_20883,N_20102,N_20482);
and U20884 (N_20884,N_20386,N_20363);
or U20885 (N_20885,N_20354,N_20198);
nand U20886 (N_20886,N_20168,N_20174);
xor U20887 (N_20887,N_20372,N_20010);
xor U20888 (N_20888,N_20233,N_20122);
nor U20889 (N_20889,N_20366,N_20040);
or U20890 (N_20890,N_20095,N_20027);
and U20891 (N_20891,N_20429,N_20035);
or U20892 (N_20892,N_20366,N_20447);
or U20893 (N_20893,N_20272,N_20432);
or U20894 (N_20894,N_20113,N_20044);
or U20895 (N_20895,N_20079,N_20085);
or U20896 (N_20896,N_20071,N_20226);
xnor U20897 (N_20897,N_20244,N_20103);
nor U20898 (N_20898,N_20343,N_20215);
nor U20899 (N_20899,N_20110,N_20303);
and U20900 (N_20900,N_20481,N_20009);
nor U20901 (N_20901,N_20290,N_20214);
nor U20902 (N_20902,N_20233,N_20067);
xor U20903 (N_20903,N_20075,N_20036);
or U20904 (N_20904,N_20385,N_20408);
nand U20905 (N_20905,N_20440,N_20107);
xnor U20906 (N_20906,N_20450,N_20369);
and U20907 (N_20907,N_20197,N_20476);
or U20908 (N_20908,N_20396,N_20313);
or U20909 (N_20909,N_20434,N_20294);
nand U20910 (N_20910,N_20490,N_20343);
and U20911 (N_20911,N_20047,N_20301);
nor U20912 (N_20912,N_20206,N_20417);
nor U20913 (N_20913,N_20061,N_20323);
xor U20914 (N_20914,N_20154,N_20031);
nor U20915 (N_20915,N_20487,N_20160);
xor U20916 (N_20916,N_20271,N_20128);
and U20917 (N_20917,N_20266,N_20174);
or U20918 (N_20918,N_20417,N_20172);
or U20919 (N_20919,N_20239,N_20030);
nand U20920 (N_20920,N_20360,N_20011);
xor U20921 (N_20921,N_20009,N_20099);
xnor U20922 (N_20922,N_20359,N_20003);
xnor U20923 (N_20923,N_20473,N_20135);
and U20924 (N_20924,N_20080,N_20402);
nor U20925 (N_20925,N_20264,N_20437);
or U20926 (N_20926,N_20324,N_20318);
and U20927 (N_20927,N_20233,N_20138);
nand U20928 (N_20928,N_20039,N_20215);
nand U20929 (N_20929,N_20377,N_20291);
and U20930 (N_20930,N_20107,N_20241);
nor U20931 (N_20931,N_20413,N_20374);
xnor U20932 (N_20932,N_20100,N_20346);
or U20933 (N_20933,N_20243,N_20318);
or U20934 (N_20934,N_20263,N_20298);
nand U20935 (N_20935,N_20396,N_20248);
nand U20936 (N_20936,N_20022,N_20097);
nor U20937 (N_20937,N_20305,N_20474);
nor U20938 (N_20938,N_20038,N_20189);
and U20939 (N_20939,N_20202,N_20350);
or U20940 (N_20940,N_20100,N_20236);
and U20941 (N_20941,N_20139,N_20245);
nand U20942 (N_20942,N_20151,N_20026);
nand U20943 (N_20943,N_20291,N_20287);
nor U20944 (N_20944,N_20355,N_20083);
and U20945 (N_20945,N_20395,N_20364);
xnor U20946 (N_20946,N_20237,N_20366);
nor U20947 (N_20947,N_20375,N_20334);
nor U20948 (N_20948,N_20058,N_20236);
nand U20949 (N_20949,N_20290,N_20352);
nor U20950 (N_20950,N_20066,N_20087);
xnor U20951 (N_20951,N_20479,N_20114);
and U20952 (N_20952,N_20196,N_20115);
or U20953 (N_20953,N_20115,N_20281);
and U20954 (N_20954,N_20225,N_20390);
nand U20955 (N_20955,N_20106,N_20173);
and U20956 (N_20956,N_20268,N_20168);
and U20957 (N_20957,N_20123,N_20074);
and U20958 (N_20958,N_20416,N_20376);
and U20959 (N_20959,N_20025,N_20303);
nand U20960 (N_20960,N_20460,N_20258);
and U20961 (N_20961,N_20080,N_20444);
nor U20962 (N_20962,N_20472,N_20177);
xnor U20963 (N_20963,N_20434,N_20101);
xnor U20964 (N_20964,N_20145,N_20167);
nor U20965 (N_20965,N_20055,N_20385);
nor U20966 (N_20966,N_20251,N_20270);
and U20967 (N_20967,N_20285,N_20136);
xor U20968 (N_20968,N_20265,N_20058);
nor U20969 (N_20969,N_20038,N_20266);
nand U20970 (N_20970,N_20119,N_20356);
nand U20971 (N_20971,N_20473,N_20166);
or U20972 (N_20972,N_20312,N_20205);
nand U20973 (N_20973,N_20392,N_20090);
nand U20974 (N_20974,N_20105,N_20069);
nor U20975 (N_20975,N_20323,N_20009);
nor U20976 (N_20976,N_20110,N_20332);
and U20977 (N_20977,N_20472,N_20356);
nand U20978 (N_20978,N_20211,N_20475);
and U20979 (N_20979,N_20308,N_20412);
or U20980 (N_20980,N_20265,N_20306);
and U20981 (N_20981,N_20079,N_20133);
xnor U20982 (N_20982,N_20055,N_20493);
nor U20983 (N_20983,N_20078,N_20443);
and U20984 (N_20984,N_20459,N_20463);
xnor U20985 (N_20985,N_20249,N_20060);
and U20986 (N_20986,N_20027,N_20258);
or U20987 (N_20987,N_20228,N_20352);
nor U20988 (N_20988,N_20431,N_20394);
or U20989 (N_20989,N_20006,N_20206);
nor U20990 (N_20990,N_20063,N_20190);
or U20991 (N_20991,N_20031,N_20249);
nor U20992 (N_20992,N_20407,N_20229);
nor U20993 (N_20993,N_20076,N_20405);
nor U20994 (N_20994,N_20043,N_20273);
xor U20995 (N_20995,N_20253,N_20249);
and U20996 (N_20996,N_20077,N_20473);
xor U20997 (N_20997,N_20277,N_20182);
nand U20998 (N_20998,N_20106,N_20049);
and U20999 (N_20999,N_20288,N_20422);
and U21000 (N_21000,N_20974,N_20946);
xnor U21001 (N_21001,N_20864,N_20569);
or U21002 (N_21002,N_20952,N_20942);
nor U21003 (N_21003,N_20763,N_20689);
nand U21004 (N_21004,N_20891,N_20806);
or U21005 (N_21005,N_20945,N_20798);
nor U21006 (N_21006,N_20516,N_20783);
nand U21007 (N_21007,N_20660,N_20838);
nand U21008 (N_21008,N_20672,N_20653);
nor U21009 (N_21009,N_20543,N_20991);
nor U21010 (N_21010,N_20764,N_20833);
and U21011 (N_21011,N_20898,N_20500);
and U21012 (N_21012,N_20614,N_20926);
nor U21013 (N_21013,N_20998,N_20828);
nand U21014 (N_21014,N_20649,N_20507);
and U21015 (N_21015,N_20884,N_20585);
and U21016 (N_21016,N_20757,N_20754);
nand U21017 (N_21017,N_20743,N_20862);
or U21018 (N_21018,N_20954,N_20613);
or U21019 (N_21019,N_20847,N_20697);
nand U21020 (N_21020,N_20785,N_20762);
and U21021 (N_21021,N_20981,N_20997);
and U21022 (N_21022,N_20963,N_20667);
and U21023 (N_21023,N_20694,N_20666);
or U21024 (N_21024,N_20524,N_20662);
nor U21025 (N_21025,N_20896,N_20531);
nor U21026 (N_21026,N_20618,N_20724);
nand U21027 (N_21027,N_20540,N_20685);
xnor U21028 (N_21028,N_20705,N_20506);
and U21029 (N_21029,N_20652,N_20753);
xor U21030 (N_21030,N_20959,N_20987);
nand U21031 (N_21031,N_20525,N_20789);
nand U21032 (N_21032,N_20835,N_20821);
or U21033 (N_21033,N_20645,N_20633);
or U21034 (N_21034,N_20573,N_20819);
or U21035 (N_21035,N_20804,N_20912);
xnor U21036 (N_21036,N_20986,N_20751);
and U21037 (N_21037,N_20583,N_20669);
and U21038 (N_21038,N_20950,N_20736);
or U21039 (N_21039,N_20608,N_20599);
or U21040 (N_21040,N_20831,N_20880);
xor U21041 (N_21041,N_20933,N_20801);
nand U21042 (N_21042,N_20809,N_20871);
or U21043 (N_21043,N_20542,N_20714);
nor U21044 (N_21044,N_20554,N_20841);
or U21045 (N_21045,N_20641,N_20853);
or U21046 (N_21046,N_20590,N_20953);
or U21047 (N_21047,N_20843,N_20834);
nor U21048 (N_21048,N_20882,N_20899);
and U21049 (N_21049,N_20577,N_20934);
nor U21050 (N_21050,N_20975,N_20519);
and U21051 (N_21051,N_20750,N_20568);
and U21052 (N_21052,N_20962,N_20990);
xor U21053 (N_21053,N_20536,N_20917);
nor U21054 (N_21054,N_20670,N_20802);
or U21055 (N_21055,N_20854,N_20676);
and U21056 (N_21056,N_20812,N_20777);
nor U21057 (N_21057,N_20772,N_20883);
and U21058 (N_21058,N_20897,N_20984);
nor U21059 (N_21059,N_20627,N_20687);
and U21060 (N_21060,N_20696,N_20948);
nand U21061 (N_21061,N_20617,N_20541);
xnor U21062 (N_21062,N_20707,N_20589);
and U21063 (N_21063,N_20730,N_20539);
nor U21064 (N_21064,N_20867,N_20513);
or U21065 (N_21065,N_20682,N_20521);
and U21066 (N_21066,N_20570,N_20745);
or U21067 (N_21067,N_20787,N_20877);
and U21068 (N_21068,N_20739,N_20992);
nor U21069 (N_21069,N_20747,N_20935);
nor U21070 (N_21070,N_20678,N_20767);
nor U21071 (N_21071,N_20983,N_20501);
nor U21072 (N_21072,N_20718,N_20994);
nor U21073 (N_21073,N_20795,N_20921);
nand U21074 (N_21074,N_20550,N_20929);
or U21075 (N_21075,N_20563,N_20927);
nand U21076 (N_21076,N_20901,N_20702);
or U21077 (N_21077,N_20559,N_20624);
xor U21078 (N_21078,N_20856,N_20961);
nor U21079 (N_21079,N_20786,N_20910);
xnor U21080 (N_21080,N_20607,N_20911);
or U21081 (N_21081,N_20596,N_20700);
and U21082 (N_21082,N_20947,N_20842);
xor U21083 (N_21083,N_20909,N_20560);
or U21084 (N_21084,N_20977,N_20870);
nand U21085 (N_21085,N_20887,N_20729);
nor U21086 (N_21086,N_20965,N_20837);
and U21087 (N_21087,N_20868,N_20879);
nor U21088 (N_21088,N_20619,N_20788);
and U21089 (N_21089,N_20936,N_20611);
nand U21090 (N_21090,N_20567,N_20744);
or U21091 (N_21091,N_20593,N_20551);
or U21092 (N_21092,N_20978,N_20527);
or U21093 (N_21093,N_20562,N_20532);
nor U21094 (N_21094,N_20858,N_20720);
and U21095 (N_21095,N_20900,N_20979);
nor U21096 (N_21096,N_20875,N_20919);
nand U21097 (N_21097,N_20646,N_20794);
or U21098 (N_21098,N_20661,N_20930);
nand U21099 (N_21099,N_20626,N_20579);
xnor U21100 (N_21100,N_20761,N_20711);
nor U21101 (N_21101,N_20612,N_20918);
or U21102 (N_21102,N_20733,N_20811);
or U21103 (N_21103,N_20874,N_20591);
xnor U21104 (N_21104,N_20615,N_20658);
xnor U21105 (N_21105,N_20985,N_20634);
xnor U21106 (N_21106,N_20640,N_20938);
xor U21107 (N_21107,N_20620,N_20647);
nand U21108 (N_21108,N_20920,N_20748);
nand U21109 (N_21109,N_20616,N_20712);
and U21110 (N_21110,N_20749,N_20972);
or U21111 (N_21111,N_20876,N_20576);
or U21112 (N_21112,N_20999,N_20903);
or U21113 (N_21113,N_20863,N_20517);
or U21114 (N_21114,N_20737,N_20564);
or U21115 (N_21115,N_20932,N_20886);
and U21116 (N_21116,N_20807,N_20957);
or U21117 (N_21117,N_20703,N_20873);
nor U21118 (N_21118,N_20504,N_20771);
xor U21119 (N_21119,N_20851,N_20755);
nand U21120 (N_21120,N_20695,N_20655);
and U21121 (N_21121,N_20547,N_20699);
nor U21122 (N_21122,N_20820,N_20818);
xor U21123 (N_21123,N_20782,N_20629);
nor U21124 (N_21124,N_20625,N_20849);
and U21125 (N_21125,N_20826,N_20578);
and U21126 (N_21126,N_20816,N_20955);
xnor U21127 (N_21127,N_20530,N_20925);
and U21128 (N_21128,N_20698,N_20905);
nor U21129 (N_21129,N_20878,N_20836);
or U21130 (N_21130,N_20769,N_20810);
and U21131 (N_21131,N_20956,N_20928);
xnor U21132 (N_21132,N_20549,N_20759);
nor U21133 (N_21133,N_20502,N_20723);
and U21134 (N_21134,N_20690,N_20722);
and U21135 (N_21135,N_20889,N_20731);
nand U21136 (N_21136,N_20916,N_20553);
or U21137 (N_21137,N_20717,N_20824);
xor U21138 (N_21138,N_20790,N_20888);
xnor U21139 (N_21139,N_20844,N_20894);
xnor U21140 (N_21140,N_20857,N_20728);
or U21141 (N_21141,N_20779,N_20859);
xor U21142 (N_21142,N_20893,N_20943);
and U21143 (N_21143,N_20631,N_20719);
xor U21144 (N_21144,N_20840,N_20555);
nand U21145 (N_21145,N_20881,N_20691);
and U21146 (N_21146,N_20522,N_20684);
nor U21147 (N_21147,N_20914,N_20587);
and U21148 (N_21148,N_20915,N_20832);
or U21149 (N_21149,N_20566,N_20904);
nor U21150 (N_21150,N_20715,N_20605);
nand U21151 (N_21151,N_20931,N_20701);
and U21152 (N_21152,N_20580,N_20738);
xnor U21153 (N_21153,N_20637,N_20970);
and U21154 (N_21154,N_20823,N_20621);
nor U21155 (N_21155,N_20581,N_20964);
nand U21156 (N_21156,N_20708,N_20855);
xnor U21157 (N_21157,N_20546,N_20815);
or U21158 (N_21158,N_20982,N_20677);
nor U21159 (N_21159,N_20575,N_20852);
and U21160 (N_21160,N_20512,N_20845);
xor U21161 (N_21161,N_20776,N_20941);
nand U21162 (N_21162,N_20528,N_20805);
nand U21163 (N_21163,N_20535,N_20969);
or U21164 (N_21164,N_20800,N_20860);
nor U21165 (N_21165,N_20907,N_20628);
nor U21166 (N_21166,N_20503,N_20830);
and U21167 (N_21167,N_20869,N_20692);
nand U21168 (N_21168,N_20780,N_20817);
and U21169 (N_21169,N_20538,N_20526);
and U21170 (N_21170,N_20598,N_20674);
xor U21171 (N_21171,N_20773,N_20681);
nor U21172 (N_21172,N_20890,N_20713);
nor U21173 (N_21173,N_20993,N_20996);
and U21174 (N_21174,N_20586,N_20924);
nand U21175 (N_21175,N_20520,N_20995);
or U21176 (N_21176,N_20545,N_20556);
xnor U21177 (N_21177,N_20534,N_20584);
or U21178 (N_21178,N_20768,N_20958);
and U21179 (N_21179,N_20727,N_20797);
or U21180 (N_21180,N_20688,N_20709);
and U21181 (N_21181,N_20537,N_20732);
and U21182 (N_21182,N_20663,N_20980);
nor U21183 (N_21183,N_20518,N_20778);
xor U21184 (N_21184,N_20650,N_20659);
and U21185 (N_21185,N_20505,N_20735);
nand U21186 (N_21186,N_20671,N_20923);
xor U21187 (N_21187,N_20572,N_20865);
nor U21188 (N_21188,N_20604,N_20508);
nor U21189 (N_21189,N_20758,N_20648);
xnor U21190 (N_21190,N_20827,N_20796);
nor U21191 (N_21191,N_20594,N_20664);
nor U21192 (N_21192,N_20511,N_20574);
or U21193 (N_21193,N_20710,N_20937);
nor U21194 (N_21194,N_20793,N_20630);
xor U21195 (N_21195,N_20951,N_20922);
nand U21196 (N_21196,N_20571,N_20639);
nor U21197 (N_21197,N_20673,N_20784);
xnor U21198 (N_21198,N_20552,N_20741);
or U21199 (N_21199,N_20746,N_20622);
xnor U21200 (N_21200,N_20726,N_20765);
and U21201 (N_21201,N_20775,N_20989);
or U21202 (N_21202,N_20734,N_20839);
xnor U21203 (N_21203,N_20940,N_20861);
and U21204 (N_21204,N_20792,N_20623);
and U21205 (N_21205,N_20668,N_20548);
or U21206 (N_21206,N_20600,N_20636);
nor U21207 (N_21207,N_20866,N_20803);
or U21208 (N_21208,N_20892,N_20610);
or U21209 (N_21209,N_20638,N_20561);
or U21210 (N_21210,N_20848,N_20635);
nor U21211 (N_21211,N_20665,N_20514);
xnor U21212 (N_21212,N_20725,N_20523);
xnor U21213 (N_21213,N_20595,N_20601);
nand U21214 (N_21214,N_20683,N_20825);
xor U21215 (N_21215,N_20971,N_20704);
xor U21216 (N_21216,N_20960,N_20814);
nor U21217 (N_21217,N_20885,N_20770);
nand U21218 (N_21218,N_20557,N_20643);
xor U21219 (N_21219,N_20654,N_20592);
or U21220 (N_21220,N_20609,N_20752);
nor U21221 (N_21221,N_20509,N_20774);
and U21222 (N_21222,N_20693,N_20515);
or U21223 (N_21223,N_20988,N_20675);
and U21224 (N_21224,N_20642,N_20606);
nor U21225 (N_21225,N_20632,N_20657);
xor U21226 (N_21226,N_20680,N_20967);
nor U21227 (N_21227,N_20902,N_20906);
nor U21228 (N_21228,N_20949,N_20742);
xnor U21229 (N_21229,N_20944,N_20968);
nand U21230 (N_21230,N_20822,N_20756);
xnor U21231 (N_21231,N_20740,N_20686);
nand U21232 (N_21232,N_20597,N_20808);
nand U21233 (N_21233,N_20644,N_20939);
and U21234 (N_21234,N_20588,N_20721);
and U21235 (N_21235,N_20813,N_20966);
nand U21236 (N_21236,N_20565,N_20706);
xnor U21237 (N_21237,N_20850,N_20760);
nor U21238 (N_21238,N_20679,N_20766);
and U21239 (N_21239,N_20651,N_20716);
or U21240 (N_21240,N_20544,N_20510);
xnor U21241 (N_21241,N_20582,N_20846);
nand U21242 (N_21242,N_20603,N_20558);
or U21243 (N_21243,N_20781,N_20529);
nand U21244 (N_21244,N_20973,N_20976);
nor U21245 (N_21245,N_20895,N_20791);
and U21246 (N_21246,N_20656,N_20829);
and U21247 (N_21247,N_20533,N_20908);
or U21248 (N_21248,N_20872,N_20799);
nor U21249 (N_21249,N_20913,N_20602);
xnor U21250 (N_21250,N_20872,N_20926);
or U21251 (N_21251,N_20957,N_20573);
or U21252 (N_21252,N_20818,N_20724);
and U21253 (N_21253,N_20882,N_20546);
nand U21254 (N_21254,N_20540,N_20558);
and U21255 (N_21255,N_20707,N_20954);
nor U21256 (N_21256,N_20708,N_20563);
or U21257 (N_21257,N_20996,N_20685);
nor U21258 (N_21258,N_20936,N_20800);
nor U21259 (N_21259,N_20710,N_20673);
or U21260 (N_21260,N_20735,N_20611);
nand U21261 (N_21261,N_20942,N_20761);
xnor U21262 (N_21262,N_20588,N_20785);
xor U21263 (N_21263,N_20807,N_20713);
or U21264 (N_21264,N_20826,N_20852);
and U21265 (N_21265,N_20502,N_20640);
and U21266 (N_21266,N_20971,N_20791);
nor U21267 (N_21267,N_20877,N_20536);
nor U21268 (N_21268,N_20561,N_20593);
xor U21269 (N_21269,N_20995,N_20579);
nor U21270 (N_21270,N_20857,N_20566);
and U21271 (N_21271,N_20577,N_20989);
nor U21272 (N_21272,N_20824,N_20705);
or U21273 (N_21273,N_20847,N_20553);
or U21274 (N_21274,N_20971,N_20867);
nand U21275 (N_21275,N_20592,N_20563);
nor U21276 (N_21276,N_20975,N_20938);
nand U21277 (N_21277,N_20601,N_20689);
and U21278 (N_21278,N_20913,N_20729);
or U21279 (N_21279,N_20917,N_20545);
and U21280 (N_21280,N_20858,N_20561);
xnor U21281 (N_21281,N_20532,N_20697);
nand U21282 (N_21282,N_20713,N_20676);
nor U21283 (N_21283,N_20982,N_20999);
nand U21284 (N_21284,N_20775,N_20922);
or U21285 (N_21285,N_20660,N_20672);
or U21286 (N_21286,N_20865,N_20645);
and U21287 (N_21287,N_20672,N_20900);
or U21288 (N_21288,N_20800,N_20708);
nor U21289 (N_21289,N_20695,N_20893);
nor U21290 (N_21290,N_20638,N_20776);
nor U21291 (N_21291,N_20591,N_20695);
nand U21292 (N_21292,N_20625,N_20812);
nand U21293 (N_21293,N_20946,N_20881);
nand U21294 (N_21294,N_20589,N_20624);
and U21295 (N_21295,N_20837,N_20579);
xnor U21296 (N_21296,N_20624,N_20564);
nand U21297 (N_21297,N_20915,N_20799);
nand U21298 (N_21298,N_20875,N_20540);
and U21299 (N_21299,N_20668,N_20740);
xor U21300 (N_21300,N_20763,N_20704);
nor U21301 (N_21301,N_20529,N_20827);
and U21302 (N_21302,N_20998,N_20814);
xor U21303 (N_21303,N_20773,N_20882);
or U21304 (N_21304,N_20592,N_20636);
and U21305 (N_21305,N_20617,N_20978);
or U21306 (N_21306,N_20899,N_20569);
or U21307 (N_21307,N_20936,N_20970);
nor U21308 (N_21308,N_20512,N_20883);
nand U21309 (N_21309,N_20575,N_20677);
and U21310 (N_21310,N_20566,N_20744);
nand U21311 (N_21311,N_20774,N_20927);
xor U21312 (N_21312,N_20869,N_20898);
nor U21313 (N_21313,N_20807,N_20614);
or U21314 (N_21314,N_20796,N_20816);
or U21315 (N_21315,N_20645,N_20844);
and U21316 (N_21316,N_20814,N_20779);
xor U21317 (N_21317,N_20715,N_20573);
nor U21318 (N_21318,N_20761,N_20661);
or U21319 (N_21319,N_20778,N_20629);
xor U21320 (N_21320,N_20882,N_20772);
nor U21321 (N_21321,N_20758,N_20733);
and U21322 (N_21322,N_20585,N_20629);
xnor U21323 (N_21323,N_20995,N_20875);
or U21324 (N_21324,N_20880,N_20927);
nand U21325 (N_21325,N_20681,N_20519);
and U21326 (N_21326,N_20732,N_20615);
or U21327 (N_21327,N_20814,N_20576);
nor U21328 (N_21328,N_20666,N_20849);
and U21329 (N_21329,N_20903,N_20737);
and U21330 (N_21330,N_20974,N_20923);
nand U21331 (N_21331,N_20507,N_20596);
or U21332 (N_21332,N_20852,N_20994);
or U21333 (N_21333,N_20877,N_20671);
or U21334 (N_21334,N_20739,N_20673);
xor U21335 (N_21335,N_20937,N_20687);
nand U21336 (N_21336,N_20836,N_20808);
xor U21337 (N_21337,N_20968,N_20982);
nor U21338 (N_21338,N_20601,N_20763);
nand U21339 (N_21339,N_20699,N_20954);
nor U21340 (N_21340,N_20883,N_20765);
xor U21341 (N_21341,N_20899,N_20677);
and U21342 (N_21342,N_20767,N_20974);
xnor U21343 (N_21343,N_20655,N_20855);
nor U21344 (N_21344,N_20662,N_20644);
and U21345 (N_21345,N_20532,N_20577);
xnor U21346 (N_21346,N_20947,N_20744);
or U21347 (N_21347,N_20897,N_20590);
nand U21348 (N_21348,N_20530,N_20890);
xnor U21349 (N_21349,N_20895,N_20985);
nor U21350 (N_21350,N_20670,N_20631);
or U21351 (N_21351,N_20784,N_20905);
nand U21352 (N_21352,N_20696,N_20639);
nor U21353 (N_21353,N_20984,N_20759);
nand U21354 (N_21354,N_20664,N_20822);
nand U21355 (N_21355,N_20929,N_20976);
nor U21356 (N_21356,N_20700,N_20953);
xor U21357 (N_21357,N_20991,N_20730);
nand U21358 (N_21358,N_20768,N_20897);
nand U21359 (N_21359,N_20998,N_20831);
xor U21360 (N_21360,N_20573,N_20997);
nand U21361 (N_21361,N_20774,N_20770);
or U21362 (N_21362,N_20848,N_20674);
nand U21363 (N_21363,N_20729,N_20619);
nor U21364 (N_21364,N_20739,N_20789);
or U21365 (N_21365,N_20669,N_20642);
nor U21366 (N_21366,N_20667,N_20628);
nand U21367 (N_21367,N_20500,N_20549);
nand U21368 (N_21368,N_20751,N_20638);
and U21369 (N_21369,N_20696,N_20905);
or U21370 (N_21370,N_20946,N_20600);
and U21371 (N_21371,N_20772,N_20754);
or U21372 (N_21372,N_20613,N_20908);
nor U21373 (N_21373,N_20950,N_20969);
or U21374 (N_21374,N_20812,N_20725);
or U21375 (N_21375,N_20782,N_20529);
and U21376 (N_21376,N_20564,N_20522);
or U21377 (N_21377,N_20519,N_20661);
xor U21378 (N_21378,N_20659,N_20856);
nor U21379 (N_21379,N_20672,N_20526);
or U21380 (N_21380,N_20669,N_20636);
nand U21381 (N_21381,N_20610,N_20678);
xnor U21382 (N_21382,N_20755,N_20680);
xnor U21383 (N_21383,N_20502,N_20518);
nor U21384 (N_21384,N_20728,N_20999);
xnor U21385 (N_21385,N_20806,N_20699);
and U21386 (N_21386,N_20575,N_20711);
or U21387 (N_21387,N_20722,N_20869);
xor U21388 (N_21388,N_20585,N_20506);
and U21389 (N_21389,N_20532,N_20738);
xor U21390 (N_21390,N_20864,N_20514);
nor U21391 (N_21391,N_20768,N_20535);
and U21392 (N_21392,N_20757,N_20730);
xor U21393 (N_21393,N_20711,N_20853);
nor U21394 (N_21394,N_20552,N_20845);
or U21395 (N_21395,N_20792,N_20679);
nor U21396 (N_21396,N_20588,N_20856);
nor U21397 (N_21397,N_20851,N_20907);
xnor U21398 (N_21398,N_20783,N_20824);
nor U21399 (N_21399,N_20503,N_20659);
or U21400 (N_21400,N_20891,N_20562);
and U21401 (N_21401,N_20627,N_20879);
xnor U21402 (N_21402,N_20949,N_20660);
nand U21403 (N_21403,N_20701,N_20722);
nand U21404 (N_21404,N_20513,N_20584);
nor U21405 (N_21405,N_20684,N_20813);
and U21406 (N_21406,N_20806,N_20695);
nor U21407 (N_21407,N_20977,N_20728);
and U21408 (N_21408,N_20740,N_20921);
or U21409 (N_21409,N_20667,N_20725);
nand U21410 (N_21410,N_20922,N_20880);
nor U21411 (N_21411,N_20880,N_20591);
nand U21412 (N_21412,N_20762,N_20943);
nor U21413 (N_21413,N_20698,N_20773);
nand U21414 (N_21414,N_20908,N_20575);
or U21415 (N_21415,N_20574,N_20891);
xnor U21416 (N_21416,N_20528,N_20619);
nand U21417 (N_21417,N_20831,N_20731);
xnor U21418 (N_21418,N_20641,N_20537);
xnor U21419 (N_21419,N_20853,N_20741);
nor U21420 (N_21420,N_20763,N_20906);
nand U21421 (N_21421,N_20836,N_20843);
nor U21422 (N_21422,N_20791,N_20615);
or U21423 (N_21423,N_20903,N_20776);
nor U21424 (N_21424,N_20595,N_20524);
and U21425 (N_21425,N_20724,N_20880);
xnor U21426 (N_21426,N_20899,N_20758);
xor U21427 (N_21427,N_20718,N_20876);
xnor U21428 (N_21428,N_20951,N_20587);
xor U21429 (N_21429,N_20560,N_20766);
or U21430 (N_21430,N_20878,N_20601);
and U21431 (N_21431,N_20711,N_20913);
xnor U21432 (N_21432,N_20600,N_20897);
or U21433 (N_21433,N_20846,N_20773);
nor U21434 (N_21434,N_20669,N_20610);
nor U21435 (N_21435,N_20885,N_20951);
nand U21436 (N_21436,N_20873,N_20714);
nand U21437 (N_21437,N_20935,N_20796);
and U21438 (N_21438,N_20699,N_20857);
nand U21439 (N_21439,N_20871,N_20748);
or U21440 (N_21440,N_20500,N_20636);
or U21441 (N_21441,N_20980,N_20910);
and U21442 (N_21442,N_20678,N_20756);
xor U21443 (N_21443,N_20960,N_20605);
nand U21444 (N_21444,N_20599,N_20547);
nand U21445 (N_21445,N_20817,N_20562);
xor U21446 (N_21446,N_20831,N_20765);
xor U21447 (N_21447,N_20519,N_20676);
or U21448 (N_21448,N_20868,N_20883);
nand U21449 (N_21449,N_20955,N_20995);
and U21450 (N_21450,N_20562,N_20690);
or U21451 (N_21451,N_20655,N_20542);
nand U21452 (N_21452,N_20812,N_20907);
xnor U21453 (N_21453,N_20785,N_20647);
xnor U21454 (N_21454,N_20755,N_20878);
or U21455 (N_21455,N_20893,N_20552);
xor U21456 (N_21456,N_20736,N_20867);
and U21457 (N_21457,N_20724,N_20649);
nand U21458 (N_21458,N_20814,N_20839);
and U21459 (N_21459,N_20617,N_20627);
and U21460 (N_21460,N_20642,N_20763);
nor U21461 (N_21461,N_20989,N_20883);
or U21462 (N_21462,N_20769,N_20842);
xor U21463 (N_21463,N_20654,N_20572);
nand U21464 (N_21464,N_20837,N_20888);
nor U21465 (N_21465,N_20627,N_20885);
nand U21466 (N_21466,N_20893,N_20842);
nand U21467 (N_21467,N_20778,N_20717);
nand U21468 (N_21468,N_20580,N_20841);
and U21469 (N_21469,N_20758,N_20951);
nor U21470 (N_21470,N_20658,N_20853);
and U21471 (N_21471,N_20542,N_20711);
or U21472 (N_21472,N_20527,N_20592);
nor U21473 (N_21473,N_20764,N_20950);
or U21474 (N_21474,N_20668,N_20841);
xor U21475 (N_21475,N_20947,N_20726);
or U21476 (N_21476,N_20971,N_20554);
or U21477 (N_21477,N_20765,N_20794);
or U21478 (N_21478,N_20940,N_20939);
and U21479 (N_21479,N_20805,N_20787);
nand U21480 (N_21480,N_20751,N_20628);
and U21481 (N_21481,N_20939,N_20983);
xnor U21482 (N_21482,N_20705,N_20561);
and U21483 (N_21483,N_20541,N_20570);
nand U21484 (N_21484,N_20769,N_20716);
and U21485 (N_21485,N_20660,N_20531);
nand U21486 (N_21486,N_20702,N_20509);
or U21487 (N_21487,N_20944,N_20847);
and U21488 (N_21488,N_20523,N_20825);
nand U21489 (N_21489,N_20532,N_20901);
nor U21490 (N_21490,N_20865,N_20996);
and U21491 (N_21491,N_20597,N_20947);
and U21492 (N_21492,N_20740,N_20518);
or U21493 (N_21493,N_20739,N_20871);
nand U21494 (N_21494,N_20915,N_20517);
xor U21495 (N_21495,N_20628,N_20549);
nor U21496 (N_21496,N_20703,N_20609);
nor U21497 (N_21497,N_20663,N_20995);
xor U21498 (N_21498,N_20854,N_20760);
and U21499 (N_21499,N_20921,N_20524);
or U21500 (N_21500,N_21291,N_21322);
nand U21501 (N_21501,N_21454,N_21311);
and U21502 (N_21502,N_21038,N_21212);
nor U21503 (N_21503,N_21470,N_21211);
xor U21504 (N_21504,N_21115,N_21191);
nor U21505 (N_21505,N_21298,N_21032);
or U21506 (N_21506,N_21175,N_21315);
nor U21507 (N_21507,N_21339,N_21067);
nand U21508 (N_21508,N_21331,N_21147);
and U21509 (N_21509,N_21114,N_21479);
or U21510 (N_21510,N_21320,N_21371);
xor U21511 (N_21511,N_21453,N_21409);
xor U21512 (N_21512,N_21113,N_21351);
nor U21513 (N_21513,N_21436,N_21194);
xor U21514 (N_21514,N_21233,N_21046);
and U21515 (N_21515,N_21309,N_21183);
xor U21516 (N_21516,N_21262,N_21145);
and U21517 (N_21517,N_21099,N_21077);
or U21518 (N_21518,N_21009,N_21310);
or U21519 (N_21519,N_21134,N_21109);
and U21520 (N_21520,N_21196,N_21429);
xnor U21521 (N_21521,N_21120,N_21078);
xnor U21522 (N_21522,N_21422,N_21079);
and U21523 (N_21523,N_21057,N_21138);
xor U21524 (N_21524,N_21345,N_21403);
xnor U21525 (N_21525,N_21283,N_21049);
and U21526 (N_21526,N_21158,N_21313);
nor U21527 (N_21527,N_21110,N_21438);
or U21528 (N_21528,N_21228,N_21102);
or U21529 (N_21529,N_21256,N_21001);
xor U21530 (N_21530,N_21463,N_21491);
or U21531 (N_21531,N_21308,N_21307);
nand U21532 (N_21532,N_21237,N_21368);
nand U21533 (N_21533,N_21035,N_21073);
or U21534 (N_21534,N_21445,N_21280);
nor U21535 (N_21535,N_21444,N_21330);
nand U21536 (N_21536,N_21384,N_21433);
nor U21537 (N_21537,N_21162,N_21467);
or U21538 (N_21538,N_21190,N_21007);
nor U21539 (N_21539,N_21495,N_21350);
xnor U21540 (N_21540,N_21085,N_21251);
nand U21541 (N_21541,N_21005,N_21231);
or U21542 (N_21542,N_21382,N_21452);
nor U21543 (N_21543,N_21225,N_21132);
nand U21544 (N_21544,N_21333,N_21480);
or U21545 (N_21545,N_21080,N_21326);
or U21546 (N_21546,N_21314,N_21494);
or U21547 (N_21547,N_21363,N_21207);
xor U21548 (N_21548,N_21277,N_21043);
and U21549 (N_21549,N_21392,N_21279);
xor U21550 (N_21550,N_21174,N_21205);
and U21551 (N_21551,N_21236,N_21413);
or U21552 (N_21552,N_21464,N_21457);
nand U21553 (N_21553,N_21179,N_21004);
nand U21554 (N_21554,N_21250,N_21224);
or U21555 (N_21555,N_21303,N_21126);
xnor U21556 (N_21556,N_21112,N_21199);
nor U21557 (N_21557,N_21354,N_21163);
nor U21558 (N_21558,N_21156,N_21447);
nor U21559 (N_21559,N_21169,N_21358);
nor U21560 (N_21560,N_21441,N_21439);
nor U21561 (N_21561,N_21337,N_21407);
xor U21562 (N_21562,N_21269,N_21244);
nor U21563 (N_21563,N_21230,N_21037);
nand U21564 (N_21564,N_21355,N_21381);
or U21565 (N_21565,N_21259,N_21400);
and U21566 (N_21566,N_21264,N_21111);
nor U21567 (N_21567,N_21149,N_21054);
or U21568 (N_21568,N_21293,N_21036);
or U21569 (N_21569,N_21496,N_21182);
nand U21570 (N_21570,N_21278,N_21411);
nand U21571 (N_21571,N_21151,N_21021);
and U21572 (N_21572,N_21288,N_21176);
and U21573 (N_21573,N_21150,N_21484);
and U21574 (N_21574,N_21472,N_21081);
xnor U21575 (N_21575,N_21152,N_21370);
or U21576 (N_21576,N_21443,N_21489);
and U21577 (N_21577,N_21458,N_21148);
and U21578 (N_21578,N_21161,N_21171);
xnor U21579 (N_21579,N_21362,N_21016);
nor U21580 (N_21580,N_21361,N_21373);
or U21581 (N_21581,N_21094,N_21393);
nor U21582 (N_21582,N_21087,N_21334);
or U21583 (N_21583,N_21220,N_21282);
nand U21584 (N_21584,N_21419,N_21258);
xnor U21585 (N_21585,N_21451,N_21316);
and U21586 (N_21586,N_21069,N_21218);
xnor U21587 (N_21587,N_21385,N_21383);
and U21588 (N_21588,N_21165,N_21240);
and U21589 (N_21589,N_21051,N_21185);
and U21590 (N_21590,N_21047,N_21033);
nand U21591 (N_21591,N_21092,N_21146);
nor U21592 (N_21592,N_21188,N_21245);
xor U21593 (N_21593,N_21082,N_21045);
and U21594 (N_21594,N_21247,N_21469);
nor U21595 (N_21595,N_21424,N_21408);
and U21596 (N_21596,N_21234,N_21125);
or U21597 (N_21597,N_21202,N_21488);
nor U21598 (N_21598,N_21093,N_21390);
or U21599 (N_21599,N_21341,N_21100);
xor U21600 (N_21600,N_21108,N_21461);
xnor U21601 (N_21601,N_21306,N_21135);
nand U21602 (N_21602,N_21086,N_21088);
and U21603 (N_21603,N_21222,N_21011);
and U21604 (N_21604,N_21030,N_21020);
nor U21605 (N_21605,N_21075,N_21039);
and U21606 (N_21606,N_21432,N_21137);
nor U21607 (N_21607,N_21375,N_21008);
xnor U21608 (N_21608,N_21249,N_21260);
or U21609 (N_21609,N_21487,N_21287);
nand U21610 (N_21610,N_21440,N_21063);
xnor U21611 (N_21611,N_21213,N_21421);
or U21612 (N_21612,N_21367,N_21000);
xor U21613 (N_21613,N_21486,N_21103);
or U21614 (N_21614,N_21083,N_21128);
or U21615 (N_21615,N_21226,N_21299);
and U21616 (N_21616,N_21241,N_21317);
nor U21617 (N_21617,N_21435,N_21117);
or U21618 (N_21618,N_21359,N_21064);
and U21619 (N_21619,N_21027,N_21062);
or U21620 (N_21620,N_21294,N_21490);
nor U21621 (N_21621,N_21232,N_21153);
or U21622 (N_21622,N_21398,N_21498);
nand U21623 (N_21623,N_21107,N_21168);
nand U21624 (N_21624,N_21365,N_21187);
or U21625 (N_21625,N_21397,N_21389);
xor U21626 (N_21626,N_21041,N_21405);
and U21627 (N_21627,N_21013,N_21023);
and U21628 (N_21628,N_21022,N_21209);
nor U21629 (N_21629,N_21297,N_21347);
nand U21630 (N_21630,N_21052,N_21360);
nand U21631 (N_21631,N_21348,N_21173);
nor U21632 (N_21632,N_21172,N_21159);
and U21633 (N_21633,N_21154,N_21380);
nand U21634 (N_21634,N_21235,N_21164);
or U21635 (N_21635,N_21263,N_21034);
or U21636 (N_21636,N_21448,N_21442);
or U21637 (N_21637,N_21136,N_21357);
nor U21638 (N_21638,N_21223,N_21428);
nand U21639 (N_21639,N_21215,N_21426);
and U21640 (N_21640,N_21332,N_21410);
or U21641 (N_21641,N_21318,N_21242);
or U21642 (N_21642,N_21338,N_21449);
nand U21643 (N_21643,N_21002,N_21065);
xor U21644 (N_21644,N_21044,N_21210);
or U21645 (N_21645,N_21074,N_21342);
nand U21646 (N_21646,N_21131,N_21122);
nand U21647 (N_21647,N_21248,N_21305);
nor U21648 (N_21648,N_21284,N_21252);
or U21649 (N_21649,N_21024,N_21456);
nor U21650 (N_21650,N_21366,N_21473);
or U21651 (N_21651,N_21418,N_21123);
nor U21652 (N_21652,N_21257,N_21143);
xnor U21653 (N_21653,N_21404,N_21056);
or U21654 (N_21654,N_21483,N_21216);
or U21655 (N_21655,N_21379,N_21208);
and U21656 (N_21656,N_21059,N_21139);
or U21657 (N_21657,N_21267,N_21296);
xor U21658 (N_21658,N_21095,N_21289);
nor U21659 (N_21659,N_21323,N_21431);
and U21660 (N_21660,N_21420,N_21376);
nor U21661 (N_21661,N_21386,N_21097);
and U21662 (N_21662,N_21127,N_21395);
xor U21663 (N_21663,N_21301,N_21221);
and U21664 (N_21664,N_21372,N_21312);
nand U21665 (N_21665,N_21304,N_21327);
nor U21666 (N_21666,N_21203,N_21072);
or U21667 (N_21667,N_21071,N_21096);
nand U21668 (N_21668,N_21499,N_21349);
xor U21669 (N_21669,N_21181,N_21466);
nor U21670 (N_21670,N_21437,N_21396);
nand U21671 (N_21671,N_21476,N_21118);
xnor U21672 (N_21672,N_21391,N_21116);
nand U21673 (N_21673,N_21227,N_21157);
or U21674 (N_21674,N_21319,N_21254);
xor U21675 (N_21675,N_21091,N_21295);
and U21676 (N_21676,N_21070,N_21214);
nor U21677 (N_21677,N_21378,N_21084);
or U21678 (N_21678,N_21481,N_21353);
and U21679 (N_21679,N_21290,N_21462);
nand U21680 (N_21680,N_21089,N_21031);
nor U21681 (N_21681,N_21058,N_21492);
nor U21682 (N_21682,N_21478,N_21399);
nor U21683 (N_21683,N_21276,N_21160);
and U21684 (N_21684,N_21204,N_21018);
or U21685 (N_21685,N_21253,N_21417);
or U21686 (N_21686,N_21155,N_21465);
nor U21687 (N_21687,N_21015,N_21477);
or U21688 (N_21688,N_21106,N_21336);
nor U21689 (N_21689,N_21340,N_21028);
xnor U21690 (N_21690,N_21292,N_21335);
or U21691 (N_21691,N_21344,N_21402);
nor U21692 (N_21692,N_21434,N_21219);
or U21693 (N_21693,N_21415,N_21029);
or U21694 (N_21694,N_21170,N_21266);
nand U21695 (N_21695,N_21019,N_21105);
or U21696 (N_21696,N_21364,N_21140);
and U21697 (N_21697,N_21130,N_21270);
xor U21698 (N_21698,N_21026,N_21014);
xor U21699 (N_21699,N_21425,N_21369);
nand U21700 (N_21700,N_21302,N_21200);
and U21701 (N_21701,N_21142,N_21133);
and U21702 (N_21702,N_21273,N_21177);
xnor U21703 (N_21703,N_21206,N_21121);
nor U21704 (N_21704,N_21300,N_21394);
and U21705 (N_21705,N_21265,N_21321);
xnor U21706 (N_21706,N_21129,N_21053);
nand U21707 (N_21707,N_21010,N_21388);
nand U21708 (N_21708,N_21406,N_21414);
nand U21709 (N_21709,N_21066,N_21272);
or U21710 (N_21710,N_21119,N_21493);
xnor U21711 (N_21711,N_21459,N_21201);
xor U21712 (N_21712,N_21167,N_21090);
xnor U21713 (N_21713,N_21356,N_21040);
or U21714 (N_21714,N_21068,N_21197);
xnor U21715 (N_21715,N_21124,N_21352);
xor U21716 (N_21716,N_21485,N_21497);
or U21717 (N_21717,N_21471,N_21189);
nor U21718 (N_21718,N_21271,N_21061);
nor U21719 (N_21719,N_21055,N_21281);
and U21720 (N_21720,N_21060,N_21238);
nor U21721 (N_21721,N_21374,N_21003);
or U21722 (N_21722,N_21450,N_21455);
or U21723 (N_21723,N_21192,N_21343);
nor U21724 (N_21724,N_21401,N_21325);
nor U21725 (N_21725,N_21048,N_21275);
and U21726 (N_21726,N_21104,N_21475);
nor U21727 (N_21727,N_21101,N_21430);
xnor U21728 (N_21728,N_21098,N_21042);
nor U21729 (N_21729,N_21144,N_21387);
or U21730 (N_21730,N_21198,N_21178);
nor U21731 (N_21731,N_21346,N_21195);
xnor U21732 (N_21732,N_21482,N_21239);
nor U21733 (N_21733,N_21141,N_21468);
nand U21734 (N_21734,N_21255,N_21261);
xnor U21735 (N_21735,N_21427,N_21025);
or U21736 (N_21736,N_21268,N_21050);
or U21737 (N_21737,N_21423,N_21006);
and U21738 (N_21738,N_21285,N_21328);
nand U21739 (N_21739,N_21166,N_21377);
nand U21740 (N_21740,N_21217,N_21324);
or U21741 (N_21741,N_21184,N_21193);
and U21742 (N_21742,N_21460,N_21243);
and U21743 (N_21743,N_21329,N_21246);
nor U21744 (N_21744,N_21412,N_21474);
or U21745 (N_21745,N_21017,N_21012);
nand U21746 (N_21746,N_21186,N_21286);
and U21747 (N_21747,N_21446,N_21076);
nand U21748 (N_21748,N_21416,N_21274);
and U21749 (N_21749,N_21180,N_21229);
and U21750 (N_21750,N_21042,N_21308);
nand U21751 (N_21751,N_21038,N_21365);
or U21752 (N_21752,N_21113,N_21191);
and U21753 (N_21753,N_21347,N_21358);
and U21754 (N_21754,N_21465,N_21373);
nand U21755 (N_21755,N_21220,N_21319);
and U21756 (N_21756,N_21250,N_21371);
xor U21757 (N_21757,N_21325,N_21248);
xnor U21758 (N_21758,N_21362,N_21381);
or U21759 (N_21759,N_21350,N_21311);
or U21760 (N_21760,N_21155,N_21489);
or U21761 (N_21761,N_21447,N_21499);
or U21762 (N_21762,N_21030,N_21034);
or U21763 (N_21763,N_21319,N_21024);
nand U21764 (N_21764,N_21062,N_21131);
and U21765 (N_21765,N_21407,N_21101);
nor U21766 (N_21766,N_21115,N_21351);
xor U21767 (N_21767,N_21317,N_21214);
nand U21768 (N_21768,N_21032,N_21184);
nand U21769 (N_21769,N_21006,N_21278);
nor U21770 (N_21770,N_21370,N_21057);
or U21771 (N_21771,N_21126,N_21187);
xnor U21772 (N_21772,N_21440,N_21098);
nor U21773 (N_21773,N_21059,N_21117);
xnor U21774 (N_21774,N_21361,N_21068);
or U21775 (N_21775,N_21396,N_21237);
xnor U21776 (N_21776,N_21223,N_21343);
nand U21777 (N_21777,N_21117,N_21086);
or U21778 (N_21778,N_21336,N_21378);
xnor U21779 (N_21779,N_21137,N_21362);
or U21780 (N_21780,N_21001,N_21331);
and U21781 (N_21781,N_21100,N_21489);
nor U21782 (N_21782,N_21152,N_21479);
nor U21783 (N_21783,N_21146,N_21493);
xnor U21784 (N_21784,N_21134,N_21476);
and U21785 (N_21785,N_21077,N_21273);
nand U21786 (N_21786,N_21211,N_21198);
nand U21787 (N_21787,N_21233,N_21238);
and U21788 (N_21788,N_21407,N_21041);
and U21789 (N_21789,N_21088,N_21074);
and U21790 (N_21790,N_21039,N_21004);
and U21791 (N_21791,N_21266,N_21113);
nand U21792 (N_21792,N_21275,N_21104);
nor U21793 (N_21793,N_21104,N_21448);
and U21794 (N_21794,N_21038,N_21339);
nor U21795 (N_21795,N_21295,N_21112);
xor U21796 (N_21796,N_21248,N_21491);
or U21797 (N_21797,N_21465,N_21486);
nand U21798 (N_21798,N_21256,N_21106);
or U21799 (N_21799,N_21132,N_21209);
nand U21800 (N_21800,N_21285,N_21082);
and U21801 (N_21801,N_21241,N_21024);
and U21802 (N_21802,N_21492,N_21255);
nand U21803 (N_21803,N_21346,N_21117);
or U21804 (N_21804,N_21340,N_21003);
nor U21805 (N_21805,N_21426,N_21411);
and U21806 (N_21806,N_21440,N_21361);
nor U21807 (N_21807,N_21292,N_21052);
xor U21808 (N_21808,N_21346,N_21499);
nor U21809 (N_21809,N_21476,N_21015);
or U21810 (N_21810,N_21239,N_21135);
nor U21811 (N_21811,N_21169,N_21032);
xor U21812 (N_21812,N_21021,N_21121);
and U21813 (N_21813,N_21280,N_21158);
nand U21814 (N_21814,N_21119,N_21059);
nor U21815 (N_21815,N_21180,N_21477);
nand U21816 (N_21816,N_21022,N_21117);
and U21817 (N_21817,N_21187,N_21299);
nand U21818 (N_21818,N_21383,N_21086);
and U21819 (N_21819,N_21175,N_21364);
and U21820 (N_21820,N_21336,N_21304);
or U21821 (N_21821,N_21238,N_21176);
nand U21822 (N_21822,N_21271,N_21284);
and U21823 (N_21823,N_21446,N_21381);
xnor U21824 (N_21824,N_21004,N_21458);
xnor U21825 (N_21825,N_21010,N_21048);
xnor U21826 (N_21826,N_21054,N_21218);
or U21827 (N_21827,N_21490,N_21406);
and U21828 (N_21828,N_21192,N_21302);
nand U21829 (N_21829,N_21388,N_21018);
nand U21830 (N_21830,N_21253,N_21412);
or U21831 (N_21831,N_21369,N_21066);
nand U21832 (N_21832,N_21159,N_21238);
nor U21833 (N_21833,N_21225,N_21054);
xnor U21834 (N_21834,N_21034,N_21246);
and U21835 (N_21835,N_21214,N_21450);
and U21836 (N_21836,N_21379,N_21039);
nor U21837 (N_21837,N_21068,N_21329);
nor U21838 (N_21838,N_21022,N_21448);
xor U21839 (N_21839,N_21129,N_21303);
nor U21840 (N_21840,N_21288,N_21231);
nand U21841 (N_21841,N_21133,N_21442);
and U21842 (N_21842,N_21375,N_21322);
xor U21843 (N_21843,N_21324,N_21248);
xor U21844 (N_21844,N_21068,N_21117);
or U21845 (N_21845,N_21121,N_21139);
or U21846 (N_21846,N_21290,N_21357);
and U21847 (N_21847,N_21368,N_21061);
xnor U21848 (N_21848,N_21340,N_21447);
or U21849 (N_21849,N_21456,N_21312);
nor U21850 (N_21850,N_21377,N_21188);
and U21851 (N_21851,N_21286,N_21188);
nand U21852 (N_21852,N_21272,N_21096);
xnor U21853 (N_21853,N_21152,N_21209);
and U21854 (N_21854,N_21195,N_21338);
nor U21855 (N_21855,N_21196,N_21465);
xnor U21856 (N_21856,N_21405,N_21310);
nor U21857 (N_21857,N_21128,N_21136);
xor U21858 (N_21858,N_21152,N_21391);
xnor U21859 (N_21859,N_21307,N_21020);
or U21860 (N_21860,N_21263,N_21321);
nor U21861 (N_21861,N_21456,N_21056);
nand U21862 (N_21862,N_21428,N_21463);
nor U21863 (N_21863,N_21203,N_21415);
nand U21864 (N_21864,N_21388,N_21355);
and U21865 (N_21865,N_21118,N_21479);
nor U21866 (N_21866,N_21199,N_21157);
nor U21867 (N_21867,N_21011,N_21284);
nor U21868 (N_21868,N_21062,N_21372);
nand U21869 (N_21869,N_21362,N_21206);
or U21870 (N_21870,N_21239,N_21117);
xor U21871 (N_21871,N_21167,N_21408);
nor U21872 (N_21872,N_21435,N_21240);
nor U21873 (N_21873,N_21008,N_21199);
or U21874 (N_21874,N_21464,N_21492);
nand U21875 (N_21875,N_21302,N_21442);
nor U21876 (N_21876,N_21052,N_21096);
or U21877 (N_21877,N_21123,N_21370);
or U21878 (N_21878,N_21113,N_21350);
or U21879 (N_21879,N_21308,N_21214);
nor U21880 (N_21880,N_21122,N_21348);
nor U21881 (N_21881,N_21453,N_21428);
or U21882 (N_21882,N_21266,N_21222);
nor U21883 (N_21883,N_21447,N_21084);
nor U21884 (N_21884,N_21233,N_21289);
nand U21885 (N_21885,N_21320,N_21375);
nor U21886 (N_21886,N_21080,N_21316);
xnor U21887 (N_21887,N_21342,N_21235);
and U21888 (N_21888,N_21032,N_21066);
nand U21889 (N_21889,N_21244,N_21043);
nand U21890 (N_21890,N_21182,N_21163);
nor U21891 (N_21891,N_21224,N_21356);
or U21892 (N_21892,N_21174,N_21181);
or U21893 (N_21893,N_21073,N_21354);
xnor U21894 (N_21894,N_21341,N_21384);
or U21895 (N_21895,N_21215,N_21031);
nand U21896 (N_21896,N_21119,N_21270);
xnor U21897 (N_21897,N_21213,N_21368);
and U21898 (N_21898,N_21432,N_21402);
xnor U21899 (N_21899,N_21376,N_21499);
nand U21900 (N_21900,N_21190,N_21082);
nor U21901 (N_21901,N_21194,N_21069);
and U21902 (N_21902,N_21170,N_21383);
nor U21903 (N_21903,N_21171,N_21298);
nor U21904 (N_21904,N_21221,N_21447);
and U21905 (N_21905,N_21103,N_21225);
nand U21906 (N_21906,N_21363,N_21495);
or U21907 (N_21907,N_21050,N_21212);
or U21908 (N_21908,N_21048,N_21425);
xnor U21909 (N_21909,N_21200,N_21484);
nor U21910 (N_21910,N_21211,N_21319);
nor U21911 (N_21911,N_21409,N_21323);
xor U21912 (N_21912,N_21490,N_21139);
or U21913 (N_21913,N_21126,N_21038);
nand U21914 (N_21914,N_21403,N_21454);
xor U21915 (N_21915,N_21139,N_21164);
nand U21916 (N_21916,N_21205,N_21457);
or U21917 (N_21917,N_21205,N_21172);
or U21918 (N_21918,N_21173,N_21278);
xnor U21919 (N_21919,N_21010,N_21235);
nand U21920 (N_21920,N_21142,N_21018);
xnor U21921 (N_21921,N_21010,N_21233);
nor U21922 (N_21922,N_21216,N_21172);
and U21923 (N_21923,N_21116,N_21152);
nor U21924 (N_21924,N_21401,N_21209);
xor U21925 (N_21925,N_21107,N_21363);
nand U21926 (N_21926,N_21219,N_21230);
xnor U21927 (N_21927,N_21388,N_21228);
or U21928 (N_21928,N_21174,N_21260);
or U21929 (N_21929,N_21325,N_21439);
nor U21930 (N_21930,N_21438,N_21456);
xor U21931 (N_21931,N_21018,N_21331);
or U21932 (N_21932,N_21141,N_21333);
or U21933 (N_21933,N_21156,N_21390);
and U21934 (N_21934,N_21148,N_21238);
xor U21935 (N_21935,N_21104,N_21250);
and U21936 (N_21936,N_21388,N_21350);
nor U21937 (N_21937,N_21382,N_21340);
or U21938 (N_21938,N_21127,N_21456);
and U21939 (N_21939,N_21021,N_21485);
and U21940 (N_21940,N_21131,N_21145);
xor U21941 (N_21941,N_21319,N_21156);
or U21942 (N_21942,N_21245,N_21480);
nand U21943 (N_21943,N_21116,N_21144);
and U21944 (N_21944,N_21491,N_21416);
or U21945 (N_21945,N_21107,N_21120);
and U21946 (N_21946,N_21313,N_21495);
xnor U21947 (N_21947,N_21449,N_21015);
or U21948 (N_21948,N_21447,N_21266);
xor U21949 (N_21949,N_21068,N_21398);
xnor U21950 (N_21950,N_21235,N_21403);
and U21951 (N_21951,N_21308,N_21488);
or U21952 (N_21952,N_21092,N_21238);
or U21953 (N_21953,N_21217,N_21446);
xnor U21954 (N_21954,N_21114,N_21318);
nor U21955 (N_21955,N_21166,N_21451);
and U21956 (N_21956,N_21327,N_21068);
nor U21957 (N_21957,N_21281,N_21157);
or U21958 (N_21958,N_21187,N_21439);
or U21959 (N_21959,N_21070,N_21192);
xnor U21960 (N_21960,N_21143,N_21085);
nor U21961 (N_21961,N_21170,N_21004);
and U21962 (N_21962,N_21419,N_21451);
nor U21963 (N_21963,N_21217,N_21058);
nand U21964 (N_21964,N_21352,N_21101);
nand U21965 (N_21965,N_21233,N_21229);
xor U21966 (N_21966,N_21323,N_21359);
xnor U21967 (N_21967,N_21096,N_21464);
xnor U21968 (N_21968,N_21327,N_21064);
and U21969 (N_21969,N_21097,N_21469);
or U21970 (N_21970,N_21197,N_21374);
nor U21971 (N_21971,N_21038,N_21370);
nor U21972 (N_21972,N_21447,N_21159);
and U21973 (N_21973,N_21307,N_21200);
and U21974 (N_21974,N_21383,N_21303);
nand U21975 (N_21975,N_21261,N_21336);
nor U21976 (N_21976,N_21191,N_21353);
nand U21977 (N_21977,N_21026,N_21263);
nand U21978 (N_21978,N_21063,N_21001);
nor U21979 (N_21979,N_21185,N_21093);
or U21980 (N_21980,N_21141,N_21354);
nor U21981 (N_21981,N_21489,N_21107);
nor U21982 (N_21982,N_21141,N_21083);
nor U21983 (N_21983,N_21202,N_21334);
or U21984 (N_21984,N_21170,N_21087);
or U21985 (N_21985,N_21220,N_21134);
xor U21986 (N_21986,N_21246,N_21224);
nand U21987 (N_21987,N_21414,N_21139);
or U21988 (N_21988,N_21042,N_21279);
xor U21989 (N_21989,N_21173,N_21228);
or U21990 (N_21990,N_21376,N_21032);
xor U21991 (N_21991,N_21378,N_21409);
or U21992 (N_21992,N_21179,N_21409);
nand U21993 (N_21993,N_21146,N_21079);
xnor U21994 (N_21994,N_21257,N_21324);
or U21995 (N_21995,N_21413,N_21162);
nand U21996 (N_21996,N_21048,N_21368);
xnor U21997 (N_21997,N_21467,N_21190);
xor U21998 (N_21998,N_21164,N_21135);
and U21999 (N_21999,N_21473,N_21377);
or U22000 (N_22000,N_21942,N_21936);
xnor U22001 (N_22001,N_21726,N_21877);
xnor U22002 (N_22002,N_21864,N_21829);
or U22003 (N_22003,N_21506,N_21976);
and U22004 (N_22004,N_21690,N_21838);
and U22005 (N_22005,N_21850,N_21841);
xor U22006 (N_22006,N_21657,N_21804);
nor U22007 (N_22007,N_21627,N_21696);
nand U22008 (N_22008,N_21884,N_21786);
nand U22009 (N_22009,N_21733,N_21730);
nand U22010 (N_22010,N_21950,N_21963);
and U22011 (N_22011,N_21734,N_21554);
or U22012 (N_22012,N_21934,N_21571);
xnor U22013 (N_22013,N_21663,N_21562);
nand U22014 (N_22014,N_21636,N_21565);
nor U22015 (N_22015,N_21731,N_21603);
or U22016 (N_22016,N_21748,N_21525);
nand U22017 (N_22017,N_21972,N_21984);
or U22018 (N_22018,N_21755,N_21533);
xor U22019 (N_22019,N_21694,N_21975);
nand U22020 (N_22020,N_21827,N_21656);
xor U22021 (N_22021,N_21575,N_21511);
and U22022 (N_22022,N_21995,N_21505);
nand U22023 (N_22023,N_21589,N_21534);
nand U22024 (N_22024,N_21668,N_21591);
or U22025 (N_22025,N_21746,N_21914);
or U22026 (N_22026,N_21553,N_21658);
xor U22027 (N_22027,N_21951,N_21903);
or U22028 (N_22028,N_21969,N_21962);
nand U22029 (N_22029,N_21773,N_21530);
or U22030 (N_22030,N_21618,N_21714);
xor U22031 (N_22031,N_21614,N_21518);
xor U22032 (N_22032,N_21549,N_21593);
nand U22033 (N_22033,N_21599,N_21788);
or U22034 (N_22034,N_21856,N_21871);
and U22035 (N_22035,N_21558,N_21686);
and U22036 (N_22036,N_21974,N_21598);
nand U22037 (N_22037,N_21846,N_21892);
nor U22038 (N_22038,N_21996,N_21768);
nand U22039 (N_22039,N_21601,N_21781);
nand U22040 (N_22040,N_21832,N_21767);
nor U22041 (N_22041,N_21954,N_21917);
nor U22042 (N_22042,N_21783,N_21808);
xor U22043 (N_22043,N_21967,N_21957);
nand U22044 (N_22044,N_21873,N_21607);
and U22045 (N_22045,N_21921,N_21784);
nor U22046 (N_22046,N_21899,N_21585);
and U22047 (N_22047,N_21582,N_21735);
and U22048 (N_22048,N_21878,N_21512);
nor U22049 (N_22049,N_21741,N_21654);
nand U22050 (N_22050,N_21681,N_21888);
or U22051 (N_22051,N_21674,N_21897);
xor U22052 (N_22052,N_21502,N_21790);
nor U22053 (N_22053,N_21749,N_21789);
nand U22054 (N_22054,N_21820,N_21826);
xnor U22055 (N_22055,N_21772,N_21794);
xor U22056 (N_22056,N_21799,N_21955);
or U22057 (N_22057,N_21870,N_21641);
xnor U22058 (N_22058,N_21766,N_21707);
and U22059 (N_22059,N_21573,N_21724);
nor U22060 (N_22060,N_21561,N_21697);
and U22061 (N_22061,N_21504,N_21959);
xor U22062 (N_22062,N_21557,N_21776);
or U22063 (N_22063,N_21718,N_21981);
or U22064 (N_22064,N_21610,N_21979);
nand U22065 (N_22065,N_21866,N_21853);
and U22066 (N_22066,N_21949,N_21765);
xor U22067 (N_22067,N_21947,N_21705);
xor U22068 (N_22068,N_21624,N_21664);
nor U22069 (N_22069,N_21721,N_21572);
nand U22070 (N_22070,N_21855,N_21513);
nand U22071 (N_22071,N_21762,N_21539);
and U22072 (N_22072,N_21991,N_21544);
nand U22073 (N_22073,N_21545,N_21527);
xor U22074 (N_22074,N_21980,N_21854);
nand U22075 (N_22075,N_21528,N_21987);
or U22076 (N_22076,N_21824,N_21524);
xnor U22077 (N_22077,N_21823,N_21570);
xnor U22078 (N_22078,N_21851,N_21898);
nor U22079 (N_22079,N_21739,N_21901);
and U22080 (N_22080,N_21716,N_21612);
or U22081 (N_22081,N_21879,N_21999);
nand U22082 (N_22082,N_21862,N_21815);
or U22083 (N_22083,N_21740,N_21777);
nor U22084 (N_22084,N_21619,N_21874);
nand U22085 (N_22085,N_21736,N_21583);
nand U22086 (N_22086,N_21863,N_21905);
nor U22087 (N_22087,N_21831,N_21509);
xor U22088 (N_22088,N_21578,N_21514);
nor U22089 (N_22089,N_21693,N_21632);
nand U22090 (N_22090,N_21737,N_21821);
and U22091 (N_22091,N_21523,N_21596);
nand U22092 (N_22092,N_21983,N_21977);
nand U22093 (N_22093,N_21791,N_21522);
nand U22094 (N_22094,N_21937,N_21617);
nand U22095 (N_22095,N_21630,N_21688);
nor U22096 (N_22096,N_21782,N_21673);
or U22097 (N_22097,N_21728,N_21845);
and U22098 (N_22098,N_21960,N_21639);
and U22099 (N_22099,N_21973,N_21891);
xor U22100 (N_22100,N_21802,N_21894);
nor U22101 (N_22101,N_21683,N_21715);
xor U22102 (N_22102,N_21590,N_21811);
nor U22103 (N_22103,N_21629,N_21952);
and U22104 (N_22104,N_21876,N_21515);
nand U22105 (N_22105,N_21633,N_21990);
nor U22106 (N_22106,N_21985,N_21836);
xor U22107 (N_22107,N_21550,N_21819);
or U22108 (N_22108,N_21989,N_21925);
or U22109 (N_22109,N_21887,N_21586);
and U22110 (N_22110,N_21764,N_21594);
xnor U22111 (N_22111,N_21889,N_21930);
or U22112 (N_22112,N_21946,N_21813);
xor U22113 (N_22113,N_21993,N_21920);
xor U22114 (N_22114,N_21595,N_21812);
nor U22115 (N_22115,N_21556,N_21638);
nor U22116 (N_22116,N_21725,N_21971);
nand U22117 (N_22117,N_21912,N_21760);
xnor U22118 (N_22118,N_21919,N_21939);
or U22119 (N_22119,N_21780,N_21759);
nor U22120 (N_22120,N_21587,N_21576);
xnor U22121 (N_22121,N_21692,N_21647);
xor U22122 (N_22122,N_21729,N_21631);
xnor U22123 (N_22123,N_21757,N_21907);
nor U22124 (N_22124,N_21703,N_21625);
nor U22125 (N_22125,N_21893,N_21540);
xor U22126 (N_22126,N_21531,N_21835);
or U22127 (N_22127,N_21613,N_21935);
and U22128 (N_22128,N_21822,N_21800);
nor U22129 (N_22129,N_21564,N_21908);
and U22130 (N_22130,N_21538,N_21666);
or U22131 (N_22131,N_21532,N_21526);
and U22132 (N_22132,N_21861,N_21992);
and U22133 (N_22133,N_21801,N_21727);
nand U22134 (N_22134,N_21695,N_21805);
nand U22135 (N_22135,N_21940,N_21560);
nor U22136 (N_22136,N_21543,N_21843);
nand U22137 (N_22137,N_21691,N_21645);
nand U22138 (N_22138,N_21644,N_21994);
nor U22139 (N_22139,N_21883,N_21916);
or U22140 (N_22140,N_21604,N_21609);
xor U22141 (N_22141,N_21902,N_21988);
nor U22142 (N_22142,N_21709,N_21941);
nor U22143 (N_22143,N_21672,N_21833);
xor U22144 (N_22144,N_21675,N_21659);
xnor U22145 (N_22145,N_21652,N_21551);
nand U22146 (N_22146,N_21842,N_21915);
or U22147 (N_22147,N_21685,N_21653);
nand U22148 (N_22148,N_21763,N_21886);
or U22149 (N_22149,N_21529,N_21643);
and U22150 (N_22150,N_21507,N_21677);
nand U22151 (N_22151,N_21535,N_21931);
and U22152 (N_22152,N_21592,N_21742);
nand U22153 (N_22153,N_21814,N_21660);
or U22154 (N_22154,N_21706,N_21542);
and U22155 (N_22155,N_21932,N_21684);
and U22156 (N_22156,N_21698,N_21834);
nor U22157 (N_22157,N_21754,N_21517);
and U22158 (N_22158,N_21758,N_21968);
nand U22159 (N_22159,N_21769,N_21849);
or U22160 (N_22160,N_21860,N_21546);
and U22161 (N_22161,N_21597,N_21918);
nor U22162 (N_22162,N_21508,N_21548);
and U22163 (N_22163,N_21655,N_21837);
or U22164 (N_22164,N_21559,N_21982);
nand U22165 (N_22165,N_21678,N_21661);
xnor U22166 (N_22166,N_21669,N_21671);
and U22167 (N_22167,N_21970,N_21956);
and U22168 (N_22168,N_21779,N_21965);
xor U22169 (N_22169,N_21615,N_21605);
nor U22170 (N_22170,N_21648,N_21938);
or U22171 (N_22171,N_21825,N_21787);
xnor U22172 (N_22172,N_21785,N_21708);
nand U22173 (N_22173,N_21521,N_21600);
xor U22174 (N_22174,N_21806,N_21699);
or U22175 (N_22175,N_21964,N_21828);
nand U22176 (N_22176,N_21774,N_21750);
nor U22177 (N_22177,N_21756,N_21717);
xor U22178 (N_22178,N_21722,N_21662);
or U22179 (N_22179,N_21606,N_21701);
xor U22180 (N_22180,N_21602,N_21563);
and U22181 (N_22181,N_21574,N_21998);
nor U22182 (N_22182,N_21628,N_21650);
and U22183 (N_22183,N_21541,N_21751);
or U22184 (N_22184,N_21651,N_21953);
nor U22185 (N_22185,N_21679,N_21616);
xnor U22186 (N_22186,N_21667,N_21961);
nand U22187 (N_22187,N_21611,N_21830);
and U22188 (N_22188,N_21520,N_21798);
and U22189 (N_22189,N_21637,N_21880);
xor U22190 (N_22190,N_21711,N_21913);
xnor U22191 (N_22191,N_21922,N_21682);
xor U22192 (N_22192,N_21933,N_21702);
xnor U22193 (N_22193,N_21700,N_21796);
or U22194 (N_22194,N_21710,N_21986);
nand U22195 (N_22195,N_21713,N_21537);
or U22196 (N_22196,N_21552,N_21577);
nor U22197 (N_22197,N_21809,N_21844);
nor U22198 (N_22198,N_21569,N_21890);
and U22199 (N_22199,N_21906,N_21875);
xor U22200 (N_22200,N_21536,N_21581);
and U22201 (N_22201,N_21797,N_21665);
and U22202 (N_22202,N_21712,N_21882);
nor U22203 (N_22203,N_21580,N_21719);
nand U22204 (N_22204,N_21817,N_21928);
nor U22205 (N_22205,N_21752,N_21634);
or U22206 (N_22206,N_21622,N_21670);
and U22207 (N_22207,N_21895,N_21778);
and U22208 (N_22208,N_21885,N_21929);
nor U22209 (N_22209,N_21868,N_21566);
nand U22210 (N_22210,N_21608,N_21948);
or U22211 (N_22211,N_21859,N_21810);
nand U22212 (N_22212,N_21881,N_21567);
and U22213 (N_22213,N_21770,N_21500);
or U22214 (N_22214,N_21753,N_21519);
xnor U22215 (N_22215,N_21904,N_21649);
or U22216 (N_22216,N_21943,N_21687);
or U22217 (N_22217,N_21503,N_21944);
nand U22218 (N_22218,N_21635,N_21723);
xor U22219 (N_22219,N_21910,N_21588);
or U22220 (N_22220,N_21620,N_21640);
nor U22221 (N_22221,N_21966,N_21626);
nor U22222 (N_22222,N_21848,N_21793);
nor U22223 (N_22223,N_21852,N_21847);
and U22224 (N_22224,N_21858,N_21555);
nand U22225 (N_22225,N_21568,N_21869);
xnor U22226 (N_22226,N_21775,N_21872);
and U22227 (N_22227,N_21926,N_21761);
and U22228 (N_22228,N_21732,N_21676);
nor U22229 (N_22229,N_21501,N_21911);
nor U22230 (N_22230,N_21803,N_21909);
and U22231 (N_22231,N_21704,N_21857);
and U22232 (N_22232,N_21900,N_21744);
nand U22233 (N_22233,N_21720,N_21816);
and U22234 (N_22234,N_21865,N_21689);
nor U22235 (N_22235,N_21945,N_21923);
nand U22236 (N_22236,N_21747,N_21896);
or U22237 (N_22237,N_21579,N_21745);
xnor U22238 (N_22238,N_21839,N_21792);
nand U22239 (N_22239,N_21738,N_21958);
nand U22240 (N_22240,N_21927,N_21997);
nor U22241 (N_22241,N_21818,N_21924);
or U22242 (N_22242,N_21867,N_21840);
xnor U22243 (N_22243,N_21795,N_21584);
nor U22244 (N_22244,N_21646,N_21547);
nand U22245 (N_22245,N_21642,N_21771);
nor U22246 (N_22246,N_21743,N_21680);
nand U22247 (N_22247,N_21623,N_21978);
nand U22248 (N_22248,N_21510,N_21621);
or U22249 (N_22249,N_21807,N_21516);
nor U22250 (N_22250,N_21934,N_21739);
nor U22251 (N_22251,N_21565,N_21906);
xor U22252 (N_22252,N_21922,N_21692);
and U22253 (N_22253,N_21595,N_21530);
nand U22254 (N_22254,N_21577,N_21969);
or U22255 (N_22255,N_21507,N_21514);
nand U22256 (N_22256,N_21807,N_21845);
nor U22257 (N_22257,N_21703,N_21750);
or U22258 (N_22258,N_21731,N_21674);
xor U22259 (N_22259,N_21659,N_21679);
nand U22260 (N_22260,N_21638,N_21787);
xor U22261 (N_22261,N_21973,N_21512);
nand U22262 (N_22262,N_21786,N_21908);
xor U22263 (N_22263,N_21995,N_21651);
nand U22264 (N_22264,N_21619,N_21666);
xor U22265 (N_22265,N_21982,N_21764);
or U22266 (N_22266,N_21807,N_21958);
and U22267 (N_22267,N_21783,N_21962);
xnor U22268 (N_22268,N_21806,N_21702);
nand U22269 (N_22269,N_21914,N_21800);
nor U22270 (N_22270,N_21782,N_21763);
or U22271 (N_22271,N_21857,N_21786);
xnor U22272 (N_22272,N_21731,N_21568);
and U22273 (N_22273,N_21535,N_21884);
nor U22274 (N_22274,N_21639,N_21794);
or U22275 (N_22275,N_21613,N_21906);
and U22276 (N_22276,N_21518,N_21854);
nor U22277 (N_22277,N_21913,N_21690);
or U22278 (N_22278,N_21574,N_21511);
xor U22279 (N_22279,N_21715,N_21826);
and U22280 (N_22280,N_21965,N_21708);
nand U22281 (N_22281,N_21903,N_21627);
nand U22282 (N_22282,N_21621,N_21701);
xor U22283 (N_22283,N_21978,N_21728);
or U22284 (N_22284,N_21929,N_21780);
nor U22285 (N_22285,N_21551,N_21775);
nor U22286 (N_22286,N_21547,N_21795);
xnor U22287 (N_22287,N_21771,N_21999);
or U22288 (N_22288,N_21830,N_21723);
nand U22289 (N_22289,N_21962,N_21699);
nor U22290 (N_22290,N_21593,N_21820);
xnor U22291 (N_22291,N_21826,N_21767);
or U22292 (N_22292,N_21831,N_21847);
or U22293 (N_22293,N_21937,N_21509);
nor U22294 (N_22294,N_21731,N_21996);
or U22295 (N_22295,N_21576,N_21539);
or U22296 (N_22296,N_21565,N_21722);
nand U22297 (N_22297,N_21590,N_21740);
and U22298 (N_22298,N_21715,N_21748);
nor U22299 (N_22299,N_21743,N_21606);
nor U22300 (N_22300,N_21863,N_21883);
nor U22301 (N_22301,N_21747,N_21906);
or U22302 (N_22302,N_21778,N_21696);
xnor U22303 (N_22303,N_21742,N_21902);
nand U22304 (N_22304,N_21856,N_21642);
nand U22305 (N_22305,N_21732,N_21663);
or U22306 (N_22306,N_21906,N_21791);
nand U22307 (N_22307,N_21556,N_21577);
and U22308 (N_22308,N_21587,N_21536);
nor U22309 (N_22309,N_21911,N_21968);
xor U22310 (N_22310,N_21730,N_21989);
nand U22311 (N_22311,N_21773,N_21844);
and U22312 (N_22312,N_21997,N_21923);
or U22313 (N_22313,N_21550,N_21639);
and U22314 (N_22314,N_21785,N_21781);
xnor U22315 (N_22315,N_21726,N_21873);
nand U22316 (N_22316,N_21711,N_21613);
or U22317 (N_22317,N_21575,N_21771);
xor U22318 (N_22318,N_21822,N_21783);
or U22319 (N_22319,N_21664,N_21709);
or U22320 (N_22320,N_21858,N_21590);
xnor U22321 (N_22321,N_21611,N_21537);
nor U22322 (N_22322,N_21950,N_21527);
or U22323 (N_22323,N_21846,N_21894);
nand U22324 (N_22324,N_21658,N_21676);
xnor U22325 (N_22325,N_21908,N_21600);
nor U22326 (N_22326,N_21530,N_21729);
and U22327 (N_22327,N_21841,N_21960);
nor U22328 (N_22328,N_21823,N_21765);
nand U22329 (N_22329,N_21589,N_21807);
and U22330 (N_22330,N_21797,N_21558);
and U22331 (N_22331,N_21853,N_21521);
and U22332 (N_22332,N_21959,N_21727);
or U22333 (N_22333,N_21704,N_21815);
nor U22334 (N_22334,N_21979,N_21662);
and U22335 (N_22335,N_21751,N_21675);
or U22336 (N_22336,N_21827,N_21720);
and U22337 (N_22337,N_21735,N_21574);
nor U22338 (N_22338,N_21845,N_21962);
or U22339 (N_22339,N_21594,N_21746);
nor U22340 (N_22340,N_21751,N_21571);
xnor U22341 (N_22341,N_21604,N_21549);
nor U22342 (N_22342,N_21669,N_21538);
xnor U22343 (N_22343,N_21552,N_21872);
xnor U22344 (N_22344,N_21667,N_21756);
or U22345 (N_22345,N_21948,N_21711);
xnor U22346 (N_22346,N_21811,N_21972);
and U22347 (N_22347,N_21501,N_21684);
nand U22348 (N_22348,N_21658,N_21593);
nand U22349 (N_22349,N_21687,N_21606);
or U22350 (N_22350,N_21713,N_21579);
or U22351 (N_22351,N_21784,N_21794);
nand U22352 (N_22352,N_21709,N_21813);
and U22353 (N_22353,N_21530,N_21682);
and U22354 (N_22354,N_21633,N_21897);
or U22355 (N_22355,N_21836,N_21992);
nor U22356 (N_22356,N_21823,N_21682);
nor U22357 (N_22357,N_21928,N_21607);
and U22358 (N_22358,N_21689,N_21682);
nor U22359 (N_22359,N_21783,N_21634);
nand U22360 (N_22360,N_21676,N_21975);
nand U22361 (N_22361,N_21736,N_21879);
and U22362 (N_22362,N_21777,N_21855);
xor U22363 (N_22363,N_21519,N_21676);
and U22364 (N_22364,N_21779,N_21881);
and U22365 (N_22365,N_21818,N_21795);
xnor U22366 (N_22366,N_21673,N_21691);
nor U22367 (N_22367,N_21504,N_21518);
nor U22368 (N_22368,N_21516,N_21556);
or U22369 (N_22369,N_21526,N_21600);
nand U22370 (N_22370,N_21736,N_21518);
and U22371 (N_22371,N_21577,N_21567);
nor U22372 (N_22372,N_21946,N_21962);
nand U22373 (N_22373,N_21599,N_21521);
xor U22374 (N_22374,N_21834,N_21880);
xnor U22375 (N_22375,N_21583,N_21690);
or U22376 (N_22376,N_21704,N_21625);
or U22377 (N_22377,N_21676,N_21597);
xnor U22378 (N_22378,N_21788,N_21860);
xor U22379 (N_22379,N_21880,N_21789);
nor U22380 (N_22380,N_21552,N_21514);
nand U22381 (N_22381,N_21512,N_21727);
nor U22382 (N_22382,N_21873,N_21736);
and U22383 (N_22383,N_21828,N_21763);
xnor U22384 (N_22384,N_21596,N_21867);
nor U22385 (N_22385,N_21972,N_21679);
nand U22386 (N_22386,N_21981,N_21947);
and U22387 (N_22387,N_21530,N_21665);
or U22388 (N_22388,N_21990,N_21688);
and U22389 (N_22389,N_21501,N_21907);
xnor U22390 (N_22390,N_21597,N_21666);
nor U22391 (N_22391,N_21862,N_21699);
nand U22392 (N_22392,N_21743,N_21790);
or U22393 (N_22393,N_21939,N_21985);
and U22394 (N_22394,N_21964,N_21536);
and U22395 (N_22395,N_21693,N_21638);
or U22396 (N_22396,N_21691,N_21803);
nor U22397 (N_22397,N_21848,N_21979);
and U22398 (N_22398,N_21809,N_21591);
or U22399 (N_22399,N_21606,N_21639);
xor U22400 (N_22400,N_21968,N_21574);
nor U22401 (N_22401,N_21865,N_21910);
nor U22402 (N_22402,N_21696,N_21713);
nor U22403 (N_22403,N_21770,N_21802);
nand U22404 (N_22404,N_21595,N_21819);
or U22405 (N_22405,N_21757,N_21975);
nand U22406 (N_22406,N_21900,N_21968);
and U22407 (N_22407,N_21705,N_21546);
nor U22408 (N_22408,N_21688,N_21720);
xor U22409 (N_22409,N_21703,N_21892);
and U22410 (N_22410,N_21906,N_21598);
nor U22411 (N_22411,N_21835,N_21608);
nor U22412 (N_22412,N_21886,N_21724);
or U22413 (N_22413,N_21945,N_21897);
nand U22414 (N_22414,N_21704,N_21812);
or U22415 (N_22415,N_21710,N_21861);
xor U22416 (N_22416,N_21810,N_21710);
or U22417 (N_22417,N_21604,N_21652);
or U22418 (N_22418,N_21507,N_21513);
nand U22419 (N_22419,N_21999,N_21569);
and U22420 (N_22420,N_21772,N_21934);
and U22421 (N_22421,N_21680,N_21794);
nor U22422 (N_22422,N_21590,N_21862);
nand U22423 (N_22423,N_21743,N_21996);
nand U22424 (N_22424,N_21706,N_21736);
nor U22425 (N_22425,N_21997,N_21720);
xnor U22426 (N_22426,N_21639,N_21845);
nor U22427 (N_22427,N_21515,N_21960);
nand U22428 (N_22428,N_21670,N_21744);
xnor U22429 (N_22429,N_21866,N_21829);
and U22430 (N_22430,N_21697,N_21526);
xnor U22431 (N_22431,N_21807,N_21741);
nor U22432 (N_22432,N_21994,N_21567);
or U22433 (N_22433,N_21937,N_21785);
xnor U22434 (N_22434,N_21520,N_21934);
nand U22435 (N_22435,N_21854,N_21726);
nor U22436 (N_22436,N_21722,N_21644);
nand U22437 (N_22437,N_21657,N_21996);
xor U22438 (N_22438,N_21811,N_21817);
or U22439 (N_22439,N_21643,N_21721);
and U22440 (N_22440,N_21548,N_21715);
or U22441 (N_22441,N_21964,N_21547);
nand U22442 (N_22442,N_21684,N_21796);
xor U22443 (N_22443,N_21939,N_21934);
nor U22444 (N_22444,N_21775,N_21960);
or U22445 (N_22445,N_21936,N_21796);
nand U22446 (N_22446,N_21716,N_21845);
and U22447 (N_22447,N_21659,N_21839);
or U22448 (N_22448,N_21975,N_21599);
nor U22449 (N_22449,N_21953,N_21768);
nand U22450 (N_22450,N_21549,N_21860);
xnor U22451 (N_22451,N_21528,N_21710);
xnor U22452 (N_22452,N_21947,N_21662);
or U22453 (N_22453,N_21543,N_21742);
nor U22454 (N_22454,N_21868,N_21963);
xnor U22455 (N_22455,N_21659,N_21513);
nand U22456 (N_22456,N_21796,N_21757);
and U22457 (N_22457,N_21851,N_21815);
nand U22458 (N_22458,N_21937,N_21726);
xor U22459 (N_22459,N_21868,N_21530);
and U22460 (N_22460,N_21588,N_21547);
nand U22461 (N_22461,N_21712,N_21586);
xnor U22462 (N_22462,N_21568,N_21760);
nand U22463 (N_22463,N_21646,N_21603);
and U22464 (N_22464,N_21844,N_21999);
or U22465 (N_22465,N_21911,N_21828);
nor U22466 (N_22466,N_21508,N_21688);
xnor U22467 (N_22467,N_21985,N_21652);
nor U22468 (N_22468,N_21582,N_21685);
and U22469 (N_22469,N_21863,N_21567);
nand U22470 (N_22470,N_21887,N_21923);
and U22471 (N_22471,N_21579,N_21509);
nor U22472 (N_22472,N_21800,N_21925);
or U22473 (N_22473,N_21691,N_21618);
nand U22474 (N_22474,N_21809,N_21767);
or U22475 (N_22475,N_21928,N_21525);
nand U22476 (N_22476,N_21554,N_21995);
nand U22477 (N_22477,N_21873,N_21796);
or U22478 (N_22478,N_21777,N_21500);
nand U22479 (N_22479,N_21809,N_21782);
nand U22480 (N_22480,N_21687,N_21772);
nor U22481 (N_22481,N_21697,N_21799);
nand U22482 (N_22482,N_21759,N_21962);
nor U22483 (N_22483,N_21933,N_21714);
nor U22484 (N_22484,N_21845,N_21952);
nor U22485 (N_22485,N_21562,N_21976);
and U22486 (N_22486,N_21985,N_21805);
nand U22487 (N_22487,N_21551,N_21766);
nor U22488 (N_22488,N_21536,N_21936);
or U22489 (N_22489,N_21514,N_21586);
nor U22490 (N_22490,N_21978,N_21510);
nor U22491 (N_22491,N_21667,N_21638);
nor U22492 (N_22492,N_21984,N_21825);
xnor U22493 (N_22493,N_21916,N_21586);
xnor U22494 (N_22494,N_21593,N_21830);
xnor U22495 (N_22495,N_21645,N_21655);
and U22496 (N_22496,N_21682,N_21620);
or U22497 (N_22497,N_21609,N_21834);
nor U22498 (N_22498,N_21611,N_21721);
nor U22499 (N_22499,N_21953,N_21962);
xor U22500 (N_22500,N_22051,N_22337);
and U22501 (N_22501,N_22346,N_22203);
nor U22502 (N_22502,N_22470,N_22303);
xor U22503 (N_22503,N_22386,N_22327);
nand U22504 (N_22504,N_22482,N_22010);
and U22505 (N_22505,N_22160,N_22366);
nor U22506 (N_22506,N_22060,N_22049);
and U22507 (N_22507,N_22493,N_22207);
nand U22508 (N_22508,N_22308,N_22024);
or U22509 (N_22509,N_22251,N_22426);
or U22510 (N_22510,N_22189,N_22157);
or U22511 (N_22511,N_22453,N_22172);
xnor U22512 (N_22512,N_22287,N_22011);
nor U22513 (N_22513,N_22293,N_22295);
xnor U22514 (N_22514,N_22107,N_22204);
and U22515 (N_22515,N_22410,N_22371);
xnor U22516 (N_22516,N_22446,N_22299);
xnor U22517 (N_22517,N_22402,N_22037);
xnor U22518 (N_22518,N_22434,N_22143);
or U22519 (N_22519,N_22377,N_22439);
nand U22520 (N_22520,N_22307,N_22005);
or U22521 (N_22521,N_22266,N_22425);
xnor U22522 (N_22522,N_22075,N_22443);
nor U22523 (N_22523,N_22267,N_22486);
and U22524 (N_22524,N_22286,N_22223);
xnor U22525 (N_22525,N_22045,N_22413);
nand U22526 (N_22526,N_22066,N_22414);
or U22527 (N_22527,N_22310,N_22492);
and U22528 (N_22528,N_22418,N_22008);
nor U22529 (N_22529,N_22082,N_22487);
nor U22530 (N_22530,N_22382,N_22319);
and U22531 (N_22531,N_22369,N_22438);
nor U22532 (N_22532,N_22451,N_22323);
or U22533 (N_22533,N_22372,N_22102);
xnor U22534 (N_22534,N_22000,N_22040);
nor U22535 (N_22535,N_22421,N_22230);
xor U22536 (N_22536,N_22096,N_22312);
or U22537 (N_22537,N_22171,N_22277);
and U22538 (N_22538,N_22103,N_22335);
or U22539 (N_22539,N_22168,N_22450);
xor U22540 (N_22540,N_22021,N_22412);
nand U22541 (N_22541,N_22198,N_22279);
and U22542 (N_22542,N_22136,N_22201);
and U22543 (N_22543,N_22396,N_22113);
nor U22544 (N_22544,N_22359,N_22114);
and U22545 (N_22545,N_22380,N_22056);
and U22546 (N_22546,N_22405,N_22119);
or U22547 (N_22547,N_22383,N_22463);
nand U22548 (N_22548,N_22229,N_22456);
or U22549 (N_22549,N_22078,N_22202);
nor U22550 (N_22550,N_22058,N_22411);
xnor U22551 (N_22551,N_22070,N_22039);
nand U22552 (N_22552,N_22241,N_22027);
xnor U22553 (N_22553,N_22181,N_22407);
or U22554 (N_22554,N_22263,N_22423);
xnor U22555 (N_22555,N_22087,N_22211);
xor U22556 (N_22556,N_22013,N_22406);
nand U22557 (N_22557,N_22080,N_22476);
nand U22558 (N_22558,N_22477,N_22022);
or U22559 (N_22559,N_22111,N_22191);
xor U22560 (N_22560,N_22466,N_22324);
or U22561 (N_22561,N_22064,N_22460);
nand U22562 (N_22562,N_22408,N_22349);
or U22563 (N_22563,N_22442,N_22375);
nor U22564 (N_22564,N_22179,N_22188);
or U22565 (N_22565,N_22393,N_22200);
xnor U22566 (N_22566,N_22081,N_22155);
xor U22567 (N_22567,N_22288,N_22130);
and U22568 (N_22568,N_22294,N_22174);
nand U22569 (N_22569,N_22326,N_22112);
nor U22570 (N_22570,N_22392,N_22355);
or U22571 (N_22571,N_22330,N_22177);
nor U22572 (N_22572,N_22419,N_22305);
nand U22573 (N_22573,N_22069,N_22395);
nand U22574 (N_22574,N_22213,N_22120);
nand U22575 (N_22575,N_22212,N_22334);
nand U22576 (N_22576,N_22398,N_22048);
and U22577 (N_22577,N_22462,N_22276);
nand U22578 (N_22578,N_22313,N_22497);
xnor U22579 (N_22579,N_22148,N_22253);
or U22580 (N_22580,N_22141,N_22445);
nor U22581 (N_22581,N_22031,N_22131);
and U22582 (N_22582,N_22135,N_22220);
or U22583 (N_22583,N_22248,N_22165);
nand U22584 (N_22584,N_22360,N_22234);
nor U22585 (N_22585,N_22199,N_22225);
or U22586 (N_22586,N_22226,N_22127);
nand U22587 (N_22587,N_22257,N_22153);
nand U22588 (N_22588,N_22218,N_22318);
nor U22589 (N_22589,N_22256,N_22317);
xnor U22590 (N_22590,N_22245,N_22014);
and U22591 (N_22591,N_22347,N_22283);
nand U22592 (N_22592,N_22457,N_22481);
or U22593 (N_22593,N_22101,N_22381);
or U22594 (N_22594,N_22321,N_22092);
nor U22595 (N_22595,N_22166,N_22314);
or U22596 (N_22596,N_22416,N_22126);
xnor U22597 (N_22597,N_22164,N_22169);
xnor U22598 (N_22598,N_22026,N_22053);
nor U22599 (N_22599,N_22015,N_22292);
xnor U22600 (N_22600,N_22154,N_22338);
or U22601 (N_22601,N_22133,N_22440);
nor U22602 (N_22602,N_22067,N_22478);
nor U22603 (N_22603,N_22361,N_22029);
nor U22604 (N_22604,N_22345,N_22271);
xor U22605 (N_22605,N_22291,N_22176);
and U22606 (N_22606,N_22259,N_22304);
nand U22607 (N_22607,N_22047,N_22054);
or U22608 (N_22608,N_22122,N_22044);
or U22609 (N_22609,N_22083,N_22163);
xor U22610 (N_22610,N_22261,N_22274);
xnor U22611 (N_22611,N_22142,N_22062);
xor U22612 (N_22612,N_22394,N_22252);
or U22613 (N_22613,N_22184,N_22296);
and U22614 (N_22614,N_22246,N_22433);
nand U22615 (N_22615,N_22461,N_22353);
nor U22616 (N_22616,N_22084,N_22185);
nor U22617 (N_22617,N_22422,N_22273);
and U22618 (N_22618,N_22221,N_22227);
or U22619 (N_22619,N_22139,N_22329);
xnor U22620 (N_22620,N_22238,N_22140);
and U22621 (N_22621,N_22437,N_22237);
or U22622 (N_22622,N_22264,N_22480);
nand U22623 (N_22623,N_22354,N_22363);
or U22624 (N_22624,N_22068,N_22384);
and U22625 (N_22625,N_22289,N_22280);
nor U22626 (N_22626,N_22452,N_22290);
and U22627 (N_22627,N_22239,N_22236);
xor U22628 (N_22628,N_22400,N_22332);
xor U22629 (N_22629,N_22182,N_22004);
xnor U22630 (N_22630,N_22025,N_22028);
or U22631 (N_22631,N_22489,N_22086);
xnor U22632 (N_22632,N_22232,N_22233);
nor U22633 (N_22633,N_22298,N_22485);
and U22634 (N_22634,N_22344,N_22228);
xnor U22635 (N_22635,N_22214,N_22195);
nor U22636 (N_22636,N_22124,N_22151);
and U22637 (N_22637,N_22357,N_22333);
or U22638 (N_22638,N_22468,N_22138);
nor U22639 (N_22639,N_22156,N_22217);
and U22640 (N_22640,N_22275,N_22018);
xnor U22641 (N_22641,N_22250,N_22073);
nor U22642 (N_22642,N_22108,N_22090);
or U22643 (N_22643,N_22301,N_22186);
and U22644 (N_22644,N_22061,N_22038);
or U22645 (N_22645,N_22210,N_22424);
nor U22646 (N_22646,N_22254,N_22474);
nand U22647 (N_22647,N_22336,N_22340);
and U22648 (N_22648,N_22429,N_22115);
xor U22649 (N_22649,N_22269,N_22149);
or U22650 (N_22650,N_22192,N_22285);
nor U22651 (N_22651,N_22311,N_22365);
xor U22652 (N_22652,N_22399,N_22041);
nand U22653 (N_22653,N_22343,N_22183);
nand U22654 (N_22654,N_22469,N_22484);
or U22655 (N_22655,N_22170,N_22465);
and U22656 (N_22656,N_22282,N_22322);
xor U22657 (N_22657,N_22494,N_22435);
or U22658 (N_22658,N_22430,N_22243);
nor U22659 (N_22659,N_22499,N_22417);
nand U22660 (N_22660,N_22428,N_22125);
nand U22661 (N_22661,N_22094,N_22328);
nor U22662 (N_22662,N_22089,N_22331);
or U22663 (N_22663,N_22215,N_22222);
nor U22664 (N_22664,N_22352,N_22196);
nor U22665 (N_22665,N_22441,N_22074);
or U22666 (N_22666,N_22093,N_22046);
or U22667 (N_22667,N_22475,N_22072);
nor U22668 (N_22668,N_22098,N_22023);
nand U22669 (N_22669,N_22284,N_22281);
or U22670 (N_22670,N_22490,N_22091);
nand U22671 (N_22671,N_22001,N_22432);
nand U22672 (N_22672,N_22231,N_22118);
and U22673 (N_22673,N_22358,N_22052);
xnor U22674 (N_22674,N_22260,N_22496);
xor U22675 (N_22675,N_22265,N_22244);
or U22676 (N_22676,N_22491,N_22187);
and U22677 (N_22677,N_22455,N_22495);
nor U22678 (N_22678,N_22444,N_22071);
and U22679 (N_22679,N_22077,N_22117);
nor U22680 (N_22680,N_22178,N_22158);
xor U22681 (N_22681,N_22309,N_22379);
and U22682 (N_22682,N_22368,N_22348);
nor U22683 (N_22683,N_22016,N_22255);
xnor U22684 (N_22684,N_22473,N_22247);
and U22685 (N_22685,N_22454,N_22272);
or U22686 (N_22686,N_22055,N_22076);
xor U22687 (N_22687,N_22162,N_22036);
nor U22688 (N_22688,N_22403,N_22144);
nand U22689 (N_22689,N_22216,N_22219);
and U22690 (N_22690,N_22009,N_22088);
or U22691 (N_22691,N_22161,N_22063);
nand U22692 (N_22692,N_22159,N_22415);
or U22693 (N_22693,N_22459,N_22110);
or U22694 (N_22694,N_22373,N_22258);
nor U22695 (N_22695,N_22409,N_22387);
and U22696 (N_22696,N_22132,N_22150);
xor U22697 (N_22697,N_22351,N_22129);
nand U22698 (N_22698,N_22034,N_22472);
nor U22699 (N_22699,N_22109,N_22471);
xnor U22700 (N_22700,N_22306,N_22370);
nor U22701 (N_22701,N_22197,N_22145);
or U22702 (N_22702,N_22033,N_22123);
or U22703 (N_22703,N_22003,N_22364);
nor U22704 (N_22704,N_22085,N_22262);
nor U22705 (N_22705,N_22106,N_22479);
nand U22706 (N_22706,N_22362,N_22240);
or U22707 (N_22707,N_22356,N_22099);
and U22708 (N_22708,N_22391,N_22374);
xor U22709 (N_22709,N_22190,N_22042);
nor U22710 (N_22710,N_22006,N_22019);
and U22711 (N_22711,N_22205,N_22390);
or U22712 (N_22712,N_22173,N_22208);
and U22713 (N_22713,N_22128,N_22137);
nor U22714 (N_22714,N_22095,N_22104);
nand U22715 (N_22715,N_22341,N_22035);
xnor U22716 (N_22716,N_22467,N_22017);
nor U22717 (N_22717,N_22079,N_22209);
xor U22718 (N_22718,N_22376,N_22134);
and U22719 (N_22719,N_22146,N_22350);
or U22720 (N_22720,N_22249,N_22397);
and U22721 (N_22721,N_22206,N_22427);
nand U22722 (N_22722,N_22235,N_22320);
nand U22723 (N_22723,N_22032,N_22447);
and U22724 (N_22724,N_22498,N_22278);
xnor U22725 (N_22725,N_22488,N_22325);
or U22726 (N_22726,N_22147,N_22002);
nor U22727 (N_22727,N_22300,N_22302);
nand U22728 (N_22728,N_22464,N_22043);
nor U22729 (N_22729,N_22224,N_22050);
or U22730 (N_22730,N_22007,N_22458);
and U22731 (N_22731,N_22097,N_22436);
or U22732 (N_22732,N_22448,N_22404);
xor U22733 (N_22733,N_22268,N_22012);
nand U22734 (N_22734,N_22389,N_22194);
nor U22735 (N_22735,N_22121,N_22242);
or U22736 (N_22736,N_22431,N_22367);
and U22737 (N_22737,N_22180,N_22449);
nand U22738 (N_22738,N_22193,N_22100);
or U22739 (N_22739,N_22059,N_22315);
nand U22740 (N_22740,N_22388,N_22270);
xor U22741 (N_22741,N_22297,N_22020);
or U22742 (N_22742,N_22483,N_22057);
xnor U22743 (N_22743,N_22167,N_22401);
or U22744 (N_22744,N_22030,N_22342);
or U22745 (N_22745,N_22339,N_22105);
and U22746 (N_22746,N_22152,N_22378);
xnor U22747 (N_22747,N_22065,N_22420);
and U22748 (N_22748,N_22316,N_22175);
nor U22749 (N_22749,N_22116,N_22385);
or U22750 (N_22750,N_22376,N_22222);
and U22751 (N_22751,N_22089,N_22453);
and U22752 (N_22752,N_22103,N_22138);
nand U22753 (N_22753,N_22475,N_22417);
xnor U22754 (N_22754,N_22266,N_22482);
nor U22755 (N_22755,N_22403,N_22239);
xor U22756 (N_22756,N_22211,N_22253);
or U22757 (N_22757,N_22211,N_22423);
or U22758 (N_22758,N_22434,N_22230);
xnor U22759 (N_22759,N_22158,N_22190);
nor U22760 (N_22760,N_22277,N_22223);
nor U22761 (N_22761,N_22448,N_22381);
or U22762 (N_22762,N_22032,N_22072);
nor U22763 (N_22763,N_22473,N_22089);
xor U22764 (N_22764,N_22443,N_22224);
or U22765 (N_22765,N_22378,N_22361);
nand U22766 (N_22766,N_22356,N_22400);
nand U22767 (N_22767,N_22384,N_22456);
and U22768 (N_22768,N_22056,N_22492);
nand U22769 (N_22769,N_22159,N_22270);
or U22770 (N_22770,N_22433,N_22448);
and U22771 (N_22771,N_22106,N_22089);
nand U22772 (N_22772,N_22242,N_22190);
nand U22773 (N_22773,N_22428,N_22115);
nand U22774 (N_22774,N_22137,N_22255);
and U22775 (N_22775,N_22104,N_22357);
or U22776 (N_22776,N_22086,N_22327);
nor U22777 (N_22777,N_22432,N_22376);
and U22778 (N_22778,N_22226,N_22009);
or U22779 (N_22779,N_22137,N_22103);
xor U22780 (N_22780,N_22395,N_22421);
nor U22781 (N_22781,N_22067,N_22332);
or U22782 (N_22782,N_22130,N_22264);
and U22783 (N_22783,N_22490,N_22071);
xnor U22784 (N_22784,N_22192,N_22434);
nor U22785 (N_22785,N_22362,N_22272);
nor U22786 (N_22786,N_22083,N_22405);
or U22787 (N_22787,N_22185,N_22474);
or U22788 (N_22788,N_22396,N_22484);
nand U22789 (N_22789,N_22413,N_22214);
xnor U22790 (N_22790,N_22196,N_22261);
and U22791 (N_22791,N_22475,N_22199);
nand U22792 (N_22792,N_22343,N_22494);
nand U22793 (N_22793,N_22080,N_22388);
nor U22794 (N_22794,N_22066,N_22305);
nand U22795 (N_22795,N_22021,N_22318);
nand U22796 (N_22796,N_22391,N_22355);
nand U22797 (N_22797,N_22091,N_22351);
and U22798 (N_22798,N_22002,N_22221);
nand U22799 (N_22799,N_22213,N_22419);
nor U22800 (N_22800,N_22247,N_22076);
and U22801 (N_22801,N_22046,N_22305);
xnor U22802 (N_22802,N_22165,N_22437);
nand U22803 (N_22803,N_22460,N_22341);
nand U22804 (N_22804,N_22458,N_22373);
and U22805 (N_22805,N_22101,N_22284);
xor U22806 (N_22806,N_22436,N_22488);
nand U22807 (N_22807,N_22399,N_22470);
nor U22808 (N_22808,N_22395,N_22477);
and U22809 (N_22809,N_22370,N_22365);
and U22810 (N_22810,N_22043,N_22354);
nand U22811 (N_22811,N_22284,N_22482);
or U22812 (N_22812,N_22495,N_22359);
and U22813 (N_22813,N_22253,N_22259);
and U22814 (N_22814,N_22026,N_22295);
nor U22815 (N_22815,N_22164,N_22059);
nor U22816 (N_22816,N_22399,N_22117);
nor U22817 (N_22817,N_22052,N_22442);
nor U22818 (N_22818,N_22045,N_22172);
nor U22819 (N_22819,N_22205,N_22461);
nor U22820 (N_22820,N_22278,N_22436);
nor U22821 (N_22821,N_22382,N_22095);
nand U22822 (N_22822,N_22281,N_22401);
or U22823 (N_22823,N_22444,N_22035);
and U22824 (N_22824,N_22011,N_22378);
xor U22825 (N_22825,N_22269,N_22303);
xnor U22826 (N_22826,N_22456,N_22275);
or U22827 (N_22827,N_22006,N_22446);
nor U22828 (N_22828,N_22147,N_22361);
and U22829 (N_22829,N_22405,N_22147);
xor U22830 (N_22830,N_22272,N_22092);
or U22831 (N_22831,N_22209,N_22328);
xor U22832 (N_22832,N_22083,N_22118);
nand U22833 (N_22833,N_22122,N_22353);
and U22834 (N_22834,N_22050,N_22295);
or U22835 (N_22835,N_22362,N_22047);
xnor U22836 (N_22836,N_22048,N_22077);
and U22837 (N_22837,N_22302,N_22409);
and U22838 (N_22838,N_22448,N_22411);
and U22839 (N_22839,N_22332,N_22435);
xnor U22840 (N_22840,N_22310,N_22317);
xnor U22841 (N_22841,N_22002,N_22375);
or U22842 (N_22842,N_22085,N_22155);
and U22843 (N_22843,N_22233,N_22369);
nand U22844 (N_22844,N_22228,N_22286);
nor U22845 (N_22845,N_22000,N_22435);
nor U22846 (N_22846,N_22098,N_22358);
nand U22847 (N_22847,N_22422,N_22194);
nor U22848 (N_22848,N_22414,N_22261);
and U22849 (N_22849,N_22262,N_22280);
and U22850 (N_22850,N_22212,N_22102);
nand U22851 (N_22851,N_22045,N_22374);
and U22852 (N_22852,N_22446,N_22321);
nor U22853 (N_22853,N_22080,N_22410);
and U22854 (N_22854,N_22324,N_22123);
nor U22855 (N_22855,N_22404,N_22325);
nor U22856 (N_22856,N_22427,N_22395);
or U22857 (N_22857,N_22214,N_22245);
and U22858 (N_22858,N_22118,N_22315);
and U22859 (N_22859,N_22276,N_22307);
or U22860 (N_22860,N_22289,N_22156);
and U22861 (N_22861,N_22234,N_22024);
nand U22862 (N_22862,N_22138,N_22433);
and U22863 (N_22863,N_22107,N_22381);
nand U22864 (N_22864,N_22459,N_22114);
nor U22865 (N_22865,N_22312,N_22153);
xor U22866 (N_22866,N_22323,N_22374);
xnor U22867 (N_22867,N_22203,N_22497);
and U22868 (N_22868,N_22333,N_22132);
and U22869 (N_22869,N_22137,N_22029);
or U22870 (N_22870,N_22435,N_22311);
xnor U22871 (N_22871,N_22494,N_22490);
xor U22872 (N_22872,N_22072,N_22439);
xnor U22873 (N_22873,N_22353,N_22294);
nand U22874 (N_22874,N_22442,N_22458);
nor U22875 (N_22875,N_22191,N_22486);
nand U22876 (N_22876,N_22291,N_22184);
and U22877 (N_22877,N_22456,N_22122);
nand U22878 (N_22878,N_22096,N_22362);
or U22879 (N_22879,N_22401,N_22341);
xor U22880 (N_22880,N_22123,N_22335);
and U22881 (N_22881,N_22174,N_22079);
nand U22882 (N_22882,N_22488,N_22250);
or U22883 (N_22883,N_22067,N_22087);
nand U22884 (N_22884,N_22103,N_22014);
and U22885 (N_22885,N_22487,N_22108);
or U22886 (N_22886,N_22157,N_22371);
and U22887 (N_22887,N_22428,N_22000);
xnor U22888 (N_22888,N_22095,N_22087);
or U22889 (N_22889,N_22286,N_22376);
xnor U22890 (N_22890,N_22099,N_22313);
xnor U22891 (N_22891,N_22095,N_22141);
xnor U22892 (N_22892,N_22290,N_22440);
and U22893 (N_22893,N_22370,N_22048);
and U22894 (N_22894,N_22109,N_22193);
and U22895 (N_22895,N_22430,N_22070);
nand U22896 (N_22896,N_22017,N_22070);
nand U22897 (N_22897,N_22294,N_22324);
xnor U22898 (N_22898,N_22461,N_22382);
and U22899 (N_22899,N_22250,N_22400);
and U22900 (N_22900,N_22440,N_22174);
nor U22901 (N_22901,N_22048,N_22180);
or U22902 (N_22902,N_22141,N_22370);
nand U22903 (N_22903,N_22113,N_22403);
nor U22904 (N_22904,N_22218,N_22459);
or U22905 (N_22905,N_22406,N_22465);
nand U22906 (N_22906,N_22026,N_22334);
and U22907 (N_22907,N_22401,N_22051);
nor U22908 (N_22908,N_22286,N_22347);
or U22909 (N_22909,N_22161,N_22474);
nor U22910 (N_22910,N_22347,N_22354);
xor U22911 (N_22911,N_22302,N_22299);
and U22912 (N_22912,N_22444,N_22318);
nor U22913 (N_22913,N_22096,N_22167);
or U22914 (N_22914,N_22348,N_22204);
or U22915 (N_22915,N_22408,N_22198);
or U22916 (N_22916,N_22348,N_22207);
nand U22917 (N_22917,N_22363,N_22287);
xnor U22918 (N_22918,N_22343,N_22481);
or U22919 (N_22919,N_22022,N_22305);
and U22920 (N_22920,N_22435,N_22056);
and U22921 (N_22921,N_22130,N_22028);
and U22922 (N_22922,N_22443,N_22472);
or U22923 (N_22923,N_22342,N_22464);
or U22924 (N_22924,N_22454,N_22260);
nor U22925 (N_22925,N_22369,N_22041);
or U22926 (N_22926,N_22248,N_22414);
nand U22927 (N_22927,N_22468,N_22276);
xnor U22928 (N_22928,N_22032,N_22283);
or U22929 (N_22929,N_22217,N_22092);
and U22930 (N_22930,N_22306,N_22212);
and U22931 (N_22931,N_22342,N_22255);
or U22932 (N_22932,N_22340,N_22186);
and U22933 (N_22933,N_22248,N_22281);
nor U22934 (N_22934,N_22310,N_22105);
and U22935 (N_22935,N_22131,N_22392);
nand U22936 (N_22936,N_22130,N_22025);
xor U22937 (N_22937,N_22335,N_22281);
nor U22938 (N_22938,N_22256,N_22265);
or U22939 (N_22939,N_22065,N_22238);
and U22940 (N_22940,N_22081,N_22291);
and U22941 (N_22941,N_22355,N_22457);
xor U22942 (N_22942,N_22307,N_22060);
or U22943 (N_22943,N_22320,N_22078);
and U22944 (N_22944,N_22343,N_22442);
xor U22945 (N_22945,N_22252,N_22051);
nand U22946 (N_22946,N_22006,N_22215);
or U22947 (N_22947,N_22257,N_22104);
nand U22948 (N_22948,N_22257,N_22487);
and U22949 (N_22949,N_22410,N_22037);
or U22950 (N_22950,N_22147,N_22160);
and U22951 (N_22951,N_22276,N_22152);
or U22952 (N_22952,N_22161,N_22483);
and U22953 (N_22953,N_22387,N_22050);
and U22954 (N_22954,N_22446,N_22285);
xnor U22955 (N_22955,N_22012,N_22048);
nand U22956 (N_22956,N_22077,N_22132);
and U22957 (N_22957,N_22194,N_22092);
nand U22958 (N_22958,N_22041,N_22156);
nor U22959 (N_22959,N_22232,N_22331);
and U22960 (N_22960,N_22499,N_22451);
or U22961 (N_22961,N_22401,N_22479);
or U22962 (N_22962,N_22391,N_22045);
nor U22963 (N_22963,N_22192,N_22145);
xnor U22964 (N_22964,N_22027,N_22152);
xor U22965 (N_22965,N_22043,N_22308);
nand U22966 (N_22966,N_22359,N_22422);
xor U22967 (N_22967,N_22494,N_22293);
xnor U22968 (N_22968,N_22492,N_22400);
nor U22969 (N_22969,N_22324,N_22204);
or U22970 (N_22970,N_22362,N_22175);
or U22971 (N_22971,N_22404,N_22180);
xor U22972 (N_22972,N_22063,N_22196);
xnor U22973 (N_22973,N_22273,N_22299);
and U22974 (N_22974,N_22409,N_22051);
and U22975 (N_22975,N_22226,N_22276);
xor U22976 (N_22976,N_22296,N_22289);
and U22977 (N_22977,N_22275,N_22293);
and U22978 (N_22978,N_22460,N_22006);
or U22979 (N_22979,N_22314,N_22104);
nor U22980 (N_22980,N_22336,N_22093);
nor U22981 (N_22981,N_22259,N_22340);
nand U22982 (N_22982,N_22147,N_22316);
nor U22983 (N_22983,N_22148,N_22340);
nor U22984 (N_22984,N_22366,N_22323);
nand U22985 (N_22985,N_22442,N_22067);
nor U22986 (N_22986,N_22294,N_22172);
or U22987 (N_22987,N_22031,N_22446);
and U22988 (N_22988,N_22356,N_22399);
or U22989 (N_22989,N_22196,N_22303);
nand U22990 (N_22990,N_22094,N_22368);
nor U22991 (N_22991,N_22459,N_22111);
xor U22992 (N_22992,N_22360,N_22335);
and U22993 (N_22993,N_22164,N_22141);
or U22994 (N_22994,N_22060,N_22320);
nand U22995 (N_22995,N_22441,N_22088);
nor U22996 (N_22996,N_22088,N_22006);
xor U22997 (N_22997,N_22133,N_22217);
nor U22998 (N_22998,N_22416,N_22264);
nand U22999 (N_22999,N_22083,N_22093);
or U23000 (N_23000,N_22929,N_22572);
and U23001 (N_23001,N_22720,N_22701);
xnor U23002 (N_23002,N_22603,N_22887);
xor U23003 (N_23003,N_22944,N_22678);
xor U23004 (N_23004,N_22522,N_22732);
or U23005 (N_23005,N_22573,N_22518);
and U23006 (N_23006,N_22948,N_22924);
nand U23007 (N_23007,N_22731,N_22846);
xnor U23008 (N_23008,N_22647,N_22875);
xnor U23009 (N_23009,N_22844,N_22801);
and U23010 (N_23010,N_22606,N_22763);
and U23011 (N_23011,N_22515,N_22639);
nor U23012 (N_23012,N_22992,N_22920);
xor U23013 (N_23013,N_22797,N_22636);
nand U23014 (N_23014,N_22661,N_22957);
or U23015 (N_23015,N_22770,N_22922);
xnor U23016 (N_23016,N_22514,N_22824);
or U23017 (N_23017,N_22857,N_22580);
xnor U23018 (N_23018,N_22987,N_22628);
or U23019 (N_23019,N_22511,N_22818);
xor U23020 (N_23020,N_22897,N_22783);
and U23021 (N_23021,N_22733,N_22809);
nand U23022 (N_23022,N_22608,N_22512);
xor U23023 (N_23023,N_22830,N_22832);
or U23024 (N_23024,N_22802,N_22510);
nand U23025 (N_23025,N_22791,N_22868);
or U23026 (N_23026,N_22549,N_22737);
or U23027 (N_23027,N_22735,N_22528);
or U23028 (N_23028,N_22727,N_22506);
nand U23029 (N_23029,N_22914,N_22590);
xor U23030 (N_23030,N_22880,N_22937);
or U23031 (N_23031,N_22805,N_22680);
nor U23032 (N_23032,N_22718,N_22691);
xnor U23033 (N_23033,N_22675,N_22671);
nor U23034 (N_23034,N_22738,N_22699);
nand U23035 (N_23035,N_22909,N_22520);
xor U23036 (N_23036,N_22531,N_22593);
xor U23037 (N_23037,N_22988,N_22625);
nand U23038 (N_23038,N_22570,N_22978);
and U23039 (N_23039,N_22577,N_22838);
xor U23040 (N_23040,N_22643,N_22670);
and U23041 (N_23041,N_22888,N_22911);
nand U23042 (N_23042,N_22503,N_22660);
nor U23043 (N_23043,N_22757,N_22779);
or U23044 (N_23044,N_22833,N_22991);
and U23045 (N_23045,N_22772,N_22652);
or U23046 (N_23046,N_22941,N_22508);
nand U23047 (N_23047,N_22672,N_22509);
or U23048 (N_23048,N_22867,N_22782);
xor U23049 (N_23049,N_22777,N_22710);
xnor U23050 (N_23050,N_22650,N_22600);
xnor U23051 (N_23051,N_22954,N_22613);
nor U23052 (N_23052,N_22778,N_22711);
or U23053 (N_23053,N_22861,N_22989);
nand U23054 (N_23054,N_22898,N_22975);
or U23055 (N_23055,N_22693,N_22624);
and U23056 (N_23056,N_22877,N_22912);
xor U23057 (N_23057,N_22513,N_22827);
or U23058 (N_23058,N_22690,N_22649);
nand U23059 (N_23059,N_22744,N_22872);
or U23060 (N_23060,N_22768,N_22984);
xor U23061 (N_23061,N_22709,N_22949);
nand U23062 (N_23062,N_22554,N_22663);
nor U23063 (N_23063,N_22794,N_22621);
nor U23064 (N_23064,N_22574,N_22705);
and U23065 (N_23065,N_22607,N_22754);
nor U23066 (N_23066,N_22773,N_22673);
or U23067 (N_23067,N_22635,N_22545);
or U23068 (N_23068,N_22592,N_22595);
nand U23069 (N_23069,N_22790,N_22740);
nand U23070 (N_23070,N_22906,N_22681);
xor U23071 (N_23071,N_22713,N_22816);
nor U23072 (N_23072,N_22622,N_22708);
or U23073 (N_23073,N_22764,N_22747);
nor U23074 (N_23074,N_22532,N_22524);
or U23075 (N_23075,N_22537,N_22535);
or U23076 (N_23076,N_22676,N_22866);
and U23077 (N_23077,N_22964,N_22615);
nor U23078 (N_23078,N_22874,N_22752);
and U23079 (N_23079,N_22891,N_22729);
and U23080 (N_23080,N_22536,N_22589);
xnor U23081 (N_23081,N_22961,N_22905);
xnor U23082 (N_23082,N_22999,N_22556);
nor U23083 (N_23083,N_22793,N_22851);
xor U23084 (N_23084,N_22565,N_22665);
nor U23085 (N_23085,N_22934,N_22677);
or U23086 (N_23086,N_22938,N_22585);
xor U23087 (N_23087,N_22553,N_22637);
nor U23088 (N_23088,N_22655,N_22835);
and U23089 (N_23089,N_22594,N_22605);
nand U23090 (N_23090,N_22766,N_22881);
xor U23091 (N_23091,N_22767,N_22576);
nor U23092 (N_23092,N_22819,N_22943);
or U23093 (N_23093,N_22958,N_22582);
and U23094 (N_23094,N_22697,N_22942);
nor U23095 (N_23095,N_22630,N_22960);
nor U23096 (N_23096,N_22684,N_22662);
xor U23097 (N_23097,N_22599,N_22979);
nor U23098 (N_23098,N_22908,N_22784);
xor U23099 (N_23099,N_22560,N_22596);
nor U23100 (N_23100,N_22631,N_22858);
xor U23101 (N_23101,N_22581,N_22762);
nand U23102 (N_23102,N_22626,N_22623);
nor U23103 (N_23103,N_22947,N_22856);
and U23104 (N_23104,N_22564,N_22946);
xnor U23105 (N_23105,N_22940,N_22583);
nand U23106 (N_23106,N_22952,N_22945);
nor U23107 (N_23107,N_22745,N_22657);
xnor U23108 (N_23108,N_22935,N_22847);
xnor U23109 (N_23109,N_22633,N_22902);
and U23110 (N_23110,N_22865,N_22561);
xor U23111 (N_23111,N_22529,N_22955);
nor U23112 (N_23112,N_22789,N_22883);
nor U23113 (N_23113,N_22656,N_22698);
or U23114 (N_23114,N_22870,N_22916);
or U23115 (N_23115,N_22559,N_22893);
xnor U23116 (N_23116,N_22533,N_22927);
xnor U23117 (N_23117,N_22602,N_22775);
xnor U23118 (N_23118,N_22640,N_22967);
or U23119 (N_23119,N_22724,N_22569);
nand U23120 (N_23120,N_22525,N_22667);
and U23121 (N_23121,N_22831,N_22892);
or U23122 (N_23122,N_22848,N_22776);
xnor U23123 (N_23123,N_22526,N_22632);
nor U23124 (N_23124,N_22546,N_22983);
or U23125 (N_23125,N_22871,N_22562);
and U23126 (N_23126,N_22849,N_22803);
xor U23127 (N_23127,N_22743,N_22540);
xor U23128 (N_23128,N_22879,N_22939);
or U23129 (N_23129,N_22800,N_22899);
or U23130 (N_23130,N_22996,N_22980);
nand U23131 (N_23131,N_22785,N_22760);
nor U23132 (N_23132,N_22959,N_22646);
nor U23133 (N_23133,N_22900,N_22811);
and U23134 (N_23134,N_22878,N_22521);
or U23135 (N_23135,N_22716,N_22627);
xnor U23136 (N_23136,N_22588,N_22771);
nand U23137 (N_23137,N_22629,N_22828);
nor U23138 (N_23138,N_22921,N_22993);
or U23139 (N_23139,N_22972,N_22923);
nor U23140 (N_23140,N_22799,N_22842);
xnor U23141 (N_23141,N_22571,N_22703);
xnor U23142 (N_23142,N_22834,N_22555);
nor U23143 (N_23143,N_22516,N_22689);
nand U23144 (N_23144,N_22704,N_22981);
and U23145 (N_23145,N_22885,N_22926);
or U23146 (N_23146,N_22931,N_22517);
nor U23147 (N_23147,N_22558,N_22541);
and U23148 (N_23148,N_22659,N_22837);
nand U23149 (N_23149,N_22601,N_22507);
or U23150 (N_23150,N_22956,N_22542);
and U23151 (N_23151,N_22820,N_22933);
nand U23152 (N_23152,N_22666,N_22829);
or U23153 (N_23153,N_22813,N_22694);
xnor U23154 (N_23154,N_22895,N_22951);
nand U23155 (N_23155,N_22527,N_22750);
or U23156 (N_23156,N_22700,N_22519);
or U23157 (N_23157,N_22758,N_22505);
nand U23158 (N_23158,N_22642,N_22557);
or U23159 (N_23159,N_22853,N_22976);
nand U23160 (N_23160,N_22994,N_22548);
xor U23161 (N_23161,N_22859,N_22714);
or U23162 (N_23162,N_22774,N_22712);
xnor U23163 (N_23163,N_22918,N_22982);
nor U23164 (N_23164,N_22917,N_22925);
nor U23165 (N_23165,N_22974,N_22502);
xnor U23166 (N_23166,N_22610,N_22688);
nor U23167 (N_23167,N_22840,N_22598);
nor U23168 (N_23168,N_22682,N_22687);
nor U23169 (N_23169,N_22668,N_22810);
and U23170 (N_23170,N_22812,N_22741);
and U23171 (N_23171,N_22932,N_22604);
xor U23172 (N_23172,N_22852,N_22616);
and U23173 (N_23173,N_22873,N_22634);
nor U23174 (N_23174,N_22806,N_22586);
or U23175 (N_23175,N_22686,N_22904);
nand U23176 (N_23176,N_22817,N_22619);
nor U23177 (N_23177,N_22567,N_22886);
nand U23178 (N_23178,N_22769,N_22910);
nand U23179 (N_23179,N_22584,N_22970);
xor U23180 (N_23180,N_22674,N_22756);
or U23181 (N_23181,N_22751,N_22845);
and U23182 (N_23182,N_22901,N_22950);
nand U23183 (N_23183,N_22651,N_22971);
or U23184 (N_23184,N_22696,N_22836);
or U23185 (N_23185,N_22882,N_22579);
or U23186 (N_23186,N_22706,N_22578);
xor U23187 (N_23187,N_22814,N_22826);
xor U23188 (N_23188,N_22587,N_22547);
and U23189 (N_23189,N_22550,N_22930);
nor U23190 (N_23190,N_22761,N_22860);
and U23191 (N_23191,N_22841,N_22614);
and U23192 (N_23192,N_22719,N_22780);
nor U23193 (N_23193,N_22692,N_22796);
and U23194 (N_23194,N_22641,N_22749);
or U23195 (N_23195,N_22739,N_22617);
nor U23196 (N_23196,N_22990,N_22968);
nor U23197 (N_23197,N_22591,N_22755);
and U23198 (N_23198,N_22855,N_22715);
or U23199 (N_23199,N_22742,N_22977);
nand U23200 (N_23200,N_22850,N_22903);
or U23201 (N_23201,N_22539,N_22753);
xnor U23202 (N_23202,N_22915,N_22620);
nor U23203 (N_23203,N_22566,N_22889);
nor U23204 (N_23204,N_22707,N_22721);
nand U23205 (N_23205,N_22736,N_22597);
nor U23206 (N_23206,N_22658,N_22965);
or U23207 (N_23207,N_22759,N_22702);
and U23208 (N_23208,N_22618,N_22876);
nor U23209 (N_23209,N_22786,N_22890);
nand U23210 (N_23210,N_22504,N_22725);
and U23211 (N_23211,N_22962,N_22534);
and U23212 (N_23212,N_22611,N_22734);
nand U23213 (N_23213,N_22685,N_22723);
or U23214 (N_23214,N_22523,N_22843);
and U23215 (N_23215,N_22501,N_22966);
and U23216 (N_23216,N_22695,N_22664);
and U23217 (N_23217,N_22612,N_22815);
nand U23218 (N_23218,N_22798,N_22995);
xor U23219 (N_23219,N_22653,N_22748);
nor U23220 (N_23220,N_22645,N_22808);
and U23221 (N_23221,N_22854,N_22969);
nor U23222 (N_23222,N_22936,N_22538);
nand U23223 (N_23223,N_22804,N_22551);
and U23224 (N_23224,N_22654,N_22973);
nand U23225 (N_23225,N_22807,N_22896);
or U23226 (N_23226,N_22869,N_22726);
and U23227 (N_23227,N_22822,N_22862);
xor U23228 (N_23228,N_22717,N_22638);
xor U23229 (N_23229,N_22679,N_22928);
nor U23230 (N_23230,N_22894,N_22543);
nand U23231 (N_23231,N_22568,N_22722);
xor U23232 (N_23232,N_22839,N_22746);
or U23233 (N_23233,N_22795,N_22644);
xnor U23234 (N_23234,N_22919,N_22864);
or U23235 (N_23235,N_22683,N_22765);
nor U23236 (N_23236,N_22730,N_22552);
xnor U23237 (N_23237,N_22985,N_22963);
and U23238 (N_23238,N_22986,N_22792);
and U23239 (N_23239,N_22787,N_22648);
or U23240 (N_23240,N_22825,N_22821);
or U23241 (N_23241,N_22823,N_22781);
nand U23242 (N_23242,N_22575,N_22544);
or U23243 (N_23243,N_22953,N_22563);
xnor U23244 (N_23244,N_22997,N_22728);
nor U23245 (N_23245,N_22500,N_22669);
nor U23246 (N_23246,N_22609,N_22863);
or U23247 (N_23247,N_22788,N_22907);
nor U23248 (N_23248,N_22913,N_22884);
nor U23249 (N_23249,N_22998,N_22530);
and U23250 (N_23250,N_22602,N_22805);
and U23251 (N_23251,N_22881,N_22807);
and U23252 (N_23252,N_22923,N_22584);
or U23253 (N_23253,N_22500,N_22546);
nand U23254 (N_23254,N_22957,N_22689);
nand U23255 (N_23255,N_22830,N_22580);
xor U23256 (N_23256,N_22864,N_22543);
nand U23257 (N_23257,N_22670,N_22836);
and U23258 (N_23258,N_22522,N_22507);
nor U23259 (N_23259,N_22599,N_22726);
or U23260 (N_23260,N_22835,N_22922);
nor U23261 (N_23261,N_22838,N_22994);
or U23262 (N_23262,N_22711,N_22871);
nand U23263 (N_23263,N_22957,N_22733);
xor U23264 (N_23264,N_22976,N_22948);
xnor U23265 (N_23265,N_22639,N_22558);
or U23266 (N_23266,N_22799,N_22538);
nand U23267 (N_23267,N_22653,N_22728);
nor U23268 (N_23268,N_22730,N_22616);
nand U23269 (N_23269,N_22545,N_22916);
xnor U23270 (N_23270,N_22594,N_22899);
and U23271 (N_23271,N_22991,N_22752);
nor U23272 (N_23272,N_22549,N_22579);
nor U23273 (N_23273,N_22915,N_22714);
nor U23274 (N_23274,N_22645,N_22720);
nand U23275 (N_23275,N_22739,N_22847);
nand U23276 (N_23276,N_22824,N_22737);
xor U23277 (N_23277,N_22993,N_22781);
or U23278 (N_23278,N_22863,N_22875);
nand U23279 (N_23279,N_22800,N_22851);
or U23280 (N_23280,N_22959,N_22759);
nor U23281 (N_23281,N_22656,N_22713);
and U23282 (N_23282,N_22724,N_22896);
or U23283 (N_23283,N_22767,N_22705);
xnor U23284 (N_23284,N_22605,N_22900);
and U23285 (N_23285,N_22873,N_22902);
nand U23286 (N_23286,N_22892,N_22797);
and U23287 (N_23287,N_22998,N_22938);
and U23288 (N_23288,N_22529,N_22891);
xnor U23289 (N_23289,N_22850,N_22623);
and U23290 (N_23290,N_22896,N_22795);
or U23291 (N_23291,N_22978,N_22685);
xor U23292 (N_23292,N_22814,N_22526);
and U23293 (N_23293,N_22556,N_22601);
xor U23294 (N_23294,N_22911,N_22935);
or U23295 (N_23295,N_22811,N_22984);
nor U23296 (N_23296,N_22680,N_22746);
xnor U23297 (N_23297,N_22744,N_22704);
and U23298 (N_23298,N_22989,N_22825);
xnor U23299 (N_23299,N_22706,N_22844);
and U23300 (N_23300,N_22568,N_22517);
nand U23301 (N_23301,N_22503,N_22929);
xnor U23302 (N_23302,N_22971,N_22801);
nor U23303 (N_23303,N_22873,N_22802);
and U23304 (N_23304,N_22716,N_22979);
and U23305 (N_23305,N_22780,N_22803);
and U23306 (N_23306,N_22949,N_22588);
and U23307 (N_23307,N_22679,N_22929);
nor U23308 (N_23308,N_22958,N_22615);
xor U23309 (N_23309,N_22531,N_22592);
and U23310 (N_23310,N_22964,N_22854);
or U23311 (N_23311,N_22778,N_22702);
xnor U23312 (N_23312,N_22997,N_22698);
and U23313 (N_23313,N_22967,N_22877);
nor U23314 (N_23314,N_22708,N_22653);
xor U23315 (N_23315,N_22607,N_22975);
nor U23316 (N_23316,N_22565,N_22980);
nand U23317 (N_23317,N_22664,N_22980);
xor U23318 (N_23318,N_22855,N_22794);
and U23319 (N_23319,N_22859,N_22565);
nor U23320 (N_23320,N_22884,N_22903);
and U23321 (N_23321,N_22962,N_22740);
and U23322 (N_23322,N_22875,N_22635);
and U23323 (N_23323,N_22530,N_22862);
and U23324 (N_23324,N_22796,N_22599);
and U23325 (N_23325,N_22989,N_22513);
nor U23326 (N_23326,N_22932,N_22506);
xor U23327 (N_23327,N_22738,N_22640);
nand U23328 (N_23328,N_22733,N_22571);
and U23329 (N_23329,N_22783,N_22552);
xnor U23330 (N_23330,N_22847,N_22558);
or U23331 (N_23331,N_22876,N_22847);
and U23332 (N_23332,N_22910,N_22772);
xnor U23333 (N_23333,N_22503,N_22717);
or U23334 (N_23334,N_22830,N_22623);
nand U23335 (N_23335,N_22984,N_22750);
and U23336 (N_23336,N_22655,N_22901);
xnor U23337 (N_23337,N_22781,N_22690);
nand U23338 (N_23338,N_22756,N_22553);
xnor U23339 (N_23339,N_22502,N_22656);
nor U23340 (N_23340,N_22876,N_22549);
xor U23341 (N_23341,N_22931,N_22546);
nor U23342 (N_23342,N_22682,N_22683);
nand U23343 (N_23343,N_22614,N_22947);
nor U23344 (N_23344,N_22649,N_22515);
xor U23345 (N_23345,N_22871,N_22950);
nand U23346 (N_23346,N_22706,N_22589);
xnor U23347 (N_23347,N_22836,N_22750);
and U23348 (N_23348,N_22831,N_22988);
nand U23349 (N_23349,N_22501,N_22964);
nor U23350 (N_23350,N_22738,N_22790);
xnor U23351 (N_23351,N_22884,N_22964);
nand U23352 (N_23352,N_22686,N_22893);
or U23353 (N_23353,N_22876,N_22566);
nor U23354 (N_23354,N_22972,N_22935);
xnor U23355 (N_23355,N_22618,N_22956);
nand U23356 (N_23356,N_22914,N_22535);
xnor U23357 (N_23357,N_22917,N_22772);
or U23358 (N_23358,N_22907,N_22919);
xnor U23359 (N_23359,N_22541,N_22987);
xnor U23360 (N_23360,N_22849,N_22809);
nand U23361 (N_23361,N_22964,N_22582);
xnor U23362 (N_23362,N_22902,N_22791);
nor U23363 (N_23363,N_22879,N_22773);
xor U23364 (N_23364,N_22531,N_22774);
nor U23365 (N_23365,N_22854,N_22966);
nand U23366 (N_23366,N_22800,N_22993);
nand U23367 (N_23367,N_22533,N_22701);
and U23368 (N_23368,N_22922,N_22821);
and U23369 (N_23369,N_22531,N_22875);
nor U23370 (N_23370,N_22695,N_22860);
and U23371 (N_23371,N_22625,N_22855);
xnor U23372 (N_23372,N_22957,N_22966);
nor U23373 (N_23373,N_22583,N_22533);
and U23374 (N_23374,N_22991,N_22668);
and U23375 (N_23375,N_22598,N_22930);
xnor U23376 (N_23376,N_22965,N_22533);
nand U23377 (N_23377,N_22673,N_22538);
xnor U23378 (N_23378,N_22646,N_22825);
nand U23379 (N_23379,N_22962,N_22696);
nand U23380 (N_23380,N_22873,N_22888);
xnor U23381 (N_23381,N_22571,N_22668);
and U23382 (N_23382,N_22829,N_22843);
xor U23383 (N_23383,N_22895,N_22712);
xnor U23384 (N_23384,N_22802,N_22958);
xnor U23385 (N_23385,N_22943,N_22842);
or U23386 (N_23386,N_22699,N_22803);
or U23387 (N_23387,N_22722,N_22574);
nor U23388 (N_23388,N_22863,N_22549);
xor U23389 (N_23389,N_22736,N_22981);
nor U23390 (N_23390,N_22987,N_22543);
xnor U23391 (N_23391,N_22507,N_22922);
xor U23392 (N_23392,N_22513,N_22702);
xnor U23393 (N_23393,N_22709,N_22635);
nor U23394 (N_23394,N_22575,N_22938);
and U23395 (N_23395,N_22792,N_22862);
xnor U23396 (N_23396,N_22975,N_22773);
nor U23397 (N_23397,N_22813,N_22986);
nand U23398 (N_23398,N_22602,N_22911);
and U23399 (N_23399,N_22540,N_22613);
and U23400 (N_23400,N_22905,N_22954);
nand U23401 (N_23401,N_22937,N_22944);
and U23402 (N_23402,N_22605,N_22984);
or U23403 (N_23403,N_22869,N_22998);
or U23404 (N_23404,N_22879,N_22564);
nand U23405 (N_23405,N_22681,N_22972);
and U23406 (N_23406,N_22799,N_22552);
nand U23407 (N_23407,N_22814,N_22986);
and U23408 (N_23408,N_22748,N_22721);
nor U23409 (N_23409,N_22684,N_22652);
nor U23410 (N_23410,N_22558,N_22781);
nor U23411 (N_23411,N_22520,N_22767);
and U23412 (N_23412,N_22508,N_22869);
and U23413 (N_23413,N_22518,N_22797);
xnor U23414 (N_23414,N_22650,N_22784);
nor U23415 (N_23415,N_22849,N_22598);
and U23416 (N_23416,N_22821,N_22858);
or U23417 (N_23417,N_22578,N_22685);
and U23418 (N_23418,N_22629,N_22946);
and U23419 (N_23419,N_22642,N_22626);
or U23420 (N_23420,N_22650,N_22762);
and U23421 (N_23421,N_22939,N_22703);
xnor U23422 (N_23422,N_22843,N_22620);
and U23423 (N_23423,N_22849,N_22662);
xor U23424 (N_23424,N_22595,N_22786);
xnor U23425 (N_23425,N_22637,N_22579);
nand U23426 (N_23426,N_22984,N_22892);
xor U23427 (N_23427,N_22530,N_22540);
or U23428 (N_23428,N_22907,N_22625);
and U23429 (N_23429,N_22578,N_22760);
and U23430 (N_23430,N_22862,N_22844);
xnor U23431 (N_23431,N_22652,N_22843);
and U23432 (N_23432,N_22893,N_22671);
nor U23433 (N_23433,N_22546,N_22837);
nand U23434 (N_23434,N_22836,N_22590);
nand U23435 (N_23435,N_22836,N_22802);
nor U23436 (N_23436,N_22936,N_22966);
xor U23437 (N_23437,N_22999,N_22944);
nor U23438 (N_23438,N_22946,N_22904);
nand U23439 (N_23439,N_22846,N_22936);
nand U23440 (N_23440,N_22648,N_22554);
xor U23441 (N_23441,N_22952,N_22521);
nand U23442 (N_23442,N_22617,N_22613);
nor U23443 (N_23443,N_22913,N_22950);
xnor U23444 (N_23444,N_22528,N_22509);
and U23445 (N_23445,N_22619,N_22912);
xor U23446 (N_23446,N_22772,N_22961);
and U23447 (N_23447,N_22658,N_22552);
nor U23448 (N_23448,N_22853,N_22673);
xor U23449 (N_23449,N_22763,N_22842);
and U23450 (N_23450,N_22855,N_22528);
nor U23451 (N_23451,N_22868,N_22563);
nor U23452 (N_23452,N_22562,N_22628);
xnor U23453 (N_23453,N_22825,N_22824);
nor U23454 (N_23454,N_22695,N_22567);
nand U23455 (N_23455,N_22707,N_22601);
nand U23456 (N_23456,N_22982,N_22536);
nor U23457 (N_23457,N_22567,N_22926);
nand U23458 (N_23458,N_22690,N_22880);
nor U23459 (N_23459,N_22652,N_22510);
and U23460 (N_23460,N_22964,N_22583);
nor U23461 (N_23461,N_22859,N_22541);
nand U23462 (N_23462,N_22929,N_22613);
nor U23463 (N_23463,N_22567,N_22528);
and U23464 (N_23464,N_22517,N_22910);
nand U23465 (N_23465,N_22950,N_22896);
nor U23466 (N_23466,N_22824,N_22574);
or U23467 (N_23467,N_22951,N_22772);
nor U23468 (N_23468,N_22985,N_22753);
and U23469 (N_23469,N_22866,N_22910);
nand U23470 (N_23470,N_22951,N_22836);
nor U23471 (N_23471,N_22696,N_22947);
xnor U23472 (N_23472,N_22580,N_22936);
or U23473 (N_23473,N_22672,N_22851);
or U23474 (N_23474,N_22897,N_22695);
xnor U23475 (N_23475,N_22683,N_22793);
nand U23476 (N_23476,N_22546,N_22804);
and U23477 (N_23477,N_22780,N_22617);
xnor U23478 (N_23478,N_22678,N_22823);
nand U23479 (N_23479,N_22938,N_22653);
xnor U23480 (N_23480,N_22717,N_22682);
xor U23481 (N_23481,N_22912,N_22580);
nand U23482 (N_23482,N_22587,N_22559);
nand U23483 (N_23483,N_22974,N_22602);
or U23484 (N_23484,N_22960,N_22598);
nor U23485 (N_23485,N_22779,N_22821);
nand U23486 (N_23486,N_22718,N_22701);
nand U23487 (N_23487,N_22623,N_22785);
xor U23488 (N_23488,N_22725,N_22950);
and U23489 (N_23489,N_22544,N_22768);
and U23490 (N_23490,N_22718,N_22607);
nor U23491 (N_23491,N_22605,N_22676);
nor U23492 (N_23492,N_22602,N_22735);
or U23493 (N_23493,N_22535,N_22852);
nor U23494 (N_23494,N_22840,N_22671);
xor U23495 (N_23495,N_22835,N_22786);
xor U23496 (N_23496,N_22840,N_22999);
xnor U23497 (N_23497,N_22842,N_22982);
nand U23498 (N_23498,N_22661,N_22590);
xnor U23499 (N_23499,N_22587,N_22740);
nand U23500 (N_23500,N_23219,N_23260);
nand U23501 (N_23501,N_23295,N_23247);
nor U23502 (N_23502,N_23455,N_23200);
xor U23503 (N_23503,N_23444,N_23440);
xor U23504 (N_23504,N_23363,N_23328);
nor U23505 (N_23505,N_23057,N_23016);
nand U23506 (N_23506,N_23040,N_23153);
xor U23507 (N_23507,N_23416,N_23139);
nor U23508 (N_23508,N_23182,N_23197);
and U23509 (N_23509,N_23356,N_23296);
xnor U23510 (N_23510,N_23134,N_23433);
nand U23511 (N_23511,N_23461,N_23249);
nor U23512 (N_23512,N_23316,N_23286);
or U23513 (N_23513,N_23272,N_23332);
and U23514 (N_23514,N_23143,N_23257);
or U23515 (N_23515,N_23305,N_23339);
nor U23516 (N_23516,N_23022,N_23268);
nor U23517 (N_23517,N_23209,N_23163);
and U23518 (N_23518,N_23179,N_23072);
or U23519 (N_23519,N_23469,N_23025);
or U23520 (N_23520,N_23447,N_23415);
xor U23521 (N_23521,N_23131,N_23288);
nor U23522 (N_23522,N_23147,N_23300);
nor U23523 (N_23523,N_23292,N_23207);
or U23524 (N_23524,N_23251,N_23385);
nand U23525 (N_23525,N_23477,N_23119);
or U23526 (N_23526,N_23196,N_23046);
or U23527 (N_23527,N_23488,N_23125);
xor U23528 (N_23528,N_23380,N_23329);
and U23529 (N_23529,N_23165,N_23347);
and U23530 (N_23530,N_23358,N_23301);
nand U23531 (N_23531,N_23441,N_23013);
or U23532 (N_23532,N_23388,N_23063);
and U23533 (N_23533,N_23011,N_23325);
nand U23534 (N_23534,N_23351,N_23041);
xnor U23535 (N_23535,N_23482,N_23122);
nor U23536 (N_23536,N_23135,N_23151);
xor U23537 (N_23537,N_23481,N_23269);
nor U23538 (N_23538,N_23105,N_23424);
nand U23539 (N_23539,N_23456,N_23335);
nand U23540 (N_23540,N_23451,N_23113);
nor U23541 (N_23541,N_23327,N_23344);
or U23542 (N_23542,N_23364,N_23452);
or U23543 (N_23543,N_23039,N_23343);
nor U23544 (N_23544,N_23483,N_23445);
xnor U23545 (N_23545,N_23127,N_23373);
xor U23546 (N_23546,N_23137,N_23308);
nand U23547 (N_23547,N_23045,N_23255);
xor U23548 (N_23548,N_23460,N_23394);
xor U23549 (N_23549,N_23211,N_23024);
xor U23550 (N_23550,N_23216,N_23067);
xor U23551 (N_23551,N_23058,N_23117);
nand U23552 (N_23552,N_23193,N_23104);
or U23553 (N_23553,N_23429,N_23284);
nor U23554 (N_23554,N_23029,N_23244);
or U23555 (N_23555,N_23309,N_23078);
xnor U23556 (N_23556,N_23256,N_23336);
or U23557 (N_23557,N_23318,N_23326);
nand U23558 (N_23558,N_23204,N_23449);
or U23559 (N_23559,N_23164,N_23273);
and U23560 (N_23560,N_23346,N_23087);
or U23561 (N_23561,N_23479,N_23263);
nand U23562 (N_23562,N_23369,N_23084);
nor U23563 (N_23563,N_23317,N_23160);
nand U23564 (N_23564,N_23458,N_23495);
and U23565 (N_23565,N_23166,N_23060);
nor U23566 (N_23566,N_23302,N_23224);
xnor U23567 (N_23567,N_23185,N_23108);
and U23568 (N_23568,N_23271,N_23395);
xor U23569 (N_23569,N_23354,N_23202);
nor U23570 (N_23570,N_23075,N_23048);
and U23571 (N_23571,N_23177,N_23285);
nor U23572 (N_23572,N_23463,N_23419);
nand U23573 (N_23573,N_23176,N_23133);
or U23574 (N_23574,N_23437,N_23240);
nand U23575 (N_23575,N_23487,N_23103);
or U23576 (N_23576,N_23299,N_23218);
or U23577 (N_23577,N_23368,N_23074);
nor U23578 (N_23578,N_23298,N_23290);
nor U23579 (N_23579,N_23223,N_23361);
and U23580 (N_23580,N_23337,N_23015);
nor U23581 (N_23581,N_23402,N_23068);
nand U23582 (N_23582,N_23457,N_23232);
and U23583 (N_23583,N_23413,N_23043);
and U23584 (N_23584,N_23228,N_23405);
nor U23585 (N_23585,N_23492,N_23367);
and U23586 (N_23586,N_23303,N_23222);
nor U23587 (N_23587,N_23167,N_23096);
nor U23588 (N_23588,N_23494,N_23435);
or U23589 (N_23589,N_23055,N_23348);
xnor U23590 (N_23590,N_23321,N_23235);
nor U23591 (N_23591,N_23054,N_23267);
nor U23592 (N_23592,N_23059,N_23007);
nand U23593 (N_23593,N_23009,N_23254);
and U23594 (N_23594,N_23192,N_23259);
nand U23595 (N_23595,N_23044,N_23323);
and U23596 (N_23596,N_23066,N_23396);
and U23597 (N_23597,N_23434,N_23019);
and U23598 (N_23598,N_23387,N_23370);
nand U23599 (N_23599,N_23426,N_23277);
or U23600 (N_23600,N_23042,N_23161);
nor U23601 (N_23601,N_23378,N_23004);
and U23602 (N_23602,N_23146,N_23474);
nand U23603 (N_23603,N_23093,N_23281);
or U23604 (N_23604,N_23485,N_23052);
nand U23605 (N_23605,N_23130,N_23341);
nor U23606 (N_23606,N_23003,N_23189);
xor U23607 (N_23607,N_23493,N_23028);
xnor U23608 (N_23608,N_23132,N_23198);
or U23609 (N_23609,N_23050,N_23436);
nor U23610 (N_23610,N_23203,N_23397);
and U23611 (N_23611,N_23486,N_23425);
nor U23612 (N_23612,N_23357,N_23386);
xnor U23613 (N_23613,N_23080,N_23069);
nand U23614 (N_23614,N_23377,N_23032);
xnor U23615 (N_23615,N_23391,N_23264);
nand U23616 (N_23616,N_23026,N_23338);
nand U23617 (N_23617,N_23002,N_23038);
and U23618 (N_23618,N_23466,N_23008);
or U23619 (N_23619,N_23306,N_23234);
or U23620 (N_23620,N_23014,N_23205);
nor U23621 (N_23621,N_23453,N_23421);
and U23622 (N_23622,N_23148,N_23170);
nor U23623 (N_23623,N_23324,N_23390);
xnor U23624 (N_23624,N_23000,N_23439);
and U23625 (N_23625,N_23417,N_23475);
nand U23626 (N_23626,N_23106,N_23304);
or U23627 (N_23627,N_23129,N_23178);
nand U23628 (N_23628,N_23095,N_23484);
or U23629 (N_23629,N_23409,N_23090);
nand U23630 (N_23630,N_23315,N_23027);
or U23631 (N_23631,N_23404,N_23162);
nor U23632 (N_23632,N_23006,N_23073);
nor U23633 (N_23633,N_23275,N_23330);
or U23634 (N_23634,N_23283,N_23238);
nor U23635 (N_23635,N_23490,N_23071);
or U23636 (N_23636,N_23156,N_23401);
xnor U23637 (N_23637,N_23340,N_23109);
and U23638 (N_23638,N_23012,N_23051);
nand U23639 (N_23639,N_23070,N_23410);
nor U23640 (N_23640,N_23010,N_23121);
or U23641 (N_23641,N_23467,N_23213);
nor U23642 (N_23642,N_23291,N_23406);
and U23643 (N_23643,N_23005,N_23110);
xor U23644 (N_23644,N_23053,N_23253);
nor U23645 (N_23645,N_23111,N_23077);
xor U23646 (N_23646,N_23199,N_23379);
nand U23647 (N_23647,N_23422,N_23086);
nor U23648 (N_23648,N_23365,N_23114);
or U23649 (N_23649,N_23159,N_23188);
or U23650 (N_23650,N_23226,N_23034);
and U23651 (N_23651,N_23242,N_23035);
nand U23652 (N_23652,N_23231,N_23289);
or U23653 (N_23653,N_23175,N_23374);
and U23654 (N_23654,N_23124,N_23088);
xnor U23655 (N_23655,N_23168,N_23215);
or U23656 (N_23656,N_23342,N_23123);
or U23657 (N_23657,N_23258,N_23100);
or U23658 (N_23658,N_23407,N_23400);
nand U23659 (N_23659,N_23017,N_23265);
nor U23660 (N_23660,N_23064,N_23172);
xor U23661 (N_23661,N_23261,N_23001);
xor U23662 (N_23662,N_23392,N_23237);
or U23663 (N_23663,N_23225,N_23061);
xnor U23664 (N_23664,N_23239,N_23089);
xor U23665 (N_23665,N_23297,N_23371);
or U23666 (N_23666,N_23126,N_23220);
nor U23667 (N_23667,N_23194,N_23206);
or U23668 (N_23668,N_23047,N_23366);
nor U23669 (N_23669,N_23152,N_23195);
and U23670 (N_23670,N_23241,N_23446);
and U23671 (N_23671,N_23149,N_23375);
and U23672 (N_23672,N_23428,N_23454);
nor U23673 (N_23673,N_23398,N_23118);
xnor U23674 (N_23674,N_23293,N_23140);
nor U23675 (N_23675,N_23138,N_23079);
or U23676 (N_23676,N_23036,N_23462);
nand U23677 (N_23677,N_23279,N_23217);
nor U23678 (N_23678,N_23476,N_23418);
or U23679 (N_23679,N_23432,N_23294);
nor U23680 (N_23680,N_23018,N_23393);
nor U23681 (N_23681,N_23107,N_23274);
and U23682 (N_23682,N_23154,N_23155);
nor U23683 (N_23683,N_23381,N_23062);
xnor U23684 (N_23684,N_23183,N_23158);
nand U23685 (N_23685,N_23414,N_23471);
nand U23686 (N_23686,N_23210,N_23169);
xor U23687 (N_23687,N_23049,N_23157);
nor U23688 (N_23688,N_23056,N_23334);
nor U23689 (N_23689,N_23360,N_23248);
and U23690 (N_23690,N_23101,N_23115);
xnor U23691 (N_23691,N_23276,N_23307);
nand U23692 (N_23692,N_23438,N_23423);
xor U23693 (N_23693,N_23229,N_23099);
and U23694 (N_23694,N_23144,N_23180);
xor U23695 (N_23695,N_23201,N_23319);
xor U23696 (N_23696,N_23411,N_23399);
nand U23697 (N_23697,N_23171,N_23280);
xnor U23698 (N_23698,N_23097,N_23278);
nor U23699 (N_23699,N_23450,N_23496);
and U23700 (N_23700,N_23252,N_23459);
or U23701 (N_23701,N_23312,N_23081);
xnor U23702 (N_23702,N_23065,N_23023);
and U23703 (N_23703,N_23091,N_23142);
xnor U23704 (N_23704,N_23362,N_23442);
xnor U23705 (N_23705,N_23473,N_23037);
nor U23706 (N_23706,N_23262,N_23353);
and U23707 (N_23707,N_23174,N_23314);
or U23708 (N_23708,N_23470,N_23350);
and U23709 (N_23709,N_23266,N_23345);
nand U23710 (N_23710,N_23465,N_23376);
and U23711 (N_23711,N_23372,N_23112);
xnor U23712 (N_23712,N_23233,N_23083);
or U23713 (N_23713,N_23141,N_23186);
xor U23714 (N_23714,N_23184,N_23359);
nand U23715 (N_23715,N_23214,N_23491);
and U23716 (N_23716,N_23020,N_23245);
or U23717 (N_23717,N_23383,N_23250);
nand U23718 (N_23718,N_23227,N_23150);
xor U23719 (N_23719,N_23191,N_23431);
xnor U23720 (N_23720,N_23033,N_23349);
xnor U23721 (N_23721,N_23430,N_23082);
or U23722 (N_23722,N_23489,N_23322);
nand U23723 (N_23723,N_23472,N_23331);
nor U23724 (N_23724,N_23173,N_23030);
nor U23725 (N_23725,N_23085,N_23102);
nand U23726 (N_23726,N_23094,N_23181);
and U23727 (N_23727,N_23098,N_23021);
nand U23728 (N_23728,N_23031,N_23420);
nor U23729 (N_23729,N_23145,N_23355);
nor U23730 (N_23730,N_23190,N_23136);
nand U23731 (N_23731,N_23221,N_23443);
xor U23732 (N_23732,N_23464,N_23287);
nor U23733 (N_23733,N_23403,N_23282);
nand U23734 (N_23734,N_23116,N_23270);
and U23735 (N_23735,N_23497,N_23468);
or U23736 (N_23736,N_23382,N_23352);
xnor U23737 (N_23737,N_23243,N_23499);
nand U23738 (N_23738,N_23120,N_23313);
and U23739 (N_23739,N_23128,N_23448);
or U23740 (N_23740,N_23311,N_23076);
xnor U23741 (N_23741,N_23092,N_23236);
and U23742 (N_23742,N_23478,N_23310);
and U23743 (N_23743,N_23389,N_23320);
nand U23744 (N_23744,N_23427,N_23412);
nor U23745 (N_23745,N_23384,N_23208);
xor U23746 (N_23746,N_23187,N_23246);
nor U23747 (N_23747,N_23480,N_23408);
nand U23748 (N_23748,N_23333,N_23212);
nand U23749 (N_23749,N_23498,N_23230);
xnor U23750 (N_23750,N_23011,N_23406);
nor U23751 (N_23751,N_23199,N_23371);
or U23752 (N_23752,N_23234,N_23001);
nand U23753 (N_23753,N_23320,N_23206);
or U23754 (N_23754,N_23128,N_23342);
nand U23755 (N_23755,N_23236,N_23142);
xnor U23756 (N_23756,N_23101,N_23132);
and U23757 (N_23757,N_23057,N_23153);
nor U23758 (N_23758,N_23405,N_23238);
and U23759 (N_23759,N_23078,N_23245);
xor U23760 (N_23760,N_23134,N_23486);
or U23761 (N_23761,N_23491,N_23302);
xor U23762 (N_23762,N_23246,N_23408);
or U23763 (N_23763,N_23495,N_23135);
nor U23764 (N_23764,N_23097,N_23140);
nand U23765 (N_23765,N_23046,N_23418);
and U23766 (N_23766,N_23457,N_23248);
xnor U23767 (N_23767,N_23444,N_23473);
nor U23768 (N_23768,N_23278,N_23255);
nand U23769 (N_23769,N_23097,N_23099);
nor U23770 (N_23770,N_23049,N_23192);
nand U23771 (N_23771,N_23143,N_23355);
nand U23772 (N_23772,N_23417,N_23241);
and U23773 (N_23773,N_23266,N_23328);
and U23774 (N_23774,N_23157,N_23105);
nor U23775 (N_23775,N_23471,N_23262);
nand U23776 (N_23776,N_23018,N_23419);
or U23777 (N_23777,N_23046,N_23134);
or U23778 (N_23778,N_23276,N_23490);
nor U23779 (N_23779,N_23403,N_23457);
and U23780 (N_23780,N_23118,N_23339);
nor U23781 (N_23781,N_23066,N_23445);
or U23782 (N_23782,N_23162,N_23225);
nand U23783 (N_23783,N_23453,N_23026);
xor U23784 (N_23784,N_23289,N_23492);
or U23785 (N_23785,N_23493,N_23468);
and U23786 (N_23786,N_23177,N_23362);
or U23787 (N_23787,N_23244,N_23180);
and U23788 (N_23788,N_23148,N_23344);
xor U23789 (N_23789,N_23176,N_23304);
and U23790 (N_23790,N_23223,N_23130);
nor U23791 (N_23791,N_23388,N_23312);
nor U23792 (N_23792,N_23196,N_23153);
nand U23793 (N_23793,N_23346,N_23301);
or U23794 (N_23794,N_23385,N_23493);
xor U23795 (N_23795,N_23020,N_23123);
nand U23796 (N_23796,N_23183,N_23040);
nor U23797 (N_23797,N_23017,N_23101);
nor U23798 (N_23798,N_23336,N_23112);
nor U23799 (N_23799,N_23369,N_23162);
xnor U23800 (N_23800,N_23361,N_23137);
xor U23801 (N_23801,N_23055,N_23028);
or U23802 (N_23802,N_23469,N_23312);
nand U23803 (N_23803,N_23327,N_23420);
nand U23804 (N_23804,N_23335,N_23068);
xnor U23805 (N_23805,N_23482,N_23188);
nor U23806 (N_23806,N_23154,N_23239);
nor U23807 (N_23807,N_23279,N_23164);
and U23808 (N_23808,N_23395,N_23402);
xnor U23809 (N_23809,N_23062,N_23167);
and U23810 (N_23810,N_23366,N_23068);
or U23811 (N_23811,N_23353,N_23405);
nor U23812 (N_23812,N_23459,N_23328);
nand U23813 (N_23813,N_23074,N_23310);
nand U23814 (N_23814,N_23036,N_23024);
xor U23815 (N_23815,N_23158,N_23270);
nor U23816 (N_23816,N_23053,N_23220);
and U23817 (N_23817,N_23472,N_23353);
and U23818 (N_23818,N_23260,N_23303);
nor U23819 (N_23819,N_23248,N_23024);
nand U23820 (N_23820,N_23322,N_23097);
nand U23821 (N_23821,N_23199,N_23404);
or U23822 (N_23822,N_23002,N_23422);
nor U23823 (N_23823,N_23200,N_23332);
xor U23824 (N_23824,N_23136,N_23254);
xnor U23825 (N_23825,N_23300,N_23382);
and U23826 (N_23826,N_23096,N_23240);
xnor U23827 (N_23827,N_23360,N_23400);
xnor U23828 (N_23828,N_23170,N_23041);
nand U23829 (N_23829,N_23146,N_23366);
nor U23830 (N_23830,N_23083,N_23104);
or U23831 (N_23831,N_23268,N_23299);
and U23832 (N_23832,N_23020,N_23447);
xnor U23833 (N_23833,N_23307,N_23364);
nand U23834 (N_23834,N_23178,N_23261);
and U23835 (N_23835,N_23446,N_23255);
nand U23836 (N_23836,N_23006,N_23224);
or U23837 (N_23837,N_23372,N_23133);
xnor U23838 (N_23838,N_23264,N_23082);
nand U23839 (N_23839,N_23319,N_23092);
nor U23840 (N_23840,N_23278,N_23266);
nand U23841 (N_23841,N_23138,N_23106);
xor U23842 (N_23842,N_23495,N_23463);
nor U23843 (N_23843,N_23271,N_23189);
nand U23844 (N_23844,N_23013,N_23354);
nand U23845 (N_23845,N_23402,N_23114);
nand U23846 (N_23846,N_23329,N_23287);
xor U23847 (N_23847,N_23310,N_23410);
nand U23848 (N_23848,N_23305,N_23225);
nor U23849 (N_23849,N_23224,N_23069);
nor U23850 (N_23850,N_23397,N_23274);
and U23851 (N_23851,N_23497,N_23026);
xor U23852 (N_23852,N_23078,N_23472);
or U23853 (N_23853,N_23050,N_23215);
or U23854 (N_23854,N_23247,N_23005);
and U23855 (N_23855,N_23132,N_23040);
nand U23856 (N_23856,N_23159,N_23178);
and U23857 (N_23857,N_23487,N_23305);
or U23858 (N_23858,N_23316,N_23150);
xnor U23859 (N_23859,N_23362,N_23445);
xnor U23860 (N_23860,N_23330,N_23210);
nor U23861 (N_23861,N_23248,N_23218);
and U23862 (N_23862,N_23284,N_23326);
xnor U23863 (N_23863,N_23087,N_23221);
nand U23864 (N_23864,N_23050,N_23022);
xor U23865 (N_23865,N_23277,N_23403);
nand U23866 (N_23866,N_23133,N_23259);
or U23867 (N_23867,N_23466,N_23209);
nor U23868 (N_23868,N_23249,N_23397);
xor U23869 (N_23869,N_23268,N_23208);
nor U23870 (N_23870,N_23417,N_23188);
and U23871 (N_23871,N_23434,N_23319);
and U23872 (N_23872,N_23091,N_23302);
nand U23873 (N_23873,N_23241,N_23187);
xor U23874 (N_23874,N_23439,N_23382);
or U23875 (N_23875,N_23469,N_23001);
nor U23876 (N_23876,N_23273,N_23246);
or U23877 (N_23877,N_23424,N_23492);
xor U23878 (N_23878,N_23490,N_23016);
nor U23879 (N_23879,N_23259,N_23358);
or U23880 (N_23880,N_23045,N_23180);
xnor U23881 (N_23881,N_23286,N_23192);
nand U23882 (N_23882,N_23095,N_23144);
or U23883 (N_23883,N_23479,N_23287);
and U23884 (N_23884,N_23341,N_23219);
nor U23885 (N_23885,N_23277,N_23351);
xor U23886 (N_23886,N_23460,N_23305);
nand U23887 (N_23887,N_23382,N_23226);
or U23888 (N_23888,N_23246,N_23174);
or U23889 (N_23889,N_23243,N_23087);
xnor U23890 (N_23890,N_23011,N_23026);
nand U23891 (N_23891,N_23302,N_23194);
xnor U23892 (N_23892,N_23007,N_23477);
and U23893 (N_23893,N_23174,N_23111);
nor U23894 (N_23894,N_23485,N_23412);
nor U23895 (N_23895,N_23398,N_23413);
or U23896 (N_23896,N_23305,N_23493);
and U23897 (N_23897,N_23287,N_23030);
nand U23898 (N_23898,N_23317,N_23301);
xor U23899 (N_23899,N_23151,N_23024);
nor U23900 (N_23900,N_23331,N_23132);
xor U23901 (N_23901,N_23327,N_23080);
xnor U23902 (N_23902,N_23161,N_23151);
or U23903 (N_23903,N_23383,N_23101);
nand U23904 (N_23904,N_23335,N_23428);
nor U23905 (N_23905,N_23048,N_23224);
and U23906 (N_23906,N_23270,N_23498);
and U23907 (N_23907,N_23074,N_23043);
nor U23908 (N_23908,N_23137,N_23154);
xnor U23909 (N_23909,N_23063,N_23440);
or U23910 (N_23910,N_23088,N_23275);
and U23911 (N_23911,N_23427,N_23096);
nor U23912 (N_23912,N_23215,N_23147);
xnor U23913 (N_23913,N_23116,N_23407);
nor U23914 (N_23914,N_23042,N_23017);
and U23915 (N_23915,N_23233,N_23064);
or U23916 (N_23916,N_23069,N_23378);
and U23917 (N_23917,N_23440,N_23340);
and U23918 (N_23918,N_23267,N_23463);
nand U23919 (N_23919,N_23085,N_23240);
or U23920 (N_23920,N_23334,N_23025);
and U23921 (N_23921,N_23366,N_23126);
and U23922 (N_23922,N_23239,N_23498);
and U23923 (N_23923,N_23271,N_23382);
nor U23924 (N_23924,N_23084,N_23281);
xor U23925 (N_23925,N_23474,N_23379);
nand U23926 (N_23926,N_23264,N_23431);
nand U23927 (N_23927,N_23098,N_23246);
xor U23928 (N_23928,N_23428,N_23320);
nand U23929 (N_23929,N_23482,N_23308);
nand U23930 (N_23930,N_23267,N_23037);
and U23931 (N_23931,N_23115,N_23322);
and U23932 (N_23932,N_23331,N_23104);
xor U23933 (N_23933,N_23140,N_23220);
xor U23934 (N_23934,N_23144,N_23379);
nor U23935 (N_23935,N_23053,N_23240);
xor U23936 (N_23936,N_23039,N_23017);
nor U23937 (N_23937,N_23131,N_23191);
nand U23938 (N_23938,N_23374,N_23213);
nor U23939 (N_23939,N_23337,N_23353);
xnor U23940 (N_23940,N_23447,N_23159);
nor U23941 (N_23941,N_23140,N_23180);
nor U23942 (N_23942,N_23383,N_23451);
nand U23943 (N_23943,N_23491,N_23355);
nor U23944 (N_23944,N_23435,N_23010);
and U23945 (N_23945,N_23362,N_23011);
or U23946 (N_23946,N_23030,N_23458);
xnor U23947 (N_23947,N_23153,N_23062);
or U23948 (N_23948,N_23064,N_23192);
or U23949 (N_23949,N_23351,N_23105);
or U23950 (N_23950,N_23478,N_23199);
or U23951 (N_23951,N_23219,N_23124);
xor U23952 (N_23952,N_23152,N_23361);
and U23953 (N_23953,N_23181,N_23085);
nor U23954 (N_23954,N_23331,N_23388);
nor U23955 (N_23955,N_23460,N_23129);
nor U23956 (N_23956,N_23077,N_23099);
nor U23957 (N_23957,N_23208,N_23389);
nor U23958 (N_23958,N_23192,N_23354);
or U23959 (N_23959,N_23320,N_23089);
or U23960 (N_23960,N_23278,N_23408);
nand U23961 (N_23961,N_23150,N_23289);
xor U23962 (N_23962,N_23448,N_23158);
nand U23963 (N_23963,N_23225,N_23451);
and U23964 (N_23964,N_23014,N_23493);
nand U23965 (N_23965,N_23080,N_23366);
or U23966 (N_23966,N_23197,N_23304);
nor U23967 (N_23967,N_23194,N_23319);
and U23968 (N_23968,N_23018,N_23214);
or U23969 (N_23969,N_23416,N_23108);
and U23970 (N_23970,N_23191,N_23038);
or U23971 (N_23971,N_23071,N_23039);
and U23972 (N_23972,N_23384,N_23028);
nor U23973 (N_23973,N_23139,N_23178);
and U23974 (N_23974,N_23457,N_23045);
nand U23975 (N_23975,N_23457,N_23203);
or U23976 (N_23976,N_23459,N_23057);
and U23977 (N_23977,N_23215,N_23196);
or U23978 (N_23978,N_23222,N_23039);
nand U23979 (N_23979,N_23042,N_23069);
or U23980 (N_23980,N_23010,N_23082);
and U23981 (N_23981,N_23048,N_23212);
xor U23982 (N_23982,N_23261,N_23168);
nand U23983 (N_23983,N_23211,N_23059);
or U23984 (N_23984,N_23323,N_23269);
nand U23985 (N_23985,N_23282,N_23216);
and U23986 (N_23986,N_23456,N_23388);
and U23987 (N_23987,N_23109,N_23390);
and U23988 (N_23988,N_23092,N_23252);
or U23989 (N_23989,N_23458,N_23246);
or U23990 (N_23990,N_23317,N_23247);
nand U23991 (N_23991,N_23068,N_23367);
nand U23992 (N_23992,N_23362,N_23053);
nor U23993 (N_23993,N_23383,N_23264);
nand U23994 (N_23994,N_23166,N_23010);
or U23995 (N_23995,N_23351,N_23448);
nor U23996 (N_23996,N_23483,N_23459);
and U23997 (N_23997,N_23319,N_23130);
nand U23998 (N_23998,N_23264,N_23061);
nand U23999 (N_23999,N_23031,N_23062);
xor U24000 (N_24000,N_23738,N_23817);
and U24001 (N_24001,N_23662,N_23951);
nor U24002 (N_24002,N_23607,N_23541);
nor U24003 (N_24003,N_23922,N_23698);
xor U24004 (N_24004,N_23562,N_23528);
xor U24005 (N_24005,N_23599,N_23623);
nand U24006 (N_24006,N_23737,N_23937);
or U24007 (N_24007,N_23886,N_23613);
nand U24008 (N_24008,N_23764,N_23678);
xnor U24009 (N_24009,N_23733,N_23992);
xnor U24010 (N_24010,N_23861,N_23934);
or U24011 (N_24011,N_23900,N_23622);
or U24012 (N_24012,N_23539,N_23593);
and U24013 (N_24013,N_23745,N_23959);
nor U24014 (N_24014,N_23556,N_23950);
nor U24015 (N_24015,N_23509,N_23869);
and U24016 (N_24016,N_23803,N_23611);
nand U24017 (N_24017,N_23693,N_23988);
nand U24018 (N_24018,N_23620,N_23808);
nand U24019 (N_24019,N_23520,N_23600);
and U24020 (N_24020,N_23812,N_23824);
xnor U24021 (N_24021,N_23834,N_23550);
or U24022 (N_24022,N_23547,N_23596);
and U24023 (N_24023,N_23521,N_23781);
nand U24024 (N_24024,N_23625,N_23574);
nor U24025 (N_24025,N_23619,N_23936);
nand U24026 (N_24026,N_23987,N_23962);
nand U24027 (N_24027,N_23699,N_23512);
nor U24028 (N_24028,N_23919,N_23788);
or U24029 (N_24029,N_23501,N_23872);
or U24030 (N_24030,N_23579,N_23971);
and U24031 (N_24031,N_23533,N_23702);
and U24032 (N_24032,N_23998,N_23975);
xnor U24033 (N_24033,N_23551,N_23825);
nand U24034 (N_24034,N_23649,N_23982);
nor U24035 (N_24035,N_23530,N_23567);
nor U24036 (N_24036,N_23914,N_23794);
nor U24037 (N_24037,N_23885,N_23798);
and U24038 (N_24038,N_23602,N_23514);
or U24039 (N_24039,N_23686,N_23773);
and U24040 (N_24040,N_23748,N_23744);
nor U24041 (N_24041,N_23641,N_23828);
and U24042 (N_24042,N_23797,N_23767);
or U24043 (N_24043,N_23854,N_23694);
nor U24044 (N_24044,N_23908,N_23814);
nor U24045 (N_24045,N_23902,N_23891);
or U24046 (N_24046,N_23713,N_23893);
or U24047 (N_24047,N_23983,N_23639);
nand U24048 (N_24048,N_23701,N_23672);
nand U24049 (N_24049,N_23525,N_23755);
and U24050 (N_24050,N_23832,N_23981);
or U24051 (N_24051,N_23532,N_23954);
xor U24052 (N_24052,N_23526,N_23795);
xor U24053 (N_24053,N_23608,N_23684);
nor U24054 (N_24054,N_23830,N_23665);
or U24055 (N_24055,N_23668,N_23617);
nand U24056 (N_24056,N_23732,N_23775);
xnor U24057 (N_24057,N_23636,N_23670);
and U24058 (N_24058,N_23881,N_23667);
xnor U24059 (N_24059,N_23839,N_23949);
and U24060 (N_24060,N_23647,N_23907);
xnor U24061 (N_24061,N_23663,N_23896);
nand U24062 (N_24062,N_23771,N_23978);
and U24063 (N_24063,N_23555,N_23882);
and U24064 (N_24064,N_23801,N_23840);
or U24065 (N_24065,N_23614,N_23973);
nor U24066 (N_24066,N_23860,N_23522);
xor U24067 (N_24067,N_23570,N_23586);
and U24068 (N_24068,N_23927,N_23892);
and U24069 (N_24069,N_23822,N_23612);
xor U24070 (N_24070,N_23718,N_23507);
or U24071 (N_24071,N_23787,N_23785);
nand U24072 (N_24072,N_23805,N_23709);
or U24073 (N_24073,N_23683,N_23564);
or U24074 (N_24074,N_23631,N_23849);
or U24075 (N_24075,N_23500,N_23603);
nand U24076 (N_24076,N_23553,N_23750);
or U24077 (N_24077,N_23754,N_23681);
or U24078 (N_24078,N_23585,N_23752);
nor U24079 (N_24079,N_23658,N_23594);
and U24080 (N_24080,N_23627,N_23844);
and U24081 (N_24081,N_23821,N_23848);
or U24082 (N_24082,N_23510,N_23763);
nand U24083 (N_24083,N_23565,N_23661);
nor U24084 (N_24084,N_23545,N_23901);
nor U24085 (N_24085,N_23943,N_23913);
nand U24086 (N_24086,N_23736,N_23536);
xnor U24087 (N_24087,N_23502,N_23855);
xor U24088 (N_24088,N_23866,N_23873);
or U24089 (N_24089,N_23967,N_23685);
nor U24090 (N_24090,N_23591,N_23899);
nor U24091 (N_24091,N_23909,N_23880);
or U24092 (N_24092,N_23876,N_23974);
nor U24093 (N_24093,N_23859,N_23990);
or U24094 (N_24094,N_23726,N_23540);
nand U24095 (N_24095,N_23637,N_23731);
or U24096 (N_24096,N_23888,N_23753);
nor U24097 (N_24097,N_23676,N_23843);
and U24098 (N_24098,N_23878,N_23955);
xor U24099 (N_24099,N_23942,N_23835);
or U24100 (N_24100,N_23995,N_23642);
or U24101 (N_24101,N_23823,N_23671);
nand U24102 (N_24102,N_23758,N_23944);
or U24103 (N_24103,N_23598,N_23833);
xor U24104 (N_24104,N_23654,N_23597);
nor U24105 (N_24105,N_23777,N_23711);
or U24106 (N_24106,N_23765,N_23956);
nand U24107 (N_24107,N_23710,N_23997);
nand U24108 (N_24108,N_23723,N_23985);
nor U24109 (N_24109,N_23519,N_23566);
xor U24110 (N_24110,N_23910,N_23609);
or U24111 (N_24111,N_23739,N_23704);
nand U24112 (N_24112,N_23646,N_23741);
xnor U24113 (N_24113,N_23581,N_23552);
xor U24114 (N_24114,N_23993,N_23904);
or U24115 (N_24115,N_23560,N_23791);
and U24116 (N_24116,N_23621,N_23604);
xor U24117 (N_24117,N_23692,N_23714);
nand U24118 (N_24118,N_23537,N_23707);
nand U24119 (N_24119,N_23538,N_23761);
and U24120 (N_24120,N_23728,N_23749);
nand U24121 (N_24121,N_23535,N_23583);
xnor U24122 (N_24122,N_23929,N_23920);
nand U24123 (N_24123,N_23529,N_23572);
nand U24124 (N_24124,N_23518,N_23687);
and U24125 (N_24125,N_23506,N_23800);
xor U24126 (N_24126,N_23563,N_23925);
and U24127 (N_24127,N_23953,N_23582);
xnor U24128 (N_24128,N_23911,N_23864);
nor U24129 (N_24129,N_23867,N_23923);
nand U24130 (N_24130,N_23769,N_23961);
and U24131 (N_24131,N_23846,N_23557);
or U24132 (N_24132,N_23584,N_23931);
xor U24133 (N_24133,N_23722,N_23802);
nand U24134 (N_24134,N_23595,N_23747);
xnor U24135 (N_24135,N_23703,N_23505);
nor U24136 (N_24136,N_23673,N_23708);
or U24137 (N_24137,N_23504,N_23695);
xnor U24138 (N_24138,N_23587,N_23879);
or U24139 (N_24139,N_23527,N_23578);
nand U24140 (N_24140,N_23930,N_23818);
or U24141 (N_24141,N_23716,N_23513);
nand U24142 (N_24142,N_23932,N_23523);
xnor U24143 (N_24143,N_23508,N_23674);
nor U24144 (N_24144,N_23735,N_23768);
or U24145 (N_24145,N_23660,N_23776);
nand U24146 (N_24146,N_23573,N_23980);
or U24147 (N_24147,N_23796,N_23724);
and U24148 (N_24148,N_23984,N_23601);
nor U24149 (N_24149,N_23895,N_23952);
nor U24150 (N_24150,N_23810,N_23850);
and U24151 (N_24151,N_23634,N_23780);
xor U24152 (N_24152,N_23793,N_23945);
nor U24153 (N_24153,N_23783,N_23877);
nor U24154 (N_24154,N_23657,N_23546);
nor U24155 (N_24155,N_23946,N_23542);
nor U24156 (N_24156,N_23940,N_23991);
or U24157 (N_24157,N_23589,N_23851);
xnor U24158 (N_24158,N_23916,N_23655);
and U24159 (N_24159,N_23675,N_23757);
nor U24160 (N_24160,N_23734,N_23948);
and U24161 (N_24161,N_23719,N_23697);
xnor U24162 (N_24162,N_23633,N_23503);
nor U24163 (N_24163,N_23610,N_23874);
nand U24164 (N_24164,N_23807,N_23548);
and U24165 (N_24165,N_23836,N_23778);
and U24166 (N_24166,N_23571,N_23632);
and U24167 (N_24167,N_23691,N_23845);
xor U24168 (N_24168,N_23669,N_23534);
xor U24169 (N_24169,N_23924,N_23559);
nand U24170 (N_24170,N_23715,N_23630);
nand U24171 (N_24171,N_23947,N_23590);
or U24172 (N_24172,N_23554,N_23790);
nor U24173 (N_24173,N_23838,N_23870);
or U24174 (N_24174,N_23721,N_23743);
nor U24175 (N_24175,N_23903,N_23811);
nor U24176 (N_24176,N_23815,N_23770);
nand U24177 (N_24177,N_23831,N_23645);
and U24178 (N_24178,N_23941,N_23827);
and U24179 (N_24179,N_23644,N_23696);
nor U24180 (N_24180,N_23871,N_23915);
and U24181 (N_24181,N_23543,N_23616);
nor U24182 (N_24182,N_23690,N_23759);
and U24183 (N_24183,N_23918,N_23935);
nand U24184 (N_24184,N_23926,N_23897);
nand U24185 (N_24185,N_23717,N_23651);
xor U24186 (N_24186,N_23730,N_23592);
nand U24187 (N_24187,N_23858,N_23853);
and U24188 (N_24188,N_23883,N_23705);
xor U24189 (N_24189,N_23569,N_23842);
xor U24190 (N_24190,N_23624,N_23568);
and U24191 (N_24191,N_23516,N_23826);
xor U24192 (N_24192,N_23751,N_23906);
and U24193 (N_24193,N_23628,N_23999);
and U24194 (N_24194,N_23894,N_23933);
or U24195 (N_24195,N_23544,N_23875);
nand U24196 (N_24196,N_23575,N_23618);
xor U24197 (N_24197,N_23958,N_23939);
xnor U24198 (N_24198,N_23979,N_23779);
xor U24199 (N_24199,N_23666,N_23515);
and U24200 (N_24200,N_23524,N_23577);
or U24201 (N_24201,N_23679,N_23966);
xor U24202 (N_24202,N_23890,N_23729);
xnor U24203 (N_24203,N_23680,N_23626);
and U24204 (N_24204,N_23996,N_23786);
nor U24205 (N_24205,N_23652,N_23725);
nor U24206 (N_24206,N_23756,N_23829);
or U24207 (N_24207,N_23588,N_23852);
nand U24208 (N_24208,N_23809,N_23863);
nand U24209 (N_24209,N_23580,N_23740);
xnor U24210 (N_24210,N_23766,N_23605);
and U24211 (N_24211,N_23689,N_23558);
xnor U24212 (N_24212,N_23742,N_23989);
nand U24213 (N_24213,N_23792,N_23977);
nor U24214 (N_24214,N_23917,N_23561);
nor U24215 (N_24215,N_23656,N_23746);
and U24216 (N_24216,N_23782,N_23517);
and U24217 (N_24217,N_23576,N_23712);
or U24218 (N_24218,N_23970,N_23720);
nor U24219 (N_24219,N_23847,N_23643);
nor U24220 (N_24220,N_23976,N_23606);
and U24221 (N_24221,N_23813,N_23912);
nor U24222 (N_24222,N_23772,N_23960);
or U24223 (N_24223,N_23820,N_23968);
nor U24224 (N_24224,N_23938,N_23921);
nand U24225 (N_24225,N_23841,N_23887);
xnor U24226 (N_24226,N_23898,N_23905);
and U24227 (N_24227,N_23964,N_23868);
nand U24228 (N_24228,N_23994,N_23856);
xnor U24229 (N_24229,N_23638,N_23865);
or U24230 (N_24230,N_23819,N_23664);
and U24231 (N_24231,N_23682,N_23816);
or U24232 (N_24232,N_23549,N_23889);
and U24233 (N_24233,N_23762,N_23804);
or U24234 (N_24234,N_23688,N_23972);
nor U24235 (N_24235,N_23677,N_23862);
nand U24236 (N_24236,N_23799,N_23965);
nand U24237 (N_24237,N_23957,N_23986);
nand U24238 (N_24238,N_23969,N_23648);
nand U24239 (N_24239,N_23531,N_23615);
nor U24240 (N_24240,N_23837,N_23635);
nor U24241 (N_24241,N_23784,N_23650);
or U24242 (N_24242,N_23789,N_23928);
xnor U24243 (N_24243,N_23659,N_23653);
nand U24244 (N_24244,N_23727,N_23511);
nand U24245 (N_24245,N_23963,N_23700);
nor U24246 (N_24246,N_23774,N_23706);
or U24247 (N_24247,N_23629,N_23806);
nor U24248 (N_24248,N_23857,N_23884);
and U24249 (N_24249,N_23760,N_23640);
and U24250 (N_24250,N_23633,N_23906);
xnor U24251 (N_24251,N_23594,N_23608);
and U24252 (N_24252,N_23987,N_23999);
nor U24253 (N_24253,N_23503,N_23613);
xor U24254 (N_24254,N_23825,N_23687);
and U24255 (N_24255,N_23696,N_23607);
nand U24256 (N_24256,N_23913,N_23706);
xor U24257 (N_24257,N_23852,N_23687);
nand U24258 (N_24258,N_23620,N_23869);
nor U24259 (N_24259,N_23928,N_23889);
nand U24260 (N_24260,N_23649,N_23776);
and U24261 (N_24261,N_23934,N_23856);
or U24262 (N_24262,N_23946,N_23533);
nand U24263 (N_24263,N_23836,N_23520);
nor U24264 (N_24264,N_23827,N_23978);
nand U24265 (N_24265,N_23850,N_23713);
or U24266 (N_24266,N_23526,N_23655);
or U24267 (N_24267,N_23634,N_23865);
and U24268 (N_24268,N_23949,N_23575);
nand U24269 (N_24269,N_23985,N_23789);
nand U24270 (N_24270,N_23668,N_23792);
xor U24271 (N_24271,N_23662,N_23877);
xor U24272 (N_24272,N_23638,N_23954);
nand U24273 (N_24273,N_23578,N_23526);
xnor U24274 (N_24274,N_23815,N_23614);
nand U24275 (N_24275,N_23556,N_23947);
nor U24276 (N_24276,N_23615,N_23961);
xnor U24277 (N_24277,N_23770,N_23725);
nor U24278 (N_24278,N_23823,N_23805);
xnor U24279 (N_24279,N_23899,N_23717);
or U24280 (N_24280,N_23948,N_23528);
nor U24281 (N_24281,N_23969,N_23663);
and U24282 (N_24282,N_23916,N_23968);
and U24283 (N_24283,N_23863,N_23659);
and U24284 (N_24284,N_23537,N_23932);
nor U24285 (N_24285,N_23755,N_23587);
nor U24286 (N_24286,N_23764,N_23846);
or U24287 (N_24287,N_23862,N_23757);
nand U24288 (N_24288,N_23826,N_23557);
nor U24289 (N_24289,N_23723,N_23783);
nor U24290 (N_24290,N_23840,N_23540);
nand U24291 (N_24291,N_23894,N_23948);
and U24292 (N_24292,N_23739,N_23588);
xor U24293 (N_24293,N_23839,N_23868);
nor U24294 (N_24294,N_23972,N_23762);
and U24295 (N_24295,N_23628,N_23767);
nor U24296 (N_24296,N_23893,N_23816);
nor U24297 (N_24297,N_23762,N_23770);
and U24298 (N_24298,N_23616,N_23783);
and U24299 (N_24299,N_23854,N_23579);
and U24300 (N_24300,N_23993,N_23644);
or U24301 (N_24301,N_23964,N_23719);
xor U24302 (N_24302,N_23897,N_23675);
xnor U24303 (N_24303,N_23989,N_23644);
or U24304 (N_24304,N_23913,N_23588);
or U24305 (N_24305,N_23760,N_23641);
nand U24306 (N_24306,N_23824,N_23551);
nor U24307 (N_24307,N_23651,N_23732);
nor U24308 (N_24308,N_23566,N_23501);
xor U24309 (N_24309,N_23859,N_23843);
nor U24310 (N_24310,N_23509,N_23924);
nand U24311 (N_24311,N_23865,N_23534);
nand U24312 (N_24312,N_23981,N_23512);
nand U24313 (N_24313,N_23657,N_23686);
and U24314 (N_24314,N_23597,N_23612);
nand U24315 (N_24315,N_23633,N_23822);
and U24316 (N_24316,N_23639,N_23606);
and U24317 (N_24317,N_23825,N_23978);
nor U24318 (N_24318,N_23995,N_23689);
nand U24319 (N_24319,N_23743,N_23766);
nand U24320 (N_24320,N_23578,N_23742);
nand U24321 (N_24321,N_23795,N_23650);
nor U24322 (N_24322,N_23729,N_23971);
nor U24323 (N_24323,N_23739,N_23930);
nor U24324 (N_24324,N_23795,N_23919);
or U24325 (N_24325,N_23892,N_23763);
and U24326 (N_24326,N_23891,N_23869);
and U24327 (N_24327,N_23590,N_23575);
and U24328 (N_24328,N_23831,N_23748);
xor U24329 (N_24329,N_23957,N_23704);
or U24330 (N_24330,N_23834,N_23731);
or U24331 (N_24331,N_23990,N_23615);
nand U24332 (N_24332,N_23632,N_23770);
nand U24333 (N_24333,N_23659,N_23560);
and U24334 (N_24334,N_23578,N_23899);
and U24335 (N_24335,N_23552,N_23847);
nor U24336 (N_24336,N_23844,N_23814);
xnor U24337 (N_24337,N_23742,N_23949);
and U24338 (N_24338,N_23818,N_23911);
or U24339 (N_24339,N_23716,N_23544);
or U24340 (N_24340,N_23761,N_23503);
and U24341 (N_24341,N_23625,N_23618);
nand U24342 (N_24342,N_23540,N_23702);
or U24343 (N_24343,N_23947,N_23647);
and U24344 (N_24344,N_23758,N_23628);
and U24345 (N_24345,N_23878,N_23534);
and U24346 (N_24346,N_23569,N_23575);
xor U24347 (N_24347,N_23707,N_23690);
and U24348 (N_24348,N_23839,N_23799);
xor U24349 (N_24349,N_23872,N_23802);
nand U24350 (N_24350,N_23603,N_23606);
nand U24351 (N_24351,N_23787,N_23603);
nand U24352 (N_24352,N_23948,N_23674);
nand U24353 (N_24353,N_23811,N_23519);
nor U24354 (N_24354,N_23939,N_23660);
nand U24355 (N_24355,N_23522,N_23505);
nor U24356 (N_24356,N_23730,N_23789);
nand U24357 (N_24357,N_23976,N_23543);
xor U24358 (N_24358,N_23528,N_23919);
nand U24359 (N_24359,N_23709,N_23560);
and U24360 (N_24360,N_23607,N_23805);
nand U24361 (N_24361,N_23527,N_23555);
nand U24362 (N_24362,N_23618,N_23772);
and U24363 (N_24363,N_23807,N_23731);
and U24364 (N_24364,N_23849,N_23916);
or U24365 (N_24365,N_23735,N_23945);
or U24366 (N_24366,N_23553,N_23535);
or U24367 (N_24367,N_23604,N_23711);
nor U24368 (N_24368,N_23836,N_23819);
and U24369 (N_24369,N_23841,N_23789);
nand U24370 (N_24370,N_23784,N_23888);
xnor U24371 (N_24371,N_23932,N_23762);
nor U24372 (N_24372,N_23680,N_23796);
nand U24373 (N_24373,N_23550,N_23651);
and U24374 (N_24374,N_23884,N_23951);
nand U24375 (N_24375,N_23647,N_23936);
or U24376 (N_24376,N_23836,N_23548);
or U24377 (N_24377,N_23903,N_23717);
and U24378 (N_24378,N_23872,N_23591);
nor U24379 (N_24379,N_23619,N_23766);
xnor U24380 (N_24380,N_23819,N_23740);
or U24381 (N_24381,N_23639,N_23550);
and U24382 (N_24382,N_23543,N_23889);
nor U24383 (N_24383,N_23670,N_23948);
xor U24384 (N_24384,N_23705,N_23660);
xor U24385 (N_24385,N_23967,N_23915);
xnor U24386 (N_24386,N_23649,N_23624);
and U24387 (N_24387,N_23977,N_23990);
nand U24388 (N_24388,N_23945,N_23543);
and U24389 (N_24389,N_23846,N_23889);
and U24390 (N_24390,N_23580,N_23779);
nor U24391 (N_24391,N_23988,N_23630);
and U24392 (N_24392,N_23682,N_23673);
nand U24393 (N_24393,N_23672,N_23930);
or U24394 (N_24394,N_23856,N_23773);
nor U24395 (N_24395,N_23944,N_23789);
and U24396 (N_24396,N_23980,N_23538);
and U24397 (N_24397,N_23626,N_23809);
and U24398 (N_24398,N_23823,N_23635);
and U24399 (N_24399,N_23612,N_23946);
or U24400 (N_24400,N_23968,N_23667);
nor U24401 (N_24401,N_23687,N_23582);
or U24402 (N_24402,N_23565,N_23525);
nand U24403 (N_24403,N_23548,N_23897);
or U24404 (N_24404,N_23709,N_23612);
or U24405 (N_24405,N_23903,N_23807);
xnor U24406 (N_24406,N_23500,N_23702);
and U24407 (N_24407,N_23907,N_23635);
or U24408 (N_24408,N_23943,N_23634);
xor U24409 (N_24409,N_23624,N_23841);
and U24410 (N_24410,N_23579,N_23816);
and U24411 (N_24411,N_23701,N_23974);
and U24412 (N_24412,N_23760,N_23751);
nor U24413 (N_24413,N_23944,N_23558);
or U24414 (N_24414,N_23939,N_23805);
and U24415 (N_24415,N_23603,N_23909);
nor U24416 (N_24416,N_23580,N_23978);
nand U24417 (N_24417,N_23505,N_23688);
nand U24418 (N_24418,N_23945,N_23997);
and U24419 (N_24419,N_23863,N_23917);
nor U24420 (N_24420,N_23932,N_23550);
nand U24421 (N_24421,N_23923,N_23967);
xnor U24422 (N_24422,N_23675,N_23602);
nand U24423 (N_24423,N_23973,N_23536);
xnor U24424 (N_24424,N_23681,N_23894);
nand U24425 (N_24425,N_23577,N_23585);
nor U24426 (N_24426,N_23551,N_23711);
and U24427 (N_24427,N_23573,N_23815);
and U24428 (N_24428,N_23878,N_23763);
or U24429 (N_24429,N_23630,N_23757);
xnor U24430 (N_24430,N_23766,N_23599);
xnor U24431 (N_24431,N_23739,N_23828);
xnor U24432 (N_24432,N_23782,N_23989);
nor U24433 (N_24433,N_23879,N_23924);
xor U24434 (N_24434,N_23675,N_23665);
nand U24435 (N_24435,N_23944,N_23974);
or U24436 (N_24436,N_23800,N_23744);
or U24437 (N_24437,N_23550,N_23682);
and U24438 (N_24438,N_23765,N_23552);
or U24439 (N_24439,N_23814,N_23769);
or U24440 (N_24440,N_23974,N_23585);
nand U24441 (N_24441,N_23969,N_23539);
xnor U24442 (N_24442,N_23671,N_23916);
nor U24443 (N_24443,N_23811,N_23705);
and U24444 (N_24444,N_23852,N_23874);
and U24445 (N_24445,N_23736,N_23835);
nor U24446 (N_24446,N_23522,N_23516);
nand U24447 (N_24447,N_23706,N_23739);
nand U24448 (N_24448,N_23568,N_23713);
or U24449 (N_24449,N_23809,N_23896);
or U24450 (N_24450,N_23959,N_23734);
or U24451 (N_24451,N_23956,N_23673);
or U24452 (N_24452,N_23948,N_23952);
or U24453 (N_24453,N_23980,N_23786);
and U24454 (N_24454,N_23986,N_23764);
xnor U24455 (N_24455,N_23857,N_23942);
or U24456 (N_24456,N_23546,N_23621);
or U24457 (N_24457,N_23713,N_23778);
or U24458 (N_24458,N_23860,N_23627);
and U24459 (N_24459,N_23866,N_23939);
nor U24460 (N_24460,N_23840,N_23884);
or U24461 (N_24461,N_23848,N_23962);
and U24462 (N_24462,N_23852,N_23606);
nand U24463 (N_24463,N_23565,N_23690);
xnor U24464 (N_24464,N_23612,N_23652);
or U24465 (N_24465,N_23843,N_23757);
and U24466 (N_24466,N_23518,N_23933);
nand U24467 (N_24467,N_23992,N_23572);
or U24468 (N_24468,N_23513,N_23793);
nand U24469 (N_24469,N_23992,N_23687);
xnor U24470 (N_24470,N_23870,N_23738);
xor U24471 (N_24471,N_23926,N_23871);
xor U24472 (N_24472,N_23662,N_23666);
and U24473 (N_24473,N_23847,N_23628);
xor U24474 (N_24474,N_23964,N_23524);
xor U24475 (N_24475,N_23547,N_23566);
nand U24476 (N_24476,N_23514,N_23948);
or U24477 (N_24477,N_23937,N_23547);
or U24478 (N_24478,N_23837,N_23773);
xor U24479 (N_24479,N_23864,N_23777);
xnor U24480 (N_24480,N_23803,N_23868);
xnor U24481 (N_24481,N_23501,N_23784);
xnor U24482 (N_24482,N_23894,N_23572);
and U24483 (N_24483,N_23909,N_23784);
nand U24484 (N_24484,N_23844,N_23616);
nor U24485 (N_24485,N_23860,N_23771);
nand U24486 (N_24486,N_23579,N_23917);
and U24487 (N_24487,N_23836,N_23782);
and U24488 (N_24488,N_23761,N_23690);
nor U24489 (N_24489,N_23977,N_23683);
nor U24490 (N_24490,N_23602,N_23519);
nor U24491 (N_24491,N_23885,N_23940);
nor U24492 (N_24492,N_23903,N_23714);
and U24493 (N_24493,N_23784,N_23588);
xnor U24494 (N_24494,N_23974,N_23821);
nor U24495 (N_24495,N_23728,N_23731);
or U24496 (N_24496,N_23856,N_23907);
and U24497 (N_24497,N_23660,N_23837);
nand U24498 (N_24498,N_23821,N_23667);
xnor U24499 (N_24499,N_23798,N_23984);
xor U24500 (N_24500,N_24400,N_24405);
nand U24501 (N_24501,N_24264,N_24169);
and U24502 (N_24502,N_24231,N_24419);
and U24503 (N_24503,N_24403,N_24379);
nor U24504 (N_24504,N_24470,N_24359);
or U24505 (N_24505,N_24257,N_24160);
and U24506 (N_24506,N_24077,N_24025);
or U24507 (N_24507,N_24316,N_24343);
xor U24508 (N_24508,N_24117,N_24095);
nand U24509 (N_24509,N_24336,N_24266);
nor U24510 (N_24510,N_24220,N_24023);
xor U24511 (N_24511,N_24021,N_24331);
nor U24512 (N_24512,N_24189,N_24158);
xnor U24513 (N_24513,N_24445,N_24057);
nand U24514 (N_24514,N_24097,N_24462);
nand U24515 (N_24515,N_24384,N_24273);
nand U24516 (N_24516,N_24486,N_24069);
nor U24517 (N_24517,N_24455,N_24146);
nor U24518 (N_24518,N_24232,N_24105);
nor U24519 (N_24519,N_24447,N_24079);
or U24520 (N_24520,N_24036,N_24153);
nand U24521 (N_24521,N_24110,N_24191);
xor U24522 (N_24522,N_24247,N_24482);
nor U24523 (N_24523,N_24087,N_24268);
nor U24524 (N_24524,N_24108,N_24281);
nand U24525 (N_24525,N_24055,N_24173);
and U24526 (N_24526,N_24370,N_24187);
or U24527 (N_24527,N_24054,N_24214);
and U24528 (N_24528,N_24468,N_24330);
and U24529 (N_24529,N_24272,N_24074);
and U24530 (N_24530,N_24234,N_24410);
xor U24531 (N_24531,N_24475,N_24377);
or U24532 (N_24532,N_24197,N_24490);
xnor U24533 (N_24533,N_24318,N_24329);
or U24534 (N_24534,N_24261,N_24496);
or U24535 (N_24535,N_24203,N_24114);
or U24536 (N_24536,N_24113,N_24358);
and U24537 (N_24537,N_24188,N_24128);
nor U24538 (N_24538,N_24430,N_24250);
or U24539 (N_24539,N_24306,N_24240);
or U24540 (N_24540,N_24417,N_24100);
nand U24541 (N_24541,N_24471,N_24165);
xnor U24542 (N_24542,N_24314,N_24335);
nor U24543 (N_24543,N_24199,N_24452);
xor U24544 (N_24544,N_24157,N_24138);
xnor U24545 (N_24545,N_24408,N_24388);
xor U24546 (N_24546,N_24399,N_24086);
and U24547 (N_24547,N_24008,N_24212);
and U24548 (N_24548,N_24211,N_24251);
or U24549 (N_24549,N_24466,N_24334);
and U24550 (N_24550,N_24141,N_24242);
nor U24551 (N_24551,N_24080,N_24164);
nand U24552 (N_24552,N_24044,N_24085);
nand U24553 (N_24553,N_24139,N_24378);
nor U24554 (N_24554,N_24416,N_24000);
xor U24555 (N_24555,N_24352,N_24207);
and U24556 (N_24556,N_24143,N_24256);
nor U24557 (N_24557,N_24383,N_24237);
nor U24558 (N_24558,N_24140,N_24047);
nand U24559 (N_24559,N_24245,N_24029);
or U24560 (N_24560,N_24222,N_24263);
and U24561 (N_24561,N_24346,N_24350);
or U24562 (N_24562,N_24323,N_24299);
and U24563 (N_24563,N_24348,N_24098);
nor U24564 (N_24564,N_24285,N_24166);
and U24565 (N_24565,N_24030,N_24026);
and U24566 (N_24566,N_24458,N_24046);
or U24567 (N_24567,N_24460,N_24287);
or U24568 (N_24568,N_24223,N_24103);
nor U24569 (N_24569,N_24254,N_24119);
and U24570 (N_24570,N_24106,N_24279);
nand U24571 (N_24571,N_24385,N_24180);
nand U24572 (N_24572,N_24305,N_24006);
xor U24573 (N_24573,N_24424,N_24413);
nand U24574 (N_24574,N_24294,N_24225);
nor U24575 (N_24575,N_24442,N_24371);
xnor U24576 (N_24576,N_24448,N_24121);
xor U24577 (N_24577,N_24196,N_24227);
nand U24578 (N_24578,N_24321,N_24089);
xor U24579 (N_24579,N_24412,N_24167);
nand U24580 (N_24580,N_24193,N_24120);
nand U24581 (N_24581,N_24498,N_24284);
nand U24582 (N_24582,N_24088,N_24485);
nor U24583 (N_24583,N_24319,N_24271);
xor U24584 (N_24584,N_24024,N_24332);
and U24585 (N_24585,N_24469,N_24300);
or U24586 (N_24586,N_24090,N_24355);
nor U24587 (N_24587,N_24073,N_24022);
xnor U24588 (N_24588,N_24286,N_24084);
xor U24589 (N_24589,N_24296,N_24288);
or U24590 (N_24590,N_24488,N_24328);
nor U24591 (N_24591,N_24267,N_24149);
nor U24592 (N_24592,N_24148,N_24204);
nor U24593 (N_24593,N_24182,N_24365);
nor U24594 (N_24594,N_24258,N_24465);
and U24595 (N_24595,N_24017,N_24317);
nand U24596 (N_24596,N_24239,N_24499);
or U24597 (N_24597,N_24393,N_24481);
nand U24598 (N_24598,N_24451,N_24324);
and U24599 (N_24599,N_24248,N_24392);
and U24600 (N_24600,N_24163,N_24489);
nor U24601 (N_24601,N_24102,N_24454);
and U24602 (N_24602,N_24048,N_24096);
or U24603 (N_24603,N_24368,N_24269);
xor U24604 (N_24604,N_24081,N_24243);
xor U24605 (N_24605,N_24374,N_24278);
and U24606 (N_24606,N_24168,N_24213);
or U24607 (N_24607,N_24221,N_24308);
xnor U24608 (N_24608,N_24274,N_24174);
and U24609 (N_24609,N_24463,N_24093);
and U24610 (N_24610,N_24342,N_24270);
or U24611 (N_24611,N_24443,N_24252);
or U24612 (N_24612,N_24293,N_24192);
nand U24613 (N_24613,N_24109,N_24124);
nor U24614 (N_24614,N_24453,N_24309);
nor U24615 (N_24615,N_24437,N_24493);
and U24616 (N_24616,N_24011,N_24491);
nand U24617 (N_24617,N_24438,N_24362);
and U24618 (N_24618,N_24397,N_24134);
xor U24619 (N_24619,N_24372,N_24421);
or U24620 (N_24620,N_24420,N_24238);
xor U24621 (N_24621,N_24115,N_24262);
and U24622 (N_24622,N_24357,N_24402);
or U24623 (N_24623,N_24156,N_24292);
nand U24624 (N_24624,N_24078,N_24492);
xor U24625 (N_24625,N_24450,N_24477);
xnor U24626 (N_24626,N_24112,N_24052);
or U24627 (N_24627,N_24367,N_24154);
xor U24628 (N_24628,N_24133,N_24027);
or U24629 (N_24629,N_24071,N_24322);
nand U24630 (N_24630,N_24068,N_24127);
or U24631 (N_24631,N_24354,N_24390);
xnor U24632 (N_24632,N_24431,N_24122);
xnor U24633 (N_24633,N_24325,N_24018);
or U24634 (N_24634,N_24484,N_24219);
xnor U24635 (N_24635,N_24064,N_24014);
xnor U24636 (N_24636,N_24444,N_24019);
and U24637 (N_24637,N_24373,N_24012);
nand U24638 (N_24638,N_24401,N_24260);
xnor U24639 (N_24639,N_24209,N_24161);
nor U24640 (N_24640,N_24456,N_24001);
nand U24641 (N_24641,N_24495,N_24175);
nor U24642 (N_24642,N_24144,N_24094);
xor U24643 (N_24643,N_24072,N_24341);
and U24644 (N_24644,N_24476,N_24404);
nand U24645 (N_24645,N_24389,N_24111);
and U24646 (N_24646,N_24432,N_24497);
or U24647 (N_24647,N_24249,N_24283);
nand U24648 (N_24648,N_24344,N_24228);
xnor U24649 (N_24649,N_24061,N_24013);
nor U24650 (N_24650,N_24190,N_24244);
and U24651 (N_24651,N_24473,N_24201);
nor U24652 (N_24652,N_24135,N_24433);
and U24653 (N_24653,N_24230,N_24171);
and U24654 (N_24654,N_24391,N_24131);
nor U24655 (N_24655,N_24015,N_24226);
and U24656 (N_24656,N_24179,N_24007);
nor U24657 (N_24657,N_24418,N_24126);
xor U24658 (N_24658,N_24041,N_24236);
or U24659 (N_24659,N_24277,N_24406);
or U24660 (N_24660,N_24099,N_24422);
xor U24661 (N_24661,N_24241,N_24033);
or U24662 (N_24662,N_24035,N_24298);
nor U24663 (N_24663,N_24337,N_24062);
xnor U24664 (N_24664,N_24415,N_24224);
nand U24665 (N_24665,N_24186,N_24202);
or U24666 (N_24666,N_24150,N_24155);
xor U24667 (N_24667,N_24461,N_24053);
xnor U24668 (N_24668,N_24028,N_24200);
and U24669 (N_24669,N_24347,N_24132);
or U24670 (N_24670,N_24031,N_24137);
and U24671 (N_24671,N_24435,N_24066);
nor U24672 (N_24672,N_24198,N_24386);
nand U24673 (N_24673,N_24206,N_24107);
or U24674 (N_24674,N_24280,N_24315);
and U24675 (N_24675,N_24446,N_24356);
nand U24676 (N_24676,N_24310,N_24276);
nand U24677 (N_24677,N_24483,N_24297);
xor U24678 (N_24678,N_24304,N_24208);
and U24679 (N_24679,N_24003,N_24345);
nor U24680 (N_24680,N_24255,N_24349);
or U24681 (N_24681,N_24375,N_24170);
and U24682 (N_24682,N_24301,N_24233);
nand U24683 (N_24683,N_24147,N_24009);
xnor U24684 (N_24684,N_24395,N_24065);
nand U24685 (N_24685,N_24032,N_24058);
nand U24686 (N_24686,N_24177,N_24381);
nand U24687 (N_24687,N_24480,N_24459);
nand U24688 (N_24688,N_24494,N_24016);
and U24689 (N_24689,N_24259,N_24313);
nor U24690 (N_24690,N_24123,N_24326);
nand U24691 (N_24691,N_24380,N_24194);
and U24692 (N_24692,N_24423,N_24142);
xor U24693 (N_24693,N_24136,N_24464);
xor U24694 (N_24694,N_24091,N_24195);
and U24695 (N_24695,N_24210,N_24361);
nor U24696 (N_24696,N_24070,N_24116);
nand U24697 (N_24697,N_24067,N_24040);
or U24698 (N_24698,N_24411,N_24457);
nor U24699 (N_24699,N_24449,N_24229);
nor U24700 (N_24700,N_24472,N_24409);
or U24701 (N_24701,N_24216,N_24183);
or U24702 (N_24702,N_24075,N_24479);
nand U24703 (N_24703,N_24056,N_24275);
or U24704 (N_24704,N_24104,N_24327);
and U24705 (N_24705,N_24043,N_24205);
and U24706 (N_24706,N_24414,N_24152);
or U24707 (N_24707,N_24050,N_24217);
and U24708 (N_24708,N_24289,N_24151);
nand U24709 (N_24709,N_24076,N_24426);
and U24710 (N_24710,N_24282,N_24474);
or U24711 (N_24711,N_24020,N_24427);
nand U24712 (N_24712,N_24092,N_24396);
nand U24713 (N_24713,N_24290,N_24176);
nand U24714 (N_24714,N_24407,N_24037);
and U24715 (N_24715,N_24311,N_24178);
nand U24716 (N_24716,N_24339,N_24353);
xor U24717 (N_24717,N_24059,N_24394);
nand U24718 (N_24718,N_24185,N_24436);
or U24719 (N_24719,N_24382,N_24082);
and U24720 (N_24720,N_24366,N_24184);
or U24721 (N_24721,N_24441,N_24295);
or U24722 (N_24722,N_24351,N_24049);
or U24723 (N_24723,N_24364,N_24478);
or U24724 (N_24724,N_24434,N_24291);
and U24725 (N_24725,N_24387,N_24303);
or U24726 (N_24726,N_24440,N_24130);
nand U24727 (N_24727,N_24083,N_24034);
and U24728 (N_24728,N_24235,N_24312);
xor U24729 (N_24729,N_24218,N_24125);
or U24730 (N_24730,N_24363,N_24340);
nor U24731 (N_24731,N_24467,N_24253);
and U24732 (N_24732,N_24101,N_24005);
nand U24733 (N_24733,N_24172,N_24246);
and U24734 (N_24734,N_24045,N_24063);
xnor U24735 (N_24735,N_24215,N_24039);
or U24736 (N_24736,N_24428,N_24425);
and U24737 (N_24737,N_24038,N_24002);
nand U24738 (N_24738,N_24320,N_24162);
xor U24739 (N_24739,N_24338,N_24060);
nand U24740 (N_24740,N_24360,N_24145);
xor U24741 (N_24741,N_24042,N_24051);
and U24742 (N_24742,N_24265,N_24129);
xor U24743 (N_24743,N_24369,N_24439);
nor U24744 (N_24744,N_24333,N_24159);
or U24745 (N_24745,N_24429,N_24010);
nor U24746 (N_24746,N_24376,N_24004);
or U24747 (N_24747,N_24487,N_24307);
and U24748 (N_24748,N_24302,N_24181);
nor U24749 (N_24749,N_24118,N_24398);
or U24750 (N_24750,N_24148,N_24000);
xnor U24751 (N_24751,N_24128,N_24139);
or U24752 (N_24752,N_24197,N_24186);
nand U24753 (N_24753,N_24260,N_24343);
nor U24754 (N_24754,N_24193,N_24260);
xnor U24755 (N_24755,N_24048,N_24417);
xnor U24756 (N_24756,N_24059,N_24357);
and U24757 (N_24757,N_24447,N_24113);
xnor U24758 (N_24758,N_24309,N_24022);
or U24759 (N_24759,N_24174,N_24138);
nand U24760 (N_24760,N_24341,N_24016);
xor U24761 (N_24761,N_24420,N_24342);
xor U24762 (N_24762,N_24477,N_24145);
xor U24763 (N_24763,N_24333,N_24470);
or U24764 (N_24764,N_24491,N_24223);
or U24765 (N_24765,N_24048,N_24253);
nand U24766 (N_24766,N_24135,N_24322);
and U24767 (N_24767,N_24417,N_24273);
nor U24768 (N_24768,N_24199,N_24497);
nor U24769 (N_24769,N_24383,N_24310);
or U24770 (N_24770,N_24063,N_24186);
and U24771 (N_24771,N_24027,N_24092);
and U24772 (N_24772,N_24051,N_24096);
nor U24773 (N_24773,N_24390,N_24196);
and U24774 (N_24774,N_24122,N_24140);
xor U24775 (N_24775,N_24372,N_24198);
xnor U24776 (N_24776,N_24422,N_24005);
or U24777 (N_24777,N_24137,N_24343);
nand U24778 (N_24778,N_24008,N_24448);
nor U24779 (N_24779,N_24241,N_24308);
or U24780 (N_24780,N_24300,N_24255);
nor U24781 (N_24781,N_24414,N_24437);
and U24782 (N_24782,N_24284,N_24061);
xnor U24783 (N_24783,N_24386,N_24067);
nor U24784 (N_24784,N_24351,N_24341);
or U24785 (N_24785,N_24266,N_24118);
nand U24786 (N_24786,N_24037,N_24464);
or U24787 (N_24787,N_24277,N_24032);
nor U24788 (N_24788,N_24247,N_24180);
or U24789 (N_24789,N_24062,N_24010);
xor U24790 (N_24790,N_24148,N_24073);
nor U24791 (N_24791,N_24475,N_24497);
nand U24792 (N_24792,N_24437,N_24488);
or U24793 (N_24793,N_24031,N_24489);
nand U24794 (N_24794,N_24182,N_24061);
or U24795 (N_24795,N_24254,N_24251);
nand U24796 (N_24796,N_24457,N_24186);
or U24797 (N_24797,N_24174,N_24461);
xnor U24798 (N_24798,N_24415,N_24400);
xnor U24799 (N_24799,N_24221,N_24100);
nand U24800 (N_24800,N_24385,N_24275);
nand U24801 (N_24801,N_24342,N_24410);
nand U24802 (N_24802,N_24041,N_24126);
xor U24803 (N_24803,N_24323,N_24038);
nand U24804 (N_24804,N_24017,N_24370);
xnor U24805 (N_24805,N_24437,N_24398);
xor U24806 (N_24806,N_24058,N_24262);
or U24807 (N_24807,N_24108,N_24251);
xnor U24808 (N_24808,N_24364,N_24489);
or U24809 (N_24809,N_24448,N_24441);
nor U24810 (N_24810,N_24254,N_24157);
nand U24811 (N_24811,N_24264,N_24208);
nor U24812 (N_24812,N_24251,N_24146);
xnor U24813 (N_24813,N_24095,N_24297);
nor U24814 (N_24814,N_24031,N_24309);
nor U24815 (N_24815,N_24220,N_24463);
or U24816 (N_24816,N_24484,N_24151);
xnor U24817 (N_24817,N_24181,N_24119);
or U24818 (N_24818,N_24178,N_24023);
nand U24819 (N_24819,N_24187,N_24403);
nand U24820 (N_24820,N_24340,N_24157);
xor U24821 (N_24821,N_24104,N_24052);
nor U24822 (N_24822,N_24114,N_24474);
xnor U24823 (N_24823,N_24093,N_24388);
xor U24824 (N_24824,N_24170,N_24376);
nor U24825 (N_24825,N_24098,N_24271);
or U24826 (N_24826,N_24092,N_24450);
nor U24827 (N_24827,N_24480,N_24140);
nor U24828 (N_24828,N_24410,N_24301);
and U24829 (N_24829,N_24297,N_24050);
nand U24830 (N_24830,N_24184,N_24062);
nor U24831 (N_24831,N_24097,N_24160);
nand U24832 (N_24832,N_24220,N_24105);
nor U24833 (N_24833,N_24248,N_24476);
and U24834 (N_24834,N_24380,N_24065);
nand U24835 (N_24835,N_24041,N_24185);
or U24836 (N_24836,N_24475,N_24343);
nor U24837 (N_24837,N_24157,N_24133);
or U24838 (N_24838,N_24363,N_24076);
and U24839 (N_24839,N_24384,N_24228);
or U24840 (N_24840,N_24300,N_24239);
xor U24841 (N_24841,N_24271,N_24303);
and U24842 (N_24842,N_24408,N_24385);
nand U24843 (N_24843,N_24481,N_24386);
or U24844 (N_24844,N_24098,N_24131);
nand U24845 (N_24845,N_24326,N_24418);
or U24846 (N_24846,N_24385,N_24071);
xnor U24847 (N_24847,N_24361,N_24018);
or U24848 (N_24848,N_24166,N_24220);
nor U24849 (N_24849,N_24484,N_24108);
nor U24850 (N_24850,N_24457,N_24388);
xor U24851 (N_24851,N_24111,N_24464);
xnor U24852 (N_24852,N_24253,N_24088);
and U24853 (N_24853,N_24055,N_24086);
nor U24854 (N_24854,N_24060,N_24021);
and U24855 (N_24855,N_24225,N_24224);
nand U24856 (N_24856,N_24173,N_24491);
and U24857 (N_24857,N_24312,N_24409);
and U24858 (N_24858,N_24385,N_24244);
nand U24859 (N_24859,N_24176,N_24283);
nand U24860 (N_24860,N_24439,N_24467);
and U24861 (N_24861,N_24193,N_24066);
nor U24862 (N_24862,N_24158,N_24412);
nand U24863 (N_24863,N_24003,N_24016);
and U24864 (N_24864,N_24270,N_24185);
xnor U24865 (N_24865,N_24305,N_24115);
or U24866 (N_24866,N_24286,N_24318);
xnor U24867 (N_24867,N_24303,N_24483);
xnor U24868 (N_24868,N_24398,N_24007);
or U24869 (N_24869,N_24348,N_24287);
nor U24870 (N_24870,N_24111,N_24359);
xnor U24871 (N_24871,N_24365,N_24019);
or U24872 (N_24872,N_24060,N_24262);
nand U24873 (N_24873,N_24009,N_24050);
nand U24874 (N_24874,N_24479,N_24205);
or U24875 (N_24875,N_24396,N_24196);
nand U24876 (N_24876,N_24109,N_24388);
or U24877 (N_24877,N_24039,N_24181);
and U24878 (N_24878,N_24294,N_24075);
or U24879 (N_24879,N_24405,N_24131);
xor U24880 (N_24880,N_24374,N_24332);
or U24881 (N_24881,N_24031,N_24486);
or U24882 (N_24882,N_24252,N_24010);
nand U24883 (N_24883,N_24146,N_24378);
xnor U24884 (N_24884,N_24164,N_24242);
or U24885 (N_24885,N_24375,N_24000);
and U24886 (N_24886,N_24493,N_24177);
xor U24887 (N_24887,N_24000,N_24107);
and U24888 (N_24888,N_24100,N_24088);
nor U24889 (N_24889,N_24484,N_24123);
nor U24890 (N_24890,N_24161,N_24094);
or U24891 (N_24891,N_24215,N_24412);
nor U24892 (N_24892,N_24347,N_24280);
nor U24893 (N_24893,N_24398,N_24257);
nand U24894 (N_24894,N_24227,N_24435);
or U24895 (N_24895,N_24141,N_24115);
nand U24896 (N_24896,N_24221,N_24282);
and U24897 (N_24897,N_24011,N_24476);
xnor U24898 (N_24898,N_24412,N_24003);
nand U24899 (N_24899,N_24340,N_24074);
xnor U24900 (N_24900,N_24379,N_24417);
nor U24901 (N_24901,N_24393,N_24396);
or U24902 (N_24902,N_24344,N_24198);
nor U24903 (N_24903,N_24247,N_24077);
xor U24904 (N_24904,N_24339,N_24298);
xor U24905 (N_24905,N_24235,N_24381);
nand U24906 (N_24906,N_24091,N_24407);
nand U24907 (N_24907,N_24163,N_24061);
xnor U24908 (N_24908,N_24016,N_24173);
and U24909 (N_24909,N_24303,N_24221);
nor U24910 (N_24910,N_24237,N_24123);
nor U24911 (N_24911,N_24145,N_24065);
and U24912 (N_24912,N_24468,N_24150);
or U24913 (N_24913,N_24011,N_24204);
or U24914 (N_24914,N_24459,N_24407);
and U24915 (N_24915,N_24326,N_24436);
nor U24916 (N_24916,N_24383,N_24495);
xor U24917 (N_24917,N_24303,N_24226);
or U24918 (N_24918,N_24047,N_24022);
or U24919 (N_24919,N_24142,N_24211);
or U24920 (N_24920,N_24355,N_24208);
and U24921 (N_24921,N_24229,N_24011);
and U24922 (N_24922,N_24007,N_24462);
or U24923 (N_24923,N_24241,N_24223);
xor U24924 (N_24924,N_24396,N_24115);
or U24925 (N_24925,N_24028,N_24085);
and U24926 (N_24926,N_24153,N_24037);
nor U24927 (N_24927,N_24341,N_24091);
xnor U24928 (N_24928,N_24018,N_24181);
or U24929 (N_24929,N_24428,N_24186);
xor U24930 (N_24930,N_24045,N_24211);
or U24931 (N_24931,N_24011,N_24114);
and U24932 (N_24932,N_24469,N_24019);
xor U24933 (N_24933,N_24155,N_24312);
xnor U24934 (N_24934,N_24019,N_24205);
or U24935 (N_24935,N_24183,N_24315);
xor U24936 (N_24936,N_24082,N_24412);
nand U24937 (N_24937,N_24204,N_24410);
xnor U24938 (N_24938,N_24329,N_24362);
nand U24939 (N_24939,N_24410,N_24250);
or U24940 (N_24940,N_24132,N_24325);
or U24941 (N_24941,N_24429,N_24417);
nor U24942 (N_24942,N_24025,N_24005);
xnor U24943 (N_24943,N_24310,N_24152);
nor U24944 (N_24944,N_24000,N_24342);
nor U24945 (N_24945,N_24125,N_24343);
or U24946 (N_24946,N_24458,N_24204);
nand U24947 (N_24947,N_24009,N_24199);
nand U24948 (N_24948,N_24298,N_24077);
xnor U24949 (N_24949,N_24420,N_24278);
and U24950 (N_24950,N_24455,N_24155);
and U24951 (N_24951,N_24425,N_24034);
or U24952 (N_24952,N_24247,N_24494);
and U24953 (N_24953,N_24086,N_24474);
nand U24954 (N_24954,N_24250,N_24358);
nor U24955 (N_24955,N_24100,N_24022);
nand U24956 (N_24956,N_24331,N_24257);
xor U24957 (N_24957,N_24455,N_24246);
and U24958 (N_24958,N_24263,N_24485);
or U24959 (N_24959,N_24491,N_24293);
nor U24960 (N_24960,N_24311,N_24125);
and U24961 (N_24961,N_24024,N_24027);
and U24962 (N_24962,N_24472,N_24252);
nand U24963 (N_24963,N_24333,N_24303);
or U24964 (N_24964,N_24413,N_24114);
nand U24965 (N_24965,N_24445,N_24021);
or U24966 (N_24966,N_24461,N_24493);
xor U24967 (N_24967,N_24100,N_24105);
and U24968 (N_24968,N_24034,N_24061);
nor U24969 (N_24969,N_24085,N_24052);
nand U24970 (N_24970,N_24457,N_24005);
nand U24971 (N_24971,N_24145,N_24175);
nor U24972 (N_24972,N_24091,N_24270);
nand U24973 (N_24973,N_24237,N_24433);
xnor U24974 (N_24974,N_24375,N_24087);
and U24975 (N_24975,N_24372,N_24374);
xor U24976 (N_24976,N_24478,N_24240);
xor U24977 (N_24977,N_24391,N_24106);
or U24978 (N_24978,N_24402,N_24270);
and U24979 (N_24979,N_24406,N_24271);
or U24980 (N_24980,N_24064,N_24291);
or U24981 (N_24981,N_24378,N_24320);
and U24982 (N_24982,N_24177,N_24208);
nand U24983 (N_24983,N_24164,N_24005);
xnor U24984 (N_24984,N_24155,N_24198);
xnor U24985 (N_24985,N_24063,N_24136);
or U24986 (N_24986,N_24374,N_24269);
or U24987 (N_24987,N_24252,N_24379);
or U24988 (N_24988,N_24119,N_24071);
nor U24989 (N_24989,N_24042,N_24412);
nor U24990 (N_24990,N_24304,N_24396);
xor U24991 (N_24991,N_24300,N_24361);
or U24992 (N_24992,N_24041,N_24474);
nand U24993 (N_24993,N_24367,N_24043);
nor U24994 (N_24994,N_24385,N_24478);
xnor U24995 (N_24995,N_24462,N_24168);
and U24996 (N_24996,N_24253,N_24016);
or U24997 (N_24997,N_24091,N_24293);
xnor U24998 (N_24998,N_24009,N_24151);
or U24999 (N_24999,N_24462,N_24484);
and U25000 (N_25000,N_24785,N_24811);
and U25001 (N_25001,N_24911,N_24578);
xnor U25002 (N_25002,N_24673,N_24694);
nand U25003 (N_25003,N_24991,N_24532);
and U25004 (N_25004,N_24516,N_24667);
or U25005 (N_25005,N_24640,N_24549);
and U25006 (N_25006,N_24876,N_24965);
or U25007 (N_25007,N_24548,N_24792);
or U25008 (N_25008,N_24599,N_24700);
and U25009 (N_25009,N_24797,N_24939);
nor U25010 (N_25010,N_24908,N_24937);
and U25011 (N_25011,N_24736,N_24696);
xnor U25012 (N_25012,N_24952,N_24517);
xor U25013 (N_25013,N_24955,N_24594);
nand U25014 (N_25014,N_24621,N_24553);
or U25015 (N_25015,N_24951,N_24721);
and U25016 (N_25016,N_24885,N_24649);
nand U25017 (N_25017,N_24817,N_24916);
nor U25018 (N_25018,N_24897,N_24718);
or U25019 (N_25019,N_24632,N_24777);
or U25020 (N_25020,N_24628,N_24539);
nand U25021 (N_25021,N_24675,N_24813);
nor U25022 (N_25022,N_24859,N_24926);
nor U25023 (N_25023,N_24783,N_24996);
and U25024 (N_25024,N_24821,N_24850);
and U25025 (N_25025,N_24636,N_24544);
or U25026 (N_25026,N_24642,N_24808);
nand U25027 (N_25027,N_24525,N_24619);
nor U25028 (N_25028,N_24954,N_24587);
or U25029 (N_25029,N_24904,N_24737);
nor U25030 (N_25030,N_24887,N_24551);
nor U25031 (N_25031,N_24570,N_24661);
nor U25032 (N_25032,N_24603,N_24614);
xnor U25033 (N_25033,N_24778,N_24574);
nor U25034 (N_25034,N_24670,N_24917);
xnor U25035 (N_25035,N_24716,N_24583);
nand U25036 (N_25036,N_24947,N_24930);
nor U25037 (N_25037,N_24689,N_24746);
or U25038 (N_25038,N_24923,N_24616);
nand U25039 (N_25039,N_24999,N_24511);
and U25040 (N_25040,N_24710,N_24961);
xnor U25041 (N_25041,N_24527,N_24862);
xor U25042 (N_25042,N_24901,N_24963);
nand U25043 (N_25043,N_24510,N_24837);
nor U25044 (N_25044,N_24514,N_24982);
xnor U25045 (N_25045,N_24757,N_24974);
and U25046 (N_25046,N_24891,N_24547);
nand U25047 (N_25047,N_24801,N_24712);
nor U25048 (N_25048,N_24683,N_24541);
xnor U25049 (N_25049,N_24713,N_24682);
and U25050 (N_25050,N_24892,N_24919);
or U25051 (N_25051,N_24877,N_24602);
nand U25052 (N_25052,N_24627,N_24723);
nand U25053 (N_25053,N_24826,N_24848);
xor U25054 (N_25054,N_24755,N_24520);
xor U25055 (N_25055,N_24781,N_24833);
nor U25056 (N_25056,N_24652,N_24905);
and U25057 (N_25057,N_24526,N_24918);
nor U25058 (N_25058,N_24935,N_24625);
and U25059 (N_25059,N_24898,N_24793);
nand U25060 (N_25060,N_24788,N_24528);
and U25061 (N_25061,N_24535,N_24856);
xor U25062 (N_25062,N_24577,N_24735);
nand U25063 (N_25063,N_24998,N_24690);
or U25064 (N_25064,N_24804,N_24537);
nor U25065 (N_25065,N_24717,N_24914);
or U25066 (N_25066,N_24769,N_24827);
or U25067 (N_25067,N_24842,N_24758);
nand U25068 (N_25068,N_24748,N_24749);
or U25069 (N_25069,N_24796,N_24960);
nand U25070 (N_25070,N_24997,N_24868);
nor U25071 (N_25071,N_24623,N_24802);
xnor U25072 (N_25072,N_24524,N_24641);
and U25073 (N_25073,N_24610,N_24882);
or U25074 (N_25074,N_24595,N_24656);
and U25075 (N_25075,N_24840,N_24671);
or U25076 (N_25076,N_24681,N_24626);
and U25077 (N_25077,N_24567,N_24503);
and U25078 (N_25078,N_24988,N_24776);
nor U25079 (N_25079,N_24835,N_24795);
and U25080 (N_25080,N_24576,N_24825);
or U25081 (N_25081,N_24958,N_24596);
or U25082 (N_25082,N_24953,N_24771);
nor U25083 (N_25083,N_24699,N_24558);
nand U25084 (N_25084,N_24845,N_24880);
or U25085 (N_25085,N_24775,N_24743);
or U25086 (N_25086,N_24809,N_24676);
nand U25087 (N_25087,N_24608,N_24924);
nor U25088 (N_25088,N_24709,N_24729);
and U25089 (N_25089,N_24762,N_24851);
nand U25090 (N_25090,N_24976,N_24853);
nor U25091 (N_25091,N_24873,N_24508);
or U25092 (N_25092,N_24669,N_24798);
nor U25093 (N_25093,N_24829,N_24580);
or U25094 (N_25094,N_24507,N_24606);
nor U25095 (N_25095,N_24715,N_24545);
nand U25096 (N_25096,N_24767,N_24692);
nand U25097 (N_25097,N_24838,N_24753);
and U25098 (N_25098,N_24546,N_24770);
nand U25099 (N_25099,N_24994,N_24772);
and U25100 (N_25100,N_24515,N_24579);
or U25101 (N_25101,N_24995,N_24847);
or U25102 (N_25102,N_24931,N_24766);
nand U25103 (N_25103,N_24942,N_24852);
nor U25104 (N_25104,N_24707,N_24720);
nand U25105 (N_25105,N_24512,N_24807);
nor U25106 (N_25106,N_24615,N_24938);
xnor U25107 (N_25107,N_24899,N_24645);
nor U25108 (N_25108,N_24861,N_24624);
nand U25109 (N_25109,N_24752,N_24653);
and U25110 (N_25110,N_24724,N_24674);
xnor U25111 (N_25111,N_24754,N_24611);
nand U25112 (N_25112,N_24725,N_24571);
and U25113 (N_25113,N_24701,N_24869);
or U25114 (N_25114,N_24784,N_24871);
nor U25115 (N_25115,N_24613,N_24909);
nand U25116 (N_25116,N_24824,N_24890);
or U25117 (N_25117,N_24945,N_24739);
nor U25118 (N_25118,N_24895,N_24894);
or U25119 (N_25119,N_24992,N_24730);
nor U25120 (N_25120,N_24839,N_24866);
nor U25121 (N_25121,N_24686,N_24538);
nand U25122 (N_25122,N_24605,N_24647);
and U25123 (N_25123,N_24933,N_24618);
nand U25124 (N_25124,N_24944,N_24819);
nand U25125 (N_25125,N_24896,N_24820);
xnor U25126 (N_25126,N_24949,N_24832);
nor U25127 (N_25127,N_24780,N_24865);
nor U25128 (N_25128,N_24860,N_24672);
nand U25129 (N_25129,N_24666,N_24874);
and U25130 (N_25130,N_24588,N_24969);
nor U25131 (N_25131,N_24657,N_24530);
nand U25132 (N_25132,N_24932,N_24759);
xor U25133 (N_25133,N_24983,N_24872);
xor U25134 (N_25134,N_24989,N_24814);
xnor U25135 (N_25135,N_24658,N_24663);
xor U25136 (N_25136,N_24774,N_24654);
and U25137 (N_25137,N_24646,N_24855);
xor U25138 (N_25138,N_24986,N_24593);
and U25139 (N_25139,N_24846,N_24831);
and U25140 (N_25140,N_24810,N_24591);
nor U25141 (N_25141,N_24505,N_24822);
nand U25142 (N_25142,N_24893,N_24590);
and U25143 (N_25143,N_24849,N_24834);
xnor U25144 (N_25144,N_24633,N_24706);
xor U25145 (N_25145,N_24702,N_24863);
xor U25146 (N_25146,N_24695,N_24643);
xor U25147 (N_25147,N_24765,N_24815);
and U25148 (N_25148,N_24883,N_24962);
and U25149 (N_25149,N_24987,N_24568);
or U25150 (N_25150,N_24773,N_24751);
xnor U25151 (N_25151,N_24662,N_24907);
nand U25152 (N_25152,N_24823,N_24604);
nor U25153 (N_25153,N_24742,N_24540);
xor U25154 (N_25154,N_24943,N_24557);
nand U25155 (N_25155,N_24782,N_24727);
nand U25156 (N_25156,N_24794,N_24858);
or U25157 (N_25157,N_24513,N_24950);
nand U25158 (N_25158,N_24738,N_24879);
nor U25159 (N_25159,N_24878,N_24745);
nand U25160 (N_25160,N_24889,N_24806);
nand U25161 (N_25161,N_24504,N_24529);
nor U25162 (N_25162,N_24660,N_24592);
and U25163 (N_25163,N_24726,N_24564);
xor U25164 (N_25164,N_24925,N_24678);
nor U25165 (N_25165,N_24597,N_24728);
nor U25166 (N_25166,N_24586,N_24854);
or U25167 (N_25167,N_24900,N_24964);
nor U25168 (N_25168,N_24502,N_24668);
nand U25169 (N_25169,N_24764,N_24830);
nor U25170 (N_25170,N_24521,N_24687);
xor U25171 (N_25171,N_24648,N_24799);
xnor U25172 (N_25172,N_24867,N_24518);
xnor U25173 (N_25173,N_24556,N_24978);
xor U25174 (N_25174,N_24857,N_24966);
nand U25175 (N_25175,N_24722,N_24920);
or U25176 (N_25176,N_24875,N_24970);
or U25177 (N_25177,N_24812,N_24573);
and U25178 (N_25178,N_24816,N_24934);
nor U25179 (N_25179,N_24786,N_24985);
nor U25180 (N_25180,N_24688,N_24651);
xnor U25181 (N_25181,N_24828,N_24554);
nand U25182 (N_25182,N_24971,N_24693);
and U25183 (N_25183,N_24644,N_24552);
or U25184 (N_25184,N_24630,N_24768);
nor U25185 (N_25185,N_24993,N_24650);
and U25186 (N_25186,N_24569,N_24956);
and U25187 (N_25187,N_24582,N_24921);
nor U25188 (N_25188,N_24881,N_24679);
and U25189 (N_25189,N_24601,N_24732);
nor U25190 (N_25190,N_24779,N_24731);
and U25191 (N_25191,N_24543,N_24967);
nand U25192 (N_25192,N_24763,N_24888);
nand U25193 (N_25193,N_24789,N_24634);
or U25194 (N_25194,N_24929,N_24697);
xor U25195 (N_25195,N_24536,N_24609);
nand U25196 (N_25196,N_24928,N_24844);
and U25197 (N_25197,N_24760,N_24550);
or U25198 (N_25198,N_24665,N_24680);
xor U25199 (N_25199,N_24622,N_24719);
nand U25200 (N_25200,N_24744,N_24977);
nand U25201 (N_25201,N_24585,N_24531);
nand U25202 (N_25202,N_24941,N_24704);
nor U25203 (N_25203,N_24589,N_24555);
and U25204 (N_25204,N_24581,N_24620);
xor U25205 (N_25205,N_24836,N_24957);
nand U25206 (N_25206,N_24980,N_24635);
nor U25207 (N_25207,N_24708,N_24703);
nand U25208 (N_25208,N_24803,N_24714);
nor U25209 (N_25209,N_24685,N_24990);
or U25210 (N_25210,N_24740,N_24747);
nand U25211 (N_25211,N_24790,N_24981);
and U25212 (N_25212,N_24638,N_24684);
or U25213 (N_25213,N_24902,N_24572);
xor U25214 (N_25214,N_24913,N_24559);
xnor U25215 (N_25215,N_24607,N_24973);
and U25216 (N_25216,N_24968,N_24959);
or U25217 (N_25217,N_24912,N_24979);
nand U25218 (N_25218,N_24805,N_24677);
nand U25219 (N_25219,N_24584,N_24659);
or U25220 (N_25220,N_24506,N_24927);
xnor U25221 (N_25221,N_24922,N_24519);
nor U25222 (N_25222,N_24761,N_24906);
xor U25223 (N_25223,N_24734,N_24629);
xnor U25224 (N_25224,N_24903,N_24561);
and U25225 (N_25225,N_24522,N_24617);
or U25226 (N_25226,N_24940,N_24533);
or U25227 (N_25227,N_24560,N_24639);
and U25228 (N_25228,N_24631,N_24946);
and U25229 (N_25229,N_24637,N_24500);
and U25230 (N_25230,N_24542,N_24698);
or U25231 (N_25231,N_24534,N_24756);
nand U25232 (N_25232,N_24972,N_24501);
and U25233 (N_25233,N_24886,N_24818);
or U25234 (N_25234,N_24870,N_24787);
nor U25235 (N_25235,N_24563,N_24509);
nand U25236 (N_25236,N_24750,N_24733);
nand U25237 (N_25237,N_24655,N_24691);
nor U25238 (N_25238,N_24711,N_24948);
xnor U25239 (N_25239,N_24800,N_24741);
and U25240 (N_25240,N_24841,N_24612);
xor U25241 (N_25241,N_24864,N_24562);
and U25242 (N_25242,N_24910,N_24600);
xor U25243 (N_25243,N_24566,N_24936);
xor U25244 (N_25244,N_24523,N_24598);
nand U25245 (N_25245,N_24565,N_24664);
or U25246 (N_25246,N_24705,N_24915);
nor U25247 (N_25247,N_24975,N_24791);
nand U25248 (N_25248,N_24843,N_24575);
or U25249 (N_25249,N_24984,N_24884);
nand U25250 (N_25250,N_24975,N_24532);
nor U25251 (N_25251,N_24965,N_24955);
xor U25252 (N_25252,N_24787,N_24576);
and U25253 (N_25253,N_24863,N_24561);
or U25254 (N_25254,N_24990,N_24554);
xor U25255 (N_25255,N_24661,N_24827);
nor U25256 (N_25256,N_24511,N_24827);
nand U25257 (N_25257,N_24982,N_24763);
and U25258 (N_25258,N_24959,N_24859);
nand U25259 (N_25259,N_24889,N_24787);
or U25260 (N_25260,N_24690,N_24701);
xor U25261 (N_25261,N_24750,N_24842);
xor U25262 (N_25262,N_24934,N_24755);
or U25263 (N_25263,N_24628,N_24738);
nor U25264 (N_25264,N_24584,N_24856);
nand U25265 (N_25265,N_24824,N_24539);
xnor U25266 (N_25266,N_24642,N_24950);
xnor U25267 (N_25267,N_24608,N_24659);
nand U25268 (N_25268,N_24966,N_24968);
xnor U25269 (N_25269,N_24805,N_24640);
nand U25270 (N_25270,N_24511,N_24962);
or U25271 (N_25271,N_24599,N_24838);
and U25272 (N_25272,N_24862,N_24670);
and U25273 (N_25273,N_24928,N_24949);
nand U25274 (N_25274,N_24988,N_24658);
nand U25275 (N_25275,N_24740,N_24977);
nor U25276 (N_25276,N_24926,N_24881);
nor U25277 (N_25277,N_24720,N_24716);
nor U25278 (N_25278,N_24724,N_24965);
nor U25279 (N_25279,N_24874,N_24599);
or U25280 (N_25280,N_24664,N_24761);
xor U25281 (N_25281,N_24824,N_24653);
or U25282 (N_25282,N_24567,N_24559);
xor U25283 (N_25283,N_24860,N_24758);
and U25284 (N_25284,N_24921,N_24524);
or U25285 (N_25285,N_24571,N_24946);
or U25286 (N_25286,N_24765,N_24574);
nor U25287 (N_25287,N_24807,N_24781);
xnor U25288 (N_25288,N_24977,N_24657);
xor U25289 (N_25289,N_24934,N_24968);
nor U25290 (N_25290,N_24999,N_24555);
xnor U25291 (N_25291,N_24538,N_24732);
or U25292 (N_25292,N_24737,N_24648);
nand U25293 (N_25293,N_24519,N_24777);
nor U25294 (N_25294,N_24661,N_24992);
or U25295 (N_25295,N_24962,N_24932);
and U25296 (N_25296,N_24602,N_24578);
xor U25297 (N_25297,N_24649,N_24937);
nor U25298 (N_25298,N_24892,N_24519);
nor U25299 (N_25299,N_24839,N_24564);
and U25300 (N_25300,N_24764,N_24801);
xnor U25301 (N_25301,N_24754,N_24875);
or U25302 (N_25302,N_24694,N_24840);
nor U25303 (N_25303,N_24822,N_24538);
or U25304 (N_25304,N_24569,N_24736);
nor U25305 (N_25305,N_24866,N_24728);
or U25306 (N_25306,N_24508,N_24938);
or U25307 (N_25307,N_24709,N_24897);
and U25308 (N_25308,N_24577,N_24660);
and U25309 (N_25309,N_24808,N_24721);
and U25310 (N_25310,N_24990,N_24907);
nand U25311 (N_25311,N_24572,N_24893);
and U25312 (N_25312,N_24707,N_24695);
or U25313 (N_25313,N_24897,N_24908);
or U25314 (N_25314,N_24553,N_24765);
nor U25315 (N_25315,N_24860,N_24646);
or U25316 (N_25316,N_24669,N_24696);
nor U25317 (N_25317,N_24839,N_24812);
xnor U25318 (N_25318,N_24866,N_24582);
nand U25319 (N_25319,N_24571,N_24867);
and U25320 (N_25320,N_24758,N_24519);
xnor U25321 (N_25321,N_24902,N_24640);
nor U25322 (N_25322,N_24529,N_24749);
or U25323 (N_25323,N_24966,N_24626);
xor U25324 (N_25324,N_24726,N_24712);
and U25325 (N_25325,N_24918,N_24926);
nor U25326 (N_25326,N_24982,N_24630);
nor U25327 (N_25327,N_24712,N_24785);
or U25328 (N_25328,N_24594,N_24687);
nor U25329 (N_25329,N_24557,N_24607);
xnor U25330 (N_25330,N_24519,N_24664);
nand U25331 (N_25331,N_24848,N_24527);
xor U25332 (N_25332,N_24633,N_24896);
and U25333 (N_25333,N_24631,N_24624);
and U25334 (N_25334,N_24705,N_24914);
and U25335 (N_25335,N_24918,N_24717);
nor U25336 (N_25336,N_24955,N_24603);
nand U25337 (N_25337,N_24679,N_24931);
or U25338 (N_25338,N_24692,N_24561);
and U25339 (N_25339,N_24629,N_24758);
nor U25340 (N_25340,N_24864,N_24614);
nand U25341 (N_25341,N_24918,N_24871);
nand U25342 (N_25342,N_24655,N_24683);
xor U25343 (N_25343,N_24918,N_24544);
nand U25344 (N_25344,N_24808,N_24616);
nor U25345 (N_25345,N_24941,N_24701);
nand U25346 (N_25346,N_24711,N_24763);
nor U25347 (N_25347,N_24919,N_24874);
or U25348 (N_25348,N_24596,N_24780);
and U25349 (N_25349,N_24805,N_24582);
xor U25350 (N_25350,N_24555,N_24710);
and U25351 (N_25351,N_24865,N_24814);
xnor U25352 (N_25352,N_24866,N_24967);
nor U25353 (N_25353,N_24907,N_24721);
and U25354 (N_25354,N_24641,N_24920);
nor U25355 (N_25355,N_24546,N_24525);
or U25356 (N_25356,N_24954,N_24870);
and U25357 (N_25357,N_24683,N_24705);
and U25358 (N_25358,N_24562,N_24985);
nand U25359 (N_25359,N_24689,N_24624);
xor U25360 (N_25360,N_24523,N_24845);
xor U25361 (N_25361,N_24771,N_24920);
and U25362 (N_25362,N_24679,N_24742);
xnor U25363 (N_25363,N_24585,N_24771);
nor U25364 (N_25364,N_24812,N_24755);
nor U25365 (N_25365,N_24720,N_24575);
nand U25366 (N_25366,N_24889,N_24721);
nor U25367 (N_25367,N_24771,N_24717);
or U25368 (N_25368,N_24780,N_24831);
and U25369 (N_25369,N_24741,N_24852);
nand U25370 (N_25370,N_24902,N_24511);
or U25371 (N_25371,N_24853,N_24508);
and U25372 (N_25372,N_24845,N_24908);
nor U25373 (N_25373,N_24544,N_24910);
and U25374 (N_25374,N_24620,N_24779);
or U25375 (N_25375,N_24820,N_24634);
nand U25376 (N_25376,N_24659,N_24620);
nor U25377 (N_25377,N_24787,N_24674);
nor U25378 (N_25378,N_24764,N_24802);
nand U25379 (N_25379,N_24944,N_24710);
nor U25380 (N_25380,N_24737,N_24684);
xnor U25381 (N_25381,N_24864,N_24902);
nor U25382 (N_25382,N_24857,N_24603);
nand U25383 (N_25383,N_24676,N_24889);
nand U25384 (N_25384,N_24613,N_24892);
or U25385 (N_25385,N_24527,N_24815);
xor U25386 (N_25386,N_24912,N_24621);
xnor U25387 (N_25387,N_24888,N_24646);
or U25388 (N_25388,N_24819,N_24773);
xor U25389 (N_25389,N_24715,N_24769);
nor U25390 (N_25390,N_24755,N_24913);
nand U25391 (N_25391,N_24682,N_24743);
and U25392 (N_25392,N_24720,N_24753);
nand U25393 (N_25393,N_24597,N_24712);
nor U25394 (N_25394,N_24720,N_24747);
and U25395 (N_25395,N_24852,N_24668);
or U25396 (N_25396,N_24521,N_24957);
or U25397 (N_25397,N_24698,N_24945);
nor U25398 (N_25398,N_24787,N_24693);
xnor U25399 (N_25399,N_24547,N_24996);
xnor U25400 (N_25400,N_24867,N_24660);
and U25401 (N_25401,N_24973,N_24762);
or U25402 (N_25402,N_24835,N_24893);
and U25403 (N_25403,N_24814,N_24963);
nand U25404 (N_25404,N_24710,N_24741);
nand U25405 (N_25405,N_24803,N_24723);
and U25406 (N_25406,N_24576,N_24898);
and U25407 (N_25407,N_24647,N_24528);
or U25408 (N_25408,N_24545,N_24953);
and U25409 (N_25409,N_24785,N_24927);
nand U25410 (N_25410,N_24744,N_24645);
and U25411 (N_25411,N_24552,N_24558);
and U25412 (N_25412,N_24914,N_24984);
nand U25413 (N_25413,N_24613,N_24914);
nand U25414 (N_25414,N_24823,N_24905);
and U25415 (N_25415,N_24677,N_24914);
nor U25416 (N_25416,N_24587,N_24891);
or U25417 (N_25417,N_24849,N_24974);
or U25418 (N_25418,N_24639,N_24860);
xnor U25419 (N_25419,N_24793,N_24685);
or U25420 (N_25420,N_24936,N_24661);
xor U25421 (N_25421,N_24764,N_24522);
xor U25422 (N_25422,N_24655,N_24908);
and U25423 (N_25423,N_24873,N_24682);
and U25424 (N_25424,N_24724,N_24559);
or U25425 (N_25425,N_24535,N_24969);
nand U25426 (N_25426,N_24604,N_24856);
nor U25427 (N_25427,N_24512,N_24531);
nand U25428 (N_25428,N_24660,N_24757);
nand U25429 (N_25429,N_24930,N_24944);
nand U25430 (N_25430,N_24532,N_24843);
or U25431 (N_25431,N_24966,N_24520);
xnor U25432 (N_25432,N_24583,N_24835);
and U25433 (N_25433,N_24990,N_24926);
and U25434 (N_25434,N_24705,N_24950);
xnor U25435 (N_25435,N_24688,N_24679);
xnor U25436 (N_25436,N_24610,N_24697);
or U25437 (N_25437,N_24844,N_24791);
and U25438 (N_25438,N_24628,N_24682);
xor U25439 (N_25439,N_24548,N_24830);
or U25440 (N_25440,N_24642,N_24526);
and U25441 (N_25441,N_24990,N_24510);
nor U25442 (N_25442,N_24697,N_24770);
nand U25443 (N_25443,N_24871,N_24611);
nor U25444 (N_25444,N_24851,N_24809);
nor U25445 (N_25445,N_24753,N_24992);
and U25446 (N_25446,N_24549,N_24996);
nor U25447 (N_25447,N_24886,N_24650);
xor U25448 (N_25448,N_24885,N_24625);
or U25449 (N_25449,N_24974,N_24508);
nor U25450 (N_25450,N_24984,N_24873);
or U25451 (N_25451,N_24641,N_24826);
nand U25452 (N_25452,N_24537,N_24512);
or U25453 (N_25453,N_24981,N_24749);
xnor U25454 (N_25454,N_24610,N_24928);
or U25455 (N_25455,N_24941,N_24968);
and U25456 (N_25456,N_24843,N_24570);
nand U25457 (N_25457,N_24560,N_24997);
nand U25458 (N_25458,N_24940,N_24929);
and U25459 (N_25459,N_24954,N_24781);
xnor U25460 (N_25460,N_24800,N_24634);
and U25461 (N_25461,N_24978,N_24877);
xnor U25462 (N_25462,N_24817,N_24904);
nor U25463 (N_25463,N_24908,N_24516);
and U25464 (N_25464,N_24969,N_24878);
nand U25465 (N_25465,N_24620,N_24770);
or U25466 (N_25466,N_24817,N_24940);
or U25467 (N_25467,N_24981,N_24999);
nand U25468 (N_25468,N_24802,N_24714);
and U25469 (N_25469,N_24913,N_24573);
nand U25470 (N_25470,N_24581,N_24560);
xor U25471 (N_25471,N_24859,N_24605);
nand U25472 (N_25472,N_24858,N_24671);
xnor U25473 (N_25473,N_24930,N_24646);
or U25474 (N_25474,N_24947,N_24586);
nand U25475 (N_25475,N_24819,N_24562);
nand U25476 (N_25476,N_24647,N_24949);
nand U25477 (N_25477,N_24571,N_24548);
nand U25478 (N_25478,N_24823,N_24642);
nand U25479 (N_25479,N_24625,N_24581);
nand U25480 (N_25480,N_24567,N_24797);
nor U25481 (N_25481,N_24607,N_24959);
xor U25482 (N_25482,N_24915,N_24967);
and U25483 (N_25483,N_24561,N_24992);
and U25484 (N_25484,N_24534,N_24721);
or U25485 (N_25485,N_24530,N_24774);
nor U25486 (N_25486,N_24895,N_24786);
or U25487 (N_25487,N_24780,N_24611);
nand U25488 (N_25488,N_24859,N_24764);
xor U25489 (N_25489,N_24749,N_24855);
or U25490 (N_25490,N_24713,N_24642);
nand U25491 (N_25491,N_24978,N_24532);
xnor U25492 (N_25492,N_24690,N_24833);
and U25493 (N_25493,N_24711,N_24828);
and U25494 (N_25494,N_24641,N_24530);
xnor U25495 (N_25495,N_24788,N_24589);
or U25496 (N_25496,N_24734,N_24631);
and U25497 (N_25497,N_24531,N_24757);
nor U25498 (N_25498,N_24694,N_24585);
nand U25499 (N_25499,N_24894,N_24795);
nor U25500 (N_25500,N_25494,N_25011);
and U25501 (N_25501,N_25418,N_25099);
and U25502 (N_25502,N_25284,N_25301);
nand U25503 (N_25503,N_25277,N_25161);
xor U25504 (N_25504,N_25241,N_25168);
nor U25505 (N_25505,N_25475,N_25405);
and U25506 (N_25506,N_25134,N_25028);
xor U25507 (N_25507,N_25497,N_25047);
nand U25508 (N_25508,N_25156,N_25376);
nand U25509 (N_25509,N_25281,N_25345);
xnor U25510 (N_25510,N_25231,N_25216);
or U25511 (N_25511,N_25226,N_25076);
nand U25512 (N_25512,N_25178,N_25157);
and U25513 (N_25513,N_25308,N_25370);
xor U25514 (N_25514,N_25015,N_25430);
and U25515 (N_25515,N_25489,N_25233);
nor U25516 (N_25516,N_25184,N_25062);
xnor U25517 (N_25517,N_25374,N_25278);
nand U25518 (N_25518,N_25142,N_25371);
or U25519 (N_25519,N_25442,N_25427);
or U25520 (N_25520,N_25154,N_25411);
nor U25521 (N_25521,N_25103,N_25252);
nand U25522 (N_25522,N_25219,N_25486);
nand U25523 (N_25523,N_25038,N_25004);
or U25524 (N_25524,N_25434,N_25147);
or U25525 (N_25525,N_25443,N_25144);
nor U25526 (N_25526,N_25106,N_25111);
nand U25527 (N_25527,N_25132,N_25385);
nor U25528 (N_25528,N_25209,N_25212);
xnor U25529 (N_25529,N_25478,N_25139);
nand U25530 (N_25530,N_25173,N_25265);
nor U25531 (N_25531,N_25090,N_25325);
and U25532 (N_25532,N_25008,N_25328);
nand U25533 (N_25533,N_25449,N_25229);
xnor U25534 (N_25534,N_25210,N_25181);
and U25535 (N_25535,N_25203,N_25254);
and U25536 (N_25536,N_25477,N_25125);
xor U25537 (N_25537,N_25448,N_25179);
nand U25538 (N_25538,N_25051,N_25109);
and U25539 (N_25539,N_25373,N_25034);
xnor U25540 (N_25540,N_25159,N_25259);
or U25541 (N_25541,N_25469,N_25270);
nor U25542 (N_25542,N_25010,N_25042);
and U25543 (N_25543,N_25414,N_25018);
or U25544 (N_25544,N_25030,N_25117);
xor U25545 (N_25545,N_25045,N_25316);
nor U25546 (N_25546,N_25176,N_25289);
nor U25547 (N_25547,N_25432,N_25061);
nor U25548 (N_25548,N_25399,N_25349);
and U25549 (N_25549,N_25452,N_25266);
xor U25550 (N_25550,N_25150,N_25146);
and U25551 (N_25551,N_25148,N_25221);
or U25552 (N_25552,N_25271,N_25243);
and U25553 (N_25553,N_25391,N_25075);
nand U25554 (N_25554,N_25499,N_25367);
nand U25555 (N_25555,N_25086,N_25394);
nor U25556 (N_25556,N_25364,N_25165);
nor U25557 (N_25557,N_25121,N_25407);
nor U25558 (N_25558,N_25361,N_25329);
or U25559 (N_25559,N_25072,N_25446);
and U25560 (N_25560,N_25114,N_25175);
nor U25561 (N_25561,N_25459,N_25136);
or U25562 (N_25562,N_25151,N_25110);
or U25563 (N_25563,N_25353,N_25298);
nor U25564 (N_25564,N_25077,N_25380);
or U25565 (N_25565,N_25048,N_25493);
or U25566 (N_25566,N_25050,N_25081);
and U25567 (N_25567,N_25365,N_25273);
nor U25568 (N_25568,N_25122,N_25052);
and U25569 (N_25569,N_25300,N_25333);
xnor U25570 (N_25570,N_25247,N_25182);
nand U25571 (N_25571,N_25059,N_25388);
and U25572 (N_25572,N_25098,N_25332);
or U25573 (N_25573,N_25423,N_25055);
xor U25574 (N_25574,N_25401,N_25234);
and U25575 (N_25575,N_25064,N_25304);
nand U25576 (N_25576,N_25029,N_25196);
and U25577 (N_25577,N_25009,N_25433);
or U25578 (N_25578,N_25400,N_25381);
nor U25579 (N_25579,N_25261,N_25007);
nand U25580 (N_25580,N_25354,N_25303);
and U25581 (N_25581,N_25260,N_25063);
xnor U25582 (N_25582,N_25360,N_25180);
nand U25583 (N_25583,N_25438,N_25451);
nand U25584 (N_25584,N_25412,N_25492);
or U25585 (N_25585,N_25250,N_25293);
xnor U25586 (N_25586,N_25172,N_25108);
xnor U25587 (N_25587,N_25246,N_25338);
xor U25588 (N_25588,N_25352,N_25205);
xor U25589 (N_25589,N_25272,N_25197);
and U25590 (N_25590,N_25436,N_25145);
and U25591 (N_25591,N_25129,N_25235);
and U25592 (N_25592,N_25428,N_25395);
nand U25593 (N_25593,N_25363,N_25074);
nor U25594 (N_25594,N_25208,N_25291);
nor U25595 (N_25595,N_25054,N_25041);
xor U25596 (N_25596,N_25190,N_25100);
and U25597 (N_25597,N_25276,N_25022);
nand U25598 (N_25598,N_25222,N_25128);
and U25599 (N_25599,N_25162,N_25027);
xor U25600 (N_25600,N_25236,N_25105);
and U25601 (N_25601,N_25457,N_25375);
and U25602 (N_25602,N_25366,N_25044);
xor U25603 (N_25603,N_25014,N_25126);
xnor U25604 (N_25604,N_25138,N_25140);
and U25605 (N_25605,N_25116,N_25039);
nand U25606 (N_25606,N_25384,N_25262);
or U25607 (N_25607,N_25113,N_25461);
nand U25608 (N_25608,N_25101,N_25248);
xor U25609 (N_25609,N_25169,N_25368);
xor U25610 (N_25610,N_25033,N_25115);
nor U25611 (N_25611,N_25214,N_25285);
nand U25612 (N_25612,N_25013,N_25420);
or U25613 (N_25613,N_25192,N_25194);
and U25614 (N_25614,N_25068,N_25288);
or U25615 (N_25615,N_25141,N_25143);
or U25616 (N_25616,N_25080,N_25408);
xnor U25617 (N_25617,N_25085,N_25417);
xor U25618 (N_25618,N_25253,N_25357);
or U25619 (N_25619,N_25347,N_25065);
and U25620 (N_25620,N_25046,N_25403);
nand U25621 (N_25621,N_25267,N_25379);
and U25622 (N_25622,N_25326,N_25387);
nor U25623 (N_25623,N_25318,N_25232);
nor U25624 (N_25624,N_25133,N_25153);
xnor U25625 (N_25625,N_25239,N_25372);
and U25626 (N_25626,N_25305,N_25482);
or U25627 (N_25627,N_25204,N_25450);
and U25628 (N_25628,N_25066,N_25470);
or U25629 (N_25629,N_25263,N_25067);
and U25630 (N_25630,N_25498,N_25421);
or U25631 (N_25631,N_25218,N_25369);
or U25632 (N_25632,N_25257,N_25415);
nand U25633 (N_25633,N_25280,N_25104);
and U25634 (N_25634,N_25224,N_25017);
and U25635 (N_25635,N_25317,N_25206);
xnor U25636 (N_25636,N_25458,N_25484);
or U25637 (N_25637,N_25220,N_25053);
nor U25638 (N_25638,N_25036,N_25392);
nor U25639 (N_25639,N_25227,N_25118);
nand U25640 (N_25640,N_25269,N_25426);
nand U25641 (N_25641,N_25057,N_25035);
and U25642 (N_25642,N_25188,N_25312);
nor U25643 (N_25643,N_25472,N_25336);
and U25644 (N_25644,N_25406,N_25092);
xor U25645 (N_25645,N_25230,N_25495);
nor U25646 (N_25646,N_25127,N_25023);
nand U25647 (N_25647,N_25348,N_25012);
nor U25648 (N_25648,N_25283,N_25225);
nand U25649 (N_25649,N_25211,N_25016);
or U25650 (N_25650,N_25350,N_25464);
nand U25651 (N_25651,N_25321,N_25485);
nand U25652 (N_25652,N_25341,N_25213);
nand U25653 (N_25653,N_25286,N_25037);
nand U25654 (N_25654,N_25342,N_25158);
or U25655 (N_25655,N_25191,N_25093);
nand U25656 (N_25656,N_25130,N_25073);
nand U25657 (N_25657,N_25382,N_25335);
or U25658 (N_25658,N_25199,N_25240);
nor U25659 (N_25659,N_25299,N_25202);
and U25660 (N_25660,N_25195,N_25327);
xor U25661 (N_25661,N_25290,N_25019);
or U25662 (N_25662,N_25390,N_25362);
xnor U25663 (N_25663,N_25445,N_25307);
xor U25664 (N_25664,N_25334,N_25160);
and U25665 (N_25665,N_25454,N_25473);
or U25666 (N_25666,N_25091,N_25083);
and U25667 (N_25667,N_25003,N_25024);
nor U25668 (N_25668,N_25337,N_25389);
nand U25669 (N_25669,N_25201,N_25331);
or U25670 (N_25670,N_25359,N_25386);
nand U25671 (N_25671,N_25095,N_25274);
and U25672 (N_25672,N_25149,N_25324);
nor U25673 (N_25673,N_25152,N_25483);
nand U25674 (N_25674,N_25437,N_25119);
xor U25675 (N_25675,N_25481,N_25185);
nand U25676 (N_25676,N_25397,N_25413);
nand U25677 (N_25677,N_25096,N_25319);
and U25678 (N_25678,N_25167,N_25163);
nand U25679 (N_25679,N_25058,N_25460);
or U25680 (N_25680,N_25404,N_25088);
nor U25681 (N_25681,N_25295,N_25135);
xor U25682 (N_25682,N_25242,N_25431);
xor U25683 (N_25683,N_25292,N_25463);
and U25684 (N_25684,N_25006,N_25409);
xnor U25685 (N_25685,N_25444,N_25238);
and U25686 (N_25686,N_25021,N_25453);
nand U25687 (N_25687,N_25177,N_25071);
and U25688 (N_25688,N_25056,N_25294);
or U25689 (N_25689,N_25049,N_25425);
or U25690 (N_25690,N_25087,N_25466);
xnor U25691 (N_25691,N_25383,N_25309);
or U25692 (N_25692,N_25001,N_25025);
nand U25693 (N_25693,N_25060,N_25496);
nand U25694 (N_25694,N_25200,N_25000);
nand U25695 (N_25695,N_25429,N_25410);
or U25696 (N_25696,N_25440,N_25102);
or U25697 (N_25697,N_25296,N_25323);
and U25698 (N_25698,N_25124,N_25170);
or U25699 (N_25699,N_25237,N_25097);
and U25700 (N_25700,N_25002,N_25120);
nor U25701 (N_25701,N_25287,N_25164);
and U25702 (N_25702,N_25439,N_25356);
and U25703 (N_25703,N_25166,N_25302);
or U25704 (N_25704,N_25084,N_25079);
or U25705 (N_25705,N_25031,N_25189);
or U25706 (N_25706,N_25320,N_25215);
nand U25707 (N_25707,N_25488,N_25487);
or U25708 (N_25708,N_25174,N_25020);
and U25709 (N_25709,N_25402,N_25217);
and U25710 (N_25710,N_25297,N_25416);
and U25711 (N_25711,N_25310,N_25339);
and U25712 (N_25712,N_25223,N_25183);
or U25713 (N_25713,N_25476,N_25491);
or U25714 (N_25714,N_25468,N_25358);
nor U25715 (N_25715,N_25490,N_25343);
or U25716 (N_25716,N_25279,N_25255);
nand U25717 (N_25717,N_25131,N_25474);
and U25718 (N_25718,N_25465,N_25377);
or U25719 (N_25719,N_25314,N_25123);
and U25720 (N_25720,N_25193,N_25424);
xor U25721 (N_25721,N_25393,N_25275);
nor U25722 (N_25722,N_25351,N_25089);
xnor U25723 (N_25723,N_25112,N_25155);
nand U25724 (N_25724,N_25245,N_25228);
nor U25725 (N_25725,N_25078,N_25422);
and U25726 (N_25726,N_25005,N_25378);
and U25727 (N_25727,N_25069,N_25282);
nand U25728 (N_25728,N_25171,N_25306);
nor U25729 (N_25729,N_25344,N_25258);
nand U25730 (N_25730,N_25480,N_25187);
nor U25731 (N_25731,N_25355,N_25456);
xnor U25732 (N_25732,N_25256,N_25251);
and U25733 (N_25733,N_25094,N_25315);
xnor U25734 (N_25734,N_25322,N_25070);
xnor U25735 (N_25735,N_25082,N_25455);
nand U25736 (N_25736,N_25040,N_25462);
nor U25737 (N_25737,N_25330,N_25107);
xnor U25738 (N_25738,N_25435,N_25340);
xor U25739 (N_25739,N_25447,N_25032);
nor U25740 (N_25740,N_25026,N_25398);
or U25741 (N_25741,N_25264,N_25441);
nor U25742 (N_25742,N_25268,N_25471);
or U25743 (N_25743,N_25207,N_25419);
and U25744 (N_25744,N_25249,N_25479);
nor U25745 (N_25745,N_25244,N_25186);
nand U25746 (N_25746,N_25043,N_25311);
nor U25747 (N_25747,N_25137,N_25396);
nand U25748 (N_25748,N_25198,N_25467);
xnor U25749 (N_25749,N_25346,N_25313);
and U25750 (N_25750,N_25489,N_25288);
or U25751 (N_25751,N_25074,N_25007);
or U25752 (N_25752,N_25019,N_25111);
and U25753 (N_25753,N_25219,N_25422);
nor U25754 (N_25754,N_25110,N_25468);
nor U25755 (N_25755,N_25213,N_25089);
xnor U25756 (N_25756,N_25360,N_25076);
nor U25757 (N_25757,N_25292,N_25483);
and U25758 (N_25758,N_25482,N_25488);
nand U25759 (N_25759,N_25475,N_25338);
xnor U25760 (N_25760,N_25196,N_25360);
nand U25761 (N_25761,N_25197,N_25340);
nor U25762 (N_25762,N_25072,N_25230);
xnor U25763 (N_25763,N_25234,N_25191);
xor U25764 (N_25764,N_25101,N_25420);
and U25765 (N_25765,N_25092,N_25366);
nor U25766 (N_25766,N_25116,N_25073);
nand U25767 (N_25767,N_25216,N_25463);
or U25768 (N_25768,N_25111,N_25483);
and U25769 (N_25769,N_25069,N_25437);
or U25770 (N_25770,N_25346,N_25064);
nor U25771 (N_25771,N_25133,N_25495);
nor U25772 (N_25772,N_25246,N_25358);
nand U25773 (N_25773,N_25047,N_25059);
xor U25774 (N_25774,N_25283,N_25129);
nand U25775 (N_25775,N_25101,N_25369);
or U25776 (N_25776,N_25109,N_25227);
nand U25777 (N_25777,N_25320,N_25026);
nand U25778 (N_25778,N_25061,N_25381);
nor U25779 (N_25779,N_25482,N_25220);
nor U25780 (N_25780,N_25177,N_25271);
or U25781 (N_25781,N_25230,N_25378);
nand U25782 (N_25782,N_25423,N_25141);
nand U25783 (N_25783,N_25140,N_25306);
and U25784 (N_25784,N_25433,N_25113);
and U25785 (N_25785,N_25023,N_25472);
and U25786 (N_25786,N_25207,N_25038);
nand U25787 (N_25787,N_25363,N_25147);
and U25788 (N_25788,N_25480,N_25098);
or U25789 (N_25789,N_25157,N_25168);
nand U25790 (N_25790,N_25037,N_25084);
nor U25791 (N_25791,N_25182,N_25134);
and U25792 (N_25792,N_25316,N_25174);
nand U25793 (N_25793,N_25233,N_25100);
nand U25794 (N_25794,N_25382,N_25428);
and U25795 (N_25795,N_25444,N_25429);
nor U25796 (N_25796,N_25295,N_25102);
nand U25797 (N_25797,N_25004,N_25231);
or U25798 (N_25798,N_25407,N_25150);
or U25799 (N_25799,N_25270,N_25072);
nor U25800 (N_25800,N_25266,N_25454);
nor U25801 (N_25801,N_25322,N_25139);
or U25802 (N_25802,N_25067,N_25450);
nand U25803 (N_25803,N_25233,N_25428);
or U25804 (N_25804,N_25235,N_25267);
xnor U25805 (N_25805,N_25164,N_25159);
nor U25806 (N_25806,N_25299,N_25458);
nor U25807 (N_25807,N_25370,N_25019);
or U25808 (N_25808,N_25233,N_25306);
or U25809 (N_25809,N_25428,N_25290);
xor U25810 (N_25810,N_25209,N_25026);
nand U25811 (N_25811,N_25372,N_25351);
xor U25812 (N_25812,N_25000,N_25052);
xor U25813 (N_25813,N_25468,N_25180);
and U25814 (N_25814,N_25026,N_25231);
nand U25815 (N_25815,N_25316,N_25307);
xor U25816 (N_25816,N_25029,N_25077);
and U25817 (N_25817,N_25354,N_25470);
and U25818 (N_25818,N_25093,N_25025);
nand U25819 (N_25819,N_25037,N_25085);
and U25820 (N_25820,N_25091,N_25415);
nor U25821 (N_25821,N_25124,N_25333);
xor U25822 (N_25822,N_25423,N_25038);
and U25823 (N_25823,N_25326,N_25301);
nor U25824 (N_25824,N_25100,N_25438);
or U25825 (N_25825,N_25089,N_25400);
nand U25826 (N_25826,N_25232,N_25474);
nand U25827 (N_25827,N_25286,N_25315);
nand U25828 (N_25828,N_25424,N_25241);
xor U25829 (N_25829,N_25401,N_25295);
or U25830 (N_25830,N_25411,N_25362);
nand U25831 (N_25831,N_25140,N_25315);
nor U25832 (N_25832,N_25482,N_25204);
nand U25833 (N_25833,N_25196,N_25131);
and U25834 (N_25834,N_25245,N_25169);
nand U25835 (N_25835,N_25467,N_25150);
nor U25836 (N_25836,N_25442,N_25437);
and U25837 (N_25837,N_25471,N_25202);
xnor U25838 (N_25838,N_25313,N_25499);
xnor U25839 (N_25839,N_25167,N_25046);
xnor U25840 (N_25840,N_25226,N_25102);
xnor U25841 (N_25841,N_25153,N_25323);
xnor U25842 (N_25842,N_25409,N_25495);
xnor U25843 (N_25843,N_25461,N_25227);
xnor U25844 (N_25844,N_25156,N_25409);
and U25845 (N_25845,N_25065,N_25045);
xnor U25846 (N_25846,N_25163,N_25196);
nor U25847 (N_25847,N_25249,N_25046);
and U25848 (N_25848,N_25218,N_25343);
xnor U25849 (N_25849,N_25398,N_25374);
or U25850 (N_25850,N_25135,N_25072);
xnor U25851 (N_25851,N_25342,N_25051);
xor U25852 (N_25852,N_25366,N_25177);
or U25853 (N_25853,N_25080,N_25059);
or U25854 (N_25854,N_25156,N_25391);
nor U25855 (N_25855,N_25434,N_25045);
or U25856 (N_25856,N_25146,N_25487);
and U25857 (N_25857,N_25298,N_25265);
nor U25858 (N_25858,N_25285,N_25452);
nor U25859 (N_25859,N_25173,N_25177);
nor U25860 (N_25860,N_25397,N_25422);
nor U25861 (N_25861,N_25399,N_25493);
and U25862 (N_25862,N_25272,N_25497);
xor U25863 (N_25863,N_25465,N_25400);
nor U25864 (N_25864,N_25407,N_25393);
nand U25865 (N_25865,N_25019,N_25007);
and U25866 (N_25866,N_25233,N_25287);
and U25867 (N_25867,N_25277,N_25021);
xnor U25868 (N_25868,N_25205,N_25045);
xnor U25869 (N_25869,N_25328,N_25329);
nand U25870 (N_25870,N_25004,N_25055);
and U25871 (N_25871,N_25283,N_25074);
nor U25872 (N_25872,N_25195,N_25017);
xnor U25873 (N_25873,N_25294,N_25456);
nand U25874 (N_25874,N_25005,N_25060);
and U25875 (N_25875,N_25204,N_25182);
or U25876 (N_25876,N_25448,N_25027);
or U25877 (N_25877,N_25416,N_25245);
or U25878 (N_25878,N_25011,N_25020);
nor U25879 (N_25879,N_25085,N_25239);
nand U25880 (N_25880,N_25045,N_25377);
nand U25881 (N_25881,N_25367,N_25140);
nand U25882 (N_25882,N_25320,N_25242);
or U25883 (N_25883,N_25392,N_25158);
or U25884 (N_25884,N_25453,N_25327);
and U25885 (N_25885,N_25099,N_25333);
and U25886 (N_25886,N_25159,N_25287);
or U25887 (N_25887,N_25157,N_25408);
xor U25888 (N_25888,N_25415,N_25296);
or U25889 (N_25889,N_25213,N_25429);
and U25890 (N_25890,N_25277,N_25101);
and U25891 (N_25891,N_25487,N_25484);
nor U25892 (N_25892,N_25218,N_25392);
nand U25893 (N_25893,N_25325,N_25153);
nand U25894 (N_25894,N_25043,N_25467);
and U25895 (N_25895,N_25287,N_25324);
xor U25896 (N_25896,N_25397,N_25002);
nor U25897 (N_25897,N_25340,N_25476);
xnor U25898 (N_25898,N_25118,N_25254);
nand U25899 (N_25899,N_25175,N_25486);
and U25900 (N_25900,N_25252,N_25357);
or U25901 (N_25901,N_25215,N_25437);
or U25902 (N_25902,N_25174,N_25199);
nor U25903 (N_25903,N_25348,N_25093);
nand U25904 (N_25904,N_25127,N_25128);
xnor U25905 (N_25905,N_25024,N_25091);
and U25906 (N_25906,N_25313,N_25099);
nor U25907 (N_25907,N_25213,N_25012);
nor U25908 (N_25908,N_25388,N_25375);
nand U25909 (N_25909,N_25155,N_25345);
and U25910 (N_25910,N_25432,N_25411);
xor U25911 (N_25911,N_25192,N_25132);
nand U25912 (N_25912,N_25362,N_25300);
nand U25913 (N_25913,N_25173,N_25043);
xnor U25914 (N_25914,N_25059,N_25179);
nand U25915 (N_25915,N_25245,N_25471);
xnor U25916 (N_25916,N_25267,N_25449);
nor U25917 (N_25917,N_25404,N_25120);
xnor U25918 (N_25918,N_25325,N_25299);
xnor U25919 (N_25919,N_25412,N_25238);
nand U25920 (N_25920,N_25234,N_25224);
nand U25921 (N_25921,N_25143,N_25480);
nor U25922 (N_25922,N_25089,N_25441);
xnor U25923 (N_25923,N_25346,N_25052);
nor U25924 (N_25924,N_25021,N_25201);
nand U25925 (N_25925,N_25335,N_25207);
or U25926 (N_25926,N_25099,N_25155);
nand U25927 (N_25927,N_25310,N_25303);
and U25928 (N_25928,N_25359,N_25160);
nand U25929 (N_25929,N_25208,N_25447);
nand U25930 (N_25930,N_25214,N_25470);
nor U25931 (N_25931,N_25094,N_25006);
and U25932 (N_25932,N_25293,N_25162);
or U25933 (N_25933,N_25074,N_25320);
or U25934 (N_25934,N_25212,N_25091);
xnor U25935 (N_25935,N_25469,N_25130);
nor U25936 (N_25936,N_25419,N_25136);
nand U25937 (N_25937,N_25359,N_25423);
nor U25938 (N_25938,N_25490,N_25369);
or U25939 (N_25939,N_25166,N_25412);
nor U25940 (N_25940,N_25446,N_25303);
or U25941 (N_25941,N_25060,N_25020);
nor U25942 (N_25942,N_25363,N_25415);
nor U25943 (N_25943,N_25134,N_25139);
xor U25944 (N_25944,N_25475,N_25263);
nor U25945 (N_25945,N_25153,N_25263);
or U25946 (N_25946,N_25420,N_25352);
or U25947 (N_25947,N_25359,N_25043);
nor U25948 (N_25948,N_25128,N_25139);
nand U25949 (N_25949,N_25395,N_25079);
or U25950 (N_25950,N_25032,N_25406);
xor U25951 (N_25951,N_25163,N_25313);
nor U25952 (N_25952,N_25079,N_25140);
or U25953 (N_25953,N_25256,N_25396);
xor U25954 (N_25954,N_25375,N_25142);
nand U25955 (N_25955,N_25094,N_25412);
nand U25956 (N_25956,N_25280,N_25071);
nor U25957 (N_25957,N_25359,N_25208);
or U25958 (N_25958,N_25095,N_25030);
nand U25959 (N_25959,N_25111,N_25328);
nand U25960 (N_25960,N_25370,N_25073);
nand U25961 (N_25961,N_25016,N_25188);
xnor U25962 (N_25962,N_25475,N_25106);
nand U25963 (N_25963,N_25053,N_25374);
xor U25964 (N_25964,N_25431,N_25480);
and U25965 (N_25965,N_25486,N_25325);
and U25966 (N_25966,N_25218,N_25009);
and U25967 (N_25967,N_25348,N_25234);
nand U25968 (N_25968,N_25232,N_25432);
or U25969 (N_25969,N_25473,N_25161);
xor U25970 (N_25970,N_25247,N_25267);
nand U25971 (N_25971,N_25462,N_25234);
nand U25972 (N_25972,N_25302,N_25391);
xor U25973 (N_25973,N_25013,N_25165);
nand U25974 (N_25974,N_25069,N_25016);
nand U25975 (N_25975,N_25343,N_25031);
xor U25976 (N_25976,N_25225,N_25020);
nand U25977 (N_25977,N_25094,N_25261);
nor U25978 (N_25978,N_25127,N_25482);
or U25979 (N_25979,N_25006,N_25303);
nand U25980 (N_25980,N_25003,N_25475);
xnor U25981 (N_25981,N_25272,N_25401);
nand U25982 (N_25982,N_25389,N_25374);
and U25983 (N_25983,N_25116,N_25381);
or U25984 (N_25984,N_25038,N_25465);
xor U25985 (N_25985,N_25095,N_25010);
and U25986 (N_25986,N_25102,N_25167);
xor U25987 (N_25987,N_25317,N_25282);
nor U25988 (N_25988,N_25263,N_25329);
nor U25989 (N_25989,N_25044,N_25362);
and U25990 (N_25990,N_25224,N_25420);
nor U25991 (N_25991,N_25432,N_25499);
nand U25992 (N_25992,N_25110,N_25192);
and U25993 (N_25993,N_25060,N_25120);
nor U25994 (N_25994,N_25383,N_25102);
or U25995 (N_25995,N_25110,N_25235);
or U25996 (N_25996,N_25246,N_25177);
xnor U25997 (N_25997,N_25145,N_25341);
nor U25998 (N_25998,N_25485,N_25103);
nor U25999 (N_25999,N_25007,N_25029);
and U26000 (N_26000,N_25882,N_25660);
or U26001 (N_26001,N_25588,N_25535);
xor U26002 (N_26002,N_25567,N_25598);
nor U26003 (N_26003,N_25619,N_25876);
and U26004 (N_26004,N_25538,N_25667);
nor U26005 (N_26005,N_25819,N_25825);
nand U26006 (N_26006,N_25738,N_25557);
or U26007 (N_26007,N_25569,N_25613);
nand U26008 (N_26008,N_25663,N_25893);
xnor U26009 (N_26009,N_25665,N_25718);
and U26010 (N_26010,N_25706,N_25890);
nor U26011 (N_26011,N_25549,N_25818);
and U26012 (N_26012,N_25510,N_25631);
or U26013 (N_26013,N_25776,N_25673);
or U26014 (N_26014,N_25836,N_25935);
xor U26015 (N_26015,N_25753,N_25903);
nand U26016 (N_26016,N_25958,N_25519);
xnor U26017 (N_26017,N_25912,N_25957);
and U26018 (N_26018,N_25642,N_25700);
nor U26019 (N_26019,N_25733,N_25998);
or U26020 (N_26020,N_25769,N_25944);
nor U26021 (N_26021,N_25921,N_25953);
nand U26022 (N_26022,N_25961,N_25950);
xor U26023 (N_26023,N_25584,N_25879);
nor U26024 (N_26024,N_25767,N_25575);
nor U26025 (N_26025,N_25737,N_25990);
and U26026 (N_26026,N_25938,N_25609);
xnor U26027 (N_26027,N_25726,N_25620);
and U26028 (N_26028,N_25621,N_25864);
nor U26029 (N_26029,N_25989,N_25765);
and U26030 (N_26030,N_25856,N_25860);
nand U26031 (N_26031,N_25565,N_25992);
and U26032 (N_26032,N_25949,N_25698);
xor U26033 (N_26033,N_25604,N_25951);
or U26034 (N_26034,N_25833,N_25994);
and U26035 (N_26035,N_25537,N_25979);
xor U26036 (N_26036,N_25791,N_25750);
or U26037 (N_26037,N_25740,N_25822);
or U26038 (N_26038,N_25830,N_25746);
or U26039 (N_26039,N_25674,N_25939);
and U26040 (N_26040,N_25911,N_25517);
nand U26041 (N_26041,N_25555,N_25647);
and U26042 (N_26042,N_25947,N_25844);
nand U26043 (N_26043,N_25869,N_25579);
nor U26044 (N_26044,N_25832,N_25601);
xnor U26045 (N_26045,N_25919,N_25716);
nor U26046 (N_26046,N_25834,N_25861);
or U26047 (N_26047,N_25697,N_25996);
or U26048 (N_26048,N_25801,N_25850);
and U26049 (N_26049,N_25816,N_25880);
nor U26050 (N_26050,N_25679,N_25845);
and U26051 (N_26051,N_25997,N_25981);
nor U26052 (N_26052,N_25523,N_25884);
nand U26053 (N_26053,N_25595,N_25914);
or U26054 (N_26054,N_25973,N_25752);
and U26055 (N_26055,N_25954,N_25702);
nand U26056 (N_26056,N_25943,N_25648);
and U26057 (N_26057,N_25751,N_25859);
xnor U26058 (N_26058,N_25960,N_25886);
nand U26059 (N_26059,N_25562,N_25932);
xor U26060 (N_26060,N_25657,N_25993);
xnor U26061 (N_26061,N_25787,N_25682);
xor U26062 (N_26062,N_25675,N_25683);
xnor U26063 (N_26063,N_25605,N_25867);
nand U26064 (N_26064,N_25590,N_25587);
or U26065 (N_26065,N_25863,N_25942);
nor U26066 (N_26066,N_25891,N_25540);
nand U26067 (N_26067,N_25550,N_25536);
nor U26068 (N_26068,N_25570,N_25785);
xor U26069 (N_26069,N_25987,N_25909);
nor U26070 (N_26070,N_25573,N_25518);
or U26071 (N_26071,N_25759,N_25501);
xor U26072 (N_26072,N_25731,N_25813);
nand U26073 (N_26073,N_25678,N_25762);
nand U26074 (N_26074,N_25611,N_25786);
nor U26075 (N_26075,N_25623,N_25976);
or U26076 (N_26076,N_25862,N_25883);
nand U26077 (N_26077,N_25999,N_25824);
or U26078 (N_26078,N_25927,N_25758);
and U26079 (N_26079,N_25815,N_25618);
or U26080 (N_26080,N_25991,N_25571);
or U26081 (N_26081,N_25548,N_25881);
and U26082 (N_26082,N_25946,N_25616);
and U26083 (N_26083,N_25659,N_25610);
nand U26084 (N_26084,N_25676,N_25553);
xnor U26085 (N_26085,N_25877,N_25823);
and U26086 (N_26086,N_25761,N_25800);
nand U26087 (N_26087,N_25736,N_25608);
or U26088 (N_26088,N_25978,N_25624);
xnor U26089 (N_26089,N_25809,N_25520);
nor U26090 (N_26090,N_25617,N_25808);
nor U26091 (N_26091,N_25664,N_25905);
or U26092 (N_26092,N_25709,N_25757);
nor U26093 (N_26093,N_25637,N_25839);
nor U26094 (N_26094,N_25546,N_25693);
xor U26095 (N_26095,N_25730,N_25628);
xor U26096 (N_26096,N_25748,N_25975);
nand U26097 (N_26097,N_25929,N_25955);
or U26098 (N_26098,N_25967,N_25796);
xnor U26099 (N_26099,N_25645,N_25739);
nand U26100 (N_26100,N_25928,N_25783);
nand U26101 (N_26101,N_25687,N_25849);
and U26102 (N_26102,N_25710,N_25962);
xor U26103 (N_26103,N_25560,N_25626);
and U26104 (N_26104,N_25715,N_25545);
and U26105 (N_26105,N_25968,N_25666);
or U26106 (N_26106,N_25717,N_25980);
nand U26107 (N_26107,N_25896,N_25803);
nor U26108 (N_26108,N_25853,N_25887);
nand U26109 (N_26109,N_25904,N_25742);
or U26110 (N_26110,N_25743,N_25846);
xnor U26111 (N_26111,N_25556,N_25554);
and U26112 (N_26112,N_25577,N_25649);
nor U26113 (N_26113,N_25685,N_25827);
nor U26114 (N_26114,N_25531,N_25563);
nor U26115 (N_26115,N_25582,N_25744);
xnor U26116 (N_26116,N_25564,N_25872);
nand U26117 (N_26117,N_25515,N_25894);
or U26118 (N_26118,N_25977,N_25782);
or U26119 (N_26119,N_25747,N_25754);
nand U26120 (N_26120,N_25603,N_25910);
xor U26121 (N_26121,N_25964,N_25671);
xnor U26122 (N_26122,N_25866,N_25541);
and U26123 (N_26123,N_25734,N_25615);
xnor U26124 (N_26124,N_25724,N_25695);
and U26125 (N_26125,N_25639,N_25897);
nor U26126 (N_26126,N_25551,N_25918);
or U26127 (N_26127,N_25773,N_25574);
nor U26128 (N_26128,N_25692,N_25995);
or U26129 (N_26129,N_25811,N_25865);
nand U26130 (N_26130,N_25719,N_25511);
nand U26131 (N_26131,N_25804,N_25526);
and U26132 (N_26132,N_25802,N_25646);
or U26133 (N_26133,N_25841,N_25922);
or U26134 (N_26134,N_25707,N_25542);
xor U26135 (N_26135,N_25721,N_25847);
and U26136 (N_26136,N_25771,N_25788);
xnor U26137 (N_26137,N_25636,N_25908);
or U26138 (N_26138,N_25656,N_25745);
nor U26139 (N_26139,N_25677,N_25712);
xnor U26140 (N_26140,N_25505,N_25901);
xor U26141 (N_26141,N_25622,N_25766);
and U26142 (N_26142,N_25874,N_25680);
xor U26143 (N_26143,N_25798,N_25760);
xor U26144 (N_26144,N_25727,N_25848);
nand U26145 (N_26145,N_25627,N_25583);
and U26146 (N_26146,N_25855,N_25539);
nand U26147 (N_26147,N_25755,N_25774);
xnor U26148 (N_26148,N_25530,N_25658);
xnor U26149 (N_26149,N_25831,N_25696);
nand U26150 (N_26150,N_25516,N_25508);
nand U26151 (N_26151,N_25934,N_25749);
xor U26152 (N_26152,N_25597,N_25820);
nand U26153 (N_26153,N_25593,N_25906);
or U26154 (N_26154,N_25889,N_25524);
nor U26155 (N_26155,N_25789,N_25728);
nor U26156 (N_26156,N_25837,N_25966);
xnor U26157 (N_26157,N_25821,N_25925);
nand U26158 (N_26158,N_25913,N_25552);
xor U26159 (N_26159,N_25795,N_25689);
and U26160 (N_26160,N_25591,N_25888);
nor U26161 (N_26161,N_25948,N_25703);
and U26162 (N_26162,N_25580,N_25655);
or U26163 (N_26163,N_25875,N_25920);
or U26164 (N_26164,N_25956,N_25654);
and U26165 (N_26165,N_25629,N_25506);
and U26166 (N_26166,N_25878,N_25561);
xor U26167 (N_26167,N_25529,N_25917);
nand U26168 (N_26168,N_25971,N_25694);
xnor U26169 (N_26169,N_25784,N_25500);
or U26170 (N_26170,N_25858,N_25568);
and U26171 (N_26171,N_25764,N_25982);
xnor U26172 (N_26172,N_25756,N_25638);
nor U26173 (N_26173,N_25547,N_25525);
and U26174 (N_26174,N_25777,N_25514);
and U26175 (N_26175,N_25916,N_25793);
nand U26176 (N_26176,N_25691,N_25732);
and U26177 (N_26177,N_25632,N_25681);
nand U26178 (N_26178,N_25959,N_25868);
nand U26179 (N_26179,N_25504,N_25662);
nor U26180 (N_26180,N_25670,N_25870);
nand U26181 (N_26181,N_25974,N_25779);
nand U26182 (N_26182,N_25576,N_25794);
and U26183 (N_26183,N_25594,N_25528);
nor U26184 (N_26184,N_25521,N_25701);
nand U26185 (N_26185,N_25778,N_25988);
nor U26186 (N_26186,N_25634,N_25838);
nand U26187 (N_26187,N_25507,N_25902);
nor U26188 (N_26188,N_25720,N_25690);
nor U26189 (N_26189,N_25923,N_25814);
and U26190 (N_26190,N_25614,N_25599);
nand U26191 (N_26191,N_25713,N_25699);
or U26192 (N_26192,N_25805,N_25770);
nor U26193 (N_26193,N_25945,N_25892);
xnor U26194 (N_26194,N_25963,N_25635);
nand U26195 (N_26195,N_25899,N_25533);
nand U26196 (N_26196,N_25503,N_25711);
nor U26197 (N_26197,N_25607,N_25790);
and U26198 (N_26198,N_25596,N_25653);
or U26199 (N_26199,N_25527,N_25566);
and U26200 (N_26200,N_25741,N_25926);
nor U26201 (N_26201,N_25592,N_25723);
nand U26202 (N_26202,N_25797,N_25852);
xor U26203 (N_26203,N_25768,N_25842);
or U26204 (N_26204,N_25650,N_25984);
xnor U26205 (N_26205,N_25781,N_25885);
nand U26206 (N_26206,N_25644,N_25807);
and U26207 (N_26207,N_25986,N_25985);
or U26208 (N_26208,N_25581,N_25600);
xnor U26209 (N_26209,N_25625,N_25602);
nor U26210 (N_26210,N_25606,N_25651);
xnor U26211 (N_26211,N_25895,N_25806);
nor U26212 (N_26212,N_25840,N_25970);
xnor U26213 (N_26213,N_25729,N_25969);
xor U26214 (N_26214,N_25633,N_25502);
and U26215 (N_26215,N_25708,N_25792);
nor U26216 (N_26216,N_25915,N_25672);
and U26217 (N_26217,N_25668,N_25688);
and U26218 (N_26218,N_25835,N_25725);
xnor U26219 (N_26219,N_25640,N_25965);
and U26220 (N_26220,N_25763,N_25643);
nand U26221 (N_26221,N_25686,N_25843);
nor U26222 (N_26222,N_25936,N_25543);
nand U26223 (N_26223,N_25854,N_25873);
or U26224 (N_26224,N_25705,N_25829);
xor U26225 (N_26225,N_25810,N_25930);
xnor U26226 (N_26226,N_25534,N_25722);
and U26227 (N_26227,N_25585,N_25612);
and U26228 (N_26228,N_25513,N_25817);
nand U26229 (N_26229,N_25669,N_25772);
nand U26230 (N_26230,N_25558,N_25972);
nand U26231 (N_26231,N_25812,N_25544);
and U26232 (N_26232,N_25589,N_25684);
nor U26233 (N_26233,N_25907,N_25780);
and U26234 (N_26234,N_25871,N_25559);
xnor U26235 (N_26235,N_25641,N_25826);
nand U26236 (N_26236,N_25704,N_25952);
xor U26237 (N_26237,N_25983,N_25898);
and U26238 (N_26238,N_25940,N_25522);
xor U26239 (N_26239,N_25652,N_25735);
or U26240 (N_26240,N_25828,N_25851);
or U26241 (N_26241,N_25900,N_25775);
or U26242 (N_26242,N_25509,N_25924);
nand U26243 (N_26243,N_25661,N_25799);
nand U26244 (N_26244,N_25586,N_25578);
or U26245 (N_26245,N_25572,N_25933);
xor U26246 (N_26246,N_25857,N_25630);
nor U26247 (N_26247,N_25714,N_25931);
and U26248 (N_26248,N_25937,N_25512);
or U26249 (N_26249,N_25532,N_25941);
xnor U26250 (N_26250,N_25794,N_25748);
nor U26251 (N_26251,N_25563,N_25656);
nand U26252 (N_26252,N_25504,N_25908);
xnor U26253 (N_26253,N_25532,N_25602);
or U26254 (N_26254,N_25572,N_25941);
nand U26255 (N_26255,N_25504,N_25511);
and U26256 (N_26256,N_25884,N_25588);
xnor U26257 (N_26257,N_25922,N_25979);
xor U26258 (N_26258,N_25980,N_25783);
and U26259 (N_26259,N_25756,N_25836);
xnor U26260 (N_26260,N_25891,N_25855);
or U26261 (N_26261,N_25557,N_25943);
nand U26262 (N_26262,N_25603,N_25999);
and U26263 (N_26263,N_25832,N_25735);
xnor U26264 (N_26264,N_25666,N_25835);
or U26265 (N_26265,N_25693,N_25695);
nor U26266 (N_26266,N_25829,N_25633);
xnor U26267 (N_26267,N_25518,N_25881);
and U26268 (N_26268,N_25943,N_25812);
nor U26269 (N_26269,N_25861,N_25958);
or U26270 (N_26270,N_25709,N_25616);
and U26271 (N_26271,N_25869,N_25714);
or U26272 (N_26272,N_25655,N_25530);
or U26273 (N_26273,N_25967,N_25756);
nand U26274 (N_26274,N_25666,N_25920);
and U26275 (N_26275,N_25682,N_25987);
xor U26276 (N_26276,N_25730,N_25792);
or U26277 (N_26277,N_25780,N_25594);
and U26278 (N_26278,N_25931,N_25948);
and U26279 (N_26279,N_25607,N_25535);
or U26280 (N_26280,N_25740,N_25627);
and U26281 (N_26281,N_25933,N_25581);
and U26282 (N_26282,N_25838,N_25763);
xnor U26283 (N_26283,N_25654,N_25865);
nor U26284 (N_26284,N_25971,N_25671);
or U26285 (N_26285,N_25571,N_25939);
or U26286 (N_26286,N_25533,N_25977);
nand U26287 (N_26287,N_25610,N_25560);
xor U26288 (N_26288,N_25676,N_25873);
or U26289 (N_26289,N_25901,N_25947);
nand U26290 (N_26290,N_25987,N_25976);
nor U26291 (N_26291,N_25865,N_25771);
and U26292 (N_26292,N_25926,N_25716);
nor U26293 (N_26293,N_25705,N_25614);
nand U26294 (N_26294,N_25951,N_25699);
or U26295 (N_26295,N_25931,N_25538);
nor U26296 (N_26296,N_25836,N_25875);
nand U26297 (N_26297,N_25690,N_25898);
or U26298 (N_26298,N_25927,N_25503);
nand U26299 (N_26299,N_25842,N_25612);
nor U26300 (N_26300,N_25563,N_25607);
or U26301 (N_26301,N_25868,N_25513);
xor U26302 (N_26302,N_25530,N_25721);
xor U26303 (N_26303,N_25510,N_25647);
nor U26304 (N_26304,N_25947,N_25509);
or U26305 (N_26305,N_25572,N_25612);
nor U26306 (N_26306,N_25849,N_25708);
nor U26307 (N_26307,N_25659,N_25609);
nor U26308 (N_26308,N_25755,N_25794);
or U26309 (N_26309,N_25701,N_25733);
nand U26310 (N_26310,N_25882,N_25520);
nor U26311 (N_26311,N_25731,N_25702);
and U26312 (N_26312,N_25968,N_25665);
and U26313 (N_26313,N_25563,N_25707);
xnor U26314 (N_26314,N_25976,N_25700);
and U26315 (N_26315,N_25969,N_25697);
nand U26316 (N_26316,N_25720,N_25933);
xor U26317 (N_26317,N_25753,N_25795);
nand U26318 (N_26318,N_25515,N_25544);
nor U26319 (N_26319,N_25632,N_25849);
nor U26320 (N_26320,N_25848,N_25990);
and U26321 (N_26321,N_25792,N_25987);
and U26322 (N_26322,N_25671,N_25847);
nor U26323 (N_26323,N_25726,N_25982);
nand U26324 (N_26324,N_25795,N_25737);
nand U26325 (N_26325,N_25647,N_25716);
or U26326 (N_26326,N_25559,N_25982);
nand U26327 (N_26327,N_25626,N_25999);
xnor U26328 (N_26328,N_25641,N_25643);
nor U26329 (N_26329,N_25591,N_25554);
or U26330 (N_26330,N_25693,N_25774);
nor U26331 (N_26331,N_25948,N_25541);
xnor U26332 (N_26332,N_25951,N_25961);
or U26333 (N_26333,N_25666,N_25755);
or U26334 (N_26334,N_25981,N_25719);
or U26335 (N_26335,N_25950,N_25908);
xnor U26336 (N_26336,N_25515,N_25920);
nor U26337 (N_26337,N_25551,N_25871);
xnor U26338 (N_26338,N_25676,N_25661);
xor U26339 (N_26339,N_25887,N_25975);
and U26340 (N_26340,N_25856,N_25984);
xnor U26341 (N_26341,N_25651,N_25891);
xor U26342 (N_26342,N_25917,N_25889);
and U26343 (N_26343,N_25752,N_25646);
nor U26344 (N_26344,N_25831,N_25794);
and U26345 (N_26345,N_25645,N_25512);
nand U26346 (N_26346,N_25524,N_25684);
and U26347 (N_26347,N_25848,N_25711);
or U26348 (N_26348,N_25821,N_25904);
nand U26349 (N_26349,N_25766,N_25733);
xnor U26350 (N_26350,N_25973,N_25993);
nor U26351 (N_26351,N_25590,N_25766);
and U26352 (N_26352,N_25831,N_25892);
and U26353 (N_26353,N_25859,N_25934);
xor U26354 (N_26354,N_25943,N_25878);
and U26355 (N_26355,N_25536,N_25698);
nor U26356 (N_26356,N_25807,N_25761);
or U26357 (N_26357,N_25723,N_25747);
xor U26358 (N_26358,N_25735,N_25640);
and U26359 (N_26359,N_25867,N_25838);
and U26360 (N_26360,N_25899,N_25894);
nor U26361 (N_26361,N_25707,N_25526);
and U26362 (N_26362,N_25524,N_25716);
xor U26363 (N_26363,N_25769,N_25592);
or U26364 (N_26364,N_25995,N_25940);
nand U26365 (N_26365,N_25570,N_25782);
nand U26366 (N_26366,N_25769,N_25945);
or U26367 (N_26367,N_25664,N_25768);
or U26368 (N_26368,N_25843,N_25764);
or U26369 (N_26369,N_25898,N_25560);
nor U26370 (N_26370,N_25532,N_25694);
xor U26371 (N_26371,N_25928,N_25551);
or U26372 (N_26372,N_25543,N_25540);
xor U26373 (N_26373,N_25518,N_25542);
or U26374 (N_26374,N_25725,N_25574);
and U26375 (N_26375,N_25673,N_25572);
and U26376 (N_26376,N_25868,N_25728);
nand U26377 (N_26377,N_25543,N_25750);
nor U26378 (N_26378,N_25615,N_25948);
xnor U26379 (N_26379,N_25776,N_25771);
nand U26380 (N_26380,N_25697,N_25731);
nor U26381 (N_26381,N_25666,N_25689);
nand U26382 (N_26382,N_25980,N_25765);
nor U26383 (N_26383,N_25945,N_25934);
and U26384 (N_26384,N_25710,N_25842);
and U26385 (N_26385,N_25608,N_25652);
and U26386 (N_26386,N_25651,N_25586);
and U26387 (N_26387,N_25895,N_25840);
nand U26388 (N_26388,N_25937,N_25616);
nor U26389 (N_26389,N_25612,N_25795);
nor U26390 (N_26390,N_25746,N_25736);
nor U26391 (N_26391,N_25603,N_25917);
and U26392 (N_26392,N_25774,N_25606);
or U26393 (N_26393,N_25832,N_25992);
xnor U26394 (N_26394,N_25658,N_25951);
xor U26395 (N_26395,N_25536,N_25879);
nor U26396 (N_26396,N_25648,N_25535);
or U26397 (N_26397,N_25678,N_25917);
xor U26398 (N_26398,N_25557,N_25734);
nor U26399 (N_26399,N_25761,N_25693);
and U26400 (N_26400,N_25657,N_25953);
nor U26401 (N_26401,N_25948,N_25737);
nand U26402 (N_26402,N_25685,N_25830);
and U26403 (N_26403,N_25722,N_25936);
nor U26404 (N_26404,N_25732,N_25839);
nor U26405 (N_26405,N_25515,N_25649);
or U26406 (N_26406,N_25568,N_25971);
and U26407 (N_26407,N_25524,N_25544);
nand U26408 (N_26408,N_25519,N_25866);
xor U26409 (N_26409,N_25563,N_25890);
nor U26410 (N_26410,N_25923,N_25505);
or U26411 (N_26411,N_25993,N_25671);
or U26412 (N_26412,N_25959,N_25696);
and U26413 (N_26413,N_25705,N_25761);
nand U26414 (N_26414,N_25915,N_25650);
nand U26415 (N_26415,N_25908,N_25881);
nand U26416 (N_26416,N_25820,N_25579);
and U26417 (N_26417,N_25725,N_25874);
and U26418 (N_26418,N_25938,N_25661);
nand U26419 (N_26419,N_25582,N_25680);
and U26420 (N_26420,N_25856,N_25876);
nand U26421 (N_26421,N_25844,N_25572);
and U26422 (N_26422,N_25962,N_25931);
and U26423 (N_26423,N_25821,N_25823);
or U26424 (N_26424,N_25992,N_25748);
nor U26425 (N_26425,N_25569,N_25573);
nand U26426 (N_26426,N_25808,N_25541);
xor U26427 (N_26427,N_25812,N_25999);
xor U26428 (N_26428,N_25685,N_25515);
and U26429 (N_26429,N_25502,N_25877);
xnor U26430 (N_26430,N_25713,N_25512);
or U26431 (N_26431,N_25808,N_25640);
nand U26432 (N_26432,N_25516,N_25776);
and U26433 (N_26433,N_25604,N_25684);
or U26434 (N_26434,N_25801,N_25585);
nor U26435 (N_26435,N_25644,N_25843);
and U26436 (N_26436,N_25882,N_25608);
nor U26437 (N_26437,N_25707,N_25792);
nor U26438 (N_26438,N_25840,N_25774);
nor U26439 (N_26439,N_25769,N_25635);
or U26440 (N_26440,N_25669,N_25644);
and U26441 (N_26441,N_25835,N_25994);
or U26442 (N_26442,N_25553,N_25826);
xnor U26443 (N_26443,N_25621,N_25529);
nand U26444 (N_26444,N_25941,N_25948);
or U26445 (N_26445,N_25634,N_25833);
nor U26446 (N_26446,N_25996,N_25910);
xnor U26447 (N_26447,N_25678,N_25649);
and U26448 (N_26448,N_25529,N_25655);
and U26449 (N_26449,N_25645,N_25692);
xnor U26450 (N_26450,N_25510,N_25541);
or U26451 (N_26451,N_25756,N_25615);
and U26452 (N_26452,N_25980,N_25876);
xnor U26453 (N_26453,N_25544,N_25953);
xnor U26454 (N_26454,N_25520,N_25582);
and U26455 (N_26455,N_25730,N_25715);
and U26456 (N_26456,N_25768,N_25765);
xor U26457 (N_26457,N_25967,N_25844);
and U26458 (N_26458,N_25656,N_25742);
or U26459 (N_26459,N_25535,N_25668);
nand U26460 (N_26460,N_25957,N_25654);
and U26461 (N_26461,N_25869,N_25912);
nor U26462 (N_26462,N_25991,N_25523);
nand U26463 (N_26463,N_25693,N_25960);
xnor U26464 (N_26464,N_25678,N_25916);
or U26465 (N_26465,N_25915,N_25929);
xnor U26466 (N_26466,N_25813,N_25922);
or U26467 (N_26467,N_25734,N_25981);
and U26468 (N_26468,N_25649,N_25847);
nand U26469 (N_26469,N_25556,N_25502);
nand U26470 (N_26470,N_25876,N_25972);
xor U26471 (N_26471,N_25780,N_25547);
or U26472 (N_26472,N_25930,N_25929);
and U26473 (N_26473,N_25710,N_25886);
xnor U26474 (N_26474,N_25721,N_25537);
nor U26475 (N_26475,N_25754,N_25689);
and U26476 (N_26476,N_25608,N_25708);
or U26477 (N_26477,N_25838,N_25759);
nor U26478 (N_26478,N_25721,N_25697);
or U26479 (N_26479,N_25538,N_25985);
xnor U26480 (N_26480,N_25788,N_25761);
nor U26481 (N_26481,N_25852,N_25939);
xor U26482 (N_26482,N_25874,N_25786);
or U26483 (N_26483,N_25827,N_25923);
or U26484 (N_26484,N_25658,N_25725);
nand U26485 (N_26485,N_25780,N_25679);
nor U26486 (N_26486,N_25978,N_25810);
nand U26487 (N_26487,N_25982,N_25716);
nor U26488 (N_26488,N_25593,N_25813);
and U26489 (N_26489,N_25547,N_25832);
nand U26490 (N_26490,N_25935,N_25621);
nand U26491 (N_26491,N_25585,N_25641);
or U26492 (N_26492,N_25682,N_25799);
nand U26493 (N_26493,N_25555,N_25649);
xor U26494 (N_26494,N_25551,N_25990);
nor U26495 (N_26495,N_25528,N_25522);
and U26496 (N_26496,N_25862,N_25788);
xnor U26497 (N_26497,N_25519,N_25859);
nand U26498 (N_26498,N_25620,N_25998);
xor U26499 (N_26499,N_25700,N_25873);
or U26500 (N_26500,N_26238,N_26225);
xnor U26501 (N_26501,N_26207,N_26143);
nor U26502 (N_26502,N_26179,N_26233);
nor U26503 (N_26503,N_26312,N_26182);
nor U26504 (N_26504,N_26253,N_26363);
and U26505 (N_26505,N_26132,N_26329);
and U26506 (N_26506,N_26416,N_26126);
nand U26507 (N_26507,N_26339,N_26055);
or U26508 (N_26508,N_26473,N_26311);
xnor U26509 (N_26509,N_26345,N_26064);
nor U26510 (N_26510,N_26136,N_26069);
nor U26511 (N_26511,N_26034,N_26153);
nor U26512 (N_26512,N_26445,N_26455);
or U26513 (N_26513,N_26171,N_26172);
and U26514 (N_26514,N_26111,N_26092);
nor U26515 (N_26515,N_26277,N_26439);
nand U26516 (N_26516,N_26062,N_26291);
and U26517 (N_26517,N_26008,N_26467);
nor U26518 (N_26518,N_26086,N_26316);
or U26519 (N_26519,N_26141,N_26364);
nand U26520 (N_26520,N_26059,N_26293);
nand U26521 (N_26521,N_26476,N_26429);
or U26522 (N_26522,N_26303,N_26283);
or U26523 (N_26523,N_26464,N_26302);
and U26524 (N_26524,N_26498,N_26217);
nand U26525 (N_26525,N_26334,N_26355);
nor U26526 (N_26526,N_26343,N_26084);
or U26527 (N_26527,N_26076,N_26367);
or U26528 (N_26528,N_26384,N_26251);
nor U26529 (N_26529,N_26139,N_26221);
nand U26530 (N_26530,N_26072,N_26266);
xnor U26531 (N_26531,N_26351,N_26104);
nand U26532 (N_26532,N_26397,N_26317);
nand U26533 (N_26533,N_26360,N_26336);
xor U26534 (N_26534,N_26109,N_26160);
nor U26535 (N_26535,N_26054,N_26427);
or U26536 (N_26536,N_26030,N_26256);
nand U26537 (N_26537,N_26041,N_26080);
nor U26538 (N_26538,N_26057,N_26169);
xnor U26539 (N_26539,N_26197,N_26496);
nor U26540 (N_26540,N_26257,N_26484);
or U26541 (N_26541,N_26070,N_26003);
nand U26542 (N_26542,N_26088,N_26142);
nand U26543 (N_26543,N_26382,N_26078);
nor U26544 (N_26544,N_26394,N_26258);
nor U26545 (N_26545,N_26438,N_26051);
or U26546 (N_26546,N_26465,N_26434);
nand U26547 (N_26547,N_26457,N_26239);
or U26548 (N_26548,N_26131,N_26102);
or U26549 (N_26549,N_26009,N_26292);
nand U26550 (N_26550,N_26278,N_26396);
and U26551 (N_26551,N_26101,N_26375);
xor U26552 (N_26552,N_26175,N_26401);
nand U26553 (N_26553,N_26499,N_26214);
nand U26554 (N_26554,N_26468,N_26341);
nor U26555 (N_26555,N_26288,N_26349);
nor U26556 (N_26556,N_26323,N_26006);
nor U26557 (N_26557,N_26276,N_26268);
or U26558 (N_26558,N_26218,N_26342);
or U26559 (N_26559,N_26249,N_26108);
and U26560 (N_26560,N_26454,N_26133);
nand U26561 (N_26561,N_26184,N_26494);
xor U26562 (N_26562,N_26358,N_26315);
nand U26563 (N_26563,N_26155,N_26081);
nand U26564 (N_26564,N_26159,N_26227);
xnor U26565 (N_26565,N_26428,N_26065);
xnor U26566 (N_26566,N_26408,N_26318);
xnor U26567 (N_26567,N_26196,N_26486);
and U26568 (N_26568,N_26448,N_26449);
or U26569 (N_26569,N_26422,N_26463);
or U26570 (N_26570,N_26226,N_26340);
or U26571 (N_26571,N_26407,N_26058);
and U26572 (N_26572,N_26071,N_26432);
nand U26573 (N_26573,N_26451,N_26387);
and U26574 (N_26574,N_26304,N_26223);
xnor U26575 (N_26575,N_26335,N_26123);
or U26576 (N_26576,N_26301,N_26314);
or U26577 (N_26577,N_26279,N_26442);
xnor U26578 (N_26578,N_26150,N_26014);
xnor U26579 (N_26579,N_26391,N_26145);
or U26580 (N_26580,N_26435,N_26048);
nand U26581 (N_26581,N_26286,N_26440);
nor U26582 (N_26582,N_26362,N_26479);
xor U26583 (N_26583,N_26491,N_26074);
xnor U26584 (N_26584,N_26452,N_26043);
or U26585 (N_26585,N_26294,N_26471);
or U26586 (N_26586,N_26200,N_26398);
or U26587 (N_26587,N_26211,N_26322);
or U26588 (N_26588,N_26299,N_26489);
and U26589 (N_26589,N_26333,N_26002);
xnor U26590 (N_26590,N_26296,N_26114);
and U26591 (N_26591,N_26356,N_26320);
or U26592 (N_26592,N_26147,N_26120);
and U26593 (N_26593,N_26068,N_26377);
and U26594 (N_26594,N_26230,N_26017);
or U26595 (N_26595,N_26488,N_26269);
xor U26596 (N_26596,N_26426,N_26411);
xor U26597 (N_26597,N_26099,N_26388);
xnor U26598 (N_26598,N_26161,N_26485);
xor U26599 (N_26599,N_26441,N_26117);
and U26600 (N_26600,N_26115,N_26157);
xnor U26601 (N_26601,N_26348,N_26273);
and U26602 (N_26602,N_26052,N_26004);
xnor U26603 (N_26603,N_26414,N_26378);
nor U26604 (N_26604,N_26310,N_26459);
or U26605 (N_26605,N_26274,N_26024);
nor U26606 (N_26606,N_26324,N_26393);
nand U26607 (N_26607,N_26492,N_26462);
xor U26608 (N_26608,N_26045,N_26361);
xor U26609 (N_26609,N_26077,N_26331);
xor U26610 (N_26610,N_26167,N_26490);
nand U26611 (N_26611,N_26130,N_26298);
or U26612 (N_26612,N_26020,N_26146);
nand U26613 (N_26613,N_26206,N_26144);
nand U26614 (N_26614,N_26419,N_26118);
nand U26615 (N_26615,N_26235,N_26208);
nor U26616 (N_26616,N_26033,N_26357);
nand U26617 (N_26617,N_26372,N_26290);
or U26618 (N_26618,N_26073,N_26313);
nor U26619 (N_26619,N_26229,N_26007);
or U26620 (N_26620,N_26297,N_26106);
xnor U26621 (N_26621,N_26029,N_26129);
and U26622 (N_26622,N_26189,N_26035);
nor U26623 (N_26623,N_26373,N_26176);
nand U26624 (N_26624,N_26151,N_26272);
nand U26625 (N_26625,N_26365,N_26493);
nand U26626 (N_26626,N_26083,N_26047);
xor U26627 (N_26627,N_26281,N_26480);
or U26628 (N_26628,N_26075,N_26212);
xnor U26629 (N_26629,N_26477,N_26354);
nor U26630 (N_26630,N_26113,N_26410);
and U26631 (N_26631,N_26385,N_26415);
nor U26632 (N_26632,N_26112,N_26420);
nor U26633 (N_26633,N_26237,N_26470);
xnor U26634 (N_26634,N_26032,N_26450);
nor U26635 (N_26635,N_26063,N_26236);
nor U26636 (N_26636,N_26287,N_26307);
xor U26637 (N_26637,N_26250,N_26119);
nor U26638 (N_26638,N_26246,N_26152);
nand U26639 (N_26639,N_26039,N_26110);
xnor U26640 (N_26640,N_26203,N_26260);
and U26641 (N_26641,N_26050,N_26263);
or U26642 (N_26642,N_26380,N_26379);
or U26643 (N_26643,N_26330,N_26240);
and U26644 (N_26644,N_26166,N_26164);
and U26645 (N_26645,N_26121,N_26245);
xor U26646 (N_26646,N_26368,N_26201);
xnor U26647 (N_26647,N_26234,N_26284);
and U26648 (N_26648,N_26305,N_26162);
or U26649 (N_26649,N_26027,N_26216);
and U26650 (N_26650,N_26285,N_26466);
nor U26651 (N_26651,N_26309,N_26386);
nand U26652 (N_26652,N_26173,N_26156);
nand U26653 (N_26653,N_26295,N_26138);
or U26654 (N_26654,N_26013,N_26178);
or U26655 (N_26655,N_26022,N_26232);
xnor U26656 (N_26656,N_26347,N_26321);
xor U26657 (N_26657,N_26497,N_26353);
nand U26658 (N_26658,N_26220,N_26198);
nor U26659 (N_26659,N_26424,N_26280);
nor U26660 (N_26660,N_26389,N_26231);
or U26661 (N_26661,N_26423,N_26079);
nand U26662 (N_26662,N_26275,N_26289);
nand U26663 (N_26663,N_26127,N_26134);
or U26664 (N_26664,N_26395,N_26163);
nor U26665 (N_26665,N_26067,N_26037);
and U26666 (N_26666,N_26018,N_26483);
xor U26667 (N_26667,N_26267,N_26252);
and U26668 (N_26668,N_26195,N_26222);
nor U26669 (N_26669,N_26025,N_26149);
or U26670 (N_26670,N_26103,N_26400);
and U26671 (N_26671,N_26191,N_26031);
and U26672 (N_26672,N_26095,N_26447);
or U26673 (N_26673,N_26308,N_26412);
nor U26674 (N_26674,N_26482,N_26093);
or U26675 (N_26675,N_26028,N_26352);
and U26676 (N_26676,N_26433,N_26481);
nand U26677 (N_26677,N_26261,N_26219);
nand U26678 (N_26678,N_26264,N_26213);
nand U26679 (N_26679,N_26431,N_26038);
nand U26680 (N_26680,N_26461,N_26383);
or U26681 (N_26681,N_26011,N_26089);
xnor U26682 (N_26682,N_26012,N_26000);
or U26683 (N_26683,N_26469,N_26049);
and U26684 (N_26684,N_26019,N_26332);
nand U26685 (N_26685,N_26174,N_26053);
nor U26686 (N_26686,N_26199,N_26306);
or U26687 (N_26687,N_26087,N_26366);
nor U26688 (N_26688,N_26404,N_26192);
xor U26689 (N_26689,N_26271,N_26346);
nand U26690 (N_26690,N_26085,N_26376);
nand U26691 (N_26691,N_26425,N_26060);
nor U26692 (N_26692,N_26460,N_26044);
and U26693 (N_26693,N_26344,N_26350);
xor U26694 (N_26694,N_26338,N_26061);
nor U26695 (N_26695,N_26168,N_26406);
nor U26696 (N_26696,N_26243,N_26188);
nand U26697 (N_26697,N_26056,N_26325);
xnor U26698 (N_26698,N_26437,N_26193);
xnor U26699 (N_26699,N_26405,N_26209);
nand U26700 (N_26700,N_26248,N_26458);
nor U26701 (N_26701,N_26371,N_26116);
nor U26702 (N_26702,N_26370,N_26403);
xor U26703 (N_26703,N_26475,N_26265);
nand U26704 (N_26704,N_26456,N_26259);
xnor U26705 (N_26705,N_26337,N_26107);
xnor U26706 (N_26706,N_26137,N_26015);
nor U26707 (N_26707,N_26487,N_26392);
xnor U26708 (N_26708,N_26381,N_26202);
xnor U26709 (N_26709,N_26270,N_26100);
and U26710 (N_26710,N_26021,N_26026);
or U26711 (N_26711,N_26158,N_26124);
xnor U26712 (N_26712,N_26241,N_26097);
nand U26713 (N_26713,N_26036,N_26300);
nand U26714 (N_26714,N_26430,N_26224);
or U26715 (N_26715,N_26242,N_26254);
or U26716 (N_26716,N_26170,N_26478);
and U26717 (N_26717,N_26183,N_26154);
nor U26718 (N_26718,N_26010,N_26185);
and U26719 (N_26719,N_26443,N_26005);
xor U26720 (N_26720,N_26327,N_26181);
or U26721 (N_26721,N_26105,N_26023);
xor U26722 (N_26722,N_26413,N_26495);
nor U26723 (N_26723,N_26016,N_26436);
and U26724 (N_26724,N_26262,N_26165);
xnor U26725 (N_26725,N_26255,N_26204);
nor U26726 (N_26726,N_26177,N_26205);
and U26727 (N_26727,N_26098,N_26210);
and U26728 (N_26728,N_26446,N_26444);
and U26729 (N_26729,N_26402,N_26180);
xor U26730 (N_26730,N_26244,N_26328);
and U26731 (N_26731,N_26374,N_26128);
nor U26732 (N_26732,N_26215,N_26042);
nand U26733 (N_26733,N_26090,N_26094);
and U26734 (N_26734,N_26046,N_26190);
and U26735 (N_26735,N_26186,N_26453);
nand U26736 (N_26736,N_26359,N_26040);
xor U26737 (N_26737,N_26369,N_26122);
and U26738 (N_26738,N_26135,N_26082);
nor U26739 (N_26739,N_26417,N_26194);
xnor U26740 (N_26740,N_26409,N_26474);
and U26741 (N_26741,N_26319,N_26096);
nor U26742 (N_26742,N_26125,N_26187);
and U26743 (N_26743,N_26148,N_26421);
and U26744 (N_26744,N_26001,N_26228);
and U26745 (N_26745,N_26282,N_26390);
xor U26746 (N_26746,N_26399,N_26472);
nand U26747 (N_26747,N_26091,N_26326);
and U26748 (N_26748,N_26140,N_26418);
or U26749 (N_26749,N_26066,N_26247);
nor U26750 (N_26750,N_26480,N_26185);
xor U26751 (N_26751,N_26059,N_26203);
xor U26752 (N_26752,N_26359,N_26070);
nand U26753 (N_26753,N_26374,N_26176);
nor U26754 (N_26754,N_26314,N_26169);
or U26755 (N_26755,N_26307,N_26251);
nand U26756 (N_26756,N_26007,N_26043);
xor U26757 (N_26757,N_26145,N_26323);
xor U26758 (N_26758,N_26472,N_26341);
or U26759 (N_26759,N_26075,N_26087);
xor U26760 (N_26760,N_26424,N_26064);
nor U26761 (N_26761,N_26478,N_26041);
nor U26762 (N_26762,N_26232,N_26483);
nor U26763 (N_26763,N_26444,N_26386);
xnor U26764 (N_26764,N_26383,N_26329);
and U26765 (N_26765,N_26418,N_26362);
and U26766 (N_26766,N_26057,N_26436);
or U26767 (N_26767,N_26350,N_26236);
nor U26768 (N_26768,N_26285,N_26067);
nand U26769 (N_26769,N_26265,N_26435);
or U26770 (N_26770,N_26417,N_26418);
and U26771 (N_26771,N_26431,N_26122);
nor U26772 (N_26772,N_26092,N_26444);
nand U26773 (N_26773,N_26310,N_26353);
and U26774 (N_26774,N_26418,N_26320);
nor U26775 (N_26775,N_26004,N_26107);
or U26776 (N_26776,N_26473,N_26134);
nand U26777 (N_26777,N_26376,N_26214);
nor U26778 (N_26778,N_26248,N_26168);
nor U26779 (N_26779,N_26400,N_26057);
nor U26780 (N_26780,N_26378,N_26099);
nor U26781 (N_26781,N_26137,N_26226);
and U26782 (N_26782,N_26253,N_26496);
or U26783 (N_26783,N_26459,N_26142);
or U26784 (N_26784,N_26360,N_26266);
or U26785 (N_26785,N_26384,N_26018);
or U26786 (N_26786,N_26259,N_26010);
and U26787 (N_26787,N_26029,N_26437);
nand U26788 (N_26788,N_26226,N_26223);
and U26789 (N_26789,N_26418,N_26238);
or U26790 (N_26790,N_26331,N_26266);
xor U26791 (N_26791,N_26425,N_26193);
nand U26792 (N_26792,N_26247,N_26485);
xor U26793 (N_26793,N_26191,N_26426);
nor U26794 (N_26794,N_26006,N_26325);
and U26795 (N_26795,N_26001,N_26213);
nand U26796 (N_26796,N_26218,N_26022);
nand U26797 (N_26797,N_26226,N_26062);
xnor U26798 (N_26798,N_26310,N_26024);
nor U26799 (N_26799,N_26422,N_26074);
xor U26800 (N_26800,N_26464,N_26497);
nand U26801 (N_26801,N_26377,N_26232);
xor U26802 (N_26802,N_26024,N_26238);
nand U26803 (N_26803,N_26475,N_26487);
xor U26804 (N_26804,N_26220,N_26372);
or U26805 (N_26805,N_26010,N_26029);
nor U26806 (N_26806,N_26008,N_26298);
nand U26807 (N_26807,N_26144,N_26337);
xnor U26808 (N_26808,N_26364,N_26020);
and U26809 (N_26809,N_26177,N_26054);
nand U26810 (N_26810,N_26165,N_26101);
xor U26811 (N_26811,N_26499,N_26445);
nand U26812 (N_26812,N_26134,N_26208);
nor U26813 (N_26813,N_26178,N_26089);
xor U26814 (N_26814,N_26494,N_26163);
nand U26815 (N_26815,N_26361,N_26093);
nand U26816 (N_26816,N_26247,N_26232);
nor U26817 (N_26817,N_26364,N_26060);
or U26818 (N_26818,N_26340,N_26044);
nand U26819 (N_26819,N_26060,N_26203);
nor U26820 (N_26820,N_26481,N_26460);
and U26821 (N_26821,N_26456,N_26248);
xnor U26822 (N_26822,N_26191,N_26154);
nand U26823 (N_26823,N_26284,N_26013);
nor U26824 (N_26824,N_26450,N_26106);
xor U26825 (N_26825,N_26466,N_26458);
and U26826 (N_26826,N_26340,N_26259);
nor U26827 (N_26827,N_26197,N_26236);
nor U26828 (N_26828,N_26145,N_26013);
or U26829 (N_26829,N_26363,N_26021);
nand U26830 (N_26830,N_26333,N_26238);
nand U26831 (N_26831,N_26211,N_26038);
nand U26832 (N_26832,N_26499,N_26393);
and U26833 (N_26833,N_26415,N_26437);
and U26834 (N_26834,N_26234,N_26296);
and U26835 (N_26835,N_26251,N_26488);
nor U26836 (N_26836,N_26350,N_26289);
nand U26837 (N_26837,N_26452,N_26002);
nor U26838 (N_26838,N_26010,N_26224);
xor U26839 (N_26839,N_26013,N_26204);
nand U26840 (N_26840,N_26039,N_26222);
or U26841 (N_26841,N_26231,N_26258);
nor U26842 (N_26842,N_26398,N_26146);
nor U26843 (N_26843,N_26366,N_26216);
nand U26844 (N_26844,N_26012,N_26249);
nor U26845 (N_26845,N_26065,N_26402);
xnor U26846 (N_26846,N_26244,N_26137);
nand U26847 (N_26847,N_26156,N_26259);
nor U26848 (N_26848,N_26433,N_26365);
nor U26849 (N_26849,N_26264,N_26437);
and U26850 (N_26850,N_26437,N_26365);
nand U26851 (N_26851,N_26097,N_26413);
nor U26852 (N_26852,N_26014,N_26184);
or U26853 (N_26853,N_26043,N_26460);
nor U26854 (N_26854,N_26286,N_26407);
or U26855 (N_26855,N_26418,N_26342);
or U26856 (N_26856,N_26402,N_26324);
or U26857 (N_26857,N_26476,N_26051);
xnor U26858 (N_26858,N_26395,N_26124);
xnor U26859 (N_26859,N_26171,N_26367);
nand U26860 (N_26860,N_26153,N_26189);
xnor U26861 (N_26861,N_26341,N_26351);
and U26862 (N_26862,N_26062,N_26158);
nand U26863 (N_26863,N_26372,N_26016);
xor U26864 (N_26864,N_26031,N_26371);
nor U26865 (N_26865,N_26137,N_26312);
nand U26866 (N_26866,N_26303,N_26459);
xor U26867 (N_26867,N_26100,N_26302);
and U26868 (N_26868,N_26440,N_26406);
or U26869 (N_26869,N_26134,N_26395);
nor U26870 (N_26870,N_26265,N_26080);
nor U26871 (N_26871,N_26001,N_26118);
xnor U26872 (N_26872,N_26341,N_26172);
xor U26873 (N_26873,N_26376,N_26299);
or U26874 (N_26874,N_26255,N_26478);
xnor U26875 (N_26875,N_26234,N_26329);
nor U26876 (N_26876,N_26432,N_26336);
nor U26877 (N_26877,N_26057,N_26198);
xor U26878 (N_26878,N_26226,N_26025);
and U26879 (N_26879,N_26165,N_26138);
nor U26880 (N_26880,N_26227,N_26241);
nor U26881 (N_26881,N_26210,N_26291);
nand U26882 (N_26882,N_26113,N_26091);
or U26883 (N_26883,N_26439,N_26352);
and U26884 (N_26884,N_26465,N_26228);
xor U26885 (N_26885,N_26494,N_26301);
nand U26886 (N_26886,N_26386,N_26301);
nor U26887 (N_26887,N_26207,N_26244);
xnor U26888 (N_26888,N_26495,N_26134);
nand U26889 (N_26889,N_26127,N_26028);
nand U26890 (N_26890,N_26456,N_26100);
xor U26891 (N_26891,N_26390,N_26289);
xor U26892 (N_26892,N_26011,N_26154);
nor U26893 (N_26893,N_26255,N_26496);
or U26894 (N_26894,N_26000,N_26133);
nor U26895 (N_26895,N_26308,N_26457);
nand U26896 (N_26896,N_26406,N_26206);
xnor U26897 (N_26897,N_26029,N_26136);
nor U26898 (N_26898,N_26220,N_26457);
nor U26899 (N_26899,N_26493,N_26151);
nor U26900 (N_26900,N_26021,N_26047);
xnor U26901 (N_26901,N_26395,N_26227);
and U26902 (N_26902,N_26153,N_26011);
nand U26903 (N_26903,N_26420,N_26311);
nor U26904 (N_26904,N_26444,N_26053);
and U26905 (N_26905,N_26086,N_26361);
or U26906 (N_26906,N_26115,N_26081);
nor U26907 (N_26907,N_26393,N_26167);
nor U26908 (N_26908,N_26294,N_26238);
nor U26909 (N_26909,N_26060,N_26267);
nor U26910 (N_26910,N_26040,N_26241);
nor U26911 (N_26911,N_26127,N_26453);
xnor U26912 (N_26912,N_26060,N_26254);
nor U26913 (N_26913,N_26206,N_26111);
xnor U26914 (N_26914,N_26276,N_26233);
nand U26915 (N_26915,N_26116,N_26305);
xor U26916 (N_26916,N_26052,N_26132);
nand U26917 (N_26917,N_26480,N_26357);
nor U26918 (N_26918,N_26030,N_26002);
nor U26919 (N_26919,N_26302,N_26458);
nand U26920 (N_26920,N_26044,N_26041);
xor U26921 (N_26921,N_26471,N_26414);
nor U26922 (N_26922,N_26115,N_26452);
or U26923 (N_26923,N_26450,N_26387);
and U26924 (N_26924,N_26140,N_26015);
and U26925 (N_26925,N_26423,N_26100);
nor U26926 (N_26926,N_26249,N_26381);
xnor U26927 (N_26927,N_26481,N_26327);
nor U26928 (N_26928,N_26050,N_26247);
and U26929 (N_26929,N_26439,N_26270);
xnor U26930 (N_26930,N_26194,N_26447);
nand U26931 (N_26931,N_26376,N_26379);
nand U26932 (N_26932,N_26434,N_26427);
and U26933 (N_26933,N_26447,N_26342);
and U26934 (N_26934,N_26116,N_26123);
nor U26935 (N_26935,N_26383,N_26458);
nor U26936 (N_26936,N_26126,N_26223);
and U26937 (N_26937,N_26294,N_26322);
or U26938 (N_26938,N_26109,N_26238);
nand U26939 (N_26939,N_26060,N_26295);
and U26940 (N_26940,N_26013,N_26158);
or U26941 (N_26941,N_26317,N_26469);
or U26942 (N_26942,N_26496,N_26314);
and U26943 (N_26943,N_26405,N_26196);
and U26944 (N_26944,N_26184,N_26433);
nor U26945 (N_26945,N_26324,N_26291);
nor U26946 (N_26946,N_26414,N_26446);
or U26947 (N_26947,N_26402,N_26190);
nand U26948 (N_26948,N_26143,N_26011);
nand U26949 (N_26949,N_26080,N_26183);
nand U26950 (N_26950,N_26323,N_26398);
nand U26951 (N_26951,N_26139,N_26148);
nor U26952 (N_26952,N_26260,N_26442);
or U26953 (N_26953,N_26002,N_26126);
and U26954 (N_26954,N_26073,N_26164);
or U26955 (N_26955,N_26434,N_26415);
nand U26956 (N_26956,N_26249,N_26475);
nand U26957 (N_26957,N_26068,N_26145);
nor U26958 (N_26958,N_26237,N_26360);
xnor U26959 (N_26959,N_26102,N_26045);
nor U26960 (N_26960,N_26454,N_26278);
nand U26961 (N_26961,N_26093,N_26247);
nand U26962 (N_26962,N_26418,N_26368);
or U26963 (N_26963,N_26043,N_26357);
and U26964 (N_26964,N_26194,N_26109);
or U26965 (N_26965,N_26310,N_26232);
nor U26966 (N_26966,N_26023,N_26147);
xor U26967 (N_26967,N_26329,N_26237);
and U26968 (N_26968,N_26440,N_26305);
nand U26969 (N_26969,N_26488,N_26213);
nand U26970 (N_26970,N_26266,N_26212);
xor U26971 (N_26971,N_26468,N_26404);
xor U26972 (N_26972,N_26124,N_26355);
or U26973 (N_26973,N_26444,N_26372);
nor U26974 (N_26974,N_26424,N_26115);
nor U26975 (N_26975,N_26349,N_26285);
and U26976 (N_26976,N_26444,N_26254);
and U26977 (N_26977,N_26423,N_26153);
nor U26978 (N_26978,N_26150,N_26477);
nor U26979 (N_26979,N_26319,N_26396);
nor U26980 (N_26980,N_26465,N_26200);
and U26981 (N_26981,N_26102,N_26088);
nor U26982 (N_26982,N_26102,N_26252);
nand U26983 (N_26983,N_26433,N_26499);
nand U26984 (N_26984,N_26413,N_26090);
and U26985 (N_26985,N_26158,N_26192);
nand U26986 (N_26986,N_26291,N_26221);
xor U26987 (N_26987,N_26036,N_26070);
nand U26988 (N_26988,N_26449,N_26489);
nor U26989 (N_26989,N_26435,N_26438);
and U26990 (N_26990,N_26261,N_26059);
and U26991 (N_26991,N_26310,N_26474);
and U26992 (N_26992,N_26198,N_26358);
xor U26993 (N_26993,N_26074,N_26377);
nor U26994 (N_26994,N_26353,N_26184);
xor U26995 (N_26995,N_26385,N_26344);
xnor U26996 (N_26996,N_26488,N_26288);
nor U26997 (N_26997,N_26347,N_26463);
or U26998 (N_26998,N_26342,N_26242);
xnor U26999 (N_26999,N_26161,N_26216);
nand U27000 (N_27000,N_26618,N_26701);
and U27001 (N_27001,N_26865,N_26646);
nor U27002 (N_27002,N_26539,N_26657);
xnor U27003 (N_27003,N_26891,N_26585);
xor U27004 (N_27004,N_26830,N_26674);
or U27005 (N_27005,N_26906,N_26981);
xnor U27006 (N_27006,N_26792,N_26856);
xor U27007 (N_27007,N_26999,N_26630);
nand U27008 (N_27008,N_26864,N_26968);
nor U27009 (N_27009,N_26652,N_26501);
and U27010 (N_27010,N_26880,N_26500);
nor U27011 (N_27011,N_26598,N_26606);
and U27012 (N_27012,N_26791,N_26963);
xor U27013 (N_27013,N_26793,N_26971);
and U27014 (N_27014,N_26945,N_26928);
nand U27015 (N_27015,N_26577,N_26680);
and U27016 (N_27016,N_26907,N_26746);
nand U27017 (N_27017,N_26867,N_26751);
nand U27018 (N_27018,N_26616,N_26862);
and U27019 (N_27019,N_26878,N_26550);
or U27020 (N_27020,N_26825,N_26507);
or U27021 (N_27021,N_26816,N_26578);
and U27022 (N_27022,N_26765,N_26782);
or U27023 (N_27023,N_26540,N_26957);
nand U27024 (N_27024,N_26951,N_26892);
and U27025 (N_27025,N_26966,N_26715);
or U27026 (N_27026,N_26883,N_26575);
or U27027 (N_27027,N_26557,N_26595);
nor U27028 (N_27028,N_26534,N_26528);
xnor U27029 (N_27029,N_26953,N_26978);
nor U27030 (N_27030,N_26609,N_26817);
xor U27031 (N_27031,N_26572,N_26529);
xnor U27032 (N_27032,N_26622,N_26705);
or U27033 (N_27033,N_26837,N_26810);
nand U27034 (N_27034,N_26863,N_26836);
and U27035 (N_27035,N_26697,N_26689);
or U27036 (N_27036,N_26502,N_26513);
xnor U27037 (N_27037,N_26904,N_26738);
xor U27038 (N_27038,N_26620,N_26667);
or U27039 (N_27039,N_26624,N_26911);
or U27040 (N_27040,N_26954,N_26861);
xor U27041 (N_27041,N_26613,N_26794);
and U27042 (N_27042,N_26656,N_26619);
and U27043 (N_27043,N_26716,N_26744);
and U27044 (N_27044,N_26859,N_26986);
and U27045 (N_27045,N_26987,N_26920);
and U27046 (N_27046,N_26972,N_26617);
xnor U27047 (N_27047,N_26860,N_26602);
nor U27048 (N_27048,N_26506,N_26714);
nand U27049 (N_27049,N_26665,N_26866);
xor U27050 (N_27050,N_26787,N_26958);
and U27051 (N_27051,N_26903,N_26541);
nand U27052 (N_27052,N_26873,N_26815);
nand U27053 (N_27053,N_26976,N_26589);
nor U27054 (N_27054,N_26583,N_26879);
nand U27055 (N_27055,N_26722,N_26661);
and U27056 (N_27056,N_26902,N_26658);
or U27057 (N_27057,N_26611,N_26962);
nor U27058 (N_27058,N_26659,N_26641);
nor U27059 (N_27059,N_26594,N_26605);
xor U27060 (N_27060,N_26875,N_26844);
or U27061 (N_27061,N_26764,N_26566);
nand U27062 (N_27062,N_26635,N_26779);
nand U27063 (N_27063,N_26579,N_26947);
nor U27064 (N_27064,N_26930,N_26530);
nand U27065 (N_27065,N_26668,N_26973);
nand U27066 (N_27066,N_26993,N_26524);
nor U27067 (N_27067,N_26766,N_26802);
xnor U27068 (N_27068,N_26762,N_26559);
xor U27069 (N_27069,N_26974,N_26789);
xor U27070 (N_27070,N_26803,N_26564);
nor U27071 (N_27071,N_26581,N_26670);
xor U27072 (N_27072,N_26832,N_26702);
xnor U27073 (N_27073,N_26678,N_26704);
and U27074 (N_27074,N_26874,N_26869);
and U27075 (N_27075,N_26743,N_26654);
nand U27076 (N_27076,N_26742,N_26767);
xor U27077 (N_27077,N_26568,N_26621);
or U27078 (N_27078,N_26956,N_26600);
and U27079 (N_27079,N_26982,N_26587);
nand U27080 (N_27080,N_26948,N_26852);
or U27081 (N_27081,N_26774,N_26690);
or U27082 (N_27082,N_26756,N_26666);
or U27083 (N_27083,N_26887,N_26545);
nor U27084 (N_27084,N_26515,N_26912);
xnor U27085 (N_27085,N_26748,N_26649);
or U27086 (N_27086,N_26770,N_26626);
nor U27087 (N_27087,N_26687,N_26809);
xor U27088 (N_27088,N_26822,N_26675);
nor U27089 (N_27089,N_26845,N_26709);
or U27090 (N_27090,N_26854,N_26660);
nor U27091 (N_27091,N_26796,N_26644);
and U27092 (N_27092,N_26995,N_26551);
and U27093 (N_27093,N_26959,N_26970);
xor U27094 (N_27094,N_26939,N_26848);
nand U27095 (N_27095,N_26706,N_26824);
xnor U27096 (N_27096,N_26908,N_26538);
and U27097 (N_27097,N_26596,N_26745);
xnor U27098 (N_27098,N_26698,N_26576);
xnor U27099 (N_27099,N_26521,N_26897);
nor U27100 (N_27100,N_26691,N_26719);
xor U27101 (N_27101,N_26607,N_26749);
or U27102 (N_27102,N_26610,N_26943);
nand U27103 (N_27103,N_26909,N_26727);
nand U27104 (N_27104,N_26553,N_26946);
nand U27105 (N_27105,N_26663,N_26855);
xor U27106 (N_27106,N_26634,N_26707);
nor U27107 (N_27107,N_26898,N_26812);
and U27108 (N_27108,N_26673,N_26664);
nand U27109 (N_27109,N_26662,N_26868);
or U27110 (N_27110,N_26843,N_26808);
xor U27111 (N_27111,N_26893,N_26542);
nand U27112 (N_27112,N_26795,N_26776);
or U27113 (N_27113,N_26916,N_26643);
or U27114 (N_27114,N_26653,N_26571);
and U27115 (N_27115,N_26952,N_26710);
nor U27116 (N_27116,N_26556,N_26877);
nand U27117 (N_27117,N_26728,N_26633);
and U27118 (N_27118,N_26771,N_26931);
and U27119 (N_27119,N_26682,N_26516);
and U27120 (N_27120,N_26693,N_26934);
or U27121 (N_27121,N_26736,N_26784);
or U27122 (N_27122,N_26631,N_26536);
nor U27123 (N_27123,N_26900,N_26980);
xor U27124 (N_27124,N_26990,N_26526);
xnor U27125 (N_27125,N_26798,N_26828);
or U27126 (N_27126,N_26692,N_26872);
xor U27127 (N_27127,N_26944,N_26758);
nand U27128 (N_27128,N_26615,N_26735);
xor U27129 (N_27129,N_26820,N_26881);
or U27130 (N_27130,N_26681,N_26555);
nand U27131 (N_27131,N_26558,N_26679);
nor U27132 (N_27132,N_26781,N_26601);
xnor U27133 (N_27133,N_26938,N_26785);
xnor U27134 (N_27134,N_26642,N_26713);
or U27135 (N_27135,N_26807,N_26942);
nor U27136 (N_27136,N_26905,N_26819);
xnor U27137 (N_27137,N_26842,N_26741);
nor U27138 (N_27138,N_26591,N_26997);
nand U27139 (N_27139,N_26772,N_26512);
nand U27140 (N_27140,N_26737,N_26780);
and U27141 (N_27141,N_26531,N_26778);
and U27142 (N_27142,N_26546,N_26645);
xnor U27143 (N_27143,N_26969,N_26923);
and U27144 (N_27144,N_26632,N_26975);
nand U27145 (N_27145,N_26783,N_26732);
xnor U27146 (N_27146,N_26629,N_26569);
or U27147 (N_27147,N_26851,N_26965);
or U27148 (N_27148,N_26608,N_26818);
nand U27149 (N_27149,N_26739,N_26805);
or U27150 (N_27150,N_26740,N_26926);
xnor U27151 (N_27151,N_26763,N_26977);
nor U27152 (N_27152,N_26899,N_26929);
nor U27153 (N_27153,N_26655,N_26989);
xnor U27154 (N_27154,N_26543,N_26597);
or U27155 (N_27155,N_26549,N_26720);
nor U27156 (N_27156,N_26806,N_26669);
nor U27157 (N_27157,N_26850,N_26777);
or U27158 (N_27158,N_26725,N_26733);
nor U27159 (N_27159,N_26623,N_26588);
xnor U27160 (N_27160,N_26677,N_26533);
or U27161 (N_27161,N_26554,N_26671);
xnor U27162 (N_27162,N_26979,N_26518);
or U27163 (N_27163,N_26901,N_26857);
and U27164 (N_27164,N_26650,N_26580);
and U27165 (N_27165,N_26888,N_26582);
nand U27166 (N_27166,N_26695,N_26603);
nor U27167 (N_27167,N_26961,N_26636);
xor U27168 (N_27168,N_26846,N_26940);
nand U27169 (N_27169,N_26984,N_26853);
or U27170 (N_27170,N_26941,N_26520);
nand U27171 (N_27171,N_26730,N_26639);
and U27172 (N_27172,N_26834,N_26552);
or U27173 (N_27173,N_26648,N_26996);
xor U27174 (N_27174,N_26734,N_26922);
nor U27175 (N_27175,N_26882,N_26858);
nand U27176 (N_27176,N_26884,N_26933);
and U27177 (N_27177,N_26827,N_26769);
xnor U27178 (N_27178,N_26685,N_26960);
and U27179 (N_27179,N_26625,N_26768);
nand U27180 (N_27180,N_26889,N_26988);
xor U27181 (N_27181,N_26752,N_26573);
xnor U27182 (N_27182,N_26829,N_26804);
nand U27183 (N_27183,N_26786,N_26921);
xnor U27184 (N_27184,N_26895,N_26561);
and U27185 (N_27185,N_26567,N_26686);
nor U27186 (N_27186,N_26932,N_26915);
nand U27187 (N_27187,N_26994,N_26522);
nand U27188 (N_27188,N_26731,N_26544);
nor U27189 (N_27189,N_26599,N_26985);
nand U27190 (N_27190,N_26992,N_26560);
nand U27191 (N_27191,N_26797,N_26724);
xnor U27192 (N_27192,N_26627,N_26562);
nor U27193 (N_27193,N_26755,N_26509);
nor U27194 (N_27194,N_26894,N_26950);
xor U27195 (N_27195,N_26592,N_26750);
nor U27196 (N_27196,N_26801,N_26517);
and U27197 (N_27197,N_26910,N_26532);
xnor U27198 (N_27198,N_26918,N_26676);
or U27199 (N_27199,N_26925,N_26699);
nand U27200 (N_27200,N_26723,N_26504);
xor U27201 (N_27201,N_26590,N_26565);
nand U27202 (N_27202,N_26647,N_26628);
and U27203 (N_27203,N_26831,N_26913);
nand U27204 (N_27204,N_26964,N_26505);
and U27205 (N_27205,N_26563,N_26840);
nand U27206 (N_27206,N_26708,N_26638);
and U27207 (N_27207,N_26510,N_26890);
nor U27208 (N_27208,N_26514,N_26841);
nor U27209 (N_27209,N_26593,N_26800);
nand U27210 (N_27210,N_26811,N_26760);
nand U27211 (N_27211,N_26503,N_26604);
xnor U27212 (N_27212,N_26790,N_26523);
or U27213 (N_27213,N_26729,N_26935);
xnor U27214 (N_27214,N_26721,N_26821);
xor U27215 (N_27215,N_26547,N_26788);
nand U27216 (N_27216,N_26871,N_26773);
nand U27217 (N_27217,N_26936,N_26927);
nor U27218 (N_27218,N_26839,N_26937);
nor U27219 (N_27219,N_26833,N_26525);
nand U27220 (N_27220,N_26949,N_26684);
nor U27221 (N_27221,N_26726,N_26703);
or U27222 (N_27222,N_26876,N_26847);
and U27223 (N_27223,N_26640,N_26574);
or U27224 (N_27224,N_26637,N_26519);
nand U27225 (N_27225,N_26511,N_26955);
and U27226 (N_27226,N_26508,N_26570);
and U27227 (N_27227,N_26917,N_26761);
nand U27228 (N_27228,N_26718,N_26688);
nor U27229 (N_27229,N_26823,N_26919);
and U27230 (N_27230,N_26983,N_26754);
nand U27231 (N_27231,N_26548,N_26694);
nand U27232 (N_27232,N_26991,N_26813);
and U27233 (N_27233,N_26914,N_26757);
xnor U27234 (N_27234,N_26535,N_26967);
nor U27235 (N_27235,N_26886,N_26683);
nor U27236 (N_27236,N_26838,N_26799);
nand U27237 (N_27237,N_26651,N_26826);
nand U27238 (N_27238,N_26896,N_26814);
and U27239 (N_27239,N_26924,N_26717);
and U27240 (N_27240,N_26998,N_26870);
xnor U27241 (N_27241,N_26747,N_26711);
xnor U27242 (N_27242,N_26775,N_26672);
or U27243 (N_27243,N_26849,N_26835);
nand U27244 (N_27244,N_26586,N_26584);
nand U27245 (N_27245,N_26696,N_26753);
nor U27246 (N_27246,N_26885,N_26614);
and U27247 (N_27247,N_26700,N_26759);
xor U27248 (N_27248,N_26527,N_26712);
xor U27249 (N_27249,N_26537,N_26612);
or U27250 (N_27250,N_26642,N_26857);
nor U27251 (N_27251,N_26963,N_26767);
xor U27252 (N_27252,N_26932,N_26990);
nand U27253 (N_27253,N_26840,N_26539);
xnor U27254 (N_27254,N_26963,N_26940);
or U27255 (N_27255,N_26992,N_26653);
xnor U27256 (N_27256,N_26612,N_26619);
or U27257 (N_27257,N_26606,N_26974);
nor U27258 (N_27258,N_26731,N_26667);
nor U27259 (N_27259,N_26524,N_26945);
nand U27260 (N_27260,N_26811,N_26780);
xnor U27261 (N_27261,N_26510,N_26934);
nor U27262 (N_27262,N_26854,N_26631);
xor U27263 (N_27263,N_26659,N_26952);
or U27264 (N_27264,N_26717,N_26750);
and U27265 (N_27265,N_26732,N_26594);
nand U27266 (N_27266,N_26821,N_26661);
xor U27267 (N_27267,N_26745,N_26914);
or U27268 (N_27268,N_26797,N_26690);
xor U27269 (N_27269,N_26687,N_26662);
nor U27270 (N_27270,N_26798,N_26573);
nand U27271 (N_27271,N_26711,N_26505);
and U27272 (N_27272,N_26521,N_26701);
or U27273 (N_27273,N_26940,N_26977);
and U27274 (N_27274,N_26963,N_26824);
nand U27275 (N_27275,N_26559,N_26672);
nand U27276 (N_27276,N_26598,N_26522);
or U27277 (N_27277,N_26827,N_26860);
nand U27278 (N_27278,N_26846,N_26821);
nor U27279 (N_27279,N_26656,N_26626);
and U27280 (N_27280,N_26810,N_26864);
xnor U27281 (N_27281,N_26612,N_26601);
nor U27282 (N_27282,N_26642,N_26911);
or U27283 (N_27283,N_26720,N_26523);
and U27284 (N_27284,N_26622,N_26512);
nand U27285 (N_27285,N_26570,N_26857);
or U27286 (N_27286,N_26797,N_26632);
or U27287 (N_27287,N_26595,N_26846);
nor U27288 (N_27288,N_26594,N_26868);
nand U27289 (N_27289,N_26963,N_26560);
nor U27290 (N_27290,N_26553,N_26784);
nand U27291 (N_27291,N_26787,N_26885);
xnor U27292 (N_27292,N_26946,N_26710);
nor U27293 (N_27293,N_26902,N_26779);
nor U27294 (N_27294,N_26688,N_26533);
xor U27295 (N_27295,N_26516,N_26659);
nand U27296 (N_27296,N_26850,N_26948);
nand U27297 (N_27297,N_26980,N_26732);
nand U27298 (N_27298,N_26552,N_26768);
xnor U27299 (N_27299,N_26675,N_26866);
or U27300 (N_27300,N_26836,N_26795);
or U27301 (N_27301,N_26998,N_26824);
xor U27302 (N_27302,N_26606,N_26896);
xor U27303 (N_27303,N_26814,N_26500);
xor U27304 (N_27304,N_26591,N_26530);
nor U27305 (N_27305,N_26542,N_26706);
nand U27306 (N_27306,N_26817,N_26811);
xor U27307 (N_27307,N_26839,N_26806);
nand U27308 (N_27308,N_26534,N_26775);
and U27309 (N_27309,N_26546,N_26587);
nor U27310 (N_27310,N_26924,N_26606);
and U27311 (N_27311,N_26538,N_26787);
nor U27312 (N_27312,N_26863,N_26927);
or U27313 (N_27313,N_26827,N_26765);
nor U27314 (N_27314,N_26538,N_26900);
or U27315 (N_27315,N_26588,N_26997);
or U27316 (N_27316,N_26835,N_26708);
or U27317 (N_27317,N_26622,N_26598);
or U27318 (N_27318,N_26697,N_26510);
xnor U27319 (N_27319,N_26829,N_26803);
nand U27320 (N_27320,N_26808,N_26521);
or U27321 (N_27321,N_26819,N_26924);
and U27322 (N_27322,N_26540,N_26838);
nand U27323 (N_27323,N_26596,N_26562);
nor U27324 (N_27324,N_26651,N_26897);
and U27325 (N_27325,N_26855,N_26892);
xnor U27326 (N_27326,N_26978,N_26735);
xnor U27327 (N_27327,N_26996,N_26709);
or U27328 (N_27328,N_26855,N_26885);
or U27329 (N_27329,N_26505,N_26511);
and U27330 (N_27330,N_26578,N_26707);
or U27331 (N_27331,N_26780,N_26617);
nor U27332 (N_27332,N_26866,N_26963);
nand U27333 (N_27333,N_26939,N_26675);
and U27334 (N_27334,N_26743,N_26969);
or U27335 (N_27335,N_26684,N_26861);
xor U27336 (N_27336,N_26812,N_26614);
nand U27337 (N_27337,N_26901,N_26841);
nand U27338 (N_27338,N_26517,N_26605);
nor U27339 (N_27339,N_26991,N_26960);
xnor U27340 (N_27340,N_26521,N_26730);
nand U27341 (N_27341,N_26846,N_26607);
or U27342 (N_27342,N_26555,N_26801);
or U27343 (N_27343,N_26596,N_26890);
xor U27344 (N_27344,N_26599,N_26872);
and U27345 (N_27345,N_26784,N_26591);
and U27346 (N_27346,N_26685,N_26853);
and U27347 (N_27347,N_26722,N_26790);
or U27348 (N_27348,N_26706,N_26914);
nor U27349 (N_27349,N_26796,N_26631);
nor U27350 (N_27350,N_26595,N_26646);
xor U27351 (N_27351,N_26690,N_26831);
and U27352 (N_27352,N_26833,N_26531);
nand U27353 (N_27353,N_26861,N_26931);
or U27354 (N_27354,N_26518,N_26850);
nor U27355 (N_27355,N_26798,N_26521);
or U27356 (N_27356,N_26986,N_26549);
nand U27357 (N_27357,N_26906,N_26803);
nand U27358 (N_27358,N_26545,N_26916);
and U27359 (N_27359,N_26782,N_26757);
or U27360 (N_27360,N_26955,N_26844);
xnor U27361 (N_27361,N_26674,N_26809);
or U27362 (N_27362,N_26656,N_26737);
or U27363 (N_27363,N_26932,N_26991);
or U27364 (N_27364,N_26981,N_26638);
xnor U27365 (N_27365,N_26701,N_26861);
xor U27366 (N_27366,N_26919,N_26821);
nand U27367 (N_27367,N_26937,N_26922);
xor U27368 (N_27368,N_26689,N_26714);
nor U27369 (N_27369,N_26889,N_26531);
or U27370 (N_27370,N_26977,N_26882);
or U27371 (N_27371,N_26900,N_26611);
or U27372 (N_27372,N_26870,N_26762);
xor U27373 (N_27373,N_26712,N_26785);
or U27374 (N_27374,N_26586,N_26603);
xnor U27375 (N_27375,N_26531,N_26939);
xnor U27376 (N_27376,N_26703,N_26812);
nand U27377 (N_27377,N_26773,N_26823);
nor U27378 (N_27378,N_26951,N_26760);
nand U27379 (N_27379,N_26845,N_26923);
and U27380 (N_27380,N_26683,N_26937);
nand U27381 (N_27381,N_26881,N_26962);
xnor U27382 (N_27382,N_26799,N_26747);
xnor U27383 (N_27383,N_26857,N_26572);
nand U27384 (N_27384,N_26769,N_26736);
xor U27385 (N_27385,N_26595,N_26713);
or U27386 (N_27386,N_26853,N_26755);
and U27387 (N_27387,N_26596,N_26642);
nor U27388 (N_27388,N_26565,N_26503);
nor U27389 (N_27389,N_26645,N_26660);
nor U27390 (N_27390,N_26733,N_26691);
and U27391 (N_27391,N_26653,N_26694);
nor U27392 (N_27392,N_26861,N_26699);
nor U27393 (N_27393,N_26879,N_26796);
nand U27394 (N_27394,N_26563,N_26663);
nand U27395 (N_27395,N_26820,N_26683);
nor U27396 (N_27396,N_26735,N_26659);
and U27397 (N_27397,N_26987,N_26505);
xor U27398 (N_27398,N_26904,N_26968);
or U27399 (N_27399,N_26745,N_26834);
nor U27400 (N_27400,N_26669,N_26750);
xnor U27401 (N_27401,N_26800,N_26663);
or U27402 (N_27402,N_26715,N_26771);
or U27403 (N_27403,N_26628,N_26684);
and U27404 (N_27404,N_26893,N_26612);
and U27405 (N_27405,N_26854,N_26598);
or U27406 (N_27406,N_26837,N_26961);
or U27407 (N_27407,N_26743,N_26551);
and U27408 (N_27408,N_26732,N_26758);
nand U27409 (N_27409,N_26874,N_26666);
nand U27410 (N_27410,N_26864,N_26920);
and U27411 (N_27411,N_26618,N_26899);
and U27412 (N_27412,N_26639,N_26840);
and U27413 (N_27413,N_26569,N_26730);
nand U27414 (N_27414,N_26691,N_26842);
xor U27415 (N_27415,N_26596,N_26830);
nor U27416 (N_27416,N_26604,N_26724);
nand U27417 (N_27417,N_26753,N_26786);
and U27418 (N_27418,N_26976,N_26777);
nor U27419 (N_27419,N_26921,N_26549);
nor U27420 (N_27420,N_26571,N_26712);
nor U27421 (N_27421,N_26716,N_26761);
nand U27422 (N_27422,N_26911,N_26744);
xor U27423 (N_27423,N_26625,N_26634);
xnor U27424 (N_27424,N_26620,N_26889);
nand U27425 (N_27425,N_26987,N_26659);
nand U27426 (N_27426,N_26874,N_26846);
nand U27427 (N_27427,N_26702,N_26883);
or U27428 (N_27428,N_26826,N_26666);
and U27429 (N_27429,N_26810,N_26561);
nand U27430 (N_27430,N_26985,N_26826);
and U27431 (N_27431,N_26733,N_26578);
and U27432 (N_27432,N_26647,N_26526);
and U27433 (N_27433,N_26952,N_26866);
nand U27434 (N_27434,N_26912,N_26899);
nor U27435 (N_27435,N_26775,N_26665);
nand U27436 (N_27436,N_26743,N_26621);
xnor U27437 (N_27437,N_26683,N_26901);
or U27438 (N_27438,N_26623,N_26612);
nand U27439 (N_27439,N_26954,N_26943);
nand U27440 (N_27440,N_26982,N_26905);
nor U27441 (N_27441,N_26721,N_26996);
and U27442 (N_27442,N_26829,N_26701);
nand U27443 (N_27443,N_26987,N_26955);
nor U27444 (N_27444,N_26562,N_26743);
or U27445 (N_27445,N_26740,N_26932);
nand U27446 (N_27446,N_26654,N_26773);
or U27447 (N_27447,N_26597,N_26601);
and U27448 (N_27448,N_26975,N_26927);
nand U27449 (N_27449,N_26910,N_26902);
xor U27450 (N_27450,N_26940,N_26960);
xnor U27451 (N_27451,N_26609,N_26773);
or U27452 (N_27452,N_26606,N_26828);
and U27453 (N_27453,N_26902,N_26908);
xor U27454 (N_27454,N_26756,N_26572);
and U27455 (N_27455,N_26912,N_26625);
and U27456 (N_27456,N_26777,N_26695);
nand U27457 (N_27457,N_26819,N_26675);
nor U27458 (N_27458,N_26842,N_26509);
or U27459 (N_27459,N_26716,N_26755);
nor U27460 (N_27460,N_26656,N_26888);
or U27461 (N_27461,N_26694,N_26952);
nor U27462 (N_27462,N_26912,N_26839);
nand U27463 (N_27463,N_26583,N_26741);
nand U27464 (N_27464,N_26748,N_26811);
and U27465 (N_27465,N_26874,N_26517);
nand U27466 (N_27466,N_26826,N_26742);
xnor U27467 (N_27467,N_26558,N_26997);
or U27468 (N_27468,N_26560,N_26620);
xor U27469 (N_27469,N_26801,N_26639);
and U27470 (N_27470,N_26924,N_26614);
and U27471 (N_27471,N_26517,N_26659);
xnor U27472 (N_27472,N_26951,N_26706);
and U27473 (N_27473,N_26952,N_26772);
xnor U27474 (N_27474,N_26736,N_26646);
nor U27475 (N_27475,N_26813,N_26953);
nand U27476 (N_27476,N_26655,N_26657);
nand U27477 (N_27477,N_26747,N_26772);
xor U27478 (N_27478,N_26683,N_26529);
xnor U27479 (N_27479,N_26738,N_26955);
xnor U27480 (N_27480,N_26857,N_26613);
or U27481 (N_27481,N_26801,N_26802);
nand U27482 (N_27482,N_26615,N_26940);
nand U27483 (N_27483,N_26607,N_26932);
or U27484 (N_27484,N_26920,N_26852);
nand U27485 (N_27485,N_26981,N_26685);
xnor U27486 (N_27486,N_26795,N_26714);
or U27487 (N_27487,N_26661,N_26921);
or U27488 (N_27488,N_26763,N_26598);
or U27489 (N_27489,N_26965,N_26709);
or U27490 (N_27490,N_26984,N_26631);
xor U27491 (N_27491,N_26518,N_26858);
xnor U27492 (N_27492,N_26714,N_26692);
or U27493 (N_27493,N_26605,N_26950);
nor U27494 (N_27494,N_26501,N_26969);
nand U27495 (N_27495,N_26612,N_26843);
nand U27496 (N_27496,N_26814,N_26719);
and U27497 (N_27497,N_26564,N_26501);
xor U27498 (N_27498,N_26905,N_26855);
nor U27499 (N_27499,N_26665,N_26661);
nand U27500 (N_27500,N_27382,N_27011);
xnor U27501 (N_27501,N_27368,N_27328);
nand U27502 (N_27502,N_27111,N_27360);
nand U27503 (N_27503,N_27491,N_27374);
xor U27504 (N_27504,N_27054,N_27377);
xor U27505 (N_27505,N_27334,N_27286);
xnor U27506 (N_27506,N_27469,N_27242);
and U27507 (N_27507,N_27065,N_27346);
xor U27508 (N_27508,N_27265,N_27117);
and U27509 (N_27509,N_27338,N_27320);
nor U27510 (N_27510,N_27272,N_27262);
nor U27511 (N_27511,N_27051,N_27135);
or U27512 (N_27512,N_27427,N_27247);
and U27513 (N_27513,N_27191,N_27058);
nor U27514 (N_27514,N_27288,N_27433);
nor U27515 (N_27515,N_27268,N_27486);
and U27516 (N_27516,N_27497,N_27040);
nor U27517 (N_27517,N_27012,N_27182);
or U27518 (N_27518,N_27141,N_27251);
nor U27519 (N_27519,N_27132,N_27110);
or U27520 (N_27520,N_27294,N_27077);
nand U27521 (N_27521,N_27425,N_27416);
and U27522 (N_27522,N_27487,N_27366);
and U27523 (N_27523,N_27059,N_27315);
and U27524 (N_27524,N_27094,N_27130);
nand U27525 (N_27525,N_27003,N_27035);
nand U27526 (N_27526,N_27140,N_27047);
nor U27527 (N_27527,N_27475,N_27006);
or U27528 (N_27528,N_27109,N_27206);
xor U27529 (N_27529,N_27498,N_27235);
nor U27530 (N_27530,N_27436,N_27052);
or U27531 (N_27531,N_27091,N_27169);
and U27532 (N_27532,N_27093,N_27402);
and U27533 (N_27533,N_27451,N_27125);
nor U27534 (N_27534,N_27038,N_27420);
and U27535 (N_27535,N_27490,N_27144);
nor U27536 (N_27536,N_27361,N_27337);
nor U27537 (N_27537,N_27120,N_27378);
nand U27538 (N_27538,N_27319,N_27055);
or U27539 (N_27539,N_27018,N_27325);
and U27540 (N_27540,N_27285,N_27134);
nand U27541 (N_27541,N_27356,N_27151);
and U27542 (N_27542,N_27423,N_27230);
or U27543 (N_27543,N_27303,N_27183);
or U27544 (N_27544,N_27260,N_27193);
xnor U27545 (N_27545,N_27195,N_27063);
and U27546 (N_27546,N_27188,N_27042);
or U27547 (N_27547,N_27309,N_27215);
nor U27548 (N_27548,N_27343,N_27062);
xor U27549 (N_27549,N_27074,N_27253);
nor U27550 (N_27550,N_27176,N_27269);
xnor U27551 (N_27551,N_27305,N_27161);
or U27552 (N_27552,N_27331,N_27186);
or U27553 (N_27553,N_27118,N_27192);
nand U27554 (N_27554,N_27019,N_27148);
nor U27555 (N_27555,N_27421,N_27385);
and U27556 (N_27556,N_27217,N_27221);
and U27557 (N_27557,N_27129,N_27409);
and U27558 (N_27558,N_27267,N_27258);
or U27559 (N_27559,N_27293,N_27126);
xnor U27560 (N_27560,N_27399,N_27101);
xor U27561 (N_27561,N_27102,N_27085);
and U27562 (N_27562,N_27311,N_27313);
or U27563 (N_27563,N_27204,N_27446);
and U27564 (N_27564,N_27170,N_27185);
nand U27565 (N_27565,N_27310,N_27297);
nor U27566 (N_27566,N_27166,N_27457);
nand U27567 (N_27567,N_27428,N_27456);
xor U27568 (N_27568,N_27381,N_27424);
and U27569 (N_27569,N_27154,N_27034);
or U27570 (N_27570,N_27033,N_27452);
xor U27571 (N_27571,N_27316,N_27061);
and U27572 (N_27572,N_27112,N_27292);
and U27573 (N_27573,N_27239,N_27139);
nand U27574 (N_27574,N_27228,N_27043);
xor U27575 (N_27575,N_27367,N_27454);
xnor U27576 (N_27576,N_27435,N_27296);
xor U27577 (N_27577,N_27150,N_27280);
nor U27578 (N_27578,N_27004,N_27276);
nor U27579 (N_27579,N_27460,N_27392);
nor U27580 (N_27580,N_27159,N_27282);
nand U27581 (N_27581,N_27224,N_27256);
and U27582 (N_27582,N_27008,N_27037);
or U27583 (N_27583,N_27429,N_27283);
and U27584 (N_27584,N_27225,N_27445);
nand U27585 (N_27585,N_27016,N_27149);
or U27586 (N_27586,N_27273,N_27359);
xnor U27587 (N_27587,N_27244,N_27173);
nor U27588 (N_27588,N_27390,N_27133);
and U27589 (N_27589,N_27413,N_27370);
and U27590 (N_27590,N_27398,N_27455);
xnor U27591 (N_27591,N_27027,N_27279);
or U27592 (N_27592,N_27180,N_27086);
nor U27593 (N_27593,N_27495,N_27029);
nor U27594 (N_27594,N_27187,N_27128);
or U27595 (N_27595,N_27291,N_27137);
nand U27596 (N_27596,N_27259,N_27394);
and U27597 (N_27597,N_27252,N_27344);
nor U27598 (N_27598,N_27300,N_27417);
nor U27599 (N_27599,N_27348,N_27005);
nand U27600 (N_27600,N_27321,N_27278);
xnor U27601 (N_27601,N_27347,N_27009);
nand U27602 (N_27602,N_27241,N_27067);
and U27603 (N_27603,N_27340,N_27422);
and U27604 (N_27604,N_27226,N_27389);
xnor U27605 (N_27605,N_27301,N_27463);
xor U27606 (N_27606,N_27156,N_27468);
nor U27607 (N_27607,N_27318,N_27127);
nor U27608 (N_27608,N_27393,N_27122);
and U27609 (N_27609,N_27198,N_27240);
nor U27610 (N_27610,N_27254,N_27071);
nand U27611 (N_27611,N_27165,N_27082);
or U27612 (N_27612,N_27326,N_27358);
nand U27613 (N_27613,N_27053,N_27200);
or U27614 (N_27614,N_27017,N_27023);
nand U27615 (N_27615,N_27025,N_27243);
or U27616 (N_27616,N_27474,N_27201);
nand U27617 (N_27617,N_27068,N_27146);
and U27618 (N_27618,N_27371,N_27069);
and U27619 (N_27619,N_27307,N_27073);
and U27620 (N_27620,N_27190,N_27332);
or U27621 (N_27621,N_27284,N_27163);
and U27622 (N_27622,N_27057,N_27412);
nor U27623 (N_27623,N_27369,N_27222);
xnor U27624 (N_27624,N_27229,N_27046);
nand U27625 (N_27625,N_27196,N_27345);
nand U27626 (N_27626,N_27401,N_27335);
nand U27627 (N_27627,N_27103,N_27066);
and U27628 (N_27628,N_27461,N_27096);
and U27629 (N_27629,N_27442,N_27080);
xnor U27630 (N_27630,N_27208,N_27314);
or U27631 (N_27631,N_27266,N_27197);
nor U27632 (N_27632,N_27174,N_27261);
nand U27633 (N_27633,N_27375,N_27383);
xnor U27634 (N_27634,N_27362,N_27105);
and U27635 (N_27635,N_27030,N_27339);
nand U27636 (N_27636,N_27324,N_27031);
nand U27637 (N_27637,N_27396,N_27124);
or U27638 (N_27638,N_27289,N_27171);
xor U27639 (N_27639,N_27471,N_27199);
and U27640 (N_27640,N_27142,N_27090);
nor U27641 (N_27641,N_27323,N_27353);
nand U27642 (N_27642,N_27079,N_27364);
or U27643 (N_27643,N_27218,N_27431);
and U27644 (N_27644,N_27352,N_27365);
nand U27645 (N_27645,N_27322,N_27021);
nor U27646 (N_27646,N_27441,N_27257);
or U27647 (N_27647,N_27041,N_27231);
and U27648 (N_27648,N_27084,N_27060);
or U27649 (N_27649,N_27363,N_27449);
nand U27650 (N_27650,N_27184,N_27189);
xor U27651 (N_27651,N_27216,N_27249);
or U27652 (N_27652,N_27181,N_27440);
or U27653 (N_27653,N_27404,N_27317);
or U27654 (N_27654,N_27237,N_27472);
nor U27655 (N_27655,N_27175,N_27210);
xnor U27656 (N_27656,N_27083,N_27312);
and U27657 (N_27657,N_27426,N_27414);
xor U27658 (N_27658,N_27407,N_27081);
nor U27659 (N_27659,N_27354,N_27290);
xnor U27660 (N_27660,N_27341,N_27333);
or U27661 (N_27661,N_27443,N_27476);
and U27662 (N_27662,N_27271,N_27114);
nor U27663 (N_27663,N_27419,N_27095);
or U27664 (N_27664,N_27403,N_27075);
or U27665 (N_27665,N_27167,N_27306);
nor U27666 (N_27666,N_27482,N_27357);
xor U27667 (N_27667,N_27119,N_27088);
xor U27668 (N_27668,N_27207,N_27178);
nor U27669 (N_27669,N_27478,N_27388);
xor U27670 (N_27670,N_27108,N_27342);
or U27671 (N_27671,N_27349,N_27479);
or U27672 (N_27672,N_27145,N_27212);
nand U27673 (N_27673,N_27430,N_27202);
xor U27674 (N_27674,N_27131,N_27097);
nand U27675 (N_27675,N_27026,N_27405);
nor U27676 (N_27676,N_27287,N_27466);
xnor U27677 (N_27677,N_27400,N_27032);
or U27678 (N_27678,N_27411,N_27219);
nand U27679 (N_27679,N_27483,N_27010);
nand U27680 (N_27680,N_27234,N_27379);
and U27681 (N_27681,N_27233,N_27014);
or U27682 (N_27682,N_27078,N_27000);
nand U27683 (N_27683,N_27263,N_27158);
and U27684 (N_27684,N_27499,N_27387);
nor U27685 (N_27685,N_27488,N_27064);
and U27686 (N_27686,N_27213,N_27056);
nand U27687 (N_27687,N_27232,N_27121);
nand U27688 (N_27688,N_27104,N_27329);
nor U27689 (N_27689,N_27152,N_27236);
xor U27690 (N_27690,N_27432,N_27299);
and U27691 (N_27691,N_27327,N_27238);
xnor U27692 (N_27692,N_27157,N_27462);
nand U27693 (N_27693,N_27408,N_27113);
and U27694 (N_27694,N_27143,N_27098);
nand U27695 (N_27695,N_27194,N_27415);
xnor U27696 (N_27696,N_27087,N_27048);
xnor U27697 (N_27697,N_27485,N_27281);
nor U27698 (N_27698,N_27264,N_27489);
nand U27699 (N_27699,N_27172,N_27211);
nor U27700 (N_27700,N_27391,N_27050);
nand U27701 (N_27701,N_27450,N_27464);
nor U27702 (N_27702,N_27410,N_27336);
xnor U27703 (N_27703,N_27028,N_27024);
nand U27704 (N_27704,N_27484,N_27355);
or U27705 (N_27705,N_27439,N_27274);
or U27706 (N_27706,N_27155,N_27162);
xor U27707 (N_27707,N_27448,N_27123);
xnor U27708 (N_27708,N_27397,N_27275);
nor U27709 (N_27709,N_27384,N_27138);
or U27710 (N_27710,N_27480,N_27380);
or U27711 (N_27711,N_27160,N_27115);
nand U27712 (N_27712,N_27007,N_27295);
nor U27713 (N_27713,N_27100,N_27467);
nand U27714 (N_27714,N_27330,N_27036);
nand U27715 (N_27715,N_27001,N_27020);
nor U27716 (N_27716,N_27248,N_27089);
nor U27717 (N_27717,N_27227,N_27153);
or U27718 (N_27718,N_27406,N_27044);
xor U27719 (N_27719,N_27434,N_27350);
and U27720 (N_27720,N_27473,N_27458);
or U27721 (N_27721,N_27106,N_27039);
xor U27722 (N_27722,N_27372,N_27465);
nor U27723 (N_27723,N_27255,N_27304);
nand U27724 (N_27724,N_27099,N_27013);
and U27725 (N_27725,N_27002,N_27444);
nand U27726 (N_27726,N_27092,N_27214);
and U27727 (N_27727,N_27220,N_27493);
nor U27728 (N_27728,N_27246,N_27250);
nand U27729 (N_27729,N_27076,N_27308);
or U27730 (N_27730,N_27245,N_27437);
or U27731 (N_27731,N_27179,N_27072);
or U27732 (N_27732,N_27136,N_27386);
xnor U27733 (N_27733,N_27070,N_27022);
nor U27734 (N_27734,N_27107,N_27209);
and U27735 (N_27735,N_27438,N_27277);
or U27736 (N_27736,N_27177,N_27418);
or U27737 (N_27737,N_27168,N_27302);
or U27738 (N_27738,N_27223,N_27015);
nand U27739 (N_27739,N_27270,N_27494);
nand U27740 (N_27740,N_27470,N_27395);
and U27741 (N_27741,N_27351,N_27049);
xor U27742 (N_27742,N_27203,N_27481);
and U27743 (N_27743,N_27147,N_27298);
and U27744 (N_27744,N_27459,N_27373);
and U27745 (N_27745,N_27453,N_27447);
and U27746 (N_27746,N_27116,N_27477);
and U27747 (N_27747,N_27496,N_27164);
nand U27748 (N_27748,N_27045,N_27376);
nor U27749 (N_27749,N_27205,N_27492);
nor U27750 (N_27750,N_27186,N_27352);
and U27751 (N_27751,N_27145,N_27207);
and U27752 (N_27752,N_27214,N_27037);
or U27753 (N_27753,N_27006,N_27061);
nand U27754 (N_27754,N_27330,N_27103);
or U27755 (N_27755,N_27424,N_27251);
xor U27756 (N_27756,N_27333,N_27198);
or U27757 (N_27757,N_27413,N_27331);
or U27758 (N_27758,N_27166,N_27168);
nand U27759 (N_27759,N_27152,N_27001);
xor U27760 (N_27760,N_27405,N_27262);
xor U27761 (N_27761,N_27072,N_27042);
nand U27762 (N_27762,N_27335,N_27454);
nor U27763 (N_27763,N_27468,N_27037);
or U27764 (N_27764,N_27088,N_27046);
or U27765 (N_27765,N_27313,N_27376);
and U27766 (N_27766,N_27392,N_27479);
or U27767 (N_27767,N_27277,N_27358);
and U27768 (N_27768,N_27442,N_27282);
nor U27769 (N_27769,N_27051,N_27130);
xnor U27770 (N_27770,N_27262,N_27080);
nor U27771 (N_27771,N_27227,N_27076);
and U27772 (N_27772,N_27172,N_27368);
and U27773 (N_27773,N_27140,N_27432);
xnor U27774 (N_27774,N_27409,N_27232);
xnor U27775 (N_27775,N_27012,N_27202);
nor U27776 (N_27776,N_27036,N_27233);
xor U27777 (N_27777,N_27261,N_27316);
xnor U27778 (N_27778,N_27281,N_27092);
or U27779 (N_27779,N_27477,N_27311);
and U27780 (N_27780,N_27108,N_27456);
nor U27781 (N_27781,N_27333,N_27063);
xor U27782 (N_27782,N_27046,N_27441);
xnor U27783 (N_27783,N_27473,N_27322);
xor U27784 (N_27784,N_27360,N_27029);
nand U27785 (N_27785,N_27394,N_27182);
xnor U27786 (N_27786,N_27480,N_27175);
nand U27787 (N_27787,N_27242,N_27292);
nor U27788 (N_27788,N_27045,N_27001);
or U27789 (N_27789,N_27443,N_27195);
xnor U27790 (N_27790,N_27104,N_27406);
nand U27791 (N_27791,N_27123,N_27217);
nor U27792 (N_27792,N_27281,N_27066);
and U27793 (N_27793,N_27392,N_27349);
and U27794 (N_27794,N_27355,N_27174);
nand U27795 (N_27795,N_27030,N_27078);
or U27796 (N_27796,N_27433,N_27182);
and U27797 (N_27797,N_27229,N_27422);
nand U27798 (N_27798,N_27472,N_27151);
or U27799 (N_27799,N_27480,N_27424);
nand U27800 (N_27800,N_27402,N_27465);
xor U27801 (N_27801,N_27017,N_27270);
nand U27802 (N_27802,N_27468,N_27191);
nand U27803 (N_27803,N_27026,N_27453);
and U27804 (N_27804,N_27096,N_27201);
xnor U27805 (N_27805,N_27400,N_27172);
or U27806 (N_27806,N_27166,N_27381);
nand U27807 (N_27807,N_27344,N_27496);
xor U27808 (N_27808,N_27423,N_27357);
or U27809 (N_27809,N_27132,N_27498);
and U27810 (N_27810,N_27499,N_27157);
nor U27811 (N_27811,N_27251,N_27202);
nand U27812 (N_27812,N_27489,N_27105);
nor U27813 (N_27813,N_27027,N_27249);
or U27814 (N_27814,N_27476,N_27172);
and U27815 (N_27815,N_27388,N_27046);
nand U27816 (N_27816,N_27038,N_27395);
or U27817 (N_27817,N_27359,N_27027);
or U27818 (N_27818,N_27084,N_27100);
and U27819 (N_27819,N_27149,N_27105);
or U27820 (N_27820,N_27460,N_27053);
and U27821 (N_27821,N_27446,N_27054);
or U27822 (N_27822,N_27333,N_27220);
and U27823 (N_27823,N_27028,N_27123);
or U27824 (N_27824,N_27053,N_27159);
nor U27825 (N_27825,N_27293,N_27170);
nand U27826 (N_27826,N_27434,N_27156);
nand U27827 (N_27827,N_27156,N_27028);
nor U27828 (N_27828,N_27493,N_27494);
nor U27829 (N_27829,N_27381,N_27476);
nand U27830 (N_27830,N_27179,N_27446);
nand U27831 (N_27831,N_27447,N_27307);
or U27832 (N_27832,N_27110,N_27489);
or U27833 (N_27833,N_27052,N_27207);
and U27834 (N_27834,N_27088,N_27332);
nand U27835 (N_27835,N_27475,N_27312);
xnor U27836 (N_27836,N_27494,N_27139);
and U27837 (N_27837,N_27437,N_27417);
nand U27838 (N_27838,N_27248,N_27075);
nand U27839 (N_27839,N_27234,N_27097);
or U27840 (N_27840,N_27004,N_27123);
nand U27841 (N_27841,N_27145,N_27425);
or U27842 (N_27842,N_27186,N_27433);
nand U27843 (N_27843,N_27152,N_27184);
nand U27844 (N_27844,N_27363,N_27481);
nor U27845 (N_27845,N_27008,N_27166);
nand U27846 (N_27846,N_27282,N_27141);
nor U27847 (N_27847,N_27301,N_27167);
and U27848 (N_27848,N_27371,N_27286);
xor U27849 (N_27849,N_27080,N_27276);
nor U27850 (N_27850,N_27310,N_27183);
xor U27851 (N_27851,N_27430,N_27184);
and U27852 (N_27852,N_27158,N_27017);
xor U27853 (N_27853,N_27189,N_27129);
xor U27854 (N_27854,N_27110,N_27441);
and U27855 (N_27855,N_27021,N_27163);
nor U27856 (N_27856,N_27363,N_27273);
xnor U27857 (N_27857,N_27085,N_27333);
nand U27858 (N_27858,N_27288,N_27242);
nor U27859 (N_27859,N_27275,N_27112);
nor U27860 (N_27860,N_27084,N_27043);
nor U27861 (N_27861,N_27016,N_27046);
and U27862 (N_27862,N_27269,N_27246);
nand U27863 (N_27863,N_27193,N_27288);
xnor U27864 (N_27864,N_27334,N_27371);
or U27865 (N_27865,N_27210,N_27250);
and U27866 (N_27866,N_27009,N_27173);
and U27867 (N_27867,N_27322,N_27062);
nand U27868 (N_27868,N_27293,N_27295);
and U27869 (N_27869,N_27175,N_27453);
or U27870 (N_27870,N_27036,N_27039);
and U27871 (N_27871,N_27173,N_27405);
or U27872 (N_27872,N_27157,N_27098);
nor U27873 (N_27873,N_27157,N_27432);
nor U27874 (N_27874,N_27245,N_27344);
or U27875 (N_27875,N_27029,N_27178);
or U27876 (N_27876,N_27317,N_27174);
xor U27877 (N_27877,N_27461,N_27305);
xor U27878 (N_27878,N_27327,N_27381);
and U27879 (N_27879,N_27402,N_27429);
nand U27880 (N_27880,N_27151,N_27110);
xnor U27881 (N_27881,N_27154,N_27038);
nor U27882 (N_27882,N_27450,N_27442);
nor U27883 (N_27883,N_27005,N_27421);
nand U27884 (N_27884,N_27433,N_27205);
xnor U27885 (N_27885,N_27312,N_27026);
or U27886 (N_27886,N_27400,N_27134);
xnor U27887 (N_27887,N_27385,N_27418);
and U27888 (N_27888,N_27032,N_27135);
nor U27889 (N_27889,N_27066,N_27387);
and U27890 (N_27890,N_27221,N_27218);
or U27891 (N_27891,N_27433,N_27467);
nor U27892 (N_27892,N_27399,N_27428);
nand U27893 (N_27893,N_27470,N_27027);
or U27894 (N_27894,N_27137,N_27133);
nand U27895 (N_27895,N_27360,N_27231);
nor U27896 (N_27896,N_27124,N_27386);
and U27897 (N_27897,N_27184,N_27123);
nor U27898 (N_27898,N_27116,N_27226);
or U27899 (N_27899,N_27059,N_27378);
nand U27900 (N_27900,N_27076,N_27005);
or U27901 (N_27901,N_27217,N_27102);
or U27902 (N_27902,N_27157,N_27421);
nor U27903 (N_27903,N_27325,N_27112);
xnor U27904 (N_27904,N_27108,N_27000);
or U27905 (N_27905,N_27463,N_27012);
nor U27906 (N_27906,N_27038,N_27442);
or U27907 (N_27907,N_27387,N_27095);
and U27908 (N_27908,N_27333,N_27203);
or U27909 (N_27909,N_27260,N_27186);
or U27910 (N_27910,N_27075,N_27301);
or U27911 (N_27911,N_27270,N_27020);
and U27912 (N_27912,N_27478,N_27274);
or U27913 (N_27913,N_27274,N_27315);
nand U27914 (N_27914,N_27128,N_27169);
or U27915 (N_27915,N_27012,N_27153);
xnor U27916 (N_27916,N_27124,N_27428);
or U27917 (N_27917,N_27055,N_27068);
or U27918 (N_27918,N_27431,N_27329);
xnor U27919 (N_27919,N_27393,N_27044);
and U27920 (N_27920,N_27480,N_27061);
or U27921 (N_27921,N_27060,N_27370);
or U27922 (N_27922,N_27200,N_27401);
nand U27923 (N_27923,N_27285,N_27313);
nand U27924 (N_27924,N_27377,N_27325);
xor U27925 (N_27925,N_27487,N_27243);
nor U27926 (N_27926,N_27425,N_27275);
and U27927 (N_27927,N_27294,N_27307);
xor U27928 (N_27928,N_27250,N_27364);
xnor U27929 (N_27929,N_27067,N_27007);
or U27930 (N_27930,N_27320,N_27457);
xnor U27931 (N_27931,N_27226,N_27424);
or U27932 (N_27932,N_27340,N_27196);
nor U27933 (N_27933,N_27430,N_27152);
nand U27934 (N_27934,N_27229,N_27261);
and U27935 (N_27935,N_27062,N_27391);
or U27936 (N_27936,N_27231,N_27222);
nand U27937 (N_27937,N_27153,N_27302);
nor U27938 (N_27938,N_27340,N_27090);
xnor U27939 (N_27939,N_27193,N_27026);
nor U27940 (N_27940,N_27009,N_27239);
xor U27941 (N_27941,N_27385,N_27067);
nand U27942 (N_27942,N_27425,N_27189);
nor U27943 (N_27943,N_27084,N_27452);
xor U27944 (N_27944,N_27116,N_27054);
nor U27945 (N_27945,N_27494,N_27252);
xor U27946 (N_27946,N_27266,N_27193);
or U27947 (N_27947,N_27062,N_27183);
or U27948 (N_27948,N_27134,N_27327);
xnor U27949 (N_27949,N_27373,N_27236);
xor U27950 (N_27950,N_27058,N_27451);
nand U27951 (N_27951,N_27028,N_27247);
and U27952 (N_27952,N_27250,N_27451);
nor U27953 (N_27953,N_27035,N_27141);
nand U27954 (N_27954,N_27344,N_27482);
xor U27955 (N_27955,N_27211,N_27338);
xnor U27956 (N_27956,N_27105,N_27183);
nand U27957 (N_27957,N_27203,N_27383);
nand U27958 (N_27958,N_27320,N_27478);
and U27959 (N_27959,N_27174,N_27246);
nand U27960 (N_27960,N_27060,N_27489);
nand U27961 (N_27961,N_27168,N_27358);
and U27962 (N_27962,N_27187,N_27426);
nor U27963 (N_27963,N_27036,N_27306);
nor U27964 (N_27964,N_27283,N_27167);
xnor U27965 (N_27965,N_27475,N_27216);
nand U27966 (N_27966,N_27255,N_27368);
xor U27967 (N_27967,N_27257,N_27416);
xor U27968 (N_27968,N_27331,N_27165);
or U27969 (N_27969,N_27177,N_27176);
nor U27970 (N_27970,N_27469,N_27048);
or U27971 (N_27971,N_27152,N_27371);
or U27972 (N_27972,N_27087,N_27107);
or U27973 (N_27973,N_27191,N_27156);
and U27974 (N_27974,N_27494,N_27019);
xnor U27975 (N_27975,N_27234,N_27290);
and U27976 (N_27976,N_27064,N_27435);
or U27977 (N_27977,N_27004,N_27381);
or U27978 (N_27978,N_27492,N_27152);
nor U27979 (N_27979,N_27115,N_27293);
and U27980 (N_27980,N_27439,N_27038);
xnor U27981 (N_27981,N_27366,N_27355);
nand U27982 (N_27982,N_27058,N_27089);
xnor U27983 (N_27983,N_27028,N_27175);
nor U27984 (N_27984,N_27375,N_27313);
nand U27985 (N_27985,N_27423,N_27488);
and U27986 (N_27986,N_27480,N_27497);
nor U27987 (N_27987,N_27496,N_27343);
or U27988 (N_27988,N_27131,N_27243);
or U27989 (N_27989,N_27264,N_27150);
nand U27990 (N_27990,N_27416,N_27333);
nor U27991 (N_27991,N_27033,N_27095);
nor U27992 (N_27992,N_27051,N_27347);
or U27993 (N_27993,N_27328,N_27225);
or U27994 (N_27994,N_27166,N_27296);
nor U27995 (N_27995,N_27166,N_27171);
or U27996 (N_27996,N_27389,N_27180);
nand U27997 (N_27997,N_27391,N_27448);
nor U27998 (N_27998,N_27098,N_27284);
nor U27999 (N_27999,N_27355,N_27203);
and U28000 (N_28000,N_27851,N_27584);
nor U28001 (N_28001,N_27788,N_27801);
nor U28002 (N_28002,N_27704,N_27543);
xnor U28003 (N_28003,N_27809,N_27917);
nand U28004 (N_28004,N_27511,N_27746);
and U28005 (N_28005,N_27762,N_27818);
nand U28006 (N_28006,N_27982,N_27840);
or U28007 (N_28007,N_27806,N_27789);
xnor U28008 (N_28008,N_27872,N_27923);
or U28009 (N_28009,N_27862,N_27524);
nor U28010 (N_28010,N_27767,N_27539);
xnor U28011 (N_28011,N_27516,N_27696);
nand U28012 (N_28012,N_27864,N_27514);
nor U28013 (N_28013,N_27920,N_27608);
nand U28014 (N_28014,N_27780,N_27568);
nand U28015 (N_28015,N_27937,N_27705);
nor U28016 (N_28016,N_27783,N_27531);
nor U28017 (N_28017,N_27737,N_27817);
nand U28018 (N_28018,N_27689,N_27976);
xor U28019 (N_28019,N_27763,N_27580);
or U28020 (N_28020,N_27638,N_27834);
nor U28021 (N_28021,N_27880,N_27756);
nand U28022 (N_28022,N_27552,N_27882);
and U28023 (N_28023,N_27983,N_27790);
and U28024 (N_28024,N_27869,N_27897);
and U28025 (N_28025,N_27969,N_27883);
or U28026 (N_28026,N_27861,N_27632);
xnor U28027 (N_28027,N_27706,N_27691);
and U28028 (N_28028,N_27835,N_27606);
xor U28029 (N_28029,N_27905,N_27595);
or U28030 (N_28030,N_27813,N_27570);
and U28031 (N_28031,N_27744,N_27957);
or U28032 (N_28032,N_27940,N_27826);
nor U28033 (N_28033,N_27959,N_27645);
xnor U28034 (N_28034,N_27932,N_27769);
xor U28035 (N_28035,N_27676,N_27623);
nor U28036 (N_28036,N_27874,N_27658);
or U28037 (N_28037,N_27863,N_27707);
and U28038 (N_28038,N_27942,N_27977);
nand U28039 (N_28039,N_27564,N_27906);
or U28040 (N_28040,N_27802,N_27992);
xnor U28041 (N_28041,N_27566,N_27655);
and U28042 (N_28042,N_27928,N_27505);
or U28043 (N_28043,N_27963,N_27934);
or U28044 (N_28044,N_27731,N_27815);
nor U28045 (N_28045,N_27948,N_27830);
nand U28046 (N_28046,N_27657,N_27824);
nor U28047 (N_28047,N_27919,N_27592);
nand U28048 (N_28048,N_27823,N_27804);
xnor U28049 (N_28049,N_27891,N_27654);
nand U28050 (N_28050,N_27641,N_27520);
and U28051 (N_28051,N_27816,N_27962);
and U28052 (N_28052,N_27659,N_27719);
xor U28053 (N_28053,N_27821,N_27873);
and U28054 (N_28054,N_27661,N_27598);
nand U28055 (N_28055,N_27681,N_27546);
or U28056 (N_28056,N_27986,N_27774);
and U28057 (N_28057,N_27832,N_27672);
nor U28058 (N_28058,N_27971,N_27582);
nor U28059 (N_28059,N_27683,N_27727);
xor U28060 (N_28060,N_27587,N_27601);
nand U28061 (N_28061,N_27793,N_27939);
nor U28062 (N_28062,N_27602,N_27833);
nand U28063 (N_28063,N_27604,N_27922);
and U28064 (N_28064,N_27911,N_27925);
or U28065 (N_28065,N_27717,N_27904);
or U28066 (N_28066,N_27618,N_27798);
and U28067 (N_28067,N_27627,N_27664);
and U28068 (N_28068,N_27579,N_27663);
nand U28069 (N_28069,N_27677,N_27775);
nor U28070 (N_28070,N_27799,N_27504);
nor U28071 (N_28071,N_27513,N_27611);
nand U28072 (N_28072,N_27693,N_27590);
xor U28073 (N_28073,N_27692,N_27567);
nand U28074 (N_28074,N_27770,N_27886);
nand U28075 (N_28075,N_27711,N_27892);
or U28076 (N_28076,N_27895,N_27558);
nand U28077 (N_28077,N_27837,N_27665);
xor U28078 (N_28078,N_27915,N_27577);
nand U28079 (N_28079,N_27966,N_27916);
and U28080 (N_28080,N_27822,N_27903);
nand U28081 (N_28081,N_27749,N_27617);
or U28082 (N_28082,N_27854,N_27831);
xnor U28083 (N_28083,N_27888,N_27860);
nor U28084 (N_28084,N_27684,N_27525);
and U28085 (N_28085,N_27984,N_27648);
xnor U28086 (N_28086,N_27954,N_27941);
or U28087 (N_28087,N_27550,N_27572);
nand U28088 (N_28088,N_27878,N_27967);
and U28089 (N_28089,N_27521,N_27970);
xnor U28090 (N_28090,N_27615,N_27896);
xor U28091 (N_28091,N_27929,N_27968);
and U28092 (N_28092,N_27686,N_27666);
nor U28093 (N_28093,N_27679,N_27800);
xor U28094 (N_28094,N_27597,N_27838);
nand U28095 (N_28095,N_27740,N_27865);
and U28096 (N_28096,N_27777,N_27752);
xnor U28097 (N_28097,N_27947,N_27633);
nor U28098 (N_28098,N_27739,N_27562);
xnor U28099 (N_28099,N_27760,N_27715);
and U28100 (N_28100,N_27527,N_27561);
nand U28101 (N_28101,N_27974,N_27755);
or U28102 (N_28102,N_27535,N_27678);
nand U28103 (N_28103,N_27507,N_27709);
and U28104 (N_28104,N_27674,N_27536);
and U28105 (N_28105,N_27803,N_27768);
and U28106 (N_28106,N_27605,N_27951);
or U28107 (N_28107,N_27742,N_27508);
xnor U28108 (N_28108,N_27845,N_27574);
nand U28109 (N_28109,N_27910,N_27829);
or U28110 (N_28110,N_27563,N_27975);
nand U28111 (N_28111,N_27553,N_27625);
xor U28112 (N_28112,N_27810,N_27997);
xor U28113 (N_28113,N_27581,N_27675);
nand U28114 (N_28114,N_27551,N_27773);
xor U28115 (N_28115,N_27856,N_27781);
or U28116 (N_28116,N_27725,N_27526);
nand U28117 (N_28117,N_27782,N_27640);
and U28118 (N_28118,N_27701,N_27771);
or U28119 (N_28119,N_27698,N_27877);
nor U28120 (N_28120,N_27635,N_27643);
xor U28121 (N_28121,N_27764,N_27662);
nor U28122 (N_28122,N_27629,N_27560);
or U28123 (N_28123,N_27700,N_27933);
or U28124 (N_28124,N_27667,N_27894);
and U28125 (N_28125,N_27616,N_27952);
xor U28126 (N_28126,N_27875,N_27549);
nor U28127 (N_28127,N_27607,N_27981);
nor U28128 (N_28128,N_27515,N_27668);
or U28129 (N_28129,N_27855,N_27708);
and U28130 (N_28130,N_27733,N_27573);
and U28131 (N_28131,N_27868,N_27841);
or U28132 (N_28132,N_27533,N_27797);
nor U28133 (N_28133,N_27785,N_27702);
and U28134 (N_28134,N_27887,N_27814);
or U28135 (N_28135,N_27517,N_27900);
xor U28136 (N_28136,N_27902,N_27820);
or U28137 (N_28137,N_27898,N_27879);
and U28138 (N_28138,N_27936,N_27890);
nor U28139 (N_28139,N_27688,N_27518);
or U28140 (N_28140,N_27921,N_27870);
xor U28141 (N_28141,N_27588,N_27885);
nand U28142 (N_28142,N_27649,N_27512);
xor U28143 (N_28143,N_27642,N_27853);
or U28144 (N_28144,N_27949,N_27669);
nand U28145 (N_28145,N_27964,N_27909);
nor U28146 (N_28146,N_27650,N_27631);
or U28147 (N_28147,N_27946,N_27547);
nand U28148 (N_28148,N_27586,N_27794);
and U28149 (N_28149,N_27858,N_27914);
nor U28150 (N_28150,N_27556,N_27808);
nor U28151 (N_28151,N_27938,N_27594);
and U28152 (N_28152,N_27995,N_27844);
nor U28153 (N_28153,N_27989,N_27843);
and U28154 (N_28154,N_27961,N_27652);
and U28155 (N_28155,N_27754,N_27998);
nor U28156 (N_28156,N_27509,N_27747);
nand U28157 (N_28157,N_27559,N_27718);
or U28158 (N_28158,N_27541,N_27908);
nor U28159 (N_28159,N_27791,N_27812);
and U28160 (N_28160,N_27622,N_27502);
nor U28161 (N_28161,N_27557,N_27685);
nor U28162 (N_28162,N_27990,N_27847);
nor U28163 (N_28163,N_27958,N_27593);
xnor U28164 (N_28164,N_27716,N_27726);
nand U28165 (N_28165,N_27720,N_27999);
xnor U28166 (N_28166,N_27653,N_27772);
nor U28167 (N_28167,N_27736,N_27646);
nor U28168 (N_28168,N_27996,N_27660);
nand U28169 (N_28169,N_27935,N_27673);
xor U28170 (N_28170,N_27857,N_27965);
or U28171 (N_28171,N_27766,N_27578);
or U28172 (N_28172,N_27751,N_27828);
nand U28173 (N_28173,N_27697,N_27786);
or U28174 (N_28174,N_27960,N_27866);
nor U28175 (N_28175,N_27703,N_27912);
nand U28176 (N_28176,N_27519,N_27907);
nor U28177 (N_28177,N_27884,N_27944);
nor U28178 (N_28178,N_27889,N_27656);
xnor U28179 (N_28179,N_27721,N_27687);
xor U28180 (N_28180,N_27795,N_27811);
and U28181 (N_28181,N_27723,N_27585);
nor U28182 (N_28182,N_27569,N_27651);
nor U28183 (N_28183,N_27544,N_27729);
nand U28184 (N_28184,N_27955,N_27722);
nand U28185 (N_28185,N_27619,N_27827);
or U28186 (N_28186,N_27510,N_27589);
nand U28187 (N_28187,N_27630,N_27542);
nor U28188 (N_28188,N_27600,N_27523);
or U28189 (N_28189,N_27724,N_27624);
and U28190 (N_28190,N_27712,N_27738);
and U28191 (N_28191,N_27596,N_27620);
or U28192 (N_28192,N_27836,N_27565);
or U28193 (N_28193,N_27988,N_27614);
and U28194 (N_28194,N_27695,N_27927);
xnor U28195 (N_28195,N_27876,N_27846);
nor U28196 (N_28196,N_27714,N_27530);
nor U28197 (N_28197,N_27500,N_27612);
nand U28198 (N_28198,N_27973,N_27859);
and U28199 (N_28199,N_27682,N_27972);
or U28200 (N_28200,N_27636,N_27555);
and U28201 (N_28201,N_27529,N_27699);
or U28202 (N_28202,N_27987,N_27893);
nor U28203 (N_28203,N_27647,N_27501);
nor U28204 (N_28204,N_27694,N_27765);
xor U28205 (N_28205,N_27787,N_27931);
xnor U28206 (N_28206,N_27839,N_27576);
nand U28207 (N_28207,N_27609,N_27621);
or U28208 (N_28208,N_27732,N_27849);
and U28209 (N_28209,N_27522,N_27901);
or U28210 (N_28210,N_27784,N_27603);
nand U28211 (N_28211,N_27758,N_27825);
xnor U28212 (N_28212,N_27730,N_27796);
nor U28213 (N_28213,N_27745,N_27956);
and U28214 (N_28214,N_27540,N_27628);
nand U28215 (N_28215,N_27980,N_27792);
nand U28216 (N_28216,N_27842,N_27528);
xor U28217 (N_28217,N_27591,N_27850);
nor U28218 (N_28218,N_27750,N_27978);
nand U28219 (N_28219,N_27626,N_27985);
nor U28220 (N_28220,N_27637,N_27537);
nand U28221 (N_28221,N_27819,N_27759);
xor U28222 (N_28222,N_27741,N_27613);
nor U28223 (N_28223,N_27753,N_27994);
or U28224 (N_28224,N_27583,N_27503);
nand U28225 (N_28225,N_27852,N_27538);
nor U28226 (N_28226,N_27871,N_27735);
xor U28227 (N_28227,N_27610,N_27945);
nor U28228 (N_28228,N_27575,N_27532);
and U28229 (N_28229,N_27757,N_27913);
and U28230 (N_28230,N_27599,N_27776);
nand U28231 (N_28231,N_27710,N_27867);
nor U28232 (N_28232,N_27778,N_27639);
xor U28233 (N_28233,N_27548,N_27918);
or U28234 (N_28234,N_27734,N_27991);
nand U28235 (N_28235,N_27671,N_27924);
nand U28236 (N_28236,N_27713,N_27881);
and U28237 (N_28237,N_27545,N_27748);
and U28238 (N_28238,N_27953,N_27680);
nand U28239 (N_28239,N_27805,N_27534);
and U28240 (N_28240,N_27899,N_27943);
and U28241 (N_28241,N_27670,N_27634);
or U28242 (N_28242,N_27993,N_27690);
nor U28243 (N_28243,N_27506,N_27728);
or U28244 (N_28244,N_27554,N_27979);
or U28245 (N_28245,N_27926,N_27950);
nand U28246 (N_28246,N_27779,N_27644);
nor U28247 (N_28247,N_27571,N_27743);
nand U28248 (N_28248,N_27807,N_27930);
and U28249 (N_28249,N_27848,N_27761);
xor U28250 (N_28250,N_27721,N_27995);
nand U28251 (N_28251,N_27722,N_27577);
nor U28252 (N_28252,N_27802,N_27722);
nand U28253 (N_28253,N_27941,N_27670);
or U28254 (N_28254,N_27567,N_27913);
and U28255 (N_28255,N_27837,N_27768);
and U28256 (N_28256,N_27690,N_27630);
nor U28257 (N_28257,N_27672,N_27983);
or U28258 (N_28258,N_27902,N_27726);
or U28259 (N_28259,N_27943,N_27848);
nand U28260 (N_28260,N_27674,N_27913);
nand U28261 (N_28261,N_27604,N_27766);
nand U28262 (N_28262,N_27504,N_27635);
and U28263 (N_28263,N_27942,N_27595);
or U28264 (N_28264,N_27978,N_27970);
nor U28265 (N_28265,N_27524,N_27708);
xor U28266 (N_28266,N_27937,N_27933);
or U28267 (N_28267,N_27898,N_27528);
or U28268 (N_28268,N_27785,N_27585);
nor U28269 (N_28269,N_27737,N_27861);
nor U28270 (N_28270,N_27748,N_27638);
nand U28271 (N_28271,N_27661,N_27517);
and U28272 (N_28272,N_27555,N_27909);
xnor U28273 (N_28273,N_27559,N_27911);
xnor U28274 (N_28274,N_27577,N_27900);
nand U28275 (N_28275,N_27993,N_27664);
or U28276 (N_28276,N_27870,N_27828);
nand U28277 (N_28277,N_27738,N_27573);
xnor U28278 (N_28278,N_27690,N_27973);
nand U28279 (N_28279,N_27786,N_27919);
nand U28280 (N_28280,N_27630,N_27661);
and U28281 (N_28281,N_27990,N_27546);
xor U28282 (N_28282,N_27535,N_27980);
and U28283 (N_28283,N_27997,N_27719);
nand U28284 (N_28284,N_27909,N_27960);
and U28285 (N_28285,N_27510,N_27556);
or U28286 (N_28286,N_27914,N_27682);
or U28287 (N_28287,N_27595,N_27726);
xnor U28288 (N_28288,N_27790,N_27599);
and U28289 (N_28289,N_27540,N_27899);
nor U28290 (N_28290,N_27580,N_27998);
and U28291 (N_28291,N_27924,N_27711);
xnor U28292 (N_28292,N_27890,N_27591);
or U28293 (N_28293,N_27536,N_27616);
nand U28294 (N_28294,N_27602,N_27692);
and U28295 (N_28295,N_27672,N_27902);
or U28296 (N_28296,N_27605,N_27658);
nor U28297 (N_28297,N_27773,N_27853);
nand U28298 (N_28298,N_27876,N_27637);
xnor U28299 (N_28299,N_27941,N_27809);
xnor U28300 (N_28300,N_27976,N_27504);
and U28301 (N_28301,N_27785,N_27986);
nand U28302 (N_28302,N_27892,N_27508);
xnor U28303 (N_28303,N_27727,N_27771);
and U28304 (N_28304,N_27727,N_27757);
nor U28305 (N_28305,N_27633,N_27889);
nor U28306 (N_28306,N_27947,N_27550);
nor U28307 (N_28307,N_27527,N_27562);
and U28308 (N_28308,N_27804,N_27612);
xor U28309 (N_28309,N_27667,N_27577);
and U28310 (N_28310,N_27504,N_27604);
xor U28311 (N_28311,N_27659,N_27663);
and U28312 (N_28312,N_27675,N_27928);
nor U28313 (N_28313,N_27769,N_27852);
or U28314 (N_28314,N_27875,N_27539);
xor U28315 (N_28315,N_27516,N_27675);
and U28316 (N_28316,N_27715,N_27844);
nand U28317 (N_28317,N_27855,N_27844);
or U28318 (N_28318,N_27677,N_27698);
nand U28319 (N_28319,N_27984,N_27744);
or U28320 (N_28320,N_27603,N_27535);
nand U28321 (N_28321,N_27717,N_27571);
nor U28322 (N_28322,N_27611,N_27894);
and U28323 (N_28323,N_27709,N_27596);
nor U28324 (N_28324,N_27877,N_27834);
or U28325 (N_28325,N_27809,N_27528);
xor U28326 (N_28326,N_27689,N_27998);
nand U28327 (N_28327,N_27717,N_27567);
xnor U28328 (N_28328,N_27829,N_27844);
or U28329 (N_28329,N_27849,N_27596);
nor U28330 (N_28330,N_27880,N_27524);
nor U28331 (N_28331,N_27897,N_27757);
nand U28332 (N_28332,N_27608,N_27935);
nor U28333 (N_28333,N_27501,N_27707);
nor U28334 (N_28334,N_27686,N_27953);
or U28335 (N_28335,N_27818,N_27827);
nand U28336 (N_28336,N_27939,N_27690);
or U28337 (N_28337,N_27690,N_27666);
or U28338 (N_28338,N_27905,N_27861);
nor U28339 (N_28339,N_27506,N_27758);
nor U28340 (N_28340,N_27855,N_27988);
or U28341 (N_28341,N_27549,N_27660);
or U28342 (N_28342,N_27774,N_27577);
nand U28343 (N_28343,N_27731,N_27521);
nor U28344 (N_28344,N_27734,N_27624);
xor U28345 (N_28345,N_27812,N_27765);
nand U28346 (N_28346,N_27517,N_27846);
nor U28347 (N_28347,N_27769,N_27896);
nand U28348 (N_28348,N_27907,N_27991);
nand U28349 (N_28349,N_27580,N_27788);
nor U28350 (N_28350,N_27703,N_27614);
nor U28351 (N_28351,N_27648,N_27775);
nand U28352 (N_28352,N_27693,N_27741);
nor U28353 (N_28353,N_27835,N_27577);
and U28354 (N_28354,N_27834,N_27980);
nor U28355 (N_28355,N_27501,N_27636);
or U28356 (N_28356,N_27749,N_27571);
nand U28357 (N_28357,N_27719,N_27658);
nand U28358 (N_28358,N_27911,N_27646);
and U28359 (N_28359,N_27822,N_27872);
or U28360 (N_28360,N_27522,N_27811);
xnor U28361 (N_28361,N_27942,N_27964);
nand U28362 (N_28362,N_27651,N_27742);
and U28363 (N_28363,N_27738,N_27741);
and U28364 (N_28364,N_27626,N_27810);
or U28365 (N_28365,N_27515,N_27591);
and U28366 (N_28366,N_27828,N_27634);
nand U28367 (N_28367,N_27889,N_27587);
xnor U28368 (N_28368,N_27761,N_27542);
nor U28369 (N_28369,N_27953,N_27685);
or U28370 (N_28370,N_27580,N_27857);
or U28371 (N_28371,N_27577,N_27948);
or U28372 (N_28372,N_27770,N_27709);
nand U28373 (N_28373,N_27872,N_27859);
or U28374 (N_28374,N_27777,N_27525);
or U28375 (N_28375,N_27854,N_27560);
xor U28376 (N_28376,N_27916,N_27539);
nand U28377 (N_28377,N_27766,N_27688);
nor U28378 (N_28378,N_27940,N_27719);
and U28379 (N_28379,N_27524,N_27546);
nor U28380 (N_28380,N_27990,N_27946);
or U28381 (N_28381,N_27894,N_27724);
and U28382 (N_28382,N_27870,N_27779);
nor U28383 (N_28383,N_27771,N_27645);
nor U28384 (N_28384,N_27772,N_27640);
or U28385 (N_28385,N_27900,N_27531);
nand U28386 (N_28386,N_27711,N_27615);
nand U28387 (N_28387,N_27527,N_27987);
xor U28388 (N_28388,N_27811,N_27553);
and U28389 (N_28389,N_27852,N_27735);
nand U28390 (N_28390,N_27927,N_27954);
or U28391 (N_28391,N_27932,N_27540);
nor U28392 (N_28392,N_27664,N_27968);
xor U28393 (N_28393,N_27813,N_27711);
or U28394 (N_28394,N_27677,N_27563);
or U28395 (N_28395,N_27906,N_27759);
xnor U28396 (N_28396,N_27723,N_27613);
xnor U28397 (N_28397,N_27665,N_27836);
xor U28398 (N_28398,N_27887,N_27921);
nand U28399 (N_28399,N_27911,N_27503);
xnor U28400 (N_28400,N_27551,N_27734);
or U28401 (N_28401,N_27629,N_27567);
xnor U28402 (N_28402,N_27917,N_27952);
nor U28403 (N_28403,N_27759,N_27655);
nand U28404 (N_28404,N_27693,N_27784);
nand U28405 (N_28405,N_27571,N_27601);
or U28406 (N_28406,N_27919,N_27569);
or U28407 (N_28407,N_27850,N_27902);
or U28408 (N_28408,N_27854,N_27616);
and U28409 (N_28409,N_27548,N_27980);
or U28410 (N_28410,N_27549,N_27748);
xnor U28411 (N_28411,N_27983,N_27665);
xor U28412 (N_28412,N_27766,N_27593);
and U28413 (N_28413,N_27685,N_27724);
or U28414 (N_28414,N_27670,N_27616);
nand U28415 (N_28415,N_27730,N_27666);
xnor U28416 (N_28416,N_27920,N_27873);
nand U28417 (N_28417,N_27561,N_27649);
nand U28418 (N_28418,N_27654,N_27876);
or U28419 (N_28419,N_27731,N_27766);
xor U28420 (N_28420,N_27594,N_27629);
nand U28421 (N_28421,N_27579,N_27700);
xnor U28422 (N_28422,N_27630,N_27699);
nand U28423 (N_28423,N_27520,N_27941);
or U28424 (N_28424,N_27555,N_27634);
nor U28425 (N_28425,N_27672,N_27859);
nand U28426 (N_28426,N_27775,N_27783);
nand U28427 (N_28427,N_27552,N_27716);
and U28428 (N_28428,N_27959,N_27632);
or U28429 (N_28429,N_27695,N_27530);
xnor U28430 (N_28430,N_27675,N_27916);
or U28431 (N_28431,N_27530,N_27857);
nor U28432 (N_28432,N_27819,N_27996);
nand U28433 (N_28433,N_27521,N_27728);
nand U28434 (N_28434,N_27608,N_27521);
xnor U28435 (N_28435,N_27941,N_27826);
or U28436 (N_28436,N_27817,N_27909);
and U28437 (N_28437,N_27886,N_27655);
nand U28438 (N_28438,N_27866,N_27766);
nand U28439 (N_28439,N_27659,N_27676);
nor U28440 (N_28440,N_27797,N_27566);
nor U28441 (N_28441,N_27748,N_27820);
xor U28442 (N_28442,N_27767,N_27618);
nor U28443 (N_28443,N_27927,N_27601);
nor U28444 (N_28444,N_27986,N_27903);
and U28445 (N_28445,N_27752,N_27674);
or U28446 (N_28446,N_27954,N_27786);
nand U28447 (N_28447,N_27978,N_27769);
nand U28448 (N_28448,N_27760,N_27635);
xor U28449 (N_28449,N_27673,N_27721);
xnor U28450 (N_28450,N_27796,N_27722);
xor U28451 (N_28451,N_27869,N_27550);
nor U28452 (N_28452,N_27867,N_27885);
nand U28453 (N_28453,N_27637,N_27783);
and U28454 (N_28454,N_27582,N_27862);
xor U28455 (N_28455,N_27797,N_27952);
xor U28456 (N_28456,N_27552,N_27803);
nor U28457 (N_28457,N_27833,N_27923);
and U28458 (N_28458,N_27881,N_27821);
or U28459 (N_28459,N_27654,N_27661);
or U28460 (N_28460,N_27572,N_27918);
nor U28461 (N_28461,N_27655,N_27914);
and U28462 (N_28462,N_27983,N_27752);
nand U28463 (N_28463,N_27855,N_27525);
or U28464 (N_28464,N_27530,N_27840);
xor U28465 (N_28465,N_27603,N_27823);
nor U28466 (N_28466,N_27501,N_27976);
nor U28467 (N_28467,N_27937,N_27854);
nand U28468 (N_28468,N_27624,N_27554);
xor U28469 (N_28469,N_27503,N_27886);
nand U28470 (N_28470,N_27649,N_27788);
nand U28471 (N_28471,N_27532,N_27760);
or U28472 (N_28472,N_27925,N_27732);
and U28473 (N_28473,N_27748,N_27812);
or U28474 (N_28474,N_27755,N_27745);
nand U28475 (N_28475,N_27864,N_27509);
nor U28476 (N_28476,N_27801,N_27557);
xor U28477 (N_28477,N_27777,N_27625);
nor U28478 (N_28478,N_27892,N_27978);
or U28479 (N_28479,N_27537,N_27738);
xor U28480 (N_28480,N_27515,N_27657);
nor U28481 (N_28481,N_27811,N_27862);
nand U28482 (N_28482,N_27933,N_27525);
nor U28483 (N_28483,N_27914,N_27728);
or U28484 (N_28484,N_27541,N_27514);
or U28485 (N_28485,N_27564,N_27755);
or U28486 (N_28486,N_27938,N_27877);
nor U28487 (N_28487,N_27585,N_27686);
or U28488 (N_28488,N_27952,N_27716);
or U28489 (N_28489,N_27992,N_27706);
xor U28490 (N_28490,N_27786,N_27685);
xnor U28491 (N_28491,N_27905,N_27719);
and U28492 (N_28492,N_27775,N_27562);
and U28493 (N_28493,N_27539,N_27901);
nor U28494 (N_28494,N_27703,N_27517);
nand U28495 (N_28495,N_27549,N_27638);
nand U28496 (N_28496,N_27988,N_27677);
xor U28497 (N_28497,N_27645,N_27516);
xor U28498 (N_28498,N_27934,N_27841);
nand U28499 (N_28499,N_27682,N_27564);
nor U28500 (N_28500,N_28026,N_28310);
nand U28501 (N_28501,N_28020,N_28126);
nand U28502 (N_28502,N_28340,N_28034);
nor U28503 (N_28503,N_28191,N_28050);
and U28504 (N_28504,N_28183,N_28291);
and U28505 (N_28505,N_28012,N_28290);
nand U28506 (N_28506,N_28145,N_28348);
nand U28507 (N_28507,N_28327,N_28159);
xnor U28508 (N_28508,N_28392,N_28429);
nor U28509 (N_28509,N_28275,N_28390);
or U28510 (N_28510,N_28141,N_28023);
xnor U28511 (N_28511,N_28323,N_28198);
or U28512 (N_28512,N_28060,N_28481);
and U28513 (N_28513,N_28421,N_28367);
or U28514 (N_28514,N_28425,N_28428);
xor U28515 (N_28515,N_28469,N_28068);
nand U28516 (N_28516,N_28160,N_28167);
nand U28517 (N_28517,N_28357,N_28358);
xor U28518 (N_28518,N_28250,N_28240);
nor U28519 (N_28519,N_28235,N_28248);
and U28520 (N_28520,N_28402,N_28157);
and U28521 (N_28521,N_28496,N_28094);
nand U28522 (N_28522,N_28144,N_28150);
nand U28523 (N_28523,N_28405,N_28093);
nand U28524 (N_28524,N_28032,N_28387);
and U28525 (N_28525,N_28484,N_28115);
nand U28526 (N_28526,N_28133,N_28437);
or U28527 (N_28527,N_28120,N_28128);
and U28528 (N_28528,N_28081,N_28065);
nand U28529 (N_28529,N_28307,N_28097);
or U28530 (N_28530,N_28360,N_28488);
nor U28531 (N_28531,N_28018,N_28001);
and U28532 (N_28532,N_28195,N_28478);
or U28533 (N_28533,N_28100,N_28146);
and U28534 (N_28534,N_28113,N_28444);
and U28535 (N_28535,N_28336,N_28422);
nor U28536 (N_28536,N_28276,N_28021);
nor U28537 (N_28537,N_28420,N_28416);
xnor U28538 (N_28538,N_28401,N_28349);
or U28539 (N_28539,N_28197,N_28089);
xor U28540 (N_28540,N_28326,N_28272);
or U28541 (N_28541,N_28102,N_28029);
and U28542 (N_28542,N_28062,N_28077);
nand U28543 (N_28543,N_28281,N_28019);
nor U28544 (N_28544,N_28121,N_28229);
nor U28545 (N_28545,N_28479,N_28284);
or U28546 (N_28546,N_28136,N_28178);
nand U28547 (N_28547,N_28361,N_28118);
and U28548 (N_28548,N_28389,N_28005);
nor U28549 (N_28549,N_28066,N_28354);
nor U28550 (N_28550,N_28155,N_28236);
nor U28551 (N_28551,N_28043,N_28038);
xnor U28552 (N_28552,N_28449,N_28329);
and U28553 (N_28553,N_28110,N_28364);
nor U28554 (N_28554,N_28243,N_28302);
and U28555 (N_28555,N_28423,N_28024);
or U28556 (N_28556,N_28164,N_28414);
or U28557 (N_28557,N_28378,N_28088);
nand U28558 (N_28558,N_28177,N_28438);
nand U28559 (N_28559,N_28186,N_28385);
nand U28560 (N_28560,N_28245,N_28173);
xnor U28561 (N_28561,N_28418,N_28015);
xor U28562 (N_28562,N_28296,N_28440);
xor U28563 (N_28563,N_28413,N_28069);
nor U28564 (N_28564,N_28111,N_28063);
or U28565 (N_28565,N_28239,N_28176);
nor U28566 (N_28566,N_28084,N_28353);
or U28567 (N_28567,N_28473,N_28158);
nor U28568 (N_28568,N_28230,N_28028);
nor U28569 (N_28569,N_28388,N_28036);
and U28570 (N_28570,N_28218,N_28199);
nand U28571 (N_28571,N_28080,N_28295);
and U28572 (N_28572,N_28451,N_28262);
xnor U28573 (N_28573,N_28112,N_28461);
or U28574 (N_28574,N_28312,N_28242);
nand U28575 (N_28575,N_28187,N_28285);
nand U28576 (N_28576,N_28274,N_28193);
nand U28577 (N_28577,N_28007,N_28134);
nor U28578 (N_28578,N_28182,N_28376);
nand U28579 (N_28579,N_28225,N_28249);
xnor U28580 (N_28580,N_28202,N_28256);
and U28581 (N_28581,N_28303,N_28000);
nor U28582 (N_28582,N_28424,N_28417);
or U28583 (N_28583,N_28099,N_28064);
or U28584 (N_28584,N_28338,N_28237);
or U28585 (N_28585,N_28053,N_28471);
and U28586 (N_28586,N_28466,N_28127);
and U28587 (N_28587,N_28131,N_28465);
and U28588 (N_28588,N_28170,N_28044);
or U28589 (N_28589,N_28238,N_28103);
nor U28590 (N_28590,N_28221,N_28482);
or U28591 (N_28591,N_28076,N_28233);
or U28592 (N_28592,N_28072,N_28278);
nand U28593 (N_28593,N_28459,N_28228);
nor U28594 (N_28594,N_28129,N_28171);
xnor U28595 (N_28595,N_28075,N_28495);
or U28596 (N_28596,N_28209,N_28101);
or U28597 (N_28597,N_28460,N_28351);
nor U28598 (N_28598,N_28445,N_28122);
nand U28599 (N_28599,N_28286,N_28332);
nor U28600 (N_28600,N_28253,N_28415);
xnor U28601 (N_28601,N_28013,N_28404);
nor U28602 (N_28602,N_28067,N_28244);
xnor U28603 (N_28603,N_28304,N_28396);
nor U28604 (N_28604,N_28092,N_28457);
xor U28605 (N_28605,N_28047,N_28061);
and U28606 (N_28606,N_28095,N_28319);
xnor U28607 (N_28607,N_28328,N_28048);
xnor U28608 (N_28608,N_28030,N_28430);
nor U28609 (N_28609,N_28306,N_28395);
nor U28610 (N_28610,N_28027,N_28411);
and U28611 (N_28611,N_28222,N_28251);
and U28612 (N_28612,N_28317,N_28365);
or U28613 (N_28613,N_28431,N_28282);
nand U28614 (N_28614,N_28375,N_28196);
or U28615 (N_28615,N_28476,N_28483);
nor U28616 (N_28616,N_28217,N_28189);
nand U28617 (N_28617,N_28107,N_28079);
nand U28618 (N_28618,N_28241,N_28419);
and U28619 (N_28619,N_28450,N_28246);
nor U28620 (N_28620,N_28070,N_28147);
and U28621 (N_28621,N_28059,N_28381);
and U28622 (N_28622,N_28258,N_28016);
and U28623 (N_28623,N_28152,N_28309);
and U28624 (N_28624,N_28305,N_28223);
nand U28625 (N_28625,N_28379,N_28403);
nand U28626 (N_28626,N_28316,N_28219);
xnor U28627 (N_28627,N_28138,N_28252);
or U28628 (N_28628,N_28394,N_28114);
and U28629 (N_28629,N_28435,N_28458);
or U28630 (N_28630,N_28022,N_28453);
and U28631 (N_28631,N_28398,N_28382);
nor U28632 (N_28632,N_28267,N_28393);
nand U28633 (N_28633,N_28434,N_28071);
and U28634 (N_28634,N_28301,N_28494);
or U28635 (N_28635,N_28330,N_28117);
nor U28636 (N_28636,N_28298,N_28498);
nor U28637 (N_28637,N_28266,N_28049);
and U28638 (N_28638,N_28490,N_28003);
and U28639 (N_28639,N_28083,N_28412);
nand U28640 (N_28640,N_28492,N_28359);
nand U28641 (N_28641,N_28087,N_28212);
nand U28642 (N_28642,N_28265,N_28192);
or U28643 (N_28643,N_28078,N_28172);
nand U28644 (N_28644,N_28057,N_28470);
nand U28645 (N_28645,N_28369,N_28355);
xor U28646 (N_28646,N_28485,N_28487);
nand U28647 (N_28647,N_28210,N_28188);
nor U28648 (N_28648,N_28427,N_28194);
nor U28649 (N_28649,N_28153,N_28148);
and U28650 (N_28650,N_28407,N_28497);
and U28651 (N_28651,N_28366,N_28255);
nand U28652 (N_28652,N_28090,N_28154);
or U28653 (N_28653,N_28311,N_28308);
and U28654 (N_28654,N_28464,N_28106);
nand U28655 (N_28655,N_28283,N_28216);
xnor U28656 (N_28656,N_28037,N_28335);
nand U28657 (N_28657,N_28104,N_28264);
nand U28658 (N_28658,N_28313,N_28124);
xor U28659 (N_28659,N_28175,N_28139);
nor U28660 (N_28660,N_28039,N_28207);
nand U28661 (N_28661,N_28333,N_28014);
nand U28662 (N_28662,N_28343,N_28091);
or U28663 (N_28663,N_28374,N_28108);
or U28664 (N_28664,N_28324,N_28004);
nand U28665 (N_28665,N_28321,N_28181);
nor U28666 (N_28666,N_28455,N_28206);
and U28667 (N_28667,N_28074,N_28475);
or U28668 (N_28668,N_28214,N_28010);
nand U28669 (N_28669,N_28205,N_28085);
or U28670 (N_28670,N_28149,N_28273);
nand U28671 (N_28671,N_28344,N_28371);
and U28672 (N_28672,N_28468,N_28271);
xor U28673 (N_28673,N_28140,N_28399);
nand U28674 (N_28674,N_28372,N_28169);
nand U28675 (N_28675,N_28098,N_28287);
and U28676 (N_28676,N_28345,N_28315);
nand U28677 (N_28677,N_28185,N_28463);
nand U28678 (N_28678,N_28368,N_28356);
nor U28679 (N_28679,N_28200,N_28439);
and U28680 (N_28680,N_28082,N_28052);
nor U28681 (N_28681,N_28017,N_28448);
and U28682 (N_28682,N_28269,N_28161);
and U28683 (N_28683,N_28130,N_28341);
xnor U28684 (N_28684,N_28289,N_28190);
nor U28685 (N_28685,N_28096,N_28163);
and U28686 (N_28686,N_28268,N_28204);
xor U28687 (N_28687,N_28179,N_28474);
nor U28688 (N_28688,N_28409,N_28493);
and U28689 (N_28689,N_28334,N_28105);
and U28690 (N_28690,N_28215,N_28031);
nand U28691 (N_28691,N_28480,N_28132);
nand U28692 (N_28692,N_28446,N_28119);
xor U28693 (N_28693,N_28410,N_28362);
nand U28694 (N_28694,N_28035,N_28055);
nor U28695 (N_28695,N_28432,N_28033);
xnor U28696 (N_28696,N_28383,N_28442);
or U28697 (N_28697,N_28297,N_28135);
nor U28698 (N_28698,N_28447,N_28180);
nor U28699 (N_28699,N_28318,N_28350);
and U28700 (N_28700,N_28456,N_28292);
nor U28701 (N_28701,N_28234,N_28211);
or U28702 (N_28702,N_28009,N_28168);
nor U28703 (N_28703,N_28352,N_28280);
xor U28704 (N_28704,N_28254,N_28257);
xor U28705 (N_28705,N_28486,N_28184);
or U28706 (N_28706,N_28051,N_28300);
and U28707 (N_28707,N_28040,N_28325);
nand U28708 (N_28708,N_28046,N_28322);
nor U28709 (N_28709,N_28008,N_28041);
xor U28710 (N_28710,N_28156,N_28116);
xor U28711 (N_28711,N_28166,N_28220);
nor U28712 (N_28712,N_28086,N_28489);
nand U28713 (N_28713,N_28441,N_28231);
or U28714 (N_28714,N_28433,N_28143);
and U28715 (N_28715,N_28056,N_28443);
and U28716 (N_28716,N_28386,N_28462);
nor U28717 (N_28717,N_28397,N_28400);
xnor U28718 (N_28718,N_28142,N_28314);
or U28719 (N_28719,N_28226,N_28045);
xor U28720 (N_28720,N_28261,N_28213);
xnor U28721 (N_28721,N_28011,N_28260);
or U28722 (N_28722,N_28277,N_28002);
and U28723 (N_28723,N_28042,N_28279);
nor U28724 (N_28724,N_28224,N_28203);
xor U28725 (N_28725,N_28299,N_28337);
or U28726 (N_28726,N_28054,N_28436);
or U28727 (N_28727,N_28377,N_28151);
nand U28728 (N_28728,N_28123,N_28293);
xnor U28729 (N_28729,N_28232,N_28006);
nand U28730 (N_28730,N_28346,N_28294);
and U28731 (N_28731,N_28259,N_28270);
and U28732 (N_28732,N_28347,N_28125);
xor U28733 (N_28733,N_28165,N_28342);
xor U28734 (N_28734,N_28499,N_28025);
xor U28735 (N_28735,N_28452,N_28477);
or U28736 (N_28736,N_28201,N_28391);
or U28737 (N_28737,N_28331,N_28454);
and U28738 (N_28738,N_28363,N_28467);
nand U28739 (N_28739,N_28073,N_28227);
xor U28740 (N_28740,N_28380,N_28320);
or U28741 (N_28741,N_28263,N_28370);
nand U28742 (N_28742,N_28208,N_28408);
and U28743 (N_28743,N_28426,N_28058);
or U28744 (N_28744,N_28472,N_28174);
and U28745 (N_28745,N_28406,N_28373);
nand U28746 (N_28746,N_28247,N_28162);
or U28747 (N_28747,N_28288,N_28491);
nor U28748 (N_28748,N_28109,N_28137);
nand U28749 (N_28749,N_28384,N_28339);
and U28750 (N_28750,N_28092,N_28354);
and U28751 (N_28751,N_28379,N_28310);
or U28752 (N_28752,N_28366,N_28232);
xor U28753 (N_28753,N_28140,N_28287);
or U28754 (N_28754,N_28142,N_28448);
or U28755 (N_28755,N_28046,N_28311);
or U28756 (N_28756,N_28307,N_28028);
nor U28757 (N_28757,N_28318,N_28243);
nand U28758 (N_28758,N_28187,N_28332);
or U28759 (N_28759,N_28042,N_28217);
xnor U28760 (N_28760,N_28088,N_28157);
xnor U28761 (N_28761,N_28211,N_28229);
or U28762 (N_28762,N_28034,N_28462);
and U28763 (N_28763,N_28104,N_28180);
nand U28764 (N_28764,N_28217,N_28309);
nor U28765 (N_28765,N_28122,N_28124);
or U28766 (N_28766,N_28336,N_28106);
or U28767 (N_28767,N_28158,N_28121);
xnor U28768 (N_28768,N_28451,N_28427);
nor U28769 (N_28769,N_28452,N_28057);
or U28770 (N_28770,N_28082,N_28499);
or U28771 (N_28771,N_28275,N_28036);
or U28772 (N_28772,N_28235,N_28121);
xnor U28773 (N_28773,N_28024,N_28388);
and U28774 (N_28774,N_28231,N_28030);
xnor U28775 (N_28775,N_28468,N_28116);
nor U28776 (N_28776,N_28233,N_28146);
or U28777 (N_28777,N_28179,N_28212);
nand U28778 (N_28778,N_28241,N_28032);
nand U28779 (N_28779,N_28438,N_28319);
nor U28780 (N_28780,N_28219,N_28395);
or U28781 (N_28781,N_28292,N_28040);
nor U28782 (N_28782,N_28020,N_28437);
nor U28783 (N_28783,N_28279,N_28308);
or U28784 (N_28784,N_28222,N_28073);
nor U28785 (N_28785,N_28135,N_28231);
xor U28786 (N_28786,N_28191,N_28069);
nor U28787 (N_28787,N_28128,N_28428);
nor U28788 (N_28788,N_28210,N_28211);
xor U28789 (N_28789,N_28343,N_28445);
or U28790 (N_28790,N_28181,N_28315);
and U28791 (N_28791,N_28404,N_28144);
nor U28792 (N_28792,N_28448,N_28042);
and U28793 (N_28793,N_28386,N_28140);
nand U28794 (N_28794,N_28456,N_28167);
xor U28795 (N_28795,N_28291,N_28378);
or U28796 (N_28796,N_28099,N_28341);
nor U28797 (N_28797,N_28028,N_28193);
nor U28798 (N_28798,N_28041,N_28005);
nand U28799 (N_28799,N_28396,N_28369);
nand U28800 (N_28800,N_28451,N_28219);
or U28801 (N_28801,N_28196,N_28360);
or U28802 (N_28802,N_28450,N_28368);
nand U28803 (N_28803,N_28220,N_28173);
nor U28804 (N_28804,N_28392,N_28027);
or U28805 (N_28805,N_28227,N_28368);
and U28806 (N_28806,N_28047,N_28360);
or U28807 (N_28807,N_28425,N_28377);
or U28808 (N_28808,N_28421,N_28032);
and U28809 (N_28809,N_28294,N_28329);
nand U28810 (N_28810,N_28485,N_28151);
xor U28811 (N_28811,N_28499,N_28100);
xnor U28812 (N_28812,N_28456,N_28374);
xor U28813 (N_28813,N_28277,N_28013);
nor U28814 (N_28814,N_28252,N_28304);
or U28815 (N_28815,N_28110,N_28036);
nand U28816 (N_28816,N_28182,N_28485);
nand U28817 (N_28817,N_28068,N_28422);
nand U28818 (N_28818,N_28099,N_28232);
xor U28819 (N_28819,N_28484,N_28163);
xor U28820 (N_28820,N_28054,N_28046);
or U28821 (N_28821,N_28325,N_28367);
or U28822 (N_28822,N_28040,N_28340);
nand U28823 (N_28823,N_28157,N_28333);
xnor U28824 (N_28824,N_28316,N_28265);
or U28825 (N_28825,N_28027,N_28470);
or U28826 (N_28826,N_28207,N_28051);
and U28827 (N_28827,N_28332,N_28305);
and U28828 (N_28828,N_28170,N_28448);
or U28829 (N_28829,N_28206,N_28237);
nand U28830 (N_28830,N_28499,N_28359);
xor U28831 (N_28831,N_28084,N_28415);
and U28832 (N_28832,N_28210,N_28171);
or U28833 (N_28833,N_28117,N_28096);
and U28834 (N_28834,N_28149,N_28117);
nor U28835 (N_28835,N_28254,N_28481);
nand U28836 (N_28836,N_28125,N_28286);
nand U28837 (N_28837,N_28305,N_28010);
xor U28838 (N_28838,N_28274,N_28270);
or U28839 (N_28839,N_28441,N_28040);
and U28840 (N_28840,N_28412,N_28387);
xor U28841 (N_28841,N_28237,N_28137);
nand U28842 (N_28842,N_28227,N_28437);
nand U28843 (N_28843,N_28280,N_28174);
or U28844 (N_28844,N_28430,N_28117);
nor U28845 (N_28845,N_28106,N_28198);
xor U28846 (N_28846,N_28363,N_28348);
xor U28847 (N_28847,N_28038,N_28154);
and U28848 (N_28848,N_28093,N_28229);
xnor U28849 (N_28849,N_28138,N_28416);
nor U28850 (N_28850,N_28423,N_28458);
xor U28851 (N_28851,N_28395,N_28019);
nand U28852 (N_28852,N_28206,N_28438);
and U28853 (N_28853,N_28379,N_28241);
nor U28854 (N_28854,N_28151,N_28084);
nand U28855 (N_28855,N_28479,N_28143);
or U28856 (N_28856,N_28201,N_28016);
nand U28857 (N_28857,N_28250,N_28261);
nor U28858 (N_28858,N_28375,N_28228);
or U28859 (N_28859,N_28287,N_28124);
and U28860 (N_28860,N_28341,N_28222);
nor U28861 (N_28861,N_28260,N_28054);
or U28862 (N_28862,N_28113,N_28399);
or U28863 (N_28863,N_28091,N_28480);
and U28864 (N_28864,N_28084,N_28221);
nand U28865 (N_28865,N_28484,N_28388);
and U28866 (N_28866,N_28209,N_28323);
xnor U28867 (N_28867,N_28435,N_28398);
nor U28868 (N_28868,N_28467,N_28309);
or U28869 (N_28869,N_28376,N_28417);
and U28870 (N_28870,N_28041,N_28241);
or U28871 (N_28871,N_28271,N_28404);
and U28872 (N_28872,N_28373,N_28356);
and U28873 (N_28873,N_28035,N_28285);
xor U28874 (N_28874,N_28211,N_28228);
nand U28875 (N_28875,N_28129,N_28405);
or U28876 (N_28876,N_28340,N_28342);
and U28877 (N_28877,N_28281,N_28283);
nor U28878 (N_28878,N_28047,N_28215);
or U28879 (N_28879,N_28105,N_28024);
and U28880 (N_28880,N_28168,N_28087);
and U28881 (N_28881,N_28166,N_28054);
and U28882 (N_28882,N_28164,N_28057);
nor U28883 (N_28883,N_28122,N_28177);
xor U28884 (N_28884,N_28332,N_28474);
xor U28885 (N_28885,N_28091,N_28332);
nand U28886 (N_28886,N_28276,N_28147);
and U28887 (N_28887,N_28211,N_28272);
and U28888 (N_28888,N_28498,N_28438);
nand U28889 (N_28889,N_28349,N_28265);
nand U28890 (N_28890,N_28285,N_28380);
and U28891 (N_28891,N_28348,N_28465);
nor U28892 (N_28892,N_28131,N_28115);
nor U28893 (N_28893,N_28028,N_28005);
nand U28894 (N_28894,N_28081,N_28340);
or U28895 (N_28895,N_28365,N_28462);
nor U28896 (N_28896,N_28055,N_28153);
and U28897 (N_28897,N_28304,N_28014);
xnor U28898 (N_28898,N_28130,N_28226);
xor U28899 (N_28899,N_28000,N_28328);
nand U28900 (N_28900,N_28474,N_28122);
and U28901 (N_28901,N_28120,N_28102);
xnor U28902 (N_28902,N_28447,N_28409);
or U28903 (N_28903,N_28437,N_28420);
and U28904 (N_28904,N_28157,N_28349);
or U28905 (N_28905,N_28185,N_28437);
and U28906 (N_28906,N_28327,N_28497);
nor U28907 (N_28907,N_28224,N_28287);
and U28908 (N_28908,N_28218,N_28217);
nor U28909 (N_28909,N_28285,N_28228);
and U28910 (N_28910,N_28079,N_28466);
or U28911 (N_28911,N_28091,N_28335);
and U28912 (N_28912,N_28498,N_28142);
xnor U28913 (N_28913,N_28295,N_28340);
or U28914 (N_28914,N_28184,N_28203);
or U28915 (N_28915,N_28085,N_28107);
nor U28916 (N_28916,N_28418,N_28452);
xor U28917 (N_28917,N_28160,N_28086);
or U28918 (N_28918,N_28117,N_28226);
nand U28919 (N_28919,N_28197,N_28228);
or U28920 (N_28920,N_28472,N_28397);
xor U28921 (N_28921,N_28229,N_28461);
xnor U28922 (N_28922,N_28048,N_28212);
xor U28923 (N_28923,N_28094,N_28178);
nand U28924 (N_28924,N_28287,N_28475);
xnor U28925 (N_28925,N_28215,N_28377);
or U28926 (N_28926,N_28495,N_28378);
xnor U28927 (N_28927,N_28137,N_28448);
nand U28928 (N_28928,N_28387,N_28175);
and U28929 (N_28929,N_28169,N_28277);
xnor U28930 (N_28930,N_28327,N_28133);
or U28931 (N_28931,N_28412,N_28155);
nor U28932 (N_28932,N_28008,N_28011);
xnor U28933 (N_28933,N_28224,N_28351);
and U28934 (N_28934,N_28087,N_28452);
and U28935 (N_28935,N_28313,N_28423);
nor U28936 (N_28936,N_28086,N_28233);
nor U28937 (N_28937,N_28202,N_28038);
or U28938 (N_28938,N_28013,N_28158);
nand U28939 (N_28939,N_28320,N_28495);
nor U28940 (N_28940,N_28193,N_28114);
xnor U28941 (N_28941,N_28218,N_28126);
nand U28942 (N_28942,N_28036,N_28452);
nor U28943 (N_28943,N_28190,N_28218);
nand U28944 (N_28944,N_28357,N_28435);
and U28945 (N_28945,N_28291,N_28418);
and U28946 (N_28946,N_28066,N_28290);
or U28947 (N_28947,N_28308,N_28352);
nand U28948 (N_28948,N_28177,N_28090);
and U28949 (N_28949,N_28215,N_28200);
xnor U28950 (N_28950,N_28232,N_28026);
nand U28951 (N_28951,N_28373,N_28000);
xor U28952 (N_28952,N_28090,N_28105);
nand U28953 (N_28953,N_28082,N_28312);
nand U28954 (N_28954,N_28093,N_28356);
nand U28955 (N_28955,N_28292,N_28331);
nand U28956 (N_28956,N_28089,N_28007);
nor U28957 (N_28957,N_28089,N_28386);
and U28958 (N_28958,N_28364,N_28332);
xor U28959 (N_28959,N_28186,N_28259);
xor U28960 (N_28960,N_28102,N_28068);
xnor U28961 (N_28961,N_28257,N_28025);
nor U28962 (N_28962,N_28046,N_28095);
nor U28963 (N_28963,N_28403,N_28290);
and U28964 (N_28964,N_28494,N_28417);
xor U28965 (N_28965,N_28080,N_28399);
xnor U28966 (N_28966,N_28314,N_28326);
and U28967 (N_28967,N_28449,N_28385);
or U28968 (N_28968,N_28189,N_28127);
or U28969 (N_28969,N_28019,N_28253);
or U28970 (N_28970,N_28288,N_28287);
nor U28971 (N_28971,N_28034,N_28226);
nor U28972 (N_28972,N_28213,N_28094);
nor U28973 (N_28973,N_28419,N_28299);
nor U28974 (N_28974,N_28065,N_28019);
or U28975 (N_28975,N_28368,N_28385);
xor U28976 (N_28976,N_28183,N_28024);
nor U28977 (N_28977,N_28084,N_28187);
nand U28978 (N_28978,N_28233,N_28136);
nor U28979 (N_28979,N_28258,N_28099);
xnor U28980 (N_28980,N_28365,N_28036);
nand U28981 (N_28981,N_28186,N_28404);
nor U28982 (N_28982,N_28123,N_28010);
xnor U28983 (N_28983,N_28051,N_28255);
nand U28984 (N_28984,N_28429,N_28329);
or U28985 (N_28985,N_28443,N_28060);
or U28986 (N_28986,N_28175,N_28334);
xor U28987 (N_28987,N_28305,N_28012);
xor U28988 (N_28988,N_28198,N_28125);
and U28989 (N_28989,N_28412,N_28088);
xor U28990 (N_28990,N_28127,N_28359);
xnor U28991 (N_28991,N_28451,N_28287);
nor U28992 (N_28992,N_28167,N_28482);
nor U28993 (N_28993,N_28051,N_28474);
nand U28994 (N_28994,N_28226,N_28264);
xnor U28995 (N_28995,N_28152,N_28024);
and U28996 (N_28996,N_28071,N_28255);
nand U28997 (N_28997,N_28499,N_28172);
and U28998 (N_28998,N_28013,N_28264);
and U28999 (N_28999,N_28072,N_28322);
nor U29000 (N_29000,N_28972,N_28830);
xor U29001 (N_29001,N_28825,N_28881);
and U29002 (N_29002,N_28517,N_28924);
xnor U29003 (N_29003,N_28501,N_28723);
xnor U29004 (N_29004,N_28533,N_28522);
and U29005 (N_29005,N_28564,N_28959);
or U29006 (N_29006,N_28795,N_28935);
and U29007 (N_29007,N_28856,N_28728);
nor U29008 (N_29008,N_28609,N_28668);
xnor U29009 (N_29009,N_28610,N_28908);
nand U29010 (N_29010,N_28743,N_28587);
xor U29011 (N_29011,N_28513,N_28799);
nor U29012 (N_29012,N_28787,N_28788);
nor U29013 (N_29013,N_28640,N_28709);
nor U29014 (N_29014,N_28819,N_28714);
nor U29015 (N_29015,N_28572,N_28603);
nand U29016 (N_29016,N_28551,N_28857);
or U29017 (N_29017,N_28689,N_28629);
nor U29018 (N_29018,N_28654,N_28778);
and U29019 (N_29019,N_28917,N_28535);
nor U29020 (N_29020,N_28984,N_28641);
nand U29021 (N_29021,N_28593,N_28910);
xnor U29022 (N_29022,N_28636,N_28814);
nor U29023 (N_29023,N_28979,N_28659);
and U29024 (N_29024,N_28866,N_28744);
nor U29025 (N_29025,N_28573,N_28800);
nand U29026 (N_29026,N_28763,N_28941);
or U29027 (N_29027,N_28889,N_28607);
xor U29028 (N_29028,N_28504,N_28567);
or U29029 (N_29029,N_28677,N_28989);
xnor U29030 (N_29030,N_28975,N_28988);
or U29031 (N_29031,N_28638,N_28818);
xor U29032 (N_29032,N_28813,N_28530);
nand U29033 (N_29033,N_28816,N_28859);
nand U29034 (N_29034,N_28927,N_28536);
xor U29035 (N_29035,N_28971,N_28934);
or U29036 (N_29036,N_28582,N_28698);
and U29037 (N_29037,N_28790,N_28700);
xor U29038 (N_29038,N_28751,N_28727);
and U29039 (N_29039,N_28597,N_28735);
nor U29040 (N_29040,N_28688,N_28733);
xnor U29041 (N_29041,N_28717,N_28683);
nor U29042 (N_29042,N_28652,N_28999);
xnor U29043 (N_29043,N_28899,N_28938);
nor U29044 (N_29044,N_28948,N_28754);
xor U29045 (N_29045,N_28594,N_28949);
nor U29046 (N_29046,N_28792,N_28973);
xnor U29047 (N_29047,N_28651,N_28841);
or U29048 (N_29048,N_28863,N_28645);
nand U29049 (N_29049,N_28514,N_28552);
xnor U29050 (N_29050,N_28621,N_28703);
nand U29051 (N_29051,N_28776,N_28905);
or U29052 (N_29052,N_28696,N_28561);
nand U29053 (N_29053,N_28872,N_28851);
nor U29054 (N_29054,N_28721,N_28581);
xnor U29055 (N_29055,N_28690,N_28920);
xnor U29056 (N_29056,N_28674,N_28632);
and U29057 (N_29057,N_28981,N_28749);
xor U29058 (N_29058,N_28624,N_28817);
and U29059 (N_29059,N_28590,N_28642);
xor U29060 (N_29060,N_28794,N_28967);
xor U29061 (N_29061,N_28962,N_28619);
xnor U29062 (N_29062,N_28879,N_28867);
and U29063 (N_29063,N_28676,N_28943);
xnor U29064 (N_29064,N_28767,N_28635);
or U29065 (N_29065,N_28848,N_28861);
xor U29066 (N_29066,N_28606,N_28906);
xor U29067 (N_29067,N_28604,N_28970);
or U29068 (N_29068,N_28930,N_28528);
nand U29069 (N_29069,N_28832,N_28876);
or U29070 (N_29070,N_28768,N_28901);
xor U29071 (N_29071,N_28770,N_28686);
and U29072 (N_29072,N_28831,N_28664);
and U29073 (N_29073,N_28873,N_28803);
or U29074 (N_29074,N_28571,N_28942);
xor U29075 (N_29075,N_28622,N_28715);
nor U29076 (N_29076,N_28968,N_28925);
nand U29077 (N_29077,N_28783,N_28961);
nand U29078 (N_29078,N_28769,N_28534);
and U29079 (N_29079,N_28804,N_28998);
nor U29080 (N_29080,N_28570,N_28592);
xnor U29081 (N_29081,N_28560,N_28978);
nor U29082 (N_29082,N_28837,N_28780);
nor U29083 (N_29083,N_28982,N_28725);
nor U29084 (N_29084,N_28589,N_28634);
and U29085 (N_29085,N_28952,N_28608);
or U29086 (N_29086,N_28752,N_28555);
nor U29087 (N_29087,N_28945,N_28772);
nor U29088 (N_29088,N_28936,N_28734);
and U29089 (N_29089,N_28868,N_28985);
nor U29090 (N_29090,N_28569,N_28875);
and U29091 (N_29091,N_28614,N_28809);
nand U29092 (N_29092,N_28631,N_28523);
and U29093 (N_29093,N_28923,N_28894);
nand U29094 (N_29094,N_28870,N_28630);
nor U29095 (N_29095,N_28877,N_28500);
and U29096 (N_29096,N_28869,N_28615);
xnor U29097 (N_29097,N_28627,N_28599);
and U29098 (N_29098,N_28503,N_28963);
nand U29099 (N_29099,N_28983,N_28613);
nor U29100 (N_29100,N_28974,N_28931);
nor U29101 (N_29101,N_28986,N_28926);
or U29102 (N_29102,N_28779,N_28525);
or U29103 (N_29103,N_28656,N_28933);
and U29104 (N_29104,N_28519,N_28616);
or U29105 (N_29105,N_28529,N_28588);
nand U29106 (N_29106,N_28977,N_28520);
or U29107 (N_29107,N_28612,N_28584);
nand U29108 (N_29108,N_28987,N_28737);
xnor U29109 (N_29109,N_28846,N_28543);
and U29110 (N_29110,N_28824,N_28531);
and U29111 (N_29111,N_28665,N_28958);
xor U29112 (N_29112,N_28777,N_28996);
xnor U29113 (N_29113,N_28742,N_28644);
nor U29114 (N_29114,N_28577,N_28946);
or U29115 (N_29115,N_28748,N_28722);
and U29116 (N_29116,N_28579,N_28785);
xnor U29117 (N_29117,N_28704,N_28853);
xnor U29118 (N_29118,N_28719,N_28990);
or U29119 (N_29119,N_28566,N_28565);
xor U29120 (N_29120,N_28833,N_28960);
xor U29121 (N_29121,N_28643,N_28550);
and U29122 (N_29122,N_28991,N_28549);
or U29123 (N_29123,N_28812,N_28626);
and U29124 (N_29124,N_28667,N_28810);
and U29125 (N_29125,N_28746,N_28912);
nor U29126 (N_29126,N_28883,N_28964);
nand U29127 (N_29127,N_28844,N_28670);
xor U29128 (N_29128,N_28789,N_28611);
nand U29129 (N_29129,N_28647,N_28822);
nor U29130 (N_29130,N_28796,N_28661);
xnor U29131 (N_29131,N_28541,N_28586);
xor U29132 (N_29132,N_28658,N_28653);
nor U29133 (N_29133,N_28563,N_28580);
nand U29134 (N_29134,N_28811,N_28835);
nand U29135 (N_29135,N_28865,N_28807);
and U29136 (N_29136,N_28864,N_28827);
or U29137 (N_29137,N_28838,N_28764);
nand U29138 (N_29138,N_28623,N_28639);
nand U29139 (N_29139,N_28605,N_28692);
and U29140 (N_29140,N_28966,N_28617);
or U29141 (N_29141,N_28730,N_28801);
nor U29142 (N_29142,N_28562,N_28557);
nand U29143 (N_29143,N_28532,N_28687);
nor U29144 (N_29144,N_28542,N_28907);
nand U29145 (N_29145,N_28750,N_28874);
nor U29146 (N_29146,N_28583,N_28578);
nor U29147 (N_29147,N_28598,N_28671);
and U29148 (N_29148,N_28657,N_28739);
nand U29149 (N_29149,N_28928,N_28922);
or U29150 (N_29150,N_28951,N_28937);
nor U29151 (N_29151,N_28965,N_28860);
and U29152 (N_29152,N_28548,N_28518);
xor U29153 (N_29153,N_28956,N_28705);
xnor U29154 (N_29154,N_28655,N_28871);
nor U29155 (N_29155,N_28862,N_28511);
and U29156 (N_29156,N_28798,N_28904);
nor U29157 (N_29157,N_28663,N_28762);
or U29158 (N_29158,N_28940,N_28736);
and U29159 (N_29159,N_28887,N_28637);
xnor U29160 (N_29160,N_28673,N_28539);
and U29161 (N_29161,N_28547,N_28679);
nor U29162 (N_29162,N_28911,N_28891);
nand U29163 (N_29163,N_28898,N_28699);
nor U29164 (N_29164,N_28516,N_28995);
or U29165 (N_29165,N_28620,N_28980);
nand U29166 (N_29166,N_28757,N_28808);
or U29167 (N_29167,N_28765,N_28708);
nand U29168 (N_29168,N_28618,N_28732);
nand U29169 (N_29169,N_28896,N_28680);
xor U29170 (N_29170,N_28758,N_28527);
nand U29171 (N_29171,N_28747,N_28755);
and U29172 (N_29172,N_28650,N_28784);
xor U29173 (N_29173,N_28903,N_28888);
xor U29174 (N_29174,N_28815,N_28600);
nor U29175 (N_29175,N_28718,N_28852);
xnor U29176 (N_29176,N_28895,N_28855);
and U29177 (N_29177,N_28756,N_28575);
or U29178 (N_29178,N_28741,N_28955);
nor U29179 (N_29179,N_28802,N_28694);
nor U29180 (N_29180,N_28720,N_28766);
nand U29181 (N_29181,N_28662,N_28505);
or U29182 (N_29182,N_28900,N_28914);
and U29183 (N_29183,N_28753,N_28726);
nand U29184 (N_29184,N_28921,N_28745);
xnor U29185 (N_29185,N_28997,N_28502);
nor U29186 (N_29186,N_28994,N_28897);
xnor U29187 (N_29187,N_28843,N_28697);
and U29188 (N_29188,N_28524,N_28919);
nor U29189 (N_29189,N_28646,N_28932);
or U29190 (N_29190,N_28740,N_28711);
xor U29191 (N_29191,N_28947,N_28836);
nor U29192 (N_29192,N_28880,N_28691);
nor U29193 (N_29193,N_28976,N_28797);
and U29194 (N_29194,N_28854,N_28537);
or U29195 (N_29195,N_28585,N_28771);
and U29196 (N_29196,N_28669,N_28916);
nand U29197 (N_29197,N_28805,N_28909);
and U29198 (N_29198,N_28885,N_28666);
nor U29199 (N_29199,N_28939,N_28759);
and U29200 (N_29200,N_28782,N_28545);
xor U29201 (N_29201,N_28675,N_28512);
nand U29202 (N_29202,N_28992,N_28918);
or U29203 (N_29203,N_28712,N_28521);
nor U29204 (N_29204,N_28701,N_28595);
and U29205 (N_29205,N_28969,N_28559);
and U29206 (N_29206,N_28882,N_28628);
xor U29207 (N_29207,N_28954,N_28929);
xor U29208 (N_29208,N_28944,N_28793);
nand U29209 (N_29209,N_28774,N_28707);
nor U29210 (N_29210,N_28893,N_28892);
or U29211 (N_29211,N_28724,N_28884);
or U29212 (N_29212,N_28602,N_28915);
and U29213 (N_29213,N_28760,N_28506);
nand U29214 (N_29214,N_28702,N_28950);
nor U29215 (N_29215,N_28713,N_28845);
nor U29216 (N_29216,N_28553,N_28546);
nor U29217 (N_29217,N_28706,N_28574);
or U29218 (N_29218,N_28710,N_28509);
nor U29219 (N_29219,N_28821,N_28842);
xnor U29220 (N_29220,N_28695,N_28649);
xor U29221 (N_29221,N_28693,N_28554);
xnor U29222 (N_29222,N_28781,N_28596);
or U29223 (N_29223,N_28558,N_28840);
and U29224 (N_29224,N_28544,N_28526);
nand U29225 (N_29225,N_28913,N_28773);
and U29226 (N_29226,N_28568,N_28738);
nand U29227 (N_29227,N_28761,N_28820);
xnor U29228 (N_29228,N_28556,N_28678);
nand U29229 (N_29229,N_28850,N_28672);
nor U29230 (N_29230,N_28681,N_28953);
nor U29231 (N_29231,N_28993,N_28957);
xnor U29232 (N_29232,N_28902,N_28890);
nor U29233 (N_29233,N_28849,N_28508);
or U29234 (N_29234,N_28806,N_28823);
xnor U29235 (N_29235,N_28839,N_28858);
nor U29236 (N_29236,N_28786,N_28847);
nor U29237 (N_29237,N_28775,N_28791);
nor U29238 (N_29238,N_28716,N_28540);
xor U29239 (N_29239,N_28828,N_28538);
and U29240 (N_29240,N_28507,N_28685);
and U29241 (N_29241,N_28878,N_28829);
or U29242 (N_29242,N_28826,N_28729);
and U29243 (N_29243,N_28510,N_28515);
or U29244 (N_29244,N_28731,N_28660);
or U29245 (N_29245,N_28684,N_28633);
or U29246 (N_29246,N_28682,N_28576);
xor U29247 (N_29247,N_28886,N_28591);
or U29248 (N_29248,N_28834,N_28625);
nand U29249 (N_29249,N_28648,N_28601);
nor U29250 (N_29250,N_28984,N_28887);
xor U29251 (N_29251,N_28685,N_28852);
xor U29252 (N_29252,N_28669,N_28610);
nor U29253 (N_29253,N_28803,N_28841);
and U29254 (N_29254,N_28857,N_28926);
and U29255 (N_29255,N_28565,N_28946);
and U29256 (N_29256,N_28569,N_28728);
nor U29257 (N_29257,N_28530,N_28604);
or U29258 (N_29258,N_28718,N_28710);
and U29259 (N_29259,N_28780,N_28826);
nor U29260 (N_29260,N_28827,N_28500);
and U29261 (N_29261,N_28662,N_28868);
or U29262 (N_29262,N_28769,N_28784);
nor U29263 (N_29263,N_28693,N_28815);
and U29264 (N_29264,N_28758,N_28845);
and U29265 (N_29265,N_28768,N_28554);
and U29266 (N_29266,N_28782,N_28682);
xnor U29267 (N_29267,N_28764,N_28955);
nor U29268 (N_29268,N_28730,N_28709);
or U29269 (N_29269,N_28632,N_28849);
xnor U29270 (N_29270,N_28668,N_28885);
xor U29271 (N_29271,N_28826,N_28984);
nor U29272 (N_29272,N_28830,N_28510);
xnor U29273 (N_29273,N_28622,N_28667);
nand U29274 (N_29274,N_28740,N_28937);
nor U29275 (N_29275,N_28865,N_28830);
xor U29276 (N_29276,N_28635,N_28569);
xnor U29277 (N_29277,N_28507,N_28869);
nor U29278 (N_29278,N_28500,N_28934);
or U29279 (N_29279,N_28808,N_28735);
nor U29280 (N_29280,N_28881,N_28975);
or U29281 (N_29281,N_28764,N_28826);
nand U29282 (N_29282,N_28822,N_28940);
nand U29283 (N_29283,N_28645,N_28729);
nand U29284 (N_29284,N_28761,N_28603);
and U29285 (N_29285,N_28863,N_28897);
or U29286 (N_29286,N_28814,N_28920);
xor U29287 (N_29287,N_28855,N_28568);
nand U29288 (N_29288,N_28662,N_28679);
or U29289 (N_29289,N_28534,N_28544);
nand U29290 (N_29290,N_28950,N_28928);
nand U29291 (N_29291,N_28717,N_28652);
or U29292 (N_29292,N_28791,N_28649);
and U29293 (N_29293,N_28977,N_28673);
xnor U29294 (N_29294,N_28610,N_28670);
nor U29295 (N_29295,N_28889,N_28613);
xor U29296 (N_29296,N_28742,N_28896);
or U29297 (N_29297,N_28809,N_28913);
and U29298 (N_29298,N_28512,N_28651);
or U29299 (N_29299,N_28691,N_28907);
nor U29300 (N_29300,N_28676,N_28641);
xnor U29301 (N_29301,N_28950,N_28667);
nand U29302 (N_29302,N_28687,N_28674);
nor U29303 (N_29303,N_28927,N_28615);
xor U29304 (N_29304,N_28776,N_28921);
nand U29305 (N_29305,N_28660,N_28502);
xor U29306 (N_29306,N_28979,N_28763);
or U29307 (N_29307,N_28601,N_28991);
and U29308 (N_29308,N_28685,N_28698);
nand U29309 (N_29309,N_28593,N_28841);
nand U29310 (N_29310,N_28527,N_28738);
and U29311 (N_29311,N_28806,N_28888);
xnor U29312 (N_29312,N_28562,N_28609);
nand U29313 (N_29313,N_28504,N_28937);
nand U29314 (N_29314,N_28595,N_28936);
xor U29315 (N_29315,N_28668,N_28638);
nor U29316 (N_29316,N_28716,N_28794);
or U29317 (N_29317,N_28920,N_28616);
or U29318 (N_29318,N_28614,N_28851);
and U29319 (N_29319,N_28957,N_28544);
or U29320 (N_29320,N_28649,N_28823);
nor U29321 (N_29321,N_28848,N_28841);
and U29322 (N_29322,N_28863,N_28889);
nor U29323 (N_29323,N_28995,N_28599);
xor U29324 (N_29324,N_28858,N_28994);
nand U29325 (N_29325,N_28618,N_28624);
and U29326 (N_29326,N_28781,N_28779);
xnor U29327 (N_29327,N_28639,N_28642);
xor U29328 (N_29328,N_28904,N_28599);
and U29329 (N_29329,N_28533,N_28758);
and U29330 (N_29330,N_28518,N_28712);
and U29331 (N_29331,N_28710,N_28884);
or U29332 (N_29332,N_28825,N_28569);
or U29333 (N_29333,N_28620,N_28916);
xnor U29334 (N_29334,N_28647,N_28725);
nor U29335 (N_29335,N_28596,N_28581);
or U29336 (N_29336,N_28708,N_28697);
and U29337 (N_29337,N_28662,N_28725);
xnor U29338 (N_29338,N_28698,N_28504);
xor U29339 (N_29339,N_28949,N_28819);
or U29340 (N_29340,N_28831,N_28567);
and U29341 (N_29341,N_28879,N_28749);
nor U29342 (N_29342,N_28547,N_28688);
and U29343 (N_29343,N_28545,N_28562);
xnor U29344 (N_29344,N_28728,N_28733);
or U29345 (N_29345,N_28502,N_28897);
or U29346 (N_29346,N_28934,N_28554);
xor U29347 (N_29347,N_28604,N_28517);
nand U29348 (N_29348,N_28838,N_28980);
nand U29349 (N_29349,N_28704,N_28549);
nor U29350 (N_29350,N_28613,N_28691);
or U29351 (N_29351,N_28505,N_28639);
xnor U29352 (N_29352,N_28697,N_28590);
or U29353 (N_29353,N_28693,N_28796);
and U29354 (N_29354,N_28917,N_28668);
and U29355 (N_29355,N_28536,N_28547);
or U29356 (N_29356,N_28547,N_28968);
and U29357 (N_29357,N_28924,N_28645);
nand U29358 (N_29358,N_28720,N_28675);
nor U29359 (N_29359,N_28694,N_28885);
or U29360 (N_29360,N_28781,N_28526);
and U29361 (N_29361,N_28943,N_28607);
or U29362 (N_29362,N_28794,N_28819);
xnor U29363 (N_29363,N_28835,N_28680);
nand U29364 (N_29364,N_28649,N_28537);
and U29365 (N_29365,N_28531,N_28573);
nor U29366 (N_29366,N_28801,N_28704);
nand U29367 (N_29367,N_28611,N_28646);
nor U29368 (N_29368,N_28588,N_28955);
nor U29369 (N_29369,N_28704,N_28795);
nor U29370 (N_29370,N_28596,N_28875);
xnor U29371 (N_29371,N_28764,N_28952);
nand U29372 (N_29372,N_28940,N_28911);
xnor U29373 (N_29373,N_28965,N_28700);
or U29374 (N_29374,N_28773,N_28933);
xnor U29375 (N_29375,N_28718,N_28886);
xor U29376 (N_29376,N_28889,N_28977);
and U29377 (N_29377,N_28674,N_28536);
xor U29378 (N_29378,N_28807,N_28515);
nor U29379 (N_29379,N_28961,N_28833);
nand U29380 (N_29380,N_28632,N_28959);
or U29381 (N_29381,N_28790,N_28702);
nor U29382 (N_29382,N_28541,N_28897);
nand U29383 (N_29383,N_28580,N_28633);
nor U29384 (N_29384,N_28865,N_28855);
nand U29385 (N_29385,N_28907,N_28884);
nor U29386 (N_29386,N_28651,N_28650);
xor U29387 (N_29387,N_28666,N_28578);
nor U29388 (N_29388,N_28808,N_28925);
nor U29389 (N_29389,N_28637,N_28963);
or U29390 (N_29390,N_28814,N_28690);
nor U29391 (N_29391,N_28816,N_28593);
xor U29392 (N_29392,N_28720,N_28737);
nand U29393 (N_29393,N_28602,N_28629);
nand U29394 (N_29394,N_28985,N_28613);
nor U29395 (N_29395,N_28812,N_28775);
and U29396 (N_29396,N_28839,N_28561);
nand U29397 (N_29397,N_28898,N_28819);
xnor U29398 (N_29398,N_28846,N_28845);
nand U29399 (N_29399,N_28777,N_28524);
nor U29400 (N_29400,N_28954,N_28594);
xnor U29401 (N_29401,N_28836,N_28846);
xor U29402 (N_29402,N_28841,N_28821);
nor U29403 (N_29403,N_28886,N_28874);
and U29404 (N_29404,N_28903,N_28841);
xor U29405 (N_29405,N_28867,N_28846);
and U29406 (N_29406,N_28892,N_28575);
and U29407 (N_29407,N_28800,N_28660);
nand U29408 (N_29408,N_28633,N_28504);
nand U29409 (N_29409,N_28965,N_28659);
nor U29410 (N_29410,N_28588,N_28647);
nor U29411 (N_29411,N_28920,N_28740);
nor U29412 (N_29412,N_28935,N_28639);
and U29413 (N_29413,N_28554,N_28929);
xor U29414 (N_29414,N_28900,N_28570);
xnor U29415 (N_29415,N_28775,N_28703);
nand U29416 (N_29416,N_28810,N_28602);
and U29417 (N_29417,N_28839,N_28711);
xnor U29418 (N_29418,N_28969,N_28847);
nand U29419 (N_29419,N_28568,N_28892);
or U29420 (N_29420,N_28761,N_28849);
xnor U29421 (N_29421,N_28800,N_28571);
or U29422 (N_29422,N_28599,N_28680);
xor U29423 (N_29423,N_28829,N_28635);
nand U29424 (N_29424,N_28599,N_28869);
xor U29425 (N_29425,N_28987,N_28907);
nor U29426 (N_29426,N_28865,N_28887);
or U29427 (N_29427,N_28817,N_28811);
and U29428 (N_29428,N_28617,N_28582);
nand U29429 (N_29429,N_28504,N_28561);
nand U29430 (N_29430,N_28638,N_28718);
xor U29431 (N_29431,N_28752,N_28704);
and U29432 (N_29432,N_28679,N_28503);
xnor U29433 (N_29433,N_28781,N_28620);
nor U29434 (N_29434,N_28593,N_28564);
and U29435 (N_29435,N_28641,N_28577);
xor U29436 (N_29436,N_28792,N_28951);
and U29437 (N_29437,N_28974,N_28642);
and U29438 (N_29438,N_28678,N_28582);
nand U29439 (N_29439,N_28813,N_28946);
nor U29440 (N_29440,N_28833,N_28511);
nor U29441 (N_29441,N_28568,N_28930);
nor U29442 (N_29442,N_28659,N_28682);
nor U29443 (N_29443,N_28608,N_28841);
nor U29444 (N_29444,N_28581,N_28890);
or U29445 (N_29445,N_28507,N_28973);
and U29446 (N_29446,N_28631,N_28914);
and U29447 (N_29447,N_28870,N_28583);
and U29448 (N_29448,N_28908,N_28622);
xor U29449 (N_29449,N_28779,N_28874);
or U29450 (N_29450,N_28513,N_28613);
nand U29451 (N_29451,N_28903,N_28914);
or U29452 (N_29452,N_28729,N_28599);
or U29453 (N_29453,N_28973,N_28728);
nand U29454 (N_29454,N_28648,N_28894);
nand U29455 (N_29455,N_28821,N_28791);
nand U29456 (N_29456,N_28945,N_28691);
and U29457 (N_29457,N_28934,N_28647);
xnor U29458 (N_29458,N_28976,N_28659);
or U29459 (N_29459,N_28960,N_28548);
and U29460 (N_29460,N_28519,N_28986);
nand U29461 (N_29461,N_28554,N_28980);
and U29462 (N_29462,N_28523,N_28894);
nand U29463 (N_29463,N_28510,N_28724);
or U29464 (N_29464,N_28759,N_28897);
nor U29465 (N_29465,N_28822,N_28592);
nand U29466 (N_29466,N_28646,N_28858);
and U29467 (N_29467,N_28573,N_28551);
nor U29468 (N_29468,N_28900,N_28812);
and U29469 (N_29469,N_28759,N_28541);
nand U29470 (N_29470,N_28898,N_28838);
nor U29471 (N_29471,N_28867,N_28843);
nand U29472 (N_29472,N_28610,N_28558);
or U29473 (N_29473,N_28676,N_28824);
nand U29474 (N_29474,N_28793,N_28991);
nor U29475 (N_29475,N_28515,N_28803);
nand U29476 (N_29476,N_28809,N_28747);
nand U29477 (N_29477,N_28909,N_28809);
nand U29478 (N_29478,N_28619,N_28789);
nor U29479 (N_29479,N_28831,N_28602);
or U29480 (N_29480,N_28535,N_28986);
and U29481 (N_29481,N_28955,N_28839);
xor U29482 (N_29482,N_28685,N_28642);
and U29483 (N_29483,N_28896,N_28826);
and U29484 (N_29484,N_28534,N_28987);
or U29485 (N_29485,N_28907,N_28974);
nor U29486 (N_29486,N_28573,N_28878);
and U29487 (N_29487,N_28992,N_28646);
nor U29488 (N_29488,N_28957,N_28689);
nor U29489 (N_29489,N_28635,N_28509);
nor U29490 (N_29490,N_28859,N_28727);
or U29491 (N_29491,N_28504,N_28978);
or U29492 (N_29492,N_28739,N_28724);
nor U29493 (N_29493,N_28982,N_28680);
and U29494 (N_29494,N_28935,N_28542);
or U29495 (N_29495,N_28620,N_28521);
xor U29496 (N_29496,N_28646,N_28994);
xor U29497 (N_29497,N_28579,N_28756);
and U29498 (N_29498,N_28638,N_28573);
nor U29499 (N_29499,N_28784,N_28698);
nand U29500 (N_29500,N_29088,N_29388);
xnor U29501 (N_29501,N_29331,N_29314);
nand U29502 (N_29502,N_29470,N_29361);
nand U29503 (N_29503,N_29087,N_29397);
and U29504 (N_29504,N_29146,N_29144);
and U29505 (N_29505,N_29080,N_29190);
and U29506 (N_29506,N_29234,N_29276);
xnor U29507 (N_29507,N_29124,N_29206);
or U29508 (N_29508,N_29041,N_29297);
or U29509 (N_29509,N_29201,N_29373);
xnor U29510 (N_29510,N_29465,N_29005);
or U29511 (N_29511,N_29494,N_29447);
xor U29512 (N_29512,N_29018,N_29192);
or U29513 (N_29513,N_29301,N_29377);
and U29514 (N_29514,N_29093,N_29236);
nor U29515 (N_29515,N_29467,N_29347);
and U29516 (N_29516,N_29395,N_29405);
xnor U29517 (N_29517,N_29267,N_29382);
xor U29518 (N_29518,N_29360,N_29111);
nand U29519 (N_29519,N_29460,N_29158);
or U29520 (N_29520,N_29300,N_29261);
nand U29521 (N_29521,N_29274,N_29439);
and U29522 (N_29522,N_29351,N_29463);
nor U29523 (N_29523,N_29108,N_29004);
and U29524 (N_29524,N_29283,N_29168);
nor U29525 (N_29525,N_29161,N_29040);
xor U29526 (N_29526,N_29119,N_29231);
xnor U29527 (N_29527,N_29256,N_29086);
nand U29528 (N_29528,N_29091,N_29246);
nor U29529 (N_29529,N_29245,N_29065);
nand U29530 (N_29530,N_29468,N_29047);
nor U29531 (N_29531,N_29042,N_29226);
nand U29532 (N_29532,N_29436,N_29238);
or U29533 (N_29533,N_29356,N_29324);
and U29534 (N_29534,N_29056,N_29384);
xnor U29535 (N_29535,N_29400,N_29071);
nand U29536 (N_29536,N_29413,N_29118);
xnor U29537 (N_29537,N_29346,N_29403);
nor U29538 (N_29538,N_29315,N_29044);
xnor U29539 (N_29539,N_29126,N_29099);
nand U29540 (N_29540,N_29480,N_29054);
or U29541 (N_29541,N_29123,N_29140);
xnor U29542 (N_29542,N_29440,N_29374);
nor U29543 (N_29543,N_29489,N_29112);
and U29544 (N_29544,N_29273,N_29375);
xor U29545 (N_29545,N_29433,N_29461);
nor U29546 (N_29546,N_29213,N_29335);
nand U29547 (N_29547,N_29391,N_29365);
xnor U29548 (N_29548,N_29372,N_29390);
and U29549 (N_29549,N_29370,N_29142);
nand U29550 (N_29550,N_29265,N_29302);
nand U29551 (N_29551,N_29223,N_29442);
and U29552 (N_29552,N_29452,N_29036);
or U29553 (N_29553,N_29176,N_29287);
nor U29554 (N_29554,N_29415,N_29114);
or U29555 (N_29555,N_29007,N_29279);
and U29556 (N_29556,N_29116,N_29425);
and U29557 (N_29557,N_29414,N_29420);
nor U29558 (N_29558,N_29232,N_29340);
nand U29559 (N_29559,N_29253,N_29145);
nand U29560 (N_29560,N_29032,N_29345);
nor U29561 (N_29561,N_29185,N_29457);
or U29562 (N_29562,N_29311,N_29416);
and U29563 (N_29563,N_29288,N_29318);
nand U29564 (N_29564,N_29089,N_29187);
or U29565 (N_29565,N_29157,N_29476);
nor U29566 (N_29566,N_29182,N_29312);
and U29567 (N_29567,N_29410,N_29320);
nand U29568 (N_29568,N_29241,N_29083);
nand U29569 (N_29569,N_29205,N_29497);
and U29570 (N_29570,N_29230,N_29202);
and U29571 (N_29571,N_29034,N_29474);
nor U29572 (N_29572,N_29159,N_29125);
xnor U29573 (N_29573,N_29155,N_29254);
xor U29574 (N_29574,N_29115,N_29191);
and U29575 (N_29575,N_29020,N_29131);
xor U29576 (N_29576,N_29475,N_29334);
or U29577 (N_29577,N_29399,N_29063);
nand U29578 (N_29578,N_29010,N_29045);
nor U29579 (N_29579,N_29015,N_29257);
or U29580 (N_29580,N_29035,N_29250);
or U29581 (N_29581,N_29082,N_29174);
nor U29582 (N_29582,N_29444,N_29477);
nand U29583 (N_29583,N_29291,N_29290);
nand U29584 (N_29584,N_29298,N_29396);
nand U29585 (N_29585,N_29195,N_29059);
nand U29586 (N_29586,N_29104,N_29184);
and U29587 (N_29587,N_29423,N_29098);
nor U29588 (N_29588,N_29130,N_29012);
nand U29589 (N_29589,N_29451,N_29198);
nand U29590 (N_29590,N_29242,N_29352);
xnor U29591 (N_29591,N_29379,N_29408);
and U29592 (N_29592,N_29404,N_29364);
and U29593 (N_29593,N_29357,N_29081);
nor U29594 (N_29594,N_29342,N_29211);
and U29595 (N_29595,N_29027,N_29271);
nand U29596 (N_29596,N_29469,N_29259);
nor U29597 (N_29597,N_29350,N_29322);
or U29598 (N_29598,N_29438,N_29449);
nor U29599 (N_29599,N_29492,N_29165);
and U29600 (N_29600,N_29147,N_29325);
xor U29601 (N_29601,N_29432,N_29359);
and U29602 (N_29602,N_29085,N_29493);
nand U29603 (N_29603,N_29478,N_29269);
xnor U29604 (N_29604,N_29150,N_29128);
or U29605 (N_29605,N_29178,N_29249);
nor U29606 (N_29606,N_29096,N_29075);
xnor U29607 (N_29607,N_29456,N_29337);
nor U29608 (N_29608,N_29272,N_29479);
xnor U29609 (N_29609,N_29049,N_29260);
nor U29610 (N_29610,N_29304,N_29417);
xnor U29611 (N_29611,N_29367,N_29109);
or U29612 (N_29612,N_29022,N_29220);
or U29613 (N_29613,N_29455,N_29316);
xor U29614 (N_29614,N_29207,N_29028);
xor U29615 (N_29615,N_29485,N_29310);
xnor U29616 (N_29616,N_29381,N_29362);
xnor U29617 (N_29617,N_29107,N_29426);
or U29618 (N_29618,N_29393,N_29030);
or U29619 (N_29619,N_29333,N_29499);
nand U29620 (N_29620,N_29329,N_29151);
and U29621 (N_29621,N_29053,N_29336);
and U29622 (N_29622,N_29358,N_29039);
and U29623 (N_29623,N_29102,N_29348);
xor U29624 (N_29624,N_29180,N_29203);
nor U29625 (N_29625,N_29077,N_29305);
and U29626 (N_29626,N_29349,N_29422);
or U29627 (N_29627,N_29255,N_29453);
nand U29628 (N_29628,N_29094,N_29406);
and U29629 (N_29629,N_29369,N_29058);
nand U29630 (N_29630,N_29219,N_29371);
nor U29631 (N_29631,N_29378,N_29106);
nor U29632 (N_29632,N_29275,N_29401);
nor U29633 (N_29633,N_29014,N_29355);
nand U29634 (N_29634,N_29189,N_29194);
xnor U29635 (N_29635,N_29498,N_29224);
or U29636 (N_29636,N_29023,N_29445);
nand U29637 (N_29637,N_29363,N_29026);
or U29638 (N_29638,N_29200,N_29076);
or U29639 (N_29639,N_29166,N_29172);
nand U29640 (N_29640,N_29171,N_29286);
and U29641 (N_29641,N_29216,N_29306);
nand U29642 (N_29642,N_29001,N_29120);
and U29643 (N_29643,N_29321,N_29454);
and U29644 (N_29644,N_29092,N_29137);
nor U29645 (N_29645,N_29326,N_29285);
and U29646 (N_29646,N_29354,N_29046);
xnor U29647 (N_29647,N_29199,N_29067);
and U29648 (N_29648,N_29308,N_29394);
xor U29649 (N_29649,N_29330,N_29487);
nand U29650 (N_29650,N_29295,N_29409);
or U29651 (N_29651,N_29490,N_29013);
xnor U29652 (N_29652,N_29252,N_29196);
and U29653 (N_29653,N_29138,N_29133);
nand U29654 (N_29654,N_29025,N_29280);
nor U29655 (N_29655,N_29069,N_29074);
xor U29656 (N_29656,N_29011,N_29412);
or U29657 (N_29657,N_29338,N_29443);
or U29658 (N_29658,N_29418,N_29353);
xnor U29659 (N_29659,N_29495,N_29227);
and U29660 (N_29660,N_29188,N_29385);
or U29661 (N_29661,N_29411,N_29132);
xor U29662 (N_29662,N_29033,N_29141);
nand U29663 (N_29663,N_29428,N_29429);
and U29664 (N_29664,N_29263,N_29343);
nor U29665 (N_29665,N_29268,N_29068);
and U29666 (N_29666,N_29421,N_29292);
nand U29667 (N_29667,N_29204,N_29072);
and U29668 (N_29668,N_29486,N_29278);
xnor U29669 (N_29669,N_29079,N_29127);
or U29670 (N_29670,N_29215,N_29459);
or U29671 (N_29671,N_29113,N_29167);
and U29672 (N_29672,N_29031,N_29100);
or U29673 (N_29673,N_29491,N_29193);
or U29674 (N_29674,N_29217,N_29024);
or U29675 (N_29675,N_29446,N_29294);
xnor U29676 (N_29676,N_29152,N_29386);
or U29677 (N_29677,N_29328,N_29052);
nand U29678 (N_29678,N_29368,N_29472);
and U29679 (N_29679,N_29170,N_29208);
nand U29680 (N_29680,N_29062,N_29117);
xor U29681 (N_29681,N_29389,N_29248);
nor U29682 (N_29682,N_29148,N_29175);
nor U29683 (N_29683,N_29037,N_29209);
or U29684 (N_29684,N_29073,N_29222);
nor U29685 (N_29685,N_29319,N_29139);
xor U29686 (N_29686,N_29303,N_29048);
xor U29687 (N_29687,N_29437,N_29392);
or U29688 (N_29688,N_29462,N_29299);
xor U29689 (N_29689,N_29229,N_29380);
and U29690 (N_29690,N_29339,N_29435);
nand U29691 (N_29691,N_29473,N_29021);
or U29692 (N_29692,N_29317,N_29247);
nand U29693 (N_29693,N_29235,N_29376);
nor U29694 (N_29694,N_29050,N_29450);
xnor U29695 (N_29695,N_29481,N_29055);
xor U29696 (N_29696,N_29323,N_29090);
and U29697 (N_29697,N_29136,N_29095);
nor U29698 (N_29698,N_29434,N_29262);
nand U29699 (N_29699,N_29129,N_29218);
xor U29700 (N_29700,N_29233,N_29424);
nor U29701 (N_29701,N_29164,N_29344);
or U29702 (N_29702,N_29496,N_29122);
nand U29703 (N_29703,N_29270,N_29110);
nor U29704 (N_29704,N_29264,N_29017);
xnor U29705 (N_29705,N_29078,N_29289);
and U29706 (N_29706,N_29327,N_29097);
nand U29707 (N_29707,N_29006,N_29019);
nor U29708 (N_29708,N_29135,N_29186);
nor U29709 (N_29709,N_29134,N_29070);
and U29710 (N_29710,N_29313,N_29366);
nor U29711 (N_29711,N_29441,N_29103);
or U29712 (N_29712,N_29427,N_29064);
nand U29713 (N_29713,N_29458,N_29228);
xnor U29714 (N_29714,N_29009,N_29029);
nand U29715 (N_29715,N_29177,N_29179);
xnor U29716 (N_29716,N_29149,N_29471);
nor U29717 (N_29717,N_29307,N_29183);
nor U29718 (N_29718,N_29084,N_29282);
or U29719 (N_29719,N_29284,N_29221);
and U29720 (N_29720,N_29482,N_29060);
nand U29721 (N_29721,N_29402,N_29483);
xor U29722 (N_29722,N_29464,N_29156);
xor U29723 (N_29723,N_29153,N_29243);
nor U29724 (N_29724,N_29066,N_29258);
nand U29725 (N_29725,N_29002,N_29383);
xnor U29726 (N_29726,N_29105,N_29225);
or U29727 (N_29727,N_29387,N_29101);
nor U29728 (N_29728,N_29484,N_29173);
nor U29729 (N_29729,N_29162,N_29281);
or U29730 (N_29730,N_29277,N_29181);
and U29731 (N_29731,N_29212,N_29466);
nand U29732 (N_29732,N_29296,N_29121);
nor U29733 (N_29733,N_29309,N_29239);
and U29734 (N_29734,N_29431,N_29003);
xor U29735 (N_29735,N_29154,N_29051);
xnor U29736 (N_29736,N_29143,N_29043);
nor U29737 (N_29737,N_29000,N_29240);
xnor U29738 (N_29738,N_29214,N_29341);
nand U29739 (N_29739,N_29169,N_29160);
and U29740 (N_29740,N_29016,N_29244);
and U29741 (N_29741,N_29057,N_29210);
nor U29742 (N_29742,N_29163,N_29266);
nor U29743 (N_29743,N_29008,N_29448);
or U29744 (N_29744,N_29419,N_29430);
and U29745 (N_29745,N_29407,N_29293);
and U29746 (N_29746,N_29061,N_29038);
and U29747 (N_29747,N_29398,N_29332);
nor U29748 (N_29748,N_29197,N_29488);
or U29749 (N_29749,N_29251,N_29237);
nor U29750 (N_29750,N_29430,N_29209);
nor U29751 (N_29751,N_29023,N_29398);
or U29752 (N_29752,N_29204,N_29355);
and U29753 (N_29753,N_29171,N_29334);
xor U29754 (N_29754,N_29360,N_29248);
nor U29755 (N_29755,N_29233,N_29314);
or U29756 (N_29756,N_29043,N_29012);
xnor U29757 (N_29757,N_29377,N_29275);
xor U29758 (N_29758,N_29099,N_29054);
xor U29759 (N_29759,N_29417,N_29425);
xnor U29760 (N_29760,N_29315,N_29105);
and U29761 (N_29761,N_29130,N_29150);
and U29762 (N_29762,N_29408,N_29436);
xnor U29763 (N_29763,N_29323,N_29235);
and U29764 (N_29764,N_29315,N_29203);
nor U29765 (N_29765,N_29330,N_29205);
or U29766 (N_29766,N_29488,N_29473);
nor U29767 (N_29767,N_29414,N_29496);
nor U29768 (N_29768,N_29045,N_29028);
nand U29769 (N_29769,N_29499,N_29272);
and U29770 (N_29770,N_29331,N_29266);
and U29771 (N_29771,N_29348,N_29406);
nor U29772 (N_29772,N_29207,N_29379);
nor U29773 (N_29773,N_29406,N_29463);
nor U29774 (N_29774,N_29441,N_29270);
xor U29775 (N_29775,N_29014,N_29476);
nand U29776 (N_29776,N_29124,N_29089);
or U29777 (N_29777,N_29338,N_29087);
xor U29778 (N_29778,N_29237,N_29286);
xnor U29779 (N_29779,N_29097,N_29463);
nor U29780 (N_29780,N_29015,N_29077);
or U29781 (N_29781,N_29245,N_29047);
and U29782 (N_29782,N_29045,N_29005);
nor U29783 (N_29783,N_29138,N_29469);
xnor U29784 (N_29784,N_29234,N_29383);
nor U29785 (N_29785,N_29146,N_29317);
xor U29786 (N_29786,N_29357,N_29023);
nand U29787 (N_29787,N_29253,N_29355);
nand U29788 (N_29788,N_29284,N_29347);
nor U29789 (N_29789,N_29450,N_29002);
nand U29790 (N_29790,N_29105,N_29201);
xnor U29791 (N_29791,N_29298,N_29165);
nand U29792 (N_29792,N_29223,N_29369);
nand U29793 (N_29793,N_29004,N_29482);
nand U29794 (N_29794,N_29328,N_29021);
and U29795 (N_29795,N_29288,N_29234);
or U29796 (N_29796,N_29277,N_29234);
nor U29797 (N_29797,N_29161,N_29237);
or U29798 (N_29798,N_29100,N_29385);
nor U29799 (N_29799,N_29180,N_29060);
nand U29800 (N_29800,N_29039,N_29129);
or U29801 (N_29801,N_29056,N_29253);
nand U29802 (N_29802,N_29029,N_29290);
xnor U29803 (N_29803,N_29186,N_29107);
or U29804 (N_29804,N_29493,N_29433);
xor U29805 (N_29805,N_29236,N_29177);
xor U29806 (N_29806,N_29312,N_29269);
xnor U29807 (N_29807,N_29483,N_29268);
nor U29808 (N_29808,N_29002,N_29201);
or U29809 (N_29809,N_29310,N_29096);
or U29810 (N_29810,N_29134,N_29006);
and U29811 (N_29811,N_29052,N_29267);
or U29812 (N_29812,N_29142,N_29390);
or U29813 (N_29813,N_29435,N_29136);
nand U29814 (N_29814,N_29174,N_29191);
or U29815 (N_29815,N_29168,N_29044);
or U29816 (N_29816,N_29119,N_29039);
xnor U29817 (N_29817,N_29313,N_29280);
or U29818 (N_29818,N_29447,N_29222);
nand U29819 (N_29819,N_29183,N_29401);
xor U29820 (N_29820,N_29247,N_29122);
and U29821 (N_29821,N_29493,N_29432);
nand U29822 (N_29822,N_29454,N_29277);
and U29823 (N_29823,N_29191,N_29077);
or U29824 (N_29824,N_29082,N_29107);
nor U29825 (N_29825,N_29138,N_29496);
nand U29826 (N_29826,N_29179,N_29297);
xnor U29827 (N_29827,N_29199,N_29053);
nor U29828 (N_29828,N_29250,N_29019);
nand U29829 (N_29829,N_29250,N_29234);
xnor U29830 (N_29830,N_29060,N_29179);
nand U29831 (N_29831,N_29219,N_29049);
nand U29832 (N_29832,N_29445,N_29311);
nor U29833 (N_29833,N_29263,N_29394);
and U29834 (N_29834,N_29389,N_29058);
xnor U29835 (N_29835,N_29046,N_29011);
nor U29836 (N_29836,N_29104,N_29407);
xor U29837 (N_29837,N_29414,N_29343);
nor U29838 (N_29838,N_29103,N_29242);
or U29839 (N_29839,N_29269,N_29294);
or U29840 (N_29840,N_29137,N_29485);
or U29841 (N_29841,N_29458,N_29113);
and U29842 (N_29842,N_29303,N_29461);
nand U29843 (N_29843,N_29135,N_29388);
and U29844 (N_29844,N_29447,N_29042);
nor U29845 (N_29845,N_29210,N_29000);
xor U29846 (N_29846,N_29290,N_29052);
nor U29847 (N_29847,N_29461,N_29362);
and U29848 (N_29848,N_29036,N_29380);
and U29849 (N_29849,N_29262,N_29197);
xnor U29850 (N_29850,N_29395,N_29375);
nor U29851 (N_29851,N_29359,N_29441);
nor U29852 (N_29852,N_29363,N_29017);
nand U29853 (N_29853,N_29282,N_29280);
and U29854 (N_29854,N_29402,N_29382);
or U29855 (N_29855,N_29156,N_29082);
nor U29856 (N_29856,N_29145,N_29112);
or U29857 (N_29857,N_29423,N_29402);
nand U29858 (N_29858,N_29365,N_29310);
nand U29859 (N_29859,N_29474,N_29144);
nor U29860 (N_29860,N_29119,N_29241);
nand U29861 (N_29861,N_29454,N_29343);
nor U29862 (N_29862,N_29286,N_29323);
nand U29863 (N_29863,N_29089,N_29043);
and U29864 (N_29864,N_29150,N_29010);
nor U29865 (N_29865,N_29047,N_29446);
and U29866 (N_29866,N_29001,N_29403);
nand U29867 (N_29867,N_29057,N_29075);
nand U29868 (N_29868,N_29061,N_29249);
or U29869 (N_29869,N_29055,N_29315);
and U29870 (N_29870,N_29488,N_29310);
xor U29871 (N_29871,N_29275,N_29404);
nand U29872 (N_29872,N_29059,N_29132);
and U29873 (N_29873,N_29498,N_29031);
and U29874 (N_29874,N_29317,N_29246);
nor U29875 (N_29875,N_29201,N_29235);
and U29876 (N_29876,N_29480,N_29381);
and U29877 (N_29877,N_29369,N_29422);
or U29878 (N_29878,N_29437,N_29140);
and U29879 (N_29879,N_29089,N_29383);
and U29880 (N_29880,N_29489,N_29428);
xnor U29881 (N_29881,N_29421,N_29149);
or U29882 (N_29882,N_29395,N_29482);
nand U29883 (N_29883,N_29178,N_29318);
and U29884 (N_29884,N_29372,N_29275);
or U29885 (N_29885,N_29427,N_29334);
or U29886 (N_29886,N_29470,N_29317);
and U29887 (N_29887,N_29308,N_29243);
or U29888 (N_29888,N_29192,N_29360);
or U29889 (N_29889,N_29145,N_29336);
xnor U29890 (N_29890,N_29087,N_29035);
and U29891 (N_29891,N_29225,N_29279);
nand U29892 (N_29892,N_29289,N_29486);
xor U29893 (N_29893,N_29370,N_29221);
and U29894 (N_29894,N_29428,N_29108);
nand U29895 (N_29895,N_29380,N_29087);
xor U29896 (N_29896,N_29263,N_29281);
nand U29897 (N_29897,N_29274,N_29244);
nand U29898 (N_29898,N_29304,N_29265);
xnor U29899 (N_29899,N_29022,N_29481);
nand U29900 (N_29900,N_29018,N_29084);
or U29901 (N_29901,N_29081,N_29372);
nor U29902 (N_29902,N_29264,N_29209);
nor U29903 (N_29903,N_29438,N_29018);
xnor U29904 (N_29904,N_29152,N_29342);
nor U29905 (N_29905,N_29120,N_29170);
or U29906 (N_29906,N_29015,N_29177);
nand U29907 (N_29907,N_29153,N_29313);
and U29908 (N_29908,N_29472,N_29437);
xor U29909 (N_29909,N_29461,N_29302);
or U29910 (N_29910,N_29352,N_29214);
nor U29911 (N_29911,N_29283,N_29305);
xor U29912 (N_29912,N_29048,N_29137);
nand U29913 (N_29913,N_29242,N_29055);
nand U29914 (N_29914,N_29141,N_29441);
nand U29915 (N_29915,N_29266,N_29385);
or U29916 (N_29916,N_29414,N_29429);
or U29917 (N_29917,N_29177,N_29228);
xor U29918 (N_29918,N_29417,N_29050);
nand U29919 (N_29919,N_29332,N_29038);
and U29920 (N_29920,N_29433,N_29275);
nand U29921 (N_29921,N_29147,N_29446);
nor U29922 (N_29922,N_29427,N_29250);
or U29923 (N_29923,N_29385,N_29355);
xnor U29924 (N_29924,N_29164,N_29016);
xor U29925 (N_29925,N_29188,N_29378);
or U29926 (N_29926,N_29227,N_29039);
nor U29927 (N_29927,N_29403,N_29232);
xnor U29928 (N_29928,N_29459,N_29234);
or U29929 (N_29929,N_29487,N_29461);
and U29930 (N_29930,N_29193,N_29452);
or U29931 (N_29931,N_29481,N_29452);
or U29932 (N_29932,N_29063,N_29402);
or U29933 (N_29933,N_29340,N_29198);
and U29934 (N_29934,N_29119,N_29065);
nor U29935 (N_29935,N_29360,N_29270);
and U29936 (N_29936,N_29087,N_29299);
xor U29937 (N_29937,N_29239,N_29066);
nor U29938 (N_29938,N_29317,N_29422);
nand U29939 (N_29939,N_29213,N_29112);
nor U29940 (N_29940,N_29131,N_29066);
or U29941 (N_29941,N_29088,N_29056);
xnor U29942 (N_29942,N_29168,N_29374);
or U29943 (N_29943,N_29265,N_29192);
or U29944 (N_29944,N_29330,N_29391);
xnor U29945 (N_29945,N_29404,N_29271);
xor U29946 (N_29946,N_29462,N_29304);
nand U29947 (N_29947,N_29318,N_29030);
or U29948 (N_29948,N_29094,N_29234);
xnor U29949 (N_29949,N_29035,N_29337);
nand U29950 (N_29950,N_29391,N_29064);
xor U29951 (N_29951,N_29371,N_29301);
nand U29952 (N_29952,N_29398,N_29331);
xor U29953 (N_29953,N_29348,N_29469);
xnor U29954 (N_29954,N_29273,N_29297);
xnor U29955 (N_29955,N_29406,N_29303);
and U29956 (N_29956,N_29162,N_29069);
nor U29957 (N_29957,N_29301,N_29473);
nand U29958 (N_29958,N_29314,N_29463);
and U29959 (N_29959,N_29075,N_29217);
nor U29960 (N_29960,N_29425,N_29334);
xor U29961 (N_29961,N_29387,N_29288);
nor U29962 (N_29962,N_29379,N_29310);
nor U29963 (N_29963,N_29032,N_29216);
xnor U29964 (N_29964,N_29239,N_29182);
and U29965 (N_29965,N_29362,N_29082);
nand U29966 (N_29966,N_29423,N_29293);
nor U29967 (N_29967,N_29172,N_29332);
xnor U29968 (N_29968,N_29095,N_29101);
and U29969 (N_29969,N_29116,N_29100);
or U29970 (N_29970,N_29033,N_29464);
xor U29971 (N_29971,N_29354,N_29264);
or U29972 (N_29972,N_29379,N_29158);
and U29973 (N_29973,N_29149,N_29355);
and U29974 (N_29974,N_29395,N_29181);
or U29975 (N_29975,N_29360,N_29359);
and U29976 (N_29976,N_29203,N_29160);
and U29977 (N_29977,N_29089,N_29049);
xor U29978 (N_29978,N_29406,N_29286);
and U29979 (N_29979,N_29417,N_29062);
or U29980 (N_29980,N_29345,N_29382);
and U29981 (N_29981,N_29026,N_29282);
or U29982 (N_29982,N_29060,N_29347);
or U29983 (N_29983,N_29205,N_29286);
and U29984 (N_29984,N_29199,N_29090);
xnor U29985 (N_29985,N_29048,N_29046);
or U29986 (N_29986,N_29007,N_29091);
nand U29987 (N_29987,N_29239,N_29107);
and U29988 (N_29988,N_29049,N_29246);
nand U29989 (N_29989,N_29499,N_29093);
and U29990 (N_29990,N_29331,N_29420);
nor U29991 (N_29991,N_29418,N_29451);
and U29992 (N_29992,N_29071,N_29263);
or U29993 (N_29993,N_29350,N_29116);
xor U29994 (N_29994,N_29224,N_29405);
and U29995 (N_29995,N_29197,N_29270);
nand U29996 (N_29996,N_29099,N_29355);
nand U29997 (N_29997,N_29289,N_29326);
nor U29998 (N_29998,N_29166,N_29263);
and U29999 (N_29999,N_29129,N_29485);
xnor U30000 (N_30000,N_29553,N_29936);
nor U30001 (N_30001,N_29649,N_29776);
and U30002 (N_30002,N_29904,N_29581);
and U30003 (N_30003,N_29505,N_29849);
nand U30004 (N_30004,N_29819,N_29755);
xnor U30005 (N_30005,N_29870,N_29863);
nand U30006 (N_30006,N_29631,N_29844);
and U30007 (N_30007,N_29998,N_29509);
nand U30008 (N_30008,N_29657,N_29661);
and U30009 (N_30009,N_29513,N_29851);
nor U30010 (N_30010,N_29674,N_29650);
xnor U30011 (N_30011,N_29628,N_29602);
nor U30012 (N_30012,N_29501,N_29635);
and U30013 (N_30013,N_29732,N_29880);
xor U30014 (N_30014,N_29556,N_29830);
nand U30015 (N_30015,N_29775,N_29921);
nor U30016 (N_30016,N_29905,N_29652);
xnor U30017 (N_30017,N_29687,N_29865);
xnor U30018 (N_30018,N_29818,N_29504);
nand U30019 (N_30019,N_29860,N_29566);
or U30020 (N_30020,N_29666,N_29537);
xnor U30021 (N_30021,N_29894,N_29976);
xnor U30022 (N_30022,N_29945,N_29757);
xor U30023 (N_30023,N_29788,N_29845);
nor U30024 (N_30024,N_29580,N_29774);
nand U30025 (N_30025,N_29989,N_29878);
nand U30026 (N_30026,N_29611,N_29591);
and U30027 (N_30027,N_29761,N_29705);
and U30028 (N_30028,N_29586,N_29767);
nor U30029 (N_30029,N_29503,N_29970);
nor U30030 (N_30030,N_29876,N_29911);
nand U30031 (N_30031,N_29886,N_29500);
xor U30032 (N_30032,N_29653,N_29744);
nand U30033 (N_30033,N_29733,N_29575);
nand U30034 (N_30034,N_29670,N_29809);
and U30035 (N_30035,N_29803,N_29632);
xor U30036 (N_30036,N_29655,N_29615);
and U30037 (N_30037,N_29869,N_29986);
nand U30038 (N_30038,N_29668,N_29742);
nand U30039 (N_30039,N_29510,N_29827);
nand U30040 (N_30040,N_29974,N_29559);
and U30041 (N_30041,N_29808,N_29939);
nor U30042 (N_30042,N_29579,N_29952);
and U30043 (N_30043,N_29917,N_29654);
nand U30044 (N_30044,N_29892,N_29571);
xor U30045 (N_30045,N_29965,N_29890);
nor U30046 (N_30046,N_29791,N_29638);
or U30047 (N_30047,N_29684,N_29531);
and U30048 (N_30048,N_29707,N_29660);
xnor U30049 (N_30049,N_29836,N_29561);
nor U30050 (N_30050,N_29528,N_29873);
nand U30051 (N_30051,N_29679,N_29919);
nor U30052 (N_30052,N_29837,N_29762);
nand U30053 (N_30053,N_29642,N_29949);
or U30054 (N_30054,N_29981,N_29884);
and U30055 (N_30055,N_29843,N_29942);
or U30056 (N_30056,N_29856,N_29754);
and U30057 (N_30057,N_29734,N_29585);
or U30058 (N_30058,N_29646,N_29685);
and U30059 (N_30059,N_29619,N_29539);
nor U30060 (N_30060,N_29736,N_29583);
nor U30061 (N_30061,N_29588,N_29549);
or U30062 (N_30062,N_29532,N_29621);
nor U30063 (N_30063,N_29534,N_29888);
and U30064 (N_30064,N_29766,N_29922);
xnor U30065 (N_30065,N_29798,N_29709);
and U30066 (N_30066,N_29868,N_29946);
nand U30067 (N_30067,N_29797,N_29712);
or U30068 (N_30068,N_29608,N_29748);
xor U30069 (N_30069,N_29955,N_29716);
nand U30070 (N_30070,N_29741,N_29786);
and U30071 (N_30071,N_29519,N_29665);
xor U30072 (N_30072,N_29992,N_29926);
and U30073 (N_30073,N_29658,N_29593);
or U30074 (N_30074,N_29882,N_29625);
and U30075 (N_30075,N_29753,N_29721);
nor U30076 (N_30076,N_29542,N_29815);
and U30077 (N_30077,N_29855,N_29787);
and U30078 (N_30078,N_29715,N_29524);
nand U30079 (N_30079,N_29906,N_29810);
or U30080 (N_30080,N_29622,N_29959);
or U30081 (N_30081,N_29948,N_29614);
and U30082 (N_30082,N_29515,N_29781);
or U30083 (N_30083,N_29979,N_29599);
nand U30084 (N_30084,N_29565,N_29897);
or U30085 (N_30085,N_29700,N_29745);
and U30086 (N_30086,N_29769,N_29617);
xor U30087 (N_30087,N_29915,N_29821);
and U30088 (N_30088,N_29900,N_29592);
or U30089 (N_30089,N_29640,N_29910);
nor U30090 (N_30090,N_29828,N_29941);
nor U30091 (N_30091,N_29541,N_29895);
and U30092 (N_30092,N_29993,N_29907);
or U30093 (N_30093,N_29796,N_29594);
and U30094 (N_30094,N_29935,N_29723);
xnor U30095 (N_30095,N_29545,N_29834);
or U30096 (N_30096,N_29823,N_29609);
xor U30097 (N_30097,N_29714,N_29572);
or U30098 (N_30098,N_29804,N_29963);
nor U30099 (N_30099,N_29648,N_29852);
nand U30100 (N_30100,N_29813,N_29726);
nor U30101 (N_30101,N_29782,N_29618);
or U30102 (N_30102,N_29692,N_29569);
nor U30103 (N_30103,N_29518,N_29535);
nand U30104 (N_30104,N_29643,N_29820);
and U30105 (N_30105,N_29957,N_29752);
or U30106 (N_30106,N_29574,N_29792);
nor U30107 (N_30107,N_29706,N_29756);
or U30108 (N_30108,N_29990,N_29682);
nor U30109 (N_30109,N_29520,N_29842);
nand U30110 (N_30110,N_29931,N_29693);
and U30111 (N_30111,N_29698,N_29691);
and U30112 (N_30112,N_29947,N_29639);
xor U30113 (N_30113,N_29848,N_29710);
xnor U30114 (N_30114,N_29987,N_29590);
or U30115 (N_30115,N_29996,N_29943);
or U30116 (N_30116,N_29630,N_29578);
nand U30117 (N_30117,N_29862,N_29896);
xnor U30118 (N_30118,N_29740,N_29514);
and U30119 (N_30119,N_29724,N_29918);
nand U30120 (N_30120,N_29883,N_29547);
or U30121 (N_30121,N_29601,N_29551);
or U30122 (N_30122,N_29672,N_29749);
nor U30123 (N_30123,N_29839,N_29929);
nand U30124 (N_30124,N_29623,N_29871);
and U30125 (N_30125,N_29557,N_29814);
nand U30126 (N_30126,N_29962,N_29634);
xnor U30127 (N_30127,N_29759,N_29811);
or U30128 (N_30128,N_29800,N_29982);
nor U30129 (N_30129,N_29909,N_29738);
xor U30130 (N_30130,N_29984,N_29764);
nand U30131 (N_30131,N_29527,N_29746);
nand U30132 (N_30132,N_29879,N_29967);
and U30133 (N_30133,N_29728,N_29743);
nand U30134 (N_30134,N_29595,N_29872);
nor U30135 (N_30135,N_29552,N_29951);
nor U30136 (N_30136,N_29995,N_29711);
nand U30137 (N_30137,N_29903,N_29824);
and U30138 (N_30138,N_29584,N_29678);
and U30139 (N_30139,N_29859,N_29780);
nor U30140 (N_30140,N_29636,N_29713);
or U30141 (N_30141,N_29677,N_29567);
nand U30142 (N_30142,N_29972,N_29536);
nand U30143 (N_30143,N_29663,N_29902);
or U30144 (N_30144,N_29597,N_29676);
nand U30145 (N_30145,N_29598,N_29645);
nand U30146 (N_30146,N_29794,N_29928);
or U30147 (N_30147,N_29731,N_29913);
nor U30148 (N_30148,N_29779,N_29525);
or U30149 (N_30149,N_29908,N_29554);
xor U30150 (N_30150,N_29881,N_29603);
nand U30151 (N_30151,N_29717,N_29973);
nor U30152 (N_30152,N_29983,N_29874);
nand U30153 (N_30153,N_29656,N_29563);
nor U30154 (N_30154,N_29971,N_29673);
nand U30155 (N_30155,N_29667,N_29866);
xor U30156 (N_30156,N_29562,N_29765);
xor U30157 (N_30157,N_29994,N_29933);
and U30158 (N_30158,N_29944,N_29522);
and U30159 (N_30159,N_29506,N_29833);
nor U30160 (N_30160,N_29644,N_29502);
or U30161 (N_30161,N_29826,N_29688);
xor U30162 (N_30162,N_29954,N_29938);
or U30163 (N_30163,N_29699,N_29517);
xor U30164 (N_30164,N_29893,N_29671);
nor U30165 (N_30165,N_29530,N_29916);
or U30166 (N_30166,N_29600,N_29772);
nor U30167 (N_30167,N_29953,N_29576);
and U30168 (N_30168,N_29546,N_29829);
nor U30169 (N_30169,N_29763,N_29850);
xnor U30170 (N_30170,N_29737,N_29771);
xnor U30171 (N_30171,N_29778,N_29891);
nand U30172 (N_30172,N_29932,N_29694);
or U30173 (N_30173,N_29806,N_29784);
nor U30174 (N_30174,N_29612,N_29980);
or U30175 (N_30175,N_29977,N_29832);
xor U30176 (N_30176,N_29695,N_29596);
nand U30177 (N_30177,N_29912,N_29960);
and U30178 (N_30178,N_29950,N_29613);
nand U30179 (N_30179,N_29548,N_29651);
nor U30180 (N_30180,N_29773,N_29577);
and U30181 (N_30181,N_29508,N_29633);
xnor U30182 (N_30182,N_29573,N_29793);
nor U30183 (N_30183,N_29605,N_29877);
xor U30184 (N_30184,N_29835,N_29923);
or U30185 (N_30185,N_29587,N_29560);
or U30186 (N_30186,N_29961,N_29624);
nand U30187 (N_30187,N_29968,N_29533);
or U30188 (N_30188,N_29680,N_29568);
nand U30189 (N_30189,N_29924,N_29889);
nor U30190 (N_30190,N_29555,N_29822);
nand U30191 (N_30191,N_29795,N_29683);
nor U30192 (N_30192,N_29790,N_29747);
and U30193 (N_30193,N_29729,N_29768);
or U30194 (N_30194,N_29841,N_29975);
xor U30195 (N_30195,N_29512,N_29544);
nor U30196 (N_30196,N_29861,N_29543);
or U30197 (N_30197,N_29785,N_29898);
nand U30198 (N_30198,N_29690,N_29610);
or U30199 (N_30199,N_29526,N_29540);
xor U30200 (N_30200,N_29920,N_29704);
and U30201 (N_30201,N_29616,N_29831);
and U30202 (N_30202,N_29550,N_29529);
xnor U30203 (N_30203,N_29991,N_29978);
xnor U30204 (N_30204,N_29607,N_29686);
and U30205 (N_30205,N_29664,N_29854);
xnor U30206 (N_30206,N_29799,N_29697);
nor U30207 (N_30207,N_29681,N_29641);
and U30208 (N_30208,N_29825,N_29858);
xnor U30209 (N_30209,N_29838,N_29801);
nand U30210 (N_30210,N_29538,N_29722);
or U30211 (N_30211,N_29606,N_29720);
nand U30212 (N_30212,N_29988,N_29802);
xor U30213 (N_30213,N_29805,N_29727);
xnor U30214 (N_30214,N_29647,N_29840);
and U30215 (N_30215,N_29718,N_29864);
and U30216 (N_30216,N_29626,N_29582);
and U30217 (N_30217,N_29783,N_29604);
nand U30218 (N_30218,N_29659,N_29751);
or U30219 (N_30219,N_29558,N_29523);
xor U30220 (N_30220,N_29570,N_29999);
nand U30221 (N_30221,N_29760,N_29901);
and U30222 (N_30222,N_29940,N_29985);
nor U30223 (N_30223,N_29750,N_29846);
nor U30224 (N_30224,N_29853,N_29708);
nand U30225 (N_30225,N_29696,N_29964);
xnor U30226 (N_30226,N_29885,N_29867);
nand U30227 (N_30227,N_29934,N_29927);
or U30228 (N_30228,N_29564,N_29847);
or U30229 (N_30229,N_29637,N_29511);
nand U30230 (N_30230,N_29770,N_29956);
and U30231 (N_30231,N_29789,N_29689);
or U30232 (N_30232,N_29507,N_29521);
nand U30233 (N_30233,N_29807,N_29777);
or U30234 (N_30234,N_29966,N_29620);
xnor U30235 (N_30235,N_29589,N_29719);
or U30236 (N_30236,N_29702,N_29675);
nor U30237 (N_30237,N_29516,N_29925);
xor U30238 (N_30238,N_29662,N_29958);
nor U30239 (N_30239,N_29629,N_29725);
xnor U30240 (N_30240,N_29701,N_29812);
nand U30241 (N_30241,N_29735,N_29730);
nor U30242 (N_30242,N_29627,N_29875);
xor U30243 (N_30243,N_29857,N_29887);
or U30244 (N_30244,N_29969,N_29899);
nor U30245 (N_30245,N_29703,N_29817);
nand U30246 (N_30246,N_29997,N_29669);
or U30247 (N_30247,N_29914,N_29937);
nor U30248 (N_30248,N_29930,N_29758);
and U30249 (N_30249,N_29816,N_29739);
and U30250 (N_30250,N_29782,N_29700);
or U30251 (N_30251,N_29599,N_29580);
nand U30252 (N_30252,N_29805,N_29766);
nand U30253 (N_30253,N_29587,N_29977);
and U30254 (N_30254,N_29694,N_29879);
nand U30255 (N_30255,N_29544,N_29672);
and U30256 (N_30256,N_29767,N_29813);
and U30257 (N_30257,N_29627,N_29886);
or U30258 (N_30258,N_29561,N_29539);
and U30259 (N_30259,N_29504,N_29761);
or U30260 (N_30260,N_29671,N_29920);
or U30261 (N_30261,N_29862,N_29955);
and U30262 (N_30262,N_29612,N_29650);
nand U30263 (N_30263,N_29892,N_29655);
nor U30264 (N_30264,N_29587,N_29999);
and U30265 (N_30265,N_29550,N_29798);
xnor U30266 (N_30266,N_29652,N_29849);
xor U30267 (N_30267,N_29761,N_29988);
and U30268 (N_30268,N_29994,N_29686);
xor U30269 (N_30269,N_29861,N_29829);
and U30270 (N_30270,N_29790,N_29930);
nand U30271 (N_30271,N_29705,N_29906);
nand U30272 (N_30272,N_29969,N_29541);
nand U30273 (N_30273,N_29946,N_29975);
xor U30274 (N_30274,N_29937,N_29879);
nor U30275 (N_30275,N_29553,N_29584);
nor U30276 (N_30276,N_29684,N_29754);
or U30277 (N_30277,N_29567,N_29680);
nand U30278 (N_30278,N_29656,N_29804);
or U30279 (N_30279,N_29643,N_29641);
and U30280 (N_30280,N_29765,N_29741);
nor U30281 (N_30281,N_29533,N_29817);
xor U30282 (N_30282,N_29817,N_29909);
xor U30283 (N_30283,N_29761,N_29962);
nor U30284 (N_30284,N_29975,N_29855);
xor U30285 (N_30285,N_29960,N_29771);
and U30286 (N_30286,N_29934,N_29837);
nand U30287 (N_30287,N_29594,N_29633);
nand U30288 (N_30288,N_29894,N_29773);
nor U30289 (N_30289,N_29560,N_29917);
nor U30290 (N_30290,N_29522,N_29736);
nor U30291 (N_30291,N_29796,N_29826);
nand U30292 (N_30292,N_29865,N_29659);
and U30293 (N_30293,N_29681,N_29584);
xor U30294 (N_30294,N_29554,N_29785);
nand U30295 (N_30295,N_29638,N_29993);
xnor U30296 (N_30296,N_29598,N_29579);
nor U30297 (N_30297,N_29982,N_29758);
or U30298 (N_30298,N_29710,N_29617);
and U30299 (N_30299,N_29972,N_29692);
or U30300 (N_30300,N_29840,N_29972);
nor U30301 (N_30301,N_29916,N_29580);
nor U30302 (N_30302,N_29622,N_29672);
or U30303 (N_30303,N_29771,N_29749);
nand U30304 (N_30304,N_29660,N_29687);
nand U30305 (N_30305,N_29710,N_29797);
nand U30306 (N_30306,N_29707,N_29685);
nand U30307 (N_30307,N_29942,N_29917);
nor U30308 (N_30308,N_29908,N_29719);
or U30309 (N_30309,N_29560,N_29607);
nor U30310 (N_30310,N_29750,N_29718);
and U30311 (N_30311,N_29913,N_29858);
or U30312 (N_30312,N_29682,N_29837);
and U30313 (N_30313,N_29629,N_29612);
and U30314 (N_30314,N_29940,N_29922);
xnor U30315 (N_30315,N_29920,N_29773);
nor U30316 (N_30316,N_29826,N_29701);
or U30317 (N_30317,N_29609,N_29846);
and U30318 (N_30318,N_29685,N_29952);
xor U30319 (N_30319,N_29610,N_29781);
xor U30320 (N_30320,N_29768,N_29739);
xnor U30321 (N_30321,N_29773,N_29778);
nand U30322 (N_30322,N_29540,N_29972);
nand U30323 (N_30323,N_29767,N_29948);
xnor U30324 (N_30324,N_29969,N_29946);
nand U30325 (N_30325,N_29953,N_29903);
nor U30326 (N_30326,N_29733,N_29547);
and U30327 (N_30327,N_29607,N_29911);
xnor U30328 (N_30328,N_29519,N_29549);
or U30329 (N_30329,N_29843,N_29923);
and U30330 (N_30330,N_29523,N_29905);
nand U30331 (N_30331,N_29764,N_29604);
or U30332 (N_30332,N_29636,N_29831);
or U30333 (N_30333,N_29683,N_29654);
nand U30334 (N_30334,N_29510,N_29720);
or U30335 (N_30335,N_29554,N_29784);
nor U30336 (N_30336,N_29668,N_29585);
and U30337 (N_30337,N_29933,N_29623);
nand U30338 (N_30338,N_29619,N_29962);
nand U30339 (N_30339,N_29701,N_29868);
nor U30340 (N_30340,N_29826,N_29564);
xnor U30341 (N_30341,N_29822,N_29864);
xor U30342 (N_30342,N_29902,N_29589);
nand U30343 (N_30343,N_29847,N_29603);
or U30344 (N_30344,N_29623,N_29954);
or U30345 (N_30345,N_29622,N_29603);
and U30346 (N_30346,N_29574,N_29946);
xor U30347 (N_30347,N_29874,N_29525);
nor U30348 (N_30348,N_29774,N_29920);
and U30349 (N_30349,N_29908,N_29979);
and U30350 (N_30350,N_29613,N_29517);
nand U30351 (N_30351,N_29822,N_29585);
or U30352 (N_30352,N_29680,N_29663);
and U30353 (N_30353,N_29642,N_29809);
nor U30354 (N_30354,N_29807,N_29889);
nand U30355 (N_30355,N_29814,N_29964);
and U30356 (N_30356,N_29672,N_29782);
or U30357 (N_30357,N_29708,N_29604);
or U30358 (N_30358,N_29506,N_29943);
and U30359 (N_30359,N_29829,N_29597);
nor U30360 (N_30360,N_29621,N_29834);
nor U30361 (N_30361,N_29926,N_29560);
nor U30362 (N_30362,N_29731,N_29585);
nor U30363 (N_30363,N_29618,N_29981);
xor U30364 (N_30364,N_29608,N_29656);
and U30365 (N_30365,N_29688,N_29854);
and U30366 (N_30366,N_29936,N_29540);
and U30367 (N_30367,N_29970,N_29779);
and U30368 (N_30368,N_29678,N_29697);
or U30369 (N_30369,N_29801,N_29861);
and U30370 (N_30370,N_29676,N_29870);
nor U30371 (N_30371,N_29788,N_29983);
nand U30372 (N_30372,N_29599,N_29634);
nor U30373 (N_30373,N_29608,N_29967);
nor U30374 (N_30374,N_29906,N_29646);
and U30375 (N_30375,N_29918,N_29921);
nor U30376 (N_30376,N_29695,N_29599);
nand U30377 (N_30377,N_29770,N_29885);
and U30378 (N_30378,N_29618,N_29659);
or U30379 (N_30379,N_29901,N_29686);
and U30380 (N_30380,N_29743,N_29836);
nor U30381 (N_30381,N_29598,N_29781);
xor U30382 (N_30382,N_29751,N_29705);
nand U30383 (N_30383,N_29557,N_29629);
nand U30384 (N_30384,N_29504,N_29688);
or U30385 (N_30385,N_29982,N_29612);
nand U30386 (N_30386,N_29529,N_29668);
xor U30387 (N_30387,N_29765,N_29829);
nor U30388 (N_30388,N_29937,N_29847);
or U30389 (N_30389,N_29771,N_29981);
and U30390 (N_30390,N_29864,N_29663);
nor U30391 (N_30391,N_29855,N_29768);
nand U30392 (N_30392,N_29858,N_29685);
or U30393 (N_30393,N_29800,N_29527);
and U30394 (N_30394,N_29588,N_29989);
and U30395 (N_30395,N_29734,N_29976);
nand U30396 (N_30396,N_29927,N_29516);
xor U30397 (N_30397,N_29741,N_29506);
and U30398 (N_30398,N_29983,N_29827);
nand U30399 (N_30399,N_29919,N_29972);
xnor U30400 (N_30400,N_29754,N_29588);
xor U30401 (N_30401,N_29637,N_29574);
and U30402 (N_30402,N_29655,N_29933);
nor U30403 (N_30403,N_29810,N_29525);
nor U30404 (N_30404,N_29954,N_29893);
and U30405 (N_30405,N_29508,N_29522);
or U30406 (N_30406,N_29795,N_29721);
or U30407 (N_30407,N_29776,N_29598);
and U30408 (N_30408,N_29693,N_29965);
nor U30409 (N_30409,N_29955,N_29596);
xnor U30410 (N_30410,N_29545,N_29935);
or U30411 (N_30411,N_29543,N_29629);
nor U30412 (N_30412,N_29931,N_29871);
or U30413 (N_30413,N_29738,N_29863);
or U30414 (N_30414,N_29942,N_29895);
or U30415 (N_30415,N_29980,N_29511);
xor U30416 (N_30416,N_29980,N_29706);
nor U30417 (N_30417,N_29709,N_29505);
xnor U30418 (N_30418,N_29714,N_29639);
and U30419 (N_30419,N_29758,N_29964);
or U30420 (N_30420,N_29790,N_29510);
nand U30421 (N_30421,N_29903,N_29864);
nor U30422 (N_30422,N_29537,N_29933);
xnor U30423 (N_30423,N_29786,N_29688);
xnor U30424 (N_30424,N_29862,N_29681);
nand U30425 (N_30425,N_29917,N_29892);
nor U30426 (N_30426,N_29945,N_29734);
or U30427 (N_30427,N_29933,N_29816);
xor U30428 (N_30428,N_29764,N_29637);
and U30429 (N_30429,N_29597,N_29691);
nand U30430 (N_30430,N_29707,N_29745);
nand U30431 (N_30431,N_29816,N_29884);
nor U30432 (N_30432,N_29699,N_29512);
xnor U30433 (N_30433,N_29723,N_29667);
xnor U30434 (N_30434,N_29884,N_29960);
xnor U30435 (N_30435,N_29814,N_29724);
xnor U30436 (N_30436,N_29747,N_29520);
and U30437 (N_30437,N_29633,N_29507);
xor U30438 (N_30438,N_29554,N_29788);
nor U30439 (N_30439,N_29792,N_29942);
xor U30440 (N_30440,N_29625,N_29697);
and U30441 (N_30441,N_29751,N_29939);
nand U30442 (N_30442,N_29977,N_29912);
xnor U30443 (N_30443,N_29841,N_29643);
xnor U30444 (N_30444,N_29955,N_29527);
xor U30445 (N_30445,N_29865,N_29678);
and U30446 (N_30446,N_29858,N_29994);
and U30447 (N_30447,N_29693,N_29733);
nand U30448 (N_30448,N_29690,N_29631);
nor U30449 (N_30449,N_29597,N_29840);
or U30450 (N_30450,N_29860,N_29906);
xor U30451 (N_30451,N_29629,N_29576);
and U30452 (N_30452,N_29930,N_29835);
xnor U30453 (N_30453,N_29778,N_29838);
xnor U30454 (N_30454,N_29511,N_29746);
xnor U30455 (N_30455,N_29621,N_29901);
xnor U30456 (N_30456,N_29707,N_29539);
nor U30457 (N_30457,N_29579,N_29616);
and U30458 (N_30458,N_29547,N_29880);
nor U30459 (N_30459,N_29602,N_29631);
xnor U30460 (N_30460,N_29703,N_29989);
nand U30461 (N_30461,N_29565,N_29684);
nor U30462 (N_30462,N_29542,N_29988);
or U30463 (N_30463,N_29784,N_29511);
nor U30464 (N_30464,N_29669,N_29539);
xnor U30465 (N_30465,N_29750,N_29588);
xnor U30466 (N_30466,N_29979,N_29868);
nand U30467 (N_30467,N_29993,N_29531);
and U30468 (N_30468,N_29860,N_29593);
xor U30469 (N_30469,N_29847,N_29948);
nor U30470 (N_30470,N_29774,N_29655);
xnor U30471 (N_30471,N_29748,N_29985);
or U30472 (N_30472,N_29534,N_29703);
nor U30473 (N_30473,N_29594,N_29683);
nor U30474 (N_30474,N_29684,N_29718);
nand U30475 (N_30475,N_29725,N_29823);
nand U30476 (N_30476,N_29571,N_29936);
or U30477 (N_30477,N_29877,N_29903);
and U30478 (N_30478,N_29691,N_29986);
nor U30479 (N_30479,N_29818,N_29716);
nand U30480 (N_30480,N_29644,N_29929);
and U30481 (N_30481,N_29624,N_29910);
and U30482 (N_30482,N_29753,N_29881);
or U30483 (N_30483,N_29791,N_29877);
xnor U30484 (N_30484,N_29603,N_29730);
or U30485 (N_30485,N_29801,N_29973);
xnor U30486 (N_30486,N_29635,N_29722);
nor U30487 (N_30487,N_29835,N_29541);
nor U30488 (N_30488,N_29531,N_29544);
or U30489 (N_30489,N_29721,N_29933);
nand U30490 (N_30490,N_29829,N_29529);
xnor U30491 (N_30491,N_29792,N_29635);
nand U30492 (N_30492,N_29902,N_29544);
and U30493 (N_30493,N_29893,N_29632);
nand U30494 (N_30494,N_29939,N_29717);
and U30495 (N_30495,N_29660,N_29967);
nor U30496 (N_30496,N_29739,N_29984);
nor U30497 (N_30497,N_29594,N_29709);
xnor U30498 (N_30498,N_29738,N_29996);
nor U30499 (N_30499,N_29658,N_29928);
nor U30500 (N_30500,N_30472,N_30104);
xor U30501 (N_30501,N_30232,N_30471);
xor U30502 (N_30502,N_30329,N_30301);
or U30503 (N_30503,N_30206,N_30400);
nand U30504 (N_30504,N_30088,N_30045);
xor U30505 (N_30505,N_30079,N_30346);
or U30506 (N_30506,N_30057,N_30441);
nor U30507 (N_30507,N_30489,N_30164);
or U30508 (N_30508,N_30001,N_30221);
or U30509 (N_30509,N_30408,N_30024);
or U30510 (N_30510,N_30302,N_30437);
and U30511 (N_30511,N_30092,N_30117);
nand U30512 (N_30512,N_30429,N_30373);
or U30513 (N_30513,N_30319,N_30043);
xor U30514 (N_30514,N_30436,N_30038);
nand U30515 (N_30515,N_30287,N_30332);
and U30516 (N_30516,N_30184,N_30245);
or U30517 (N_30517,N_30390,N_30280);
nand U30518 (N_30518,N_30047,N_30014);
nand U30519 (N_30519,N_30403,N_30303);
nand U30520 (N_30520,N_30106,N_30101);
xnor U30521 (N_30521,N_30359,N_30476);
xor U30522 (N_30522,N_30034,N_30064);
xnor U30523 (N_30523,N_30149,N_30278);
and U30524 (N_30524,N_30007,N_30285);
nor U30525 (N_30525,N_30353,N_30158);
or U30526 (N_30526,N_30208,N_30192);
nor U30527 (N_30527,N_30139,N_30161);
nor U30528 (N_30528,N_30115,N_30248);
or U30529 (N_30529,N_30312,N_30250);
and U30530 (N_30530,N_30456,N_30182);
xor U30531 (N_30531,N_30442,N_30237);
or U30532 (N_30532,N_30316,N_30173);
or U30533 (N_30533,N_30496,N_30228);
and U30534 (N_30534,N_30027,N_30167);
xor U30535 (N_30535,N_30255,N_30444);
and U30536 (N_30536,N_30454,N_30314);
and U30537 (N_30537,N_30410,N_30416);
or U30538 (N_30538,N_30077,N_30053);
and U30539 (N_30539,N_30483,N_30217);
nand U30540 (N_30540,N_30487,N_30011);
and U30541 (N_30541,N_30129,N_30130);
and U30542 (N_30542,N_30062,N_30016);
xor U30543 (N_30543,N_30465,N_30426);
and U30544 (N_30544,N_30058,N_30434);
nand U30545 (N_30545,N_30290,N_30012);
nor U30546 (N_30546,N_30428,N_30417);
nor U30547 (N_30547,N_30291,N_30181);
nor U30548 (N_30548,N_30404,N_30041);
xnor U30549 (N_30549,N_30275,N_30296);
and U30550 (N_30550,N_30451,N_30387);
xnor U30551 (N_30551,N_30455,N_30499);
nand U30552 (N_30552,N_30121,N_30449);
and U30553 (N_30553,N_30243,N_30003);
nand U30554 (N_30554,N_30087,N_30098);
nor U30555 (N_30555,N_30218,N_30289);
nor U30556 (N_30556,N_30485,N_30393);
nand U30557 (N_30557,N_30475,N_30055);
or U30558 (N_30558,N_30096,N_30462);
or U30559 (N_30559,N_30376,N_30137);
and U30560 (N_30560,N_30239,N_30249);
and U30561 (N_30561,N_30153,N_30481);
nand U30562 (N_30562,N_30190,N_30086);
xnor U30563 (N_30563,N_30262,N_30059);
or U30564 (N_30564,N_30424,N_30411);
nand U30565 (N_30565,N_30107,N_30398);
xor U30566 (N_30566,N_30174,N_30150);
or U30567 (N_30567,N_30259,N_30395);
and U30568 (N_30568,N_30268,N_30327);
xnor U30569 (N_30569,N_30131,N_30214);
nand U30570 (N_30570,N_30421,N_30030);
nand U30571 (N_30571,N_30060,N_30308);
xnor U30572 (N_30572,N_30478,N_30226);
or U30573 (N_30573,N_30051,N_30028);
and U30574 (N_30574,N_30464,N_30215);
nor U30575 (N_30575,N_30343,N_30169);
and U30576 (N_30576,N_30136,N_30486);
nor U30577 (N_30577,N_30374,N_30467);
xnor U30578 (N_30578,N_30317,N_30271);
or U30579 (N_30579,N_30146,N_30324);
and U30580 (N_30580,N_30432,N_30273);
nand U30581 (N_30581,N_30363,N_30349);
nand U30582 (N_30582,N_30490,N_30364);
and U30583 (N_30583,N_30369,N_30004);
nand U30584 (N_30584,N_30293,N_30365);
nand U30585 (N_30585,N_30281,N_30265);
and U30586 (N_30586,N_30254,N_30144);
and U30587 (N_30587,N_30207,N_30492);
or U30588 (N_30588,N_30128,N_30223);
or U30589 (N_30589,N_30361,N_30070);
xor U30590 (N_30590,N_30341,N_30307);
and U30591 (N_30591,N_30187,N_30396);
nand U30592 (N_30592,N_30105,N_30066);
nor U30593 (N_30593,N_30233,N_30216);
nor U30594 (N_30594,N_30103,N_30344);
nor U30595 (N_30595,N_30056,N_30443);
xor U30596 (N_30596,N_30019,N_30141);
xor U30597 (N_30597,N_30170,N_30331);
or U30598 (N_30598,N_30219,N_30160);
and U30599 (N_30599,N_30298,N_30340);
xor U30600 (N_30600,N_30292,N_30241);
xor U30601 (N_30601,N_30222,N_30247);
nor U30602 (N_30602,N_30147,N_30392);
xor U30603 (N_30603,N_30017,N_30163);
and U30604 (N_30604,N_30383,N_30031);
and U30605 (N_30605,N_30042,N_30157);
or U30606 (N_30606,N_30176,N_30350);
and U30607 (N_30607,N_30380,N_30360);
and U30608 (N_30608,N_30235,N_30334);
or U30609 (N_30609,N_30162,N_30430);
nand U30610 (N_30610,N_30382,N_30282);
or U30611 (N_30611,N_30013,N_30304);
xor U30612 (N_30612,N_30212,N_30457);
xor U30613 (N_30613,N_30269,N_30132);
or U30614 (N_30614,N_30246,N_30305);
and U30615 (N_30615,N_30102,N_30109);
and U30616 (N_30616,N_30253,N_30354);
nor U30617 (N_30617,N_30185,N_30209);
or U30618 (N_30618,N_30491,N_30110);
nor U30619 (N_30619,N_30021,N_30286);
xnor U30620 (N_30620,N_30084,N_30463);
or U30621 (N_30621,N_30321,N_30357);
nand U30622 (N_30622,N_30439,N_30193);
nor U30623 (N_30623,N_30069,N_30065);
and U30624 (N_30624,N_30116,N_30094);
nand U30625 (N_30625,N_30122,N_30493);
or U30626 (N_30626,N_30099,N_30119);
nor U30627 (N_30627,N_30347,N_30333);
or U30628 (N_30628,N_30072,N_30126);
and U30629 (N_30629,N_30389,N_30358);
xnor U30630 (N_30630,N_30201,N_30111);
nand U30631 (N_30631,N_30191,N_30440);
nand U30632 (N_30632,N_30309,N_30022);
xnor U30633 (N_30633,N_30166,N_30260);
nand U30634 (N_30634,N_30234,N_30171);
or U30635 (N_30635,N_30469,N_30238);
xor U30636 (N_30636,N_30211,N_30230);
xor U30637 (N_30637,N_30198,N_30488);
and U30638 (N_30638,N_30048,N_30446);
and U30639 (N_30639,N_30095,N_30155);
or U30640 (N_30640,N_30325,N_30251);
nand U30641 (N_30641,N_30406,N_30080);
nand U30642 (N_30642,N_30023,N_30152);
or U30643 (N_30643,N_30090,N_30330);
xor U30644 (N_30644,N_30431,N_30040);
or U30645 (N_30645,N_30118,N_30458);
xnor U30646 (N_30646,N_30412,N_30256);
xor U30647 (N_30647,N_30477,N_30267);
xnor U30648 (N_30648,N_30100,N_30480);
nand U30649 (N_30649,N_30039,N_30266);
and U30650 (N_30650,N_30140,N_30336);
or U30651 (N_30651,N_30474,N_30366);
or U30652 (N_30652,N_30371,N_30177);
nor U30653 (N_30653,N_30220,N_30264);
nor U30654 (N_30654,N_30037,N_30370);
or U30655 (N_30655,N_30401,N_30295);
nand U30656 (N_30656,N_30120,N_30470);
and U30657 (N_30657,N_30397,N_30418);
or U30658 (N_30658,N_30448,N_30438);
nand U30659 (N_30659,N_30355,N_30083);
or U30660 (N_30660,N_30097,N_30414);
nor U30661 (N_30661,N_30026,N_30338);
nor U30662 (N_30662,N_30089,N_30135);
nand U30663 (N_30663,N_30091,N_30288);
nor U30664 (N_30664,N_30468,N_30068);
and U30665 (N_30665,N_30323,N_30210);
and U30666 (N_30666,N_30378,N_30172);
or U30667 (N_30667,N_30335,N_30032);
or U30668 (N_30668,N_30213,N_30018);
nor U30669 (N_30669,N_30420,N_30054);
nor U30670 (N_30670,N_30284,N_30180);
and U30671 (N_30671,N_30061,N_30033);
nand U30672 (N_30672,N_30000,N_30294);
or U30673 (N_30673,N_30276,N_30050);
and U30674 (N_30674,N_30459,N_30231);
nand U30675 (N_30675,N_30482,N_30452);
and U30676 (N_30676,N_30081,N_30203);
and U30677 (N_30677,N_30405,N_30071);
nor U30678 (N_30678,N_30339,N_30460);
or U30679 (N_30679,N_30311,N_30367);
xor U30680 (N_30680,N_30461,N_30299);
and U30681 (N_30681,N_30386,N_30020);
or U30682 (N_30682,N_30076,N_30318);
and U30683 (N_30683,N_30466,N_30379);
and U30684 (N_30684,N_30138,N_30008);
and U30685 (N_30685,N_30252,N_30029);
or U30686 (N_30686,N_30010,N_30204);
or U30687 (N_30687,N_30052,N_30124);
xnor U30688 (N_30688,N_30375,N_30112);
xor U30689 (N_30689,N_30326,N_30306);
xnor U30690 (N_30690,N_30188,N_30377);
xor U30691 (N_30691,N_30315,N_30351);
and U30692 (N_30692,N_30345,N_30189);
or U30693 (N_30693,N_30384,N_30399);
and U30694 (N_30694,N_30168,N_30224);
and U30695 (N_30695,N_30283,N_30391);
nand U30696 (N_30696,N_30409,N_30046);
nor U30697 (N_30697,N_30372,N_30356);
nand U30698 (N_30698,N_30009,N_30342);
nand U30699 (N_30699,N_30320,N_30242);
xor U30700 (N_30700,N_30073,N_30183);
and U30701 (N_30701,N_30422,N_30229);
and U30702 (N_30702,N_30415,N_30368);
and U30703 (N_30703,N_30049,N_30297);
nand U30704 (N_30704,N_30082,N_30423);
and U30705 (N_30705,N_30225,N_30125);
nor U30706 (N_30706,N_30165,N_30258);
nor U30707 (N_30707,N_30322,N_30175);
or U30708 (N_30708,N_30093,N_30044);
xnor U30709 (N_30709,N_30453,N_30145);
and U30710 (N_30710,N_30002,N_30337);
nand U30711 (N_30711,N_30148,N_30435);
nor U30712 (N_30712,N_30447,N_30194);
or U30713 (N_30713,N_30114,N_30272);
and U30714 (N_30714,N_30133,N_30200);
xor U30715 (N_30715,N_30075,N_30108);
nor U30716 (N_30716,N_30036,N_30006);
and U30717 (N_30717,N_30279,N_30202);
or U30718 (N_30718,N_30310,N_30479);
xor U30719 (N_30719,N_30085,N_30199);
xor U30720 (N_30720,N_30413,N_30328);
xor U30721 (N_30721,N_30484,N_30419);
nor U30722 (N_30722,N_30227,N_30261);
xor U30723 (N_30723,N_30352,N_30427);
xnor U30724 (N_30724,N_30074,N_30381);
nor U30725 (N_30725,N_30154,N_30196);
and U30726 (N_30726,N_30394,N_30425);
nor U30727 (N_30727,N_30388,N_30300);
xnor U30728 (N_30728,N_30186,N_30494);
xnor U30729 (N_30729,N_30005,N_30159);
nor U30730 (N_30730,N_30134,N_30277);
nand U30731 (N_30731,N_30362,N_30450);
xnor U30732 (N_30732,N_30495,N_30195);
nor U30733 (N_30733,N_30113,N_30078);
nor U30734 (N_30734,N_30156,N_30143);
xor U30735 (N_30735,N_30123,N_30240);
nand U30736 (N_30736,N_30385,N_30263);
nor U30737 (N_30737,N_30015,N_30270);
or U30738 (N_30738,N_30205,N_30473);
nor U30739 (N_30739,N_30445,N_30348);
and U30740 (N_30740,N_30274,N_30063);
and U30741 (N_30741,N_30151,N_30498);
or U30742 (N_30742,N_30179,N_30257);
or U30743 (N_30743,N_30035,N_30236);
nor U30744 (N_30744,N_30067,N_30025);
or U30745 (N_30745,N_30197,N_30407);
or U30746 (N_30746,N_30433,N_30127);
xnor U30747 (N_30747,N_30497,N_30178);
or U30748 (N_30748,N_30142,N_30402);
or U30749 (N_30749,N_30313,N_30244);
or U30750 (N_30750,N_30288,N_30013);
nor U30751 (N_30751,N_30427,N_30046);
and U30752 (N_30752,N_30313,N_30044);
xor U30753 (N_30753,N_30204,N_30328);
and U30754 (N_30754,N_30152,N_30142);
and U30755 (N_30755,N_30147,N_30315);
nor U30756 (N_30756,N_30133,N_30272);
nand U30757 (N_30757,N_30282,N_30236);
or U30758 (N_30758,N_30213,N_30056);
nand U30759 (N_30759,N_30160,N_30339);
and U30760 (N_30760,N_30469,N_30286);
xnor U30761 (N_30761,N_30331,N_30095);
nor U30762 (N_30762,N_30225,N_30373);
nand U30763 (N_30763,N_30388,N_30430);
nand U30764 (N_30764,N_30325,N_30178);
and U30765 (N_30765,N_30064,N_30202);
nor U30766 (N_30766,N_30380,N_30191);
or U30767 (N_30767,N_30300,N_30420);
and U30768 (N_30768,N_30265,N_30296);
and U30769 (N_30769,N_30108,N_30492);
and U30770 (N_30770,N_30483,N_30015);
or U30771 (N_30771,N_30071,N_30284);
nand U30772 (N_30772,N_30305,N_30465);
nor U30773 (N_30773,N_30028,N_30341);
nand U30774 (N_30774,N_30414,N_30357);
and U30775 (N_30775,N_30238,N_30141);
nor U30776 (N_30776,N_30128,N_30098);
or U30777 (N_30777,N_30382,N_30150);
and U30778 (N_30778,N_30076,N_30445);
and U30779 (N_30779,N_30100,N_30450);
or U30780 (N_30780,N_30293,N_30130);
nor U30781 (N_30781,N_30097,N_30270);
nor U30782 (N_30782,N_30194,N_30176);
nand U30783 (N_30783,N_30140,N_30292);
xor U30784 (N_30784,N_30053,N_30150);
nor U30785 (N_30785,N_30183,N_30110);
xor U30786 (N_30786,N_30495,N_30135);
or U30787 (N_30787,N_30012,N_30388);
nor U30788 (N_30788,N_30212,N_30047);
and U30789 (N_30789,N_30002,N_30498);
and U30790 (N_30790,N_30453,N_30431);
nand U30791 (N_30791,N_30141,N_30194);
nor U30792 (N_30792,N_30050,N_30265);
nor U30793 (N_30793,N_30214,N_30154);
nor U30794 (N_30794,N_30255,N_30009);
or U30795 (N_30795,N_30419,N_30400);
nor U30796 (N_30796,N_30309,N_30358);
and U30797 (N_30797,N_30328,N_30375);
xnor U30798 (N_30798,N_30483,N_30054);
nand U30799 (N_30799,N_30045,N_30466);
nand U30800 (N_30800,N_30421,N_30474);
xnor U30801 (N_30801,N_30152,N_30089);
or U30802 (N_30802,N_30326,N_30068);
xor U30803 (N_30803,N_30350,N_30175);
nand U30804 (N_30804,N_30488,N_30265);
nor U30805 (N_30805,N_30216,N_30304);
or U30806 (N_30806,N_30229,N_30268);
or U30807 (N_30807,N_30269,N_30172);
nand U30808 (N_30808,N_30127,N_30149);
xnor U30809 (N_30809,N_30135,N_30269);
nand U30810 (N_30810,N_30090,N_30365);
nor U30811 (N_30811,N_30305,N_30079);
nor U30812 (N_30812,N_30238,N_30495);
and U30813 (N_30813,N_30398,N_30000);
xnor U30814 (N_30814,N_30466,N_30012);
nor U30815 (N_30815,N_30455,N_30211);
and U30816 (N_30816,N_30339,N_30158);
nor U30817 (N_30817,N_30141,N_30197);
and U30818 (N_30818,N_30441,N_30433);
xnor U30819 (N_30819,N_30207,N_30050);
xnor U30820 (N_30820,N_30047,N_30498);
nor U30821 (N_30821,N_30248,N_30250);
nor U30822 (N_30822,N_30395,N_30332);
xor U30823 (N_30823,N_30157,N_30230);
xor U30824 (N_30824,N_30435,N_30483);
xor U30825 (N_30825,N_30164,N_30066);
nand U30826 (N_30826,N_30130,N_30349);
nor U30827 (N_30827,N_30386,N_30153);
nand U30828 (N_30828,N_30001,N_30383);
and U30829 (N_30829,N_30044,N_30365);
nand U30830 (N_30830,N_30042,N_30420);
nand U30831 (N_30831,N_30268,N_30142);
nand U30832 (N_30832,N_30436,N_30141);
xor U30833 (N_30833,N_30030,N_30266);
xnor U30834 (N_30834,N_30114,N_30463);
or U30835 (N_30835,N_30113,N_30233);
or U30836 (N_30836,N_30086,N_30361);
nor U30837 (N_30837,N_30422,N_30277);
nand U30838 (N_30838,N_30427,N_30268);
nand U30839 (N_30839,N_30312,N_30290);
and U30840 (N_30840,N_30005,N_30332);
nand U30841 (N_30841,N_30377,N_30261);
nand U30842 (N_30842,N_30223,N_30377);
nor U30843 (N_30843,N_30192,N_30137);
or U30844 (N_30844,N_30298,N_30147);
nor U30845 (N_30845,N_30408,N_30417);
and U30846 (N_30846,N_30062,N_30297);
xnor U30847 (N_30847,N_30119,N_30141);
nand U30848 (N_30848,N_30018,N_30493);
or U30849 (N_30849,N_30126,N_30004);
or U30850 (N_30850,N_30221,N_30241);
xnor U30851 (N_30851,N_30175,N_30362);
and U30852 (N_30852,N_30490,N_30290);
or U30853 (N_30853,N_30356,N_30261);
xor U30854 (N_30854,N_30040,N_30338);
nor U30855 (N_30855,N_30258,N_30379);
xor U30856 (N_30856,N_30076,N_30222);
xnor U30857 (N_30857,N_30412,N_30350);
nor U30858 (N_30858,N_30395,N_30169);
nand U30859 (N_30859,N_30223,N_30050);
or U30860 (N_30860,N_30307,N_30412);
xor U30861 (N_30861,N_30227,N_30319);
nand U30862 (N_30862,N_30053,N_30327);
or U30863 (N_30863,N_30429,N_30296);
and U30864 (N_30864,N_30063,N_30302);
nor U30865 (N_30865,N_30204,N_30129);
and U30866 (N_30866,N_30348,N_30371);
nand U30867 (N_30867,N_30219,N_30190);
or U30868 (N_30868,N_30010,N_30370);
and U30869 (N_30869,N_30077,N_30333);
xor U30870 (N_30870,N_30049,N_30339);
and U30871 (N_30871,N_30029,N_30270);
and U30872 (N_30872,N_30407,N_30257);
xor U30873 (N_30873,N_30191,N_30491);
and U30874 (N_30874,N_30143,N_30034);
nor U30875 (N_30875,N_30361,N_30416);
and U30876 (N_30876,N_30171,N_30064);
nor U30877 (N_30877,N_30025,N_30338);
and U30878 (N_30878,N_30286,N_30237);
and U30879 (N_30879,N_30055,N_30300);
or U30880 (N_30880,N_30067,N_30240);
or U30881 (N_30881,N_30438,N_30014);
nand U30882 (N_30882,N_30387,N_30465);
nor U30883 (N_30883,N_30040,N_30441);
or U30884 (N_30884,N_30419,N_30161);
and U30885 (N_30885,N_30458,N_30256);
nand U30886 (N_30886,N_30264,N_30077);
nand U30887 (N_30887,N_30023,N_30334);
nand U30888 (N_30888,N_30126,N_30095);
nor U30889 (N_30889,N_30328,N_30490);
nor U30890 (N_30890,N_30254,N_30420);
and U30891 (N_30891,N_30243,N_30211);
and U30892 (N_30892,N_30397,N_30161);
and U30893 (N_30893,N_30187,N_30233);
nand U30894 (N_30894,N_30111,N_30084);
nand U30895 (N_30895,N_30316,N_30250);
and U30896 (N_30896,N_30388,N_30345);
xnor U30897 (N_30897,N_30277,N_30184);
nand U30898 (N_30898,N_30100,N_30291);
nand U30899 (N_30899,N_30179,N_30383);
and U30900 (N_30900,N_30350,N_30232);
nand U30901 (N_30901,N_30052,N_30485);
or U30902 (N_30902,N_30265,N_30298);
and U30903 (N_30903,N_30183,N_30118);
or U30904 (N_30904,N_30273,N_30277);
xnor U30905 (N_30905,N_30296,N_30452);
xor U30906 (N_30906,N_30023,N_30292);
and U30907 (N_30907,N_30300,N_30123);
and U30908 (N_30908,N_30364,N_30273);
or U30909 (N_30909,N_30242,N_30172);
or U30910 (N_30910,N_30002,N_30299);
or U30911 (N_30911,N_30336,N_30077);
nand U30912 (N_30912,N_30364,N_30226);
or U30913 (N_30913,N_30005,N_30091);
nand U30914 (N_30914,N_30055,N_30134);
and U30915 (N_30915,N_30364,N_30463);
xnor U30916 (N_30916,N_30395,N_30436);
and U30917 (N_30917,N_30291,N_30251);
nor U30918 (N_30918,N_30377,N_30139);
nor U30919 (N_30919,N_30030,N_30454);
nand U30920 (N_30920,N_30384,N_30260);
xnor U30921 (N_30921,N_30488,N_30371);
nand U30922 (N_30922,N_30193,N_30057);
xor U30923 (N_30923,N_30444,N_30026);
nand U30924 (N_30924,N_30420,N_30096);
and U30925 (N_30925,N_30257,N_30482);
and U30926 (N_30926,N_30427,N_30244);
xnor U30927 (N_30927,N_30020,N_30093);
nor U30928 (N_30928,N_30426,N_30072);
or U30929 (N_30929,N_30352,N_30268);
or U30930 (N_30930,N_30361,N_30137);
nand U30931 (N_30931,N_30420,N_30076);
nand U30932 (N_30932,N_30032,N_30417);
or U30933 (N_30933,N_30134,N_30213);
and U30934 (N_30934,N_30370,N_30109);
or U30935 (N_30935,N_30059,N_30136);
nor U30936 (N_30936,N_30246,N_30239);
and U30937 (N_30937,N_30233,N_30011);
nand U30938 (N_30938,N_30329,N_30244);
or U30939 (N_30939,N_30071,N_30417);
xor U30940 (N_30940,N_30175,N_30078);
xnor U30941 (N_30941,N_30430,N_30449);
nor U30942 (N_30942,N_30316,N_30353);
nand U30943 (N_30943,N_30195,N_30430);
nor U30944 (N_30944,N_30360,N_30024);
nor U30945 (N_30945,N_30466,N_30078);
nor U30946 (N_30946,N_30327,N_30304);
and U30947 (N_30947,N_30283,N_30261);
xor U30948 (N_30948,N_30289,N_30132);
xor U30949 (N_30949,N_30217,N_30233);
and U30950 (N_30950,N_30103,N_30405);
or U30951 (N_30951,N_30493,N_30274);
and U30952 (N_30952,N_30077,N_30419);
and U30953 (N_30953,N_30381,N_30329);
or U30954 (N_30954,N_30188,N_30257);
and U30955 (N_30955,N_30008,N_30201);
xnor U30956 (N_30956,N_30121,N_30212);
xor U30957 (N_30957,N_30184,N_30291);
and U30958 (N_30958,N_30231,N_30228);
nand U30959 (N_30959,N_30290,N_30268);
xnor U30960 (N_30960,N_30485,N_30266);
nor U30961 (N_30961,N_30253,N_30431);
and U30962 (N_30962,N_30491,N_30188);
xnor U30963 (N_30963,N_30117,N_30405);
nand U30964 (N_30964,N_30360,N_30431);
nand U30965 (N_30965,N_30115,N_30351);
nand U30966 (N_30966,N_30264,N_30207);
and U30967 (N_30967,N_30275,N_30328);
and U30968 (N_30968,N_30303,N_30323);
xor U30969 (N_30969,N_30380,N_30246);
xnor U30970 (N_30970,N_30082,N_30113);
nor U30971 (N_30971,N_30428,N_30092);
or U30972 (N_30972,N_30270,N_30475);
or U30973 (N_30973,N_30266,N_30282);
xnor U30974 (N_30974,N_30335,N_30250);
nand U30975 (N_30975,N_30010,N_30387);
nor U30976 (N_30976,N_30488,N_30340);
or U30977 (N_30977,N_30209,N_30061);
or U30978 (N_30978,N_30039,N_30099);
and U30979 (N_30979,N_30415,N_30310);
xor U30980 (N_30980,N_30332,N_30447);
nand U30981 (N_30981,N_30087,N_30052);
nand U30982 (N_30982,N_30185,N_30155);
nand U30983 (N_30983,N_30428,N_30258);
or U30984 (N_30984,N_30341,N_30365);
xor U30985 (N_30985,N_30011,N_30144);
and U30986 (N_30986,N_30244,N_30199);
nor U30987 (N_30987,N_30383,N_30233);
nand U30988 (N_30988,N_30027,N_30499);
nand U30989 (N_30989,N_30031,N_30085);
xor U30990 (N_30990,N_30173,N_30180);
nand U30991 (N_30991,N_30407,N_30387);
and U30992 (N_30992,N_30304,N_30391);
or U30993 (N_30993,N_30497,N_30442);
nand U30994 (N_30994,N_30220,N_30122);
nand U30995 (N_30995,N_30171,N_30053);
nand U30996 (N_30996,N_30255,N_30388);
nand U30997 (N_30997,N_30121,N_30464);
nor U30998 (N_30998,N_30214,N_30262);
xnor U30999 (N_30999,N_30173,N_30124);
xor U31000 (N_31000,N_30570,N_30974);
nand U31001 (N_31001,N_30559,N_30923);
and U31002 (N_31002,N_30549,N_30599);
and U31003 (N_31003,N_30536,N_30734);
nand U31004 (N_31004,N_30689,N_30768);
nor U31005 (N_31005,N_30504,N_30997);
nor U31006 (N_31006,N_30982,N_30968);
nor U31007 (N_31007,N_30830,N_30765);
xor U31008 (N_31008,N_30674,N_30732);
and U31009 (N_31009,N_30616,N_30727);
or U31010 (N_31010,N_30591,N_30722);
or U31011 (N_31011,N_30720,N_30726);
xnor U31012 (N_31012,N_30645,N_30524);
xnor U31013 (N_31013,N_30764,N_30541);
nand U31014 (N_31014,N_30603,N_30613);
nand U31015 (N_31015,N_30823,N_30756);
and U31016 (N_31016,N_30833,N_30539);
nand U31017 (N_31017,N_30803,N_30593);
nand U31018 (N_31018,N_30635,N_30902);
or U31019 (N_31019,N_30828,N_30790);
or U31020 (N_31020,N_30670,N_30943);
xor U31021 (N_31021,N_30681,N_30761);
or U31022 (N_31022,N_30912,N_30954);
or U31023 (N_31023,N_30522,N_30839);
xnor U31024 (N_31024,N_30711,N_30975);
xor U31025 (N_31025,N_30994,N_30957);
xor U31026 (N_31026,N_30944,N_30762);
and U31027 (N_31027,N_30696,N_30852);
nand U31028 (N_31028,N_30614,N_30820);
xnor U31029 (N_31029,N_30985,N_30791);
nand U31030 (N_31030,N_30700,N_30573);
xor U31031 (N_31031,N_30905,N_30901);
nand U31032 (N_31032,N_30889,N_30742);
or U31033 (N_31033,N_30855,N_30684);
and U31034 (N_31034,N_30740,N_30775);
or U31035 (N_31035,N_30962,N_30723);
nor U31036 (N_31036,N_30940,N_30825);
and U31037 (N_31037,N_30891,N_30597);
xor U31038 (N_31038,N_30648,N_30995);
and U31039 (N_31039,N_30562,N_30611);
and U31040 (N_31040,N_30637,N_30675);
and U31041 (N_31041,N_30904,N_30717);
nand U31042 (N_31042,N_30697,N_30777);
nand U31043 (N_31043,N_30942,N_30592);
or U31044 (N_31044,N_30622,N_30744);
xnor U31045 (N_31045,N_30837,N_30709);
xor U31046 (N_31046,N_30693,N_30881);
or U31047 (N_31047,N_30518,N_30773);
nor U31048 (N_31048,N_30511,N_30920);
or U31049 (N_31049,N_30890,N_30529);
nor U31050 (N_31050,N_30626,N_30565);
or U31051 (N_31051,N_30770,N_30757);
nand U31052 (N_31052,N_30991,N_30615);
and U31053 (N_31053,N_30772,N_30908);
nand U31054 (N_31054,N_30651,N_30575);
xnor U31055 (N_31055,N_30832,N_30763);
nor U31056 (N_31056,N_30784,N_30937);
nand U31057 (N_31057,N_30953,N_30785);
nor U31058 (N_31058,N_30682,N_30864);
xor U31059 (N_31059,N_30643,N_30745);
nand U31060 (N_31060,N_30896,N_30551);
nor U31061 (N_31061,N_30640,N_30818);
xnor U31062 (N_31062,N_30922,N_30862);
nand U31063 (N_31063,N_30600,N_30548);
and U31064 (N_31064,N_30941,N_30503);
nand U31065 (N_31065,N_30581,N_30660);
or U31066 (N_31066,N_30885,N_30679);
or U31067 (N_31067,N_30736,N_30574);
nor U31068 (N_31068,N_30703,N_30911);
or U31069 (N_31069,N_30786,N_30808);
or U31070 (N_31070,N_30520,N_30986);
and U31071 (N_31071,N_30633,N_30984);
and U31072 (N_31072,N_30708,N_30882);
nor U31073 (N_31073,N_30654,N_30620);
nand U31074 (N_31074,N_30850,N_30535);
xnor U31075 (N_31075,N_30624,N_30866);
nand U31076 (N_31076,N_30959,N_30743);
xor U31077 (N_31077,N_30979,N_30571);
or U31078 (N_31078,N_30945,N_30560);
and U31079 (N_31079,N_30563,N_30630);
xnor U31080 (N_31080,N_30605,N_30827);
or U31081 (N_31081,N_30809,N_30967);
or U31082 (N_31082,N_30609,N_30965);
and U31083 (N_31083,N_30956,N_30795);
nor U31084 (N_31084,N_30884,N_30917);
nand U31085 (N_31085,N_30646,N_30678);
xnor U31086 (N_31086,N_30586,N_30787);
nor U31087 (N_31087,N_30776,N_30733);
and U31088 (N_31088,N_30576,N_30702);
nor U31089 (N_31089,N_30993,N_30596);
nor U31090 (N_31090,N_30972,N_30558);
nand U31091 (N_31091,N_30999,N_30612);
or U31092 (N_31092,N_30952,N_30841);
nand U31093 (N_31093,N_30686,N_30750);
xnor U31094 (N_31094,N_30934,N_30590);
xnor U31095 (N_31095,N_30948,N_30706);
and U31096 (N_31096,N_30582,N_30634);
xnor U31097 (N_31097,N_30883,N_30564);
and U31098 (N_31098,N_30928,N_30771);
or U31099 (N_31099,N_30521,N_30567);
nand U31100 (N_31100,N_30871,N_30751);
nand U31101 (N_31101,N_30836,N_30666);
and U31102 (N_31102,N_30794,N_30780);
or U31103 (N_31103,N_30816,N_30960);
or U31104 (N_31104,N_30545,N_30936);
and U31105 (N_31105,N_30653,N_30664);
nand U31106 (N_31106,N_30519,N_30533);
or U31107 (N_31107,N_30888,N_30919);
nor U31108 (N_31108,N_30505,N_30766);
nor U31109 (N_31109,N_30628,N_30623);
nor U31110 (N_31110,N_30621,N_30625);
xnor U31111 (N_31111,N_30918,N_30588);
and U31112 (N_31112,N_30716,N_30749);
or U31113 (N_31113,N_30741,N_30969);
and U31114 (N_31114,N_30644,N_30608);
nor U31115 (N_31115,N_30528,N_30699);
and U31116 (N_31116,N_30859,N_30935);
and U31117 (N_31117,N_30981,N_30792);
xor U31118 (N_31118,N_30851,N_30789);
nand U31119 (N_31119,N_30817,N_30510);
nor U31120 (N_31120,N_30739,N_30556);
or U31121 (N_31121,N_30758,N_30577);
nand U31122 (N_31122,N_30854,N_30691);
nor U31123 (N_31123,N_30754,N_30983);
and U31124 (N_31124,N_30602,N_30829);
nor U31125 (N_31125,N_30879,N_30755);
and U31126 (N_31126,N_30887,N_30595);
nand U31127 (N_31127,N_30970,N_30725);
and U31128 (N_31128,N_30822,N_30638);
xor U31129 (N_31129,N_30729,N_30857);
or U31130 (N_31130,N_30641,N_30987);
xnor U31131 (N_31131,N_30988,N_30894);
nand U31132 (N_31132,N_30710,N_30821);
xnor U31133 (N_31133,N_30868,N_30973);
and U31134 (N_31134,N_30719,N_30671);
or U31135 (N_31135,N_30667,N_30844);
nand U31136 (N_31136,N_30966,N_30655);
xor U31137 (N_31137,N_30712,N_30998);
nand U31138 (N_31138,N_30523,N_30869);
xnor U31139 (N_31139,N_30826,N_30589);
nand U31140 (N_31140,N_30811,N_30788);
and U31141 (N_31141,N_30730,N_30840);
xnor U31142 (N_31142,N_30753,N_30517);
or U31143 (N_31143,N_30799,N_30931);
xnor U31144 (N_31144,N_30698,N_30673);
nor U31145 (N_31145,N_30873,N_30815);
and U31146 (N_31146,N_30713,N_30735);
nand U31147 (N_31147,N_30662,N_30752);
and U31148 (N_31148,N_30793,N_30961);
or U31149 (N_31149,N_30661,N_30507);
xnor U31150 (N_31150,N_30915,N_30618);
or U31151 (N_31151,N_30876,N_30508);
xnor U31152 (N_31152,N_30796,N_30632);
and U31153 (N_31153,N_30627,N_30715);
xnor U31154 (N_31154,N_30909,N_30658);
nand U31155 (N_31155,N_30701,N_30685);
xnor U31156 (N_31156,N_30619,N_30669);
xnor U31157 (N_31157,N_30601,N_30977);
nor U31158 (N_31158,N_30865,N_30527);
nor U31159 (N_31159,N_30897,N_30668);
and U31160 (N_31160,N_30561,N_30672);
nand U31161 (N_31161,N_30950,N_30695);
nand U31162 (N_31162,N_30949,N_30933);
xnor U31163 (N_31163,N_30677,N_30604);
nor U31164 (N_31164,N_30812,N_30579);
nor U31165 (N_31165,N_30705,N_30939);
nor U31166 (N_31166,N_30946,N_30834);
or U31167 (N_31167,N_30683,N_30810);
xor U31168 (N_31168,N_30848,N_30797);
and U31169 (N_31169,N_30578,N_30500);
nand U31170 (N_31170,N_30747,N_30778);
or U31171 (N_31171,N_30926,N_30930);
xor U31172 (N_31172,N_30584,N_30553);
xnor U31173 (N_31173,N_30886,N_30783);
and U31174 (N_31174,N_30870,N_30801);
nand U31175 (N_31175,N_30652,N_30631);
or U31176 (N_31176,N_30831,N_30858);
nand U31177 (N_31177,N_30774,N_30714);
or U31178 (N_31178,N_30537,N_30629);
or U31179 (N_31179,N_30921,N_30639);
or U31180 (N_31180,N_30585,N_30779);
nor U31181 (N_31181,N_30587,N_30849);
nor U31182 (N_31182,N_30552,N_30824);
nand U31183 (N_31183,N_30538,N_30769);
and U31184 (N_31184,N_30996,N_30512);
nand U31185 (N_31185,N_30867,N_30690);
nand U31186 (N_31186,N_30963,N_30814);
nand U31187 (N_31187,N_30929,N_30924);
xor U31188 (N_31188,N_30557,N_30805);
xnor U31189 (N_31189,N_30903,N_30976);
xnor U31190 (N_31190,N_30636,N_30525);
xor U31191 (N_31191,N_30748,N_30760);
and U31192 (N_31192,N_30704,N_30721);
nor U31193 (N_31193,N_30707,N_30980);
nor U31194 (N_31194,N_30899,N_30737);
nand U31195 (N_31195,N_30532,N_30759);
xor U31196 (N_31196,N_30514,N_30663);
or U31197 (N_31197,N_30798,N_30544);
xor U31198 (N_31198,N_30680,N_30880);
xor U31199 (N_31199,N_30893,N_30800);
and U31200 (N_31200,N_30835,N_30842);
xor U31201 (N_31201,N_30746,N_30513);
nand U31202 (N_31202,N_30555,N_30501);
nand U31203 (N_31203,N_30878,N_30568);
xnor U31204 (N_31204,N_30877,N_30958);
or U31205 (N_31205,N_30971,N_30906);
or U31206 (N_31206,N_30892,N_30566);
xor U31207 (N_31207,N_30978,N_30860);
and U31208 (N_31208,N_30895,N_30688);
nor U31209 (N_31209,N_30992,N_30659);
or U31210 (N_31210,N_30516,N_30606);
nand U31211 (N_31211,N_30509,N_30718);
and U31212 (N_31212,N_30657,N_30990);
nor U31213 (N_31213,N_30910,N_30863);
nand U31214 (N_31214,N_30534,N_30951);
nand U31215 (N_31215,N_30838,N_30898);
nor U31216 (N_31216,N_30728,N_30649);
xor U31217 (N_31217,N_30650,N_30554);
or U31218 (N_31218,N_30531,N_30767);
nand U31219 (N_31219,N_30676,N_30914);
nand U31220 (N_31220,N_30583,N_30819);
and U31221 (N_31221,N_30647,N_30506);
or U31222 (N_31222,N_30550,N_30547);
or U31223 (N_31223,N_30542,N_30925);
and U31224 (N_31224,N_30964,N_30913);
xor U31225 (N_31225,N_30806,N_30802);
xnor U31226 (N_31226,N_30502,N_30853);
or U31227 (N_31227,N_30813,N_30846);
and U31228 (N_31228,N_30569,N_30738);
and U31229 (N_31229,N_30874,N_30665);
xnor U31230 (N_31230,N_30932,N_30916);
xnor U31231 (N_31231,N_30781,N_30656);
or U31232 (N_31232,N_30847,N_30938);
xnor U31233 (N_31233,N_30875,N_30856);
and U31234 (N_31234,N_30580,N_30540);
nor U31235 (N_31235,N_30607,N_30861);
and U31236 (N_31236,N_30947,N_30543);
nor U31237 (N_31237,N_30804,N_30843);
nor U31238 (N_31238,N_30900,N_30515);
nor U31239 (N_31239,N_30807,N_30598);
and U31240 (N_31240,N_30594,N_30694);
nand U31241 (N_31241,N_30872,N_30642);
or U31242 (N_31242,N_30572,N_30989);
nand U31243 (N_31243,N_30687,N_30692);
and U31244 (N_31244,N_30617,N_30907);
or U31245 (N_31245,N_30546,N_30955);
or U31246 (N_31246,N_30526,N_30610);
nand U31247 (N_31247,N_30724,N_30845);
xnor U31248 (N_31248,N_30927,N_30782);
or U31249 (N_31249,N_30530,N_30731);
or U31250 (N_31250,N_30832,N_30526);
and U31251 (N_31251,N_30517,N_30901);
xor U31252 (N_31252,N_30850,N_30601);
nand U31253 (N_31253,N_30866,N_30787);
nor U31254 (N_31254,N_30527,N_30931);
and U31255 (N_31255,N_30821,N_30675);
and U31256 (N_31256,N_30562,N_30586);
xor U31257 (N_31257,N_30746,N_30564);
nor U31258 (N_31258,N_30814,N_30629);
nand U31259 (N_31259,N_30767,N_30949);
xnor U31260 (N_31260,N_30973,N_30729);
nor U31261 (N_31261,N_30891,N_30543);
nor U31262 (N_31262,N_30680,N_30525);
and U31263 (N_31263,N_30546,N_30994);
and U31264 (N_31264,N_30512,N_30883);
xnor U31265 (N_31265,N_30830,N_30968);
nor U31266 (N_31266,N_30727,N_30957);
nand U31267 (N_31267,N_30752,N_30660);
or U31268 (N_31268,N_30536,N_30568);
nand U31269 (N_31269,N_30864,N_30782);
and U31270 (N_31270,N_30921,N_30668);
nand U31271 (N_31271,N_30780,N_30782);
and U31272 (N_31272,N_30529,N_30703);
or U31273 (N_31273,N_30698,N_30755);
xnor U31274 (N_31274,N_30677,N_30879);
xnor U31275 (N_31275,N_30502,N_30936);
nand U31276 (N_31276,N_30673,N_30928);
xnor U31277 (N_31277,N_30861,N_30664);
or U31278 (N_31278,N_30571,N_30996);
xnor U31279 (N_31279,N_30824,N_30598);
or U31280 (N_31280,N_30508,N_30756);
xor U31281 (N_31281,N_30956,N_30661);
or U31282 (N_31282,N_30997,N_30640);
xor U31283 (N_31283,N_30703,N_30746);
xnor U31284 (N_31284,N_30550,N_30603);
nor U31285 (N_31285,N_30890,N_30666);
nor U31286 (N_31286,N_30619,N_30697);
and U31287 (N_31287,N_30538,N_30681);
nand U31288 (N_31288,N_30610,N_30806);
xnor U31289 (N_31289,N_30531,N_30848);
nor U31290 (N_31290,N_30667,N_30859);
xor U31291 (N_31291,N_30646,N_30624);
nand U31292 (N_31292,N_30883,N_30624);
xor U31293 (N_31293,N_30786,N_30662);
or U31294 (N_31294,N_30765,N_30941);
nor U31295 (N_31295,N_30523,N_30882);
or U31296 (N_31296,N_30768,N_30609);
or U31297 (N_31297,N_30538,N_30632);
or U31298 (N_31298,N_30773,N_30743);
nor U31299 (N_31299,N_30891,N_30880);
nor U31300 (N_31300,N_30697,N_30971);
or U31301 (N_31301,N_30782,N_30920);
or U31302 (N_31302,N_30870,N_30680);
xnor U31303 (N_31303,N_30992,N_30855);
nand U31304 (N_31304,N_30791,N_30908);
nand U31305 (N_31305,N_30771,N_30548);
and U31306 (N_31306,N_30578,N_30706);
nor U31307 (N_31307,N_30674,N_30951);
or U31308 (N_31308,N_30936,N_30848);
xnor U31309 (N_31309,N_30665,N_30772);
nand U31310 (N_31310,N_30704,N_30595);
or U31311 (N_31311,N_30716,N_30520);
and U31312 (N_31312,N_30718,N_30839);
nor U31313 (N_31313,N_30688,N_30702);
nor U31314 (N_31314,N_30566,N_30888);
xnor U31315 (N_31315,N_30902,N_30679);
or U31316 (N_31316,N_30594,N_30615);
and U31317 (N_31317,N_30649,N_30920);
nand U31318 (N_31318,N_30960,N_30508);
nor U31319 (N_31319,N_30998,N_30693);
nor U31320 (N_31320,N_30822,N_30666);
or U31321 (N_31321,N_30761,N_30585);
or U31322 (N_31322,N_30865,N_30656);
nand U31323 (N_31323,N_30584,N_30772);
and U31324 (N_31324,N_30537,N_30691);
and U31325 (N_31325,N_30769,N_30589);
nor U31326 (N_31326,N_30549,N_30813);
xnor U31327 (N_31327,N_30540,N_30636);
and U31328 (N_31328,N_30759,N_30977);
xnor U31329 (N_31329,N_30534,N_30637);
and U31330 (N_31330,N_30902,N_30664);
nand U31331 (N_31331,N_30650,N_30728);
nand U31332 (N_31332,N_30939,N_30906);
and U31333 (N_31333,N_30824,N_30569);
nand U31334 (N_31334,N_30661,N_30882);
xnor U31335 (N_31335,N_30580,N_30763);
or U31336 (N_31336,N_30741,N_30815);
nor U31337 (N_31337,N_30668,N_30846);
or U31338 (N_31338,N_30817,N_30598);
and U31339 (N_31339,N_30861,N_30554);
nor U31340 (N_31340,N_30562,N_30977);
nor U31341 (N_31341,N_30825,N_30762);
nor U31342 (N_31342,N_30714,N_30884);
xor U31343 (N_31343,N_30678,N_30983);
xnor U31344 (N_31344,N_30949,N_30754);
and U31345 (N_31345,N_30903,N_30640);
and U31346 (N_31346,N_30817,N_30918);
or U31347 (N_31347,N_30723,N_30718);
nand U31348 (N_31348,N_30536,N_30562);
or U31349 (N_31349,N_30867,N_30623);
nor U31350 (N_31350,N_30872,N_30662);
nor U31351 (N_31351,N_30729,N_30711);
nor U31352 (N_31352,N_30871,N_30675);
and U31353 (N_31353,N_30537,N_30545);
xor U31354 (N_31354,N_30589,N_30793);
nand U31355 (N_31355,N_30654,N_30802);
nand U31356 (N_31356,N_30526,N_30638);
xor U31357 (N_31357,N_30849,N_30956);
nand U31358 (N_31358,N_30548,N_30706);
xnor U31359 (N_31359,N_30694,N_30531);
and U31360 (N_31360,N_30588,N_30874);
xor U31361 (N_31361,N_30820,N_30510);
xnor U31362 (N_31362,N_30688,N_30753);
nor U31363 (N_31363,N_30647,N_30629);
nor U31364 (N_31364,N_30534,N_30529);
nand U31365 (N_31365,N_30737,N_30642);
nand U31366 (N_31366,N_30611,N_30833);
and U31367 (N_31367,N_30642,N_30591);
nand U31368 (N_31368,N_30879,N_30618);
nor U31369 (N_31369,N_30901,N_30760);
nand U31370 (N_31370,N_30705,N_30747);
nor U31371 (N_31371,N_30781,N_30621);
or U31372 (N_31372,N_30943,N_30583);
nand U31373 (N_31373,N_30615,N_30825);
and U31374 (N_31374,N_30834,N_30844);
and U31375 (N_31375,N_30992,N_30984);
or U31376 (N_31376,N_30508,N_30765);
nand U31377 (N_31377,N_30783,N_30541);
nor U31378 (N_31378,N_30719,N_30669);
or U31379 (N_31379,N_30501,N_30558);
and U31380 (N_31380,N_30964,N_30901);
nand U31381 (N_31381,N_30558,N_30844);
nor U31382 (N_31382,N_30890,N_30889);
or U31383 (N_31383,N_30557,N_30653);
nand U31384 (N_31384,N_30803,N_30963);
and U31385 (N_31385,N_30846,N_30736);
and U31386 (N_31386,N_30504,N_30954);
xor U31387 (N_31387,N_30645,N_30754);
nand U31388 (N_31388,N_30890,N_30689);
nand U31389 (N_31389,N_30850,N_30948);
and U31390 (N_31390,N_30740,N_30967);
xnor U31391 (N_31391,N_30907,N_30954);
or U31392 (N_31392,N_30866,N_30612);
and U31393 (N_31393,N_30905,N_30878);
or U31394 (N_31394,N_30666,N_30598);
xor U31395 (N_31395,N_30534,N_30644);
and U31396 (N_31396,N_30634,N_30825);
nor U31397 (N_31397,N_30979,N_30937);
nor U31398 (N_31398,N_30758,N_30986);
or U31399 (N_31399,N_30617,N_30775);
and U31400 (N_31400,N_30717,N_30528);
and U31401 (N_31401,N_30601,N_30701);
or U31402 (N_31402,N_30503,N_30849);
nand U31403 (N_31403,N_30546,N_30579);
nor U31404 (N_31404,N_30869,N_30722);
nor U31405 (N_31405,N_30847,N_30708);
or U31406 (N_31406,N_30906,N_30970);
nor U31407 (N_31407,N_30858,N_30780);
xnor U31408 (N_31408,N_30611,N_30544);
nor U31409 (N_31409,N_30647,N_30945);
and U31410 (N_31410,N_30898,N_30853);
xnor U31411 (N_31411,N_30570,N_30529);
and U31412 (N_31412,N_30983,N_30656);
nand U31413 (N_31413,N_30777,N_30742);
nor U31414 (N_31414,N_30919,N_30895);
xor U31415 (N_31415,N_30691,N_30695);
and U31416 (N_31416,N_30950,N_30789);
or U31417 (N_31417,N_30995,N_30899);
or U31418 (N_31418,N_30547,N_30688);
nand U31419 (N_31419,N_30878,N_30740);
or U31420 (N_31420,N_30623,N_30610);
nand U31421 (N_31421,N_30591,N_30954);
or U31422 (N_31422,N_30716,N_30695);
or U31423 (N_31423,N_30665,N_30959);
nand U31424 (N_31424,N_30553,N_30810);
xor U31425 (N_31425,N_30777,N_30891);
xnor U31426 (N_31426,N_30581,N_30810);
xnor U31427 (N_31427,N_30732,N_30856);
xor U31428 (N_31428,N_30737,N_30589);
nand U31429 (N_31429,N_30971,N_30849);
nor U31430 (N_31430,N_30645,N_30793);
nor U31431 (N_31431,N_30824,N_30826);
nand U31432 (N_31432,N_30681,N_30528);
or U31433 (N_31433,N_30512,N_30679);
nor U31434 (N_31434,N_30506,N_30714);
or U31435 (N_31435,N_30869,N_30585);
xor U31436 (N_31436,N_30714,N_30960);
and U31437 (N_31437,N_30631,N_30851);
or U31438 (N_31438,N_30692,N_30530);
or U31439 (N_31439,N_30522,N_30740);
nand U31440 (N_31440,N_30803,N_30757);
xnor U31441 (N_31441,N_30579,N_30500);
or U31442 (N_31442,N_30820,N_30537);
or U31443 (N_31443,N_30791,N_30526);
and U31444 (N_31444,N_30949,N_30836);
nor U31445 (N_31445,N_30675,N_30619);
and U31446 (N_31446,N_30802,N_30777);
nand U31447 (N_31447,N_30851,N_30792);
xor U31448 (N_31448,N_30955,N_30993);
nand U31449 (N_31449,N_30647,N_30560);
and U31450 (N_31450,N_30690,N_30620);
or U31451 (N_31451,N_30799,N_30976);
or U31452 (N_31452,N_30909,N_30791);
nor U31453 (N_31453,N_30654,N_30854);
and U31454 (N_31454,N_30656,N_30968);
xor U31455 (N_31455,N_30681,N_30592);
nand U31456 (N_31456,N_30626,N_30702);
nor U31457 (N_31457,N_30562,N_30982);
nor U31458 (N_31458,N_30775,N_30796);
or U31459 (N_31459,N_30988,N_30821);
and U31460 (N_31460,N_30575,N_30671);
nand U31461 (N_31461,N_30541,N_30777);
or U31462 (N_31462,N_30830,N_30931);
nor U31463 (N_31463,N_30797,N_30641);
and U31464 (N_31464,N_30754,N_30575);
or U31465 (N_31465,N_30923,N_30619);
and U31466 (N_31466,N_30701,N_30993);
nand U31467 (N_31467,N_30686,N_30500);
nand U31468 (N_31468,N_30674,N_30856);
and U31469 (N_31469,N_30866,N_30752);
xor U31470 (N_31470,N_30912,N_30898);
xor U31471 (N_31471,N_30600,N_30657);
xor U31472 (N_31472,N_30704,N_30956);
xor U31473 (N_31473,N_30577,N_30781);
or U31474 (N_31474,N_30948,N_30765);
or U31475 (N_31475,N_30568,N_30794);
nand U31476 (N_31476,N_30677,N_30883);
nor U31477 (N_31477,N_30642,N_30528);
nor U31478 (N_31478,N_30635,N_30892);
nand U31479 (N_31479,N_30894,N_30933);
or U31480 (N_31480,N_30560,N_30671);
nor U31481 (N_31481,N_30631,N_30532);
or U31482 (N_31482,N_30927,N_30806);
and U31483 (N_31483,N_30962,N_30865);
or U31484 (N_31484,N_30768,N_30998);
nor U31485 (N_31485,N_30757,N_30880);
and U31486 (N_31486,N_30761,N_30866);
or U31487 (N_31487,N_30946,N_30527);
nor U31488 (N_31488,N_30777,N_30790);
xnor U31489 (N_31489,N_30562,N_30937);
or U31490 (N_31490,N_30549,N_30943);
or U31491 (N_31491,N_30991,N_30742);
xor U31492 (N_31492,N_30797,N_30631);
and U31493 (N_31493,N_30914,N_30552);
nand U31494 (N_31494,N_30724,N_30582);
and U31495 (N_31495,N_30862,N_30506);
nand U31496 (N_31496,N_30890,N_30756);
nand U31497 (N_31497,N_30620,N_30947);
or U31498 (N_31498,N_30945,N_30554);
or U31499 (N_31499,N_30812,N_30714);
xnor U31500 (N_31500,N_31210,N_31137);
nor U31501 (N_31501,N_31268,N_31220);
and U31502 (N_31502,N_31190,N_31253);
nand U31503 (N_31503,N_31313,N_31192);
nor U31504 (N_31504,N_31219,N_31301);
nand U31505 (N_31505,N_31425,N_31150);
xnor U31506 (N_31506,N_31432,N_31485);
or U31507 (N_31507,N_31047,N_31168);
xnor U31508 (N_31508,N_31354,N_31246);
xor U31509 (N_31509,N_31453,N_31142);
xor U31510 (N_31510,N_31036,N_31351);
nand U31511 (N_31511,N_31228,N_31067);
and U31512 (N_31512,N_31431,N_31125);
or U31513 (N_31513,N_31325,N_31381);
xnor U31514 (N_31514,N_31378,N_31048);
xor U31515 (N_31515,N_31202,N_31315);
and U31516 (N_31516,N_31327,N_31018);
xor U31517 (N_31517,N_31127,N_31222);
nor U31518 (N_31518,N_31306,N_31387);
nand U31519 (N_31519,N_31177,N_31410);
nand U31520 (N_31520,N_31011,N_31349);
nand U31521 (N_31521,N_31272,N_31195);
nand U31522 (N_31522,N_31469,N_31424);
nor U31523 (N_31523,N_31496,N_31476);
and U31524 (N_31524,N_31462,N_31377);
nand U31525 (N_31525,N_31383,N_31136);
xor U31526 (N_31526,N_31474,N_31198);
xnor U31527 (N_31527,N_31110,N_31356);
or U31528 (N_31528,N_31031,N_31010);
nor U31529 (N_31529,N_31433,N_31045);
and U31530 (N_31530,N_31115,N_31174);
xor U31531 (N_31531,N_31131,N_31412);
and U31532 (N_31532,N_31364,N_31188);
nand U31533 (N_31533,N_31266,N_31418);
nor U31534 (N_31534,N_31012,N_31102);
and U31535 (N_31535,N_31229,N_31014);
and U31536 (N_31536,N_31173,N_31430);
or U31537 (N_31537,N_31186,N_31061);
and U31538 (N_31538,N_31120,N_31434);
nor U31539 (N_31539,N_31256,N_31106);
xnor U31540 (N_31540,N_31399,N_31237);
nor U31541 (N_31541,N_31450,N_31487);
nor U31542 (N_31542,N_31429,N_31024);
or U31543 (N_31543,N_31322,N_31262);
and U31544 (N_31544,N_31078,N_31232);
nor U31545 (N_31545,N_31282,N_31263);
nand U31546 (N_31546,N_31160,N_31300);
and U31547 (N_31547,N_31352,N_31422);
nand U31548 (N_31548,N_31339,N_31231);
and U31549 (N_31549,N_31404,N_31182);
xnor U31550 (N_31550,N_31307,N_31426);
or U31551 (N_31551,N_31440,N_31119);
nor U31552 (N_31552,N_31355,N_31209);
xor U31553 (N_31553,N_31112,N_31166);
xnor U31554 (N_31554,N_31050,N_31278);
or U31555 (N_31555,N_31075,N_31326);
xor U31556 (N_31556,N_31242,N_31408);
or U31557 (N_31557,N_31324,N_31259);
nor U31558 (N_31558,N_31459,N_31403);
nor U31559 (N_31559,N_31206,N_31118);
xnor U31560 (N_31560,N_31214,N_31309);
nand U31561 (N_31561,N_31489,N_31104);
nor U31562 (N_31562,N_31499,N_31235);
nand U31563 (N_31563,N_31409,N_31491);
and U31564 (N_31564,N_31252,N_31191);
xnor U31565 (N_31565,N_31197,N_31490);
nor U31566 (N_31566,N_31271,N_31297);
xor U31567 (N_31567,N_31287,N_31405);
and U31568 (N_31568,N_31091,N_31436);
nand U31569 (N_31569,N_31342,N_31042);
and U31570 (N_31570,N_31157,N_31138);
xor U31571 (N_31571,N_31132,N_31143);
nand U31572 (N_31572,N_31133,N_31420);
xor U31573 (N_31573,N_31054,N_31467);
nor U31574 (N_31574,N_31486,N_31391);
nand U31575 (N_31575,N_31465,N_31402);
xor U31576 (N_31576,N_31261,N_31294);
xor U31577 (N_31577,N_31189,N_31081);
nand U31578 (N_31578,N_31323,N_31006);
nor U31579 (N_31579,N_31396,N_31308);
xnor U31580 (N_31580,N_31480,N_31375);
and U31581 (N_31581,N_31376,N_31265);
nand U31582 (N_31582,N_31251,N_31066);
xor U31583 (N_31583,N_31350,N_31097);
and U31584 (N_31584,N_31318,N_31371);
or U31585 (N_31585,N_31033,N_31034);
and U31586 (N_31586,N_31359,N_31448);
or U31587 (N_31587,N_31084,N_31076);
nor U31588 (N_31588,N_31303,N_31370);
and U31589 (N_31589,N_31362,N_31041);
nand U31590 (N_31590,N_31390,N_31479);
nand U31591 (N_31591,N_31279,N_31395);
xnor U31592 (N_31592,N_31204,N_31095);
nand U31593 (N_31593,N_31105,N_31365);
or U31594 (N_31594,N_31003,N_31407);
nand U31595 (N_31595,N_31338,N_31427);
or U31596 (N_31596,N_31452,N_31464);
nor U31597 (N_31597,N_31181,N_31471);
or U31598 (N_31598,N_31366,N_31329);
nand U31599 (N_31599,N_31072,N_31027);
nor U31600 (N_31600,N_31472,N_31124);
and U31601 (N_31601,N_31037,N_31461);
or U31602 (N_31602,N_31245,N_31099);
nand U31603 (N_31603,N_31281,N_31293);
nand U31604 (N_31604,N_31147,N_31056);
nand U31605 (N_31605,N_31092,N_31164);
or U31606 (N_31606,N_31416,N_31139);
xor U31607 (N_31607,N_31032,N_31217);
and U31608 (N_31608,N_31457,N_31126);
xor U31609 (N_31609,N_31234,N_31015);
nand U31610 (N_31610,N_31473,N_31101);
or U31611 (N_31611,N_31269,N_31247);
nand U31612 (N_31612,N_31270,N_31317);
nor U31613 (N_31613,N_31302,N_31108);
and U31614 (N_31614,N_31064,N_31477);
or U31615 (N_31615,N_31156,N_31392);
and U31616 (N_31616,N_31074,N_31098);
nand U31617 (N_31617,N_31346,N_31154);
nand U31618 (N_31618,N_31211,N_31428);
or U31619 (N_31619,N_31414,N_31347);
or U31620 (N_31620,N_31208,N_31030);
xor U31621 (N_31621,N_31215,N_31152);
and U31622 (N_31622,N_31288,N_31025);
or U31623 (N_31623,N_31069,N_31141);
nand U31624 (N_31624,N_31070,N_31236);
xor U31625 (N_31625,N_31248,N_31004);
or U31626 (N_31626,N_31413,N_31382);
nand U31627 (N_31627,N_31466,N_31226);
and U31628 (N_31628,N_31332,N_31162);
nand U31629 (N_31629,N_31002,N_31176);
nand U31630 (N_31630,N_31135,N_31335);
nand U31631 (N_31631,N_31249,N_31239);
and U31632 (N_31632,N_31344,N_31345);
and U31633 (N_31633,N_31028,N_31212);
nor U31634 (N_31634,N_31216,N_31223);
nand U31635 (N_31635,N_31053,N_31257);
xor U31636 (N_31636,N_31167,N_31320);
nor U31637 (N_31637,N_31494,N_31008);
xor U31638 (N_31638,N_31421,N_31470);
and U31639 (N_31639,N_31123,N_31052);
nor U31640 (N_31640,N_31039,N_31254);
nand U31641 (N_31641,N_31017,N_31079);
xnor U31642 (N_31642,N_31178,N_31170);
or U31643 (N_31643,N_31080,N_31495);
nand U31644 (N_31644,N_31196,N_31085);
nand U31645 (N_31645,N_31063,N_31284);
nor U31646 (N_31646,N_31199,N_31130);
or U31647 (N_31647,N_31417,N_31423);
and U31648 (N_31648,N_31446,N_31264);
nor U31649 (N_31649,N_31291,N_31384);
nor U31650 (N_31650,N_31458,N_31393);
nor U31651 (N_31651,N_31116,N_31273);
nand U31652 (N_31652,N_31140,N_31087);
and U31653 (N_31653,N_31218,N_31488);
xor U31654 (N_31654,N_31155,N_31463);
nand U31655 (N_31655,N_31107,N_31275);
or U31656 (N_31656,N_31337,N_31035);
or U31657 (N_31657,N_31043,N_31029);
nor U31658 (N_31658,N_31333,N_31305);
nand U31659 (N_31659,N_31238,N_31439);
and U31660 (N_31660,N_31055,N_31073);
or U31661 (N_31661,N_31368,N_31314);
nand U31662 (N_31662,N_31086,N_31169);
nand U31663 (N_31663,N_31049,N_31159);
nor U31664 (N_31664,N_31353,N_31059);
nand U31665 (N_31665,N_31482,N_31373);
nand U31666 (N_31666,N_31398,N_31367);
xnor U31667 (N_31667,N_31369,N_31000);
xnor U31668 (N_31668,N_31372,N_31388);
or U31669 (N_31669,N_31447,N_31267);
xor U31670 (N_31670,N_31207,N_31258);
xor U31671 (N_31671,N_31151,N_31013);
nand U31672 (N_31672,N_31437,N_31241);
nand U31673 (N_31673,N_31386,N_31094);
xor U31674 (N_31674,N_31274,N_31401);
or U31675 (N_31675,N_31243,N_31230);
and U31676 (N_31676,N_31451,N_31153);
xor U31677 (N_31677,N_31492,N_31065);
and U31678 (N_31678,N_31148,N_31146);
nand U31679 (N_31679,N_31255,N_31385);
xnor U31680 (N_31680,N_31109,N_31163);
and U31681 (N_31681,N_31497,N_31400);
xnor U31682 (N_31682,N_31319,N_31128);
or U31683 (N_31683,N_31312,N_31158);
nor U31684 (N_31684,N_31244,N_31454);
xnor U31685 (N_31685,N_31062,N_31460);
xor U31686 (N_31686,N_31172,N_31129);
xnor U31687 (N_31687,N_31295,N_31280);
nor U31688 (N_31688,N_31357,N_31225);
and U31689 (N_31689,N_31203,N_31290);
and U31690 (N_31690,N_31213,N_31483);
nand U31691 (N_31691,N_31016,N_31456);
xor U31692 (N_31692,N_31185,N_31304);
nand U31693 (N_31693,N_31082,N_31088);
xor U31694 (N_31694,N_31096,N_31009);
nand U31695 (N_31695,N_31201,N_31227);
xnor U31696 (N_31696,N_31221,N_31090);
or U31697 (N_31697,N_31144,N_31089);
nand U31698 (N_31698,N_31361,N_31276);
or U31699 (N_31699,N_31277,N_31334);
xor U31700 (N_31700,N_31077,N_31071);
or U31701 (N_31701,N_31057,N_31114);
or U31702 (N_31702,N_31493,N_31374);
nand U31703 (N_31703,N_31475,N_31444);
or U31704 (N_31704,N_31449,N_31233);
or U31705 (N_31705,N_31438,N_31184);
nand U31706 (N_31706,N_31468,N_31111);
and U31707 (N_31707,N_31310,N_31283);
xor U31708 (N_31708,N_31358,N_31117);
xor U31709 (N_31709,N_31328,N_31187);
or U31710 (N_31710,N_31060,N_31321);
nand U31711 (N_31711,N_31165,N_31341);
xor U31712 (N_31712,N_31296,N_31193);
or U31713 (N_31713,N_31455,N_31481);
xor U31714 (N_31714,N_31134,N_31478);
or U31715 (N_31715,N_31113,N_31360);
or U31716 (N_31716,N_31442,N_31380);
nor U31717 (N_31717,N_31331,N_31100);
xor U31718 (N_31718,N_31044,N_31046);
xor U31719 (N_31719,N_31415,N_31183);
nand U31720 (N_31720,N_31122,N_31058);
or U31721 (N_31721,N_31498,N_31180);
or U31722 (N_31722,N_31411,N_31224);
nand U31723 (N_31723,N_31161,N_31419);
nor U31724 (N_31724,N_31336,N_31394);
and U31725 (N_31725,N_31260,N_31441);
nand U31726 (N_31726,N_31397,N_31194);
or U31727 (N_31727,N_31007,N_31145);
nor U31728 (N_31728,N_31240,N_31068);
and U31729 (N_31729,N_31250,N_31020);
and U31730 (N_31730,N_31484,N_31363);
or U31731 (N_31731,N_31340,N_31040);
nor U31732 (N_31732,N_31083,N_31026);
nand U31733 (N_31733,N_31389,N_31298);
nor U31734 (N_31734,N_31289,N_31292);
nand U31735 (N_31735,N_31443,N_31286);
or U31736 (N_31736,N_31379,N_31175);
nand U31737 (N_31737,N_31093,N_31435);
xnor U31738 (N_31738,N_31022,N_31445);
nand U31739 (N_31739,N_31200,N_31001);
or U31740 (N_31740,N_31299,N_31316);
and U31741 (N_31741,N_31103,N_31051);
and U31742 (N_31742,N_31330,N_31121);
nor U31743 (N_31743,N_31023,N_31348);
nand U31744 (N_31744,N_31406,N_31019);
or U31745 (N_31745,N_31343,N_31005);
nand U31746 (N_31746,N_31021,N_31038);
xor U31747 (N_31747,N_31179,N_31285);
nand U31748 (N_31748,N_31205,N_31149);
and U31749 (N_31749,N_31171,N_31311);
nand U31750 (N_31750,N_31395,N_31380);
or U31751 (N_31751,N_31022,N_31376);
or U31752 (N_31752,N_31233,N_31322);
nor U31753 (N_31753,N_31270,N_31304);
xnor U31754 (N_31754,N_31011,N_31295);
xnor U31755 (N_31755,N_31460,N_31318);
nor U31756 (N_31756,N_31207,N_31159);
nor U31757 (N_31757,N_31273,N_31344);
or U31758 (N_31758,N_31427,N_31317);
or U31759 (N_31759,N_31233,N_31205);
and U31760 (N_31760,N_31166,N_31248);
and U31761 (N_31761,N_31154,N_31130);
nand U31762 (N_31762,N_31076,N_31003);
or U31763 (N_31763,N_31122,N_31277);
and U31764 (N_31764,N_31379,N_31151);
nor U31765 (N_31765,N_31299,N_31015);
or U31766 (N_31766,N_31309,N_31339);
and U31767 (N_31767,N_31038,N_31117);
and U31768 (N_31768,N_31359,N_31001);
xnor U31769 (N_31769,N_31182,N_31376);
xor U31770 (N_31770,N_31485,N_31147);
and U31771 (N_31771,N_31222,N_31369);
nor U31772 (N_31772,N_31142,N_31290);
and U31773 (N_31773,N_31374,N_31039);
or U31774 (N_31774,N_31053,N_31447);
xor U31775 (N_31775,N_31427,N_31460);
and U31776 (N_31776,N_31266,N_31462);
or U31777 (N_31777,N_31101,N_31456);
nor U31778 (N_31778,N_31150,N_31022);
nor U31779 (N_31779,N_31238,N_31050);
and U31780 (N_31780,N_31402,N_31220);
nor U31781 (N_31781,N_31152,N_31375);
and U31782 (N_31782,N_31276,N_31174);
and U31783 (N_31783,N_31328,N_31022);
or U31784 (N_31784,N_31457,N_31398);
and U31785 (N_31785,N_31094,N_31260);
or U31786 (N_31786,N_31369,N_31034);
or U31787 (N_31787,N_31378,N_31052);
xnor U31788 (N_31788,N_31453,N_31036);
nand U31789 (N_31789,N_31407,N_31178);
nand U31790 (N_31790,N_31280,N_31089);
or U31791 (N_31791,N_31207,N_31160);
nor U31792 (N_31792,N_31053,N_31448);
or U31793 (N_31793,N_31110,N_31497);
nor U31794 (N_31794,N_31462,N_31147);
or U31795 (N_31795,N_31371,N_31274);
xnor U31796 (N_31796,N_31143,N_31255);
xor U31797 (N_31797,N_31226,N_31052);
nor U31798 (N_31798,N_31241,N_31338);
nand U31799 (N_31799,N_31230,N_31456);
xor U31800 (N_31800,N_31445,N_31389);
and U31801 (N_31801,N_31104,N_31422);
and U31802 (N_31802,N_31293,N_31373);
nor U31803 (N_31803,N_31453,N_31126);
and U31804 (N_31804,N_31384,N_31482);
and U31805 (N_31805,N_31495,N_31374);
or U31806 (N_31806,N_31166,N_31168);
or U31807 (N_31807,N_31445,N_31194);
or U31808 (N_31808,N_31231,N_31452);
xnor U31809 (N_31809,N_31155,N_31012);
nand U31810 (N_31810,N_31208,N_31056);
and U31811 (N_31811,N_31306,N_31272);
xnor U31812 (N_31812,N_31123,N_31159);
xnor U31813 (N_31813,N_31443,N_31192);
nand U31814 (N_31814,N_31158,N_31291);
nand U31815 (N_31815,N_31049,N_31202);
or U31816 (N_31816,N_31166,N_31303);
nor U31817 (N_31817,N_31081,N_31071);
xnor U31818 (N_31818,N_31405,N_31107);
xnor U31819 (N_31819,N_31117,N_31468);
and U31820 (N_31820,N_31422,N_31426);
xor U31821 (N_31821,N_31126,N_31367);
nor U31822 (N_31822,N_31477,N_31126);
or U31823 (N_31823,N_31192,N_31123);
nand U31824 (N_31824,N_31235,N_31378);
nor U31825 (N_31825,N_31220,N_31099);
or U31826 (N_31826,N_31442,N_31131);
xnor U31827 (N_31827,N_31451,N_31189);
nor U31828 (N_31828,N_31460,N_31395);
nor U31829 (N_31829,N_31381,N_31362);
or U31830 (N_31830,N_31101,N_31111);
xnor U31831 (N_31831,N_31415,N_31095);
xnor U31832 (N_31832,N_31057,N_31471);
nand U31833 (N_31833,N_31141,N_31034);
and U31834 (N_31834,N_31314,N_31311);
nand U31835 (N_31835,N_31468,N_31019);
and U31836 (N_31836,N_31313,N_31152);
xnor U31837 (N_31837,N_31222,N_31364);
and U31838 (N_31838,N_31338,N_31102);
and U31839 (N_31839,N_31214,N_31191);
nand U31840 (N_31840,N_31087,N_31124);
or U31841 (N_31841,N_31029,N_31416);
nor U31842 (N_31842,N_31277,N_31430);
and U31843 (N_31843,N_31376,N_31038);
xnor U31844 (N_31844,N_31170,N_31452);
xor U31845 (N_31845,N_31144,N_31340);
or U31846 (N_31846,N_31179,N_31168);
xor U31847 (N_31847,N_31324,N_31085);
nand U31848 (N_31848,N_31274,N_31033);
and U31849 (N_31849,N_31013,N_31263);
and U31850 (N_31850,N_31253,N_31427);
xnor U31851 (N_31851,N_31128,N_31285);
and U31852 (N_31852,N_31370,N_31019);
or U31853 (N_31853,N_31267,N_31152);
nand U31854 (N_31854,N_31301,N_31302);
nand U31855 (N_31855,N_31412,N_31289);
and U31856 (N_31856,N_31457,N_31323);
nor U31857 (N_31857,N_31246,N_31009);
and U31858 (N_31858,N_31359,N_31273);
nor U31859 (N_31859,N_31357,N_31052);
nand U31860 (N_31860,N_31347,N_31443);
and U31861 (N_31861,N_31245,N_31345);
nand U31862 (N_31862,N_31012,N_31174);
nor U31863 (N_31863,N_31435,N_31136);
and U31864 (N_31864,N_31279,N_31104);
xnor U31865 (N_31865,N_31486,N_31207);
and U31866 (N_31866,N_31099,N_31345);
or U31867 (N_31867,N_31349,N_31002);
and U31868 (N_31868,N_31408,N_31048);
and U31869 (N_31869,N_31063,N_31050);
or U31870 (N_31870,N_31326,N_31263);
xor U31871 (N_31871,N_31259,N_31263);
nand U31872 (N_31872,N_31022,N_31087);
nand U31873 (N_31873,N_31102,N_31121);
or U31874 (N_31874,N_31431,N_31231);
nand U31875 (N_31875,N_31299,N_31251);
or U31876 (N_31876,N_31228,N_31289);
or U31877 (N_31877,N_31032,N_31143);
and U31878 (N_31878,N_31376,N_31037);
nand U31879 (N_31879,N_31314,N_31427);
and U31880 (N_31880,N_31249,N_31129);
xnor U31881 (N_31881,N_31245,N_31457);
xnor U31882 (N_31882,N_31239,N_31213);
and U31883 (N_31883,N_31043,N_31233);
nand U31884 (N_31884,N_31442,N_31460);
xnor U31885 (N_31885,N_31253,N_31205);
and U31886 (N_31886,N_31473,N_31278);
xnor U31887 (N_31887,N_31004,N_31443);
xor U31888 (N_31888,N_31350,N_31034);
nor U31889 (N_31889,N_31474,N_31410);
and U31890 (N_31890,N_31191,N_31329);
and U31891 (N_31891,N_31024,N_31433);
nor U31892 (N_31892,N_31062,N_31212);
and U31893 (N_31893,N_31354,N_31346);
and U31894 (N_31894,N_31482,N_31281);
nand U31895 (N_31895,N_31040,N_31399);
or U31896 (N_31896,N_31193,N_31079);
and U31897 (N_31897,N_31228,N_31438);
or U31898 (N_31898,N_31473,N_31266);
nor U31899 (N_31899,N_31418,N_31438);
nand U31900 (N_31900,N_31123,N_31346);
nand U31901 (N_31901,N_31462,N_31287);
and U31902 (N_31902,N_31012,N_31489);
nand U31903 (N_31903,N_31337,N_31147);
and U31904 (N_31904,N_31440,N_31364);
or U31905 (N_31905,N_31448,N_31183);
nand U31906 (N_31906,N_31013,N_31008);
or U31907 (N_31907,N_31255,N_31002);
nand U31908 (N_31908,N_31229,N_31172);
or U31909 (N_31909,N_31206,N_31354);
nand U31910 (N_31910,N_31015,N_31344);
nor U31911 (N_31911,N_31468,N_31498);
nor U31912 (N_31912,N_31471,N_31009);
nand U31913 (N_31913,N_31060,N_31086);
or U31914 (N_31914,N_31061,N_31379);
xor U31915 (N_31915,N_31147,N_31313);
and U31916 (N_31916,N_31136,N_31391);
xnor U31917 (N_31917,N_31039,N_31068);
or U31918 (N_31918,N_31097,N_31433);
nand U31919 (N_31919,N_31226,N_31043);
nand U31920 (N_31920,N_31311,N_31039);
xor U31921 (N_31921,N_31208,N_31045);
nor U31922 (N_31922,N_31356,N_31052);
or U31923 (N_31923,N_31442,N_31476);
nor U31924 (N_31924,N_31056,N_31429);
nand U31925 (N_31925,N_31215,N_31450);
and U31926 (N_31926,N_31434,N_31106);
nor U31927 (N_31927,N_31021,N_31347);
and U31928 (N_31928,N_31120,N_31212);
and U31929 (N_31929,N_31230,N_31462);
xnor U31930 (N_31930,N_31488,N_31007);
nand U31931 (N_31931,N_31311,N_31477);
xor U31932 (N_31932,N_31323,N_31153);
and U31933 (N_31933,N_31176,N_31145);
nor U31934 (N_31934,N_31318,N_31400);
xnor U31935 (N_31935,N_31062,N_31109);
or U31936 (N_31936,N_31333,N_31078);
or U31937 (N_31937,N_31459,N_31445);
xnor U31938 (N_31938,N_31320,N_31145);
xor U31939 (N_31939,N_31437,N_31143);
nand U31940 (N_31940,N_31375,N_31432);
nor U31941 (N_31941,N_31005,N_31297);
nand U31942 (N_31942,N_31236,N_31480);
and U31943 (N_31943,N_31075,N_31227);
nand U31944 (N_31944,N_31076,N_31330);
xnor U31945 (N_31945,N_31128,N_31490);
nand U31946 (N_31946,N_31482,N_31476);
nor U31947 (N_31947,N_31084,N_31040);
nor U31948 (N_31948,N_31261,N_31034);
xnor U31949 (N_31949,N_31194,N_31335);
nand U31950 (N_31950,N_31002,N_31441);
and U31951 (N_31951,N_31151,N_31015);
and U31952 (N_31952,N_31257,N_31281);
xnor U31953 (N_31953,N_31199,N_31296);
nand U31954 (N_31954,N_31391,N_31301);
nand U31955 (N_31955,N_31328,N_31167);
xnor U31956 (N_31956,N_31018,N_31027);
and U31957 (N_31957,N_31470,N_31464);
nor U31958 (N_31958,N_31361,N_31421);
and U31959 (N_31959,N_31221,N_31010);
and U31960 (N_31960,N_31007,N_31071);
xnor U31961 (N_31961,N_31359,N_31014);
nand U31962 (N_31962,N_31401,N_31272);
and U31963 (N_31963,N_31068,N_31247);
nand U31964 (N_31964,N_31452,N_31026);
or U31965 (N_31965,N_31041,N_31319);
nor U31966 (N_31966,N_31271,N_31451);
or U31967 (N_31967,N_31023,N_31180);
nand U31968 (N_31968,N_31453,N_31344);
xor U31969 (N_31969,N_31388,N_31454);
xor U31970 (N_31970,N_31052,N_31263);
and U31971 (N_31971,N_31036,N_31461);
nand U31972 (N_31972,N_31474,N_31100);
nor U31973 (N_31973,N_31132,N_31066);
nor U31974 (N_31974,N_31118,N_31426);
xnor U31975 (N_31975,N_31151,N_31318);
nor U31976 (N_31976,N_31031,N_31340);
xnor U31977 (N_31977,N_31216,N_31079);
and U31978 (N_31978,N_31239,N_31363);
xor U31979 (N_31979,N_31491,N_31450);
nor U31980 (N_31980,N_31386,N_31002);
xnor U31981 (N_31981,N_31457,N_31054);
and U31982 (N_31982,N_31002,N_31167);
or U31983 (N_31983,N_31226,N_31078);
nand U31984 (N_31984,N_31252,N_31389);
nand U31985 (N_31985,N_31294,N_31243);
or U31986 (N_31986,N_31238,N_31123);
or U31987 (N_31987,N_31105,N_31492);
nor U31988 (N_31988,N_31148,N_31186);
nand U31989 (N_31989,N_31157,N_31241);
xnor U31990 (N_31990,N_31352,N_31373);
nand U31991 (N_31991,N_31321,N_31460);
or U31992 (N_31992,N_31146,N_31020);
nor U31993 (N_31993,N_31134,N_31206);
nor U31994 (N_31994,N_31483,N_31402);
or U31995 (N_31995,N_31018,N_31227);
and U31996 (N_31996,N_31336,N_31366);
or U31997 (N_31997,N_31399,N_31179);
nand U31998 (N_31998,N_31246,N_31492);
xor U31999 (N_31999,N_31052,N_31171);
nand U32000 (N_32000,N_31770,N_31870);
and U32001 (N_32001,N_31590,N_31962);
or U32002 (N_32002,N_31974,N_31919);
nand U32003 (N_32003,N_31698,N_31936);
or U32004 (N_32004,N_31914,N_31737);
or U32005 (N_32005,N_31857,N_31676);
xor U32006 (N_32006,N_31742,N_31834);
and U32007 (N_32007,N_31838,N_31901);
nor U32008 (N_32008,N_31598,N_31675);
and U32009 (N_32009,N_31509,N_31597);
and U32010 (N_32010,N_31904,N_31721);
nand U32011 (N_32011,N_31532,N_31640);
xnor U32012 (N_32012,N_31589,N_31554);
and U32013 (N_32013,N_31650,N_31712);
xnor U32014 (N_32014,N_31806,N_31989);
nand U32015 (N_32015,N_31651,N_31607);
nand U32016 (N_32016,N_31922,N_31969);
nor U32017 (N_32017,N_31735,N_31937);
or U32018 (N_32018,N_31622,N_31624);
and U32019 (N_32019,N_31580,N_31998);
xor U32020 (N_32020,N_31821,N_31811);
or U32021 (N_32021,N_31574,N_31959);
xnor U32022 (N_32022,N_31911,N_31978);
nand U32023 (N_32023,N_31601,N_31536);
nand U32024 (N_32024,N_31957,N_31505);
xor U32025 (N_32025,N_31518,N_31513);
xor U32026 (N_32026,N_31813,N_31582);
xnor U32027 (N_32027,N_31700,N_31592);
xor U32028 (N_32028,N_31760,N_31584);
and U32029 (N_32029,N_31875,N_31689);
xnor U32030 (N_32030,N_31858,N_31855);
or U32031 (N_32031,N_31779,N_31555);
and U32032 (N_32032,N_31940,N_31500);
nor U32033 (N_32033,N_31780,N_31568);
and U32034 (N_32034,N_31877,N_31548);
and U32035 (N_32035,N_31688,N_31757);
or U32036 (N_32036,N_31845,N_31611);
nor U32037 (N_32037,N_31741,N_31558);
xor U32038 (N_32038,N_31625,N_31943);
nand U32039 (N_32039,N_31502,N_31679);
and U32040 (N_32040,N_31774,N_31523);
and U32041 (N_32041,N_31852,N_31831);
or U32042 (N_32042,N_31881,N_31748);
nor U32043 (N_32043,N_31733,N_31690);
nor U32044 (N_32044,N_31933,N_31667);
or U32045 (N_32045,N_31983,N_31599);
nor U32046 (N_32046,N_31678,N_31950);
nand U32047 (N_32047,N_31645,N_31866);
or U32048 (N_32048,N_31850,N_31999);
nor U32049 (N_32049,N_31872,N_31653);
and U32050 (N_32050,N_31562,N_31784);
nand U32051 (N_32051,N_31517,N_31749);
nor U32052 (N_32052,N_31656,N_31594);
xor U32053 (N_32053,N_31843,N_31539);
or U32054 (N_32054,N_31844,N_31766);
nor U32055 (N_32055,N_31665,N_31932);
xnor U32056 (N_32056,N_31588,N_31612);
nor U32057 (N_32057,N_31994,N_31930);
nand U32058 (N_32058,N_31777,N_31764);
xor U32059 (N_32059,N_31934,N_31731);
nor U32060 (N_32060,N_31706,N_31958);
nor U32061 (N_32061,N_31711,N_31863);
xnor U32062 (N_32062,N_31802,N_31514);
nor U32063 (N_32063,N_31918,N_31761);
xor U32064 (N_32064,N_31931,N_31893);
xnor U32065 (N_32065,N_31644,N_31797);
xor U32066 (N_32066,N_31605,N_31684);
or U32067 (N_32067,N_31672,N_31842);
nand U32068 (N_32068,N_31729,N_31623);
and U32069 (N_32069,N_31864,N_31659);
or U32070 (N_32070,N_31544,N_31745);
or U32071 (N_32071,N_31683,N_31907);
nand U32072 (N_32072,N_31669,N_31738);
xor U32073 (N_32073,N_31878,N_31686);
and U32074 (N_32074,N_31581,N_31586);
xor U32075 (N_32075,N_31719,N_31890);
nand U32076 (N_32076,N_31677,N_31680);
and U32077 (N_32077,N_31552,N_31995);
xor U32078 (N_32078,N_31848,N_31786);
nor U32079 (N_32079,N_31519,N_31693);
or U32080 (N_32080,N_31810,N_31723);
nand U32081 (N_32081,N_31655,N_31867);
nor U32082 (N_32082,N_31746,N_31968);
or U32083 (N_32083,N_31906,N_31840);
nand U32084 (N_32084,N_31501,N_31992);
nor U32085 (N_32085,N_31533,N_31946);
nor U32086 (N_32086,N_31527,N_31649);
nand U32087 (N_32087,N_31977,N_31908);
and U32088 (N_32088,N_31530,N_31986);
xnor U32089 (N_32089,N_31829,N_31614);
xnor U32090 (N_32090,N_31814,N_31639);
and U32091 (N_32091,N_31824,N_31879);
and U32092 (N_32092,N_31565,N_31726);
xor U32093 (N_32093,N_31947,N_31615);
xnor U32094 (N_32094,N_31982,N_31902);
or U32095 (N_32095,N_31661,N_31817);
and U32096 (N_32096,N_31516,N_31572);
xor U32097 (N_32097,N_31851,N_31788);
nor U32098 (N_32098,N_31534,N_31541);
or U32099 (N_32099,N_31778,N_31634);
nor U32100 (N_32100,N_31671,N_31874);
or U32101 (N_32101,N_31713,N_31799);
or U32102 (N_32102,N_31510,N_31979);
nor U32103 (N_32103,N_31951,N_31961);
nor U32104 (N_32104,N_31809,N_31724);
or U32105 (N_32105,N_31646,N_31553);
and U32106 (N_32106,N_31576,N_31567);
nand U32107 (N_32107,N_31805,N_31663);
and U32108 (N_32108,N_31709,N_31755);
nor U32109 (N_32109,N_31954,N_31892);
nor U32110 (N_32110,N_31604,N_31620);
nor U32111 (N_32111,N_31522,N_31561);
and U32112 (N_32112,N_31984,N_31702);
and U32113 (N_32113,N_31616,N_31728);
or U32114 (N_32114,N_31920,N_31585);
or U32115 (N_32115,N_31791,N_31503);
or U32116 (N_32116,N_31573,N_31606);
xnor U32117 (N_32117,N_31915,N_31751);
or U32118 (N_32118,N_31769,N_31662);
nand U32119 (N_32119,N_31538,N_31826);
or U32120 (N_32120,N_31743,N_31990);
nor U32121 (N_32121,N_31781,N_31971);
nor U32122 (N_32122,N_31765,N_31900);
nor U32123 (N_32123,N_31832,N_31658);
or U32124 (N_32124,N_31550,N_31626);
xnor U32125 (N_32125,N_31525,N_31638);
nand U32126 (N_32126,N_31839,N_31570);
xnor U32127 (N_32127,N_31705,N_31627);
xor U32128 (N_32128,N_31520,N_31593);
xor U32129 (N_32129,N_31512,N_31822);
or U32130 (N_32130,N_31528,N_31825);
and U32131 (N_32131,N_31710,N_31642);
nand U32132 (N_32132,N_31944,N_31886);
xor U32133 (N_32133,N_31960,N_31707);
or U32134 (N_32134,N_31635,N_31889);
nor U32135 (N_32135,N_31563,N_31673);
or U32136 (N_32136,N_31691,N_31583);
nand U32137 (N_32137,N_31542,N_31682);
and U32138 (N_32138,N_31966,N_31579);
xnor U32139 (N_32139,N_31602,N_31785);
and U32140 (N_32140,N_31942,N_31714);
xnor U32141 (N_32141,N_31657,N_31637);
nand U32142 (N_32142,N_31955,N_31923);
and U32143 (N_32143,N_31758,N_31648);
or U32144 (N_32144,N_31718,N_31894);
nand U32145 (N_32145,N_31981,N_31609);
or U32146 (N_32146,N_31701,N_31964);
nor U32147 (N_32147,N_31692,N_31985);
and U32148 (N_32148,N_31796,N_31652);
nor U32149 (N_32149,N_31571,N_31792);
or U32150 (N_32150,N_31628,N_31587);
or U32151 (N_32151,N_31703,N_31569);
or U32152 (N_32152,N_31747,N_31980);
nand U32153 (N_32153,N_31849,N_31762);
or U32154 (N_32154,N_31595,N_31647);
xor U32155 (N_32155,N_31883,N_31861);
nor U32156 (N_32156,N_31921,N_31704);
and U32157 (N_32157,N_31660,N_31750);
or U32158 (N_32158,N_31540,N_31754);
and U32159 (N_32159,N_31631,N_31896);
xor U32160 (N_32160,N_31506,N_31965);
and U32161 (N_32161,N_31551,N_31722);
or U32162 (N_32162,N_31531,N_31591);
nor U32163 (N_32163,N_31827,N_31508);
xor U32164 (N_32164,N_31521,N_31577);
or U32165 (N_32165,N_31939,N_31629);
and U32166 (N_32166,N_31716,N_31815);
nor U32167 (N_32167,N_31670,N_31860);
nand U32168 (N_32168,N_31790,N_31546);
xor U32169 (N_32169,N_31812,N_31991);
or U32170 (N_32170,N_31800,N_31873);
nor U32171 (N_32171,N_31876,N_31732);
nor U32172 (N_32172,N_31668,N_31756);
or U32173 (N_32173,N_31524,N_31925);
xnor U32174 (N_32174,N_31898,N_31888);
or U32175 (N_32175,N_31636,N_31697);
nor U32176 (N_32176,N_31818,N_31808);
nand U32177 (N_32177,N_31807,N_31948);
nor U32178 (N_32178,N_31507,N_31926);
and U32179 (N_32179,N_31578,N_31763);
nand U32180 (N_32180,N_31734,N_31853);
xnor U32181 (N_32181,N_31776,N_31783);
or U32182 (N_32182,N_31730,N_31854);
or U32183 (N_32183,N_31847,N_31643);
xor U32184 (N_32184,N_31856,N_31909);
xor U32185 (N_32185,N_31720,N_31833);
xor U32186 (N_32186,N_31685,N_31841);
and U32187 (N_32187,N_31967,N_31752);
xor U32188 (N_32188,N_31696,N_31596);
and U32189 (N_32189,N_31687,N_31988);
nor U32190 (N_32190,N_31794,N_31801);
or U32191 (N_32191,N_31529,N_31767);
and U32192 (N_32192,N_31972,N_31976);
nand U32193 (N_32193,N_31740,N_31666);
nand U32194 (N_32194,N_31941,N_31997);
xor U32195 (N_32195,N_31559,N_31793);
nand U32196 (N_32196,N_31816,N_31771);
or U32197 (N_32197,N_31880,N_31935);
nor U32198 (N_32198,N_31547,N_31803);
and U32199 (N_32199,N_31905,N_31526);
and U32200 (N_32200,N_31557,N_31613);
nor U32201 (N_32201,N_31975,N_31913);
xnor U32202 (N_32202,N_31782,N_31535);
and U32203 (N_32203,N_31820,N_31927);
or U32204 (N_32204,N_31600,N_31887);
xor U32205 (N_32205,N_31694,N_31798);
nor U32206 (N_32206,N_31775,N_31895);
nand U32207 (N_32207,N_31910,N_31549);
nor U32208 (N_32208,N_31917,N_31836);
nor U32209 (N_32209,N_31772,N_31543);
xnor U32210 (N_32210,N_31884,N_31823);
and U32211 (N_32211,N_31768,N_31759);
nor U32212 (N_32212,N_31504,N_31556);
or U32213 (N_32213,N_31727,N_31871);
and U32214 (N_32214,N_31787,N_31511);
nor U32215 (N_32215,N_31610,N_31725);
and U32216 (N_32216,N_31903,N_31885);
or U32217 (N_32217,N_31633,N_31545);
nand U32218 (N_32218,N_31868,N_31912);
and U32219 (N_32219,N_31753,N_31828);
or U32220 (N_32220,N_31938,N_31564);
xor U32221 (N_32221,N_31630,N_31744);
or U32222 (N_32222,N_31862,N_31891);
nor U32223 (N_32223,N_31928,N_31945);
nor U32224 (N_32224,N_31952,N_31956);
xor U32225 (N_32225,N_31865,N_31537);
nor U32226 (N_32226,N_31654,N_31869);
and U32227 (N_32227,N_31789,N_31996);
or U32228 (N_32228,N_31708,N_31603);
nor U32229 (N_32229,N_31575,N_31882);
nor U32230 (N_32230,N_31773,N_31859);
and U32231 (N_32231,N_31681,N_31899);
or U32232 (N_32232,N_31804,N_31560);
nand U32233 (N_32233,N_31715,N_31963);
nor U32234 (N_32234,N_31664,N_31739);
nor U32235 (N_32235,N_31617,N_31897);
or U32236 (N_32236,N_31916,N_31970);
or U32237 (N_32237,N_31717,N_31674);
or U32238 (N_32238,N_31987,N_31566);
or U32239 (N_32239,N_31641,N_31993);
nor U32240 (N_32240,N_31608,N_31830);
or U32241 (N_32241,N_31846,N_31929);
xor U32242 (N_32242,N_31949,N_31632);
or U32243 (N_32243,N_31619,N_31924);
or U32244 (N_32244,N_31736,N_31837);
or U32245 (N_32245,N_31695,N_31515);
or U32246 (N_32246,N_31819,N_31953);
and U32247 (N_32247,N_31795,N_31618);
and U32248 (N_32248,N_31699,N_31621);
or U32249 (N_32249,N_31835,N_31973);
nand U32250 (N_32250,N_31970,N_31898);
nand U32251 (N_32251,N_31652,N_31722);
nor U32252 (N_32252,N_31734,N_31935);
xor U32253 (N_32253,N_31889,N_31624);
nor U32254 (N_32254,N_31731,N_31709);
and U32255 (N_32255,N_31901,N_31965);
or U32256 (N_32256,N_31500,N_31955);
nor U32257 (N_32257,N_31908,N_31781);
or U32258 (N_32258,N_31561,N_31739);
nor U32259 (N_32259,N_31543,N_31719);
and U32260 (N_32260,N_31878,N_31895);
xnor U32261 (N_32261,N_31542,N_31666);
or U32262 (N_32262,N_31991,N_31536);
or U32263 (N_32263,N_31814,N_31753);
xnor U32264 (N_32264,N_31501,N_31559);
xnor U32265 (N_32265,N_31677,N_31947);
xor U32266 (N_32266,N_31910,N_31810);
nand U32267 (N_32267,N_31714,N_31542);
xnor U32268 (N_32268,N_31932,N_31754);
nand U32269 (N_32269,N_31538,N_31784);
and U32270 (N_32270,N_31903,N_31978);
xor U32271 (N_32271,N_31871,N_31512);
xor U32272 (N_32272,N_31889,N_31816);
xnor U32273 (N_32273,N_31984,N_31830);
nand U32274 (N_32274,N_31650,N_31537);
xor U32275 (N_32275,N_31937,N_31796);
and U32276 (N_32276,N_31583,N_31555);
nor U32277 (N_32277,N_31548,N_31966);
nor U32278 (N_32278,N_31659,N_31874);
and U32279 (N_32279,N_31984,N_31562);
xor U32280 (N_32280,N_31741,N_31738);
nand U32281 (N_32281,N_31845,N_31968);
nor U32282 (N_32282,N_31982,N_31977);
nor U32283 (N_32283,N_31809,N_31582);
nand U32284 (N_32284,N_31839,N_31840);
xor U32285 (N_32285,N_31558,N_31675);
and U32286 (N_32286,N_31683,N_31617);
nor U32287 (N_32287,N_31719,N_31562);
xor U32288 (N_32288,N_31568,N_31561);
nor U32289 (N_32289,N_31773,N_31839);
nand U32290 (N_32290,N_31513,N_31912);
or U32291 (N_32291,N_31524,N_31644);
xnor U32292 (N_32292,N_31805,N_31831);
nor U32293 (N_32293,N_31702,N_31968);
and U32294 (N_32294,N_31739,N_31988);
nor U32295 (N_32295,N_31593,N_31708);
xnor U32296 (N_32296,N_31585,N_31940);
xnor U32297 (N_32297,N_31980,N_31876);
nand U32298 (N_32298,N_31817,N_31789);
xor U32299 (N_32299,N_31655,N_31651);
xor U32300 (N_32300,N_31506,N_31514);
and U32301 (N_32301,N_31863,N_31898);
or U32302 (N_32302,N_31965,N_31578);
or U32303 (N_32303,N_31550,N_31796);
or U32304 (N_32304,N_31906,N_31525);
nor U32305 (N_32305,N_31859,N_31791);
nand U32306 (N_32306,N_31563,N_31893);
or U32307 (N_32307,N_31846,N_31925);
or U32308 (N_32308,N_31698,N_31956);
nor U32309 (N_32309,N_31985,N_31897);
nor U32310 (N_32310,N_31885,N_31952);
and U32311 (N_32311,N_31993,N_31866);
or U32312 (N_32312,N_31663,N_31917);
nor U32313 (N_32313,N_31629,N_31971);
nand U32314 (N_32314,N_31502,N_31727);
nand U32315 (N_32315,N_31794,N_31769);
or U32316 (N_32316,N_31908,N_31823);
nor U32317 (N_32317,N_31669,N_31736);
and U32318 (N_32318,N_31791,N_31679);
xnor U32319 (N_32319,N_31686,N_31576);
and U32320 (N_32320,N_31610,N_31582);
or U32321 (N_32321,N_31554,N_31588);
nor U32322 (N_32322,N_31577,N_31716);
nor U32323 (N_32323,N_31774,N_31635);
or U32324 (N_32324,N_31858,N_31950);
or U32325 (N_32325,N_31762,N_31657);
nor U32326 (N_32326,N_31718,N_31849);
and U32327 (N_32327,N_31851,N_31844);
xnor U32328 (N_32328,N_31697,N_31634);
nand U32329 (N_32329,N_31952,N_31740);
nor U32330 (N_32330,N_31524,N_31994);
nand U32331 (N_32331,N_31920,N_31708);
and U32332 (N_32332,N_31628,N_31570);
nor U32333 (N_32333,N_31960,N_31592);
nor U32334 (N_32334,N_31543,N_31628);
nand U32335 (N_32335,N_31513,N_31968);
nor U32336 (N_32336,N_31905,N_31848);
nor U32337 (N_32337,N_31516,N_31721);
nand U32338 (N_32338,N_31787,N_31843);
or U32339 (N_32339,N_31823,N_31631);
nor U32340 (N_32340,N_31807,N_31782);
xnor U32341 (N_32341,N_31684,N_31755);
nor U32342 (N_32342,N_31677,N_31860);
nor U32343 (N_32343,N_31989,N_31593);
nand U32344 (N_32344,N_31911,N_31636);
nand U32345 (N_32345,N_31959,N_31504);
nand U32346 (N_32346,N_31700,N_31600);
nand U32347 (N_32347,N_31592,N_31604);
nor U32348 (N_32348,N_31585,N_31824);
nor U32349 (N_32349,N_31661,N_31505);
and U32350 (N_32350,N_31926,N_31710);
nor U32351 (N_32351,N_31718,N_31722);
xnor U32352 (N_32352,N_31665,N_31734);
and U32353 (N_32353,N_31696,N_31521);
xnor U32354 (N_32354,N_31635,N_31695);
xor U32355 (N_32355,N_31507,N_31722);
nor U32356 (N_32356,N_31519,N_31836);
and U32357 (N_32357,N_31998,N_31886);
nand U32358 (N_32358,N_31765,N_31761);
nand U32359 (N_32359,N_31807,N_31825);
nand U32360 (N_32360,N_31753,N_31767);
or U32361 (N_32361,N_31854,N_31501);
nor U32362 (N_32362,N_31931,N_31607);
or U32363 (N_32363,N_31921,N_31634);
xor U32364 (N_32364,N_31819,N_31603);
xor U32365 (N_32365,N_31596,N_31587);
or U32366 (N_32366,N_31544,N_31539);
xnor U32367 (N_32367,N_31672,N_31694);
nand U32368 (N_32368,N_31518,N_31605);
nand U32369 (N_32369,N_31812,N_31565);
or U32370 (N_32370,N_31844,N_31703);
xnor U32371 (N_32371,N_31634,N_31625);
nand U32372 (N_32372,N_31972,N_31705);
and U32373 (N_32373,N_31969,N_31517);
or U32374 (N_32374,N_31925,N_31872);
xor U32375 (N_32375,N_31667,N_31609);
and U32376 (N_32376,N_31973,N_31505);
and U32377 (N_32377,N_31773,N_31842);
and U32378 (N_32378,N_31601,N_31835);
xor U32379 (N_32379,N_31983,N_31914);
or U32380 (N_32380,N_31640,N_31916);
xnor U32381 (N_32381,N_31970,N_31859);
nand U32382 (N_32382,N_31587,N_31941);
nand U32383 (N_32383,N_31771,N_31531);
and U32384 (N_32384,N_31570,N_31798);
or U32385 (N_32385,N_31572,N_31635);
xnor U32386 (N_32386,N_31718,N_31855);
nor U32387 (N_32387,N_31555,N_31569);
and U32388 (N_32388,N_31736,N_31853);
nand U32389 (N_32389,N_31910,N_31957);
nor U32390 (N_32390,N_31716,N_31978);
nor U32391 (N_32391,N_31813,N_31627);
nor U32392 (N_32392,N_31898,N_31870);
and U32393 (N_32393,N_31826,N_31573);
and U32394 (N_32394,N_31746,N_31558);
xor U32395 (N_32395,N_31934,N_31985);
xor U32396 (N_32396,N_31828,N_31611);
and U32397 (N_32397,N_31933,N_31736);
and U32398 (N_32398,N_31781,N_31518);
nand U32399 (N_32399,N_31571,N_31749);
xor U32400 (N_32400,N_31775,N_31713);
xor U32401 (N_32401,N_31593,N_31628);
xor U32402 (N_32402,N_31629,N_31889);
or U32403 (N_32403,N_31813,N_31844);
and U32404 (N_32404,N_31833,N_31672);
and U32405 (N_32405,N_31702,N_31677);
or U32406 (N_32406,N_31690,N_31794);
or U32407 (N_32407,N_31854,N_31909);
xnor U32408 (N_32408,N_31750,N_31549);
and U32409 (N_32409,N_31742,N_31999);
xor U32410 (N_32410,N_31597,N_31943);
and U32411 (N_32411,N_31591,N_31583);
nor U32412 (N_32412,N_31904,N_31866);
and U32413 (N_32413,N_31905,N_31558);
and U32414 (N_32414,N_31772,N_31553);
nand U32415 (N_32415,N_31517,N_31689);
or U32416 (N_32416,N_31896,N_31740);
nor U32417 (N_32417,N_31726,N_31949);
nand U32418 (N_32418,N_31905,N_31941);
xnor U32419 (N_32419,N_31966,N_31992);
nor U32420 (N_32420,N_31920,N_31754);
nor U32421 (N_32421,N_31613,N_31956);
nor U32422 (N_32422,N_31773,N_31709);
nand U32423 (N_32423,N_31740,N_31598);
nand U32424 (N_32424,N_31851,N_31688);
or U32425 (N_32425,N_31902,N_31930);
xnor U32426 (N_32426,N_31617,N_31942);
nor U32427 (N_32427,N_31646,N_31783);
nor U32428 (N_32428,N_31920,N_31987);
nand U32429 (N_32429,N_31788,N_31549);
or U32430 (N_32430,N_31880,N_31675);
or U32431 (N_32431,N_31551,N_31903);
xnor U32432 (N_32432,N_31865,N_31553);
xnor U32433 (N_32433,N_31605,N_31997);
nor U32434 (N_32434,N_31882,N_31614);
nand U32435 (N_32435,N_31825,N_31868);
nand U32436 (N_32436,N_31866,N_31872);
or U32437 (N_32437,N_31645,N_31915);
nor U32438 (N_32438,N_31802,N_31713);
nand U32439 (N_32439,N_31761,N_31904);
nor U32440 (N_32440,N_31694,N_31815);
nor U32441 (N_32441,N_31879,N_31909);
nand U32442 (N_32442,N_31898,N_31668);
and U32443 (N_32443,N_31981,N_31665);
or U32444 (N_32444,N_31861,N_31547);
or U32445 (N_32445,N_31970,N_31567);
nor U32446 (N_32446,N_31511,N_31615);
xor U32447 (N_32447,N_31737,N_31893);
xor U32448 (N_32448,N_31843,N_31752);
or U32449 (N_32449,N_31672,N_31914);
xor U32450 (N_32450,N_31526,N_31698);
and U32451 (N_32451,N_31573,N_31865);
or U32452 (N_32452,N_31726,N_31881);
xor U32453 (N_32453,N_31821,N_31682);
xor U32454 (N_32454,N_31976,N_31768);
or U32455 (N_32455,N_31667,N_31915);
nand U32456 (N_32456,N_31706,N_31736);
and U32457 (N_32457,N_31572,N_31894);
nand U32458 (N_32458,N_31862,N_31598);
and U32459 (N_32459,N_31875,N_31739);
and U32460 (N_32460,N_31954,N_31811);
or U32461 (N_32461,N_31518,N_31614);
xor U32462 (N_32462,N_31729,N_31796);
nand U32463 (N_32463,N_31969,N_31981);
xnor U32464 (N_32464,N_31778,N_31676);
nor U32465 (N_32465,N_31680,N_31692);
nand U32466 (N_32466,N_31936,N_31974);
or U32467 (N_32467,N_31996,N_31652);
xnor U32468 (N_32468,N_31740,N_31597);
xnor U32469 (N_32469,N_31995,N_31912);
or U32470 (N_32470,N_31930,N_31628);
or U32471 (N_32471,N_31824,N_31819);
nor U32472 (N_32472,N_31523,N_31741);
xor U32473 (N_32473,N_31779,N_31531);
or U32474 (N_32474,N_31649,N_31831);
or U32475 (N_32475,N_31985,N_31674);
and U32476 (N_32476,N_31577,N_31617);
and U32477 (N_32477,N_31565,N_31512);
and U32478 (N_32478,N_31674,N_31514);
nand U32479 (N_32479,N_31965,N_31898);
xor U32480 (N_32480,N_31963,N_31833);
nor U32481 (N_32481,N_31798,N_31587);
and U32482 (N_32482,N_31893,N_31761);
nand U32483 (N_32483,N_31796,N_31785);
and U32484 (N_32484,N_31919,N_31571);
or U32485 (N_32485,N_31954,N_31840);
nor U32486 (N_32486,N_31791,N_31905);
xor U32487 (N_32487,N_31761,N_31537);
nand U32488 (N_32488,N_31891,N_31666);
xnor U32489 (N_32489,N_31967,N_31821);
and U32490 (N_32490,N_31624,N_31593);
nor U32491 (N_32491,N_31899,N_31683);
and U32492 (N_32492,N_31544,N_31893);
and U32493 (N_32493,N_31781,N_31564);
xor U32494 (N_32494,N_31698,N_31651);
nand U32495 (N_32495,N_31583,N_31782);
xnor U32496 (N_32496,N_31817,N_31814);
and U32497 (N_32497,N_31949,N_31951);
xnor U32498 (N_32498,N_31972,N_31654);
nor U32499 (N_32499,N_31775,N_31677);
and U32500 (N_32500,N_32055,N_32290);
nand U32501 (N_32501,N_32469,N_32415);
nor U32502 (N_32502,N_32205,N_32067);
and U32503 (N_32503,N_32381,N_32107);
xnor U32504 (N_32504,N_32320,N_32074);
nand U32505 (N_32505,N_32121,N_32164);
or U32506 (N_32506,N_32468,N_32158);
or U32507 (N_32507,N_32224,N_32457);
nand U32508 (N_32508,N_32431,N_32222);
or U32509 (N_32509,N_32418,N_32004);
nor U32510 (N_32510,N_32408,N_32313);
or U32511 (N_32511,N_32422,N_32407);
nand U32512 (N_32512,N_32272,N_32363);
xnor U32513 (N_32513,N_32209,N_32101);
and U32514 (N_32514,N_32474,N_32297);
xor U32515 (N_32515,N_32356,N_32192);
nor U32516 (N_32516,N_32479,N_32384);
nand U32517 (N_32517,N_32033,N_32119);
xor U32518 (N_32518,N_32355,N_32047);
or U32519 (N_32519,N_32338,N_32174);
or U32520 (N_32520,N_32375,N_32348);
xnor U32521 (N_32521,N_32476,N_32044);
or U32522 (N_32522,N_32060,N_32030);
nand U32523 (N_32523,N_32072,N_32271);
and U32524 (N_32524,N_32050,N_32152);
and U32525 (N_32525,N_32211,N_32478);
nor U32526 (N_32526,N_32210,N_32143);
nor U32527 (N_32527,N_32185,N_32423);
xnor U32528 (N_32528,N_32166,N_32439);
nor U32529 (N_32529,N_32245,N_32347);
or U32530 (N_32530,N_32230,N_32144);
and U32531 (N_32531,N_32082,N_32485);
nor U32532 (N_32532,N_32481,N_32462);
nand U32533 (N_32533,N_32279,N_32006);
or U32534 (N_32534,N_32295,N_32373);
nor U32535 (N_32535,N_32333,N_32294);
xor U32536 (N_32536,N_32369,N_32339);
nand U32537 (N_32537,N_32093,N_32013);
xnor U32538 (N_32538,N_32089,N_32366);
nor U32539 (N_32539,N_32113,N_32496);
nor U32540 (N_32540,N_32206,N_32054);
nand U32541 (N_32541,N_32497,N_32332);
or U32542 (N_32542,N_32103,N_32216);
and U32543 (N_32543,N_32259,N_32377);
nor U32544 (N_32544,N_32094,N_32203);
nor U32545 (N_32545,N_32023,N_32043);
nor U32546 (N_32546,N_32424,N_32383);
or U32547 (N_32547,N_32123,N_32201);
xor U32548 (N_32548,N_32360,N_32213);
nand U32549 (N_32549,N_32343,N_32005);
xnor U32550 (N_32550,N_32122,N_32168);
and U32551 (N_32551,N_32191,N_32065);
or U32552 (N_32552,N_32039,N_32437);
and U32553 (N_32553,N_32076,N_32127);
or U32554 (N_32554,N_32414,N_32098);
nand U32555 (N_32555,N_32133,N_32025);
nor U32556 (N_32556,N_32287,N_32268);
or U32557 (N_32557,N_32417,N_32198);
nand U32558 (N_32558,N_32329,N_32058);
and U32559 (N_32559,N_32466,N_32326);
or U32560 (N_32560,N_32077,N_32021);
or U32561 (N_32561,N_32003,N_32063);
nand U32562 (N_32562,N_32483,N_32260);
and U32563 (N_32563,N_32099,N_32432);
nor U32564 (N_32564,N_32292,N_32264);
xor U32565 (N_32565,N_32492,N_32386);
or U32566 (N_32566,N_32017,N_32342);
nand U32567 (N_32567,N_32188,N_32455);
and U32568 (N_32568,N_32199,N_32438);
xnor U32569 (N_32569,N_32250,N_32440);
xnor U32570 (N_32570,N_32461,N_32036);
and U32571 (N_32571,N_32079,N_32112);
nor U32572 (N_32572,N_32219,N_32404);
xor U32573 (N_32573,N_32037,N_32235);
or U32574 (N_32574,N_32499,N_32467);
or U32575 (N_32575,N_32080,N_32236);
or U32576 (N_32576,N_32128,N_32350);
nand U32577 (N_32577,N_32001,N_32181);
nand U32578 (N_32578,N_32117,N_32477);
and U32579 (N_32579,N_32396,N_32011);
and U32580 (N_32580,N_32317,N_32471);
nand U32581 (N_32581,N_32125,N_32393);
and U32582 (N_32582,N_32159,N_32090);
or U32583 (N_32583,N_32177,N_32406);
and U32584 (N_32584,N_32040,N_32301);
or U32585 (N_32585,N_32064,N_32286);
xnor U32586 (N_32586,N_32412,N_32374);
xnor U32587 (N_32587,N_32311,N_32097);
nor U32588 (N_32588,N_32325,N_32156);
nand U32589 (N_32589,N_32026,N_32436);
nand U32590 (N_32590,N_32204,N_32042);
nor U32591 (N_32591,N_32397,N_32298);
nor U32592 (N_32592,N_32134,N_32251);
nor U32593 (N_32593,N_32232,N_32020);
nand U32594 (N_32594,N_32456,N_32187);
xor U32595 (N_32595,N_32458,N_32172);
nor U32596 (N_32596,N_32409,N_32029);
and U32597 (N_32597,N_32255,N_32129);
nor U32598 (N_32598,N_32150,N_32429);
nor U32599 (N_32599,N_32357,N_32114);
and U32600 (N_32600,N_32370,N_32394);
nand U32601 (N_32601,N_32131,N_32028);
or U32602 (N_32602,N_32009,N_32254);
xor U32603 (N_32603,N_32487,N_32304);
and U32604 (N_32604,N_32484,N_32282);
xnor U32605 (N_32605,N_32000,N_32179);
and U32606 (N_32606,N_32249,N_32486);
or U32607 (N_32607,N_32240,N_32330);
or U32608 (N_32608,N_32274,N_32170);
nand U32609 (N_32609,N_32163,N_32053);
nor U32610 (N_32610,N_32390,N_32454);
nor U32611 (N_32611,N_32277,N_32184);
nor U32612 (N_32612,N_32175,N_32038);
or U32613 (N_32613,N_32482,N_32388);
nor U32614 (N_32614,N_32139,N_32078);
or U32615 (N_32615,N_32402,N_32176);
xor U32616 (N_32616,N_32108,N_32171);
xor U32617 (N_32617,N_32262,N_32495);
or U32618 (N_32618,N_32307,N_32096);
nor U32619 (N_32619,N_32244,N_32195);
xor U32620 (N_32620,N_32346,N_32489);
or U32621 (N_32621,N_32391,N_32361);
nor U32622 (N_32622,N_32315,N_32389);
nand U32623 (N_32623,N_32155,N_32084);
nand U32624 (N_32624,N_32303,N_32449);
or U32625 (N_32625,N_32318,N_32442);
and U32626 (N_32626,N_32413,N_32257);
or U32627 (N_32627,N_32085,N_32196);
nor U32628 (N_32628,N_32376,N_32447);
nand U32629 (N_32629,N_32126,N_32365);
and U32630 (N_32630,N_32073,N_32289);
or U32631 (N_32631,N_32288,N_32241);
and U32632 (N_32632,N_32226,N_32443);
xnor U32633 (N_32633,N_32448,N_32340);
and U32634 (N_32634,N_32352,N_32265);
or U32635 (N_32635,N_32411,N_32403);
nor U32636 (N_32636,N_32451,N_32016);
or U32637 (N_32637,N_32308,N_32372);
nand U32638 (N_32638,N_32248,N_32385);
and U32639 (N_32639,N_32327,N_32247);
and U32640 (N_32640,N_32334,N_32091);
xor U32641 (N_32641,N_32463,N_32331);
and U32642 (N_32642,N_32312,N_32452);
nor U32643 (N_32643,N_32136,N_32349);
nand U32644 (N_32644,N_32086,N_32162);
nand U32645 (N_32645,N_32237,N_32428);
xnor U32646 (N_32646,N_32269,N_32066);
nand U32647 (N_32647,N_32056,N_32441);
or U32648 (N_32648,N_32305,N_32273);
xor U32649 (N_32649,N_32284,N_32057);
xor U32650 (N_32650,N_32378,N_32225);
xnor U32651 (N_32651,N_32253,N_32464);
or U32652 (N_32652,N_32088,N_32182);
or U32653 (N_32653,N_32336,N_32212);
nand U32654 (N_32654,N_32425,N_32316);
xor U32655 (N_32655,N_32100,N_32138);
or U32656 (N_32656,N_32008,N_32256);
and U32657 (N_32657,N_32239,N_32296);
xnor U32658 (N_32658,N_32102,N_32032);
or U32659 (N_32659,N_32190,N_32223);
xnor U32660 (N_32660,N_32193,N_32052);
and U32661 (N_32661,N_32281,N_32049);
xor U32662 (N_32662,N_32221,N_32142);
nor U32663 (N_32663,N_32323,N_32218);
or U32664 (N_32664,N_32135,N_32387);
xnor U32665 (N_32665,N_32285,N_32460);
or U32666 (N_32666,N_32227,N_32141);
nand U32667 (N_32667,N_32246,N_32427);
xor U32668 (N_32668,N_32252,N_32202);
or U32669 (N_32669,N_32335,N_32291);
nand U32670 (N_32670,N_32401,N_32214);
nor U32671 (N_32671,N_32220,N_32328);
or U32672 (N_32672,N_32034,N_32434);
and U32673 (N_32673,N_32270,N_32398);
and U32674 (N_32674,N_32014,N_32261);
nand U32675 (N_32675,N_32341,N_32278);
nor U32676 (N_32676,N_32153,N_32233);
nor U32677 (N_32677,N_32083,N_32022);
and U32678 (N_32678,N_32475,N_32145);
nand U32679 (N_32679,N_32061,N_32228);
nand U32680 (N_32680,N_32324,N_32491);
or U32681 (N_32681,N_32367,N_32071);
and U32682 (N_32682,N_32070,N_32490);
xnor U32683 (N_32683,N_32263,N_32149);
xor U32684 (N_32684,N_32051,N_32189);
or U32685 (N_32685,N_32106,N_32095);
and U32686 (N_32686,N_32368,N_32018);
nand U32687 (N_32687,N_32059,N_32002);
or U32688 (N_32688,N_32124,N_32132);
and U32689 (N_32689,N_32069,N_32045);
and U32690 (N_32690,N_32154,N_32371);
and U32691 (N_32691,N_32161,N_32031);
nor U32692 (N_32692,N_32358,N_32147);
xnor U32693 (N_32693,N_32151,N_32280);
xor U32694 (N_32694,N_32160,N_32087);
xnor U32695 (N_32695,N_32207,N_32110);
or U32696 (N_32696,N_32180,N_32062);
nand U32697 (N_32697,N_32465,N_32118);
xor U32698 (N_32698,N_32419,N_32494);
and U32699 (N_32699,N_32362,N_32109);
xor U32700 (N_32700,N_32276,N_32146);
xor U32701 (N_32701,N_32167,N_32293);
nand U32702 (N_32702,N_32379,N_32012);
nor U32703 (N_32703,N_32231,N_32473);
nor U32704 (N_32704,N_32010,N_32445);
nand U32705 (N_32705,N_32321,N_32420);
nor U32706 (N_32706,N_32186,N_32183);
nor U32707 (N_32707,N_32024,N_32104);
and U32708 (N_32708,N_32488,N_32299);
nand U32709 (N_32709,N_32173,N_32019);
xnor U32710 (N_32710,N_32493,N_32364);
nor U32711 (N_32711,N_32410,N_32498);
nor U32712 (N_32712,N_32433,N_32048);
nor U32713 (N_32713,N_32140,N_32120);
or U32714 (N_32714,N_32353,N_32130);
nand U32715 (N_32715,N_32306,N_32359);
and U32716 (N_32716,N_32229,N_32238);
nand U32717 (N_32717,N_32450,N_32314);
nor U32718 (N_32718,N_32395,N_32007);
nor U32719 (N_32719,N_32148,N_32351);
nand U32720 (N_32720,N_32157,N_32275);
nor U32721 (N_32721,N_32243,N_32446);
and U32722 (N_32722,N_32075,N_32234);
and U32723 (N_32723,N_32068,N_32027);
and U32724 (N_32724,N_32194,N_32453);
and U32725 (N_32725,N_32242,N_32421);
nor U32726 (N_32726,N_32430,N_32435);
or U32727 (N_32727,N_32345,N_32300);
and U32728 (N_32728,N_32283,N_32041);
nor U32729 (N_32729,N_32215,N_32416);
or U32730 (N_32730,N_32399,N_32480);
nand U32731 (N_32731,N_32472,N_32459);
nor U32732 (N_32732,N_32116,N_32165);
nand U32733 (N_32733,N_32309,N_32382);
nand U32734 (N_32734,N_32105,N_32258);
or U32735 (N_32735,N_32111,N_32267);
nand U32736 (N_32736,N_32137,N_32405);
nand U32737 (N_32737,N_32197,N_32319);
xnor U32738 (N_32738,N_32444,N_32208);
and U32739 (N_32739,N_32266,N_32092);
and U32740 (N_32740,N_32426,N_32302);
nor U32741 (N_32741,N_32344,N_32046);
or U32742 (N_32742,N_32015,N_32115);
or U32743 (N_32743,N_32337,N_32081);
nand U32744 (N_32744,N_32354,N_32200);
or U32745 (N_32745,N_32392,N_32310);
nor U32746 (N_32746,N_32400,N_32169);
and U32747 (N_32747,N_32380,N_32217);
xor U32748 (N_32748,N_32178,N_32035);
nor U32749 (N_32749,N_32322,N_32470);
nor U32750 (N_32750,N_32452,N_32118);
or U32751 (N_32751,N_32274,N_32011);
nand U32752 (N_32752,N_32345,N_32125);
nand U32753 (N_32753,N_32138,N_32041);
xnor U32754 (N_32754,N_32437,N_32213);
and U32755 (N_32755,N_32041,N_32218);
and U32756 (N_32756,N_32198,N_32253);
xnor U32757 (N_32757,N_32134,N_32230);
nor U32758 (N_32758,N_32091,N_32243);
nand U32759 (N_32759,N_32083,N_32107);
or U32760 (N_32760,N_32200,N_32385);
xnor U32761 (N_32761,N_32324,N_32081);
nand U32762 (N_32762,N_32038,N_32497);
nor U32763 (N_32763,N_32491,N_32382);
xor U32764 (N_32764,N_32388,N_32351);
nand U32765 (N_32765,N_32373,N_32078);
xor U32766 (N_32766,N_32405,N_32218);
nand U32767 (N_32767,N_32036,N_32027);
or U32768 (N_32768,N_32002,N_32397);
and U32769 (N_32769,N_32111,N_32044);
xor U32770 (N_32770,N_32263,N_32352);
nand U32771 (N_32771,N_32026,N_32316);
and U32772 (N_32772,N_32483,N_32107);
nand U32773 (N_32773,N_32022,N_32473);
and U32774 (N_32774,N_32357,N_32137);
or U32775 (N_32775,N_32261,N_32224);
or U32776 (N_32776,N_32215,N_32134);
nand U32777 (N_32777,N_32399,N_32285);
nor U32778 (N_32778,N_32063,N_32075);
or U32779 (N_32779,N_32217,N_32465);
and U32780 (N_32780,N_32208,N_32073);
xor U32781 (N_32781,N_32339,N_32226);
and U32782 (N_32782,N_32238,N_32398);
nor U32783 (N_32783,N_32283,N_32070);
nor U32784 (N_32784,N_32295,N_32284);
nand U32785 (N_32785,N_32224,N_32035);
nand U32786 (N_32786,N_32054,N_32072);
nor U32787 (N_32787,N_32311,N_32397);
xnor U32788 (N_32788,N_32089,N_32298);
nand U32789 (N_32789,N_32357,N_32245);
or U32790 (N_32790,N_32090,N_32031);
and U32791 (N_32791,N_32229,N_32060);
or U32792 (N_32792,N_32339,N_32050);
xnor U32793 (N_32793,N_32308,N_32118);
nor U32794 (N_32794,N_32026,N_32036);
and U32795 (N_32795,N_32145,N_32191);
and U32796 (N_32796,N_32325,N_32076);
nor U32797 (N_32797,N_32063,N_32267);
or U32798 (N_32798,N_32033,N_32276);
xor U32799 (N_32799,N_32250,N_32089);
nor U32800 (N_32800,N_32320,N_32318);
or U32801 (N_32801,N_32209,N_32051);
and U32802 (N_32802,N_32462,N_32261);
nand U32803 (N_32803,N_32083,N_32389);
nand U32804 (N_32804,N_32230,N_32115);
or U32805 (N_32805,N_32210,N_32173);
nand U32806 (N_32806,N_32205,N_32386);
nor U32807 (N_32807,N_32242,N_32299);
or U32808 (N_32808,N_32456,N_32446);
and U32809 (N_32809,N_32374,N_32415);
nand U32810 (N_32810,N_32016,N_32414);
and U32811 (N_32811,N_32278,N_32445);
and U32812 (N_32812,N_32290,N_32114);
nor U32813 (N_32813,N_32259,N_32379);
or U32814 (N_32814,N_32286,N_32115);
and U32815 (N_32815,N_32090,N_32052);
nor U32816 (N_32816,N_32303,N_32271);
and U32817 (N_32817,N_32204,N_32330);
nor U32818 (N_32818,N_32156,N_32097);
nor U32819 (N_32819,N_32419,N_32491);
and U32820 (N_32820,N_32402,N_32366);
xor U32821 (N_32821,N_32182,N_32196);
nand U32822 (N_32822,N_32131,N_32255);
or U32823 (N_32823,N_32247,N_32417);
and U32824 (N_32824,N_32031,N_32003);
nor U32825 (N_32825,N_32334,N_32190);
or U32826 (N_32826,N_32289,N_32147);
nor U32827 (N_32827,N_32434,N_32407);
and U32828 (N_32828,N_32467,N_32324);
or U32829 (N_32829,N_32208,N_32280);
xnor U32830 (N_32830,N_32026,N_32240);
nor U32831 (N_32831,N_32236,N_32432);
nand U32832 (N_32832,N_32297,N_32122);
nor U32833 (N_32833,N_32370,N_32254);
or U32834 (N_32834,N_32085,N_32146);
nand U32835 (N_32835,N_32443,N_32187);
nand U32836 (N_32836,N_32163,N_32455);
and U32837 (N_32837,N_32498,N_32258);
and U32838 (N_32838,N_32176,N_32182);
nand U32839 (N_32839,N_32258,N_32319);
xnor U32840 (N_32840,N_32095,N_32129);
nand U32841 (N_32841,N_32393,N_32241);
and U32842 (N_32842,N_32014,N_32451);
nand U32843 (N_32843,N_32030,N_32126);
xor U32844 (N_32844,N_32483,N_32448);
xor U32845 (N_32845,N_32498,N_32163);
or U32846 (N_32846,N_32447,N_32495);
or U32847 (N_32847,N_32232,N_32023);
xor U32848 (N_32848,N_32016,N_32153);
nand U32849 (N_32849,N_32414,N_32151);
nor U32850 (N_32850,N_32173,N_32156);
and U32851 (N_32851,N_32451,N_32447);
nand U32852 (N_32852,N_32041,N_32073);
xnor U32853 (N_32853,N_32297,N_32081);
nor U32854 (N_32854,N_32272,N_32033);
nor U32855 (N_32855,N_32489,N_32235);
xor U32856 (N_32856,N_32182,N_32303);
nand U32857 (N_32857,N_32268,N_32332);
or U32858 (N_32858,N_32268,N_32214);
or U32859 (N_32859,N_32046,N_32053);
nand U32860 (N_32860,N_32260,N_32174);
xor U32861 (N_32861,N_32374,N_32248);
nor U32862 (N_32862,N_32193,N_32209);
xnor U32863 (N_32863,N_32458,N_32456);
or U32864 (N_32864,N_32383,N_32327);
or U32865 (N_32865,N_32319,N_32478);
and U32866 (N_32866,N_32119,N_32281);
xor U32867 (N_32867,N_32274,N_32042);
xor U32868 (N_32868,N_32054,N_32113);
xor U32869 (N_32869,N_32222,N_32488);
nor U32870 (N_32870,N_32132,N_32470);
or U32871 (N_32871,N_32022,N_32210);
nor U32872 (N_32872,N_32342,N_32020);
xor U32873 (N_32873,N_32377,N_32309);
or U32874 (N_32874,N_32310,N_32499);
and U32875 (N_32875,N_32473,N_32044);
nand U32876 (N_32876,N_32302,N_32425);
and U32877 (N_32877,N_32498,N_32102);
or U32878 (N_32878,N_32036,N_32035);
nor U32879 (N_32879,N_32472,N_32288);
nand U32880 (N_32880,N_32120,N_32436);
xnor U32881 (N_32881,N_32131,N_32321);
xnor U32882 (N_32882,N_32423,N_32126);
xor U32883 (N_32883,N_32295,N_32317);
or U32884 (N_32884,N_32248,N_32147);
xnor U32885 (N_32885,N_32126,N_32221);
or U32886 (N_32886,N_32433,N_32103);
xor U32887 (N_32887,N_32363,N_32307);
nand U32888 (N_32888,N_32040,N_32482);
xnor U32889 (N_32889,N_32279,N_32396);
nand U32890 (N_32890,N_32041,N_32326);
and U32891 (N_32891,N_32446,N_32391);
and U32892 (N_32892,N_32416,N_32424);
nand U32893 (N_32893,N_32206,N_32439);
nand U32894 (N_32894,N_32115,N_32032);
and U32895 (N_32895,N_32408,N_32306);
or U32896 (N_32896,N_32463,N_32237);
nand U32897 (N_32897,N_32259,N_32403);
nor U32898 (N_32898,N_32439,N_32123);
and U32899 (N_32899,N_32133,N_32224);
and U32900 (N_32900,N_32287,N_32009);
nand U32901 (N_32901,N_32409,N_32147);
nand U32902 (N_32902,N_32367,N_32102);
and U32903 (N_32903,N_32383,N_32192);
nand U32904 (N_32904,N_32006,N_32352);
nand U32905 (N_32905,N_32475,N_32130);
and U32906 (N_32906,N_32175,N_32221);
nand U32907 (N_32907,N_32100,N_32113);
and U32908 (N_32908,N_32062,N_32258);
nand U32909 (N_32909,N_32387,N_32277);
nand U32910 (N_32910,N_32200,N_32125);
xor U32911 (N_32911,N_32235,N_32334);
nor U32912 (N_32912,N_32312,N_32276);
xor U32913 (N_32913,N_32106,N_32150);
and U32914 (N_32914,N_32069,N_32089);
xnor U32915 (N_32915,N_32095,N_32080);
or U32916 (N_32916,N_32270,N_32113);
and U32917 (N_32917,N_32477,N_32234);
nor U32918 (N_32918,N_32388,N_32035);
or U32919 (N_32919,N_32085,N_32313);
or U32920 (N_32920,N_32219,N_32479);
xor U32921 (N_32921,N_32391,N_32131);
nor U32922 (N_32922,N_32366,N_32054);
xnor U32923 (N_32923,N_32384,N_32483);
nand U32924 (N_32924,N_32190,N_32002);
nand U32925 (N_32925,N_32399,N_32052);
and U32926 (N_32926,N_32211,N_32047);
xor U32927 (N_32927,N_32488,N_32434);
and U32928 (N_32928,N_32295,N_32473);
and U32929 (N_32929,N_32400,N_32066);
xnor U32930 (N_32930,N_32241,N_32047);
and U32931 (N_32931,N_32307,N_32443);
and U32932 (N_32932,N_32307,N_32287);
nor U32933 (N_32933,N_32159,N_32221);
xor U32934 (N_32934,N_32342,N_32468);
xor U32935 (N_32935,N_32382,N_32245);
nand U32936 (N_32936,N_32389,N_32386);
and U32937 (N_32937,N_32233,N_32038);
nor U32938 (N_32938,N_32001,N_32358);
and U32939 (N_32939,N_32254,N_32297);
or U32940 (N_32940,N_32496,N_32373);
nand U32941 (N_32941,N_32071,N_32085);
and U32942 (N_32942,N_32304,N_32166);
nor U32943 (N_32943,N_32324,N_32142);
and U32944 (N_32944,N_32326,N_32458);
nor U32945 (N_32945,N_32046,N_32028);
nor U32946 (N_32946,N_32029,N_32447);
or U32947 (N_32947,N_32174,N_32312);
nand U32948 (N_32948,N_32415,N_32020);
nor U32949 (N_32949,N_32304,N_32246);
nor U32950 (N_32950,N_32056,N_32329);
xor U32951 (N_32951,N_32152,N_32228);
or U32952 (N_32952,N_32056,N_32233);
and U32953 (N_32953,N_32057,N_32475);
xor U32954 (N_32954,N_32023,N_32438);
and U32955 (N_32955,N_32368,N_32330);
xnor U32956 (N_32956,N_32218,N_32077);
nor U32957 (N_32957,N_32085,N_32188);
nor U32958 (N_32958,N_32039,N_32240);
nor U32959 (N_32959,N_32474,N_32069);
xor U32960 (N_32960,N_32410,N_32303);
or U32961 (N_32961,N_32043,N_32076);
nand U32962 (N_32962,N_32152,N_32424);
nand U32963 (N_32963,N_32455,N_32419);
or U32964 (N_32964,N_32071,N_32448);
and U32965 (N_32965,N_32432,N_32139);
and U32966 (N_32966,N_32302,N_32360);
or U32967 (N_32967,N_32188,N_32149);
or U32968 (N_32968,N_32429,N_32436);
nand U32969 (N_32969,N_32335,N_32208);
and U32970 (N_32970,N_32186,N_32331);
nand U32971 (N_32971,N_32400,N_32154);
nor U32972 (N_32972,N_32401,N_32191);
xnor U32973 (N_32973,N_32381,N_32158);
or U32974 (N_32974,N_32067,N_32010);
nand U32975 (N_32975,N_32334,N_32498);
nor U32976 (N_32976,N_32317,N_32283);
nor U32977 (N_32977,N_32203,N_32195);
or U32978 (N_32978,N_32018,N_32404);
nor U32979 (N_32979,N_32342,N_32211);
and U32980 (N_32980,N_32420,N_32014);
nand U32981 (N_32981,N_32086,N_32294);
or U32982 (N_32982,N_32014,N_32377);
xor U32983 (N_32983,N_32215,N_32224);
nor U32984 (N_32984,N_32157,N_32394);
nand U32985 (N_32985,N_32198,N_32438);
and U32986 (N_32986,N_32235,N_32385);
nand U32987 (N_32987,N_32203,N_32078);
or U32988 (N_32988,N_32319,N_32104);
xnor U32989 (N_32989,N_32099,N_32468);
and U32990 (N_32990,N_32127,N_32259);
and U32991 (N_32991,N_32313,N_32357);
or U32992 (N_32992,N_32338,N_32465);
nand U32993 (N_32993,N_32424,N_32207);
nor U32994 (N_32994,N_32280,N_32091);
and U32995 (N_32995,N_32088,N_32087);
nand U32996 (N_32996,N_32125,N_32394);
and U32997 (N_32997,N_32007,N_32261);
xnor U32998 (N_32998,N_32499,N_32390);
nand U32999 (N_32999,N_32411,N_32027);
xnor U33000 (N_33000,N_32821,N_32852);
xnor U33001 (N_33001,N_32938,N_32587);
xnor U33002 (N_33002,N_32675,N_32897);
or U33003 (N_33003,N_32997,N_32905);
nand U33004 (N_33004,N_32509,N_32971);
and U33005 (N_33005,N_32985,N_32607);
xnor U33006 (N_33006,N_32686,N_32989);
or U33007 (N_33007,N_32708,N_32809);
xor U33008 (N_33008,N_32755,N_32746);
and U33009 (N_33009,N_32858,N_32593);
xor U33010 (N_33010,N_32550,N_32830);
xor U33011 (N_33011,N_32653,N_32690);
or U33012 (N_33012,N_32518,N_32964);
nor U33013 (N_33013,N_32854,N_32887);
and U33014 (N_33014,N_32707,N_32720);
nand U33015 (N_33015,N_32669,N_32974);
and U33016 (N_33016,N_32867,N_32959);
nand U33017 (N_33017,N_32922,N_32912);
nand U33018 (N_33018,N_32845,N_32898);
xnor U33019 (N_33019,N_32967,N_32694);
nor U33020 (N_33020,N_32711,N_32975);
and U33021 (N_33021,N_32635,N_32716);
xnor U33022 (N_33022,N_32725,N_32535);
or U33023 (N_33023,N_32642,N_32512);
xnor U33024 (N_33024,N_32882,N_32949);
nand U33025 (N_33025,N_32981,N_32689);
nand U33026 (N_33026,N_32552,N_32870);
and U33027 (N_33027,N_32932,N_32778);
or U33028 (N_33028,N_32775,N_32818);
xnor U33029 (N_33029,N_32968,N_32822);
or U33030 (N_33030,N_32749,N_32637);
nand U33031 (N_33031,N_32978,N_32756);
nand U33032 (N_33032,N_32874,N_32754);
xor U33033 (N_33033,N_32914,N_32526);
or U33034 (N_33034,N_32947,N_32761);
or U33035 (N_33035,N_32666,N_32534);
nand U33036 (N_33036,N_32737,N_32643);
nor U33037 (N_33037,N_32929,N_32983);
nand U33038 (N_33038,N_32957,N_32931);
and U33039 (N_33039,N_32736,N_32780);
or U33040 (N_33040,N_32621,N_32656);
nor U33041 (N_33041,N_32941,N_32727);
xnor U33042 (N_33042,N_32561,N_32895);
nand U33043 (N_33043,N_32995,N_32565);
and U33044 (N_33044,N_32699,N_32814);
and U33045 (N_33045,N_32551,N_32815);
xor U33046 (N_33046,N_32976,N_32702);
nor U33047 (N_33047,N_32906,N_32612);
and U33048 (N_33048,N_32624,N_32663);
nand U33049 (N_33049,N_32794,N_32641);
nor U33050 (N_33050,N_32576,N_32626);
and U33051 (N_33051,N_32970,N_32730);
xor U33052 (N_33052,N_32659,N_32807);
and U33053 (N_33053,N_32980,N_32903);
nand U33054 (N_33054,N_32578,N_32573);
or U33055 (N_33055,N_32577,N_32951);
xnor U33056 (N_33056,N_32881,N_32705);
xnor U33057 (N_33057,N_32523,N_32984);
nor U33058 (N_33058,N_32937,N_32793);
xor U33059 (N_33059,N_32602,N_32800);
xor U33060 (N_33060,N_32942,N_32605);
and U33061 (N_33061,N_32998,N_32836);
nor U33062 (N_33062,N_32560,N_32734);
or U33063 (N_33063,N_32660,N_32664);
nand U33064 (N_33064,N_32779,N_32839);
xnor U33065 (N_33065,N_32876,N_32961);
xnor U33066 (N_33066,N_32559,N_32851);
nand U33067 (N_33067,N_32528,N_32955);
xnor U33068 (N_33068,N_32501,N_32553);
nand U33069 (N_33069,N_32927,N_32894);
nor U33070 (N_33070,N_32585,N_32884);
or U33071 (N_33071,N_32634,N_32525);
nor U33072 (N_33072,N_32652,N_32787);
nand U33073 (N_33073,N_32805,N_32703);
nor U33074 (N_33074,N_32855,N_32685);
nand U33075 (N_33075,N_32570,N_32783);
or U33076 (N_33076,N_32540,N_32748);
or U33077 (N_33077,N_32522,N_32714);
xor U33078 (N_33078,N_32917,N_32670);
or U33079 (N_33079,N_32994,N_32798);
or U33080 (N_33080,N_32722,N_32549);
xnor U33081 (N_33081,N_32788,N_32568);
or U33082 (N_33082,N_32524,N_32806);
nor U33083 (N_33083,N_32883,N_32682);
and U33084 (N_33084,N_32519,N_32655);
or U33085 (N_33085,N_32515,N_32517);
or U33086 (N_33086,N_32902,N_32674);
nor U33087 (N_33087,N_32963,N_32604);
or U33088 (N_33088,N_32557,N_32592);
xnor U33089 (N_33089,N_32763,N_32996);
nor U33090 (N_33090,N_32766,N_32547);
or U33091 (N_33091,N_32583,N_32594);
nor U33092 (N_33092,N_32796,N_32657);
or U33093 (N_33093,N_32733,N_32639);
or U33094 (N_33094,N_32662,N_32507);
xor U33095 (N_33095,N_32891,N_32511);
nand U33096 (N_33096,N_32960,N_32786);
nand U33097 (N_33097,N_32841,N_32740);
nand U33098 (N_33098,N_32582,N_32923);
nand U33099 (N_33099,N_32622,N_32530);
xor U33100 (N_33100,N_32908,N_32834);
or U33101 (N_33101,N_32833,N_32772);
nand U33102 (N_33102,N_32829,N_32958);
nand U33103 (N_33103,N_32606,N_32965);
or U33104 (N_33104,N_32926,N_32948);
or U33105 (N_33105,N_32972,N_32599);
nand U33106 (N_33106,N_32679,N_32513);
xnor U33107 (N_33107,N_32886,N_32930);
or U33108 (N_33108,N_32979,N_32673);
xor U33109 (N_33109,N_32828,N_32591);
xor U33110 (N_33110,N_32514,N_32724);
xor U33111 (N_33111,N_32849,N_32645);
nand U33112 (N_33112,N_32777,N_32795);
nor U33113 (N_33113,N_32668,N_32921);
and U33114 (N_33114,N_32747,N_32567);
and U33115 (N_33115,N_32885,N_32562);
nor U33116 (N_33116,N_32899,N_32860);
or U33117 (N_33117,N_32584,N_32677);
or U33118 (N_33118,N_32610,N_32596);
and U33119 (N_33119,N_32878,N_32700);
and U33120 (N_33120,N_32840,N_32545);
nor U33121 (N_33121,N_32789,N_32865);
nand U33122 (N_33122,N_32799,N_32910);
and U33123 (N_33123,N_32817,N_32623);
or U33124 (N_33124,N_32993,N_32676);
nand U33125 (N_33125,N_32629,N_32940);
or U33126 (N_33126,N_32712,N_32919);
nor U33127 (N_33127,N_32719,N_32857);
nor U33128 (N_33128,N_32757,N_32539);
nor U33129 (N_33129,N_32521,N_32658);
xor U33130 (N_33130,N_32717,N_32811);
and U33131 (N_33131,N_32632,N_32832);
nand U33132 (N_33132,N_32618,N_32684);
nor U33133 (N_33133,N_32579,N_32536);
xnor U33134 (N_33134,N_32880,N_32743);
and U33135 (N_33135,N_32558,N_32826);
or U33136 (N_33136,N_32548,N_32866);
xnor U33137 (N_33137,N_32531,N_32896);
nor U33138 (N_33138,N_32864,N_32850);
xor U33139 (N_33139,N_32750,N_32603);
and U33140 (N_33140,N_32619,N_32966);
nor U33141 (N_33141,N_32802,N_32544);
or U33142 (N_33142,N_32831,N_32742);
and U33143 (N_33143,N_32934,N_32546);
nand U33144 (N_33144,N_32868,N_32769);
and U33145 (N_33145,N_32782,N_32933);
or U33146 (N_33146,N_32647,N_32827);
or U33147 (N_33147,N_32500,N_32628);
and U33148 (N_33148,N_32566,N_32973);
nor U33149 (N_33149,N_32991,N_32680);
and U33150 (N_33150,N_32752,N_32726);
xor U33151 (N_33151,N_32649,N_32729);
xnor U33152 (N_33152,N_32890,N_32879);
and U33153 (N_33153,N_32999,N_32542);
xor U33154 (N_33154,N_32556,N_32687);
and U33155 (N_33155,N_32510,N_32872);
nor U33156 (N_33156,N_32835,N_32928);
or U33157 (N_33157,N_32801,N_32693);
nor U33158 (N_33158,N_32816,N_32581);
and U33159 (N_33159,N_32665,N_32848);
nand U33160 (N_33160,N_32590,N_32913);
or U33161 (N_33161,N_32751,N_32838);
and U33162 (N_33162,N_32861,N_32698);
nor U33163 (N_33163,N_32696,N_32631);
nor U33164 (N_33164,N_32554,N_32900);
xor U33165 (N_33165,N_32555,N_32586);
or U33166 (N_33166,N_32721,N_32810);
nor U33167 (N_33167,N_32875,N_32907);
and U33168 (N_33168,N_32580,N_32744);
or U33169 (N_33169,N_32695,N_32506);
and U33170 (N_33170,N_32633,N_32505);
nor U33171 (N_33171,N_32701,N_32681);
and U33172 (N_33172,N_32538,N_32767);
nor U33173 (N_33173,N_32646,N_32889);
or U33174 (N_33174,N_32797,N_32946);
nor U33175 (N_33175,N_32600,N_32837);
xor U33176 (N_33176,N_32503,N_32638);
and U33177 (N_33177,N_32819,N_32601);
and U33178 (N_33178,N_32723,N_32574);
and U33179 (N_33179,N_32823,N_32785);
xor U33180 (N_33180,N_32732,N_32630);
and U33181 (N_33181,N_32710,N_32758);
xnor U33182 (N_33182,N_32651,N_32564);
nand U33183 (N_33183,N_32715,N_32532);
nor U33184 (N_33184,N_32648,N_32920);
xor U33185 (N_33185,N_32842,N_32944);
nor U33186 (N_33186,N_32697,N_32969);
nand U33187 (N_33187,N_32936,N_32768);
and U33188 (N_33188,N_32853,N_32589);
nor U33189 (N_33189,N_32713,N_32988);
nor U33190 (N_33190,N_32892,N_32611);
nor U33191 (N_33191,N_32625,N_32950);
xor U33192 (N_33192,N_32654,N_32911);
and U33193 (N_33193,N_32871,N_32706);
nor U33194 (N_33194,N_32987,N_32945);
or U33195 (N_33195,N_32924,N_32925);
nor U33196 (N_33196,N_32533,N_32990);
nor U33197 (N_33197,N_32986,N_32667);
xnor U33198 (N_33198,N_32943,N_32962);
xnor U33199 (N_33199,N_32620,N_32543);
and U33200 (N_33200,N_32846,N_32537);
nand U33201 (N_33201,N_32615,N_32644);
nand U33202 (N_33202,N_32597,N_32953);
and U33203 (N_33203,N_32508,N_32909);
nand U33204 (N_33204,N_32728,N_32901);
and U33205 (N_33205,N_32863,N_32709);
or U33206 (N_33206,N_32640,N_32731);
nand U33207 (N_33207,N_32765,N_32627);
or U33208 (N_33208,N_32753,N_32764);
or U33209 (N_33209,N_32650,N_32844);
or U33210 (N_33210,N_32824,N_32563);
nor U33211 (N_33211,N_32572,N_32843);
nand U33212 (N_33212,N_32575,N_32738);
nor U33213 (N_33213,N_32862,N_32762);
xnor U33214 (N_33214,N_32672,N_32784);
and U33215 (N_33215,N_32893,N_32718);
and U33216 (N_33216,N_32571,N_32688);
and U33217 (N_33217,N_32877,N_32588);
nand U33218 (N_33218,N_32790,N_32598);
nor U33219 (N_33219,N_32520,N_32502);
or U33220 (N_33220,N_32792,N_32859);
nor U33221 (N_33221,N_32992,N_32954);
nor U33222 (N_33222,N_32616,N_32812);
nand U33223 (N_33223,N_32569,N_32504);
or U33224 (N_33224,N_32856,N_32678);
nand U33225 (N_33225,N_32683,N_32661);
nor U33226 (N_33226,N_32741,N_32541);
and U33227 (N_33227,N_32771,N_32760);
nor U33228 (N_33228,N_32952,N_32608);
nor U33229 (N_33229,N_32825,N_32691);
nor U33230 (N_33230,N_32617,N_32774);
nand U33231 (N_33231,N_32904,N_32636);
or U33232 (N_33232,N_32529,N_32804);
and U33233 (N_33233,N_32803,N_32915);
and U33234 (N_33234,N_32791,N_32759);
nand U33235 (N_33235,N_32692,N_32956);
nand U33236 (N_33236,N_32773,N_32781);
and U33237 (N_33237,N_32847,N_32813);
nor U33238 (N_33238,N_32671,N_32939);
nor U33239 (N_33239,N_32770,N_32739);
xnor U33240 (N_33240,N_32745,N_32595);
or U33241 (N_33241,N_32609,N_32527);
and U33242 (N_33242,N_32888,N_32869);
or U33243 (N_33243,N_32704,N_32918);
nor U33244 (N_33244,N_32613,N_32935);
and U33245 (N_33245,N_32982,N_32735);
or U33246 (N_33246,N_32820,N_32873);
nand U33247 (N_33247,N_32776,N_32516);
xor U33248 (N_33248,N_32977,N_32614);
and U33249 (N_33249,N_32808,N_32916);
or U33250 (N_33250,N_32829,N_32520);
nor U33251 (N_33251,N_32561,N_32673);
or U33252 (N_33252,N_32854,N_32576);
and U33253 (N_33253,N_32917,N_32961);
nor U33254 (N_33254,N_32501,N_32532);
nand U33255 (N_33255,N_32783,N_32825);
xor U33256 (N_33256,N_32518,N_32849);
xor U33257 (N_33257,N_32528,N_32974);
xor U33258 (N_33258,N_32927,N_32718);
nand U33259 (N_33259,N_32691,N_32603);
nand U33260 (N_33260,N_32945,N_32882);
nand U33261 (N_33261,N_32535,N_32540);
xnor U33262 (N_33262,N_32668,N_32998);
nor U33263 (N_33263,N_32924,N_32571);
nand U33264 (N_33264,N_32790,N_32986);
or U33265 (N_33265,N_32870,N_32816);
xor U33266 (N_33266,N_32665,N_32702);
xnor U33267 (N_33267,N_32711,N_32594);
and U33268 (N_33268,N_32554,N_32814);
nor U33269 (N_33269,N_32600,N_32726);
nand U33270 (N_33270,N_32747,N_32891);
nand U33271 (N_33271,N_32725,N_32994);
nor U33272 (N_33272,N_32733,N_32658);
nand U33273 (N_33273,N_32665,N_32854);
nand U33274 (N_33274,N_32827,N_32532);
nand U33275 (N_33275,N_32913,N_32983);
and U33276 (N_33276,N_32653,N_32598);
and U33277 (N_33277,N_32899,N_32830);
or U33278 (N_33278,N_32532,N_32888);
or U33279 (N_33279,N_32714,N_32965);
nand U33280 (N_33280,N_32718,N_32539);
xor U33281 (N_33281,N_32776,N_32687);
or U33282 (N_33282,N_32618,N_32992);
xnor U33283 (N_33283,N_32910,N_32576);
or U33284 (N_33284,N_32642,N_32944);
nand U33285 (N_33285,N_32947,N_32818);
nand U33286 (N_33286,N_32800,N_32544);
xnor U33287 (N_33287,N_32535,N_32964);
nand U33288 (N_33288,N_32546,N_32592);
or U33289 (N_33289,N_32929,N_32641);
xor U33290 (N_33290,N_32604,N_32560);
nand U33291 (N_33291,N_32512,N_32567);
nor U33292 (N_33292,N_32627,N_32815);
or U33293 (N_33293,N_32992,N_32700);
nand U33294 (N_33294,N_32627,N_32513);
xor U33295 (N_33295,N_32870,N_32955);
and U33296 (N_33296,N_32711,N_32586);
nand U33297 (N_33297,N_32755,N_32729);
xnor U33298 (N_33298,N_32547,N_32979);
nand U33299 (N_33299,N_32772,N_32995);
nand U33300 (N_33300,N_32683,N_32707);
nor U33301 (N_33301,N_32625,N_32517);
or U33302 (N_33302,N_32626,N_32888);
or U33303 (N_33303,N_32716,N_32925);
and U33304 (N_33304,N_32644,N_32871);
and U33305 (N_33305,N_32898,N_32872);
and U33306 (N_33306,N_32932,N_32801);
nand U33307 (N_33307,N_32950,N_32586);
nor U33308 (N_33308,N_32895,N_32962);
xor U33309 (N_33309,N_32524,N_32550);
nand U33310 (N_33310,N_32965,N_32545);
nand U33311 (N_33311,N_32950,N_32915);
xor U33312 (N_33312,N_32884,N_32933);
nand U33313 (N_33313,N_32834,N_32584);
xor U33314 (N_33314,N_32574,N_32524);
or U33315 (N_33315,N_32517,N_32957);
or U33316 (N_33316,N_32925,N_32756);
nor U33317 (N_33317,N_32779,N_32627);
nor U33318 (N_33318,N_32773,N_32953);
and U33319 (N_33319,N_32889,N_32977);
nor U33320 (N_33320,N_32963,N_32632);
nand U33321 (N_33321,N_32525,N_32527);
nor U33322 (N_33322,N_32714,N_32539);
xnor U33323 (N_33323,N_32982,N_32766);
nand U33324 (N_33324,N_32594,N_32980);
or U33325 (N_33325,N_32519,N_32804);
or U33326 (N_33326,N_32670,N_32612);
nand U33327 (N_33327,N_32977,N_32890);
or U33328 (N_33328,N_32548,N_32811);
nor U33329 (N_33329,N_32748,N_32812);
xnor U33330 (N_33330,N_32879,N_32672);
or U33331 (N_33331,N_32819,N_32952);
xnor U33332 (N_33332,N_32583,N_32936);
or U33333 (N_33333,N_32821,N_32632);
and U33334 (N_33334,N_32991,N_32962);
xor U33335 (N_33335,N_32623,N_32963);
and U33336 (N_33336,N_32814,N_32809);
nand U33337 (N_33337,N_32779,N_32553);
or U33338 (N_33338,N_32591,N_32624);
nand U33339 (N_33339,N_32889,N_32862);
nor U33340 (N_33340,N_32513,N_32921);
nand U33341 (N_33341,N_32623,N_32825);
and U33342 (N_33342,N_32525,N_32619);
and U33343 (N_33343,N_32757,N_32557);
nand U33344 (N_33344,N_32977,N_32715);
or U33345 (N_33345,N_32869,N_32871);
or U33346 (N_33346,N_32927,N_32708);
or U33347 (N_33347,N_32531,N_32801);
nor U33348 (N_33348,N_32668,N_32962);
nor U33349 (N_33349,N_32849,N_32803);
nand U33350 (N_33350,N_32932,N_32980);
and U33351 (N_33351,N_32867,N_32984);
xor U33352 (N_33352,N_32863,N_32618);
and U33353 (N_33353,N_32871,N_32553);
nor U33354 (N_33354,N_32552,N_32829);
nor U33355 (N_33355,N_32862,N_32627);
xnor U33356 (N_33356,N_32720,N_32952);
nor U33357 (N_33357,N_32978,N_32735);
nor U33358 (N_33358,N_32757,N_32640);
xnor U33359 (N_33359,N_32912,N_32510);
nand U33360 (N_33360,N_32950,N_32532);
xor U33361 (N_33361,N_32863,N_32786);
and U33362 (N_33362,N_32680,N_32946);
and U33363 (N_33363,N_32647,N_32563);
or U33364 (N_33364,N_32939,N_32943);
or U33365 (N_33365,N_32694,N_32818);
nand U33366 (N_33366,N_32949,N_32579);
nand U33367 (N_33367,N_32952,N_32835);
nand U33368 (N_33368,N_32544,N_32857);
xor U33369 (N_33369,N_32996,N_32805);
or U33370 (N_33370,N_32680,N_32878);
and U33371 (N_33371,N_32814,N_32898);
or U33372 (N_33372,N_32945,N_32923);
nand U33373 (N_33373,N_32716,N_32690);
nor U33374 (N_33374,N_32593,N_32807);
xor U33375 (N_33375,N_32648,N_32943);
nor U33376 (N_33376,N_32893,N_32858);
nand U33377 (N_33377,N_32727,N_32972);
xor U33378 (N_33378,N_32574,N_32611);
or U33379 (N_33379,N_32675,N_32545);
nand U33380 (N_33380,N_32566,N_32697);
nor U33381 (N_33381,N_32692,N_32537);
nand U33382 (N_33382,N_32848,N_32720);
nor U33383 (N_33383,N_32744,N_32973);
or U33384 (N_33384,N_32850,N_32655);
and U33385 (N_33385,N_32866,N_32670);
xor U33386 (N_33386,N_32723,N_32761);
and U33387 (N_33387,N_32635,N_32970);
xnor U33388 (N_33388,N_32941,N_32976);
or U33389 (N_33389,N_32567,N_32607);
nand U33390 (N_33390,N_32711,N_32527);
nor U33391 (N_33391,N_32565,N_32677);
xnor U33392 (N_33392,N_32599,N_32710);
xor U33393 (N_33393,N_32532,N_32524);
nand U33394 (N_33394,N_32835,N_32976);
nor U33395 (N_33395,N_32955,N_32646);
nand U33396 (N_33396,N_32614,N_32582);
nor U33397 (N_33397,N_32958,N_32999);
or U33398 (N_33398,N_32785,N_32984);
nor U33399 (N_33399,N_32751,N_32672);
or U33400 (N_33400,N_32799,N_32964);
or U33401 (N_33401,N_32717,N_32916);
nand U33402 (N_33402,N_32563,N_32706);
xnor U33403 (N_33403,N_32722,N_32953);
nand U33404 (N_33404,N_32616,N_32513);
or U33405 (N_33405,N_32903,N_32512);
or U33406 (N_33406,N_32946,N_32745);
or U33407 (N_33407,N_32700,N_32871);
and U33408 (N_33408,N_32996,N_32708);
xor U33409 (N_33409,N_32751,N_32629);
nand U33410 (N_33410,N_32736,N_32913);
nand U33411 (N_33411,N_32514,N_32561);
or U33412 (N_33412,N_32842,N_32947);
xor U33413 (N_33413,N_32793,N_32851);
and U33414 (N_33414,N_32777,N_32971);
and U33415 (N_33415,N_32684,N_32820);
or U33416 (N_33416,N_32716,N_32542);
xor U33417 (N_33417,N_32878,N_32704);
xnor U33418 (N_33418,N_32896,N_32940);
nor U33419 (N_33419,N_32527,N_32532);
xor U33420 (N_33420,N_32601,N_32869);
xnor U33421 (N_33421,N_32985,N_32504);
nor U33422 (N_33422,N_32772,N_32679);
and U33423 (N_33423,N_32753,N_32592);
and U33424 (N_33424,N_32792,N_32809);
nor U33425 (N_33425,N_32510,N_32700);
nand U33426 (N_33426,N_32870,N_32856);
nand U33427 (N_33427,N_32958,N_32812);
xor U33428 (N_33428,N_32558,N_32955);
xnor U33429 (N_33429,N_32602,N_32677);
nor U33430 (N_33430,N_32937,N_32714);
xor U33431 (N_33431,N_32557,N_32955);
and U33432 (N_33432,N_32604,N_32867);
nor U33433 (N_33433,N_32543,N_32769);
nor U33434 (N_33434,N_32658,N_32866);
nor U33435 (N_33435,N_32849,N_32634);
and U33436 (N_33436,N_32503,N_32627);
and U33437 (N_33437,N_32844,N_32802);
and U33438 (N_33438,N_32793,N_32520);
or U33439 (N_33439,N_32514,N_32994);
and U33440 (N_33440,N_32942,N_32853);
xnor U33441 (N_33441,N_32825,N_32881);
or U33442 (N_33442,N_32910,N_32671);
and U33443 (N_33443,N_32976,N_32713);
xnor U33444 (N_33444,N_32521,N_32532);
nor U33445 (N_33445,N_32708,N_32584);
and U33446 (N_33446,N_32639,N_32941);
nor U33447 (N_33447,N_32961,N_32539);
nand U33448 (N_33448,N_32671,N_32973);
and U33449 (N_33449,N_32588,N_32899);
nand U33450 (N_33450,N_32840,N_32547);
nand U33451 (N_33451,N_32917,N_32699);
nand U33452 (N_33452,N_32987,N_32622);
and U33453 (N_33453,N_32803,N_32726);
and U33454 (N_33454,N_32659,N_32512);
and U33455 (N_33455,N_32516,N_32945);
or U33456 (N_33456,N_32507,N_32877);
or U33457 (N_33457,N_32581,N_32604);
xnor U33458 (N_33458,N_32558,N_32679);
nor U33459 (N_33459,N_32527,N_32662);
or U33460 (N_33460,N_32879,N_32774);
nor U33461 (N_33461,N_32913,N_32713);
nor U33462 (N_33462,N_32660,N_32676);
or U33463 (N_33463,N_32828,N_32771);
nor U33464 (N_33464,N_32755,N_32926);
nor U33465 (N_33465,N_32813,N_32877);
nor U33466 (N_33466,N_32808,N_32955);
xor U33467 (N_33467,N_32790,N_32807);
and U33468 (N_33468,N_32778,N_32861);
xor U33469 (N_33469,N_32954,N_32960);
or U33470 (N_33470,N_32931,N_32986);
nor U33471 (N_33471,N_32841,N_32917);
or U33472 (N_33472,N_32907,N_32698);
nand U33473 (N_33473,N_32605,N_32790);
nand U33474 (N_33474,N_32628,N_32857);
nand U33475 (N_33475,N_32628,N_32952);
or U33476 (N_33476,N_32736,N_32841);
nor U33477 (N_33477,N_32994,N_32527);
nor U33478 (N_33478,N_32886,N_32998);
or U33479 (N_33479,N_32719,N_32890);
nor U33480 (N_33480,N_32942,N_32900);
or U33481 (N_33481,N_32585,N_32770);
nand U33482 (N_33482,N_32729,N_32646);
xnor U33483 (N_33483,N_32799,N_32716);
or U33484 (N_33484,N_32998,N_32977);
and U33485 (N_33485,N_32532,N_32910);
nand U33486 (N_33486,N_32722,N_32807);
or U33487 (N_33487,N_32564,N_32957);
and U33488 (N_33488,N_32507,N_32622);
nor U33489 (N_33489,N_32603,N_32898);
xor U33490 (N_33490,N_32762,N_32603);
xnor U33491 (N_33491,N_32896,N_32656);
and U33492 (N_33492,N_32929,N_32802);
and U33493 (N_33493,N_32931,N_32554);
nor U33494 (N_33494,N_32675,N_32571);
nor U33495 (N_33495,N_32503,N_32874);
nor U33496 (N_33496,N_32646,N_32687);
and U33497 (N_33497,N_32690,N_32853);
xor U33498 (N_33498,N_32810,N_32961);
or U33499 (N_33499,N_32639,N_32891);
or U33500 (N_33500,N_33153,N_33063);
or U33501 (N_33501,N_33358,N_33350);
xor U33502 (N_33502,N_33091,N_33206);
nand U33503 (N_33503,N_33159,N_33378);
or U33504 (N_33504,N_33347,N_33208);
and U33505 (N_33505,N_33324,N_33064);
or U33506 (N_33506,N_33038,N_33062);
and U33507 (N_33507,N_33284,N_33126);
or U33508 (N_33508,N_33454,N_33387);
and U33509 (N_33509,N_33496,N_33459);
xnor U33510 (N_33510,N_33162,N_33123);
or U33511 (N_33511,N_33109,N_33216);
xnor U33512 (N_33512,N_33340,N_33356);
and U33513 (N_33513,N_33086,N_33410);
or U33514 (N_33514,N_33453,N_33083);
or U33515 (N_33515,N_33369,N_33140);
xnor U33516 (N_33516,N_33367,N_33413);
xnor U33517 (N_33517,N_33059,N_33081);
and U33518 (N_33518,N_33499,N_33401);
xnor U33519 (N_33519,N_33327,N_33446);
nand U33520 (N_33520,N_33074,N_33136);
nor U33521 (N_33521,N_33305,N_33178);
nor U33522 (N_33522,N_33049,N_33161);
and U33523 (N_33523,N_33402,N_33285);
and U33524 (N_33524,N_33412,N_33060);
nor U33525 (N_33525,N_33095,N_33471);
xor U33526 (N_33526,N_33357,N_33498);
and U33527 (N_33527,N_33089,N_33235);
or U33528 (N_33528,N_33271,N_33295);
or U33529 (N_33529,N_33363,N_33465);
nand U33530 (N_33530,N_33112,N_33449);
nor U33531 (N_33531,N_33041,N_33335);
xnor U33532 (N_33532,N_33400,N_33272);
nor U33533 (N_33533,N_33082,N_33396);
and U33534 (N_33534,N_33328,N_33461);
nor U33535 (N_33535,N_33390,N_33468);
nand U33536 (N_33536,N_33224,N_33039);
nor U33537 (N_33537,N_33115,N_33418);
xor U33538 (N_33538,N_33462,N_33119);
or U33539 (N_33539,N_33379,N_33419);
or U33540 (N_33540,N_33194,N_33120);
or U33541 (N_33541,N_33157,N_33076);
nor U33542 (N_33542,N_33259,N_33332);
nand U33543 (N_33543,N_33096,N_33022);
and U33544 (N_33544,N_33024,N_33457);
nand U33545 (N_33545,N_33443,N_33056);
xnor U33546 (N_33546,N_33085,N_33128);
and U33547 (N_33547,N_33190,N_33210);
xor U33548 (N_33548,N_33493,N_33179);
or U33549 (N_33549,N_33051,N_33246);
or U33550 (N_33550,N_33058,N_33351);
nand U33551 (N_33551,N_33290,N_33135);
xnor U33552 (N_33552,N_33042,N_33139);
xor U33553 (N_33553,N_33349,N_33491);
nor U33554 (N_33554,N_33006,N_33146);
nor U33555 (N_33555,N_33289,N_33155);
nor U33556 (N_33556,N_33470,N_33223);
and U33557 (N_33557,N_33197,N_33301);
nand U33558 (N_33558,N_33245,N_33341);
xor U33559 (N_33559,N_33186,N_33473);
nor U33560 (N_33560,N_33099,N_33050);
and U33561 (N_33561,N_33477,N_33043);
xnor U33562 (N_33562,N_33143,N_33071);
nand U33563 (N_33563,N_33452,N_33116);
nor U33564 (N_33564,N_33376,N_33388);
and U33565 (N_33565,N_33079,N_33469);
or U33566 (N_33566,N_33492,N_33027);
and U33567 (N_33567,N_33297,N_33372);
and U33568 (N_33568,N_33072,N_33467);
or U33569 (N_33569,N_33325,N_33320);
or U33570 (N_33570,N_33167,N_33094);
or U33571 (N_33571,N_33100,N_33067);
nand U33572 (N_33572,N_33293,N_33066);
nand U33573 (N_33573,N_33150,N_33003);
nand U33574 (N_33574,N_33311,N_33075);
xor U33575 (N_33575,N_33415,N_33125);
or U33576 (N_33576,N_33444,N_33010);
xor U33577 (N_33577,N_33277,N_33337);
and U33578 (N_33578,N_33145,N_33348);
nand U33579 (N_33579,N_33486,N_33373);
xnor U33580 (N_33580,N_33458,N_33087);
and U33581 (N_33581,N_33101,N_33474);
or U33582 (N_33582,N_33409,N_33366);
nor U33583 (N_33583,N_33152,N_33193);
nand U33584 (N_33584,N_33346,N_33487);
nand U33585 (N_33585,N_33445,N_33334);
or U33586 (N_33586,N_33181,N_33209);
nor U33587 (N_33587,N_33433,N_33069);
nor U33588 (N_33588,N_33138,N_33338);
xor U33589 (N_33589,N_33171,N_33303);
and U33590 (N_33590,N_33191,N_33423);
xor U33591 (N_33591,N_33479,N_33030);
or U33592 (N_33592,N_33287,N_33264);
and U33593 (N_33593,N_33355,N_33319);
nor U33594 (N_33594,N_33275,N_33312);
or U33595 (N_33595,N_33025,N_33326);
nand U33596 (N_33596,N_33219,N_33288);
or U33597 (N_33597,N_33118,N_33196);
and U33598 (N_33598,N_33361,N_33013);
and U33599 (N_33599,N_33053,N_33489);
and U33600 (N_33600,N_33426,N_33173);
nand U33601 (N_33601,N_33226,N_33280);
and U33602 (N_33602,N_33286,N_33317);
nand U33603 (N_33603,N_33306,N_33456);
and U33604 (N_33604,N_33472,N_33476);
nand U33605 (N_33605,N_33198,N_33192);
or U33606 (N_33606,N_33427,N_33252);
nor U33607 (N_33607,N_33424,N_33273);
xnor U33608 (N_33608,N_33149,N_33183);
nand U33609 (N_33609,N_33466,N_33124);
nor U33610 (N_33610,N_33214,N_33184);
and U33611 (N_33611,N_33266,N_33154);
and U33612 (N_33612,N_33032,N_33090);
xor U33613 (N_33613,N_33263,N_33195);
xnor U33614 (N_33614,N_33227,N_33028);
xor U33615 (N_33615,N_33104,N_33004);
nand U33616 (N_33616,N_33403,N_33254);
nand U33617 (N_33617,N_33047,N_33088);
nor U33618 (N_33618,N_33336,N_33405);
nor U33619 (N_33619,N_33036,N_33478);
nor U33620 (N_33620,N_33234,N_33439);
and U33621 (N_33621,N_33151,N_33213);
nor U33622 (N_33622,N_33108,N_33310);
nand U33623 (N_33623,N_33132,N_33260);
or U33624 (N_33624,N_33230,N_33014);
nand U33625 (N_33625,N_33238,N_33428);
nand U33626 (N_33626,N_33141,N_33250);
nand U33627 (N_33627,N_33045,N_33451);
xor U33628 (N_33628,N_33111,N_33165);
nor U33629 (N_33629,N_33352,N_33029);
and U33630 (N_33630,N_33057,N_33037);
nand U33631 (N_33631,N_33353,N_33429);
xnor U33632 (N_33632,N_33239,N_33256);
xor U33633 (N_33633,N_33343,N_33211);
nor U33634 (N_33634,N_33368,N_33169);
xor U33635 (N_33635,N_33331,N_33441);
or U33636 (N_33636,N_33204,N_33065);
nand U33637 (N_33637,N_33205,N_33318);
nand U33638 (N_33638,N_33242,N_33134);
or U33639 (N_33639,N_33435,N_33251);
and U33640 (N_33640,N_33342,N_33438);
nand U33641 (N_33641,N_33437,N_33265);
nor U33642 (N_33642,N_33258,N_33483);
nand U33643 (N_33643,N_33011,N_33330);
and U33644 (N_33644,N_33207,N_33333);
nand U33645 (N_33645,N_33026,N_33222);
nor U33646 (N_33646,N_33323,N_33005);
nor U33647 (N_33647,N_33117,N_33255);
nand U33648 (N_33648,N_33130,N_33127);
or U33649 (N_33649,N_33148,N_33278);
xnor U33650 (N_33650,N_33016,N_33302);
nand U33651 (N_33651,N_33276,N_33281);
or U33652 (N_33652,N_33001,N_33370);
or U33653 (N_33653,N_33202,N_33292);
xor U33654 (N_33654,N_33158,N_33034);
nor U33655 (N_33655,N_33431,N_33495);
or U33656 (N_33656,N_33354,N_33488);
and U33657 (N_33657,N_33164,N_33322);
nand U33658 (N_33658,N_33172,N_33144);
xnor U33659 (N_33659,N_33364,N_33061);
xor U33660 (N_33660,N_33023,N_33314);
nand U33661 (N_33661,N_33033,N_33073);
or U33662 (N_33662,N_33414,N_33236);
nor U33663 (N_33663,N_33233,N_33359);
nand U33664 (N_33664,N_33484,N_33105);
or U33665 (N_33665,N_33309,N_33411);
nor U33666 (N_33666,N_33170,N_33298);
and U33667 (N_33667,N_33385,N_33048);
and U33668 (N_33668,N_33360,N_33068);
nand U33669 (N_33669,N_33274,N_33247);
or U33670 (N_33670,N_33114,N_33078);
nand U33671 (N_33671,N_33147,N_33482);
and U33672 (N_33672,N_33267,N_33160);
nor U33673 (N_33673,N_33383,N_33241);
and U33674 (N_33674,N_33375,N_33422);
nor U33675 (N_33675,N_33215,N_33244);
nand U33676 (N_33676,N_33188,N_33232);
nor U33677 (N_33677,N_33249,N_33009);
and U33678 (N_33678,N_33485,N_33291);
xnor U33679 (N_33679,N_33382,N_33054);
or U33680 (N_33680,N_33046,N_33417);
or U33681 (N_33681,N_33404,N_33077);
or U33682 (N_33682,N_33240,N_33221);
and U33683 (N_33683,N_33253,N_33294);
nand U33684 (N_33684,N_33447,N_33182);
or U33685 (N_33685,N_33296,N_33374);
or U33686 (N_33686,N_33175,N_33200);
or U33687 (N_33687,N_33102,N_33279);
and U33688 (N_33688,N_33450,N_33377);
xor U33689 (N_33689,N_33440,N_33044);
xor U33690 (N_33690,N_33237,N_33380);
or U33691 (N_33691,N_33156,N_33389);
or U33692 (N_33692,N_33339,N_33008);
xnor U33693 (N_33693,N_33494,N_33397);
nand U33694 (N_33694,N_33299,N_33460);
and U33695 (N_33695,N_33040,N_33018);
and U33696 (N_33696,N_33217,N_33425);
nor U33697 (N_33697,N_33228,N_33345);
or U33698 (N_33698,N_33399,N_33110);
nand U33699 (N_33699,N_33344,N_33185);
or U33700 (N_33700,N_33248,N_33092);
nor U33701 (N_33701,N_33365,N_33229);
and U33702 (N_33702,N_33231,N_33002);
and U33703 (N_33703,N_33407,N_33307);
xor U33704 (N_33704,N_33199,N_33017);
and U33705 (N_33705,N_33189,N_33269);
and U33706 (N_33706,N_33371,N_33329);
and U33707 (N_33707,N_33097,N_33093);
or U33708 (N_33708,N_33007,N_33315);
nand U33709 (N_33709,N_33168,N_33163);
xor U33710 (N_33710,N_33308,N_33464);
or U33711 (N_33711,N_33392,N_33133);
xor U33712 (N_33712,N_33395,N_33052);
xor U33713 (N_33713,N_33420,N_33321);
nor U33714 (N_33714,N_33177,N_33225);
nor U33715 (N_33715,N_33243,N_33035);
nor U33716 (N_33716,N_33268,N_33384);
and U33717 (N_33717,N_33262,N_33406);
nand U33718 (N_33718,N_33019,N_33261);
or U33719 (N_33719,N_33490,N_33129);
or U33720 (N_33720,N_33080,N_33012);
nor U33721 (N_33721,N_33201,N_33497);
nand U33722 (N_33722,N_33416,N_33203);
or U33723 (N_33723,N_33000,N_33282);
nand U33724 (N_33724,N_33174,N_33176);
nand U33725 (N_33725,N_33106,N_33131);
or U33726 (N_33726,N_33455,N_33362);
nand U33727 (N_33727,N_33218,N_33300);
nor U33728 (N_33728,N_33391,N_33393);
and U33729 (N_33729,N_33430,N_33103);
nand U33730 (N_33730,N_33121,N_33070);
and U33731 (N_33731,N_33257,N_33448);
nand U33732 (N_33732,N_33055,N_33084);
nor U33733 (N_33733,N_33398,N_33434);
or U33734 (N_33734,N_33394,N_33098);
or U33735 (N_33735,N_33212,N_33316);
nand U33736 (N_33736,N_33432,N_33107);
nand U33737 (N_33737,N_33020,N_33304);
nand U33738 (N_33738,N_33220,N_33180);
and U33739 (N_33739,N_33187,N_33166);
nand U33740 (N_33740,N_33015,N_33122);
and U33741 (N_33741,N_33480,N_33031);
xnor U33742 (N_33742,N_33283,N_33386);
nand U33743 (N_33743,N_33463,N_33142);
and U33744 (N_33744,N_33481,N_33408);
nor U33745 (N_33745,N_33113,N_33475);
and U33746 (N_33746,N_33381,N_33021);
xor U33747 (N_33747,N_33436,N_33442);
xor U33748 (N_33748,N_33421,N_33137);
xor U33749 (N_33749,N_33270,N_33313);
nor U33750 (N_33750,N_33474,N_33216);
and U33751 (N_33751,N_33307,N_33476);
nor U33752 (N_33752,N_33318,N_33461);
and U33753 (N_33753,N_33108,N_33203);
nand U33754 (N_33754,N_33467,N_33017);
and U33755 (N_33755,N_33073,N_33486);
nor U33756 (N_33756,N_33209,N_33374);
nor U33757 (N_33757,N_33003,N_33462);
and U33758 (N_33758,N_33239,N_33037);
nor U33759 (N_33759,N_33326,N_33252);
and U33760 (N_33760,N_33318,N_33432);
nor U33761 (N_33761,N_33037,N_33299);
and U33762 (N_33762,N_33011,N_33157);
and U33763 (N_33763,N_33384,N_33370);
xor U33764 (N_33764,N_33220,N_33109);
and U33765 (N_33765,N_33017,N_33064);
and U33766 (N_33766,N_33293,N_33155);
nand U33767 (N_33767,N_33412,N_33206);
nor U33768 (N_33768,N_33003,N_33308);
xnor U33769 (N_33769,N_33077,N_33377);
xnor U33770 (N_33770,N_33201,N_33012);
nand U33771 (N_33771,N_33075,N_33443);
nand U33772 (N_33772,N_33053,N_33276);
nor U33773 (N_33773,N_33025,N_33021);
xor U33774 (N_33774,N_33349,N_33220);
nand U33775 (N_33775,N_33030,N_33381);
or U33776 (N_33776,N_33290,N_33178);
nand U33777 (N_33777,N_33033,N_33095);
and U33778 (N_33778,N_33156,N_33248);
or U33779 (N_33779,N_33394,N_33127);
or U33780 (N_33780,N_33172,N_33222);
or U33781 (N_33781,N_33002,N_33456);
xor U33782 (N_33782,N_33255,N_33290);
xor U33783 (N_33783,N_33092,N_33407);
nand U33784 (N_33784,N_33262,N_33169);
xor U33785 (N_33785,N_33238,N_33000);
nor U33786 (N_33786,N_33403,N_33245);
nor U33787 (N_33787,N_33401,N_33129);
nand U33788 (N_33788,N_33262,N_33037);
and U33789 (N_33789,N_33252,N_33232);
nor U33790 (N_33790,N_33048,N_33308);
nor U33791 (N_33791,N_33391,N_33369);
nor U33792 (N_33792,N_33207,N_33015);
or U33793 (N_33793,N_33265,N_33299);
or U33794 (N_33794,N_33103,N_33116);
or U33795 (N_33795,N_33237,N_33337);
nor U33796 (N_33796,N_33273,N_33421);
or U33797 (N_33797,N_33244,N_33176);
or U33798 (N_33798,N_33199,N_33366);
xor U33799 (N_33799,N_33496,N_33127);
nand U33800 (N_33800,N_33409,N_33027);
or U33801 (N_33801,N_33346,N_33197);
nand U33802 (N_33802,N_33363,N_33414);
and U33803 (N_33803,N_33319,N_33375);
and U33804 (N_33804,N_33308,N_33395);
or U33805 (N_33805,N_33326,N_33283);
nand U33806 (N_33806,N_33332,N_33384);
nor U33807 (N_33807,N_33143,N_33369);
xor U33808 (N_33808,N_33052,N_33391);
nand U33809 (N_33809,N_33087,N_33072);
xor U33810 (N_33810,N_33278,N_33112);
nand U33811 (N_33811,N_33319,N_33228);
or U33812 (N_33812,N_33207,N_33451);
and U33813 (N_33813,N_33429,N_33391);
xnor U33814 (N_33814,N_33082,N_33244);
nor U33815 (N_33815,N_33492,N_33229);
nand U33816 (N_33816,N_33480,N_33173);
nand U33817 (N_33817,N_33149,N_33302);
nor U33818 (N_33818,N_33282,N_33431);
nor U33819 (N_33819,N_33132,N_33316);
nor U33820 (N_33820,N_33164,N_33168);
or U33821 (N_33821,N_33158,N_33232);
or U33822 (N_33822,N_33287,N_33444);
xor U33823 (N_33823,N_33443,N_33286);
or U33824 (N_33824,N_33440,N_33331);
and U33825 (N_33825,N_33172,N_33110);
xor U33826 (N_33826,N_33405,N_33006);
nor U33827 (N_33827,N_33140,N_33043);
nand U33828 (N_33828,N_33261,N_33478);
nor U33829 (N_33829,N_33203,N_33217);
and U33830 (N_33830,N_33354,N_33201);
xnor U33831 (N_33831,N_33076,N_33214);
nand U33832 (N_33832,N_33307,N_33050);
nand U33833 (N_33833,N_33400,N_33225);
nand U33834 (N_33834,N_33438,N_33429);
xor U33835 (N_33835,N_33393,N_33379);
nor U33836 (N_33836,N_33116,N_33378);
xnor U33837 (N_33837,N_33187,N_33155);
nor U33838 (N_33838,N_33073,N_33498);
xnor U33839 (N_33839,N_33161,N_33284);
or U33840 (N_33840,N_33230,N_33352);
or U33841 (N_33841,N_33392,N_33085);
or U33842 (N_33842,N_33464,N_33274);
nand U33843 (N_33843,N_33187,N_33338);
xor U33844 (N_33844,N_33480,N_33442);
nand U33845 (N_33845,N_33167,N_33269);
nor U33846 (N_33846,N_33094,N_33260);
nand U33847 (N_33847,N_33052,N_33462);
xor U33848 (N_33848,N_33275,N_33236);
or U33849 (N_33849,N_33048,N_33000);
and U33850 (N_33850,N_33478,N_33277);
nor U33851 (N_33851,N_33436,N_33144);
or U33852 (N_33852,N_33108,N_33279);
nand U33853 (N_33853,N_33418,N_33070);
nor U33854 (N_33854,N_33156,N_33088);
or U33855 (N_33855,N_33429,N_33018);
xnor U33856 (N_33856,N_33029,N_33056);
xnor U33857 (N_33857,N_33264,N_33012);
nand U33858 (N_33858,N_33154,N_33214);
or U33859 (N_33859,N_33132,N_33096);
and U33860 (N_33860,N_33314,N_33214);
or U33861 (N_33861,N_33497,N_33046);
nor U33862 (N_33862,N_33319,N_33219);
and U33863 (N_33863,N_33258,N_33409);
nor U33864 (N_33864,N_33045,N_33014);
xnor U33865 (N_33865,N_33082,N_33067);
xor U33866 (N_33866,N_33216,N_33467);
nor U33867 (N_33867,N_33161,N_33118);
xnor U33868 (N_33868,N_33202,N_33275);
or U33869 (N_33869,N_33061,N_33116);
nor U33870 (N_33870,N_33355,N_33359);
nand U33871 (N_33871,N_33076,N_33411);
or U33872 (N_33872,N_33178,N_33315);
xnor U33873 (N_33873,N_33311,N_33478);
nor U33874 (N_33874,N_33475,N_33080);
and U33875 (N_33875,N_33270,N_33421);
nor U33876 (N_33876,N_33429,N_33270);
or U33877 (N_33877,N_33343,N_33405);
or U33878 (N_33878,N_33490,N_33280);
nand U33879 (N_33879,N_33444,N_33265);
nand U33880 (N_33880,N_33164,N_33196);
nand U33881 (N_33881,N_33491,N_33322);
and U33882 (N_33882,N_33276,N_33127);
xor U33883 (N_33883,N_33275,N_33470);
xor U33884 (N_33884,N_33368,N_33303);
or U33885 (N_33885,N_33426,N_33210);
nor U33886 (N_33886,N_33067,N_33318);
and U33887 (N_33887,N_33200,N_33181);
or U33888 (N_33888,N_33139,N_33096);
nand U33889 (N_33889,N_33187,N_33079);
xnor U33890 (N_33890,N_33171,N_33046);
nand U33891 (N_33891,N_33345,N_33053);
and U33892 (N_33892,N_33305,N_33449);
or U33893 (N_33893,N_33011,N_33382);
nand U33894 (N_33894,N_33396,N_33420);
and U33895 (N_33895,N_33116,N_33044);
nor U33896 (N_33896,N_33375,N_33386);
nor U33897 (N_33897,N_33140,N_33236);
and U33898 (N_33898,N_33376,N_33158);
or U33899 (N_33899,N_33487,N_33012);
and U33900 (N_33900,N_33094,N_33446);
and U33901 (N_33901,N_33218,N_33009);
nand U33902 (N_33902,N_33488,N_33349);
xnor U33903 (N_33903,N_33275,N_33139);
nand U33904 (N_33904,N_33202,N_33102);
and U33905 (N_33905,N_33267,N_33481);
nor U33906 (N_33906,N_33154,N_33494);
and U33907 (N_33907,N_33396,N_33303);
and U33908 (N_33908,N_33280,N_33440);
and U33909 (N_33909,N_33197,N_33147);
nor U33910 (N_33910,N_33301,N_33408);
xor U33911 (N_33911,N_33201,N_33217);
or U33912 (N_33912,N_33037,N_33192);
and U33913 (N_33913,N_33162,N_33380);
nand U33914 (N_33914,N_33006,N_33353);
nand U33915 (N_33915,N_33072,N_33369);
nor U33916 (N_33916,N_33028,N_33128);
nor U33917 (N_33917,N_33151,N_33100);
nor U33918 (N_33918,N_33274,N_33483);
or U33919 (N_33919,N_33028,N_33311);
xor U33920 (N_33920,N_33028,N_33022);
xnor U33921 (N_33921,N_33199,N_33051);
nor U33922 (N_33922,N_33138,N_33381);
and U33923 (N_33923,N_33220,N_33183);
xnor U33924 (N_33924,N_33218,N_33383);
or U33925 (N_33925,N_33254,N_33308);
and U33926 (N_33926,N_33256,N_33328);
and U33927 (N_33927,N_33395,N_33242);
and U33928 (N_33928,N_33427,N_33153);
and U33929 (N_33929,N_33329,N_33231);
nand U33930 (N_33930,N_33373,N_33210);
xnor U33931 (N_33931,N_33345,N_33047);
xnor U33932 (N_33932,N_33146,N_33083);
xor U33933 (N_33933,N_33163,N_33151);
nor U33934 (N_33934,N_33116,N_33167);
and U33935 (N_33935,N_33427,N_33365);
nand U33936 (N_33936,N_33043,N_33413);
or U33937 (N_33937,N_33299,N_33221);
and U33938 (N_33938,N_33019,N_33314);
and U33939 (N_33939,N_33383,N_33068);
xnor U33940 (N_33940,N_33127,N_33476);
and U33941 (N_33941,N_33198,N_33446);
and U33942 (N_33942,N_33236,N_33420);
nand U33943 (N_33943,N_33474,N_33196);
xor U33944 (N_33944,N_33256,N_33123);
and U33945 (N_33945,N_33042,N_33227);
and U33946 (N_33946,N_33435,N_33293);
and U33947 (N_33947,N_33380,N_33462);
xnor U33948 (N_33948,N_33347,N_33386);
or U33949 (N_33949,N_33296,N_33278);
or U33950 (N_33950,N_33223,N_33415);
and U33951 (N_33951,N_33219,N_33158);
xnor U33952 (N_33952,N_33035,N_33054);
or U33953 (N_33953,N_33279,N_33442);
and U33954 (N_33954,N_33289,N_33436);
xor U33955 (N_33955,N_33455,N_33051);
and U33956 (N_33956,N_33323,N_33387);
nor U33957 (N_33957,N_33095,N_33006);
or U33958 (N_33958,N_33492,N_33020);
nand U33959 (N_33959,N_33241,N_33393);
xor U33960 (N_33960,N_33445,N_33372);
or U33961 (N_33961,N_33021,N_33240);
or U33962 (N_33962,N_33050,N_33047);
nand U33963 (N_33963,N_33184,N_33451);
xnor U33964 (N_33964,N_33331,N_33098);
xor U33965 (N_33965,N_33416,N_33111);
and U33966 (N_33966,N_33498,N_33135);
or U33967 (N_33967,N_33073,N_33006);
or U33968 (N_33968,N_33211,N_33172);
and U33969 (N_33969,N_33089,N_33127);
and U33970 (N_33970,N_33497,N_33356);
xnor U33971 (N_33971,N_33061,N_33343);
or U33972 (N_33972,N_33341,N_33129);
nor U33973 (N_33973,N_33348,N_33401);
and U33974 (N_33974,N_33242,N_33154);
xnor U33975 (N_33975,N_33122,N_33493);
xor U33976 (N_33976,N_33106,N_33387);
nor U33977 (N_33977,N_33174,N_33427);
or U33978 (N_33978,N_33331,N_33494);
and U33979 (N_33979,N_33116,N_33366);
xor U33980 (N_33980,N_33459,N_33140);
and U33981 (N_33981,N_33115,N_33459);
xnor U33982 (N_33982,N_33261,N_33355);
nand U33983 (N_33983,N_33453,N_33318);
or U33984 (N_33984,N_33263,N_33186);
nand U33985 (N_33985,N_33472,N_33320);
nand U33986 (N_33986,N_33222,N_33204);
nand U33987 (N_33987,N_33357,N_33071);
or U33988 (N_33988,N_33225,N_33328);
or U33989 (N_33989,N_33163,N_33110);
nand U33990 (N_33990,N_33462,N_33441);
and U33991 (N_33991,N_33215,N_33383);
and U33992 (N_33992,N_33462,N_33002);
nor U33993 (N_33993,N_33355,N_33200);
nor U33994 (N_33994,N_33265,N_33056);
or U33995 (N_33995,N_33088,N_33146);
xor U33996 (N_33996,N_33305,N_33073);
nand U33997 (N_33997,N_33375,N_33434);
xnor U33998 (N_33998,N_33106,N_33322);
and U33999 (N_33999,N_33221,N_33056);
and U34000 (N_34000,N_33628,N_33856);
nor U34001 (N_34001,N_33645,N_33984);
xnor U34002 (N_34002,N_33740,N_33608);
nor U34003 (N_34003,N_33950,N_33842);
and U34004 (N_34004,N_33992,N_33962);
xor U34005 (N_34005,N_33864,N_33785);
nand U34006 (N_34006,N_33771,N_33937);
nand U34007 (N_34007,N_33516,N_33668);
xnor U34008 (N_34008,N_33996,N_33784);
nor U34009 (N_34009,N_33923,N_33692);
nor U34010 (N_34010,N_33582,N_33916);
nor U34011 (N_34011,N_33929,N_33625);
or U34012 (N_34012,N_33698,N_33725);
or U34013 (N_34013,N_33732,N_33726);
xnor U34014 (N_34014,N_33972,N_33642);
nand U34015 (N_34015,N_33769,N_33670);
nor U34016 (N_34016,N_33956,N_33612);
or U34017 (N_34017,N_33700,N_33559);
and U34018 (N_34018,N_33677,N_33696);
nor U34019 (N_34019,N_33540,N_33720);
and U34020 (N_34020,N_33606,N_33714);
nand U34021 (N_34021,N_33886,N_33795);
or U34022 (N_34022,N_33835,N_33525);
or U34023 (N_34023,N_33613,N_33605);
xor U34024 (N_34024,N_33805,N_33709);
xnor U34025 (N_34025,N_33837,N_33686);
xnor U34026 (N_34026,N_33596,N_33581);
and U34027 (N_34027,N_33979,N_33858);
xor U34028 (N_34028,N_33727,N_33601);
nor U34029 (N_34029,N_33533,N_33825);
or U34030 (N_34030,N_33846,N_33555);
xnor U34031 (N_34031,N_33913,N_33764);
and U34032 (N_34032,N_33500,N_33621);
nand U34033 (N_34033,N_33942,N_33620);
and U34034 (N_34034,N_33813,N_33724);
or U34035 (N_34035,N_33821,N_33501);
or U34036 (N_34036,N_33954,N_33607);
nand U34037 (N_34037,N_33797,N_33713);
and U34038 (N_34038,N_33861,N_33780);
or U34039 (N_34039,N_33800,N_33891);
nor U34040 (N_34040,N_33566,N_33745);
nand U34041 (N_34041,N_33624,N_33952);
nor U34042 (N_34042,N_33752,N_33778);
or U34043 (N_34043,N_33883,N_33591);
nand U34044 (N_34044,N_33505,N_33770);
nand U34045 (N_34045,N_33884,N_33747);
and U34046 (N_34046,N_33548,N_33875);
or U34047 (N_34047,N_33661,N_33594);
and U34048 (N_34048,N_33760,N_33834);
or U34049 (N_34049,N_33958,N_33993);
nor U34050 (N_34050,N_33863,N_33564);
xnor U34051 (N_34051,N_33640,N_33666);
nor U34052 (N_34052,N_33663,N_33574);
nor U34053 (N_34053,N_33838,N_33552);
and U34054 (N_34054,N_33761,N_33911);
nor U34055 (N_34055,N_33506,N_33918);
nand U34056 (N_34056,N_33791,N_33964);
or U34057 (N_34057,N_33966,N_33694);
nor U34058 (N_34058,N_33828,N_33810);
or U34059 (N_34059,N_33908,N_33741);
and U34060 (N_34060,N_33792,N_33815);
and U34061 (N_34061,N_33998,N_33939);
and U34062 (N_34062,N_33748,N_33907);
or U34063 (N_34063,N_33866,N_33789);
xnor U34064 (N_34064,N_33894,N_33901);
nor U34065 (N_34065,N_33699,N_33547);
nand U34066 (N_34066,N_33757,N_33961);
nor U34067 (N_34067,N_33573,N_33804);
and U34068 (N_34068,N_33563,N_33836);
xnor U34069 (N_34069,N_33655,N_33653);
nor U34070 (N_34070,N_33708,N_33600);
and U34071 (N_34071,N_33779,N_33603);
nor U34072 (N_34072,N_33595,N_33922);
xnor U34073 (N_34073,N_33584,N_33976);
xnor U34074 (N_34074,N_33627,N_33843);
xnor U34075 (N_34075,N_33841,N_33744);
or U34076 (N_34076,N_33638,N_33963);
nand U34077 (N_34077,N_33514,N_33746);
nand U34078 (N_34078,N_33722,N_33840);
xor U34079 (N_34079,N_33987,N_33953);
and U34080 (N_34080,N_33615,N_33545);
xor U34081 (N_34081,N_33572,N_33560);
or U34082 (N_34082,N_33577,N_33951);
or U34083 (N_34083,N_33991,N_33524);
or U34084 (N_34084,N_33737,N_33799);
or U34085 (N_34085,N_33848,N_33537);
and U34086 (N_34086,N_33710,N_33728);
nand U34087 (N_34087,N_33860,N_33845);
nand U34088 (N_34088,N_33788,N_33915);
or U34089 (N_34089,N_33862,N_33729);
nor U34090 (N_34090,N_33753,N_33721);
and U34091 (N_34091,N_33510,N_33672);
and U34092 (N_34092,N_33902,N_33676);
nand U34093 (N_34093,N_33733,N_33990);
xor U34094 (N_34094,N_33597,N_33775);
nor U34095 (N_34095,N_33543,N_33647);
xor U34096 (N_34096,N_33716,N_33635);
nand U34097 (N_34097,N_33509,N_33656);
nand U34098 (N_34098,N_33568,N_33890);
xor U34099 (N_34099,N_33882,N_33830);
nor U34100 (N_34100,N_33602,N_33521);
xor U34101 (N_34101,N_33691,N_33852);
nor U34102 (N_34102,N_33895,N_33933);
xnor U34103 (N_34103,N_33684,N_33742);
xor U34104 (N_34104,N_33783,N_33580);
nor U34105 (N_34105,N_33946,N_33558);
xnor U34106 (N_34106,N_33518,N_33865);
xor U34107 (N_34107,N_33925,N_33641);
nor U34108 (N_34108,N_33616,N_33879);
nand U34109 (N_34109,N_33871,N_33812);
and U34110 (N_34110,N_33829,N_33735);
xor U34111 (N_34111,N_33850,N_33701);
or U34112 (N_34112,N_33697,N_33773);
xor U34113 (N_34113,N_33648,N_33934);
and U34114 (N_34114,N_33685,N_33639);
or U34115 (N_34115,N_33989,N_33578);
nand U34116 (N_34116,N_33553,N_33738);
nand U34117 (N_34117,N_33534,N_33502);
nand U34118 (N_34118,N_33557,N_33816);
xor U34119 (N_34119,N_33867,N_33680);
nor U34120 (N_34120,N_33675,N_33973);
xor U34121 (N_34121,N_33554,N_33960);
or U34122 (N_34122,N_33579,N_33588);
and U34123 (N_34123,N_33814,N_33693);
nor U34124 (N_34124,N_33702,N_33712);
or U34125 (N_34125,N_33983,N_33539);
and U34126 (N_34126,N_33535,N_33567);
or U34127 (N_34127,N_33823,N_33622);
nor U34128 (N_34128,N_33549,N_33619);
or U34129 (N_34129,N_33767,N_33528);
nor U34130 (N_34130,N_33889,N_33774);
and U34131 (N_34131,N_33936,N_33633);
and U34132 (N_34132,N_33681,N_33519);
or U34133 (N_34133,N_33985,N_33855);
xnor U34134 (N_34134,N_33530,N_33590);
nor U34135 (N_34135,N_33811,N_33669);
nand U34136 (N_34136,N_33561,N_33806);
or U34137 (N_34137,N_33965,N_33718);
nor U34138 (N_34138,N_33526,N_33919);
and U34139 (N_34139,N_33957,N_33935);
or U34140 (N_34140,N_33776,N_33585);
nand U34141 (N_34141,N_33978,N_33515);
xnor U34142 (N_34142,N_33593,N_33654);
and U34143 (N_34143,N_33796,N_33874);
nor U34144 (N_34144,N_33927,N_33562);
nor U34145 (N_34145,N_33538,N_33660);
or U34146 (N_34146,N_33872,N_33614);
and U34147 (N_34147,N_33751,N_33731);
nor U34148 (N_34148,N_33833,N_33587);
nor U34149 (N_34149,N_33772,N_33794);
and U34150 (N_34150,N_33906,N_33920);
and U34151 (N_34151,N_33904,N_33926);
nor U34152 (N_34152,N_33623,N_33903);
nor U34153 (N_34153,N_33977,N_33598);
nand U34154 (N_34154,N_33687,N_33610);
nor U34155 (N_34155,N_33592,N_33730);
nor U34156 (N_34156,N_33707,N_33532);
or U34157 (N_34157,N_33604,N_33636);
nand U34158 (N_34158,N_33690,N_33632);
xnor U34159 (N_34159,N_33754,N_33831);
and U34160 (N_34160,N_33766,N_33899);
nor U34161 (N_34161,N_33881,N_33523);
nand U34162 (N_34162,N_33763,N_33544);
nand U34163 (N_34163,N_33999,N_33893);
nor U34164 (N_34164,N_33947,N_33576);
xnor U34165 (N_34165,N_33705,N_33885);
nor U34166 (N_34166,N_33695,N_33798);
nor U34167 (N_34167,N_33912,N_33851);
and U34168 (N_34168,N_33659,N_33717);
and U34169 (N_34169,N_33898,N_33917);
or U34170 (N_34170,N_33542,N_33704);
xnor U34171 (N_34171,N_33749,N_33529);
xor U34172 (N_34172,N_33887,N_33611);
or U34173 (N_34173,N_33793,N_33631);
and U34174 (N_34174,N_33928,N_33507);
xnor U34175 (N_34175,N_33880,N_33630);
and U34176 (N_34176,N_33508,N_33643);
nor U34177 (N_34177,N_33981,N_33674);
xor U34178 (N_34178,N_33940,N_33988);
nor U34179 (N_34179,N_33967,N_33678);
xor U34180 (N_34180,N_33679,N_33536);
or U34181 (N_34181,N_33671,N_33877);
nand U34182 (N_34182,N_33503,N_33897);
nand U34183 (N_34183,N_33667,N_33808);
xnor U34184 (N_34184,N_33626,N_33803);
xor U34185 (N_34185,N_33859,N_33575);
and U34186 (N_34186,N_33873,N_33959);
nand U34187 (N_34187,N_33924,N_33909);
and U34188 (N_34188,N_33504,N_33736);
nand U34189 (N_34189,N_33826,N_33646);
xor U34190 (N_34190,N_33765,N_33723);
nand U34191 (N_34191,N_33551,N_33931);
nand U34192 (N_34192,N_33629,N_33556);
nor U34193 (N_34193,N_33719,N_33520);
nand U34194 (N_34194,N_33968,N_33827);
xor U34195 (N_34195,N_33777,N_33809);
nor U34196 (N_34196,N_33900,N_33832);
nand U34197 (N_34197,N_33941,N_33652);
nor U34198 (N_34198,N_33688,N_33944);
nor U34199 (N_34199,N_33618,N_33649);
or U34200 (N_34200,N_33786,N_33673);
nor U34201 (N_34201,N_33546,N_33970);
or U34202 (N_34202,N_33715,N_33974);
and U34203 (N_34203,N_33743,N_33711);
nand U34204 (N_34204,N_33969,N_33982);
nand U34205 (N_34205,N_33787,N_33689);
nand U34206 (N_34206,N_33762,N_33822);
xnor U34207 (N_34207,N_33945,N_33802);
xnor U34208 (N_34208,N_33818,N_33876);
xor U34209 (N_34209,N_33790,N_33527);
and U34210 (N_34210,N_33869,N_33651);
xnor U34211 (N_34211,N_33955,N_33758);
xnor U34212 (N_34212,N_33910,N_33650);
xor U34213 (N_34213,N_33662,N_33657);
or U34214 (N_34214,N_33511,N_33658);
and U34215 (N_34215,N_33948,N_33522);
nand U34216 (N_34216,N_33586,N_33932);
xnor U34217 (N_34217,N_33994,N_33839);
nand U34218 (N_34218,N_33569,N_33571);
nor U34219 (N_34219,N_33820,N_33750);
nand U34220 (N_34220,N_33664,N_33782);
nand U34221 (N_34221,N_33665,N_33550);
and U34222 (N_34222,N_33755,N_33819);
or U34223 (N_34223,N_33531,N_33986);
nor U34224 (N_34224,N_33995,N_33921);
nand U34225 (N_34225,N_33541,N_33801);
or U34226 (N_34226,N_33589,N_33878);
nor U34227 (N_34227,N_33892,N_33896);
nor U34228 (N_34228,N_33570,N_33739);
nor U34229 (N_34229,N_33599,N_33609);
nand U34230 (N_34230,N_33517,N_33870);
nand U34231 (N_34231,N_33637,N_33644);
nor U34232 (N_34232,N_33854,N_33949);
and U34233 (N_34233,N_33943,N_33807);
nor U34234 (N_34234,N_33905,N_33914);
xor U34235 (N_34235,N_33682,N_33853);
or U34236 (N_34236,N_33781,N_33706);
and U34237 (N_34237,N_33512,N_33759);
or U34238 (N_34238,N_33938,N_33824);
nand U34239 (N_34239,N_33888,N_33847);
and U34240 (N_34240,N_33734,N_33844);
or U34241 (N_34241,N_33971,N_33849);
nor U34242 (N_34242,N_33997,N_33683);
or U34243 (N_34243,N_33513,N_33703);
and U34244 (N_34244,N_33768,N_33817);
xnor U34245 (N_34245,N_33930,N_33868);
nor U34246 (N_34246,N_33857,N_33565);
xor U34247 (N_34247,N_33634,N_33617);
or U34248 (N_34248,N_33975,N_33756);
and U34249 (N_34249,N_33583,N_33980);
nor U34250 (N_34250,N_33581,N_33989);
and U34251 (N_34251,N_33548,N_33768);
and U34252 (N_34252,N_33652,N_33638);
and U34253 (N_34253,N_33755,N_33510);
or U34254 (N_34254,N_33953,N_33819);
and U34255 (N_34255,N_33799,N_33683);
or U34256 (N_34256,N_33811,N_33676);
nand U34257 (N_34257,N_33717,N_33719);
nor U34258 (N_34258,N_33620,N_33560);
nor U34259 (N_34259,N_33602,N_33748);
nand U34260 (N_34260,N_33667,N_33902);
xnor U34261 (N_34261,N_33630,N_33824);
nor U34262 (N_34262,N_33650,N_33866);
nand U34263 (N_34263,N_33700,N_33514);
xnor U34264 (N_34264,N_33646,N_33592);
or U34265 (N_34265,N_33852,N_33935);
or U34266 (N_34266,N_33717,N_33684);
nand U34267 (N_34267,N_33728,N_33868);
nand U34268 (N_34268,N_33760,N_33919);
nor U34269 (N_34269,N_33988,N_33802);
or U34270 (N_34270,N_33924,N_33930);
xnor U34271 (N_34271,N_33827,N_33625);
nor U34272 (N_34272,N_33796,N_33593);
and U34273 (N_34273,N_33534,N_33607);
or U34274 (N_34274,N_33605,N_33790);
and U34275 (N_34275,N_33782,N_33565);
xnor U34276 (N_34276,N_33767,N_33703);
nor U34277 (N_34277,N_33715,N_33885);
xor U34278 (N_34278,N_33659,N_33817);
and U34279 (N_34279,N_33637,N_33709);
xnor U34280 (N_34280,N_33559,N_33952);
nand U34281 (N_34281,N_33913,N_33599);
and U34282 (N_34282,N_33931,N_33944);
and U34283 (N_34283,N_33508,N_33868);
or U34284 (N_34284,N_33768,N_33861);
or U34285 (N_34285,N_33651,N_33624);
nor U34286 (N_34286,N_33964,N_33761);
xnor U34287 (N_34287,N_33897,N_33748);
and U34288 (N_34288,N_33974,N_33609);
or U34289 (N_34289,N_33510,N_33581);
nor U34290 (N_34290,N_33689,N_33771);
and U34291 (N_34291,N_33803,N_33856);
nor U34292 (N_34292,N_33788,N_33859);
or U34293 (N_34293,N_33868,N_33621);
nor U34294 (N_34294,N_33612,N_33579);
nand U34295 (N_34295,N_33723,N_33843);
or U34296 (N_34296,N_33903,N_33608);
nand U34297 (N_34297,N_33820,N_33793);
xor U34298 (N_34298,N_33720,N_33917);
nand U34299 (N_34299,N_33844,N_33572);
nor U34300 (N_34300,N_33572,N_33912);
or U34301 (N_34301,N_33973,N_33827);
or U34302 (N_34302,N_33530,N_33695);
nor U34303 (N_34303,N_33727,N_33572);
and U34304 (N_34304,N_33713,N_33948);
nand U34305 (N_34305,N_33997,N_33988);
nand U34306 (N_34306,N_33561,N_33612);
and U34307 (N_34307,N_33651,N_33633);
nand U34308 (N_34308,N_33661,N_33835);
xnor U34309 (N_34309,N_33631,N_33807);
and U34310 (N_34310,N_33970,N_33652);
nor U34311 (N_34311,N_33555,N_33692);
and U34312 (N_34312,N_33564,N_33797);
or U34313 (N_34313,N_33861,N_33555);
or U34314 (N_34314,N_33566,N_33710);
nand U34315 (N_34315,N_33764,N_33650);
xnor U34316 (N_34316,N_33711,N_33748);
and U34317 (N_34317,N_33602,N_33610);
and U34318 (N_34318,N_33780,N_33937);
or U34319 (N_34319,N_33839,N_33503);
nor U34320 (N_34320,N_33731,N_33526);
or U34321 (N_34321,N_33750,N_33890);
or U34322 (N_34322,N_33755,N_33716);
or U34323 (N_34323,N_33632,N_33589);
or U34324 (N_34324,N_33823,N_33828);
nor U34325 (N_34325,N_33681,N_33529);
or U34326 (N_34326,N_33658,N_33600);
or U34327 (N_34327,N_33585,N_33642);
nor U34328 (N_34328,N_33724,N_33619);
nand U34329 (N_34329,N_33567,N_33834);
xnor U34330 (N_34330,N_33856,N_33604);
or U34331 (N_34331,N_33683,N_33814);
xor U34332 (N_34332,N_33881,N_33536);
xnor U34333 (N_34333,N_33683,N_33842);
or U34334 (N_34334,N_33720,N_33578);
xnor U34335 (N_34335,N_33945,N_33504);
nor U34336 (N_34336,N_33528,N_33514);
and U34337 (N_34337,N_33544,N_33898);
or U34338 (N_34338,N_33678,N_33778);
and U34339 (N_34339,N_33570,N_33861);
nor U34340 (N_34340,N_33967,N_33677);
and U34341 (N_34341,N_33612,N_33804);
xnor U34342 (N_34342,N_33960,N_33569);
or U34343 (N_34343,N_33872,N_33956);
and U34344 (N_34344,N_33755,N_33674);
or U34345 (N_34345,N_33674,N_33970);
nor U34346 (N_34346,N_33649,N_33693);
nand U34347 (N_34347,N_33766,N_33684);
xor U34348 (N_34348,N_33724,N_33679);
or U34349 (N_34349,N_33800,N_33602);
xnor U34350 (N_34350,N_33520,N_33576);
and U34351 (N_34351,N_33988,N_33916);
nand U34352 (N_34352,N_33595,N_33654);
nand U34353 (N_34353,N_33981,N_33555);
nand U34354 (N_34354,N_33548,N_33570);
nor U34355 (N_34355,N_33706,N_33812);
and U34356 (N_34356,N_33682,N_33916);
xor U34357 (N_34357,N_33566,N_33777);
xor U34358 (N_34358,N_33819,N_33530);
nor U34359 (N_34359,N_33985,N_33596);
or U34360 (N_34360,N_33847,N_33933);
nor U34361 (N_34361,N_33934,N_33979);
xnor U34362 (N_34362,N_33574,N_33680);
or U34363 (N_34363,N_33657,N_33806);
nor U34364 (N_34364,N_33919,N_33505);
nor U34365 (N_34365,N_33563,N_33603);
xnor U34366 (N_34366,N_33547,N_33741);
nor U34367 (N_34367,N_33513,N_33862);
nand U34368 (N_34368,N_33786,N_33505);
or U34369 (N_34369,N_33879,N_33932);
or U34370 (N_34370,N_33820,N_33867);
nor U34371 (N_34371,N_33581,N_33559);
and U34372 (N_34372,N_33976,N_33847);
xnor U34373 (N_34373,N_33867,N_33511);
nand U34374 (N_34374,N_33505,N_33838);
and U34375 (N_34375,N_33693,N_33636);
or U34376 (N_34376,N_33639,N_33514);
nor U34377 (N_34377,N_33908,N_33930);
nand U34378 (N_34378,N_33858,N_33944);
nor U34379 (N_34379,N_33684,N_33757);
nand U34380 (N_34380,N_33509,N_33590);
xnor U34381 (N_34381,N_33787,N_33727);
or U34382 (N_34382,N_33962,N_33931);
xor U34383 (N_34383,N_33891,N_33583);
nand U34384 (N_34384,N_33952,N_33837);
xor U34385 (N_34385,N_33575,N_33798);
nand U34386 (N_34386,N_33943,N_33671);
xnor U34387 (N_34387,N_33922,N_33525);
nand U34388 (N_34388,N_33976,N_33923);
nor U34389 (N_34389,N_33971,N_33570);
nor U34390 (N_34390,N_33513,N_33765);
and U34391 (N_34391,N_33670,N_33902);
and U34392 (N_34392,N_33591,N_33714);
nor U34393 (N_34393,N_33977,N_33874);
nand U34394 (N_34394,N_33721,N_33907);
nand U34395 (N_34395,N_33880,N_33613);
and U34396 (N_34396,N_33633,N_33582);
or U34397 (N_34397,N_33815,N_33822);
and U34398 (N_34398,N_33583,N_33503);
nor U34399 (N_34399,N_33605,N_33831);
xnor U34400 (N_34400,N_33932,N_33527);
nand U34401 (N_34401,N_33946,N_33537);
xnor U34402 (N_34402,N_33653,N_33782);
or U34403 (N_34403,N_33637,N_33511);
nand U34404 (N_34404,N_33557,N_33692);
and U34405 (N_34405,N_33999,N_33866);
nor U34406 (N_34406,N_33874,N_33802);
nand U34407 (N_34407,N_33641,N_33621);
nor U34408 (N_34408,N_33906,N_33808);
nand U34409 (N_34409,N_33682,N_33578);
or U34410 (N_34410,N_33623,N_33680);
and U34411 (N_34411,N_33562,N_33553);
nand U34412 (N_34412,N_33781,N_33646);
nor U34413 (N_34413,N_33565,N_33750);
xnor U34414 (N_34414,N_33736,N_33870);
xnor U34415 (N_34415,N_33754,N_33716);
xor U34416 (N_34416,N_33906,N_33597);
nand U34417 (N_34417,N_33776,N_33964);
nor U34418 (N_34418,N_33528,N_33545);
nand U34419 (N_34419,N_33626,N_33652);
xnor U34420 (N_34420,N_33678,N_33585);
and U34421 (N_34421,N_33688,N_33617);
nor U34422 (N_34422,N_33882,N_33609);
nand U34423 (N_34423,N_33785,N_33715);
nand U34424 (N_34424,N_33808,N_33629);
xor U34425 (N_34425,N_33582,N_33825);
nor U34426 (N_34426,N_33656,N_33811);
and U34427 (N_34427,N_33544,N_33821);
or U34428 (N_34428,N_33804,N_33604);
or U34429 (N_34429,N_33777,N_33629);
nor U34430 (N_34430,N_33881,N_33731);
xnor U34431 (N_34431,N_33857,N_33883);
or U34432 (N_34432,N_33964,N_33883);
or U34433 (N_34433,N_33732,N_33556);
xnor U34434 (N_34434,N_33523,N_33936);
and U34435 (N_34435,N_33637,N_33940);
and U34436 (N_34436,N_33785,N_33574);
or U34437 (N_34437,N_33911,N_33942);
xnor U34438 (N_34438,N_33704,N_33827);
nand U34439 (N_34439,N_33525,N_33771);
and U34440 (N_34440,N_33722,N_33916);
or U34441 (N_34441,N_33833,N_33710);
nand U34442 (N_34442,N_33851,N_33584);
or U34443 (N_34443,N_33780,N_33809);
and U34444 (N_34444,N_33977,N_33962);
xnor U34445 (N_34445,N_33540,N_33559);
or U34446 (N_34446,N_33574,N_33506);
and U34447 (N_34447,N_33931,N_33954);
or U34448 (N_34448,N_33743,N_33869);
and U34449 (N_34449,N_33701,N_33622);
nand U34450 (N_34450,N_33570,N_33559);
nand U34451 (N_34451,N_33861,N_33558);
nor U34452 (N_34452,N_33821,N_33901);
or U34453 (N_34453,N_33725,N_33821);
and U34454 (N_34454,N_33728,N_33685);
or U34455 (N_34455,N_33622,N_33948);
and U34456 (N_34456,N_33931,N_33601);
and U34457 (N_34457,N_33712,N_33856);
or U34458 (N_34458,N_33638,N_33782);
nand U34459 (N_34459,N_33762,N_33767);
xnor U34460 (N_34460,N_33873,N_33958);
nand U34461 (N_34461,N_33808,N_33647);
xnor U34462 (N_34462,N_33800,N_33610);
or U34463 (N_34463,N_33784,N_33531);
nor U34464 (N_34464,N_33571,N_33555);
or U34465 (N_34465,N_33601,N_33735);
xor U34466 (N_34466,N_33680,N_33956);
nor U34467 (N_34467,N_33653,N_33632);
nand U34468 (N_34468,N_33953,N_33715);
or U34469 (N_34469,N_33798,N_33563);
and U34470 (N_34470,N_33649,N_33790);
or U34471 (N_34471,N_33691,N_33525);
and U34472 (N_34472,N_33608,N_33995);
nand U34473 (N_34473,N_33950,N_33734);
xnor U34474 (N_34474,N_33728,N_33855);
nor U34475 (N_34475,N_33659,N_33964);
xnor U34476 (N_34476,N_33933,N_33690);
nand U34477 (N_34477,N_33573,N_33541);
nor U34478 (N_34478,N_33644,N_33782);
nand U34479 (N_34479,N_33940,N_33715);
nor U34480 (N_34480,N_33701,N_33607);
xor U34481 (N_34481,N_33533,N_33638);
nor U34482 (N_34482,N_33523,N_33513);
nand U34483 (N_34483,N_33969,N_33618);
or U34484 (N_34484,N_33629,N_33867);
and U34485 (N_34485,N_33950,N_33961);
nand U34486 (N_34486,N_33912,N_33501);
and U34487 (N_34487,N_33835,N_33507);
and U34488 (N_34488,N_33693,N_33525);
nand U34489 (N_34489,N_33504,N_33984);
xor U34490 (N_34490,N_33675,N_33895);
nor U34491 (N_34491,N_33689,N_33634);
nor U34492 (N_34492,N_33813,N_33730);
nand U34493 (N_34493,N_33519,N_33550);
and U34494 (N_34494,N_33871,N_33979);
xnor U34495 (N_34495,N_33516,N_33662);
xor U34496 (N_34496,N_33679,N_33500);
or U34497 (N_34497,N_33663,N_33754);
nand U34498 (N_34498,N_33678,N_33677);
and U34499 (N_34499,N_33598,N_33850);
or U34500 (N_34500,N_34388,N_34319);
and U34501 (N_34501,N_34241,N_34038);
or U34502 (N_34502,N_34117,N_34178);
xor U34503 (N_34503,N_34225,N_34105);
or U34504 (N_34504,N_34061,N_34018);
and U34505 (N_34505,N_34145,N_34308);
or U34506 (N_34506,N_34416,N_34402);
xnor U34507 (N_34507,N_34429,N_34498);
or U34508 (N_34508,N_34005,N_34185);
or U34509 (N_34509,N_34365,N_34484);
nand U34510 (N_34510,N_34163,N_34397);
and U34511 (N_34511,N_34435,N_34093);
xnor U34512 (N_34512,N_34266,N_34291);
nor U34513 (N_34513,N_34347,N_34286);
xor U34514 (N_34514,N_34133,N_34425);
nor U34515 (N_34515,N_34218,N_34016);
xnor U34516 (N_34516,N_34369,N_34125);
and U34517 (N_34517,N_34153,N_34334);
xnor U34518 (N_34518,N_34219,N_34022);
nand U34519 (N_34519,N_34254,N_34462);
nand U34520 (N_34520,N_34030,N_34460);
and U34521 (N_34521,N_34345,N_34231);
nand U34522 (N_34522,N_34193,N_34172);
nand U34523 (N_34523,N_34183,N_34141);
or U34524 (N_34524,N_34168,N_34344);
nand U34525 (N_34525,N_34041,N_34333);
xnor U34526 (N_34526,N_34026,N_34098);
xnor U34527 (N_34527,N_34048,N_34322);
nor U34528 (N_34528,N_34451,N_34332);
nand U34529 (N_34529,N_34027,N_34213);
or U34530 (N_34530,N_34494,N_34216);
xnor U34531 (N_34531,N_34062,N_34427);
xnor U34532 (N_34532,N_34203,N_34471);
nand U34533 (N_34533,N_34276,N_34130);
xor U34534 (N_34534,N_34326,N_34400);
or U34535 (N_34535,N_34491,N_34487);
nor U34536 (N_34536,N_34051,N_34407);
or U34537 (N_34537,N_34211,N_34055);
xor U34538 (N_34538,N_34449,N_34302);
and U34539 (N_34539,N_34077,N_34132);
and U34540 (N_34540,N_34127,N_34476);
and U34541 (N_34541,N_34012,N_34474);
nor U34542 (N_34542,N_34379,N_34088);
xnor U34543 (N_34543,N_34492,N_34089);
and U34544 (N_34544,N_34257,N_34010);
or U34545 (N_34545,N_34123,N_34238);
and U34546 (N_34546,N_34034,N_34387);
nand U34547 (N_34547,N_34318,N_34497);
or U34548 (N_34548,N_34043,N_34170);
or U34549 (N_34549,N_34057,N_34430);
or U34550 (N_34550,N_34152,N_34229);
nand U34551 (N_34551,N_34470,N_34140);
and U34552 (N_34552,N_34118,N_34066);
and U34553 (N_34553,N_34409,N_34015);
and U34554 (N_34554,N_34155,N_34299);
xor U34555 (N_34555,N_34348,N_34252);
or U34556 (N_34556,N_34280,N_34253);
nor U34557 (N_34557,N_34190,N_34174);
or U34558 (N_34558,N_34298,N_34372);
nand U34559 (N_34559,N_34068,N_34184);
nand U34560 (N_34560,N_34380,N_34354);
or U34561 (N_34561,N_34385,N_34273);
nor U34562 (N_34562,N_34272,N_34281);
or U34563 (N_34563,N_34264,N_34311);
nor U34564 (N_34564,N_34381,N_34108);
or U34565 (N_34565,N_34075,N_34176);
nand U34566 (N_34566,N_34056,N_34021);
xor U34567 (N_34567,N_34432,N_34485);
nand U34568 (N_34568,N_34410,N_34481);
or U34569 (N_34569,N_34244,N_34070);
nand U34570 (N_34570,N_34232,N_34148);
and U34571 (N_34571,N_34301,N_34074);
nor U34572 (N_34572,N_34175,N_34204);
or U34573 (N_34573,N_34182,N_34001);
nand U34574 (N_34574,N_34437,N_34292);
and U34575 (N_34575,N_34220,N_34275);
nand U34576 (N_34576,N_34064,N_34459);
and U34577 (N_34577,N_34303,N_34147);
nand U34578 (N_34578,N_34233,N_34360);
xor U34579 (N_34579,N_34134,N_34346);
nand U34580 (N_34580,N_34414,N_34124);
xor U34581 (N_34581,N_34479,N_34042);
or U34582 (N_34582,N_34161,N_34000);
or U34583 (N_34583,N_34046,N_34054);
or U34584 (N_34584,N_34404,N_34423);
or U34585 (N_34585,N_34063,N_34353);
nor U34586 (N_34586,N_34405,N_34305);
nand U34587 (N_34587,N_34463,N_34329);
xnor U34588 (N_34588,N_34300,N_34251);
and U34589 (N_34589,N_34059,N_34217);
and U34590 (N_34590,N_34448,N_34455);
nor U34591 (N_34591,N_34413,N_34428);
or U34592 (N_34592,N_34047,N_34293);
or U34593 (N_34593,N_34477,N_34031);
xor U34594 (N_34594,N_34114,N_34071);
and U34595 (N_34595,N_34079,N_34028);
nand U34596 (N_34596,N_34260,N_34446);
nor U34597 (N_34597,N_34321,N_34313);
or U34598 (N_34598,N_34396,N_34136);
or U34599 (N_34599,N_34151,N_34073);
or U34600 (N_34600,N_34106,N_34095);
nand U34601 (N_34601,N_34137,N_34436);
xor U34602 (N_34602,N_34156,N_34109);
nand U34603 (N_34603,N_34146,N_34110);
or U34604 (N_34604,N_34103,N_34149);
or U34605 (N_34605,N_34189,N_34475);
or U34606 (N_34606,N_34392,N_34165);
and U34607 (N_34607,N_34316,N_34102);
xor U34608 (N_34608,N_34008,N_34327);
and U34609 (N_34609,N_34086,N_34131);
or U34610 (N_34610,N_34119,N_34128);
xnor U34611 (N_34611,N_34227,N_34209);
nor U34612 (N_34612,N_34269,N_34235);
nor U34613 (N_34613,N_34310,N_34389);
xor U34614 (N_34614,N_34457,N_34226);
and U34615 (N_34615,N_34143,N_34004);
nand U34616 (N_34616,N_34036,N_34072);
or U34617 (N_34617,N_34014,N_34472);
nor U34618 (N_34618,N_34403,N_34371);
or U34619 (N_34619,N_34139,N_34282);
or U34620 (N_34620,N_34395,N_34297);
nor U34621 (N_34621,N_34179,N_34447);
xor U34622 (N_34622,N_34242,N_34493);
nor U34623 (N_34623,N_34285,N_34196);
nand U34624 (N_34624,N_34222,N_34386);
nor U34625 (N_34625,N_34058,N_34412);
xnor U34626 (N_34626,N_34115,N_34420);
nand U34627 (N_34627,N_34091,N_34011);
nand U34628 (N_34628,N_34100,N_34456);
and U34629 (N_34629,N_34249,N_34052);
or U34630 (N_34630,N_34339,N_34443);
xor U34631 (N_34631,N_34408,N_34374);
xnor U34632 (N_34632,N_34101,N_34158);
nand U34633 (N_34633,N_34200,N_34246);
nor U34634 (N_34634,N_34349,N_34078);
nor U34635 (N_34635,N_34169,N_34096);
nor U34636 (N_34636,N_34419,N_34421);
or U34637 (N_34637,N_34482,N_34489);
xor U34638 (N_34638,N_34035,N_34138);
nand U34639 (N_34639,N_34364,N_34069);
nor U34640 (N_34640,N_34480,N_34076);
or U34641 (N_34641,N_34129,N_34445);
xnor U34642 (N_34642,N_34186,N_34243);
xor U34643 (N_34643,N_34325,N_34007);
or U34644 (N_34644,N_34167,N_34496);
and U34645 (N_34645,N_34391,N_34331);
nand U34646 (N_34646,N_34373,N_34262);
xnor U34647 (N_34647,N_34083,N_34469);
xnor U34648 (N_34648,N_34324,N_34126);
or U34649 (N_34649,N_34320,N_34221);
and U34650 (N_34650,N_34290,N_34006);
nor U34651 (N_34651,N_34017,N_34122);
nor U34652 (N_34652,N_34278,N_34053);
and U34653 (N_34653,N_34444,N_34433);
or U34654 (N_34654,N_34092,N_34120);
or U34655 (N_34655,N_34442,N_34426);
xor U34656 (N_34656,N_34368,N_34240);
and U34657 (N_34657,N_34084,N_34314);
nand U34658 (N_34658,N_34236,N_34247);
or U34659 (N_34659,N_34341,N_34309);
and U34660 (N_34660,N_34452,N_34343);
nor U34661 (N_34661,N_34081,N_34111);
and U34662 (N_34662,N_34085,N_34488);
and U34663 (N_34663,N_34363,N_34224);
or U34664 (N_34664,N_34206,N_34037);
and U34665 (N_34665,N_34090,N_34104);
and U34666 (N_34666,N_34376,N_34112);
and U34667 (N_34667,N_34323,N_34060);
and U34668 (N_34668,N_34020,N_34306);
and U34669 (N_34669,N_34356,N_34362);
and U34670 (N_34670,N_34082,N_34289);
and U34671 (N_34671,N_34013,N_34099);
xnor U34672 (N_34672,N_34268,N_34390);
nand U34673 (N_34673,N_34359,N_34144);
nor U34674 (N_34674,N_34384,N_34050);
xnor U34675 (N_34675,N_34208,N_34044);
and U34676 (N_34676,N_34187,N_34166);
and U34677 (N_34677,N_34230,N_34003);
or U34678 (N_34678,N_34304,N_34228);
or U34679 (N_34679,N_34258,N_34202);
or U34680 (N_34680,N_34248,N_34270);
and U34681 (N_34681,N_34205,N_34094);
or U34682 (N_34682,N_34067,N_34181);
or U34683 (N_34683,N_34337,N_34024);
nor U34684 (N_34684,N_34340,N_34483);
nand U34685 (N_34685,N_34355,N_34366);
or U34686 (N_34686,N_34195,N_34032);
and U34687 (N_34687,N_34250,N_34180);
nor U34688 (N_34688,N_34335,N_34431);
nand U34689 (N_34689,N_34116,N_34361);
nand U34690 (N_34690,N_34440,N_34450);
and U34691 (N_34691,N_34065,N_34490);
nand U34692 (N_34692,N_34256,N_34214);
nand U34693 (N_34693,N_34342,N_34375);
nor U34694 (N_34694,N_34296,N_34350);
nand U34695 (N_34695,N_34192,N_34173);
xor U34696 (N_34696,N_34045,N_34411);
or U34697 (N_34697,N_34194,N_34157);
or U34698 (N_34698,N_34338,N_34422);
and U34699 (N_34699,N_34277,N_34121);
nand U34700 (N_34700,N_34191,N_34215);
or U34701 (N_34701,N_34312,N_34199);
nor U34702 (N_34702,N_34142,N_34162);
nand U34703 (N_34703,N_34415,N_34239);
and U34704 (N_34704,N_34287,N_34009);
and U34705 (N_34705,N_34439,N_34087);
or U34706 (N_34706,N_34468,N_34378);
and U34707 (N_34707,N_34033,N_34473);
nand U34708 (N_34708,N_34499,N_34466);
nand U34709 (N_34709,N_34288,N_34352);
xnor U34710 (N_34710,N_34398,N_34358);
xor U34711 (N_34711,N_34259,N_34406);
and U34712 (N_34712,N_34025,N_34164);
and U34713 (N_34713,N_34295,N_34367);
or U34714 (N_34714,N_34495,N_34255);
xor U34715 (N_34715,N_34261,N_34237);
nand U34716 (N_34716,N_34267,N_34002);
or U34717 (N_34717,N_34317,N_34461);
xnor U34718 (N_34718,N_34245,N_34434);
nor U34719 (N_34719,N_34150,N_34154);
or U34720 (N_34720,N_34464,N_34351);
nor U34721 (N_34721,N_34159,N_34486);
and U34722 (N_34722,N_34370,N_34171);
xor U34723 (N_34723,N_34188,N_34336);
or U34724 (N_34724,N_34113,N_34274);
or U34725 (N_34725,N_34198,N_34441);
xor U34726 (N_34726,N_34307,N_34418);
nand U34727 (N_34727,N_34453,N_34107);
and U34728 (N_34728,N_34284,N_34049);
and U34729 (N_34729,N_34382,N_34424);
and U34730 (N_34730,N_34330,N_34399);
nor U34731 (N_34731,N_34454,N_34315);
nand U34732 (N_34732,N_34458,N_34263);
nor U34733 (N_34733,N_34478,N_34383);
nor U34734 (N_34734,N_34283,N_34039);
xor U34735 (N_34735,N_34223,N_34357);
nand U34736 (N_34736,N_34294,N_34265);
nor U34737 (N_34737,N_34465,N_34393);
xor U34738 (N_34738,N_34040,N_34328);
nand U34739 (N_34739,N_34212,N_34177);
nand U34740 (N_34740,N_34023,N_34210);
nand U34741 (N_34741,N_34401,N_34097);
and U34742 (N_34742,N_34467,N_34377);
nand U34743 (N_34743,N_34029,N_34201);
and U34744 (N_34744,N_34160,N_34438);
and U34745 (N_34745,N_34417,N_34080);
nor U34746 (N_34746,N_34135,N_34207);
xnor U34747 (N_34747,N_34234,N_34271);
xor U34748 (N_34748,N_34019,N_34197);
and U34749 (N_34749,N_34394,N_34279);
xnor U34750 (N_34750,N_34347,N_34260);
and U34751 (N_34751,N_34333,N_34173);
nand U34752 (N_34752,N_34396,N_34117);
xnor U34753 (N_34753,N_34117,N_34429);
nor U34754 (N_34754,N_34184,N_34220);
nor U34755 (N_34755,N_34376,N_34478);
nand U34756 (N_34756,N_34300,N_34383);
and U34757 (N_34757,N_34399,N_34451);
nand U34758 (N_34758,N_34172,N_34097);
nand U34759 (N_34759,N_34484,N_34336);
nor U34760 (N_34760,N_34253,N_34000);
xnor U34761 (N_34761,N_34478,N_34270);
nor U34762 (N_34762,N_34474,N_34470);
or U34763 (N_34763,N_34037,N_34238);
or U34764 (N_34764,N_34327,N_34305);
and U34765 (N_34765,N_34305,N_34217);
or U34766 (N_34766,N_34342,N_34063);
nor U34767 (N_34767,N_34399,N_34231);
or U34768 (N_34768,N_34237,N_34319);
nand U34769 (N_34769,N_34058,N_34155);
nor U34770 (N_34770,N_34122,N_34121);
or U34771 (N_34771,N_34052,N_34427);
nor U34772 (N_34772,N_34265,N_34290);
or U34773 (N_34773,N_34234,N_34001);
nor U34774 (N_34774,N_34043,N_34461);
and U34775 (N_34775,N_34181,N_34420);
or U34776 (N_34776,N_34075,N_34358);
nor U34777 (N_34777,N_34245,N_34169);
xnor U34778 (N_34778,N_34293,N_34421);
nand U34779 (N_34779,N_34127,N_34488);
and U34780 (N_34780,N_34205,N_34426);
or U34781 (N_34781,N_34238,N_34153);
nor U34782 (N_34782,N_34071,N_34085);
or U34783 (N_34783,N_34413,N_34068);
or U34784 (N_34784,N_34193,N_34012);
nand U34785 (N_34785,N_34221,N_34443);
or U34786 (N_34786,N_34275,N_34492);
xor U34787 (N_34787,N_34124,N_34453);
and U34788 (N_34788,N_34143,N_34267);
or U34789 (N_34789,N_34342,N_34228);
nor U34790 (N_34790,N_34077,N_34235);
nor U34791 (N_34791,N_34304,N_34115);
nor U34792 (N_34792,N_34198,N_34162);
and U34793 (N_34793,N_34048,N_34098);
nand U34794 (N_34794,N_34442,N_34260);
xor U34795 (N_34795,N_34335,N_34142);
xnor U34796 (N_34796,N_34168,N_34062);
and U34797 (N_34797,N_34175,N_34178);
nand U34798 (N_34798,N_34235,N_34134);
or U34799 (N_34799,N_34481,N_34360);
nand U34800 (N_34800,N_34498,N_34334);
or U34801 (N_34801,N_34214,N_34412);
or U34802 (N_34802,N_34147,N_34100);
nand U34803 (N_34803,N_34030,N_34036);
xnor U34804 (N_34804,N_34476,N_34244);
or U34805 (N_34805,N_34490,N_34274);
nor U34806 (N_34806,N_34221,N_34099);
or U34807 (N_34807,N_34252,N_34441);
nor U34808 (N_34808,N_34218,N_34199);
nand U34809 (N_34809,N_34130,N_34413);
and U34810 (N_34810,N_34046,N_34133);
nor U34811 (N_34811,N_34266,N_34261);
or U34812 (N_34812,N_34237,N_34219);
and U34813 (N_34813,N_34068,N_34178);
nor U34814 (N_34814,N_34037,N_34358);
xor U34815 (N_34815,N_34178,N_34288);
xor U34816 (N_34816,N_34055,N_34283);
xor U34817 (N_34817,N_34297,N_34158);
nor U34818 (N_34818,N_34285,N_34151);
or U34819 (N_34819,N_34233,N_34381);
xor U34820 (N_34820,N_34085,N_34295);
and U34821 (N_34821,N_34376,N_34046);
and U34822 (N_34822,N_34184,N_34377);
or U34823 (N_34823,N_34356,N_34411);
and U34824 (N_34824,N_34080,N_34009);
xnor U34825 (N_34825,N_34344,N_34147);
nor U34826 (N_34826,N_34417,N_34098);
nand U34827 (N_34827,N_34193,N_34044);
or U34828 (N_34828,N_34397,N_34279);
and U34829 (N_34829,N_34233,N_34366);
and U34830 (N_34830,N_34181,N_34212);
and U34831 (N_34831,N_34083,N_34084);
or U34832 (N_34832,N_34247,N_34372);
or U34833 (N_34833,N_34282,N_34180);
or U34834 (N_34834,N_34065,N_34157);
nor U34835 (N_34835,N_34322,N_34397);
nand U34836 (N_34836,N_34006,N_34498);
nand U34837 (N_34837,N_34019,N_34337);
nor U34838 (N_34838,N_34034,N_34399);
or U34839 (N_34839,N_34329,N_34194);
xnor U34840 (N_34840,N_34391,N_34399);
xnor U34841 (N_34841,N_34123,N_34433);
and U34842 (N_34842,N_34369,N_34346);
or U34843 (N_34843,N_34147,N_34007);
or U34844 (N_34844,N_34385,N_34365);
xnor U34845 (N_34845,N_34318,N_34439);
or U34846 (N_34846,N_34378,N_34489);
nand U34847 (N_34847,N_34177,N_34472);
nor U34848 (N_34848,N_34083,N_34279);
nand U34849 (N_34849,N_34249,N_34224);
or U34850 (N_34850,N_34128,N_34103);
nand U34851 (N_34851,N_34078,N_34047);
or U34852 (N_34852,N_34488,N_34157);
or U34853 (N_34853,N_34366,N_34252);
or U34854 (N_34854,N_34273,N_34028);
xnor U34855 (N_34855,N_34362,N_34206);
and U34856 (N_34856,N_34064,N_34374);
xor U34857 (N_34857,N_34089,N_34431);
nand U34858 (N_34858,N_34455,N_34406);
and U34859 (N_34859,N_34397,N_34355);
nand U34860 (N_34860,N_34493,N_34024);
nor U34861 (N_34861,N_34138,N_34258);
xor U34862 (N_34862,N_34091,N_34258);
and U34863 (N_34863,N_34342,N_34469);
or U34864 (N_34864,N_34369,N_34442);
or U34865 (N_34865,N_34411,N_34228);
nor U34866 (N_34866,N_34347,N_34470);
nand U34867 (N_34867,N_34363,N_34209);
or U34868 (N_34868,N_34146,N_34325);
nand U34869 (N_34869,N_34190,N_34055);
xnor U34870 (N_34870,N_34060,N_34272);
nor U34871 (N_34871,N_34113,N_34484);
nand U34872 (N_34872,N_34080,N_34342);
nand U34873 (N_34873,N_34438,N_34487);
xor U34874 (N_34874,N_34253,N_34461);
and U34875 (N_34875,N_34305,N_34055);
nor U34876 (N_34876,N_34295,N_34002);
or U34877 (N_34877,N_34471,N_34255);
or U34878 (N_34878,N_34068,N_34275);
or U34879 (N_34879,N_34101,N_34354);
or U34880 (N_34880,N_34094,N_34482);
xnor U34881 (N_34881,N_34344,N_34491);
and U34882 (N_34882,N_34307,N_34434);
nor U34883 (N_34883,N_34353,N_34278);
xnor U34884 (N_34884,N_34365,N_34085);
xor U34885 (N_34885,N_34302,N_34181);
or U34886 (N_34886,N_34344,N_34237);
or U34887 (N_34887,N_34303,N_34270);
nand U34888 (N_34888,N_34489,N_34019);
and U34889 (N_34889,N_34384,N_34483);
or U34890 (N_34890,N_34498,N_34111);
nand U34891 (N_34891,N_34314,N_34480);
and U34892 (N_34892,N_34100,N_34027);
xnor U34893 (N_34893,N_34029,N_34495);
xnor U34894 (N_34894,N_34280,N_34078);
nor U34895 (N_34895,N_34178,N_34495);
nand U34896 (N_34896,N_34397,N_34089);
or U34897 (N_34897,N_34076,N_34359);
nor U34898 (N_34898,N_34397,N_34346);
xor U34899 (N_34899,N_34285,N_34437);
or U34900 (N_34900,N_34151,N_34421);
and U34901 (N_34901,N_34468,N_34228);
xnor U34902 (N_34902,N_34214,N_34239);
nand U34903 (N_34903,N_34072,N_34308);
nor U34904 (N_34904,N_34284,N_34153);
nand U34905 (N_34905,N_34089,N_34382);
nand U34906 (N_34906,N_34194,N_34225);
nand U34907 (N_34907,N_34327,N_34292);
or U34908 (N_34908,N_34284,N_34350);
xor U34909 (N_34909,N_34080,N_34259);
or U34910 (N_34910,N_34200,N_34261);
or U34911 (N_34911,N_34200,N_34242);
xor U34912 (N_34912,N_34277,N_34323);
nor U34913 (N_34913,N_34232,N_34367);
nand U34914 (N_34914,N_34184,N_34348);
nand U34915 (N_34915,N_34149,N_34248);
and U34916 (N_34916,N_34076,N_34416);
and U34917 (N_34917,N_34167,N_34221);
and U34918 (N_34918,N_34086,N_34429);
nand U34919 (N_34919,N_34291,N_34450);
nand U34920 (N_34920,N_34362,N_34303);
nor U34921 (N_34921,N_34341,N_34499);
nand U34922 (N_34922,N_34139,N_34008);
xor U34923 (N_34923,N_34124,N_34054);
xnor U34924 (N_34924,N_34169,N_34006);
and U34925 (N_34925,N_34260,N_34136);
nor U34926 (N_34926,N_34327,N_34155);
nand U34927 (N_34927,N_34363,N_34099);
nor U34928 (N_34928,N_34221,N_34183);
or U34929 (N_34929,N_34383,N_34258);
nand U34930 (N_34930,N_34465,N_34213);
or U34931 (N_34931,N_34189,N_34217);
and U34932 (N_34932,N_34457,N_34325);
nand U34933 (N_34933,N_34330,N_34343);
nand U34934 (N_34934,N_34016,N_34226);
or U34935 (N_34935,N_34085,N_34451);
or U34936 (N_34936,N_34189,N_34282);
or U34937 (N_34937,N_34158,N_34454);
or U34938 (N_34938,N_34266,N_34037);
nand U34939 (N_34939,N_34349,N_34347);
xnor U34940 (N_34940,N_34229,N_34261);
xnor U34941 (N_34941,N_34125,N_34016);
nor U34942 (N_34942,N_34072,N_34236);
and U34943 (N_34943,N_34477,N_34371);
xor U34944 (N_34944,N_34465,N_34377);
nor U34945 (N_34945,N_34013,N_34086);
nand U34946 (N_34946,N_34343,N_34113);
or U34947 (N_34947,N_34310,N_34453);
and U34948 (N_34948,N_34212,N_34486);
and U34949 (N_34949,N_34397,N_34140);
or U34950 (N_34950,N_34334,N_34470);
xor U34951 (N_34951,N_34044,N_34124);
nor U34952 (N_34952,N_34423,N_34362);
or U34953 (N_34953,N_34423,N_34015);
and U34954 (N_34954,N_34010,N_34253);
xor U34955 (N_34955,N_34099,N_34269);
nor U34956 (N_34956,N_34465,N_34102);
nand U34957 (N_34957,N_34304,N_34075);
nand U34958 (N_34958,N_34241,N_34451);
or U34959 (N_34959,N_34149,N_34402);
nor U34960 (N_34960,N_34169,N_34486);
and U34961 (N_34961,N_34219,N_34449);
or U34962 (N_34962,N_34100,N_34148);
nor U34963 (N_34963,N_34254,N_34027);
nor U34964 (N_34964,N_34412,N_34497);
and U34965 (N_34965,N_34397,N_34289);
xnor U34966 (N_34966,N_34036,N_34461);
and U34967 (N_34967,N_34029,N_34008);
or U34968 (N_34968,N_34406,N_34015);
nand U34969 (N_34969,N_34364,N_34025);
or U34970 (N_34970,N_34012,N_34313);
nand U34971 (N_34971,N_34417,N_34470);
and U34972 (N_34972,N_34121,N_34465);
and U34973 (N_34973,N_34224,N_34047);
and U34974 (N_34974,N_34025,N_34252);
nor U34975 (N_34975,N_34308,N_34252);
xor U34976 (N_34976,N_34448,N_34301);
xnor U34977 (N_34977,N_34433,N_34401);
nor U34978 (N_34978,N_34386,N_34478);
xnor U34979 (N_34979,N_34041,N_34363);
or U34980 (N_34980,N_34212,N_34363);
nor U34981 (N_34981,N_34197,N_34233);
nor U34982 (N_34982,N_34175,N_34196);
nor U34983 (N_34983,N_34219,N_34088);
and U34984 (N_34984,N_34045,N_34315);
nand U34985 (N_34985,N_34039,N_34128);
xnor U34986 (N_34986,N_34381,N_34488);
or U34987 (N_34987,N_34246,N_34382);
xnor U34988 (N_34988,N_34087,N_34442);
nor U34989 (N_34989,N_34403,N_34437);
nor U34990 (N_34990,N_34260,N_34216);
or U34991 (N_34991,N_34080,N_34422);
nor U34992 (N_34992,N_34394,N_34016);
and U34993 (N_34993,N_34298,N_34491);
nor U34994 (N_34994,N_34080,N_34296);
and U34995 (N_34995,N_34052,N_34252);
xnor U34996 (N_34996,N_34132,N_34293);
or U34997 (N_34997,N_34344,N_34432);
xor U34998 (N_34998,N_34109,N_34172);
nor U34999 (N_34999,N_34043,N_34428);
or U35000 (N_35000,N_34675,N_34897);
nand U35001 (N_35001,N_34545,N_34957);
and U35002 (N_35002,N_34583,N_34525);
and U35003 (N_35003,N_34782,N_34935);
and U35004 (N_35004,N_34730,N_34997);
xor U35005 (N_35005,N_34951,N_34960);
or U35006 (N_35006,N_34958,N_34631);
xnor U35007 (N_35007,N_34939,N_34885);
or U35008 (N_35008,N_34769,N_34875);
or U35009 (N_35009,N_34637,N_34509);
nand U35010 (N_35010,N_34688,N_34702);
and U35011 (N_35011,N_34975,N_34953);
xnor U35012 (N_35012,N_34766,N_34629);
nor U35013 (N_35013,N_34523,N_34536);
or U35014 (N_35014,N_34836,N_34661);
nor U35015 (N_35015,N_34589,N_34703);
nor U35016 (N_35016,N_34850,N_34669);
xnor U35017 (N_35017,N_34848,N_34639);
or U35018 (N_35018,N_34713,N_34944);
or U35019 (N_35019,N_34711,N_34548);
xor U35020 (N_35020,N_34514,N_34898);
or U35021 (N_35021,N_34526,N_34866);
or U35022 (N_35022,N_34585,N_34687);
or U35023 (N_35023,N_34858,N_34716);
or U35024 (N_35024,N_34588,N_34881);
xor U35025 (N_35025,N_34746,N_34946);
xnor U35026 (N_35026,N_34783,N_34582);
nor U35027 (N_35027,N_34749,N_34581);
or U35028 (N_35028,N_34718,N_34643);
and U35029 (N_35029,N_34814,N_34940);
nor U35030 (N_35030,N_34507,N_34872);
and U35031 (N_35031,N_34697,N_34627);
and U35032 (N_35032,N_34560,N_34715);
nand U35033 (N_35033,N_34758,N_34936);
nand U35034 (N_35034,N_34739,N_34677);
xor U35035 (N_35035,N_34787,N_34654);
nor U35036 (N_35036,N_34924,N_34923);
xnor U35037 (N_35037,N_34994,N_34541);
and U35038 (N_35038,N_34705,N_34538);
or U35039 (N_35039,N_34986,N_34554);
or U35040 (N_35040,N_34889,N_34655);
nor U35041 (N_35041,N_34645,N_34922);
nor U35042 (N_35042,N_34547,N_34807);
and U35043 (N_35043,N_34828,N_34522);
nand U35044 (N_35044,N_34999,N_34993);
nand U35045 (N_35045,N_34719,N_34860);
and U35046 (N_35046,N_34604,N_34985);
or U35047 (N_35047,N_34603,N_34616);
or U35048 (N_35048,N_34950,N_34911);
nand U35049 (N_35049,N_34597,N_34626);
or U35050 (N_35050,N_34884,N_34969);
or U35051 (N_35051,N_34930,N_34903);
nor U35052 (N_35052,N_34696,N_34537);
nand U35053 (N_35053,N_34874,N_34992);
xnor U35054 (N_35054,N_34796,N_34617);
and U35055 (N_35055,N_34891,N_34967);
xnor U35056 (N_35056,N_34651,N_34593);
and U35057 (N_35057,N_34972,N_34785);
nor U35058 (N_35058,N_34671,N_34952);
nand U35059 (N_35059,N_34750,N_34938);
nand U35060 (N_35060,N_34596,N_34945);
xnor U35061 (N_35061,N_34727,N_34744);
and U35062 (N_35062,N_34693,N_34808);
and U35063 (N_35063,N_34724,N_34592);
nor U35064 (N_35064,N_34587,N_34809);
xnor U35065 (N_35065,N_34852,N_34855);
nand U35066 (N_35066,N_34909,N_34733);
nand U35067 (N_35067,N_34558,N_34735);
and U35068 (N_35068,N_34729,N_34542);
nand U35069 (N_35069,N_34820,N_34899);
and U35070 (N_35070,N_34646,N_34919);
nand U35071 (N_35071,N_34510,N_34965);
nor U35072 (N_35072,N_34833,N_34811);
and U35073 (N_35073,N_34741,N_34608);
xor U35074 (N_35074,N_34759,N_34680);
nor U35075 (N_35075,N_34734,N_34941);
nor U35076 (N_35076,N_34664,N_34802);
or U35077 (N_35077,N_34534,N_34557);
xnor U35078 (N_35078,N_34863,N_34544);
nor U35079 (N_35079,N_34574,N_34778);
nor U35080 (N_35080,N_34980,N_34956);
xor U35081 (N_35081,N_34673,N_34672);
nor U35082 (N_35082,N_34694,N_34775);
nor U35083 (N_35083,N_34505,N_34652);
xnor U35084 (N_35084,N_34784,N_34779);
nor U35085 (N_35085,N_34754,N_34521);
nor U35086 (N_35086,N_34834,N_34932);
or U35087 (N_35087,N_34789,N_34822);
and U35088 (N_35088,N_34799,N_34798);
nor U35089 (N_35089,N_34854,N_34942);
nand U35090 (N_35090,N_34925,N_34826);
and U35091 (N_35091,N_34690,N_34998);
or U35092 (N_35092,N_34559,N_34732);
nand U35093 (N_35093,N_34600,N_34519);
nor U35094 (N_35094,N_34966,N_34678);
and U35095 (N_35095,N_34937,N_34772);
xnor U35096 (N_35096,N_34692,N_34700);
or U35097 (N_35097,N_34575,N_34663);
or U35098 (N_35098,N_34818,N_34792);
and U35099 (N_35099,N_34615,N_34609);
or U35100 (N_35100,N_34880,N_34816);
or U35101 (N_35101,N_34662,N_34791);
nor U35102 (N_35102,N_34584,N_34679);
xnor U35103 (N_35103,N_34517,N_34709);
and U35104 (N_35104,N_34786,N_34723);
nor U35105 (N_35105,N_34742,N_34862);
and U35106 (N_35106,N_34640,N_34511);
nand U35107 (N_35107,N_34949,N_34931);
or U35108 (N_35108,N_34636,N_34795);
nor U35109 (N_35109,N_34513,N_34920);
nor U35110 (N_35110,N_34685,N_34873);
and U35111 (N_35111,N_34682,N_34977);
nor U35112 (N_35112,N_34926,N_34876);
nand U35113 (N_35113,N_34856,N_34987);
nand U35114 (N_35114,N_34959,N_34883);
xnor U35115 (N_35115,N_34539,N_34890);
nor U35116 (N_35116,N_34817,N_34752);
and U35117 (N_35117,N_34757,N_34740);
xnor U35118 (N_35118,N_34983,N_34841);
nor U35119 (N_35119,N_34503,N_34824);
or U35120 (N_35120,N_34943,N_34823);
and U35121 (N_35121,N_34590,N_34964);
nor U35122 (N_35122,N_34955,N_34530);
and U35123 (N_35123,N_34812,N_34963);
or U35124 (N_35124,N_34668,N_34904);
and U35125 (N_35125,N_34568,N_34755);
or U35126 (N_35126,N_34540,N_34974);
and U35127 (N_35127,N_34586,N_34761);
or U35128 (N_35128,N_34598,N_34832);
xnor U35129 (N_35129,N_34760,N_34599);
and U35130 (N_35130,N_34815,N_34839);
nor U35131 (N_35131,N_34722,N_34861);
and U35132 (N_35132,N_34916,N_34515);
nand U35133 (N_35133,N_34606,N_34518);
xor U35134 (N_35134,N_34857,N_34928);
xor U35135 (N_35135,N_34806,N_34776);
xor U35136 (N_35136,N_34641,N_34929);
or U35137 (N_35137,N_34991,N_34948);
or U35138 (N_35138,N_34647,N_34877);
xor U35139 (N_35139,N_34656,N_34707);
xor U35140 (N_35140,N_34528,N_34632);
and U35141 (N_35141,N_34869,N_34571);
and U35142 (N_35142,N_34622,N_34767);
nor U35143 (N_35143,N_34619,N_34613);
or U35144 (N_35144,N_34895,N_34892);
xnor U35145 (N_35145,N_34610,N_34580);
xnor U35146 (N_35146,N_34745,N_34773);
and U35147 (N_35147,N_34901,N_34710);
or U35148 (N_35148,N_34914,N_34670);
or U35149 (N_35149,N_34982,N_34738);
xor U35150 (N_35150,N_34793,N_34763);
nor U35151 (N_35151,N_34971,N_34549);
or U35152 (N_35152,N_34633,N_34835);
or U35153 (N_35153,N_34804,N_34512);
nand U35154 (N_35154,N_34968,N_34847);
and U35155 (N_35155,N_34748,N_34611);
nand U35156 (N_35156,N_34551,N_34684);
nor U35157 (N_35157,N_34628,N_34658);
xor U35158 (N_35158,N_34996,N_34520);
and U35159 (N_35159,N_34506,N_34780);
nor U35160 (N_35160,N_34659,N_34879);
nand U35161 (N_35161,N_34970,N_34829);
and U35162 (N_35162,N_34726,N_34845);
nor U35163 (N_35163,N_34805,N_34915);
nand U35164 (N_35164,N_34620,N_34594);
nor U35165 (N_35165,N_34908,N_34725);
nand U35166 (N_35166,N_34988,N_34813);
or U35167 (N_35167,N_34790,N_34882);
xor U35168 (N_35168,N_34849,N_34771);
and U35169 (N_35169,N_34774,N_34502);
or U35170 (N_35170,N_34570,N_34764);
nand U35171 (N_35171,N_34720,N_34624);
or U35172 (N_35172,N_34825,N_34762);
xor U35173 (N_35173,N_34995,N_34800);
and U35174 (N_35174,N_34630,N_34644);
nor U35175 (N_35175,N_34698,N_34550);
nor U35176 (N_35176,N_34701,N_34553);
or U35177 (N_35177,N_34578,N_34844);
xnor U35178 (N_35178,N_34567,N_34918);
or U35179 (N_35179,N_34552,N_34973);
or U35180 (N_35180,N_34917,N_34921);
xor U35181 (N_35181,N_34714,N_34532);
xor U35182 (N_35182,N_34635,N_34736);
and U35183 (N_35183,N_34634,N_34712);
xor U35184 (N_35184,N_34667,N_34529);
xor U35185 (N_35185,N_34843,N_34934);
nand U35186 (N_35186,N_34913,N_34878);
and U35187 (N_35187,N_34887,N_34765);
and U35188 (N_35188,N_34660,N_34649);
nor U35189 (N_35189,N_34605,N_34572);
nor U35190 (N_35190,N_34737,N_34674);
nand U35191 (N_35191,N_34810,N_34888);
xnor U35192 (N_35192,N_34827,N_34533);
or U35193 (N_35193,N_34868,N_34867);
xor U35194 (N_35194,N_34546,N_34569);
and U35195 (N_35195,N_34781,N_34900);
xor U35196 (N_35196,N_34601,N_34704);
xnor U35197 (N_35197,N_34543,N_34981);
and U35198 (N_35198,N_34648,N_34770);
nor U35199 (N_35199,N_34556,N_34535);
nand U35200 (N_35200,N_34837,N_34691);
nor U35201 (N_35201,N_34984,N_34853);
xnor U35202 (N_35202,N_34666,N_34902);
xnor U35203 (N_35203,N_34527,N_34650);
nand U35204 (N_35204,N_34563,N_34896);
nor U35205 (N_35205,N_34642,N_34794);
xnor U35206 (N_35206,N_34595,N_34625);
and U35207 (N_35207,N_34989,N_34504);
and U35208 (N_35208,N_34508,N_34706);
and U35209 (N_35209,N_34699,N_34683);
nand U35210 (N_35210,N_34927,N_34728);
xor U35211 (N_35211,N_34905,N_34933);
nor U35212 (N_35212,N_34865,N_34747);
and U35213 (N_35213,N_34797,N_34717);
nand U35214 (N_35214,N_34954,N_34708);
nor U35215 (N_35215,N_34566,N_34821);
or U35216 (N_35216,N_34607,N_34777);
and U35217 (N_35217,N_34564,N_34689);
or U35218 (N_35218,N_34756,N_34962);
xor U35219 (N_35219,N_34819,N_34907);
nor U35220 (N_35220,N_34602,N_34579);
and U35221 (N_35221,N_34838,N_34831);
nor U35222 (N_35222,N_34576,N_34731);
xnor U35223 (N_35223,N_34686,N_34990);
xnor U35224 (N_35224,N_34681,N_34864);
xor U35225 (N_35225,N_34653,N_34591);
xnor U35226 (N_35226,N_34501,N_34638);
and U35227 (N_35227,N_34803,N_34976);
and U35228 (N_35228,N_34573,N_34614);
and U35229 (N_35229,N_34840,N_34859);
xnor U35230 (N_35230,N_34721,N_34665);
nor U35231 (N_35231,N_34516,N_34612);
xnor U35232 (N_35232,N_34531,N_34978);
xor U35233 (N_35233,N_34561,N_34618);
xnor U35234 (N_35234,N_34621,N_34893);
nand U35235 (N_35235,N_34743,N_34842);
nor U35236 (N_35236,N_34947,N_34768);
and U35237 (N_35237,N_34870,N_34524);
xor U35238 (N_35238,N_34912,N_34565);
and U35239 (N_35239,N_34830,N_34577);
xnor U35240 (N_35240,N_34753,N_34886);
xnor U35241 (N_35241,N_34695,N_34788);
or U35242 (N_35242,N_34751,N_34500);
and U35243 (N_35243,N_34623,N_34906);
nand U35244 (N_35244,N_34676,N_34801);
nand U35245 (N_35245,N_34979,N_34657);
and U35246 (N_35246,N_34894,N_34562);
xnor U35247 (N_35247,N_34851,N_34555);
nand U35248 (N_35248,N_34871,N_34910);
and U35249 (N_35249,N_34846,N_34961);
nor U35250 (N_35250,N_34685,N_34699);
nand U35251 (N_35251,N_34735,N_34907);
and U35252 (N_35252,N_34534,N_34532);
nand U35253 (N_35253,N_34533,N_34570);
and U35254 (N_35254,N_34654,N_34801);
xnor U35255 (N_35255,N_34662,N_34796);
and U35256 (N_35256,N_34640,N_34658);
or U35257 (N_35257,N_34831,N_34961);
or U35258 (N_35258,N_34766,N_34931);
and U35259 (N_35259,N_34996,N_34873);
or U35260 (N_35260,N_34991,N_34524);
and U35261 (N_35261,N_34873,N_34939);
xor U35262 (N_35262,N_34571,N_34757);
or U35263 (N_35263,N_34972,N_34545);
nor U35264 (N_35264,N_34717,N_34755);
xor U35265 (N_35265,N_34522,N_34904);
nand U35266 (N_35266,N_34804,N_34814);
and U35267 (N_35267,N_34635,N_34752);
and U35268 (N_35268,N_34873,N_34740);
nor U35269 (N_35269,N_34838,N_34902);
xor U35270 (N_35270,N_34792,N_34645);
or U35271 (N_35271,N_34505,N_34893);
xnor U35272 (N_35272,N_34886,N_34675);
xnor U35273 (N_35273,N_34741,N_34897);
and U35274 (N_35274,N_34916,N_34812);
or U35275 (N_35275,N_34862,N_34654);
or U35276 (N_35276,N_34843,N_34504);
and U35277 (N_35277,N_34741,N_34794);
or U35278 (N_35278,N_34653,N_34864);
or U35279 (N_35279,N_34992,N_34627);
xnor U35280 (N_35280,N_34538,N_34659);
or U35281 (N_35281,N_34800,N_34812);
or U35282 (N_35282,N_34940,N_34863);
nor U35283 (N_35283,N_34703,N_34637);
xnor U35284 (N_35284,N_34828,N_34796);
nor U35285 (N_35285,N_34911,N_34760);
or U35286 (N_35286,N_34668,N_34564);
nor U35287 (N_35287,N_34778,N_34684);
nor U35288 (N_35288,N_34571,N_34549);
or U35289 (N_35289,N_34912,N_34708);
and U35290 (N_35290,N_34895,N_34796);
or U35291 (N_35291,N_34510,N_34728);
or U35292 (N_35292,N_34615,N_34857);
nand U35293 (N_35293,N_34619,N_34786);
nor U35294 (N_35294,N_34899,N_34905);
xnor U35295 (N_35295,N_34829,N_34615);
nor U35296 (N_35296,N_34621,N_34851);
or U35297 (N_35297,N_34774,N_34696);
or U35298 (N_35298,N_34593,N_34712);
or U35299 (N_35299,N_34969,N_34782);
xnor U35300 (N_35300,N_34605,N_34825);
xnor U35301 (N_35301,N_34952,N_34932);
nand U35302 (N_35302,N_34692,N_34554);
or U35303 (N_35303,N_34625,N_34656);
nand U35304 (N_35304,N_34929,N_34731);
nand U35305 (N_35305,N_34634,N_34752);
nand U35306 (N_35306,N_34570,N_34848);
nand U35307 (N_35307,N_34759,N_34955);
nand U35308 (N_35308,N_34764,N_34580);
and U35309 (N_35309,N_34711,N_34668);
or U35310 (N_35310,N_34592,N_34770);
nand U35311 (N_35311,N_34939,N_34766);
nand U35312 (N_35312,N_34566,N_34925);
xnor U35313 (N_35313,N_34658,N_34540);
nand U35314 (N_35314,N_34780,N_34679);
and U35315 (N_35315,N_34767,N_34662);
and U35316 (N_35316,N_34532,N_34891);
nor U35317 (N_35317,N_34595,N_34976);
nand U35318 (N_35318,N_34929,N_34988);
nor U35319 (N_35319,N_34583,N_34941);
or U35320 (N_35320,N_34857,N_34889);
and U35321 (N_35321,N_34530,N_34672);
and U35322 (N_35322,N_34899,N_34731);
and U35323 (N_35323,N_34510,N_34817);
or U35324 (N_35324,N_34554,N_34549);
nor U35325 (N_35325,N_34546,N_34765);
xor U35326 (N_35326,N_34598,N_34716);
or U35327 (N_35327,N_34588,N_34710);
nor U35328 (N_35328,N_34600,N_34933);
xor U35329 (N_35329,N_34664,N_34974);
nand U35330 (N_35330,N_34795,N_34578);
nor U35331 (N_35331,N_34654,N_34758);
and U35332 (N_35332,N_34806,N_34894);
xor U35333 (N_35333,N_34876,N_34750);
xnor U35334 (N_35334,N_34964,N_34911);
nor U35335 (N_35335,N_34624,N_34523);
xnor U35336 (N_35336,N_34771,N_34997);
nand U35337 (N_35337,N_34815,N_34742);
nor U35338 (N_35338,N_34620,N_34912);
and U35339 (N_35339,N_34960,N_34511);
nor U35340 (N_35340,N_34657,N_34571);
xnor U35341 (N_35341,N_34548,N_34848);
or U35342 (N_35342,N_34765,N_34930);
xnor U35343 (N_35343,N_34944,N_34795);
or U35344 (N_35344,N_34787,N_34826);
xnor U35345 (N_35345,N_34758,N_34989);
xnor U35346 (N_35346,N_34644,N_34803);
and U35347 (N_35347,N_34830,N_34787);
and U35348 (N_35348,N_34606,N_34693);
xnor U35349 (N_35349,N_34716,N_34932);
xnor U35350 (N_35350,N_34510,N_34665);
or U35351 (N_35351,N_34982,N_34728);
and U35352 (N_35352,N_34919,N_34693);
and U35353 (N_35353,N_34992,N_34855);
nand U35354 (N_35354,N_34926,N_34588);
or U35355 (N_35355,N_34852,N_34530);
or U35356 (N_35356,N_34707,N_34690);
xor U35357 (N_35357,N_34549,N_34846);
or U35358 (N_35358,N_34711,N_34542);
or U35359 (N_35359,N_34994,N_34976);
and U35360 (N_35360,N_34505,N_34577);
or U35361 (N_35361,N_34952,N_34833);
nand U35362 (N_35362,N_34747,N_34563);
or U35363 (N_35363,N_34653,N_34624);
or U35364 (N_35364,N_34772,N_34899);
or U35365 (N_35365,N_34814,N_34875);
xnor U35366 (N_35366,N_34743,N_34827);
or U35367 (N_35367,N_34845,N_34633);
nor U35368 (N_35368,N_34908,N_34836);
xor U35369 (N_35369,N_34583,N_34860);
nor U35370 (N_35370,N_34934,N_34721);
and U35371 (N_35371,N_34830,N_34863);
xor U35372 (N_35372,N_34786,N_34985);
nor U35373 (N_35373,N_34853,N_34970);
or U35374 (N_35374,N_34825,N_34902);
or U35375 (N_35375,N_34933,N_34712);
or U35376 (N_35376,N_34545,N_34804);
nand U35377 (N_35377,N_34949,N_34896);
nor U35378 (N_35378,N_34794,N_34919);
nor U35379 (N_35379,N_34678,N_34557);
or U35380 (N_35380,N_34964,N_34671);
and U35381 (N_35381,N_34899,N_34522);
nand U35382 (N_35382,N_34809,N_34629);
and U35383 (N_35383,N_34997,N_34747);
nor U35384 (N_35384,N_34594,N_34713);
and U35385 (N_35385,N_34951,N_34734);
or U35386 (N_35386,N_34983,N_34964);
nor U35387 (N_35387,N_34738,N_34769);
nor U35388 (N_35388,N_34904,N_34565);
nor U35389 (N_35389,N_34734,N_34827);
or U35390 (N_35390,N_34825,N_34928);
and U35391 (N_35391,N_34751,N_34817);
nand U35392 (N_35392,N_34827,N_34665);
and U35393 (N_35393,N_34930,N_34821);
nor U35394 (N_35394,N_34898,N_34705);
xor U35395 (N_35395,N_34746,N_34874);
xnor U35396 (N_35396,N_34932,N_34624);
or U35397 (N_35397,N_34713,N_34552);
nand U35398 (N_35398,N_34776,N_34954);
xor U35399 (N_35399,N_34789,N_34889);
nand U35400 (N_35400,N_34791,N_34835);
nand U35401 (N_35401,N_34986,N_34683);
and U35402 (N_35402,N_34519,N_34558);
nand U35403 (N_35403,N_34780,N_34814);
nor U35404 (N_35404,N_34876,N_34729);
nor U35405 (N_35405,N_34797,N_34686);
or U35406 (N_35406,N_34955,N_34549);
nand U35407 (N_35407,N_34685,N_34745);
and U35408 (N_35408,N_34664,N_34940);
xor U35409 (N_35409,N_34560,N_34916);
xor U35410 (N_35410,N_34875,N_34836);
and U35411 (N_35411,N_34756,N_34535);
xor U35412 (N_35412,N_34856,N_34978);
xor U35413 (N_35413,N_34735,N_34936);
and U35414 (N_35414,N_34743,N_34944);
nor U35415 (N_35415,N_34843,N_34666);
or U35416 (N_35416,N_34902,N_34857);
nor U35417 (N_35417,N_34959,N_34748);
or U35418 (N_35418,N_34576,N_34762);
or U35419 (N_35419,N_34911,N_34934);
xnor U35420 (N_35420,N_34702,N_34931);
and U35421 (N_35421,N_34993,N_34729);
and U35422 (N_35422,N_34517,N_34567);
nor U35423 (N_35423,N_34858,N_34853);
and U35424 (N_35424,N_34757,N_34654);
and U35425 (N_35425,N_34536,N_34647);
and U35426 (N_35426,N_34500,N_34931);
and U35427 (N_35427,N_34625,N_34970);
nor U35428 (N_35428,N_34883,N_34531);
or U35429 (N_35429,N_34658,N_34680);
and U35430 (N_35430,N_34691,N_34999);
or U35431 (N_35431,N_34901,N_34696);
or U35432 (N_35432,N_34896,N_34786);
or U35433 (N_35433,N_34890,N_34728);
and U35434 (N_35434,N_34779,N_34806);
xnor U35435 (N_35435,N_34931,N_34551);
xor U35436 (N_35436,N_34720,N_34613);
or U35437 (N_35437,N_34624,N_34717);
nor U35438 (N_35438,N_34867,N_34542);
nand U35439 (N_35439,N_34690,N_34960);
xnor U35440 (N_35440,N_34872,N_34578);
and U35441 (N_35441,N_34983,N_34948);
xnor U35442 (N_35442,N_34754,N_34950);
and U35443 (N_35443,N_34591,N_34722);
nor U35444 (N_35444,N_34511,N_34893);
or U35445 (N_35445,N_34759,N_34907);
nand U35446 (N_35446,N_34882,N_34521);
or U35447 (N_35447,N_34505,N_34746);
nor U35448 (N_35448,N_34669,N_34528);
xor U35449 (N_35449,N_34960,N_34567);
nand U35450 (N_35450,N_34543,N_34526);
and U35451 (N_35451,N_34950,N_34716);
xnor U35452 (N_35452,N_34617,N_34615);
nor U35453 (N_35453,N_34796,N_34919);
and U35454 (N_35454,N_34804,N_34984);
nand U35455 (N_35455,N_34748,N_34790);
or U35456 (N_35456,N_34892,N_34713);
nand U35457 (N_35457,N_34600,N_34713);
or U35458 (N_35458,N_34581,N_34838);
nor U35459 (N_35459,N_34915,N_34846);
and U35460 (N_35460,N_34951,N_34931);
nand U35461 (N_35461,N_34923,N_34778);
nor U35462 (N_35462,N_34932,N_34961);
xor U35463 (N_35463,N_34780,N_34760);
and U35464 (N_35464,N_34801,N_34524);
or U35465 (N_35465,N_34987,N_34795);
nand U35466 (N_35466,N_34935,N_34970);
nor U35467 (N_35467,N_34693,N_34569);
and U35468 (N_35468,N_34711,N_34864);
and U35469 (N_35469,N_34774,N_34642);
and U35470 (N_35470,N_34909,N_34920);
nand U35471 (N_35471,N_34697,N_34667);
and U35472 (N_35472,N_34724,N_34878);
or U35473 (N_35473,N_34769,N_34992);
or U35474 (N_35474,N_34728,N_34720);
nor U35475 (N_35475,N_34998,N_34622);
xnor U35476 (N_35476,N_34962,N_34848);
nor U35477 (N_35477,N_34987,N_34865);
nor U35478 (N_35478,N_34656,N_34949);
nor U35479 (N_35479,N_34844,N_34761);
and U35480 (N_35480,N_34619,N_34880);
nor U35481 (N_35481,N_34884,N_34601);
and U35482 (N_35482,N_34656,N_34757);
nand U35483 (N_35483,N_34866,N_34676);
xor U35484 (N_35484,N_34760,N_34874);
and U35485 (N_35485,N_34852,N_34582);
and U35486 (N_35486,N_34961,N_34621);
or U35487 (N_35487,N_34891,N_34918);
and U35488 (N_35488,N_34642,N_34932);
nand U35489 (N_35489,N_34974,N_34824);
nor U35490 (N_35490,N_34513,N_34899);
nor U35491 (N_35491,N_34558,N_34616);
or U35492 (N_35492,N_34658,N_34853);
nor U35493 (N_35493,N_34597,N_34557);
and U35494 (N_35494,N_34803,N_34985);
xnor U35495 (N_35495,N_34904,N_34533);
and U35496 (N_35496,N_34691,N_34889);
nor U35497 (N_35497,N_34519,N_34556);
nor U35498 (N_35498,N_34701,N_34580);
xor U35499 (N_35499,N_34791,N_34822);
and U35500 (N_35500,N_35273,N_35203);
or U35501 (N_35501,N_35092,N_35190);
nor U35502 (N_35502,N_35479,N_35116);
and U35503 (N_35503,N_35216,N_35037);
nand U35504 (N_35504,N_35356,N_35221);
or U35505 (N_35505,N_35486,N_35055);
or U35506 (N_35506,N_35097,N_35394);
nand U35507 (N_35507,N_35252,N_35162);
nand U35508 (N_35508,N_35075,N_35149);
nor U35509 (N_35509,N_35316,N_35173);
xor U35510 (N_35510,N_35269,N_35485);
nand U35511 (N_35511,N_35056,N_35388);
nand U35512 (N_35512,N_35193,N_35308);
xnor U35513 (N_35513,N_35219,N_35236);
and U35514 (N_35514,N_35089,N_35279);
and U35515 (N_35515,N_35440,N_35208);
xnor U35516 (N_35516,N_35405,N_35293);
or U35517 (N_35517,N_35110,N_35147);
nor U35518 (N_35518,N_35264,N_35315);
nor U35519 (N_35519,N_35191,N_35425);
nand U35520 (N_35520,N_35298,N_35033);
xnor U35521 (N_35521,N_35074,N_35164);
nor U35522 (N_35522,N_35230,N_35048);
xnor U35523 (N_35523,N_35400,N_35233);
xor U35524 (N_35524,N_35489,N_35412);
and U35525 (N_35525,N_35014,N_35061);
xnor U35526 (N_35526,N_35439,N_35199);
xor U35527 (N_35527,N_35312,N_35389);
nor U35528 (N_35528,N_35448,N_35072);
or U35529 (N_35529,N_35091,N_35163);
or U35530 (N_35530,N_35260,N_35031);
xnor U35531 (N_35531,N_35420,N_35287);
nand U35532 (N_35532,N_35437,N_35424);
nor U35533 (N_35533,N_35416,N_35004);
or U35534 (N_35534,N_35028,N_35160);
and U35535 (N_35535,N_35244,N_35043);
nor U35536 (N_35536,N_35169,N_35143);
or U35537 (N_35537,N_35330,N_35320);
nand U35538 (N_35538,N_35076,N_35141);
and U35539 (N_35539,N_35151,N_35059);
nor U35540 (N_35540,N_35111,N_35081);
and U35541 (N_35541,N_35429,N_35000);
and U35542 (N_35542,N_35123,N_35449);
nand U35543 (N_35543,N_35197,N_35011);
nor U35544 (N_35544,N_35372,N_35274);
and U35545 (N_35545,N_35460,N_35022);
nand U35546 (N_35546,N_35218,N_35484);
and U35547 (N_35547,N_35104,N_35189);
xnor U35548 (N_35548,N_35410,N_35369);
xnor U35549 (N_35549,N_35178,N_35069);
and U35550 (N_35550,N_35324,N_35174);
nor U35551 (N_35551,N_35352,N_35185);
or U35552 (N_35552,N_35120,N_35052);
or U35553 (N_35553,N_35248,N_35237);
and U35554 (N_35554,N_35499,N_35458);
and U35555 (N_35555,N_35426,N_35328);
or U35556 (N_35556,N_35130,N_35107);
and U35557 (N_35557,N_35140,N_35177);
or U35558 (N_35558,N_35327,N_35300);
and U35559 (N_35559,N_35378,N_35006);
nand U35560 (N_35560,N_35257,N_35342);
nand U35561 (N_35561,N_35399,N_35088);
xnor U35562 (N_35562,N_35438,N_35138);
nor U35563 (N_35563,N_35434,N_35026);
xnor U35564 (N_35564,N_35148,N_35036);
or U35565 (N_35565,N_35494,N_35166);
nand U35566 (N_35566,N_35431,N_35126);
or U35567 (N_35567,N_35231,N_35192);
nand U35568 (N_35568,N_35475,N_35361);
nand U35569 (N_35569,N_35467,N_35381);
or U35570 (N_35570,N_35102,N_35165);
xnor U35571 (N_35571,N_35270,N_35477);
nand U35572 (N_35572,N_35276,N_35351);
and U35573 (N_35573,N_35474,N_35461);
or U35574 (N_35574,N_35453,N_35187);
nor U35575 (N_35575,N_35417,N_35353);
or U35576 (N_35576,N_35357,N_35395);
nor U35577 (N_35577,N_35480,N_35409);
nand U35578 (N_35578,N_35047,N_35064);
nand U35579 (N_35579,N_35262,N_35058);
and U35580 (N_35580,N_35157,N_35398);
xor U35581 (N_35581,N_35242,N_35027);
or U35582 (N_35582,N_35343,N_35232);
xor U35583 (N_35583,N_35017,N_35432);
or U35584 (N_35584,N_35172,N_35331);
nand U35585 (N_35585,N_35284,N_35376);
or U35586 (N_35586,N_35195,N_35122);
xor U35587 (N_35587,N_35358,N_35243);
nand U35588 (N_35588,N_35314,N_35085);
nor U35589 (N_35589,N_35430,N_35333);
xnor U35590 (N_35590,N_35039,N_35186);
nor U35591 (N_35591,N_35057,N_35129);
or U35592 (N_35592,N_35355,N_35490);
nand U35593 (N_35593,N_35281,N_35124);
xor U35594 (N_35594,N_35283,N_35206);
nor U35595 (N_35595,N_35167,N_35465);
or U35596 (N_35596,N_35096,N_35457);
or U35597 (N_35597,N_35068,N_35344);
and U35598 (N_35598,N_35121,N_35239);
or U35599 (N_35599,N_35240,N_35435);
and U35600 (N_35600,N_35042,N_35201);
and U35601 (N_35601,N_35019,N_35263);
or U35602 (N_35602,N_35049,N_35154);
and U35603 (N_35603,N_35084,N_35025);
nand U35604 (N_35604,N_35265,N_35476);
nand U35605 (N_35605,N_35387,N_35347);
nand U35606 (N_35606,N_35211,N_35001);
nand U35607 (N_35607,N_35456,N_35238);
nor U35608 (N_35608,N_35098,N_35051);
or U35609 (N_35609,N_35183,N_35322);
xnor U35610 (N_35610,N_35109,N_35452);
nand U35611 (N_35611,N_35127,N_35223);
nor U35612 (N_35612,N_35371,N_35018);
nor U35613 (N_35613,N_35488,N_35340);
xor U35614 (N_35614,N_35272,N_35336);
and U35615 (N_35615,N_35146,N_35278);
nor U35616 (N_35616,N_35099,N_35079);
nand U35617 (N_35617,N_35291,N_35217);
nand U35618 (N_35618,N_35466,N_35132);
xor U35619 (N_35619,N_35370,N_35133);
nand U35620 (N_35620,N_35338,N_35065);
nor U35621 (N_35621,N_35294,N_35491);
nand U35622 (N_35622,N_35415,N_35101);
xnor U35623 (N_35623,N_35297,N_35487);
or U35624 (N_35624,N_35153,N_35087);
or U35625 (N_35625,N_35118,N_35222);
nand U35626 (N_35626,N_35117,N_35176);
nor U35627 (N_35627,N_35450,N_35411);
or U35628 (N_35628,N_35402,N_35207);
xor U35629 (N_35629,N_35082,N_35241);
or U35630 (N_35630,N_35214,N_35170);
or U35631 (N_35631,N_35181,N_35478);
nand U35632 (N_35632,N_35250,N_35053);
and U35633 (N_35633,N_35015,N_35423);
and U35634 (N_35634,N_35295,N_35392);
nor U35635 (N_35635,N_35229,N_35433);
or U35636 (N_35636,N_35288,N_35073);
and U35637 (N_35637,N_35005,N_35050);
nor U35638 (N_35638,N_35246,N_35045);
and U35639 (N_35639,N_35009,N_35419);
nor U35640 (N_35640,N_35063,N_35100);
and U35641 (N_35641,N_35078,N_35215);
nand U35642 (N_35642,N_35180,N_35443);
xor U35643 (N_35643,N_35204,N_35158);
xnor U35644 (N_35644,N_35114,N_35010);
xor U35645 (N_35645,N_35285,N_35271);
nor U35646 (N_35646,N_35012,N_35194);
nor U35647 (N_35647,N_35105,N_35459);
and U35648 (N_35648,N_35003,N_35367);
or U35649 (N_35649,N_35106,N_35418);
nor U35650 (N_35650,N_35414,N_35290);
nor U35651 (N_35651,N_35307,N_35345);
and U35652 (N_35652,N_35359,N_35496);
xnor U35653 (N_35653,N_35255,N_35428);
and U35654 (N_35654,N_35311,N_35188);
nor U35655 (N_35655,N_35258,N_35482);
or U35656 (N_35656,N_35379,N_35319);
or U35657 (N_35657,N_35228,N_35032);
nor U35658 (N_35658,N_35225,N_35016);
nor U35659 (N_35659,N_35296,N_35386);
or U35660 (N_35660,N_35303,N_35339);
and U35661 (N_35661,N_35247,N_35403);
or U35662 (N_35662,N_35182,N_35391);
xnor U35663 (N_35663,N_35041,N_35483);
nand U35664 (N_35664,N_35454,N_35377);
xor U35665 (N_35665,N_35023,N_35095);
xnor U35666 (N_35666,N_35071,N_35442);
nand U35667 (N_35667,N_35396,N_35383);
nand U35668 (N_35668,N_35304,N_35226);
nand U35669 (N_35669,N_35196,N_35366);
and U35670 (N_35670,N_35472,N_35282);
and U35671 (N_35671,N_35444,N_35224);
and U35672 (N_35672,N_35234,N_35145);
nor U35673 (N_35673,N_35030,N_35038);
xnor U35674 (N_35674,N_35268,N_35408);
nand U35675 (N_35675,N_35374,N_35093);
nand U35676 (N_35676,N_35323,N_35363);
nand U35677 (N_35677,N_35393,N_35495);
nand U35678 (N_35678,N_35302,N_35112);
nand U35679 (N_35679,N_35156,N_35380);
nor U35680 (N_35680,N_35368,N_35317);
or U35681 (N_35681,N_35326,N_35086);
or U35682 (N_35682,N_35335,N_35407);
nor U35683 (N_35683,N_35447,N_35346);
nand U35684 (N_35684,N_35128,N_35002);
nor U35685 (N_35685,N_35373,N_35292);
and U35686 (N_35686,N_35404,N_35094);
nor U35687 (N_35687,N_35493,N_35364);
xor U35688 (N_35688,N_35134,N_35200);
nand U35689 (N_35689,N_35375,N_35034);
or U35690 (N_35690,N_35139,N_35220);
xor U35691 (N_35691,N_35313,N_35066);
xor U35692 (N_35692,N_35286,N_35152);
nand U35693 (N_35693,N_35062,N_35348);
xor U35694 (N_35694,N_35007,N_35468);
and U35695 (N_35695,N_35035,N_35350);
or U35696 (N_35696,N_35060,N_35390);
and U35697 (N_35697,N_35159,N_35103);
nand U35698 (N_35698,N_35384,N_35280);
nand U35699 (N_35699,N_35227,N_35266);
xnor U35700 (N_35700,N_35397,N_35362);
nand U35701 (N_35701,N_35360,N_35135);
nand U35702 (N_35702,N_35321,N_35329);
nand U35703 (N_35703,N_35337,N_35275);
or U35704 (N_35704,N_35277,N_35245);
or U35705 (N_35705,N_35013,N_35113);
nor U35706 (N_35706,N_35446,N_35213);
and U35707 (N_35707,N_35310,N_35175);
or U35708 (N_35708,N_35305,N_35259);
nand U35709 (N_35709,N_35445,N_35040);
nand U35710 (N_35710,N_35168,N_35498);
nand U35711 (N_35711,N_35401,N_35161);
xor U35712 (N_35712,N_35289,N_35070);
or U35713 (N_35713,N_35497,N_35341);
nor U35714 (N_35714,N_35254,N_35334);
nand U35715 (N_35715,N_35249,N_35253);
xnor U35716 (N_35716,N_35077,N_35090);
nor U35717 (N_35717,N_35481,N_35365);
and U35718 (N_35718,N_35131,N_35171);
or U35719 (N_35719,N_35080,N_35212);
nor U35720 (N_35720,N_35256,N_35413);
nor U35721 (N_35721,N_35422,N_35202);
and U35722 (N_35722,N_35309,N_35455);
nor U35723 (N_35723,N_35210,N_35382);
xnor U35724 (N_35724,N_35024,N_35020);
xor U35725 (N_35725,N_35299,N_35492);
or U35726 (N_35726,N_35125,N_35469);
nor U35727 (N_35727,N_35470,N_35306);
xor U35728 (N_35728,N_35451,N_35205);
and U35729 (N_35729,N_35108,N_35441);
xnor U35730 (N_35730,N_35251,N_35332);
nand U35731 (N_35731,N_35115,N_35144);
and U35732 (N_35732,N_35473,N_35044);
and U35733 (N_35733,N_35119,N_35008);
xnor U35734 (N_35734,N_35354,N_35235);
nor U35735 (N_35735,N_35046,N_35318);
xor U35736 (N_35736,N_35179,N_35427);
or U35737 (N_35737,N_35325,N_35137);
and U35738 (N_35738,N_35463,N_35136);
nand U35739 (N_35739,N_35261,N_35067);
xnor U35740 (N_35740,N_35385,N_35054);
or U35741 (N_35741,N_35301,N_35198);
and U35742 (N_35742,N_35142,N_35267);
xor U35743 (N_35743,N_35462,N_35021);
nor U35744 (N_35744,N_35155,N_35436);
nor U35745 (N_35745,N_35150,N_35421);
nand U35746 (N_35746,N_35471,N_35029);
xor U35747 (N_35747,N_35349,N_35464);
xnor U35748 (N_35748,N_35406,N_35209);
or U35749 (N_35749,N_35083,N_35184);
xor U35750 (N_35750,N_35251,N_35016);
xor U35751 (N_35751,N_35491,N_35009);
nor U35752 (N_35752,N_35410,N_35012);
nor U35753 (N_35753,N_35460,N_35279);
nand U35754 (N_35754,N_35169,N_35159);
xnor U35755 (N_35755,N_35349,N_35436);
or U35756 (N_35756,N_35378,N_35440);
nand U35757 (N_35757,N_35158,N_35051);
xor U35758 (N_35758,N_35382,N_35053);
nand U35759 (N_35759,N_35174,N_35246);
and U35760 (N_35760,N_35100,N_35447);
nand U35761 (N_35761,N_35251,N_35284);
and U35762 (N_35762,N_35102,N_35114);
nand U35763 (N_35763,N_35023,N_35166);
nor U35764 (N_35764,N_35166,N_35430);
nand U35765 (N_35765,N_35331,N_35372);
xnor U35766 (N_35766,N_35093,N_35444);
and U35767 (N_35767,N_35101,N_35198);
or U35768 (N_35768,N_35415,N_35167);
nand U35769 (N_35769,N_35492,N_35387);
xnor U35770 (N_35770,N_35221,N_35171);
nand U35771 (N_35771,N_35054,N_35055);
or U35772 (N_35772,N_35422,N_35250);
or U35773 (N_35773,N_35125,N_35259);
nand U35774 (N_35774,N_35341,N_35403);
xnor U35775 (N_35775,N_35368,N_35066);
nor U35776 (N_35776,N_35428,N_35330);
and U35777 (N_35777,N_35085,N_35049);
nor U35778 (N_35778,N_35260,N_35305);
nor U35779 (N_35779,N_35133,N_35040);
xnor U35780 (N_35780,N_35215,N_35104);
and U35781 (N_35781,N_35449,N_35290);
or U35782 (N_35782,N_35367,N_35443);
xnor U35783 (N_35783,N_35052,N_35262);
nor U35784 (N_35784,N_35196,N_35401);
xnor U35785 (N_35785,N_35020,N_35293);
nor U35786 (N_35786,N_35260,N_35258);
and U35787 (N_35787,N_35157,N_35112);
xor U35788 (N_35788,N_35337,N_35214);
nor U35789 (N_35789,N_35016,N_35363);
nor U35790 (N_35790,N_35162,N_35135);
nand U35791 (N_35791,N_35415,N_35343);
and U35792 (N_35792,N_35403,N_35286);
xnor U35793 (N_35793,N_35246,N_35063);
xnor U35794 (N_35794,N_35260,N_35158);
nor U35795 (N_35795,N_35160,N_35168);
xor U35796 (N_35796,N_35269,N_35055);
and U35797 (N_35797,N_35158,N_35041);
and U35798 (N_35798,N_35342,N_35355);
or U35799 (N_35799,N_35479,N_35038);
nand U35800 (N_35800,N_35462,N_35008);
nor U35801 (N_35801,N_35328,N_35141);
nand U35802 (N_35802,N_35282,N_35465);
nand U35803 (N_35803,N_35385,N_35059);
and U35804 (N_35804,N_35437,N_35029);
xnor U35805 (N_35805,N_35434,N_35264);
nor U35806 (N_35806,N_35335,N_35408);
xnor U35807 (N_35807,N_35252,N_35076);
nor U35808 (N_35808,N_35035,N_35435);
nor U35809 (N_35809,N_35396,N_35266);
and U35810 (N_35810,N_35261,N_35006);
xnor U35811 (N_35811,N_35257,N_35405);
xor U35812 (N_35812,N_35079,N_35152);
nand U35813 (N_35813,N_35368,N_35043);
and U35814 (N_35814,N_35310,N_35359);
and U35815 (N_35815,N_35114,N_35016);
nor U35816 (N_35816,N_35203,N_35312);
or U35817 (N_35817,N_35430,N_35361);
nand U35818 (N_35818,N_35080,N_35071);
xor U35819 (N_35819,N_35062,N_35363);
nor U35820 (N_35820,N_35331,N_35345);
xnor U35821 (N_35821,N_35319,N_35059);
and U35822 (N_35822,N_35111,N_35098);
nand U35823 (N_35823,N_35176,N_35410);
or U35824 (N_35824,N_35073,N_35065);
nand U35825 (N_35825,N_35205,N_35115);
and U35826 (N_35826,N_35351,N_35277);
and U35827 (N_35827,N_35378,N_35323);
nand U35828 (N_35828,N_35009,N_35119);
or U35829 (N_35829,N_35497,N_35470);
nand U35830 (N_35830,N_35240,N_35186);
nor U35831 (N_35831,N_35072,N_35414);
and U35832 (N_35832,N_35229,N_35449);
nand U35833 (N_35833,N_35368,N_35288);
nand U35834 (N_35834,N_35169,N_35174);
or U35835 (N_35835,N_35423,N_35451);
and U35836 (N_35836,N_35252,N_35325);
nor U35837 (N_35837,N_35413,N_35452);
xnor U35838 (N_35838,N_35360,N_35021);
or U35839 (N_35839,N_35311,N_35242);
or U35840 (N_35840,N_35415,N_35158);
nor U35841 (N_35841,N_35121,N_35043);
or U35842 (N_35842,N_35323,N_35253);
nand U35843 (N_35843,N_35211,N_35468);
nor U35844 (N_35844,N_35132,N_35089);
nor U35845 (N_35845,N_35264,N_35389);
and U35846 (N_35846,N_35401,N_35262);
nand U35847 (N_35847,N_35418,N_35055);
or U35848 (N_35848,N_35229,N_35097);
nor U35849 (N_35849,N_35333,N_35245);
or U35850 (N_35850,N_35252,N_35053);
nand U35851 (N_35851,N_35479,N_35177);
nor U35852 (N_35852,N_35188,N_35485);
nor U35853 (N_35853,N_35325,N_35277);
xor U35854 (N_35854,N_35444,N_35322);
and U35855 (N_35855,N_35107,N_35177);
or U35856 (N_35856,N_35190,N_35138);
or U35857 (N_35857,N_35154,N_35423);
nor U35858 (N_35858,N_35196,N_35425);
or U35859 (N_35859,N_35310,N_35299);
and U35860 (N_35860,N_35423,N_35107);
xor U35861 (N_35861,N_35040,N_35044);
and U35862 (N_35862,N_35322,N_35101);
nor U35863 (N_35863,N_35384,N_35244);
nand U35864 (N_35864,N_35215,N_35255);
and U35865 (N_35865,N_35362,N_35185);
nand U35866 (N_35866,N_35445,N_35411);
or U35867 (N_35867,N_35044,N_35169);
nor U35868 (N_35868,N_35307,N_35092);
nand U35869 (N_35869,N_35402,N_35233);
nand U35870 (N_35870,N_35065,N_35441);
nand U35871 (N_35871,N_35137,N_35103);
and U35872 (N_35872,N_35399,N_35036);
and U35873 (N_35873,N_35331,N_35189);
xor U35874 (N_35874,N_35102,N_35178);
or U35875 (N_35875,N_35498,N_35350);
or U35876 (N_35876,N_35228,N_35365);
nand U35877 (N_35877,N_35192,N_35122);
or U35878 (N_35878,N_35481,N_35009);
xnor U35879 (N_35879,N_35400,N_35154);
nor U35880 (N_35880,N_35342,N_35102);
or U35881 (N_35881,N_35030,N_35260);
nand U35882 (N_35882,N_35271,N_35008);
nor U35883 (N_35883,N_35128,N_35433);
xnor U35884 (N_35884,N_35075,N_35058);
xnor U35885 (N_35885,N_35288,N_35045);
or U35886 (N_35886,N_35276,N_35256);
or U35887 (N_35887,N_35013,N_35197);
xor U35888 (N_35888,N_35201,N_35398);
xnor U35889 (N_35889,N_35178,N_35262);
nor U35890 (N_35890,N_35354,N_35390);
nand U35891 (N_35891,N_35146,N_35373);
and U35892 (N_35892,N_35211,N_35168);
nor U35893 (N_35893,N_35480,N_35037);
and U35894 (N_35894,N_35172,N_35486);
xnor U35895 (N_35895,N_35284,N_35426);
or U35896 (N_35896,N_35401,N_35475);
and U35897 (N_35897,N_35174,N_35186);
and U35898 (N_35898,N_35402,N_35065);
xnor U35899 (N_35899,N_35454,N_35170);
or U35900 (N_35900,N_35001,N_35217);
nor U35901 (N_35901,N_35405,N_35253);
and U35902 (N_35902,N_35092,N_35397);
and U35903 (N_35903,N_35042,N_35112);
and U35904 (N_35904,N_35221,N_35086);
or U35905 (N_35905,N_35010,N_35070);
nand U35906 (N_35906,N_35030,N_35239);
xnor U35907 (N_35907,N_35206,N_35067);
xnor U35908 (N_35908,N_35402,N_35312);
and U35909 (N_35909,N_35307,N_35112);
or U35910 (N_35910,N_35109,N_35481);
or U35911 (N_35911,N_35210,N_35325);
nor U35912 (N_35912,N_35146,N_35132);
and U35913 (N_35913,N_35032,N_35060);
xnor U35914 (N_35914,N_35364,N_35430);
or U35915 (N_35915,N_35168,N_35053);
and U35916 (N_35916,N_35093,N_35474);
xnor U35917 (N_35917,N_35390,N_35157);
nor U35918 (N_35918,N_35441,N_35164);
nor U35919 (N_35919,N_35319,N_35174);
nand U35920 (N_35920,N_35455,N_35327);
nor U35921 (N_35921,N_35293,N_35206);
or U35922 (N_35922,N_35493,N_35286);
xnor U35923 (N_35923,N_35079,N_35159);
xor U35924 (N_35924,N_35372,N_35307);
xnor U35925 (N_35925,N_35079,N_35455);
xor U35926 (N_35926,N_35416,N_35380);
and U35927 (N_35927,N_35181,N_35235);
xor U35928 (N_35928,N_35101,N_35039);
and U35929 (N_35929,N_35467,N_35453);
nor U35930 (N_35930,N_35454,N_35171);
or U35931 (N_35931,N_35336,N_35218);
and U35932 (N_35932,N_35481,N_35071);
xor U35933 (N_35933,N_35077,N_35438);
or U35934 (N_35934,N_35341,N_35195);
or U35935 (N_35935,N_35100,N_35142);
nand U35936 (N_35936,N_35354,N_35136);
nor U35937 (N_35937,N_35221,N_35359);
or U35938 (N_35938,N_35084,N_35382);
xor U35939 (N_35939,N_35424,N_35314);
nor U35940 (N_35940,N_35102,N_35164);
nand U35941 (N_35941,N_35340,N_35178);
xnor U35942 (N_35942,N_35337,N_35131);
or U35943 (N_35943,N_35023,N_35439);
xor U35944 (N_35944,N_35006,N_35354);
and U35945 (N_35945,N_35427,N_35168);
nor U35946 (N_35946,N_35334,N_35405);
and U35947 (N_35947,N_35212,N_35323);
nand U35948 (N_35948,N_35249,N_35178);
and U35949 (N_35949,N_35308,N_35126);
and U35950 (N_35950,N_35079,N_35420);
nor U35951 (N_35951,N_35022,N_35088);
xnor U35952 (N_35952,N_35175,N_35231);
and U35953 (N_35953,N_35011,N_35023);
xnor U35954 (N_35954,N_35167,N_35252);
and U35955 (N_35955,N_35041,N_35104);
xor U35956 (N_35956,N_35385,N_35370);
and U35957 (N_35957,N_35439,N_35190);
xor U35958 (N_35958,N_35259,N_35192);
nand U35959 (N_35959,N_35404,N_35076);
or U35960 (N_35960,N_35067,N_35330);
or U35961 (N_35961,N_35457,N_35040);
nor U35962 (N_35962,N_35463,N_35043);
nand U35963 (N_35963,N_35042,N_35221);
nand U35964 (N_35964,N_35086,N_35214);
xor U35965 (N_35965,N_35317,N_35008);
nand U35966 (N_35966,N_35044,N_35020);
and U35967 (N_35967,N_35499,N_35429);
nand U35968 (N_35968,N_35171,N_35175);
nand U35969 (N_35969,N_35198,N_35376);
nor U35970 (N_35970,N_35375,N_35326);
nand U35971 (N_35971,N_35339,N_35342);
and U35972 (N_35972,N_35030,N_35141);
xor U35973 (N_35973,N_35070,N_35003);
and U35974 (N_35974,N_35301,N_35020);
and U35975 (N_35975,N_35408,N_35273);
and U35976 (N_35976,N_35447,N_35399);
nand U35977 (N_35977,N_35450,N_35492);
or U35978 (N_35978,N_35441,N_35374);
or U35979 (N_35979,N_35358,N_35407);
nand U35980 (N_35980,N_35180,N_35142);
and U35981 (N_35981,N_35158,N_35271);
xor U35982 (N_35982,N_35288,N_35379);
xor U35983 (N_35983,N_35366,N_35156);
or U35984 (N_35984,N_35371,N_35490);
nor U35985 (N_35985,N_35415,N_35173);
nor U35986 (N_35986,N_35420,N_35110);
nand U35987 (N_35987,N_35464,N_35147);
nand U35988 (N_35988,N_35035,N_35289);
and U35989 (N_35989,N_35494,N_35192);
nor U35990 (N_35990,N_35067,N_35402);
and U35991 (N_35991,N_35259,N_35484);
and U35992 (N_35992,N_35284,N_35179);
nor U35993 (N_35993,N_35426,N_35053);
or U35994 (N_35994,N_35309,N_35448);
xor U35995 (N_35995,N_35055,N_35384);
or U35996 (N_35996,N_35329,N_35360);
or U35997 (N_35997,N_35487,N_35289);
and U35998 (N_35998,N_35203,N_35476);
or U35999 (N_35999,N_35300,N_35146);
nand U36000 (N_36000,N_35571,N_35635);
nand U36001 (N_36001,N_35588,N_35940);
xor U36002 (N_36002,N_35766,N_35846);
and U36003 (N_36003,N_35779,N_35673);
nand U36004 (N_36004,N_35778,N_35761);
and U36005 (N_36005,N_35870,N_35557);
xnor U36006 (N_36006,N_35532,N_35710);
and U36007 (N_36007,N_35686,N_35567);
nor U36008 (N_36008,N_35861,N_35606);
nor U36009 (N_36009,N_35732,N_35843);
nor U36010 (N_36010,N_35845,N_35962);
xor U36011 (N_36011,N_35565,N_35738);
and U36012 (N_36012,N_35748,N_35944);
or U36013 (N_36013,N_35929,N_35867);
nand U36014 (N_36014,N_35596,N_35862);
xnor U36015 (N_36015,N_35988,N_35733);
nand U36016 (N_36016,N_35508,N_35511);
xor U36017 (N_36017,N_35628,N_35807);
xnor U36018 (N_36018,N_35801,N_35726);
nor U36019 (N_36019,N_35774,N_35966);
xnor U36020 (N_36020,N_35989,N_35872);
xor U36021 (N_36021,N_35637,N_35668);
or U36022 (N_36022,N_35873,N_35608);
xnor U36023 (N_36023,N_35936,N_35816);
nand U36024 (N_36024,N_35636,N_35947);
or U36025 (N_36025,N_35651,N_35687);
or U36026 (N_36026,N_35852,N_35893);
nand U36027 (N_36027,N_35556,N_35706);
or U36028 (N_36028,N_35715,N_35850);
xor U36029 (N_36029,N_35725,N_35786);
xnor U36030 (N_36030,N_35755,N_35613);
and U36031 (N_36031,N_35994,N_35611);
nor U36032 (N_36032,N_35593,N_35971);
nor U36033 (N_36033,N_35711,N_35827);
or U36034 (N_36034,N_35623,N_35860);
xnor U36035 (N_36035,N_35681,N_35926);
nor U36036 (N_36036,N_35770,N_35782);
and U36037 (N_36037,N_35930,N_35570);
and U36038 (N_36038,N_35544,N_35894);
nor U36039 (N_36039,N_35856,N_35704);
nand U36040 (N_36040,N_35505,N_35527);
or U36041 (N_36041,N_35718,N_35773);
xnor U36042 (N_36042,N_35908,N_35808);
or U36043 (N_36043,N_35569,N_35612);
nor U36044 (N_36044,N_35875,N_35888);
xor U36045 (N_36045,N_35982,N_35553);
or U36046 (N_36046,N_35920,N_35996);
nor U36047 (N_36047,N_35721,N_35512);
nor U36048 (N_36048,N_35661,N_35837);
nor U36049 (N_36049,N_35787,N_35534);
and U36050 (N_36050,N_35806,N_35741);
nor U36051 (N_36051,N_35735,N_35560);
nor U36052 (N_36052,N_35682,N_35825);
nor U36053 (N_36053,N_35848,N_35584);
xor U36054 (N_36054,N_35632,N_35641);
and U36055 (N_36055,N_35907,N_35969);
or U36056 (N_36056,N_35616,N_35678);
xnor U36057 (N_36057,N_35690,N_35656);
nor U36058 (N_36058,N_35603,N_35914);
xnor U36059 (N_36059,N_35762,N_35542);
nor U36060 (N_36060,N_35500,N_35780);
xnor U36061 (N_36061,N_35714,N_35645);
and U36062 (N_36062,N_35529,N_35700);
xnor U36063 (N_36063,N_35876,N_35805);
nand U36064 (N_36064,N_35540,N_35615);
nor U36065 (N_36065,N_35535,N_35979);
or U36066 (N_36066,N_35784,N_35702);
xor U36067 (N_36067,N_35980,N_35643);
xor U36068 (N_36068,N_35601,N_35857);
xnor U36069 (N_36069,N_35509,N_35520);
xor U36070 (N_36070,N_35829,N_35948);
and U36071 (N_36071,N_35555,N_35659);
nor U36072 (N_36072,N_35579,N_35865);
or U36073 (N_36073,N_35776,N_35528);
nand U36074 (N_36074,N_35953,N_35858);
nand U36075 (N_36075,N_35869,N_35941);
xor U36076 (N_36076,N_35781,N_35792);
nor U36077 (N_36077,N_35968,N_35760);
and U36078 (N_36078,N_35881,N_35594);
or U36079 (N_36079,N_35853,N_35692);
xnor U36080 (N_36080,N_35727,N_35946);
or U36081 (N_36081,N_35618,N_35712);
nor U36082 (N_36082,N_35677,N_35642);
nor U36083 (N_36083,N_35964,N_35812);
nand U36084 (N_36084,N_35660,N_35817);
nand U36085 (N_36085,N_35600,N_35831);
nor U36086 (N_36086,N_35810,N_35866);
xor U36087 (N_36087,N_35559,N_35595);
or U36088 (N_36088,N_35647,N_35871);
and U36089 (N_36089,N_35765,N_35890);
or U36090 (N_36090,N_35768,N_35609);
nand U36091 (N_36091,N_35878,N_35975);
nand U36092 (N_36092,N_35756,N_35895);
xor U36093 (N_36093,N_35684,N_35874);
or U36094 (N_36094,N_35717,N_35984);
or U36095 (N_36095,N_35833,N_35960);
or U36096 (N_36096,N_35959,N_35583);
xnor U36097 (N_36097,N_35917,N_35802);
xor U36098 (N_36098,N_35614,N_35832);
and U36099 (N_36099,N_35699,N_35904);
or U36100 (N_36100,N_35620,N_35519);
and U36101 (N_36101,N_35949,N_35950);
or U36102 (N_36102,N_35501,N_35737);
nor U36103 (N_36103,N_35887,N_35899);
nor U36104 (N_36104,N_35551,N_35646);
and U36105 (N_36105,N_35526,N_35772);
or U36106 (N_36106,N_35548,N_35558);
or U36107 (N_36107,N_35921,N_35924);
xor U36108 (N_36108,N_35785,N_35723);
nor U36109 (N_36109,N_35859,N_35739);
nand U36110 (N_36110,N_35824,N_35574);
nand U36111 (N_36111,N_35951,N_35954);
and U36112 (N_36112,N_35543,N_35884);
xor U36113 (N_36113,N_35961,N_35992);
and U36114 (N_36114,N_35967,N_35589);
xor U36115 (N_36115,N_35758,N_35877);
nor U36116 (N_36116,N_35918,N_35999);
nand U36117 (N_36117,N_35592,N_35937);
xor U36118 (N_36118,N_35942,N_35648);
xor U36119 (N_36119,N_35639,N_35803);
xnor U36120 (N_36120,N_35838,N_35743);
and U36121 (N_36121,N_35729,N_35581);
or U36122 (N_36122,N_35518,N_35549);
nand U36123 (N_36123,N_35649,N_35742);
nor U36124 (N_36124,N_35891,N_35575);
nor U36125 (N_36125,N_35834,N_35965);
and U36126 (N_36126,N_35905,N_35719);
nor U36127 (N_36127,N_35703,N_35531);
or U36128 (N_36128,N_35537,N_35550);
xnor U36129 (N_36129,N_35597,N_35516);
and U36130 (N_36130,N_35883,N_35854);
and U36131 (N_36131,N_35836,N_35906);
nor U36132 (N_36132,N_35713,N_35578);
or U36133 (N_36133,N_35669,N_35911);
xor U36134 (N_36134,N_35745,N_35902);
nor U36135 (N_36135,N_35602,N_35728);
xor U36136 (N_36136,N_35676,N_35759);
nand U36137 (N_36137,N_35985,N_35754);
nand U36138 (N_36138,N_35675,N_35724);
xor U36139 (N_36139,N_35910,N_35683);
and U36140 (N_36140,N_35913,N_35811);
and U36141 (N_36141,N_35956,N_35610);
nor U36142 (N_36142,N_35633,N_35629);
or U36143 (N_36143,N_35586,N_35698);
or U36144 (N_36144,N_35795,N_35685);
nor U36145 (N_36145,N_35749,N_35932);
and U36146 (N_36146,N_35538,N_35638);
or U36147 (N_36147,N_35835,N_35502);
or U36148 (N_36148,N_35680,N_35804);
or U36149 (N_36149,N_35892,N_35868);
and U36150 (N_36150,N_35619,N_35736);
nor U36151 (N_36151,N_35809,N_35655);
nand U36152 (N_36152,N_35644,N_35771);
nand U36153 (N_36153,N_35521,N_35672);
xor U36154 (N_36154,N_35506,N_35981);
nand U36155 (N_36155,N_35563,N_35747);
xor U36156 (N_36156,N_35577,N_35547);
and U36157 (N_36157,N_35983,N_35731);
nor U36158 (N_36158,N_35842,N_35819);
nor U36159 (N_36159,N_35815,N_35800);
or U36160 (N_36160,N_35744,N_35963);
or U36161 (N_36161,N_35821,N_35525);
xor U36162 (N_36162,N_35775,N_35752);
or U36163 (N_36163,N_35734,N_35909);
nand U36164 (N_36164,N_35794,N_35793);
or U36165 (N_36165,N_35552,N_35840);
or U36166 (N_36166,N_35561,N_35564);
nor U36167 (N_36167,N_35694,N_35697);
nand U36168 (N_36168,N_35546,N_35514);
and U36169 (N_36169,N_35777,N_35566);
nor U36170 (N_36170,N_35572,N_35716);
xnor U36171 (N_36171,N_35879,N_35851);
nand U36172 (N_36172,N_35707,N_35934);
or U36173 (N_36173,N_35849,N_35653);
nor U36174 (N_36174,N_35626,N_35976);
nand U36175 (N_36175,N_35693,N_35652);
nand U36176 (N_36176,N_35513,N_35695);
and U36177 (N_36177,N_35688,N_35701);
or U36178 (N_36178,N_35978,N_35864);
nand U36179 (N_36179,N_35767,N_35974);
or U36180 (N_36180,N_35523,N_35799);
nor U36181 (N_36181,N_35783,N_35995);
nor U36182 (N_36182,N_35885,N_35919);
and U36183 (N_36183,N_35973,N_35889);
nor U36184 (N_36184,N_35708,N_35705);
xnor U36185 (N_36185,N_35986,N_35662);
or U36186 (N_36186,N_35517,N_35666);
xnor U36187 (N_36187,N_35503,N_35998);
nand U36188 (N_36188,N_35928,N_35952);
and U36189 (N_36189,N_35958,N_35922);
or U36190 (N_36190,N_35598,N_35582);
nand U36191 (N_36191,N_35539,N_35554);
nand U36192 (N_36192,N_35625,N_35791);
nor U36193 (N_36193,N_35631,N_35763);
xnor U36194 (N_36194,N_35515,N_35826);
xnor U36195 (N_36195,N_35664,N_35790);
and U36196 (N_36196,N_35587,N_35797);
or U36197 (N_36197,N_35654,N_35663);
or U36198 (N_36198,N_35650,N_35820);
xor U36199 (N_36199,N_35634,N_35788);
nor U36200 (N_36200,N_35830,N_35576);
xor U36201 (N_36201,N_35585,N_35510);
xor U36202 (N_36202,N_35839,N_35847);
or U36203 (N_36203,N_35507,N_35696);
xor U36204 (N_36204,N_35796,N_35536);
and U36205 (N_36205,N_35822,N_35750);
or U36206 (N_36206,N_35931,N_35987);
nand U36207 (N_36207,N_35580,N_35912);
nand U36208 (N_36208,N_35740,N_35939);
and U36209 (N_36209,N_35764,N_35657);
and U36210 (N_36210,N_35671,N_35997);
and U36211 (N_36211,N_35568,N_35753);
nand U36212 (N_36212,N_35990,N_35993);
or U36213 (N_36213,N_35915,N_35769);
nor U36214 (N_36214,N_35916,N_35901);
xor U36215 (N_36215,N_35925,N_35627);
and U36216 (N_36216,N_35897,N_35903);
or U36217 (N_36217,N_35622,N_35670);
or U36218 (N_36218,N_35945,N_35972);
xor U36219 (N_36219,N_35841,N_35722);
or U36220 (N_36220,N_35640,N_35541);
nand U36221 (N_36221,N_35957,N_35573);
nor U36222 (N_36222,N_35658,N_35863);
xor U36223 (N_36223,N_35927,N_35530);
or U36224 (N_36224,N_35533,N_35746);
nor U36225 (N_36225,N_35624,N_35522);
and U36226 (N_36226,N_35818,N_35933);
nor U36227 (N_36227,N_35813,N_35674);
and U36228 (N_36228,N_35970,N_35504);
xnor U36229 (N_36229,N_35630,N_35617);
nor U36230 (N_36230,N_35900,N_35751);
or U36231 (N_36231,N_35798,N_35935);
nor U36232 (N_36232,N_35689,N_35823);
nand U36233 (N_36233,N_35923,N_35709);
and U36234 (N_36234,N_35855,N_35562);
or U36235 (N_36235,N_35828,N_35621);
and U36236 (N_36236,N_35886,N_35938);
and U36237 (N_36237,N_35607,N_35591);
xnor U36238 (N_36238,N_35604,N_35977);
nor U36239 (N_36239,N_35882,N_35665);
xor U36240 (N_36240,N_35599,N_35679);
nor U36241 (N_36241,N_35955,N_35898);
nand U36242 (N_36242,N_35757,N_35789);
or U36243 (N_36243,N_35730,N_35896);
and U36244 (N_36244,N_35590,N_35605);
nand U36245 (N_36245,N_35943,N_35880);
and U36246 (N_36246,N_35545,N_35720);
nor U36247 (N_36247,N_35814,N_35844);
and U36248 (N_36248,N_35691,N_35524);
and U36249 (N_36249,N_35667,N_35991);
or U36250 (N_36250,N_35981,N_35638);
and U36251 (N_36251,N_35775,N_35851);
xor U36252 (N_36252,N_35842,N_35658);
or U36253 (N_36253,N_35768,N_35733);
xnor U36254 (N_36254,N_35542,N_35757);
nor U36255 (N_36255,N_35748,N_35785);
nand U36256 (N_36256,N_35733,N_35867);
nor U36257 (N_36257,N_35660,N_35752);
and U36258 (N_36258,N_35843,N_35862);
nand U36259 (N_36259,N_35936,N_35791);
xor U36260 (N_36260,N_35802,N_35503);
and U36261 (N_36261,N_35619,N_35737);
nor U36262 (N_36262,N_35828,N_35909);
nand U36263 (N_36263,N_35998,N_35860);
or U36264 (N_36264,N_35918,N_35969);
nor U36265 (N_36265,N_35667,N_35631);
nand U36266 (N_36266,N_35700,N_35545);
or U36267 (N_36267,N_35839,N_35586);
or U36268 (N_36268,N_35790,N_35945);
and U36269 (N_36269,N_35677,N_35760);
or U36270 (N_36270,N_35556,N_35529);
nand U36271 (N_36271,N_35625,N_35873);
xor U36272 (N_36272,N_35526,N_35885);
nand U36273 (N_36273,N_35694,N_35515);
nand U36274 (N_36274,N_35677,N_35675);
nand U36275 (N_36275,N_35759,N_35690);
nand U36276 (N_36276,N_35956,N_35542);
and U36277 (N_36277,N_35626,N_35886);
or U36278 (N_36278,N_35746,N_35990);
xor U36279 (N_36279,N_35688,N_35722);
nand U36280 (N_36280,N_35920,N_35786);
and U36281 (N_36281,N_35909,N_35675);
xnor U36282 (N_36282,N_35626,N_35573);
xor U36283 (N_36283,N_35558,N_35923);
nor U36284 (N_36284,N_35623,N_35775);
nor U36285 (N_36285,N_35566,N_35984);
or U36286 (N_36286,N_35540,N_35884);
xnor U36287 (N_36287,N_35991,N_35587);
or U36288 (N_36288,N_35684,N_35858);
nand U36289 (N_36289,N_35755,N_35575);
xor U36290 (N_36290,N_35921,N_35699);
and U36291 (N_36291,N_35760,N_35695);
or U36292 (N_36292,N_35972,N_35624);
and U36293 (N_36293,N_35692,N_35986);
nand U36294 (N_36294,N_35972,N_35646);
nor U36295 (N_36295,N_35967,N_35580);
xnor U36296 (N_36296,N_35602,N_35778);
or U36297 (N_36297,N_35581,N_35962);
or U36298 (N_36298,N_35734,N_35978);
or U36299 (N_36299,N_35915,N_35836);
xnor U36300 (N_36300,N_35805,N_35840);
xor U36301 (N_36301,N_35584,N_35678);
nand U36302 (N_36302,N_35961,N_35813);
nor U36303 (N_36303,N_35824,N_35656);
and U36304 (N_36304,N_35638,N_35804);
or U36305 (N_36305,N_35908,N_35869);
nand U36306 (N_36306,N_35709,N_35756);
and U36307 (N_36307,N_35926,N_35619);
or U36308 (N_36308,N_35579,N_35855);
xor U36309 (N_36309,N_35514,N_35695);
xor U36310 (N_36310,N_35879,N_35844);
or U36311 (N_36311,N_35985,N_35903);
nand U36312 (N_36312,N_35544,N_35945);
or U36313 (N_36313,N_35579,N_35535);
nor U36314 (N_36314,N_35856,N_35716);
xor U36315 (N_36315,N_35582,N_35656);
nand U36316 (N_36316,N_35927,N_35841);
or U36317 (N_36317,N_35551,N_35625);
or U36318 (N_36318,N_35635,N_35890);
and U36319 (N_36319,N_35681,N_35545);
and U36320 (N_36320,N_35710,N_35866);
nor U36321 (N_36321,N_35651,N_35648);
or U36322 (N_36322,N_35862,N_35629);
xor U36323 (N_36323,N_35570,N_35696);
or U36324 (N_36324,N_35897,N_35850);
and U36325 (N_36325,N_35884,N_35806);
nor U36326 (N_36326,N_35966,N_35617);
or U36327 (N_36327,N_35817,N_35977);
and U36328 (N_36328,N_35648,N_35655);
xnor U36329 (N_36329,N_35527,N_35643);
nor U36330 (N_36330,N_35505,N_35645);
nor U36331 (N_36331,N_35966,N_35670);
xor U36332 (N_36332,N_35970,N_35795);
xor U36333 (N_36333,N_35923,N_35564);
or U36334 (N_36334,N_35572,N_35518);
xor U36335 (N_36335,N_35873,N_35734);
or U36336 (N_36336,N_35691,N_35952);
nor U36337 (N_36337,N_35674,N_35649);
or U36338 (N_36338,N_35832,N_35954);
nand U36339 (N_36339,N_35518,N_35629);
or U36340 (N_36340,N_35617,N_35529);
or U36341 (N_36341,N_35791,N_35751);
nor U36342 (N_36342,N_35717,N_35753);
nor U36343 (N_36343,N_35625,N_35787);
nor U36344 (N_36344,N_35574,N_35731);
or U36345 (N_36345,N_35597,N_35550);
or U36346 (N_36346,N_35954,N_35885);
xor U36347 (N_36347,N_35963,N_35686);
nand U36348 (N_36348,N_35617,N_35570);
nor U36349 (N_36349,N_35863,N_35970);
nor U36350 (N_36350,N_35625,N_35883);
and U36351 (N_36351,N_35617,N_35677);
xnor U36352 (N_36352,N_35730,N_35799);
nor U36353 (N_36353,N_35922,N_35546);
or U36354 (N_36354,N_35982,N_35511);
or U36355 (N_36355,N_35685,N_35652);
nand U36356 (N_36356,N_35893,N_35788);
nor U36357 (N_36357,N_35769,N_35796);
xnor U36358 (N_36358,N_35818,N_35896);
nor U36359 (N_36359,N_35609,N_35893);
and U36360 (N_36360,N_35939,N_35540);
nand U36361 (N_36361,N_35606,N_35776);
or U36362 (N_36362,N_35625,N_35710);
and U36363 (N_36363,N_35992,N_35868);
nor U36364 (N_36364,N_35859,N_35518);
and U36365 (N_36365,N_35769,N_35875);
nand U36366 (N_36366,N_35594,N_35896);
nand U36367 (N_36367,N_35556,N_35588);
xor U36368 (N_36368,N_35791,N_35624);
or U36369 (N_36369,N_35999,N_35619);
nand U36370 (N_36370,N_35725,N_35969);
nor U36371 (N_36371,N_35739,N_35814);
nand U36372 (N_36372,N_35554,N_35726);
or U36373 (N_36373,N_35655,N_35563);
xnor U36374 (N_36374,N_35613,N_35602);
xnor U36375 (N_36375,N_35706,N_35630);
and U36376 (N_36376,N_35970,N_35846);
xor U36377 (N_36377,N_35661,N_35692);
nor U36378 (N_36378,N_35709,N_35695);
or U36379 (N_36379,N_35518,N_35874);
or U36380 (N_36380,N_35525,N_35704);
and U36381 (N_36381,N_35848,N_35570);
or U36382 (N_36382,N_35669,N_35692);
xnor U36383 (N_36383,N_35575,N_35543);
and U36384 (N_36384,N_35748,N_35732);
and U36385 (N_36385,N_35571,N_35656);
nor U36386 (N_36386,N_35652,N_35828);
nand U36387 (N_36387,N_35613,N_35527);
nor U36388 (N_36388,N_35675,N_35633);
or U36389 (N_36389,N_35715,N_35762);
and U36390 (N_36390,N_35890,N_35785);
xnor U36391 (N_36391,N_35720,N_35690);
nand U36392 (N_36392,N_35934,N_35624);
and U36393 (N_36393,N_35786,N_35659);
nor U36394 (N_36394,N_35898,N_35826);
xor U36395 (N_36395,N_35750,N_35708);
or U36396 (N_36396,N_35813,N_35922);
nor U36397 (N_36397,N_35818,N_35878);
nand U36398 (N_36398,N_35761,N_35989);
nor U36399 (N_36399,N_35715,N_35790);
xnor U36400 (N_36400,N_35654,N_35845);
xor U36401 (N_36401,N_35590,N_35698);
nor U36402 (N_36402,N_35793,N_35988);
nand U36403 (N_36403,N_35929,N_35879);
xor U36404 (N_36404,N_35593,N_35701);
xor U36405 (N_36405,N_35929,N_35595);
nand U36406 (N_36406,N_35924,N_35938);
nor U36407 (N_36407,N_35699,N_35591);
or U36408 (N_36408,N_35526,N_35908);
or U36409 (N_36409,N_35656,N_35575);
nor U36410 (N_36410,N_35855,N_35720);
or U36411 (N_36411,N_35667,N_35659);
and U36412 (N_36412,N_35737,N_35819);
or U36413 (N_36413,N_35910,N_35929);
or U36414 (N_36414,N_35827,N_35610);
xnor U36415 (N_36415,N_35793,N_35959);
or U36416 (N_36416,N_35636,N_35816);
nor U36417 (N_36417,N_35665,N_35670);
or U36418 (N_36418,N_35557,N_35752);
xnor U36419 (N_36419,N_35816,N_35502);
nor U36420 (N_36420,N_35715,N_35623);
or U36421 (N_36421,N_35621,N_35518);
and U36422 (N_36422,N_35993,N_35863);
and U36423 (N_36423,N_35847,N_35964);
nand U36424 (N_36424,N_35778,N_35517);
nor U36425 (N_36425,N_35963,N_35552);
or U36426 (N_36426,N_35792,N_35575);
and U36427 (N_36427,N_35836,N_35845);
and U36428 (N_36428,N_35632,N_35973);
nand U36429 (N_36429,N_35621,N_35896);
xor U36430 (N_36430,N_35879,N_35583);
xor U36431 (N_36431,N_35934,N_35851);
nand U36432 (N_36432,N_35524,N_35931);
or U36433 (N_36433,N_35659,N_35742);
or U36434 (N_36434,N_35692,N_35861);
nand U36435 (N_36435,N_35884,N_35839);
or U36436 (N_36436,N_35648,N_35644);
nor U36437 (N_36437,N_35950,N_35879);
nand U36438 (N_36438,N_35506,N_35870);
or U36439 (N_36439,N_35872,N_35566);
or U36440 (N_36440,N_35626,N_35608);
and U36441 (N_36441,N_35900,N_35978);
xnor U36442 (N_36442,N_35700,N_35901);
nand U36443 (N_36443,N_35720,N_35541);
nand U36444 (N_36444,N_35591,N_35754);
nand U36445 (N_36445,N_35773,N_35599);
xor U36446 (N_36446,N_35709,N_35974);
xor U36447 (N_36447,N_35983,N_35603);
and U36448 (N_36448,N_35843,N_35719);
xor U36449 (N_36449,N_35981,N_35608);
or U36450 (N_36450,N_35734,N_35532);
nand U36451 (N_36451,N_35840,N_35950);
or U36452 (N_36452,N_35976,N_35811);
and U36453 (N_36453,N_35812,N_35787);
xnor U36454 (N_36454,N_35519,N_35824);
nor U36455 (N_36455,N_35558,N_35773);
or U36456 (N_36456,N_35893,N_35524);
nor U36457 (N_36457,N_35628,N_35563);
or U36458 (N_36458,N_35938,N_35596);
xor U36459 (N_36459,N_35762,N_35508);
and U36460 (N_36460,N_35608,N_35515);
nand U36461 (N_36461,N_35998,N_35935);
nand U36462 (N_36462,N_35533,N_35580);
nor U36463 (N_36463,N_35592,N_35895);
or U36464 (N_36464,N_35669,N_35747);
and U36465 (N_36465,N_35546,N_35605);
nand U36466 (N_36466,N_35669,N_35832);
and U36467 (N_36467,N_35521,N_35830);
nor U36468 (N_36468,N_35610,N_35917);
xnor U36469 (N_36469,N_35548,N_35700);
nand U36470 (N_36470,N_35964,N_35950);
nand U36471 (N_36471,N_35982,N_35932);
or U36472 (N_36472,N_35875,N_35568);
xnor U36473 (N_36473,N_35728,N_35597);
and U36474 (N_36474,N_35576,N_35833);
and U36475 (N_36475,N_35862,N_35733);
and U36476 (N_36476,N_35947,N_35958);
nand U36477 (N_36477,N_35662,N_35643);
xor U36478 (N_36478,N_35661,N_35920);
xor U36479 (N_36479,N_35599,N_35652);
and U36480 (N_36480,N_35519,N_35768);
and U36481 (N_36481,N_35536,N_35535);
or U36482 (N_36482,N_35921,N_35867);
and U36483 (N_36483,N_35956,N_35898);
and U36484 (N_36484,N_35938,N_35508);
nor U36485 (N_36485,N_35880,N_35912);
nor U36486 (N_36486,N_35731,N_35694);
nor U36487 (N_36487,N_35573,N_35854);
and U36488 (N_36488,N_35606,N_35623);
or U36489 (N_36489,N_35855,N_35889);
and U36490 (N_36490,N_35664,N_35624);
nand U36491 (N_36491,N_35706,N_35722);
or U36492 (N_36492,N_35937,N_35570);
nand U36493 (N_36493,N_35970,N_35694);
or U36494 (N_36494,N_35697,N_35910);
and U36495 (N_36495,N_35959,N_35704);
or U36496 (N_36496,N_35865,N_35626);
nor U36497 (N_36497,N_35887,N_35830);
nor U36498 (N_36498,N_35793,N_35756);
or U36499 (N_36499,N_35582,N_35918);
nand U36500 (N_36500,N_36015,N_36235);
xor U36501 (N_36501,N_36326,N_36187);
nor U36502 (N_36502,N_36372,N_36219);
and U36503 (N_36503,N_36122,N_36100);
nand U36504 (N_36504,N_36358,N_36247);
nand U36505 (N_36505,N_36249,N_36420);
nor U36506 (N_36506,N_36340,N_36485);
nor U36507 (N_36507,N_36246,N_36378);
nor U36508 (N_36508,N_36224,N_36268);
nor U36509 (N_36509,N_36415,N_36269);
nor U36510 (N_36510,N_36201,N_36162);
xnor U36511 (N_36511,N_36003,N_36085);
nor U36512 (N_36512,N_36440,N_36359);
and U36513 (N_36513,N_36321,N_36193);
nor U36514 (N_36514,N_36237,N_36091);
nand U36515 (N_36515,N_36116,N_36059);
and U36516 (N_36516,N_36203,N_36484);
and U36517 (N_36517,N_36238,N_36044);
or U36518 (N_36518,N_36006,N_36035);
nand U36519 (N_36519,N_36400,N_36087);
xnor U36520 (N_36520,N_36318,N_36094);
and U36521 (N_36521,N_36121,N_36433);
xor U36522 (N_36522,N_36153,N_36351);
nor U36523 (N_36523,N_36336,N_36478);
nand U36524 (N_36524,N_36434,N_36045);
nor U36525 (N_36525,N_36446,N_36226);
xnor U36526 (N_36526,N_36084,N_36458);
nor U36527 (N_36527,N_36215,N_36254);
nand U36528 (N_36528,N_36441,N_36324);
nor U36529 (N_36529,N_36210,N_36236);
and U36530 (N_36530,N_36171,N_36407);
nand U36531 (N_36531,N_36075,N_36480);
and U36532 (N_36532,N_36453,N_36463);
or U36533 (N_36533,N_36472,N_36342);
and U36534 (N_36534,N_36048,N_36167);
and U36535 (N_36535,N_36448,N_36209);
nor U36536 (N_36536,N_36253,N_36160);
and U36537 (N_36537,N_36142,N_36169);
nand U36538 (N_36538,N_36114,N_36239);
nand U36539 (N_36539,N_36288,N_36287);
xnor U36540 (N_36540,N_36362,N_36089);
nor U36541 (N_36541,N_36431,N_36406);
xor U36542 (N_36542,N_36289,N_36390);
and U36543 (N_36543,N_36454,N_36218);
nand U36544 (N_36544,N_36310,N_36261);
or U36545 (N_36545,N_36469,N_36341);
nor U36546 (N_36546,N_36018,N_36387);
and U36547 (N_36547,N_36056,N_36497);
nand U36548 (N_36548,N_36012,N_36216);
or U36549 (N_36549,N_36128,N_36119);
or U36550 (N_36550,N_36275,N_36135);
xor U36551 (N_36551,N_36071,N_36063);
xor U36552 (N_36552,N_36042,N_36429);
nor U36553 (N_36553,N_36147,N_36335);
nand U36554 (N_36554,N_36081,N_36284);
and U36555 (N_36555,N_36319,N_36107);
or U36556 (N_36556,N_36328,N_36248);
or U36557 (N_36557,N_36136,N_36489);
or U36558 (N_36558,N_36233,N_36205);
nand U36559 (N_36559,N_36138,N_36230);
and U36560 (N_36560,N_36240,N_36402);
nand U36561 (N_36561,N_36314,N_36461);
nor U36562 (N_36562,N_36380,N_36041);
and U36563 (N_36563,N_36047,N_36130);
nor U36564 (N_36564,N_36159,N_36143);
xnor U36565 (N_36565,N_36115,N_36439);
nor U36566 (N_36566,N_36363,N_36225);
and U36567 (N_36567,N_36192,N_36140);
nand U36568 (N_36568,N_36421,N_36376);
nor U36569 (N_36569,N_36029,N_36399);
or U36570 (N_36570,N_36197,N_36060);
nor U36571 (N_36571,N_36290,N_36090);
xnor U36572 (N_36572,N_36120,N_36105);
and U36573 (N_36573,N_36002,N_36316);
nor U36574 (N_36574,N_36255,N_36432);
or U36575 (N_36575,N_36353,N_36293);
and U36576 (N_36576,N_36021,N_36391);
xnor U36577 (N_36577,N_36086,N_36337);
nor U36578 (N_36578,N_36104,N_36493);
nand U36579 (N_36579,N_36082,N_36451);
and U36580 (N_36580,N_36212,N_36026);
nand U36581 (N_36581,N_36036,N_36334);
nor U36582 (N_36582,N_36260,N_36279);
nand U36583 (N_36583,N_36039,N_36118);
and U36584 (N_36584,N_36152,N_36103);
or U36585 (N_36585,N_36196,N_36349);
or U36586 (N_36586,N_36061,N_36250);
or U36587 (N_36587,N_36266,N_36297);
nand U36588 (N_36588,N_36070,N_36345);
nor U36589 (N_36589,N_36031,N_36179);
nand U36590 (N_36590,N_36076,N_36490);
xor U36591 (N_36591,N_36055,N_36096);
nor U36592 (N_36592,N_36329,N_36356);
and U36593 (N_36593,N_36207,N_36473);
nand U36594 (N_36594,N_36127,N_36146);
nor U36595 (N_36595,N_36355,N_36418);
nor U36596 (N_36596,N_36456,N_36397);
or U36597 (N_36597,N_36243,N_36327);
nand U36598 (N_36598,N_36113,N_36294);
nand U36599 (N_36599,N_36189,N_36264);
and U36600 (N_36600,N_36220,N_36200);
xor U36601 (N_36601,N_36457,N_36459);
and U36602 (N_36602,N_36027,N_36257);
nor U36603 (N_36603,N_36148,N_36123);
nand U36604 (N_36604,N_36270,N_36190);
nor U36605 (N_36605,N_36384,N_36483);
nor U36606 (N_36606,N_36206,N_36126);
nor U36607 (N_36607,N_36401,N_36178);
xnor U36608 (N_36608,N_36155,N_36109);
nor U36609 (N_36609,N_36424,N_36292);
xor U36610 (N_36610,N_36422,N_36038);
and U36611 (N_36611,N_36204,N_36156);
nand U36612 (N_36612,N_36168,N_36030);
and U36613 (N_36613,N_36371,N_36277);
nand U36614 (N_36614,N_36004,N_36442);
xnor U36615 (N_36615,N_36227,N_36447);
nand U36616 (N_36616,N_36022,N_36377);
nor U36617 (N_36617,N_36110,N_36487);
xnor U36618 (N_36618,N_36283,N_36419);
and U36619 (N_36619,N_36373,N_36450);
or U36620 (N_36620,N_36476,N_36049);
xnor U36621 (N_36621,N_36409,N_36182);
and U36622 (N_36622,N_36242,N_36479);
nand U36623 (N_36623,N_36317,N_36073);
xor U36624 (N_36624,N_36033,N_36217);
nor U36625 (N_36625,N_36129,N_36330);
nand U36626 (N_36626,N_36062,N_36374);
or U36627 (N_36627,N_36097,N_36028);
nor U36628 (N_36628,N_36010,N_36369);
or U36629 (N_36629,N_36477,N_36436);
or U36630 (N_36630,N_36065,N_36000);
nor U36631 (N_36631,N_36111,N_36304);
nor U36632 (N_36632,N_36396,N_36428);
nor U36633 (N_36633,N_36185,N_36364);
nand U36634 (N_36634,N_36017,N_36092);
or U36635 (N_36635,N_36339,N_36455);
or U36636 (N_36636,N_36410,N_36393);
or U36637 (N_36637,N_36106,N_36367);
xor U36638 (N_36638,N_36079,N_36306);
xor U36639 (N_36639,N_36199,N_36058);
nor U36640 (N_36640,N_36414,N_36430);
and U36641 (N_36641,N_36232,N_36214);
or U36642 (N_36642,N_36379,N_36208);
or U36643 (N_36643,N_36037,N_36361);
xnor U36644 (N_36644,N_36481,N_36053);
xor U36645 (N_36645,N_36173,N_36299);
nand U36646 (N_36646,N_36170,N_36191);
nor U36647 (N_36647,N_36005,N_36386);
nand U36648 (N_36648,N_36174,N_36176);
or U36649 (N_36649,N_36001,N_36093);
nand U36650 (N_36650,N_36050,N_36375);
nor U36651 (N_36651,N_36425,N_36144);
xnor U36652 (N_36652,N_36300,N_36470);
and U36653 (N_36653,N_36382,N_36252);
or U36654 (N_36654,N_36404,N_36282);
or U36655 (N_36655,N_36389,N_36405);
or U36656 (N_36656,N_36273,N_36009);
and U36657 (N_36657,N_36007,N_36437);
nor U36658 (N_36658,N_36271,N_36040);
and U36659 (N_36659,N_36435,N_36020);
or U36660 (N_36660,N_36354,N_36098);
nor U36661 (N_36661,N_36468,N_36417);
or U36662 (N_36662,N_36411,N_36475);
nand U36663 (N_36663,N_36262,N_36449);
xnor U36664 (N_36664,N_36496,N_36211);
and U36665 (N_36665,N_36080,N_36259);
nand U36666 (N_36666,N_36068,N_36256);
nand U36667 (N_36667,N_36149,N_36231);
or U36668 (N_36668,N_36057,N_36443);
nand U36669 (N_36669,N_36408,N_36198);
nand U36670 (N_36670,N_36278,N_36308);
nand U36671 (N_36671,N_36333,N_36108);
xor U36672 (N_36672,N_36019,N_36014);
nand U36673 (N_36673,N_36311,N_36460);
and U36674 (N_36674,N_36370,N_36072);
nor U36675 (N_36675,N_36445,N_36054);
or U36676 (N_36676,N_36423,N_36157);
and U36677 (N_36677,N_36350,N_36462);
nand U36678 (N_36678,N_36357,N_36348);
xor U36679 (N_36679,N_36325,N_36180);
and U36680 (N_36680,N_36125,N_36366);
nand U36681 (N_36681,N_36385,N_36088);
nor U36682 (N_36682,N_36141,N_36438);
nor U36683 (N_36683,N_36024,N_36352);
and U36684 (N_36684,N_36307,N_36303);
nor U36685 (N_36685,N_36474,N_36301);
xor U36686 (N_36686,N_36295,N_36222);
xor U36687 (N_36687,N_36172,N_36465);
or U36688 (N_36688,N_36427,N_36139);
or U36689 (N_36689,N_36181,N_36343);
and U36690 (N_36690,N_36360,N_36285);
nor U36691 (N_36691,N_36263,N_36154);
and U36692 (N_36692,N_36313,N_36486);
nand U36693 (N_36693,N_36046,N_36272);
nor U36694 (N_36694,N_36258,N_36016);
nand U36695 (N_36695,N_36347,N_36471);
nand U36696 (N_36696,N_36346,N_36078);
nor U36697 (N_36697,N_36467,N_36101);
and U36698 (N_36698,N_36134,N_36368);
nand U36699 (N_36699,N_36151,N_36495);
and U36700 (N_36700,N_36083,N_36499);
and U36701 (N_36701,N_36488,N_36183);
nand U36702 (N_36702,N_36395,N_36320);
or U36703 (N_36703,N_36164,N_36286);
xnor U36704 (N_36704,N_36161,N_36112);
or U36705 (N_36705,N_36145,N_36381);
and U36706 (N_36706,N_36133,N_36202);
nor U36707 (N_36707,N_36194,N_36344);
or U36708 (N_36708,N_36392,N_36426);
xor U36709 (N_36709,N_36163,N_36281);
nand U36710 (N_36710,N_36280,N_36131);
or U36711 (N_36711,N_36186,N_36265);
nor U36712 (N_36712,N_36025,N_36064);
or U36713 (N_36713,N_36195,N_36498);
nand U36714 (N_36714,N_36305,N_36452);
xnor U36715 (N_36715,N_36267,N_36365);
or U36716 (N_36716,N_36312,N_36034);
and U36717 (N_36717,N_36051,N_36464);
and U36718 (N_36718,N_36388,N_36132);
and U36719 (N_36719,N_36245,N_36221);
or U36720 (N_36720,N_36066,N_36175);
and U36721 (N_36721,N_36032,N_36077);
nand U36722 (N_36722,N_36309,N_36166);
and U36723 (N_36723,N_36332,N_36124);
nand U36724 (N_36724,N_36150,N_36315);
xnor U36725 (N_36725,N_36416,N_36492);
nor U36726 (N_36726,N_36412,N_36069);
nor U36727 (N_36727,N_36177,N_36117);
and U36728 (N_36728,N_36229,N_36067);
xor U36729 (N_36729,N_36466,N_36491);
xnor U36730 (N_36730,N_36296,N_36482);
and U36731 (N_36731,N_36234,N_36137);
nor U36732 (N_36732,N_36008,N_36095);
nand U36733 (N_36733,N_36074,N_36291);
xor U36734 (N_36734,N_36158,N_36013);
or U36735 (N_36735,N_36241,N_36188);
xnor U36736 (N_36736,N_36338,N_36276);
xnor U36737 (N_36737,N_36213,N_36444);
or U36738 (N_36738,N_36099,N_36394);
nand U36739 (N_36739,N_36494,N_36398);
or U36740 (N_36740,N_36102,N_36011);
nand U36741 (N_36741,N_36023,N_36052);
nor U36742 (N_36742,N_36403,N_36184);
nand U36743 (N_36743,N_36413,N_36043);
and U36744 (N_36744,N_36251,N_36274);
xnor U36745 (N_36745,N_36331,N_36165);
xnor U36746 (N_36746,N_36223,N_36322);
nand U36747 (N_36747,N_36244,N_36228);
or U36748 (N_36748,N_36383,N_36298);
nor U36749 (N_36749,N_36302,N_36323);
or U36750 (N_36750,N_36096,N_36471);
nor U36751 (N_36751,N_36213,N_36399);
nand U36752 (N_36752,N_36122,N_36319);
xnor U36753 (N_36753,N_36083,N_36380);
nor U36754 (N_36754,N_36123,N_36037);
nand U36755 (N_36755,N_36461,N_36409);
nor U36756 (N_36756,N_36437,N_36055);
nand U36757 (N_36757,N_36368,N_36338);
nand U36758 (N_36758,N_36305,N_36241);
nor U36759 (N_36759,N_36245,N_36124);
nor U36760 (N_36760,N_36270,N_36303);
nand U36761 (N_36761,N_36210,N_36020);
nor U36762 (N_36762,N_36080,N_36316);
nand U36763 (N_36763,N_36144,N_36361);
nand U36764 (N_36764,N_36189,N_36304);
xnor U36765 (N_36765,N_36276,N_36439);
and U36766 (N_36766,N_36129,N_36009);
nor U36767 (N_36767,N_36340,N_36002);
and U36768 (N_36768,N_36088,N_36059);
and U36769 (N_36769,N_36088,N_36294);
nor U36770 (N_36770,N_36019,N_36321);
and U36771 (N_36771,N_36007,N_36063);
xor U36772 (N_36772,N_36103,N_36049);
or U36773 (N_36773,N_36079,N_36029);
xnor U36774 (N_36774,N_36322,N_36299);
xor U36775 (N_36775,N_36322,N_36140);
nand U36776 (N_36776,N_36047,N_36166);
nor U36777 (N_36777,N_36255,N_36457);
nor U36778 (N_36778,N_36056,N_36076);
and U36779 (N_36779,N_36373,N_36214);
nor U36780 (N_36780,N_36348,N_36246);
xor U36781 (N_36781,N_36095,N_36137);
xor U36782 (N_36782,N_36235,N_36323);
nor U36783 (N_36783,N_36178,N_36461);
and U36784 (N_36784,N_36456,N_36355);
xnor U36785 (N_36785,N_36126,N_36349);
and U36786 (N_36786,N_36308,N_36198);
nand U36787 (N_36787,N_36349,N_36108);
nand U36788 (N_36788,N_36126,N_36276);
nand U36789 (N_36789,N_36352,N_36453);
nand U36790 (N_36790,N_36429,N_36408);
or U36791 (N_36791,N_36204,N_36367);
xor U36792 (N_36792,N_36029,N_36080);
or U36793 (N_36793,N_36257,N_36164);
nand U36794 (N_36794,N_36337,N_36466);
xor U36795 (N_36795,N_36107,N_36258);
or U36796 (N_36796,N_36090,N_36248);
nor U36797 (N_36797,N_36235,N_36447);
nand U36798 (N_36798,N_36291,N_36067);
nand U36799 (N_36799,N_36079,N_36350);
nor U36800 (N_36800,N_36190,N_36123);
or U36801 (N_36801,N_36281,N_36332);
or U36802 (N_36802,N_36091,N_36382);
or U36803 (N_36803,N_36079,N_36321);
xor U36804 (N_36804,N_36401,N_36303);
nor U36805 (N_36805,N_36295,N_36255);
or U36806 (N_36806,N_36390,N_36092);
xnor U36807 (N_36807,N_36450,N_36115);
xnor U36808 (N_36808,N_36368,N_36170);
nor U36809 (N_36809,N_36244,N_36140);
and U36810 (N_36810,N_36026,N_36041);
nand U36811 (N_36811,N_36150,N_36090);
or U36812 (N_36812,N_36395,N_36088);
nor U36813 (N_36813,N_36172,N_36311);
nand U36814 (N_36814,N_36063,N_36067);
or U36815 (N_36815,N_36409,N_36267);
or U36816 (N_36816,N_36292,N_36436);
or U36817 (N_36817,N_36331,N_36164);
nor U36818 (N_36818,N_36077,N_36052);
nor U36819 (N_36819,N_36373,N_36080);
nor U36820 (N_36820,N_36117,N_36340);
or U36821 (N_36821,N_36153,N_36393);
or U36822 (N_36822,N_36164,N_36387);
or U36823 (N_36823,N_36166,N_36124);
xor U36824 (N_36824,N_36490,N_36487);
nor U36825 (N_36825,N_36194,N_36461);
xor U36826 (N_36826,N_36459,N_36366);
or U36827 (N_36827,N_36336,N_36212);
nand U36828 (N_36828,N_36192,N_36406);
xnor U36829 (N_36829,N_36278,N_36256);
and U36830 (N_36830,N_36296,N_36179);
nand U36831 (N_36831,N_36073,N_36312);
xor U36832 (N_36832,N_36076,N_36302);
or U36833 (N_36833,N_36176,N_36461);
xor U36834 (N_36834,N_36059,N_36327);
nor U36835 (N_36835,N_36186,N_36445);
nand U36836 (N_36836,N_36315,N_36163);
nand U36837 (N_36837,N_36034,N_36234);
xnor U36838 (N_36838,N_36172,N_36366);
or U36839 (N_36839,N_36337,N_36228);
nand U36840 (N_36840,N_36291,N_36337);
xor U36841 (N_36841,N_36281,N_36130);
and U36842 (N_36842,N_36146,N_36423);
or U36843 (N_36843,N_36032,N_36368);
xor U36844 (N_36844,N_36429,N_36251);
or U36845 (N_36845,N_36394,N_36123);
xor U36846 (N_36846,N_36317,N_36392);
nor U36847 (N_36847,N_36024,N_36008);
xor U36848 (N_36848,N_36377,N_36275);
nor U36849 (N_36849,N_36497,N_36025);
and U36850 (N_36850,N_36299,N_36068);
nand U36851 (N_36851,N_36025,N_36029);
nor U36852 (N_36852,N_36108,N_36142);
xnor U36853 (N_36853,N_36478,N_36205);
xor U36854 (N_36854,N_36147,N_36065);
and U36855 (N_36855,N_36004,N_36308);
xnor U36856 (N_36856,N_36209,N_36410);
nand U36857 (N_36857,N_36010,N_36034);
and U36858 (N_36858,N_36344,N_36193);
nand U36859 (N_36859,N_36244,N_36452);
nor U36860 (N_36860,N_36267,N_36490);
nand U36861 (N_36861,N_36415,N_36385);
and U36862 (N_36862,N_36419,N_36238);
nor U36863 (N_36863,N_36209,N_36202);
and U36864 (N_36864,N_36349,N_36119);
nor U36865 (N_36865,N_36355,N_36251);
nor U36866 (N_36866,N_36028,N_36496);
and U36867 (N_36867,N_36365,N_36366);
xnor U36868 (N_36868,N_36460,N_36209);
nor U36869 (N_36869,N_36344,N_36348);
nand U36870 (N_36870,N_36165,N_36322);
xor U36871 (N_36871,N_36128,N_36349);
xor U36872 (N_36872,N_36220,N_36356);
or U36873 (N_36873,N_36380,N_36323);
xor U36874 (N_36874,N_36387,N_36205);
nor U36875 (N_36875,N_36040,N_36421);
or U36876 (N_36876,N_36092,N_36033);
and U36877 (N_36877,N_36112,N_36446);
nand U36878 (N_36878,N_36167,N_36161);
nand U36879 (N_36879,N_36209,N_36165);
nand U36880 (N_36880,N_36451,N_36487);
nand U36881 (N_36881,N_36001,N_36236);
nor U36882 (N_36882,N_36454,N_36248);
and U36883 (N_36883,N_36361,N_36001);
nand U36884 (N_36884,N_36038,N_36194);
or U36885 (N_36885,N_36475,N_36222);
and U36886 (N_36886,N_36350,N_36480);
nor U36887 (N_36887,N_36251,N_36473);
or U36888 (N_36888,N_36170,N_36121);
or U36889 (N_36889,N_36403,N_36365);
or U36890 (N_36890,N_36000,N_36261);
xnor U36891 (N_36891,N_36051,N_36079);
or U36892 (N_36892,N_36485,N_36433);
and U36893 (N_36893,N_36384,N_36017);
nor U36894 (N_36894,N_36151,N_36136);
xnor U36895 (N_36895,N_36478,N_36198);
xor U36896 (N_36896,N_36282,N_36102);
nor U36897 (N_36897,N_36202,N_36236);
and U36898 (N_36898,N_36114,N_36067);
xnor U36899 (N_36899,N_36158,N_36285);
or U36900 (N_36900,N_36440,N_36339);
xnor U36901 (N_36901,N_36403,N_36399);
nor U36902 (N_36902,N_36245,N_36332);
nor U36903 (N_36903,N_36371,N_36307);
nand U36904 (N_36904,N_36017,N_36388);
nor U36905 (N_36905,N_36134,N_36176);
and U36906 (N_36906,N_36310,N_36293);
and U36907 (N_36907,N_36099,N_36007);
and U36908 (N_36908,N_36092,N_36481);
or U36909 (N_36909,N_36333,N_36317);
xnor U36910 (N_36910,N_36335,N_36416);
xnor U36911 (N_36911,N_36096,N_36056);
nor U36912 (N_36912,N_36242,N_36108);
xnor U36913 (N_36913,N_36217,N_36332);
nand U36914 (N_36914,N_36458,N_36295);
nor U36915 (N_36915,N_36151,N_36177);
nand U36916 (N_36916,N_36438,N_36267);
nor U36917 (N_36917,N_36138,N_36099);
xnor U36918 (N_36918,N_36402,N_36152);
xor U36919 (N_36919,N_36238,N_36172);
nor U36920 (N_36920,N_36452,N_36462);
or U36921 (N_36921,N_36095,N_36437);
nor U36922 (N_36922,N_36444,N_36454);
xnor U36923 (N_36923,N_36178,N_36388);
or U36924 (N_36924,N_36291,N_36458);
nor U36925 (N_36925,N_36003,N_36220);
xor U36926 (N_36926,N_36005,N_36222);
and U36927 (N_36927,N_36128,N_36290);
nand U36928 (N_36928,N_36483,N_36244);
xor U36929 (N_36929,N_36463,N_36292);
nor U36930 (N_36930,N_36477,N_36160);
and U36931 (N_36931,N_36305,N_36187);
nor U36932 (N_36932,N_36050,N_36001);
and U36933 (N_36933,N_36336,N_36120);
nand U36934 (N_36934,N_36149,N_36329);
nand U36935 (N_36935,N_36193,N_36234);
nor U36936 (N_36936,N_36067,N_36253);
nand U36937 (N_36937,N_36265,N_36334);
nor U36938 (N_36938,N_36259,N_36017);
and U36939 (N_36939,N_36080,N_36062);
nand U36940 (N_36940,N_36423,N_36228);
or U36941 (N_36941,N_36113,N_36093);
xor U36942 (N_36942,N_36218,N_36281);
xor U36943 (N_36943,N_36152,N_36232);
xor U36944 (N_36944,N_36389,N_36484);
xnor U36945 (N_36945,N_36116,N_36434);
nand U36946 (N_36946,N_36162,N_36003);
xnor U36947 (N_36947,N_36179,N_36379);
nand U36948 (N_36948,N_36421,N_36186);
or U36949 (N_36949,N_36123,N_36352);
or U36950 (N_36950,N_36178,N_36298);
and U36951 (N_36951,N_36324,N_36005);
and U36952 (N_36952,N_36205,N_36487);
and U36953 (N_36953,N_36290,N_36029);
or U36954 (N_36954,N_36202,N_36210);
nor U36955 (N_36955,N_36292,N_36394);
nand U36956 (N_36956,N_36444,N_36062);
or U36957 (N_36957,N_36201,N_36494);
and U36958 (N_36958,N_36121,N_36067);
xor U36959 (N_36959,N_36213,N_36075);
nand U36960 (N_36960,N_36420,N_36202);
and U36961 (N_36961,N_36107,N_36333);
xnor U36962 (N_36962,N_36262,N_36084);
or U36963 (N_36963,N_36416,N_36021);
and U36964 (N_36964,N_36473,N_36246);
xor U36965 (N_36965,N_36009,N_36358);
nand U36966 (N_36966,N_36099,N_36336);
and U36967 (N_36967,N_36489,N_36497);
nand U36968 (N_36968,N_36094,N_36043);
nand U36969 (N_36969,N_36124,N_36071);
nor U36970 (N_36970,N_36274,N_36219);
xnor U36971 (N_36971,N_36095,N_36334);
nor U36972 (N_36972,N_36338,N_36470);
nand U36973 (N_36973,N_36435,N_36474);
nand U36974 (N_36974,N_36484,N_36078);
nand U36975 (N_36975,N_36236,N_36032);
or U36976 (N_36976,N_36460,N_36121);
xnor U36977 (N_36977,N_36181,N_36013);
or U36978 (N_36978,N_36456,N_36168);
or U36979 (N_36979,N_36190,N_36311);
or U36980 (N_36980,N_36174,N_36288);
nor U36981 (N_36981,N_36390,N_36076);
nand U36982 (N_36982,N_36461,N_36089);
nand U36983 (N_36983,N_36022,N_36440);
nor U36984 (N_36984,N_36478,N_36347);
xnor U36985 (N_36985,N_36057,N_36016);
nand U36986 (N_36986,N_36157,N_36020);
and U36987 (N_36987,N_36206,N_36396);
or U36988 (N_36988,N_36279,N_36390);
nor U36989 (N_36989,N_36055,N_36214);
or U36990 (N_36990,N_36487,N_36497);
nor U36991 (N_36991,N_36037,N_36090);
and U36992 (N_36992,N_36255,N_36267);
nor U36993 (N_36993,N_36381,N_36172);
nor U36994 (N_36994,N_36246,N_36310);
nand U36995 (N_36995,N_36097,N_36345);
xor U36996 (N_36996,N_36268,N_36305);
nand U36997 (N_36997,N_36482,N_36295);
and U36998 (N_36998,N_36372,N_36418);
and U36999 (N_36999,N_36159,N_36430);
nand U37000 (N_37000,N_36575,N_36932);
xor U37001 (N_37001,N_36755,N_36509);
xor U37002 (N_37002,N_36614,N_36597);
or U37003 (N_37003,N_36517,N_36843);
xnor U37004 (N_37004,N_36834,N_36599);
nor U37005 (N_37005,N_36865,N_36516);
and U37006 (N_37006,N_36933,N_36812);
nor U37007 (N_37007,N_36892,N_36958);
or U37008 (N_37008,N_36605,N_36805);
nor U37009 (N_37009,N_36998,N_36734);
and U37010 (N_37010,N_36901,N_36867);
nor U37011 (N_37011,N_36866,N_36642);
or U37012 (N_37012,N_36583,N_36884);
and U37013 (N_37013,N_36612,N_36502);
xor U37014 (N_37014,N_36961,N_36592);
or U37015 (N_37015,N_36766,N_36858);
nand U37016 (N_37016,N_36915,N_36674);
or U37017 (N_37017,N_36800,N_36530);
nand U37018 (N_37018,N_36780,N_36620);
and U37019 (N_37019,N_36578,N_36665);
or U37020 (N_37020,N_36666,N_36576);
and U37021 (N_37021,N_36920,N_36754);
xnor U37022 (N_37022,N_36688,N_36524);
or U37023 (N_37023,N_36720,N_36750);
xnor U37024 (N_37024,N_36567,N_36954);
or U37025 (N_37025,N_36582,N_36927);
nand U37026 (N_37026,N_36994,N_36648);
nor U37027 (N_37027,N_36551,N_36783);
nand U37028 (N_37028,N_36633,N_36893);
nor U37029 (N_37029,N_36640,N_36598);
or U37030 (N_37030,N_36637,N_36775);
or U37031 (N_37031,N_36768,N_36773);
xor U37032 (N_37032,N_36760,N_36851);
xnor U37033 (N_37033,N_36917,N_36794);
or U37034 (N_37034,N_36822,N_36986);
nor U37035 (N_37035,N_36870,N_36903);
nand U37036 (N_37036,N_36788,N_36677);
or U37037 (N_37037,N_36727,N_36584);
nand U37038 (N_37038,N_36953,N_36859);
or U37039 (N_37039,N_36676,N_36504);
xor U37040 (N_37040,N_36748,N_36738);
nor U37041 (N_37041,N_36769,N_36619);
xnor U37042 (N_37042,N_36778,N_36847);
or U37043 (N_37043,N_36790,N_36852);
xor U37044 (N_37044,N_36532,N_36538);
nand U37045 (N_37045,N_36526,N_36549);
or U37046 (N_37046,N_36574,N_36781);
xnor U37047 (N_37047,N_36692,N_36730);
nor U37048 (N_37048,N_36772,N_36774);
and U37049 (N_37049,N_36959,N_36639);
and U37050 (N_37050,N_36891,N_36546);
or U37051 (N_37051,N_36879,N_36993);
nand U37052 (N_37052,N_36912,N_36815);
and U37053 (N_37053,N_36985,N_36797);
nor U37054 (N_37054,N_36736,N_36520);
or U37055 (N_37055,N_36793,N_36579);
nand U37056 (N_37056,N_36724,N_36806);
xor U37057 (N_37057,N_36675,N_36528);
xnor U37058 (N_37058,N_36798,N_36646);
xor U37059 (N_37059,N_36745,N_36647);
or U37060 (N_37060,N_36896,N_36918);
nor U37061 (N_37061,N_36659,N_36561);
or U37062 (N_37062,N_36924,N_36876);
xnor U37063 (N_37063,N_36623,N_36719);
and U37064 (N_37064,N_36632,N_36849);
nand U37065 (N_37065,N_36501,N_36808);
nand U37066 (N_37066,N_36919,N_36681);
or U37067 (N_37067,N_36537,N_36601);
nor U37068 (N_37068,N_36694,N_36706);
nor U37069 (N_37069,N_36973,N_36635);
nand U37070 (N_37070,N_36848,N_36506);
nand U37071 (N_37071,N_36697,N_36991);
or U37072 (N_37072,N_36861,N_36535);
nand U37073 (N_37073,N_36586,N_36789);
nand U37074 (N_37074,N_36934,N_36782);
nor U37075 (N_37075,N_36641,N_36820);
nor U37076 (N_37076,N_36824,N_36702);
or U37077 (N_37077,N_36515,N_36854);
nor U37078 (N_37078,N_36943,N_36568);
and U37079 (N_37079,N_36856,N_36764);
or U37080 (N_37080,N_36823,N_36952);
xor U37081 (N_37081,N_36591,N_36705);
or U37082 (N_37082,N_36761,N_36747);
xor U37083 (N_37083,N_36937,N_36984);
xnor U37084 (N_37084,N_36542,N_36946);
nor U37085 (N_37085,N_36617,N_36655);
or U37086 (N_37086,N_36547,N_36622);
nor U37087 (N_37087,N_36531,N_36616);
nor U37088 (N_37088,N_36644,N_36678);
xnor U37089 (N_37089,N_36949,N_36587);
and U37090 (N_37090,N_36603,N_36707);
and U37091 (N_37091,N_36828,N_36510);
xnor U37092 (N_37092,N_36691,N_36631);
nand U37093 (N_37093,N_36796,N_36540);
nand U37094 (N_37094,N_36850,N_36636);
and U37095 (N_37095,N_36767,N_36762);
nor U37096 (N_37096,N_36928,N_36875);
xor U37097 (N_37097,N_36552,N_36500);
or U37098 (N_37098,N_36672,N_36906);
nor U37099 (N_37099,N_36602,N_36723);
nand U37100 (N_37100,N_36731,N_36960);
and U37101 (N_37101,N_36844,N_36758);
nor U37102 (N_37102,N_36886,N_36590);
or U37103 (N_37103,N_36687,N_36975);
and U37104 (N_37104,N_36630,N_36779);
or U37105 (N_37105,N_36735,N_36698);
nand U37106 (N_37106,N_36787,N_36753);
xnor U37107 (N_37107,N_36657,N_36803);
nor U37108 (N_37108,N_36643,N_36988);
nor U37109 (N_37109,N_36786,N_36507);
nand U37110 (N_37110,N_36714,N_36817);
nand U37111 (N_37111,N_36751,N_36556);
and U37112 (N_37112,N_36968,N_36595);
and U37113 (N_37113,N_36565,N_36818);
nand U37114 (N_37114,N_36931,N_36795);
and U37115 (N_37115,N_36792,N_36811);
nor U37116 (N_37116,N_36938,N_36871);
nor U37117 (N_37117,N_36979,N_36680);
nor U37118 (N_37118,N_36543,N_36519);
or U37119 (N_37119,N_36660,N_36580);
nor U37120 (N_37120,N_36505,N_36829);
nor U37121 (N_37121,N_36566,N_36661);
xnor U37122 (N_37122,N_36813,N_36835);
nand U37123 (N_37123,N_36732,N_36709);
nand U37124 (N_37124,N_36577,N_36511);
nor U37125 (N_37125,N_36658,N_36770);
and U37126 (N_37126,N_36801,N_36978);
nand U37127 (N_37127,N_36683,N_36771);
nand U37128 (N_37128,N_36527,N_36909);
and U37129 (N_37129,N_36971,N_36695);
or U37130 (N_37130,N_36956,N_36523);
xor U37131 (N_37131,N_36905,N_36873);
xnor U37132 (N_37132,N_36525,N_36570);
and U37133 (N_37133,N_36539,N_36846);
and U37134 (N_37134,N_36895,N_36563);
nor U37135 (N_37135,N_36594,N_36589);
nand U37136 (N_37136,N_36963,N_36651);
xnor U37137 (N_37137,N_36593,N_36977);
and U37138 (N_37138,N_36728,N_36894);
or U37139 (N_37139,N_36610,N_36541);
or U37140 (N_37140,N_36902,N_36742);
and U37141 (N_37141,N_36609,N_36741);
nor U37142 (N_37142,N_36759,N_36921);
xnor U37143 (N_37143,N_36652,N_36842);
xor U37144 (N_37144,N_36914,N_36889);
nand U37145 (N_37145,N_36571,N_36746);
and U37146 (N_37146,N_36940,N_36962);
xnor U37147 (N_37147,N_36560,N_36997);
or U37148 (N_37148,N_36650,N_36816);
and U37149 (N_37149,N_36558,N_36888);
nor U37150 (N_37150,N_36913,N_36987);
xnor U37151 (N_37151,N_36826,N_36611);
nor U37152 (N_37152,N_36878,N_36534);
or U37153 (N_37153,N_36596,N_36715);
or U37154 (N_37154,N_36853,N_36559);
and U37155 (N_37155,N_36900,N_36863);
or U37156 (N_37156,N_36948,N_36898);
xnor U37157 (N_37157,N_36743,N_36897);
or U37158 (N_37158,N_36845,N_36964);
nand U37159 (N_37159,N_36729,N_36791);
nand U37160 (N_37160,N_36830,N_36930);
and U37161 (N_37161,N_36656,N_36825);
xor U37162 (N_37162,N_36872,N_36983);
and U37163 (N_37163,N_36972,N_36992);
xor U37164 (N_37164,N_36689,N_36855);
nand U37165 (N_37165,N_36679,N_36703);
and U37166 (N_37166,N_36649,N_36554);
and U37167 (N_37167,N_36629,N_36951);
or U37168 (N_37168,N_36508,N_36922);
and U37169 (N_37169,N_36712,N_36837);
and U37170 (N_37170,N_36942,N_36550);
or U37171 (N_37171,N_36980,N_36701);
xor U37172 (N_37172,N_36799,N_36947);
nor U37173 (N_37173,N_36713,N_36669);
nor U37174 (N_37174,N_36887,N_36725);
or U37175 (N_37175,N_36757,N_36776);
nor U37176 (N_37176,N_36739,N_36819);
and U37177 (N_37177,N_36950,N_36613);
nand U37178 (N_37178,N_36615,N_36904);
xnor U37179 (N_37179,N_36545,N_36557);
nand U37180 (N_37180,N_36533,N_36882);
nand U37181 (N_37181,N_36521,N_36744);
nand U37182 (N_37182,N_36907,N_36572);
nand U37183 (N_37183,N_36733,N_36995);
and U37184 (N_37184,N_36981,N_36634);
and U37185 (N_37185,N_36700,N_36804);
or U37186 (N_37186,N_36923,N_36916);
nor U37187 (N_37187,N_36885,N_36717);
or U37188 (N_37188,N_36645,N_36690);
nand U37189 (N_37189,N_36544,N_36939);
nand U37190 (N_37190,N_36718,N_36737);
or U37191 (N_37191,N_36862,N_36604);
nor U37192 (N_37192,N_36945,N_36785);
nand U37193 (N_37193,N_36638,N_36529);
or U37194 (N_37194,N_36512,N_36562);
xor U37195 (N_37195,N_36935,N_36625);
nand U37196 (N_37196,N_36807,N_36970);
xnor U37197 (N_37197,N_36555,N_36864);
xnor U37198 (N_37198,N_36874,N_36908);
and U37199 (N_37199,N_36881,N_36699);
nand U37200 (N_37200,N_36763,N_36518);
nand U37201 (N_37201,N_36708,N_36684);
nand U37202 (N_37202,N_36513,N_36653);
xor U37203 (N_37203,N_36667,N_36925);
nor U37204 (N_37204,N_36839,N_36955);
xor U37205 (N_37205,N_36857,N_36840);
and U37206 (N_37206,N_36686,N_36503);
and U37207 (N_37207,N_36627,N_36765);
nor U37208 (N_37208,N_36607,N_36965);
and U37209 (N_37209,N_36621,N_36581);
or U37210 (N_37210,N_36841,N_36564);
nand U37211 (N_37211,N_36608,N_36827);
or U37212 (N_37212,N_36969,N_36726);
and U37213 (N_37213,N_36941,N_36654);
or U37214 (N_37214,N_36814,N_36974);
xnor U37215 (N_37215,N_36514,N_36721);
or U37216 (N_37216,N_36752,N_36989);
and U37217 (N_37217,N_36749,N_36868);
nand U37218 (N_37218,N_36869,N_36996);
or U37219 (N_37219,N_36966,N_36784);
nand U37220 (N_37220,N_36573,N_36976);
xor U37221 (N_37221,N_36821,N_36618);
and U37222 (N_37222,N_36585,N_36662);
and U37223 (N_37223,N_36838,N_36673);
nor U37224 (N_37224,N_36836,N_36522);
or U37225 (N_37225,N_36628,N_36802);
xor U37226 (N_37226,N_36957,N_36588);
or U37227 (N_37227,N_36696,N_36929);
nor U37228 (N_37228,N_36880,N_36810);
and U37229 (N_37229,N_36982,N_36990);
xor U37230 (N_37230,N_36722,N_36668);
nand U37231 (N_37231,N_36670,N_36926);
xnor U37232 (N_37232,N_36682,N_36832);
or U37233 (N_37233,N_36711,N_36877);
nor U37234 (N_37234,N_36777,N_36664);
or U37235 (N_37235,N_36833,N_36626);
nand U37236 (N_37236,N_36624,N_36685);
and U37237 (N_37237,N_36899,N_36710);
nor U37238 (N_37238,N_36890,N_36704);
nor U37239 (N_37239,N_36999,N_36756);
and U37240 (N_37240,N_36967,N_36600);
and U37241 (N_37241,N_36910,N_36548);
xnor U37242 (N_37242,N_36606,N_36569);
nor U37243 (N_37243,N_36671,N_36936);
and U37244 (N_37244,N_36716,N_36693);
nand U37245 (N_37245,N_36831,N_36860);
nor U37246 (N_37246,N_36809,N_36944);
and U37247 (N_37247,N_36536,N_36553);
nor U37248 (N_37248,N_36663,N_36740);
nor U37249 (N_37249,N_36911,N_36883);
nor U37250 (N_37250,N_36612,N_36622);
or U37251 (N_37251,N_36940,N_36873);
and U37252 (N_37252,N_36533,N_36997);
xor U37253 (N_37253,N_36578,N_36793);
and U37254 (N_37254,N_36706,N_36816);
nor U37255 (N_37255,N_36794,N_36716);
nand U37256 (N_37256,N_36986,N_36717);
or U37257 (N_37257,N_36599,N_36724);
nand U37258 (N_37258,N_36892,N_36968);
nand U37259 (N_37259,N_36709,N_36701);
nor U37260 (N_37260,N_36750,N_36988);
xor U37261 (N_37261,N_36854,N_36509);
xnor U37262 (N_37262,N_36750,N_36518);
xor U37263 (N_37263,N_36878,N_36791);
nand U37264 (N_37264,N_36871,N_36773);
and U37265 (N_37265,N_36571,N_36588);
and U37266 (N_37266,N_36501,N_36920);
or U37267 (N_37267,N_36784,N_36622);
nor U37268 (N_37268,N_36751,N_36996);
nor U37269 (N_37269,N_36777,N_36868);
or U37270 (N_37270,N_36826,N_36773);
nand U37271 (N_37271,N_36603,N_36646);
or U37272 (N_37272,N_36749,N_36801);
nand U37273 (N_37273,N_36747,N_36834);
nor U37274 (N_37274,N_36579,N_36584);
or U37275 (N_37275,N_36678,N_36863);
nor U37276 (N_37276,N_36750,N_36911);
nor U37277 (N_37277,N_36500,N_36522);
and U37278 (N_37278,N_36743,N_36831);
nand U37279 (N_37279,N_36827,N_36651);
and U37280 (N_37280,N_36929,N_36612);
nand U37281 (N_37281,N_36806,N_36935);
nand U37282 (N_37282,N_36845,N_36808);
or U37283 (N_37283,N_36515,N_36986);
or U37284 (N_37284,N_36593,N_36919);
nand U37285 (N_37285,N_36735,N_36719);
xnor U37286 (N_37286,N_36809,N_36862);
and U37287 (N_37287,N_36724,N_36980);
xnor U37288 (N_37288,N_36540,N_36960);
nand U37289 (N_37289,N_36966,N_36884);
and U37290 (N_37290,N_36970,N_36727);
xnor U37291 (N_37291,N_36732,N_36917);
xnor U37292 (N_37292,N_36730,N_36746);
nor U37293 (N_37293,N_36804,N_36984);
nor U37294 (N_37294,N_36882,N_36830);
nand U37295 (N_37295,N_36878,N_36662);
nor U37296 (N_37296,N_36822,N_36664);
nand U37297 (N_37297,N_36684,N_36980);
or U37298 (N_37298,N_36554,N_36943);
nor U37299 (N_37299,N_36871,N_36550);
nor U37300 (N_37300,N_36655,N_36502);
nand U37301 (N_37301,N_36821,N_36880);
xnor U37302 (N_37302,N_36745,N_36651);
xor U37303 (N_37303,N_36690,N_36615);
or U37304 (N_37304,N_36639,N_36776);
or U37305 (N_37305,N_36974,N_36868);
or U37306 (N_37306,N_36610,N_36741);
and U37307 (N_37307,N_36533,N_36632);
nand U37308 (N_37308,N_36752,N_36544);
nor U37309 (N_37309,N_36522,N_36774);
xnor U37310 (N_37310,N_36913,N_36962);
and U37311 (N_37311,N_36558,N_36791);
nor U37312 (N_37312,N_36785,N_36534);
nor U37313 (N_37313,N_36906,N_36577);
xor U37314 (N_37314,N_36708,N_36592);
nand U37315 (N_37315,N_36581,N_36750);
nor U37316 (N_37316,N_36707,N_36518);
or U37317 (N_37317,N_36915,N_36653);
or U37318 (N_37318,N_36647,N_36512);
xnor U37319 (N_37319,N_36557,N_36731);
xnor U37320 (N_37320,N_36984,N_36693);
nor U37321 (N_37321,N_36882,N_36647);
nor U37322 (N_37322,N_36684,N_36531);
and U37323 (N_37323,N_36796,N_36772);
nand U37324 (N_37324,N_36905,N_36651);
nor U37325 (N_37325,N_36502,N_36557);
xor U37326 (N_37326,N_36706,N_36741);
nand U37327 (N_37327,N_36712,N_36667);
or U37328 (N_37328,N_36733,N_36636);
nand U37329 (N_37329,N_36689,N_36813);
and U37330 (N_37330,N_36511,N_36916);
nor U37331 (N_37331,N_36765,N_36921);
nor U37332 (N_37332,N_36931,N_36634);
nor U37333 (N_37333,N_36645,N_36758);
nand U37334 (N_37334,N_36834,N_36820);
nor U37335 (N_37335,N_36944,N_36512);
nor U37336 (N_37336,N_36537,N_36647);
and U37337 (N_37337,N_36962,N_36983);
nor U37338 (N_37338,N_36680,N_36748);
and U37339 (N_37339,N_36996,N_36638);
xor U37340 (N_37340,N_36965,N_36774);
nor U37341 (N_37341,N_36609,N_36765);
nor U37342 (N_37342,N_36872,N_36584);
or U37343 (N_37343,N_36846,N_36914);
and U37344 (N_37344,N_36929,N_36930);
and U37345 (N_37345,N_36506,N_36597);
nand U37346 (N_37346,N_36726,N_36545);
or U37347 (N_37347,N_36572,N_36613);
xnor U37348 (N_37348,N_36529,N_36893);
or U37349 (N_37349,N_36888,N_36703);
nand U37350 (N_37350,N_36710,N_36663);
nor U37351 (N_37351,N_36919,N_36500);
xnor U37352 (N_37352,N_36805,N_36693);
nor U37353 (N_37353,N_36538,N_36924);
and U37354 (N_37354,N_36670,N_36970);
xnor U37355 (N_37355,N_36938,N_36537);
xnor U37356 (N_37356,N_36658,N_36598);
and U37357 (N_37357,N_36677,N_36507);
nand U37358 (N_37358,N_36645,N_36829);
nor U37359 (N_37359,N_36802,N_36801);
or U37360 (N_37360,N_36853,N_36998);
nor U37361 (N_37361,N_36785,N_36914);
and U37362 (N_37362,N_36842,N_36944);
xnor U37363 (N_37363,N_36924,N_36954);
nor U37364 (N_37364,N_36769,N_36661);
nor U37365 (N_37365,N_36888,N_36730);
xor U37366 (N_37366,N_36928,N_36670);
and U37367 (N_37367,N_36860,N_36798);
and U37368 (N_37368,N_36889,N_36888);
and U37369 (N_37369,N_36960,N_36618);
xnor U37370 (N_37370,N_36941,N_36630);
nand U37371 (N_37371,N_36974,N_36574);
xnor U37372 (N_37372,N_36540,N_36541);
nor U37373 (N_37373,N_36699,N_36508);
nand U37374 (N_37374,N_36811,N_36513);
and U37375 (N_37375,N_36573,N_36774);
xor U37376 (N_37376,N_36987,N_36585);
or U37377 (N_37377,N_36580,N_36847);
xnor U37378 (N_37378,N_36895,N_36529);
and U37379 (N_37379,N_36927,N_36867);
xor U37380 (N_37380,N_36953,N_36788);
or U37381 (N_37381,N_36815,N_36930);
or U37382 (N_37382,N_36803,N_36793);
nor U37383 (N_37383,N_36943,N_36882);
nand U37384 (N_37384,N_36787,N_36514);
nand U37385 (N_37385,N_36581,N_36993);
nor U37386 (N_37386,N_36887,N_36527);
or U37387 (N_37387,N_36858,N_36631);
and U37388 (N_37388,N_36670,N_36816);
or U37389 (N_37389,N_36819,N_36686);
nand U37390 (N_37390,N_36887,N_36776);
and U37391 (N_37391,N_36632,N_36774);
nor U37392 (N_37392,N_36516,N_36840);
nor U37393 (N_37393,N_36929,N_36699);
nor U37394 (N_37394,N_36695,N_36990);
nor U37395 (N_37395,N_36947,N_36923);
or U37396 (N_37396,N_36960,N_36903);
and U37397 (N_37397,N_36652,N_36833);
and U37398 (N_37398,N_36691,N_36670);
nand U37399 (N_37399,N_36737,N_36547);
or U37400 (N_37400,N_36759,N_36901);
or U37401 (N_37401,N_36831,N_36760);
nand U37402 (N_37402,N_36615,N_36945);
or U37403 (N_37403,N_36897,N_36956);
xnor U37404 (N_37404,N_36674,N_36623);
xor U37405 (N_37405,N_36691,N_36998);
xnor U37406 (N_37406,N_36600,N_36739);
or U37407 (N_37407,N_36778,N_36518);
xnor U37408 (N_37408,N_36779,N_36604);
xnor U37409 (N_37409,N_36804,N_36725);
or U37410 (N_37410,N_36987,N_36948);
nor U37411 (N_37411,N_36553,N_36976);
nand U37412 (N_37412,N_36969,N_36572);
xor U37413 (N_37413,N_36763,N_36822);
nor U37414 (N_37414,N_36770,N_36996);
xnor U37415 (N_37415,N_36683,N_36982);
and U37416 (N_37416,N_36589,N_36997);
and U37417 (N_37417,N_36906,N_36561);
nand U37418 (N_37418,N_36559,N_36633);
and U37419 (N_37419,N_36966,N_36747);
nand U37420 (N_37420,N_36568,N_36525);
or U37421 (N_37421,N_36938,N_36822);
nand U37422 (N_37422,N_36717,N_36932);
nor U37423 (N_37423,N_36875,N_36771);
xor U37424 (N_37424,N_36814,N_36978);
or U37425 (N_37425,N_36641,N_36930);
and U37426 (N_37426,N_36519,N_36637);
xor U37427 (N_37427,N_36631,N_36577);
and U37428 (N_37428,N_36674,N_36540);
nor U37429 (N_37429,N_36879,N_36877);
and U37430 (N_37430,N_36893,N_36595);
nand U37431 (N_37431,N_36564,N_36983);
or U37432 (N_37432,N_36823,N_36682);
xor U37433 (N_37433,N_36603,N_36915);
nand U37434 (N_37434,N_36663,N_36845);
and U37435 (N_37435,N_36883,N_36844);
nand U37436 (N_37436,N_36612,N_36589);
nor U37437 (N_37437,N_36553,N_36834);
nand U37438 (N_37438,N_36782,N_36649);
or U37439 (N_37439,N_36820,N_36730);
nand U37440 (N_37440,N_36753,N_36801);
xnor U37441 (N_37441,N_36763,N_36701);
nor U37442 (N_37442,N_36878,N_36757);
nand U37443 (N_37443,N_36932,N_36884);
or U37444 (N_37444,N_36656,N_36815);
nand U37445 (N_37445,N_36915,N_36849);
xnor U37446 (N_37446,N_36870,N_36995);
xnor U37447 (N_37447,N_36956,N_36838);
nor U37448 (N_37448,N_36754,N_36827);
nor U37449 (N_37449,N_36688,N_36726);
nor U37450 (N_37450,N_36555,N_36546);
nand U37451 (N_37451,N_36838,N_36965);
nand U37452 (N_37452,N_36509,N_36630);
or U37453 (N_37453,N_36910,N_36947);
xor U37454 (N_37454,N_36698,N_36820);
nand U37455 (N_37455,N_36809,N_36563);
nor U37456 (N_37456,N_36917,N_36638);
or U37457 (N_37457,N_36748,N_36535);
nor U37458 (N_37458,N_36506,N_36626);
xnor U37459 (N_37459,N_36872,N_36868);
and U37460 (N_37460,N_36768,N_36677);
nor U37461 (N_37461,N_36792,N_36609);
nor U37462 (N_37462,N_36764,N_36724);
nand U37463 (N_37463,N_36888,N_36603);
nand U37464 (N_37464,N_36964,N_36941);
and U37465 (N_37465,N_36805,N_36600);
xor U37466 (N_37466,N_36791,N_36892);
xor U37467 (N_37467,N_36851,N_36768);
xor U37468 (N_37468,N_36798,N_36774);
and U37469 (N_37469,N_36949,N_36726);
nand U37470 (N_37470,N_36964,N_36895);
nand U37471 (N_37471,N_36509,N_36825);
and U37472 (N_37472,N_36793,N_36521);
xor U37473 (N_37473,N_36650,N_36883);
or U37474 (N_37474,N_36757,N_36753);
nor U37475 (N_37475,N_36525,N_36730);
xor U37476 (N_37476,N_36569,N_36726);
and U37477 (N_37477,N_36831,N_36711);
xor U37478 (N_37478,N_36893,N_36778);
or U37479 (N_37479,N_36923,N_36535);
and U37480 (N_37480,N_36659,N_36777);
and U37481 (N_37481,N_36896,N_36991);
or U37482 (N_37482,N_36847,N_36577);
nor U37483 (N_37483,N_36807,N_36765);
xor U37484 (N_37484,N_36690,N_36619);
nor U37485 (N_37485,N_36521,N_36895);
or U37486 (N_37486,N_36680,N_36805);
xnor U37487 (N_37487,N_36943,N_36762);
and U37488 (N_37488,N_36867,N_36898);
nand U37489 (N_37489,N_36668,N_36628);
nor U37490 (N_37490,N_36706,N_36523);
xor U37491 (N_37491,N_36875,N_36946);
nor U37492 (N_37492,N_36724,N_36648);
nand U37493 (N_37493,N_36558,N_36713);
and U37494 (N_37494,N_36902,N_36890);
xor U37495 (N_37495,N_36942,N_36552);
and U37496 (N_37496,N_36786,N_36804);
xor U37497 (N_37497,N_36870,N_36966);
xor U37498 (N_37498,N_36835,N_36691);
and U37499 (N_37499,N_36751,N_36960);
and U37500 (N_37500,N_37434,N_37213);
xnor U37501 (N_37501,N_37001,N_37087);
nand U37502 (N_37502,N_37490,N_37225);
nand U37503 (N_37503,N_37493,N_37277);
xnor U37504 (N_37504,N_37004,N_37359);
nor U37505 (N_37505,N_37370,N_37125);
xor U37506 (N_37506,N_37283,N_37405);
or U37507 (N_37507,N_37058,N_37440);
or U37508 (N_37508,N_37026,N_37298);
nor U37509 (N_37509,N_37089,N_37293);
nor U37510 (N_37510,N_37074,N_37211);
or U37511 (N_37511,N_37236,N_37468);
nand U37512 (N_37512,N_37237,N_37472);
nand U37513 (N_37513,N_37176,N_37034);
nor U37514 (N_37514,N_37343,N_37301);
nand U37515 (N_37515,N_37425,N_37429);
nand U37516 (N_37516,N_37047,N_37287);
nand U37517 (N_37517,N_37349,N_37061);
nor U37518 (N_37518,N_37157,N_37187);
xnor U37519 (N_37519,N_37380,N_37284);
nor U37520 (N_37520,N_37107,N_37188);
nor U37521 (N_37521,N_37180,N_37375);
nor U37522 (N_37522,N_37433,N_37110);
xor U37523 (N_37523,N_37379,N_37009);
and U37524 (N_37524,N_37390,N_37413);
and U37525 (N_37525,N_37141,N_37191);
and U37526 (N_37526,N_37338,N_37383);
nand U37527 (N_37527,N_37443,N_37309);
or U37528 (N_37528,N_37171,N_37106);
or U37529 (N_37529,N_37037,N_37060);
nand U37530 (N_37530,N_37145,N_37486);
nand U37531 (N_37531,N_37360,N_37482);
xor U37532 (N_37532,N_37163,N_37403);
and U37533 (N_37533,N_37203,N_37181);
nor U37534 (N_37534,N_37054,N_37240);
nor U37535 (N_37535,N_37109,N_37018);
nand U37536 (N_37536,N_37400,N_37066);
nand U37537 (N_37537,N_37445,N_37049);
nor U37538 (N_37538,N_37111,N_37068);
or U37539 (N_37539,N_37408,N_37005);
nand U37540 (N_37540,N_37175,N_37285);
xor U37541 (N_37541,N_37139,N_37029);
xor U37542 (N_37542,N_37358,N_37488);
xor U37543 (N_37543,N_37348,N_37315);
or U37544 (N_37544,N_37094,N_37173);
nand U37545 (N_37545,N_37270,N_37202);
and U37546 (N_37546,N_37323,N_37392);
nor U37547 (N_37547,N_37248,N_37069);
nand U37548 (N_37548,N_37122,N_37159);
or U37549 (N_37549,N_37102,N_37414);
nand U37550 (N_37550,N_37388,N_37340);
or U37551 (N_37551,N_37124,N_37337);
and U37552 (N_37552,N_37281,N_37346);
xor U37553 (N_37553,N_37432,N_37489);
and U37554 (N_37554,N_37333,N_37010);
nand U37555 (N_37555,N_37291,N_37178);
or U37556 (N_37556,N_37154,N_37117);
nor U37557 (N_37557,N_37256,N_37057);
or U37558 (N_37558,N_37144,N_37072);
xor U37559 (N_37559,N_37282,N_37326);
nor U37560 (N_37560,N_37342,N_37231);
and U37561 (N_37561,N_37210,N_37377);
and U37562 (N_37562,N_37165,N_37243);
and U37563 (N_37563,N_37098,N_37394);
xnor U37564 (N_37564,N_37267,N_37115);
and U37565 (N_37565,N_37067,N_37322);
or U37566 (N_37566,N_37196,N_37321);
nor U37567 (N_37567,N_37142,N_37039);
nor U37568 (N_37568,N_37456,N_37201);
nor U37569 (N_37569,N_37242,N_37347);
nor U37570 (N_37570,N_37214,N_37156);
nor U37571 (N_37571,N_37480,N_37297);
xor U37572 (N_37572,N_37169,N_37369);
or U37573 (N_37573,N_37431,N_37090);
or U37574 (N_37574,N_37132,N_37320);
nand U37575 (N_37575,N_37193,N_37352);
and U37576 (N_37576,N_37198,N_37485);
or U37577 (N_37577,N_37452,N_37395);
nand U37578 (N_37578,N_37081,N_37378);
nor U37579 (N_37579,N_37092,N_37263);
and U37580 (N_37580,N_37454,N_37366);
or U37581 (N_37581,N_37462,N_37186);
and U37582 (N_37582,N_37120,N_37216);
or U37583 (N_37583,N_37444,N_37200);
xnor U37584 (N_37584,N_37238,N_37085);
nand U37585 (N_37585,N_37177,N_37424);
and U37586 (N_37586,N_37224,N_37114);
xnor U37587 (N_37587,N_37208,N_37170);
nand U37588 (N_37588,N_37253,N_37276);
and U37589 (N_37589,N_37062,N_37324);
xnor U37590 (N_37590,N_37172,N_37179);
nor U37591 (N_37591,N_37127,N_37404);
and U37592 (N_37592,N_37077,N_37084);
or U37593 (N_37593,N_37467,N_37149);
nand U37594 (N_37594,N_37271,N_37008);
nor U37595 (N_37595,N_37487,N_37461);
nand U37596 (N_37596,N_37044,N_37006);
xnor U37597 (N_37597,N_37002,N_37212);
or U37598 (N_37598,N_37235,N_37205);
xor U37599 (N_37599,N_37406,N_37448);
xnor U37600 (N_37600,N_37146,N_37464);
or U37601 (N_37601,N_37295,N_37450);
or U37602 (N_37602,N_37476,N_37245);
xnor U37603 (N_37603,N_37209,N_37020);
nor U37604 (N_37604,N_37442,N_37244);
nand U37605 (N_37605,N_37116,N_37079);
or U37606 (N_37606,N_37460,N_37415);
nor U37607 (N_37607,N_37318,N_37335);
xor U37608 (N_37608,N_37112,N_37356);
nor U37609 (N_37609,N_37185,N_37416);
xnor U37610 (N_37610,N_37140,N_37331);
nor U37611 (N_37611,N_37304,N_37045);
or U37612 (N_37612,N_37022,N_37308);
or U37613 (N_37613,N_37289,N_37466);
and U37614 (N_37614,N_37484,N_37030);
nand U37615 (N_37615,N_37025,N_37232);
xor U37616 (N_37616,N_37426,N_37036);
xnor U37617 (N_37617,N_37332,N_37311);
or U37618 (N_37618,N_37357,N_37477);
nor U37619 (N_37619,N_37459,N_37143);
xnor U37620 (N_37620,N_37217,N_37437);
and U37621 (N_37621,N_37470,N_37128);
or U37622 (N_37622,N_37197,N_37218);
xor U37623 (N_37623,N_37327,N_37409);
xnor U37624 (N_37624,N_37272,N_37003);
or U37625 (N_37625,N_37451,N_37166);
and U37626 (N_37626,N_37381,N_37474);
and U37627 (N_37627,N_37126,N_37103);
nor U37628 (N_37628,N_37307,N_37292);
xor U37629 (N_37629,N_37252,N_37155);
or U37630 (N_37630,N_37104,N_37136);
and U37631 (N_37631,N_37481,N_37046);
or U37632 (N_37632,N_37420,N_37150);
and U37633 (N_37633,N_37266,N_37078);
xor U37634 (N_37634,N_37056,N_37478);
nor U37635 (N_37635,N_37391,N_37041);
or U37636 (N_37636,N_37093,N_37096);
nor U37637 (N_37637,N_37019,N_37334);
and U37638 (N_37638,N_37279,N_37250);
nor U37639 (N_37639,N_37365,N_37354);
and U37640 (N_37640,N_37449,N_37241);
nor U37641 (N_37641,N_37167,N_37024);
nor U37642 (N_37642,N_37280,N_37399);
nand U37643 (N_37643,N_37016,N_37296);
or U37644 (N_37644,N_37227,N_37479);
nand U37645 (N_37645,N_37251,N_37255);
and U37646 (N_37646,N_37097,N_37230);
or U37647 (N_37647,N_37147,N_37286);
nand U37648 (N_37648,N_37043,N_37491);
nor U37649 (N_37649,N_37402,N_37469);
nor U37650 (N_37650,N_37364,N_37164);
nand U37651 (N_37651,N_37457,N_37325);
and U37652 (N_37652,N_37032,N_37133);
nor U37653 (N_37653,N_37316,N_37435);
and U37654 (N_37654,N_37088,N_37421);
or U37655 (N_37655,N_37300,N_37330);
or U37656 (N_37656,N_37397,N_37418);
and U37657 (N_37657,N_37494,N_37317);
and U37658 (N_37658,N_37288,N_37401);
xnor U37659 (N_37659,N_37053,N_37119);
nor U37660 (N_37660,N_37278,N_37073);
nand U37661 (N_37661,N_37314,N_37389);
nor U37662 (N_37662,N_37492,N_37051);
xnor U37663 (N_37663,N_37247,N_37310);
xor U37664 (N_37664,N_37372,N_37436);
nand U37665 (N_37665,N_37190,N_37151);
nor U37666 (N_37666,N_37312,N_37294);
nor U37667 (N_37667,N_37222,N_37194);
and U37668 (N_37668,N_37229,N_37427);
nor U37669 (N_37669,N_37455,N_37302);
nor U37670 (N_37670,N_37361,N_37233);
or U37671 (N_37671,N_37135,N_37367);
or U37672 (N_37672,N_37148,N_37123);
nor U37673 (N_37673,N_37430,N_37386);
nor U37674 (N_37674,N_37138,N_37371);
xnor U37675 (N_37675,N_37076,N_37385);
nor U37676 (N_37676,N_37265,N_37031);
nand U37677 (N_37677,N_37261,N_37207);
or U37678 (N_37678,N_37257,N_37258);
nand U37679 (N_37679,N_37355,N_37070);
and U37680 (N_37680,N_37319,N_37017);
or U37681 (N_37681,N_37306,N_37189);
nand U37682 (N_37682,N_37055,N_37059);
nand U37683 (N_37683,N_37095,N_37410);
and U37684 (N_37684,N_37384,N_37174);
xnor U37685 (N_37685,N_37422,N_37458);
nor U37686 (N_37686,N_37262,N_37099);
nand U37687 (N_37687,N_37345,N_37083);
and U37688 (N_37688,N_37038,N_37075);
nor U37689 (N_37689,N_37428,N_37042);
and U37690 (N_37690,N_37259,N_37105);
nand U37691 (N_37691,N_37160,N_37368);
and U37692 (N_37692,N_37091,N_37152);
or U37693 (N_37693,N_37305,N_37274);
and U37694 (N_37694,N_37108,N_37353);
nand U37695 (N_37695,N_37086,N_37260);
or U37696 (N_37696,N_37204,N_37411);
nand U37697 (N_37697,N_37007,N_37161);
xnor U37698 (N_37698,N_37407,N_37249);
xnor U37699 (N_37699,N_37439,N_37064);
or U37700 (N_37700,N_37195,N_37234);
xor U37701 (N_37701,N_37336,N_37021);
and U37702 (N_37702,N_37027,N_37351);
or U37703 (N_37703,N_37273,N_37498);
xor U37704 (N_37704,N_37033,N_37275);
nor U37705 (N_37705,N_37373,N_37254);
xor U37706 (N_37706,N_37417,N_37438);
xor U37707 (N_37707,N_37313,N_37184);
and U37708 (N_37708,N_37495,N_37130);
xnor U37709 (N_37709,N_37499,N_37446);
nand U37710 (N_37710,N_37050,N_37339);
nor U37711 (N_37711,N_37215,N_37040);
nand U37712 (N_37712,N_37463,N_37035);
nand U37713 (N_37713,N_37192,N_37412);
and U37714 (N_37714,N_37113,N_37471);
xor U37715 (N_37715,N_37228,N_37023);
nor U37716 (N_37716,N_37129,N_37264);
or U37717 (N_37717,N_37246,N_37419);
xnor U37718 (N_37718,N_37221,N_37137);
nand U37719 (N_37719,N_37220,N_37475);
or U37720 (N_37720,N_37269,N_37206);
or U37721 (N_37721,N_37447,N_37441);
nand U37722 (N_37722,N_37153,N_37219);
and U37723 (N_37723,N_37329,N_37028);
nor U37724 (N_37724,N_37423,N_37239);
and U37725 (N_37725,N_37393,N_37268);
nand U37726 (N_37726,N_37013,N_37134);
and U37727 (N_37727,N_37226,N_37071);
or U37728 (N_37728,N_37344,N_37496);
and U37729 (N_37729,N_37374,N_37118);
and U37730 (N_37730,N_37299,N_37082);
nand U37731 (N_37731,N_37453,N_37168);
or U37732 (N_37732,N_37328,N_37015);
nor U37733 (N_37733,N_37080,N_37101);
nor U37734 (N_37734,N_37000,N_37131);
or U37735 (N_37735,N_37473,N_37398);
and U37736 (N_37736,N_37065,N_37063);
nor U37737 (N_37737,N_37363,N_37158);
nand U37738 (N_37738,N_37290,N_37183);
nor U37739 (N_37739,N_37048,N_37350);
xnor U37740 (N_37740,N_37465,N_37223);
nand U37741 (N_37741,N_37396,N_37362);
xor U37742 (N_37742,N_37199,N_37303);
nor U37743 (N_37743,N_37162,N_37012);
or U37744 (N_37744,N_37121,N_37341);
xor U37745 (N_37745,N_37387,N_37382);
or U37746 (N_37746,N_37182,N_37497);
nor U37747 (N_37747,N_37014,N_37100);
nor U37748 (N_37748,N_37052,N_37483);
or U37749 (N_37749,N_37011,N_37376);
nand U37750 (N_37750,N_37055,N_37039);
nor U37751 (N_37751,N_37035,N_37106);
or U37752 (N_37752,N_37455,N_37038);
or U37753 (N_37753,N_37461,N_37232);
and U37754 (N_37754,N_37144,N_37099);
or U37755 (N_37755,N_37492,N_37011);
nor U37756 (N_37756,N_37278,N_37372);
or U37757 (N_37757,N_37190,N_37460);
xor U37758 (N_37758,N_37050,N_37085);
or U37759 (N_37759,N_37044,N_37406);
nor U37760 (N_37760,N_37018,N_37088);
nand U37761 (N_37761,N_37193,N_37125);
nor U37762 (N_37762,N_37472,N_37184);
nand U37763 (N_37763,N_37013,N_37299);
nor U37764 (N_37764,N_37151,N_37349);
nor U37765 (N_37765,N_37224,N_37437);
or U37766 (N_37766,N_37227,N_37268);
or U37767 (N_37767,N_37372,N_37169);
nand U37768 (N_37768,N_37364,N_37352);
xnor U37769 (N_37769,N_37330,N_37206);
or U37770 (N_37770,N_37443,N_37043);
xnor U37771 (N_37771,N_37461,N_37331);
and U37772 (N_37772,N_37216,N_37428);
or U37773 (N_37773,N_37321,N_37392);
xnor U37774 (N_37774,N_37114,N_37135);
nor U37775 (N_37775,N_37149,N_37239);
or U37776 (N_37776,N_37483,N_37401);
xor U37777 (N_37777,N_37148,N_37239);
nand U37778 (N_37778,N_37324,N_37433);
nand U37779 (N_37779,N_37279,N_37337);
xor U37780 (N_37780,N_37262,N_37158);
nand U37781 (N_37781,N_37198,N_37441);
nand U37782 (N_37782,N_37376,N_37209);
nor U37783 (N_37783,N_37480,N_37002);
or U37784 (N_37784,N_37258,N_37390);
nand U37785 (N_37785,N_37426,N_37337);
nand U37786 (N_37786,N_37228,N_37284);
nand U37787 (N_37787,N_37216,N_37458);
xnor U37788 (N_37788,N_37075,N_37224);
nand U37789 (N_37789,N_37101,N_37146);
xnor U37790 (N_37790,N_37279,N_37393);
or U37791 (N_37791,N_37103,N_37426);
and U37792 (N_37792,N_37253,N_37440);
and U37793 (N_37793,N_37219,N_37328);
or U37794 (N_37794,N_37114,N_37427);
and U37795 (N_37795,N_37272,N_37141);
nand U37796 (N_37796,N_37355,N_37094);
or U37797 (N_37797,N_37065,N_37376);
and U37798 (N_37798,N_37064,N_37161);
xor U37799 (N_37799,N_37097,N_37126);
and U37800 (N_37800,N_37348,N_37357);
or U37801 (N_37801,N_37249,N_37467);
nand U37802 (N_37802,N_37093,N_37318);
nand U37803 (N_37803,N_37229,N_37281);
or U37804 (N_37804,N_37014,N_37372);
and U37805 (N_37805,N_37179,N_37073);
or U37806 (N_37806,N_37352,N_37197);
xnor U37807 (N_37807,N_37442,N_37049);
nor U37808 (N_37808,N_37393,N_37245);
and U37809 (N_37809,N_37113,N_37212);
or U37810 (N_37810,N_37153,N_37430);
and U37811 (N_37811,N_37303,N_37220);
nor U37812 (N_37812,N_37460,N_37111);
and U37813 (N_37813,N_37225,N_37065);
and U37814 (N_37814,N_37166,N_37131);
nand U37815 (N_37815,N_37464,N_37099);
xnor U37816 (N_37816,N_37418,N_37469);
xor U37817 (N_37817,N_37084,N_37308);
xor U37818 (N_37818,N_37167,N_37453);
and U37819 (N_37819,N_37412,N_37181);
nor U37820 (N_37820,N_37267,N_37186);
xnor U37821 (N_37821,N_37225,N_37018);
nor U37822 (N_37822,N_37173,N_37310);
nand U37823 (N_37823,N_37441,N_37488);
xnor U37824 (N_37824,N_37397,N_37192);
and U37825 (N_37825,N_37214,N_37449);
xnor U37826 (N_37826,N_37475,N_37308);
and U37827 (N_37827,N_37143,N_37436);
xnor U37828 (N_37828,N_37338,N_37165);
nor U37829 (N_37829,N_37297,N_37121);
or U37830 (N_37830,N_37408,N_37350);
nand U37831 (N_37831,N_37134,N_37289);
xor U37832 (N_37832,N_37299,N_37284);
xor U37833 (N_37833,N_37491,N_37173);
xor U37834 (N_37834,N_37369,N_37349);
and U37835 (N_37835,N_37168,N_37005);
nand U37836 (N_37836,N_37146,N_37099);
and U37837 (N_37837,N_37075,N_37018);
xnor U37838 (N_37838,N_37218,N_37074);
and U37839 (N_37839,N_37354,N_37361);
xnor U37840 (N_37840,N_37326,N_37266);
xor U37841 (N_37841,N_37101,N_37250);
nand U37842 (N_37842,N_37043,N_37323);
or U37843 (N_37843,N_37043,N_37473);
nor U37844 (N_37844,N_37333,N_37132);
or U37845 (N_37845,N_37007,N_37475);
and U37846 (N_37846,N_37248,N_37348);
and U37847 (N_37847,N_37054,N_37384);
or U37848 (N_37848,N_37494,N_37159);
nand U37849 (N_37849,N_37393,N_37357);
nand U37850 (N_37850,N_37171,N_37300);
nor U37851 (N_37851,N_37015,N_37278);
nand U37852 (N_37852,N_37389,N_37352);
nor U37853 (N_37853,N_37064,N_37181);
or U37854 (N_37854,N_37174,N_37315);
or U37855 (N_37855,N_37185,N_37003);
or U37856 (N_37856,N_37455,N_37171);
xor U37857 (N_37857,N_37432,N_37174);
nand U37858 (N_37858,N_37325,N_37495);
nand U37859 (N_37859,N_37098,N_37241);
or U37860 (N_37860,N_37093,N_37079);
xor U37861 (N_37861,N_37398,N_37117);
or U37862 (N_37862,N_37189,N_37426);
xnor U37863 (N_37863,N_37443,N_37189);
nor U37864 (N_37864,N_37170,N_37452);
or U37865 (N_37865,N_37103,N_37313);
xor U37866 (N_37866,N_37330,N_37113);
nand U37867 (N_37867,N_37465,N_37441);
nand U37868 (N_37868,N_37451,N_37455);
nor U37869 (N_37869,N_37269,N_37418);
and U37870 (N_37870,N_37005,N_37391);
nand U37871 (N_37871,N_37012,N_37194);
nor U37872 (N_37872,N_37485,N_37074);
or U37873 (N_37873,N_37244,N_37301);
or U37874 (N_37874,N_37064,N_37398);
nor U37875 (N_37875,N_37306,N_37127);
and U37876 (N_37876,N_37105,N_37385);
and U37877 (N_37877,N_37456,N_37370);
xor U37878 (N_37878,N_37428,N_37126);
or U37879 (N_37879,N_37467,N_37177);
or U37880 (N_37880,N_37489,N_37009);
nor U37881 (N_37881,N_37198,N_37258);
and U37882 (N_37882,N_37127,N_37441);
nor U37883 (N_37883,N_37182,N_37026);
nand U37884 (N_37884,N_37029,N_37132);
or U37885 (N_37885,N_37264,N_37198);
nand U37886 (N_37886,N_37154,N_37342);
nor U37887 (N_37887,N_37208,N_37461);
nor U37888 (N_37888,N_37442,N_37341);
or U37889 (N_37889,N_37235,N_37001);
and U37890 (N_37890,N_37228,N_37003);
or U37891 (N_37891,N_37360,N_37325);
nand U37892 (N_37892,N_37208,N_37102);
and U37893 (N_37893,N_37191,N_37087);
nor U37894 (N_37894,N_37265,N_37012);
or U37895 (N_37895,N_37281,N_37300);
xor U37896 (N_37896,N_37462,N_37423);
and U37897 (N_37897,N_37377,N_37045);
or U37898 (N_37898,N_37455,N_37294);
xnor U37899 (N_37899,N_37011,N_37049);
nor U37900 (N_37900,N_37114,N_37325);
and U37901 (N_37901,N_37464,N_37119);
or U37902 (N_37902,N_37313,N_37166);
xor U37903 (N_37903,N_37128,N_37124);
nand U37904 (N_37904,N_37360,N_37182);
and U37905 (N_37905,N_37467,N_37138);
or U37906 (N_37906,N_37428,N_37259);
xor U37907 (N_37907,N_37486,N_37034);
xnor U37908 (N_37908,N_37344,N_37050);
nor U37909 (N_37909,N_37149,N_37368);
nand U37910 (N_37910,N_37443,N_37473);
and U37911 (N_37911,N_37420,N_37148);
or U37912 (N_37912,N_37425,N_37444);
and U37913 (N_37913,N_37162,N_37474);
nor U37914 (N_37914,N_37210,N_37477);
nor U37915 (N_37915,N_37484,N_37380);
or U37916 (N_37916,N_37081,N_37297);
xor U37917 (N_37917,N_37135,N_37153);
or U37918 (N_37918,N_37291,N_37411);
or U37919 (N_37919,N_37109,N_37016);
xnor U37920 (N_37920,N_37449,N_37325);
xor U37921 (N_37921,N_37043,N_37244);
or U37922 (N_37922,N_37231,N_37340);
nand U37923 (N_37923,N_37324,N_37424);
nand U37924 (N_37924,N_37189,N_37031);
nor U37925 (N_37925,N_37185,N_37447);
nand U37926 (N_37926,N_37361,N_37153);
and U37927 (N_37927,N_37274,N_37486);
nand U37928 (N_37928,N_37157,N_37015);
and U37929 (N_37929,N_37019,N_37435);
nor U37930 (N_37930,N_37177,N_37017);
and U37931 (N_37931,N_37053,N_37397);
or U37932 (N_37932,N_37347,N_37299);
or U37933 (N_37933,N_37315,N_37111);
or U37934 (N_37934,N_37224,N_37062);
xor U37935 (N_37935,N_37209,N_37123);
nand U37936 (N_37936,N_37275,N_37166);
xnor U37937 (N_37937,N_37103,N_37170);
nor U37938 (N_37938,N_37435,N_37437);
or U37939 (N_37939,N_37007,N_37097);
nand U37940 (N_37940,N_37230,N_37061);
nor U37941 (N_37941,N_37021,N_37242);
and U37942 (N_37942,N_37283,N_37436);
nand U37943 (N_37943,N_37412,N_37474);
xnor U37944 (N_37944,N_37408,N_37004);
nor U37945 (N_37945,N_37143,N_37077);
or U37946 (N_37946,N_37224,N_37315);
nand U37947 (N_37947,N_37079,N_37262);
or U37948 (N_37948,N_37167,N_37127);
xnor U37949 (N_37949,N_37280,N_37467);
nand U37950 (N_37950,N_37192,N_37349);
xnor U37951 (N_37951,N_37202,N_37241);
xor U37952 (N_37952,N_37135,N_37193);
nor U37953 (N_37953,N_37398,N_37320);
or U37954 (N_37954,N_37131,N_37160);
and U37955 (N_37955,N_37112,N_37373);
or U37956 (N_37956,N_37392,N_37248);
and U37957 (N_37957,N_37302,N_37385);
nand U37958 (N_37958,N_37065,N_37046);
nor U37959 (N_37959,N_37229,N_37382);
xor U37960 (N_37960,N_37355,N_37253);
and U37961 (N_37961,N_37470,N_37169);
and U37962 (N_37962,N_37445,N_37415);
or U37963 (N_37963,N_37072,N_37220);
and U37964 (N_37964,N_37199,N_37147);
xnor U37965 (N_37965,N_37104,N_37226);
nor U37966 (N_37966,N_37137,N_37167);
and U37967 (N_37967,N_37418,N_37005);
nand U37968 (N_37968,N_37114,N_37210);
xnor U37969 (N_37969,N_37330,N_37214);
nand U37970 (N_37970,N_37353,N_37477);
and U37971 (N_37971,N_37164,N_37205);
or U37972 (N_37972,N_37136,N_37484);
nand U37973 (N_37973,N_37148,N_37342);
and U37974 (N_37974,N_37475,N_37405);
or U37975 (N_37975,N_37342,N_37357);
xnor U37976 (N_37976,N_37284,N_37134);
and U37977 (N_37977,N_37481,N_37255);
and U37978 (N_37978,N_37355,N_37474);
or U37979 (N_37979,N_37246,N_37065);
nand U37980 (N_37980,N_37227,N_37259);
or U37981 (N_37981,N_37292,N_37237);
xor U37982 (N_37982,N_37325,N_37471);
or U37983 (N_37983,N_37009,N_37111);
xor U37984 (N_37984,N_37394,N_37160);
and U37985 (N_37985,N_37406,N_37120);
or U37986 (N_37986,N_37104,N_37377);
xor U37987 (N_37987,N_37466,N_37366);
or U37988 (N_37988,N_37080,N_37346);
or U37989 (N_37989,N_37495,N_37077);
and U37990 (N_37990,N_37055,N_37454);
nor U37991 (N_37991,N_37464,N_37426);
or U37992 (N_37992,N_37072,N_37104);
nand U37993 (N_37993,N_37081,N_37109);
nand U37994 (N_37994,N_37271,N_37468);
and U37995 (N_37995,N_37143,N_37138);
xor U37996 (N_37996,N_37059,N_37456);
nor U37997 (N_37997,N_37369,N_37461);
or U37998 (N_37998,N_37033,N_37366);
xor U37999 (N_37999,N_37153,N_37009);
and U38000 (N_38000,N_37949,N_37582);
nand U38001 (N_38001,N_37609,N_37667);
or U38002 (N_38002,N_37841,N_37966);
xnor U38003 (N_38003,N_37770,N_37517);
xnor U38004 (N_38004,N_37734,N_37871);
or U38005 (N_38005,N_37781,N_37808);
nand U38006 (N_38006,N_37501,N_37595);
and U38007 (N_38007,N_37535,N_37544);
xor U38008 (N_38008,N_37826,N_37888);
nand U38009 (N_38009,N_37942,N_37668);
xnor U38010 (N_38010,N_37862,N_37747);
and U38011 (N_38011,N_37900,N_37732);
or U38012 (N_38012,N_37790,N_37556);
and U38013 (N_38013,N_37776,N_37752);
nor U38014 (N_38014,N_37853,N_37682);
or U38015 (N_38015,N_37646,N_37531);
or U38016 (N_38016,N_37766,N_37746);
and U38017 (N_38017,N_37883,N_37837);
and U38018 (N_38018,N_37863,N_37519);
xor U38019 (N_38019,N_37769,N_37669);
xnor U38020 (N_38020,N_37916,N_37755);
xnor U38021 (N_38021,N_37925,N_37572);
or U38022 (N_38022,N_37675,N_37570);
or U38023 (N_38023,N_37597,N_37534);
xor U38024 (N_38024,N_37631,N_37891);
or U38025 (N_38025,N_37525,N_37867);
nand U38026 (N_38026,N_37777,N_37854);
xnor U38027 (N_38027,N_37806,N_37927);
or U38028 (N_38028,N_37635,N_37641);
xor U38029 (N_38029,N_37710,N_37948);
xnor U38030 (N_38030,N_37502,N_37923);
nor U38031 (N_38031,N_37885,N_37742);
xnor U38032 (N_38032,N_37690,N_37697);
and U38033 (N_38033,N_37823,N_37743);
xor U38034 (N_38034,N_37521,N_37912);
nand U38035 (N_38035,N_37874,N_37802);
nand U38036 (N_38036,N_37623,N_37998);
nor U38037 (N_38037,N_37593,N_37562);
xnor U38038 (N_38038,N_37657,N_37763);
xnor U38039 (N_38039,N_37993,N_37899);
and U38040 (N_38040,N_37990,N_37713);
or U38041 (N_38041,N_37721,N_37590);
xnor U38042 (N_38042,N_37584,N_37674);
nand U38043 (N_38043,N_37528,N_37602);
nor U38044 (N_38044,N_37530,N_37793);
xor U38045 (N_38045,N_37754,N_37638);
nand U38046 (N_38046,N_37678,N_37789);
xnor U38047 (N_38047,N_37594,N_37999);
or U38048 (N_38048,N_37958,N_37692);
nor U38049 (N_38049,N_37799,N_37640);
nand U38050 (N_38050,N_37851,N_37578);
nand U38051 (N_38051,N_37985,N_37717);
or U38052 (N_38052,N_37508,N_37639);
or U38053 (N_38053,N_37771,N_37928);
and U38054 (N_38054,N_37745,N_37926);
and U38055 (N_38055,N_37796,N_37726);
xor U38056 (N_38056,N_37617,N_37811);
or U38057 (N_38057,N_37991,N_37812);
or U38058 (N_38058,N_37500,N_37870);
or U38059 (N_38059,N_37551,N_37784);
or U38060 (N_38060,N_37698,N_37892);
nand U38061 (N_38061,N_37574,N_37718);
nand U38062 (N_38062,N_37797,N_37566);
or U38063 (N_38063,N_37606,N_37917);
nand U38064 (N_38064,N_37960,N_37507);
nor U38065 (N_38065,N_37872,N_37954);
xnor U38066 (N_38066,N_37976,N_37968);
xor U38067 (N_38067,N_37820,N_37670);
nand U38068 (N_38068,N_37659,N_37715);
or U38069 (N_38069,N_37695,N_37773);
nand U38070 (N_38070,N_37905,N_37704);
nand U38071 (N_38071,N_37672,N_37921);
nand U38072 (N_38072,N_37583,N_37953);
xor U38073 (N_38073,N_37895,N_37988);
and U38074 (N_38074,N_37586,N_37611);
xnor U38075 (N_38075,N_37876,N_37832);
xor U38076 (N_38076,N_37901,N_37939);
or U38077 (N_38077,N_37549,N_37973);
or U38078 (N_38078,N_37936,N_37857);
and U38079 (N_38079,N_37795,N_37569);
or U38080 (N_38080,N_37527,N_37996);
or U38081 (N_38081,N_37884,N_37767);
and U38082 (N_38082,N_37546,N_37520);
and U38083 (N_38083,N_37821,N_37780);
and U38084 (N_38084,N_37902,N_37564);
nor U38085 (N_38085,N_37585,N_37523);
nor U38086 (N_38086,N_37918,N_37533);
nand U38087 (N_38087,N_37986,N_37539);
and U38088 (N_38088,N_37577,N_37749);
nand U38089 (N_38089,N_37693,N_37757);
nor U38090 (N_38090,N_37543,N_37592);
nand U38091 (N_38091,N_37794,N_37860);
xnor U38092 (N_38092,N_37803,N_37600);
or U38093 (N_38093,N_37817,N_37937);
xor U38094 (N_38094,N_37654,N_37858);
and U38095 (N_38095,N_37861,N_37840);
or U38096 (N_38096,N_37716,N_37829);
nor U38097 (N_38097,N_37681,N_37619);
or U38098 (N_38098,N_37753,N_37506);
and U38099 (N_38099,N_37977,N_37818);
nor U38100 (N_38100,N_37529,N_37620);
or U38101 (N_38101,N_37866,N_37890);
or U38102 (N_38102,N_37589,N_37804);
nand U38103 (N_38103,N_37856,N_37736);
and U38104 (N_38104,N_37645,N_37622);
xnor U38105 (N_38105,N_37788,N_37970);
nand U38106 (N_38106,N_37587,N_37935);
nor U38107 (N_38107,N_37580,N_37558);
xnor U38108 (N_38108,N_37878,N_37538);
xnor U38109 (N_38109,N_37852,N_37706);
nand U38110 (N_38110,N_37541,N_37740);
and U38111 (N_38111,N_37768,N_37945);
or U38112 (N_38112,N_37944,N_37709);
nor U38113 (N_38113,N_37687,N_37575);
nand U38114 (N_38114,N_37838,N_37588);
xnor U38115 (N_38115,N_37624,N_37783);
and U38116 (N_38116,N_37707,N_37610);
nor U38117 (N_38117,N_37571,N_37791);
or U38118 (N_38118,N_37971,N_37887);
xor U38119 (N_38119,N_37855,N_37552);
xnor U38120 (N_38120,N_37850,N_37881);
or U38121 (N_38121,N_37689,N_37898);
nor U38122 (N_38122,N_37932,N_37772);
xor U38123 (N_38123,N_37550,N_37511);
and U38124 (N_38124,N_37762,N_37972);
or U38125 (N_38125,N_37536,N_37738);
xnor U38126 (N_38126,N_37650,N_37633);
or U38127 (N_38127,N_37975,N_37560);
or U38128 (N_38128,N_37896,N_37515);
xnor U38129 (N_38129,N_37962,N_37605);
nand U38130 (N_38130,N_37952,N_37733);
or U38131 (N_38131,N_37751,N_37813);
xor U38132 (N_38132,N_37894,N_37608);
xnor U38133 (N_38133,N_37601,N_37844);
nor U38134 (N_38134,N_37748,N_37542);
nor U38135 (N_38135,N_37642,N_37532);
nand U38136 (N_38136,N_37626,N_37613);
nor U38137 (N_38137,N_37576,N_37634);
or U38138 (N_38138,N_37628,N_37956);
xor U38139 (N_38139,N_37764,N_37505);
or U38140 (N_38140,N_37967,N_37735);
xor U38141 (N_38141,N_37603,N_37513);
or U38142 (N_38142,N_37978,N_37625);
or U38143 (N_38143,N_37940,N_37688);
nor U38144 (N_38144,N_37660,N_37636);
nand U38145 (N_38145,N_37964,N_37873);
or U38146 (N_38146,N_37537,N_37963);
and U38147 (N_38147,N_37676,N_37679);
xor U38148 (N_38148,N_37522,N_37810);
nor U38149 (N_38149,N_37904,N_37792);
or U38150 (N_38150,N_37759,N_37651);
and U38151 (N_38151,N_37699,N_37787);
and U38152 (N_38152,N_37516,N_37518);
xnor U38153 (N_38153,N_37720,N_37691);
xor U38154 (N_38154,N_37929,N_37761);
nand U38155 (N_38155,N_37714,N_37992);
nand U38156 (N_38156,N_37744,N_37995);
nor U38157 (N_38157,N_37711,N_37616);
nand U38158 (N_38158,N_37683,N_37504);
or U38159 (N_38159,N_37568,N_37630);
and U38160 (N_38160,N_37822,N_37719);
or U38161 (N_38161,N_37581,N_37545);
nand U38162 (N_38162,N_37997,N_37983);
and U38163 (N_38163,N_37938,N_37877);
xnor U38164 (N_38164,N_37758,N_37906);
and U38165 (N_38165,N_37615,N_37785);
and U38166 (N_38166,N_37700,N_37598);
or U38167 (N_38167,N_37828,N_37947);
nor U38168 (N_38168,N_37664,N_37765);
or U38169 (N_38169,N_37868,N_37644);
and U38170 (N_38170,N_37557,N_37632);
xor U38171 (N_38171,N_37591,N_37680);
nor U38172 (N_38172,N_37893,N_37725);
nor U38173 (N_38173,N_37951,N_37565);
xnor U38174 (N_38174,N_37526,N_37987);
or U38175 (N_38175,N_37774,N_37982);
nor U38176 (N_38176,N_37665,N_37547);
nand U38177 (N_38177,N_37673,N_37729);
nand U38178 (N_38178,N_37553,N_37869);
and U38179 (N_38179,N_37782,N_37661);
xnor U38180 (N_38180,N_37612,N_37607);
nor U38181 (N_38181,N_37835,N_37671);
nor U38182 (N_38182,N_37554,N_37614);
nor U38183 (N_38183,N_37737,N_37750);
or U38184 (N_38184,N_37965,N_37712);
nor U38185 (N_38185,N_37825,N_37555);
nand U38186 (N_38186,N_37658,N_37643);
nor U38187 (N_38187,N_37666,N_37662);
and U38188 (N_38188,N_37703,N_37819);
and U38189 (N_38189,N_37846,N_37723);
nand U38190 (N_38190,N_37931,N_37910);
nand U38191 (N_38191,N_37824,N_37512);
xnor U38192 (N_38192,N_37563,N_37579);
nand U38193 (N_38193,N_37875,N_37779);
xor U38194 (N_38194,N_37880,N_37637);
nor U38195 (N_38195,N_37727,N_37980);
or U38196 (N_38196,N_37897,N_37559);
xnor U38197 (N_38197,N_37724,N_37839);
nor U38198 (N_38198,N_37913,N_37778);
and U38199 (N_38199,N_37848,N_37629);
nor U38200 (N_38200,N_37920,N_37979);
nand U38201 (N_38201,N_37705,N_37969);
nor U38202 (N_38202,N_37561,N_37696);
nor U38203 (N_38203,N_37663,N_37656);
nand U38204 (N_38204,N_37908,N_37984);
nor U38205 (N_38205,N_37827,N_37903);
nor U38206 (N_38206,N_37859,N_37648);
xnor U38207 (N_38207,N_37865,N_37686);
or U38208 (N_38208,N_37836,N_37950);
xor U38209 (N_38209,N_37847,N_37694);
xor U38210 (N_38210,N_37842,N_37915);
xnor U38211 (N_38211,N_37730,N_37599);
and U38212 (N_38212,N_37959,N_37573);
or U38213 (N_38213,N_37941,N_37889);
nand U38214 (N_38214,N_37957,N_37627);
nor U38215 (N_38215,N_37981,N_37974);
nand U38216 (N_38216,N_37833,N_37798);
nand U38217 (N_38217,N_37864,N_37756);
and U38218 (N_38218,N_37786,N_37775);
nor U38219 (N_38219,N_37930,N_37816);
nor U38220 (N_38220,N_37701,N_37919);
or U38221 (N_38221,N_37909,N_37805);
or U38222 (N_38222,N_37509,N_37649);
and U38223 (N_38223,N_37955,N_37914);
nor U38224 (N_38224,N_37510,N_37514);
nand U38225 (N_38225,N_37567,N_37685);
and U38226 (N_38226,N_37924,N_37621);
nor U38227 (N_38227,N_37596,N_37845);
and U38228 (N_38228,N_37934,N_37655);
nand U38229 (N_38229,N_37524,N_37830);
xnor U38230 (N_38230,N_37831,N_37800);
nand U38231 (N_38231,N_37647,N_37604);
and U38232 (N_38232,N_37922,N_37834);
nand U38233 (N_38233,N_37708,N_37741);
or U38234 (N_38234,N_37961,N_37849);
or U38235 (N_38235,N_37907,N_37728);
xnor U38236 (N_38236,N_37815,N_37801);
nor U38237 (N_38237,N_37994,N_37503);
or U38238 (N_38238,N_37760,N_37618);
nor U38239 (N_38239,N_37653,N_37652);
nand U38240 (N_38240,N_37843,N_37809);
xnor U38241 (N_38241,N_37807,N_37814);
or U38242 (N_38242,N_37933,N_37702);
or U38243 (N_38243,N_37886,N_37677);
and U38244 (N_38244,N_37882,N_37731);
or U38245 (N_38245,N_37911,N_37540);
and U38246 (N_38246,N_37879,N_37739);
nor U38247 (N_38247,N_37684,N_37943);
nand U38248 (N_38248,N_37722,N_37946);
and U38249 (N_38249,N_37548,N_37989);
and U38250 (N_38250,N_37671,N_37784);
nand U38251 (N_38251,N_37980,N_37769);
and U38252 (N_38252,N_37544,N_37512);
xor U38253 (N_38253,N_37856,N_37721);
nand U38254 (N_38254,N_37641,N_37967);
or U38255 (N_38255,N_37915,N_37700);
or U38256 (N_38256,N_37664,N_37850);
nand U38257 (N_38257,N_37615,N_37803);
xor U38258 (N_38258,N_37760,N_37972);
nand U38259 (N_38259,N_37857,N_37931);
and U38260 (N_38260,N_37829,N_37990);
xnor U38261 (N_38261,N_37666,N_37856);
nand U38262 (N_38262,N_37818,N_37636);
nand U38263 (N_38263,N_37966,N_37891);
and U38264 (N_38264,N_37615,N_37506);
nor U38265 (N_38265,N_37670,N_37816);
or U38266 (N_38266,N_37980,N_37684);
nor U38267 (N_38267,N_37973,N_37744);
nand U38268 (N_38268,N_37702,N_37779);
nand U38269 (N_38269,N_37998,N_37690);
or U38270 (N_38270,N_37746,N_37711);
nand U38271 (N_38271,N_37554,N_37569);
nor U38272 (N_38272,N_37763,N_37541);
xor U38273 (N_38273,N_37766,N_37572);
or U38274 (N_38274,N_37545,N_37934);
xnor U38275 (N_38275,N_37771,N_37505);
and U38276 (N_38276,N_37713,N_37791);
nand U38277 (N_38277,N_37592,N_37511);
or U38278 (N_38278,N_37777,N_37948);
nor U38279 (N_38279,N_37606,N_37724);
and U38280 (N_38280,N_37783,N_37956);
nand U38281 (N_38281,N_37684,N_37512);
and U38282 (N_38282,N_37993,N_37986);
xor U38283 (N_38283,N_37885,N_37891);
nand U38284 (N_38284,N_37525,N_37797);
nor U38285 (N_38285,N_37604,N_37659);
nand U38286 (N_38286,N_37709,N_37616);
nor U38287 (N_38287,N_37519,N_37807);
nor U38288 (N_38288,N_37718,N_37799);
nor U38289 (N_38289,N_37714,N_37596);
nand U38290 (N_38290,N_37783,N_37962);
and U38291 (N_38291,N_37811,N_37521);
xor U38292 (N_38292,N_37807,N_37888);
xnor U38293 (N_38293,N_37775,N_37576);
xor U38294 (N_38294,N_37767,N_37574);
nand U38295 (N_38295,N_37800,N_37832);
and U38296 (N_38296,N_37780,N_37611);
or U38297 (N_38297,N_37720,N_37975);
nand U38298 (N_38298,N_37799,N_37973);
nand U38299 (N_38299,N_37913,N_37729);
xor U38300 (N_38300,N_37820,N_37610);
or U38301 (N_38301,N_37675,N_37987);
nor U38302 (N_38302,N_37959,N_37761);
xnor U38303 (N_38303,N_37634,N_37902);
nand U38304 (N_38304,N_37609,N_37784);
xnor U38305 (N_38305,N_37987,N_37702);
and U38306 (N_38306,N_37993,N_37996);
nor U38307 (N_38307,N_37626,N_37661);
nand U38308 (N_38308,N_37815,N_37913);
or U38309 (N_38309,N_37575,N_37605);
xor U38310 (N_38310,N_37734,N_37642);
nand U38311 (N_38311,N_37884,N_37973);
nor U38312 (N_38312,N_37643,N_37771);
or U38313 (N_38313,N_37869,N_37992);
nor U38314 (N_38314,N_37604,N_37941);
xor U38315 (N_38315,N_37578,N_37700);
and U38316 (N_38316,N_37814,N_37743);
nor U38317 (N_38317,N_37728,N_37648);
nor U38318 (N_38318,N_37854,N_37704);
nand U38319 (N_38319,N_37946,N_37872);
nand U38320 (N_38320,N_37604,N_37897);
nor U38321 (N_38321,N_37532,N_37539);
nor U38322 (N_38322,N_37525,N_37857);
and U38323 (N_38323,N_37614,N_37624);
nor U38324 (N_38324,N_37525,N_37788);
nand U38325 (N_38325,N_37766,N_37824);
xor U38326 (N_38326,N_37801,N_37612);
and U38327 (N_38327,N_37935,N_37634);
nand U38328 (N_38328,N_37787,N_37643);
or U38329 (N_38329,N_37916,N_37751);
and U38330 (N_38330,N_37829,N_37801);
nand U38331 (N_38331,N_37544,N_37965);
or U38332 (N_38332,N_37571,N_37567);
and U38333 (N_38333,N_37562,N_37517);
and U38334 (N_38334,N_37595,N_37608);
nand U38335 (N_38335,N_37933,N_37607);
and U38336 (N_38336,N_37659,N_37710);
nand U38337 (N_38337,N_37849,N_37682);
or U38338 (N_38338,N_37540,N_37937);
or U38339 (N_38339,N_37760,N_37892);
nand U38340 (N_38340,N_37608,N_37676);
nand U38341 (N_38341,N_37744,N_37586);
nand U38342 (N_38342,N_37793,N_37868);
xor U38343 (N_38343,N_37991,N_37569);
nor U38344 (N_38344,N_37630,N_37710);
or U38345 (N_38345,N_37565,N_37541);
nor U38346 (N_38346,N_37961,N_37533);
or U38347 (N_38347,N_37611,N_37926);
xor U38348 (N_38348,N_37615,N_37989);
or U38349 (N_38349,N_37708,N_37794);
or U38350 (N_38350,N_37532,N_37847);
xor U38351 (N_38351,N_37718,N_37726);
nor U38352 (N_38352,N_37752,N_37697);
nand U38353 (N_38353,N_37507,N_37769);
nor U38354 (N_38354,N_37773,N_37866);
nor U38355 (N_38355,N_37938,N_37936);
or U38356 (N_38356,N_37916,N_37740);
xor U38357 (N_38357,N_37949,N_37585);
and U38358 (N_38358,N_37508,N_37927);
nor U38359 (N_38359,N_37586,N_37703);
xor U38360 (N_38360,N_37818,N_37629);
and U38361 (N_38361,N_37827,N_37790);
and U38362 (N_38362,N_37659,N_37632);
nand U38363 (N_38363,N_37502,N_37517);
and U38364 (N_38364,N_37919,N_37691);
and U38365 (N_38365,N_37688,N_37514);
xnor U38366 (N_38366,N_37871,N_37552);
nand U38367 (N_38367,N_37610,N_37635);
xor U38368 (N_38368,N_37815,N_37748);
and U38369 (N_38369,N_37720,N_37833);
xnor U38370 (N_38370,N_37519,N_37830);
nor U38371 (N_38371,N_37611,N_37695);
or U38372 (N_38372,N_37647,N_37636);
nor U38373 (N_38373,N_37908,N_37526);
nor U38374 (N_38374,N_37520,N_37933);
or U38375 (N_38375,N_37748,N_37934);
and U38376 (N_38376,N_37775,N_37779);
xnor U38377 (N_38377,N_37873,N_37787);
or U38378 (N_38378,N_37865,N_37961);
or U38379 (N_38379,N_37534,N_37737);
nand U38380 (N_38380,N_37774,N_37696);
or U38381 (N_38381,N_37594,N_37662);
nand U38382 (N_38382,N_37976,N_37706);
or U38383 (N_38383,N_37677,N_37867);
nand U38384 (N_38384,N_37894,N_37578);
xor U38385 (N_38385,N_37970,N_37825);
or U38386 (N_38386,N_37652,N_37829);
and U38387 (N_38387,N_37603,N_37656);
and U38388 (N_38388,N_37617,N_37534);
nand U38389 (N_38389,N_37562,N_37602);
or U38390 (N_38390,N_37823,N_37856);
or U38391 (N_38391,N_37688,N_37968);
and U38392 (N_38392,N_37822,N_37956);
xor U38393 (N_38393,N_37733,N_37878);
nor U38394 (N_38394,N_37506,N_37838);
and U38395 (N_38395,N_37915,N_37792);
or U38396 (N_38396,N_37805,N_37941);
nor U38397 (N_38397,N_37731,N_37944);
or U38398 (N_38398,N_37968,N_37894);
and U38399 (N_38399,N_37733,N_37874);
xor U38400 (N_38400,N_37804,N_37697);
nand U38401 (N_38401,N_37628,N_37527);
or U38402 (N_38402,N_37915,N_37561);
xor U38403 (N_38403,N_37600,N_37642);
nor U38404 (N_38404,N_37754,N_37574);
and U38405 (N_38405,N_37560,N_37992);
xor U38406 (N_38406,N_37912,N_37626);
nand U38407 (N_38407,N_37920,N_37698);
xor U38408 (N_38408,N_37906,N_37938);
nand U38409 (N_38409,N_37732,N_37680);
nor U38410 (N_38410,N_37663,N_37817);
or U38411 (N_38411,N_37555,N_37904);
nor U38412 (N_38412,N_37688,N_37906);
xnor U38413 (N_38413,N_37947,N_37595);
and U38414 (N_38414,N_37820,N_37669);
nor U38415 (N_38415,N_37908,N_37956);
nor U38416 (N_38416,N_37533,N_37730);
nor U38417 (N_38417,N_37775,N_37923);
nand U38418 (N_38418,N_37558,N_37754);
nand U38419 (N_38419,N_37629,N_37785);
xor U38420 (N_38420,N_37973,N_37529);
nor U38421 (N_38421,N_37890,N_37736);
nor U38422 (N_38422,N_37571,N_37855);
or U38423 (N_38423,N_37700,N_37632);
and U38424 (N_38424,N_37790,N_37611);
nand U38425 (N_38425,N_37937,N_37706);
and U38426 (N_38426,N_37762,N_37831);
or U38427 (N_38427,N_37821,N_37838);
nand U38428 (N_38428,N_37635,N_37636);
nand U38429 (N_38429,N_37694,N_37517);
and U38430 (N_38430,N_37724,N_37713);
nor U38431 (N_38431,N_37516,N_37545);
or U38432 (N_38432,N_37981,N_37791);
and U38433 (N_38433,N_37833,N_37637);
and U38434 (N_38434,N_37536,N_37789);
or U38435 (N_38435,N_37599,N_37676);
nor U38436 (N_38436,N_37525,N_37952);
xor U38437 (N_38437,N_37749,N_37960);
and U38438 (N_38438,N_37981,N_37968);
xnor U38439 (N_38439,N_37861,N_37502);
and U38440 (N_38440,N_37732,N_37534);
or U38441 (N_38441,N_37661,N_37722);
xnor U38442 (N_38442,N_37871,N_37660);
xor U38443 (N_38443,N_37939,N_37774);
or U38444 (N_38444,N_37961,N_37844);
nor U38445 (N_38445,N_37539,N_37958);
or U38446 (N_38446,N_37892,N_37749);
or U38447 (N_38447,N_37638,N_37681);
and U38448 (N_38448,N_37647,N_37936);
nand U38449 (N_38449,N_37819,N_37973);
nand U38450 (N_38450,N_37864,N_37865);
xor U38451 (N_38451,N_37588,N_37951);
nor U38452 (N_38452,N_37514,N_37802);
nand U38453 (N_38453,N_37915,N_37800);
or U38454 (N_38454,N_37787,N_37909);
nor U38455 (N_38455,N_37664,N_37864);
nor U38456 (N_38456,N_37803,N_37531);
xnor U38457 (N_38457,N_37515,N_37606);
or U38458 (N_38458,N_37601,N_37876);
nor U38459 (N_38459,N_37877,N_37761);
nand U38460 (N_38460,N_37505,N_37590);
or U38461 (N_38461,N_37711,N_37511);
nor U38462 (N_38462,N_37817,N_37889);
or U38463 (N_38463,N_37751,N_37790);
nand U38464 (N_38464,N_37899,N_37690);
nor U38465 (N_38465,N_37516,N_37795);
or U38466 (N_38466,N_37955,N_37848);
nand U38467 (N_38467,N_37799,N_37544);
xnor U38468 (N_38468,N_37665,N_37669);
nand U38469 (N_38469,N_37822,N_37693);
nor U38470 (N_38470,N_37932,N_37917);
and U38471 (N_38471,N_37890,N_37615);
and U38472 (N_38472,N_37640,N_37797);
or U38473 (N_38473,N_37758,N_37923);
and U38474 (N_38474,N_37663,N_37775);
or U38475 (N_38475,N_37689,N_37603);
and U38476 (N_38476,N_37779,N_37899);
or U38477 (N_38477,N_37860,N_37905);
and U38478 (N_38478,N_37704,N_37575);
xor U38479 (N_38479,N_37554,N_37647);
and U38480 (N_38480,N_37798,N_37832);
and U38481 (N_38481,N_37739,N_37515);
nor U38482 (N_38482,N_37908,N_37631);
or U38483 (N_38483,N_37863,N_37646);
xnor U38484 (N_38484,N_37972,N_37979);
nor U38485 (N_38485,N_37616,N_37916);
or U38486 (N_38486,N_37775,N_37833);
nor U38487 (N_38487,N_37850,N_37849);
nand U38488 (N_38488,N_37607,N_37971);
or U38489 (N_38489,N_37558,N_37766);
nand U38490 (N_38490,N_37582,N_37764);
or U38491 (N_38491,N_37564,N_37888);
and U38492 (N_38492,N_37852,N_37661);
nor U38493 (N_38493,N_37987,N_37627);
xnor U38494 (N_38494,N_37805,N_37510);
nand U38495 (N_38495,N_37842,N_37905);
or U38496 (N_38496,N_37622,N_37606);
or U38497 (N_38497,N_37534,N_37645);
xor U38498 (N_38498,N_37604,N_37704);
and U38499 (N_38499,N_37917,N_37760);
and U38500 (N_38500,N_38251,N_38400);
nand U38501 (N_38501,N_38184,N_38076);
nand U38502 (N_38502,N_38351,N_38346);
nor U38503 (N_38503,N_38434,N_38454);
nor U38504 (N_38504,N_38086,N_38422);
nor U38505 (N_38505,N_38332,N_38408);
and U38506 (N_38506,N_38019,N_38231);
or U38507 (N_38507,N_38483,N_38381);
or U38508 (N_38508,N_38083,N_38432);
or U38509 (N_38509,N_38136,N_38243);
nand U38510 (N_38510,N_38016,N_38262);
and U38511 (N_38511,N_38485,N_38156);
nor U38512 (N_38512,N_38097,N_38438);
nor U38513 (N_38513,N_38134,N_38363);
or U38514 (N_38514,N_38385,N_38326);
and U38515 (N_38515,N_38224,N_38366);
or U38516 (N_38516,N_38008,N_38225);
or U38517 (N_38517,N_38190,N_38331);
or U38518 (N_38518,N_38135,N_38102);
or U38519 (N_38519,N_38461,N_38232);
or U38520 (N_38520,N_38012,N_38169);
nor U38521 (N_38521,N_38066,N_38397);
and U38522 (N_38522,N_38226,N_38374);
and U38523 (N_38523,N_38100,N_38177);
and U38524 (N_38524,N_38093,N_38072);
nor U38525 (N_38525,N_38281,N_38044);
nand U38526 (N_38526,N_38162,N_38201);
xor U38527 (N_38527,N_38234,N_38050);
nor U38528 (N_38528,N_38247,N_38452);
or U38529 (N_38529,N_38430,N_38273);
nand U38530 (N_38530,N_38294,N_38401);
nand U38531 (N_38531,N_38194,N_38200);
xor U38532 (N_38532,N_38146,N_38176);
xnor U38533 (N_38533,N_38268,N_38042);
nand U38534 (N_38534,N_38227,N_38445);
xnor U38535 (N_38535,N_38034,N_38017);
xnor U38536 (N_38536,N_38090,N_38298);
xnor U38537 (N_38537,N_38185,N_38412);
nand U38538 (N_38538,N_38478,N_38300);
xnor U38539 (N_38539,N_38143,N_38155);
or U38540 (N_38540,N_38254,N_38117);
nand U38541 (N_38541,N_38498,N_38047);
and U38542 (N_38542,N_38427,N_38203);
and U38543 (N_38543,N_38088,N_38235);
and U38544 (N_38544,N_38271,N_38046);
nor U38545 (N_38545,N_38256,N_38447);
xnor U38546 (N_38546,N_38323,N_38221);
xnor U38547 (N_38547,N_38236,N_38295);
or U38548 (N_38548,N_38015,N_38286);
nand U38549 (N_38549,N_38063,N_38239);
or U38550 (N_38550,N_38023,N_38322);
or U38551 (N_38551,N_38187,N_38101);
nor U38552 (N_38552,N_38089,N_38475);
nor U38553 (N_38553,N_38108,N_38186);
nor U38554 (N_38554,N_38278,N_38469);
xnor U38555 (N_38555,N_38440,N_38407);
nand U38556 (N_38556,N_38214,N_38104);
xnor U38557 (N_38557,N_38379,N_38010);
nor U38558 (N_38558,N_38168,N_38174);
nor U38559 (N_38559,N_38116,N_38428);
xor U38560 (N_38560,N_38065,N_38071);
and U38561 (N_38561,N_38140,N_38055);
nand U38562 (N_38562,N_38433,N_38386);
nand U38563 (N_38563,N_38314,N_38204);
and U38564 (N_38564,N_38005,N_38343);
nand U38565 (N_38565,N_38069,N_38431);
nor U38566 (N_38566,N_38474,N_38142);
nor U38567 (N_38567,N_38033,N_38161);
and U38568 (N_38568,N_38121,N_38052);
or U38569 (N_38569,N_38457,N_38098);
nand U38570 (N_38570,N_38337,N_38419);
xnor U38571 (N_38571,N_38425,N_38289);
or U38572 (N_38572,N_38127,N_38311);
and U38573 (N_38573,N_38164,N_38335);
and U38574 (N_38574,N_38391,N_38356);
xor U38575 (N_38575,N_38373,N_38287);
and U38576 (N_38576,N_38417,N_38399);
and U38577 (N_38577,N_38423,N_38338);
nor U38578 (N_38578,N_38026,N_38358);
or U38579 (N_38579,N_38499,N_38248);
or U38580 (N_38580,N_38141,N_38384);
and U38581 (N_38581,N_38077,N_38280);
xnor U38582 (N_38582,N_38021,N_38179);
or U38583 (N_38583,N_38492,N_38151);
xor U38584 (N_38584,N_38276,N_38181);
xnor U38585 (N_38585,N_38429,N_38360);
xor U38586 (N_38586,N_38370,N_38109);
nand U38587 (N_38587,N_38105,N_38094);
xor U38588 (N_38588,N_38199,N_38013);
nand U38589 (N_38589,N_38103,N_38441);
nor U38590 (N_38590,N_38389,N_38087);
or U38591 (N_38591,N_38189,N_38230);
and U38592 (N_38592,N_38306,N_38488);
nand U38593 (N_38593,N_38325,N_38067);
or U38594 (N_38594,N_38395,N_38375);
nand U38595 (N_38595,N_38303,N_38007);
and U38596 (N_38596,N_38319,N_38240);
nor U38597 (N_38597,N_38315,N_38107);
or U38598 (N_38598,N_38171,N_38345);
nor U38599 (N_38599,N_38154,N_38215);
nor U38600 (N_38600,N_38416,N_38031);
nor U38601 (N_38601,N_38341,N_38182);
nand U38602 (N_38602,N_38147,N_38367);
nand U38603 (N_38603,N_38279,N_38329);
nand U38604 (N_38604,N_38292,N_38223);
or U38605 (N_38605,N_38213,N_38470);
nor U38606 (N_38606,N_38170,N_38043);
xor U38607 (N_38607,N_38482,N_38139);
nand U38608 (N_38608,N_38450,N_38383);
xnor U38609 (N_38609,N_38006,N_38233);
xor U38610 (N_38610,N_38409,N_38150);
and U38611 (N_38611,N_38082,N_38144);
xnor U38612 (N_38612,N_38489,N_38411);
nand U38613 (N_38613,N_38002,N_38096);
nand U38614 (N_38614,N_38321,N_38263);
nand U38615 (N_38615,N_38259,N_38192);
xor U38616 (N_38616,N_38106,N_38218);
nand U38617 (N_38617,N_38282,N_38426);
nand U38618 (N_38618,N_38078,N_38152);
xnor U38619 (N_38619,N_38372,N_38133);
xnor U38620 (N_38620,N_38352,N_38443);
or U38621 (N_38621,N_38284,N_38111);
xor U38622 (N_38622,N_38403,N_38471);
nand U38623 (N_38623,N_38449,N_38039);
and U38624 (N_38624,N_38486,N_38160);
xnor U38625 (N_38625,N_38365,N_38081);
nor U38626 (N_38626,N_38264,N_38359);
and U38627 (N_38627,N_38467,N_38004);
or U38628 (N_38628,N_38491,N_38217);
and U38629 (N_38629,N_38056,N_38442);
nand U38630 (N_38630,N_38269,N_38393);
or U38631 (N_38631,N_38252,N_38421);
nor U38632 (N_38632,N_38418,N_38458);
and U38633 (N_38633,N_38355,N_38466);
nand U38634 (N_38634,N_38456,N_38420);
nor U38635 (N_38635,N_38099,N_38244);
and U38636 (N_38636,N_38377,N_38130);
nand U38637 (N_38637,N_38357,N_38413);
xnor U38638 (N_38638,N_38313,N_38333);
xnor U38639 (N_38639,N_38038,N_38241);
nand U38640 (N_38640,N_38362,N_38166);
xor U38641 (N_38641,N_38245,N_38446);
nand U38642 (N_38642,N_38030,N_38250);
nor U38643 (N_38643,N_38159,N_38301);
or U38644 (N_38644,N_38188,N_38484);
xor U38645 (N_38645,N_38493,N_38414);
nor U38646 (N_38646,N_38032,N_38029);
nor U38647 (N_38647,N_38132,N_38059);
and U38648 (N_38648,N_38037,N_38191);
or U38649 (N_38649,N_38149,N_38324);
xor U38650 (N_38650,N_38137,N_38092);
and U38651 (N_38651,N_38126,N_38095);
nand U38652 (N_38652,N_38476,N_38153);
or U38653 (N_38653,N_38451,N_38229);
and U38654 (N_38654,N_38064,N_38157);
nor U38655 (N_38655,N_38020,N_38439);
nor U38656 (N_38656,N_38291,N_38237);
xnor U38657 (N_38657,N_38158,N_38041);
nand U38658 (N_38658,N_38207,N_38062);
and U38659 (N_38659,N_38079,N_38275);
nand U38660 (N_38660,N_38304,N_38353);
xor U38661 (N_38661,N_38009,N_38261);
nor U38662 (N_38662,N_38018,N_38208);
or U38663 (N_38663,N_38260,N_38057);
or U38664 (N_38664,N_38025,N_38198);
or U38665 (N_38665,N_38496,N_38196);
nor U38666 (N_38666,N_38073,N_38435);
nor U38667 (N_38667,N_38288,N_38061);
xor U38668 (N_38668,N_38472,N_38495);
or U38669 (N_38669,N_38124,N_38197);
nor U38670 (N_38670,N_38308,N_38255);
xor U38671 (N_38671,N_38173,N_38388);
xor U38672 (N_38672,N_38129,N_38054);
nand U38673 (N_38673,N_38394,N_38001);
xor U38674 (N_38674,N_38481,N_38206);
and U38675 (N_38675,N_38115,N_38216);
and U38676 (N_38676,N_38497,N_38048);
and U38677 (N_38677,N_38336,N_38014);
nand U38678 (N_38678,N_38131,N_38340);
and U38679 (N_38679,N_38238,N_38487);
or U38680 (N_38680,N_38228,N_38285);
and U38681 (N_38681,N_38257,N_38272);
nor U38682 (N_38682,N_38479,N_38053);
nand U38683 (N_38683,N_38145,N_38113);
or U38684 (N_38684,N_38163,N_38348);
nor U38685 (N_38685,N_38328,N_38309);
or U38686 (N_38686,N_38327,N_38212);
and U38687 (N_38687,N_38410,N_38277);
nand U38688 (N_38688,N_38027,N_38220);
xor U38689 (N_38689,N_38125,N_38293);
and U38690 (N_38690,N_38468,N_38296);
nand U38691 (N_38691,N_38242,N_38070);
xor U38692 (N_38692,N_38305,N_38371);
xnor U38693 (N_38693,N_38024,N_38320);
xor U38694 (N_38694,N_38480,N_38148);
or U38695 (N_38695,N_38274,N_38354);
and U38696 (N_38696,N_38368,N_38459);
or U38697 (N_38697,N_38376,N_38219);
nand U38698 (N_38698,N_38473,N_38202);
nor U38699 (N_38699,N_38075,N_38378);
or U38700 (N_38700,N_38045,N_38364);
and U38701 (N_38701,N_38011,N_38036);
and U38702 (N_38702,N_38369,N_38302);
nand U38703 (N_38703,N_38334,N_38347);
xor U38704 (N_38704,N_38205,N_38193);
nor U38705 (N_38705,N_38380,N_38490);
xnor U38706 (N_38706,N_38477,N_38084);
xnor U38707 (N_38707,N_38265,N_38003);
nand U38708 (N_38708,N_38270,N_38119);
or U38709 (N_38709,N_38339,N_38211);
and U38710 (N_38710,N_38175,N_38316);
or U38711 (N_38711,N_38415,N_38058);
and U38712 (N_38712,N_38290,N_38349);
and U38713 (N_38713,N_38091,N_38035);
xnor U38714 (N_38714,N_38167,N_38382);
and U38715 (N_38715,N_38249,N_38222);
nand U38716 (N_38716,N_38455,N_38404);
nand U38717 (N_38717,N_38246,N_38118);
xor U38718 (N_38718,N_38494,N_38283);
nor U38719 (N_38719,N_38266,N_38460);
xor U38720 (N_38720,N_38465,N_38138);
nor U38721 (N_38721,N_38396,N_38342);
xor U38722 (N_38722,N_38317,N_38299);
nor U38723 (N_38723,N_38258,N_38398);
or U38724 (N_38724,N_38074,N_38209);
xnor U38725 (N_38725,N_38128,N_38436);
and U38726 (N_38726,N_38210,N_38444);
xnor U38727 (N_38727,N_38040,N_38405);
and U38728 (N_38728,N_38297,N_38307);
xor U38729 (N_38729,N_38028,N_38253);
nand U38730 (N_38730,N_38310,N_38267);
and U38731 (N_38731,N_38049,N_38392);
or U38732 (N_38732,N_38406,N_38463);
nand U38733 (N_38733,N_38361,N_38344);
nand U38734 (N_38734,N_38330,N_38462);
or U38735 (N_38735,N_38318,N_38448);
nand U38736 (N_38736,N_38060,N_38437);
nor U38737 (N_38737,N_38068,N_38165);
or U38738 (N_38738,N_38402,N_38112);
xor U38739 (N_38739,N_38178,N_38085);
nor U38740 (N_38740,N_38051,N_38390);
and U38741 (N_38741,N_38114,N_38022);
nor U38742 (N_38742,N_38000,N_38172);
nand U38743 (N_38743,N_38123,N_38080);
xnor U38744 (N_38744,N_38350,N_38183);
nand U38745 (N_38745,N_38120,N_38387);
and U38746 (N_38746,N_38424,N_38453);
nor U38747 (N_38747,N_38122,N_38312);
or U38748 (N_38748,N_38464,N_38180);
xor U38749 (N_38749,N_38195,N_38110);
xor U38750 (N_38750,N_38258,N_38455);
or U38751 (N_38751,N_38130,N_38059);
nor U38752 (N_38752,N_38292,N_38407);
nor U38753 (N_38753,N_38366,N_38315);
or U38754 (N_38754,N_38142,N_38459);
xor U38755 (N_38755,N_38193,N_38460);
or U38756 (N_38756,N_38224,N_38190);
and U38757 (N_38757,N_38369,N_38281);
and U38758 (N_38758,N_38468,N_38378);
xnor U38759 (N_38759,N_38007,N_38151);
and U38760 (N_38760,N_38276,N_38114);
nand U38761 (N_38761,N_38258,N_38078);
xor U38762 (N_38762,N_38076,N_38380);
nand U38763 (N_38763,N_38256,N_38090);
and U38764 (N_38764,N_38158,N_38281);
or U38765 (N_38765,N_38234,N_38090);
nor U38766 (N_38766,N_38119,N_38433);
or U38767 (N_38767,N_38411,N_38259);
nand U38768 (N_38768,N_38007,N_38228);
and U38769 (N_38769,N_38299,N_38183);
and U38770 (N_38770,N_38331,N_38322);
nand U38771 (N_38771,N_38365,N_38278);
nand U38772 (N_38772,N_38477,N_38232);
nor U38773 (N_38773,N_38277,N_38115);
or U38774 (N_38774,N_38127,N_38033);
nor U38775 (N_38775,N_38111,N_38124);
or U38776 (N_38776,N_38109,N_38013);
nand U38777 (N_38777,N_38449,N_38461);
or U38778 (N_38778,N_38463,N_38441);
or U38779 (N_38779,N_38474,N_38236);
xor U38780 (N_38780,N_38190,N_38440);
or U38781 (N_38781,N_38485,N_38212);
or U38782 (N_38782,N_38448,N_38059);
and U38783 (N_38783,N_38474,N_38081);
nor U38784 (N_38784,N_38125,N_38003);
or U38785 (N_38785,N_38077,N_38346);
xnor U38786 (N_38786,N_38193,N_38406);
nand U38787 (N_38787,N_38261,N_38295);
nor U38788 (N_38788,N_38202,N_38261);
and U38789 (N_38789,N_38273,N_38496);
and U38790 (N_38790,N_38115,N_38184);
nor U38791 (N_38791,N_38140,N_38388);
or U38792 (N_38792,N_38482,N_38454);
or U38793 (N_38793,N_38048,N_38492);
or U38794 (N_38794,N_38028,N_38120);
xnor U38795 (N_38795,N_38405,N_38323);
xor U38796 (N_38796,N_38298,N_38352);
nor U38797 (N_38797,N_38132,N_38355);
or U38798 (N_38798,N_38315,N_38378);
xnor U38799 (N_38799,N_38118,N_38343);
xnor U38800 (N_38800,N_38066,N_38385);
and U38801 (N_38801,N_38349,N_38458);
nor U38802 (N_38802,N_38326,N_38238);
xnor U38803 (N_38803,N_38129,N_38394);
xnor U38804 (N_38804,N_38339,N_38464);
and U38805 (N_38805,N_38144,N_38286);
nor U38806 (N_38806,N_38267,N_38445);
and U38807 (N_38807,N_38390,N_38431);
nor U38808 (N_38808,N_38159,N_38425);
and U38809 (N_38809,N_38323,N_38203);
and U38810 (N_38810,N_38089,N_38466);
nand U38811 (N_38811,N_38112,N_38020);
nand U38812 (N_38812,N_38276,N_38410);
or U38813 (N_38813,N_38261,N_38296);
or U38814 (N_38814,N_38372,N_38059);
or U38815 (N_38815,N_38479,N_38209);
nor U38816 (N_38816,N_38192,N_38263);
nand U38817 (N_38817,N_38380,N_38471);
xor U38818 (N_38818,N_38316,N_38071);
xnor U38819 (N_38819,N_38126,N_38294);
and U38820 (N_38820,N_38032,N_38083);
and U38821 (N_38821,N_38445,N_38131);
xor U38822 (N_38822,N_38106,N_38135);
nor U38823 (N_38823,N_38001,N_38199);
nand U38824 (N_38824,N_38276,N_38426);
nor U38825 (N_38825,N_38298,N_38136);
and U38826 (N_38826,N_38274,N_38104);
nor U38827 (N_38827,N_38122,N_38459);
xnor U38828 (N_38828,N_38071,N_38389);
nand U38829 (N_38829,N_38278,N_38114);
nor U38830 (N_38830,N_38130,N_38040);
and U38831 (N_38831,N_38268,N_38028);
nand U38832 (N_38832,N_38022,N_38045);
nand U38833 (N_38833,N_38273,N_38187);
xor U38834 (N_38834,N_38158,N_38305);
or U38835 (N_38835,N_38048,N_38076);
and U38836 (N_38836,N_38039,N_38233);
nand U38837 (N_38837,N_38190,N_38201);
nand U38838 (N_38838,N_38421,N_38189);
and U38839 (N_38839,N_38083,N_38320);
xor U38840 (N_38840,N_38332,N_38305);
or U38841 (N_38841,N_38251,N_38315);
nor U38842 (N_38842,N_38473,N_38231);
nor U38843 (N_38843,N_38187,N_38114);
and U38844 (N_38844,N_38124,N_38382);
or U38845 (N_38845,N_38179,N_38468);
xor U38846 (N_38846,N_38227,N_38133);
or U38847 (N_38847,N_38049,N_38424);
or U38848 (N_38848,N_38030,N_38426);
nor U38849 (N_38849,N_38177,N_38234);
nor U38850 (N_38850,N_38172,N_38251);
nor U38851 (N_38851,N_38245,N_38071);
and U38852 (N_38852,N_38368,N_38405);
xor U38853 (N_38853,N_38134,N_38016);
and U38854 (N_38854,N_38455,N_38062);
nor U38855 (N_38855,N_38178,N_38310);
and U38856 (N_38856,N_38311,N_38251);
nor U38857 (N_38857,N_38208,N_38050);
and U38858 (N_38858,N_38280,N_38369);
and U38859 (N_38859,N_38332,N_38272);
and U38860 (N_38860,N_38430,N_38359);
nor U38861 (N_38861,N_38478,N_38430);
xnor U38862 (N_38862,N_38172,N_38496);
nor U38863 (N_38863,N_38165,N_38361);
and U38864 (N_38864,N_38182,N_38430);
nor U38865 (N_38865,N_38237,N_38085);
or U38866 (N_38866,N_38203,N_38395);
xor U38867 (N_38867,N_38446,N_38331);
nand U38868 (N_38868,N_38074,N_38447);
nor U38869 (N_38869,N_38394,N_38033);
nor U38870 (N_38870,N_38221,N_38399);
nand U38871 (N_38871,N_38057,N_38177);
or U38872 (N_38872,N_38362,N_38306);
nand U38873 (N_38873,N_38424,N_38446);
and U38874 (N_38874,N_38316,N_38345);
or U38875 (N_38875,N_38395,N_38487);
or U38876 (N_38876,N_38314,N_38341);
nand U38877 (N_38877,N_38041,N_38324);
nor U38878 (N_38878,N_38444,N_38470);
xor U38879 (N_38879,N_38422,N_38031);
or U38880 (N_38880,N_38185,N_38294);
nand U38881 (N_38881,N_38409,N_38056);
nor U38882 (N_38882,N_38228,N_38490);
and U38883 (N_38883,N_38186,N_38486);
or U38884 (N_38884,N_38411,N_38112);
nand U38885 (N_38885,N_38354,N_38325);
nor U38886 (N_38886,N_38100,N_38354);
nand U38887 (N_38887,N_38076,N_38128);
and U38888 (N_38888,N_38445,N_38302);
nor U38889 (N_38889,N_38082,N_38352);
or U38890 (N_38890,N_38116,N_38414);
xnor U38891 (N_38891,N_38194,N_38152);
and U38892 (N_38892,N_38186,N_38433);
nor U38893 (N_38893,N_38029,N_38370);
xor U38894 (N_38894,N_38135,N_38377);
nor U38895 (N_38895,N_38133,N_38432);
nor U38896 (N_38896,N_38011,N_38089);
xor U38897 (N_38897,N_38205,N_38431);
or U38898 (N_38898,N_38449,N_38235);
nor U38899 (N_38899,N_38102,N_38473);
nand U38900 (N_38900,N_38474,N_38011);
nand U38901 (N_38901,N_38026,N_38470);
nor U38902 (N_38902,N_38446,N_38379);
nand U38903 (N_38903,N_38398,N_38151);
or U38904 (N_38904,N_38119,N_38406);
or U38905 (N_38905,N_38495,N_38414);
xnor U38906 (N_38906,N_38014,N_38060);
and U38907 (N_38907,N_38293,N_38256);
and U38908 (N_38908,N_38101,N_38369);
xnor U38909 (N_38909,N_38290,N_38119);
and U38910 (N_38910,N_38110,N_38221);
nand U38911 (N_38911,N_38063,N_38323);
nand U38912 (N_38912,N_38009,N_38052);
nand U38913 (N_38913,N_38140,N_38227);
nor U38914 (N_38914,N_38480,N_38130);
and U38915 (N_38915,N_38039,N_38196);
nor U38916 (N_38916,N_38431,N_38038);
or U38917 (N_38917,N_38188,N_38241);
and U38918 (N_38918,N_38022,N_38396);
nor U38919 (N_38919,N_38355,N_38154);
nor U38920 (N_38920,N_38301,N_38480);
nand U38921 (N_38921,N_38376,N_38020);
nor U38922 (N_38922,N_38442,N_38351);
and U38923 (N_38923,N_38165,N_38085);
xnor U38924 (N_38924,N_38147,N_38111);
xnor U38925 (N_38925,N_38050,N_38045);
nor U38926 (N_38926,N_38487,N_38232);
nor U38927 (N_38927,N_38003,N_38291);
nand U38928 (N_38928,N_38182,N_38003);
nor U38929 (N_38929,N_38329,N_38061);
nor U38930 (N_38930,N_38378,N_38427);
xnor U38931 (N_38931,N_38081,N_38055);
nand U38932 (N_38932,N_38140,N_38174);
nor U38933 (N_38933,N_38141,N_38355);
and U38934 (N_38934,N_38240,N_38303);
nor U38935 (N_38935,N_38063,N_38209);
and U38936 (N_38936,N_38368,N_38260);
and U38937 (N_38937,N_38421,N_38140);
nor U38938 (N_38938,N_38099,N_38477);
nor U38939 (N_38939,N_38470,N_38384);
xnor U38940 (N_38940,N_38248,N_38108);
or U38941 (N_38941,N_38385,N_38265);
nand U38942 (N_38942,N_38199,N_38324);
xnor U38943 (N_38943,N_38351,N_38244);
and U38944 (N_38944,N_38407,N_38155);
or U38945 (N_38945,N_38417,N_38345);
xnor U38946 (N_38946,N_38256,N_38052);
or U38947 (N_38947,N_38272,N_38363);
xnor U38948 (N_38948,N_38069,N_38446);
or U38949 (N_38949,N_38398,N_38244);
nand U38950 (N_38950,N_38408,N_38437);
xor U38951 (N_38951,N_38397,N_38428);
nor U38952 (N_38952,N_38347,N_38318);
nand U38953 (N_38953,N_38277,N_38280);
nand U38954 (N_38954,N_38363,N_38403);
or U38955 (N_38955,N_38035,N_38155);
xnor U38956 (N_38956,N_38455,N_38427);
and U38957 (N_38957,N_38299,N_38094);
or U38958 (N_38958,N_38256,N_38413);
or U38959 (N_38959,N_38199,N_38021);
xor U38960 (N_38960,N_38479,N_38392);
nor U38961 (N_38961,N_38259,N_38106);
xor U38962 (N_38962,N_38425,N_38002);
or U38963 (N_38963,N_38458,N_38234);
and U38964 (N_38964,N_38122,N_38485);
and U38965 (N_38965,N_38186,N_38488);
nand U38966 (N_38966,N_38371,N_38104);
nor U38967 (N_38967,N_38143,N_38291);
and U38968 (N_38968,N_38277,N_38164);
nor U38969 (N_38969,N_38012,N_38400);
xor U38970 (N_38970,N_38245,N_38030);
nand U38971 (N_38971,N_38017,N_38138);
nor U38972 (N_38972,N_38357,N_38158);
nor U38973 (N_38973,N_38244,N_38016);
xor U38974 (N_38974,N_38051,N_38228);
and U38975 (N_38975,N_38046,N_38488);
or U38976 (N_38976,N_38250,N_38463);
nand U38977 (N_38977,N_38181,N_38316);
or U38978 (N_38978,N_38448,N_38240);
nor U38979 (N_38979,N_38015,N_38027);
nor U38980 (N_38980,N_38412,N_38071);
nand U38981 (N_38981,N_38280,N_38379);
nand U38982 (N_38982,N_38044,N_38114);
xor U38983 (N_38983,N_38211,N_38197);
and U38984 (N_38984,N_38464,N_38149);
or U38985 (N_38985,N_38044,N_38407);
and U38986 (N_38986,N_38436,N_38067);
nor U38987 (N_38987,N_38065,N_38409);
and U38988 (N_38988,N_38454,N_38077);
nor U38989 (N_38989,N_38176,N_38245);
or U38990 (N_38990,N_38132,N_38225);
or U38991 (N_38991,N_38169,N_38139);
nor U38992 (N_38992,N_38097,N_38297);
nor U38993 (N_38993,N_38436,N_38155);
nand U38994 (N_38994,N_38304,N_38285);
nor U38995 (N_38995,N_38076,N_38482);
nor U38996 (N_38996,N_38469,N_38225);
and U38997 (N_38997,N_38107,N_38045);
nor U38998 (N_38998,N_38256,N_38257);
or U38999 (N_38999,N_38490,N_38126);
xor U39000 (N_39000,N_38632,N_38587);
nor U39001 (N_39001,N_38583,N_38575);
and U39002 (N_39002,N_38907,N_38721);
or U39003 (N_39003,N_38897,N_38935);
or U39004 (N_39004,N_38613,N_38848);
and U39005 (N_39005,N_38745,N_38875);
or U39006 (N_39006,N_38657,N_38547);
xor U39007 (N_39007,N_38685,N_38866);
xnor U39008 (N_39008,N_38682,N_38787);
and U39009 (N_39009,N_38506,N_38692);
nor U39010 (N_39010,N_38643,N_38957);
and U39011 (N_39011,N_38695,N_38654);
nor U39012 (N_39012,N_38730,N_38604);
or U39013 (N_39013,N_38983,N_38768);
and U39014 (N_39014,N_38633,N_38656);
and U39015 (N_39015,N_38681,N_38725);
or U39016 (N_39016,N_38786,N_38838);
and U39017 (N_39017,N_38647,N_38658);
and U39018 (N_39018,N_38963,N_38723);
and U39019 (N_39019,N_38781,N_38899);
nor U39020 (N_39020,N_38586,N_38828);
nor U39021 (N_39021,N_38571,N_38717);
nand U39022 (N_39022,N_38594,N_38732);
nor U39023 (N_39023,N_38758,N_38511);
and U39024 (N_39024,N_38967,N_38500);
xor U39025 (N_39025,N_38562,N_38669);
xor U39026 (N_39026,N_38520,N_38534);
xor U39027 (N_39027,N_38878,N_38573);
or U39028 (N_39028,N_38545,N_38574);
nand U39029 (N_39029,N_38955,N_38733);
nand U39030 (N_39030,N_38585,N_38936);
nor U39031 (N_39031,N_38973,N_38784);
nand U39032 (N_39032,N_38831,N_38771);
xor U39033 (N_39033,N_38942,N_38618);
nand U39034 (N_39034,N_38922,N_38515);
or U39035 (N_39035,N_38794,N_38765);
nand U39036 (N_39036,N_38990,N_38531);
and U39037 (N_39037,N_38568,N_38947);
nor U39038 (N_39038,N_38852,N_38865);
and U39039 (N_39039,N_38555,N_38505);
nor U39040 (N_39040,N_38700,N_38729);
nand U39041 (N_39041,N_38927,N_38803);
or U39042 (N_39042,N_38611,N_38739);
xor U39043 (N_39043,N_38513,N_38814);
xor U39044 (N_39044,N_38811,N_38982);
xor U39045 (N_39045,N_38903,N_38740);
and U39046 (N_39046,N_38665,N_38652);
or U39047 (N_39047,N_38761,N_38966);
and U39048 (N_39048,N_38638,N_38813);
nand U39049 (N_39049,N_38501,N_38653);
and U39050 (N_39050,N_38807,N_38661);
xor U39051 (N_39051,N_38645,N_38667);
nor U39052 (N_39052,N_38835,N_38960);
nor U39053 (N_39053,N_38524,N_38526);
or U39054 (N_39054,N_38726,N_38623);
or U39055 (N_39055,N_38854,N_38541);
or U39056 (N_39056,N_38876,N_38651);
nand U39057 (N_39057,N_38577,N_38543);
nor U39058 (N_39058,N_38671,N_38954);
or U39059 (N_39059,N_38868,N_38995);
and U39060 (N_39060,N_38754,N_38608);
nor U39061 (N_39061,N_38523,N_38715);
xor U39062 (N_39062,N_38710,N_38528);
and U39063 (N_39063,N_38840,N_38744);
or U39064 (N_39064,N_38655,N_38697);
nor U39065 (N_39065,N_38646,N_38845);
nand U39066 (N_39066,N_38614,N_38686);
nor U39067 (N_39067,N_38605,N_38998);
and U39068 (N_39068,N_38772,N_38676);
or U39069 (N_39069,N_38650,N_38801);
xor U39070 (N_39070,N_38951,N_38991);
or U39071 (N_39071,N_38833,N_38548);
nor U39072 (N_39072,N_38785,N_38620);
or U39073 (N_39073,N_38981,N_38970);
or U39074 (N_39074,N_38708,N_38797);
nand U39075 (N_39075,N_38588,N_38959);
nor U39076 (N_39076,N_38626,N_38847);
xor U39077 (N_39077,N_38802,N_38679);
nand U39078 (N_39078,N_38592,N_38727);
and U39079 (N_39079,N_38822,N_38783);
nand U39080 (N_39080,N_38841,N_38642);
xnor U39081 (N_39081,N_38634,N_38952);
xnor U39082 (N_39082,N_38962,N_38759);
nor U39083 (N_39083,N_38560,N_38815);
xnor U39084 (N_39084,N_38529,N_38775);
and U39085 (N_39085,N_38762,N_38789);
or U39086 (N_39086,N_38788,N_38664);
xnor U39087 (N_39087,N_38591,N_38793);
or U39088 (N_39088,N_38858,N_38516);
nand U39089 (N_39089,N_38826,N_38810);
and U39090 (N_39090,N_38767,N_38522);
and U39091 (N_39091,N_38684,N_38880);
nand U39092 (N_39092,N_38930,N_38752);
nor U39093 (N_39093,N_38846,N_38798);
and U39094 (N_39094,N_38870,N_38773);
and U39095 (N_39095,N_38817,N_38928);
xor U39096 (N_39096,N_38640,N_38864);
nor U39097 (N_39097,N_38994,N_38597);
and U39098 (N_39098,N_38536,N_38663);
or U39099 (N_39099,N_38943,N_38891);
xor U39100 (N_39100,N_38944,N_38712);
or U39101 (N_39101,N_38791,N_38883);
and U39102 (N_39102,N_38972,N_38734);
xor U39103 (N_39103,N_38631,N_38748);
nand U39104 (N_39104,N_38662,N_38751);
nand U39105 (N_39105,N_38938,N_38904);
and U39106 (N_39106,N_38747,N_38933);
nand U39107 (N_39107,N_38570,N_38949);
nor U39108 (N_39108,N_38923,N_38926);
xor U39109 (N_39109,N_38639,N_38680);
xnor U39110 (N_39110,N_38549,N_38757);
nor U39111 (N_39111,N_38996,N_38863);
nand U39112 (N_39112,N_38984,N_38932);
and U39113 (N_39113,N_38630,N_38504);
and U39114 (N_39114,N_38704,N_38736);
nor U39115 (N_39115,N_38746,N_38920);
nand U39116 (N_39116,N_38877,N_38827);
nor U39117 (N_39117,N_38509,N_38743);
nand U39118 (N_39118,N_38940,N_38659);
nor U39119 (N_39119,N_38709,N_38603);
and U39120 (N_39120,N_38579,N_38527);
nor U39121 (N_39121,N_38755,N_38979);
and U39122 (N_39122,N_38553,N_38964);
nor U39123 (N_39123,N_38997,N_38590);
or U39124 (N_39124,N_38619,N_38975);
or U39125 (N_39125,N_38580,N_38902);
nor U39126 (N_39126,N_38728,N_38909);
or U39127 (N_39127,N_38986,N_38830);
nor U39128 (N_39128,N_38862,N_38644);
and U39129 (N_39129,N_38546,N_38988);
and U39130 (N_39130,N_38612,N_38599);
or U39131 (N_39131,N_38939,N_38719);
nor U39132 (N_39132,N_38912,N_38888);
and U39133 (N_39133,N_38871,N_38859);
nand U39134 (N_39134,N_38578,N_38837);
xnor U39135 (N_39135,N_38950,N_38918);
nand U39136 (N_39136,N_38628,N_38919);
xor U39137 (N_39137,N_38636,N_38978);
or U39138 (N_39138,N_38617,N_38738);
xor U39139 (N_39139,N_38764,N_38576);
or U39140 (N_39140,N_38956,N_38849);
nand U39141 (N_39141,N_38699,N_38724);
nand U39142 (N_39142,N_38530,N_38673);
xor U39143 (N_39143,N_38843,N_38989);
and U39144 (N_39144,N_38806,N_38867);
nor U39145 (N_39145,N_38749,N_38689);
nor U39146 (N_39146,N_38582,N_38790);
nor U39147 (N_39147,N_38539,N_38606);
or U39148 (N_39148,N_38672,N_38987);
and U39149 (N_39149,N_38819,N_38993);
nand U39150 (N_39150,N_38741,N_38635);
and U39151 (N_39151,N_38844,N_38915);
or U39152 (N_39152,N_38561,N_38584);
nor U39153 (N_39153,N_38675,N_38853);
nand U39154 (N_39154,N_38941,N_38911);
or U39155 (N_39155,N_38533,N_38716);
and U39156 (N_39156,N_38776,N_38929);
and U39157 (N_39157,N_38857,N_38971);
nand U39158 (N_39158,N_38782,N_38948);
xor U39159 (N_39159,N_38770,N_38542);
or U39160 (N_39160,N_38799,N_38677);
and U39161 (N_39161,N_38999,N_38607);
nor U39162 (N_39162,N_38992,N_38958);
xor U39163 (N_39163,N_38514,N_38688);
or U39164 (N_39164,N_38908,N_38627);
xnor U39165 (N_39165,N_38510,N_38980);
xor U39166 (N_39166,N_38598,N_38937);
nand U39167 (N_39167,N_38885,N_38985);
or U39168 (N_39168,N_38901,N_38832);
nor U39169 (N_39169,N_38691,N_38796);
nand U39170 (N_39170,N_38753,N_38889);
and U39171 (N_39171,N_38690,N_38874);
and U39172 (N_39172,N_38742,N_38519);
nand U39173 (N_39173,N_38625,N_38969);
xor U39174 (N_39174,N_38714,N_38872);
and U39175 (N_39175,N_38881,N_38769);
or U39176 (N_39176,N_38917,N_38760);
and U39177 (N_39177,N_38774,N_38693);
nand U39178 (N_39178,N_38563,N_38953);
nand U39179 (N_39179,N_38890,N_38502);
or U39180 (N_39180,N_38976,N_38503);
and U39181 (N_39181,N_38559,N_38869);
xnor U39182 (N_39182,N_38804,N_38558);
xnor U39183 (N_39183,N_38809,N_38713);
nand U39184 (N_39184,N_38887,N_38861);
or U39185 (N_39185,N_38906,N_38884);
or U39186 (N_39186,N_38766,N_38800);
xor U39187 (N_39187,N_38720,N_38795);
nor U39188 (N_39188,N_38629,N_38921);
xor U39189 (N_39189,N_38621,N_38882);
and U39190 (N_39190,N_38517,N_38641);
nand U39191 (N_39191,N_38886,N_38839);
or U39192 (N_39192,N_38556,N_38668);
xnor U39193 (N_39193,N_38860,N_38805);
or U39194 (N_39194,N_38816,N_38856);
nand U39195 (N_39195,N_38842,N_38572);
nor U39196 (N_39196,N_38750,N_38564);
xor U39197 (N_39197,N_38602,N_38540);
or U39198 (N_39198,N_38977,N_38851);
or U39199 (N_39199,N_38694,N_38945);
or U39200 (N_39200,N_38622,N_38946);
nor U39201 (N_39201,N_38660,N_38756);
and U39202 (N_39202,N_38850,N_38565);
nor U39203 (N_39203,N_38557,N_38550);
or U39204 (N_39204,N_38896,N_38544);
and U39205 (N_39205,N_38532,N_38735);
nor U39206 (N_39206,N_38595,N_38698);
and U39207 (N_39207,N_38965,N_38521);
nor U39208 (N_39208,N_38552,N_38610);
nor U39209 (N_39209,N_38705,N_38905);
nand U39210 (N_39210,N_38707,N_38925);
or U39211 (N_39211,N_38968,N_38873);
nand U39212 (N_39212,N_38615,N_38820);
or U39213 (N_39213,N_38934,N_38507);
nor U39214 (N_39214,N_38834,N_38731);
xor U39215 (N_39215,N_38567,N_38535);
xor U39216 (N_39216,N_38779,N_38649);
xnor U39217 (N_39217,N_38778,N_38737);
or U39218 (N_39218,N_38894,N_38600);
or U39219 (N_39219,N_38670,N_38900);
or U39220 (N_39220,N_38508,N_38512);
and U39221 (N_39221,N_38780,N_38703);
or U39222 (N_39222,N_38931,N_38566);
and U39223 (N_39223,N_38538,N_38808);
xnor U39224 (N_39224,N_38593,N_38569);
nand U39225 (N_39225,N_38711,N_38914);
or U39226 (N_39226,N_38879,N_38624);
nand U39227 (N_39227,N_38525,N_38609);
nor U39228 (N_39228,N_38601,N_38961);
and U39229 (N_39229,N_38581,N_38596);
or U39230 (N_39230,N_38825,N_38792);
nor U39231 (N_39231,N_38687,N_38898);
xor U39232 (N_39232,N_38718,N_38648);
xnor U39233 (N_39233,N_38974,N_38763);
xnor U39234 (N_39234,N_38554,N_38678);
nand U39235 (N_39235,N_38616,N_38551);
and U39236 (N_39236,N_38855,N_38706);
nor U39237 (N_39237,N_38674,N_38812);
nor U39238 (N_39238,N_38892,N_38823);
and U39239 (N_39239,N_38537,N_38722);
nor U39240 (N_39240,N_38666,N_38910);
xnor U39241 (N_39241,N_38701,N_38696);
or U39242 (N_39242,N_38836,N_38913);
and U39243 (N_39243,N_38829,N_38683);
nor U39244 (N_39244,N_38518,N_38824);
and U39245 (N_39245,N_38702,N_38637);
nand U39246 (N_39246,N_38916,N_38589);
nor U39247 (N_39247,N_38924,N_38777);
and U39248 (N_39248,N_38893,N_38895);
or U39249 (N_39249,N_38818,N_38821);
or U39250 (N_39250,N_38691,N_38632);
and U39251 (N_39251,N_38986,N_38679);
nand U39252 (N_39252,N_38746,N_38969);
xnor U39253 (N_39253,N_38908,N_38868);
and U39254 (N_39254,N_38646,N_38655);
nand U39255 (N_39255,N_38707,N_38966);
nor U39256 (N_39256,N_38889,N_38620);
xor U39257 (N_39257,N_38517,N_38664);
xnor U39258 (N_39258,N_38539,N_38952);
nand U39259 (N_39259,N_38663,N_38989);
and U39260 (N_39260,N_38669,N_38699);
xor U39261 (N_39261,N_38930,N_38883);
xnor U39262 (N_39262,N_38726,N_38723);
xnor U39263 (N_39263,N_38575,N_38731);
and U39264 (N_39264,N_38570,N_38990);
xnor U39265 (N_39265,N_38777,N_38565);
nor U39266 (N_39266,N_38962,N_38766);
and U39267 (N_39267,N_38941,N_38778);
xnor U39268 (N_39268,N_38503,N_38603);
or U39269 (N_39269,N_38839,N_38997);
nand U39270 (N_39270,N_38986,N_38853);
or U39271 (N_39271,N_38790,N_38672);
xor U39272 (N_39272,N_38893,N_38705);
and U39273 (N_39273,N_38939,N_38937);
xor U39274 (N_39274,N_38671,N_38905);
or U39275 (N_39275,N_38958,N_38965);
nand U39276 (N_39276,N_38763,N_38921);
and U39277 (N_39277,N_38749,N_38790);
nor U39278 (N_39278,N_38550,N_38660);
xnor U39279 (N_39279,N_38542,N_38604);
nand U39280 (N_39280,N_38619,N_38500);
xor U39281 (N_39281,N_38755,N_38562);
nor U39282 (N_39282,N_38538,N_38680);
and U39283 (N_39283,N_38692,N_38801);
xnor U39284 (N_39284,N_38985,N_38925);
or U39285 (N_39285,N_38874,N_38754);
and U39286 (N_39286,N_38594,N_38503);
and U39287 (N_39287,N_38835,N_38967);
nor U39288 (N_39288,N_38785,N_38871);
and U39289 (N_39289,N_38533,N_38849);
and U39290 (N_39290,N_38558,N_38622);
xor U39291 (N_39291,N_38802,N_38967);
and U39292 (N_39292,N_38687,N_38594);
xnor U39293 (N_39293,N_38907,N_38757);
nand U39294 (N_39294,N_38660,N_38759);
xor U39295 (N_39295,N_38805,N_38966);
or U39296 (N_39296,N_38605,N_38791);
nand U39297 (N_39297,N_38747,N_38581);
nand U39298 (N_39298,N_38545,N_38533);
or U39299 (N_39299,N_38603,N_38777);
or U39300 (N_39300,N_38978,N_38958);
nor U39301 (N_39301,N_38534,N_38685);
nor U39302 (N_39302,N_38861,N_38835);
nand U39303 (N_39303,N_38734,N_38994);
and U39304 (N_39304,N_38949,N_38700);
and U39305 (N_39305,N_38578,N_38777);
nand U39306 (N_39306,N_38500,N_38556);
xnor U39307 (N_39307,N_38801,N_38606);
xnor U39308 (N_39308,N_38962,N_38684);
nand U39309 (N_39309,N_38740,N_38683);
xnor U39310 (N_39310,N_38661,N_38931);
or U39311 (N_39311,N_38926,N_38876);
or U39312 (N_39312,N_38804,N_38983);
nor U39313 (N_39313,N_38636,N_38887);
nand U39314 (N_39314,N_38839,N_38699);
nor U39315 (N_39315,N_38912,N_38936);
and U39316 (N_39316,N_38766,N_38865);
nand U39317 (N_39317,N_38544,N_38832);
or U39318 (N_39318,N_38936,N_38690);
xnor U39319 (N_39319,N_38568,N_38794);
nor U39320 (N_39320,N_38962,N_38666);
or U39321 (N_39321,N_38583,N_38983);
xnor U39322 (N_39322,N_38554,N_38835);
xnor U39323 (N_39323,N_38636,N_38541);
or U39324 (N_39324,N_38719,N_38699);
nand U39325 (N_39325,N_38849,N_38794);
nand U39326 (N_39326,N_38729,N_38722);
and U39327 (N_39327,N_38816,N_38619);
xnor U39328 (N_39328,N_38510,N_38880);
nand U39329 (N_39329,N_38513,N_38504);
nor U39330 (N_39330,N_38837,N_38944);
xnor U39331 (N_39331,N_38709,N_38668);
nand U39332 (N_39332,N_38681,N_38635);
and U39333 (N_39333,N_38991,N_38618);
xor U39334 (N_39334,N_38638,N_38984);
nor U39335 (N_39335,N_38891,N_38683);
xor U39336 (N_39336,N_38699,N_38758);
nand U39337 (N_39337,N_38997,N_38828);
nand U39338 (N_39338,N_38677,N_38532);
nor U39339 (N_39339,N_38893,N_38583);
nor U39340 (N_39340,N_38657,N_38587);
and U39341 (N_39341,N_38677,N_38957);
or U39342 (N_39342,N_38921,N_38749);
or U39343 (N_39343,N_38803,N_38729);
nor U39344 (N_39344,N_38572,N_38795);
nor U39345 (N_39345,N_38879,N_38646);
nand U39346 (N_39346,N_38980,N_38602);
xor U39347 (N_39347,N_38562,N_38847);
xor U39348 (N_39348,N_38654,N_38633);
nand U39349 (N_39349,N_38843,N_38544);
nor U39350 (N_39350,N_38542,N_38703);
xor U39351 (N_39351,N_38852,N_38856);
nand U39352 (N_39352,N_38769,N_38800);
nand U39353 (N_39353,N_38737,N_38644);
and U39354 (N_39354,N_38872,N_38533);
and U39355 (N_39355,N_38973,N_38855);
xor U39356 (N_39356,N_38532,N_38934);
xor U39357 (N_39357,N_38644,N_38918);
and U39358 (N_39358,N_38881,N_38978);
nor U39359 (N_39359,N_38782,N_38887);
nor U39360 (N_39360,N_38661,N_38519);
nand U39361 (N_39361,N_38530,N_38757);
nor U39362 (N_39362,N_38681,N_38963);
nand U39363 (N_39363,N_38584,N_38571);
or U39364 (N_39364,N_38691,N_38621);
nand U39365 (N_39365,N_38844,N_38906);
xor U39366 (N_39366,N_38840,N_38681);
nand U39367 (N_39367,N_38893,N_38834);
and U39368 (N_39368,N_38924,N_38857);
or U39369 (N_39369,N_38609,N_38840);
nor U39370 (N_39370,N_38733,N_38570);
and U39371 (N_39371,N_38802,N_38652);
nand U39372 (N_39372,N_38987,N_38871);
and U39373 (N_39373,N_38867,N_38700);
and U39374 (N_39374,N_38693,N_38900);
nand U39375 (N_39375,N_38845,N_38815);
xor U39376 (N_39376,N_38931,N_38644);
and U39377 (N_39377,N_38645,N_38588);
nor U39378 (N_39378,N_38584,N_38995);
or U39379 (N_39379,N_38579,N_38997);
xnor U39380 (N_39380,N_38946,N_38978);
nor U39381 (N_39381,N_38925,N_38819);
and U39382 (N_39382,N_38826,N_38713);
and U39383 (N_39383,N_38617,N_38872);
or U39384 (N_39384,N_38528,N_38862);
nor U39385 (N_39385,N_38513,N_38609);
and U39386 (N_39386,N_38509,N_38956);
nand U39387 (N_39387,N_38815,N_38663);
and U39388 (N_39388,N_38518,N_38688);
or U39389 (N_39389,N_38938,N_38674);
xor U39390 (N_39390,N_38655,N_38807);
or U39391 (N_39391,N_38867,N_38776);
nand U39392 (N_39392,N_38847,N_38660);
and U39393 (N_39393,N_38839,N_38992);
and U39394 (N_39394,N_38870,N_38660);
nand U39395 (N_39395,N_38912,N_38849);
nor U39396 (N_39396,N_38559,N_38542);
and U39397 (N_39397,N_38676,N_38937);
and U39398 (N_39398,N_38751,N_38949);
xor U39399 (N_39399,N_38997,N_38674);
nor U39400 (N_39400,N_38694,N_38523);
and U39401 (N_39401,N_38514,N_38526);
nor U39402 (N_39402,N_38745,N_38656);
or U39403 (N_39403,N_38681,N_38524);
or U39404 (N_39404,N_38950,N_38778);
nor U39405 (N_39405,N_38598,N_38646);
and U39406 (N_39406,N_38621,N_38650);
xor U39407 (N_39407,N_38565,N_38544);
xnor U39408 (N_39408,N_38981,N_38703);
nor U39409 (N_39409,N_38823,N_38791);
xnor U39410 (N_39410,N_38956,N_38872);
nor U39411 (N_39411,N_38964,N_38520);
nor U39412 (N_39412,N_38917,N_38848);
xnor U39413 (N_39413,N_38751,N_38566);
nor U39414 (N_39414,N_38767,N_38836);
or U39415 (N_39415,N_38653,N_38612);
or U39416 (N_39416,N_38912,N_38827);
xnor U39417 (N_39417,N_38971,N_38510);
nor U39418 (N_39418,N_38783,N_38996);
and U39419 (N_39419,N_38804,N_38605);
xnor U39420 (N_39420,N_38834,N_38910);
nor U39421 (N_39421,N_38708,N_38605);
and U39422 (N_39422,N_38702,N_38560);
and U39423 (N_39423,N_38678,N_38906);
nand U39424 (N_39424,N_38773,N_38735);
nor U39425 (N_39425,N_38957,N_38530);
or U39426 (N_39426,N_38614,N_38668);
nor U39427 (N_39427,N_38505,N_38695);
or U39428 (N_39428,N_38733,N_38628);
and U39429 (N_39429,N_38507,N_38802);
nor U39430 (N_39430,N_38746,N_38855);
nor U39431 (N_39431,N_38866,N_38880);
or U39432 (N_39432,N_38646,N_38644);
xnor U39433 (N_39433,N_38556,N_38549);
nor U39434 (N_39434,N_38661,N_38827);
nor U39435 (N_39435,N_38659,N_38655);
or U39436 (N_39436,N_38503,N_38553);
and U39437 (N_39437,N_38594,N_38549);
nor U39438 (N_39438,N_38560,N_38801);
and U39439 (N_39439,N_38627,N_38999);
nor U39440 (N_39440,N_38940,N_38618);
xnor U39441 (N_39441,N_38552,N_38783);
or U39442 (N_39442,N_38988,N_38779);
or U39443 (N_39443,N_38540,N_38794);
nor U39444 (N_39444,N_38976,N_38890);
nand U39445 (N_39445,N_38971,N_38973);
and U39446 (N_39446,N_38988,N_38667);
or U39447 (N_39447,N_38953,N_38945);
or U39448 (N_39448,N_38935,N_38584);
and U39449 (N_39449,N_38519,N_38627);
xnor U39450 (N_39450,N_38953,N_38726);
or U39451 (N_39451,N_38607,N_38596);
and U39452 (N_39452,N_38643,N_38900);
xor U39453 (N_39453,N_38940,N_38742);
or U39454 (N_39454,N_38573,N_38665);
and U39455 (N_39455,N_38929,N_38660);
nand U39456 (N_39456,N_38891,N_38904);
nand U39457 (N_39457,N_38755,N_38943);
xnor U39458 (N_39458,N_38555,N_38830);
nand U39459 (N_39459,N_38657,N_38922);
and U39460 (N_39460,N_38753,N_38723);
xnor U39461 (N_39461,N_38744,N_38559);
xnor U39462 (N_39462,N_38509,N_38849);
xor U39463 (N_39463,N_38642,N_38705);
nor U39464 (N_39464,N_38741,N_38630);
nand U39465 (N_39465,N_38564,N_38752);
or U39466 (N_39466,N_38547,N_38538);
or U39467 (N_39467,N_38927,N_38613);
or U39468 (N_39468,N_38980,N_38938);
and U39469 (N_39469,N_38750,N_38733);
and U39470 (N_39470,N_38781,N_38867);
xor U39471 (N_39471,N_38677,N_38948);
nand U39472 (N_39472,N_38749,N_38682);
or U39473 (N_39473,N_38557,N_38772);
nand U39474 (N_39474,N_38753,N_38568);
and U39475 (N_39475,N_38758,N_38673);
or U39476 (N_39476,N_38504,N_38575);
nor U39477 (N_39477,N_38530,N_38658);
nor U39478 (N_39478,N_38933,N_38538);
nor U39479 (N_39479,N_38560,N_38545);
and U39480 (N_39480,N_38969,N_38530);
xnor U39481 (N_39481,N_38834,N_38757);
or U39482 (N_39482,N_38609,N_38689);
and U39483 (N_39483,N_38518,N_38900);
xnor U39484 (N_39484,N_38759,N_38769);
nand U39485 (N_39485,N_38789,N_38555);
or U39486 (N_39486,N_38529,N_38956);
xor U39487 (N_39487,N_38657,N_38863);
xnor U39488 (N_39488,N_38947,N_38625);
or U39489 (N_39489,N_38543,N_38919);
nand U39490 (N_39490,N_38858,N_38633);
or U39491 (N_39491,N_38792,N_38759);
and U39492 (N_39492,N_38857,N_38560);
or U39493 (N_39493,N_38959,N_38519);
xnor U39494 (N_39494,N_38626,N_38566);
nand U39495 (N_39495,N_38631,N_38763);
xnor U39496 (N_39496,N_38959,N_38556);
xor U39497 (N_39497,N_38576,N_38828);
and U39498 (N_39498,N_38753,N_38500);
and U39499 (N_39499,N_38784,N_38828);
or U39500 (N_39500,N_39485,N_39430);
nor U39501 (N_39501,N_39466,N_39183);
nand U39502 (N_39502,N_39453,N_39068);
or U39503 (N_39503,N_39058,N_39478);
and U39504 (N_39504,N_39147,N_39332);
and U39505 (N_39505,N_39310,N_39180);
nand U39506 (N_39506,N_39169,N_39009);
nand U39507 (N_39507,N_39461,N_39188);
nand U39508 (N_39508,N_39294,N_39110);
or U39509 (N_39509,N_39102,N_39146);
nand U39510 (N_39510,N_39120,N_39211);
or U39511 (N_39511,N_39353,N_39205);
xor U39512 (N_39512,N_39074,N_39412);
and U39513 (N_39513,N_39369,N_39459);
nor U39514 (N_39514,N_39383,N_39030);
nand U39515 (N_39515,N_39252,N_39326);
and U39516 (N_39516,N_39360,N_39100);
nor U39517 (N_39517,N_39214,N_39470);
nor U39518 (N_39518,N_39007,N_39056);
nor U39519 (N_39519,N_39389,N_39038);
nand U39520 (N_39520,N_39022,N_39278);
xnor U39521 (N_39521,N_39239,N_39143);
nor U39522 (N_39522,N_39439,N_39320);
nor U39523 (N_39523,N_39125,N_39443);
nand U39524 (N_39524,N_39241,N_39329);
xor U39525 (N_39525,N_39077,N_39219);
xor U39526 (N_39526,N_39254,N_39157);
nand U39527 (N_39527,N_39233,N_39108);
nor U39528 (N_39528,N_39053,N_39171);
or U39529 (N_39529,N_39235,N_39000);
nor U39530 (N_39530,N_39119,N_39282);
nand U39531 (N_39531,N_39323,N_39398);
and U39532 (N_39532,N_39008,N_39473);
xnor U39533 (N_39533,N_39153,N_39006);
nand U39534 (N_39534,N_39250,N_39274);
nand U39535 (N_39535,N_39105,N_39440);
and U39536 (N_39536,N_39315,N_39139);
nand U39537 (N_39537,N_39213,N_39085);
or U39538 (N_39538,N_39054,N_39465);
or U39539 (N_39539,N_39408,N_39240);
xnor U39540 (N_39540,N_39474,N_39341);
nand U39541 (N_39541,N_39346,N_39327);
xor U39542 (N_39542,N_39452,N_39215);
or U39543 (N_39543,N_39486,N_39162);
nand U39544 (N_39544,N_39044,N_39194);
nand U39545 (N_39545,N_39028,N_39417);
and U39546 (N_39546,N_39073,N_39457);
and U39547 (N_39547,N_39142,N_39446);
xnor U39548 (N_39548,N_39161,N_39178);
nand U39549 (N_39549,N_39218,N_39268);
or U39550 (N_39550,N_39377,N_39356);
nor U39551 (N_39551,N_39024,N_39127);
nand U39552 (N_39552,N_39176,N_39472);
nand U39553 (N_39553,N_39445,N_39265);
nand U39554 (N_39554,N_39303,N_39253);
nand U39555 (N_39555,N_39003,N_39225);
nand U39556 (N_39556,N_39281,N_39476);
nand U39557 (N_39557,N_39393,N_39331);
and U39558 (N_39558,N_39086,N_39092);
and U39559 (N_39559,N_39104,N_39358);
nor U39560 (N_39560,N_39229,N_39141);
nor U39561 (N_39561,N_39078,N_39450);
nand U39562 (N_39562,N_39454,N_39222);
or U39563 (N_39563,N_39113,N_39001);
nor U39564 (N_39564,N_39067,N_39135);
nor U39565 (N_39565,N_39313,N_39002);
xnor U39566 (N_39566,N_39349,N_39492);
and U39567 (N_39567,N_39340,N_39280);
or U39568 (N_39568,N_39469,N_39390);
nor U39569 (N_39569,N_39374,N_39101);
nor U39570 (N_39570,N_39495,N_39015);
xor U39571 (N_39571,N_39145,N_39283);
nand U39572 (N_39572,N_39165,N_39122);
and U39573 (N_39573,N_39080,N_39043);
nand U39574 (N_39574,N_39410,N_39375);
xor U39575 (N_39575,N_39425,N_39487);
and U39576 (N_39576,N_39350,N_39150);
xor U39577 (N_39577,N_39034,N_39447);
xnor U39578 (N_39578,N_39304,N_39031);
and U39579 (N_39579,N_39202,N_39126);
nand U39580 (N_39580,N_39246,N_39091);
or U39581 (N_39581,N_39255,N_39232);
and U39582 (N_39582,N_39103,N_39048);
and U39583 (N_39583,N_39491,N_39267);
xnor U39584 (N_39584,N_39168,N_39464);
and U39585 (N_39585,N_39012,N_39134);
nand U39586 (N_39586,N_39394,N_39065);
xnor U39587 (N_39587,N_39471,N_39039);
nor U39588 (N_39588,N_39387,N_39160);
xor U39589 (N_39589,N_39373,N_39212);
nand U39590 (N_39590,N_39223,N_39385);
nor U39591 (N_39591,N_39069,N_39115);
and U39592 (N_39592,N_39025,N_39249);
and U39593 (N_39593,N_39409,N_39499);
xnor U39594 (N_39594,N_39462,N_39449);
or U39595 (N_39595,N_39489,N_39203);
or U39596 (N_39596,N_39033,N_39285);
xor U39597 (N_39597,N_39455,N_39192);
nor U39598 (N_39598,N_39224,N_39437);
xor U39599 (N_39599,N_39338,N_39251);
or U39600 (N_39600,N_39128,N_39075);
nor U39601 (N_39601,N_39070,N_39339);
or U39602 (N_39602,N_39302,N_39010);
or U39603 (N_39603,N_39089,N_39289);
or U39604 (N_39604,N_39190,N_39081);
and U39605 (N_39605,N_39016,N_39264);
or U39606 (N_39606,N_39245,N_39426);
nor U39607 (N_39607,N_39296,N_39291);
or U39608 (N_39608,N_39483,N_39045);
xor U39609 (N_39609,N_39191,N_39221);
nand U39610 (N_39610,N_39413,N_39272);
and U39611 (N_39611,N_39336,N_39234);
nor U39612 (N_39612,N_39121,N_39328);
nor U39613 (N_39613,N_39481,N_39170);
nor U39614 (N_39614,N_39064,N_39076);
and U39615 (N_39615,N_39114,N_39405);
xnor U39616 (N_39616,N_39484,N_39419);
nor U39617 (N_39617,N_39456,N_39384);
nor U39618 (N_39618,N_39181,N_39388);
and U39619 (N_39619,N_39248,N_39309);
nand U39620 (N_39620,N_39227,N_39208);
or U39621 (N_39621,N_39163,N_39187);
xnor U39622 (N_39622,N_39036,N_39293);
xnor U39623 (N_39623,N_39014,N_39195);
or U39624 (N_39624,N_39386,N_39316);
xnor U39625 (N_39625,N_39244,N_39279);
nand U39626 (N_39626,N_39155,N_39111);
or U39627 (N_39627,N_39441,N_39175);
and U39628 (N_39628,N_39396,N_39347);
or U39629 (N_39629,N_39357,N_39217);
nor U39630 (N_39630,N_39460,N_39026);
nor U39631 (N_39631,N_39037,N_39324);
xor U39632 (N_39632,N_39082,N_39432);
nor U39633 (N_39633,N_39206,N_39062);
nand U39634 (N_39634,N_39050,N_39395);
nand U39635 (N_39635,N_39237,N_39429);
xnor U39636 (N_39636,N_39379,N_39260);
nor U39637 (N_39637,N_39005,N_39345);
xor U39638 (N_39638,N_39365,N_39173);
and U39639 (N_39639,N_39403,N_39311);
or U39640 (N_39640,N_39414,N_39094);
and U39641 (N_39641,N_39059,N_39342);
or U39642 (N_39642,N_39061,N_39090);
or U39643 (N_39643,N_39148,N_39368);
xor U39644 (N_39644,N_39020,N_39318);
or U39645 (N_39645,N_39416,N_39262);
nor U39646 (N_39646,N_39186,N_39182);
or U39647 (N_39647,N_39266,N_39494);
nor U39648 (N_39648,N_39210,N_39431);
xor U39649 (N_39649,N_39297,N_39072);
or U39650 (N_39650,N_39133,N_39438);
nand U39651 (N_39651,N_39199,N_39164);
nand U39652 (N_39652,N_39138,N_39354);
and U39653 (N_39653,N_39193,N_39172);
nor U39654 (N_39654,N_39132,N_39201);
xnor U39655 (N_39655,N_39179,N_39325);
xor U39656 (N_39656,N_39391,N_39256);
nor U39657 (N_39657,N_39372,N_39238);
nand U39658 (N_39658,N_39380,N_39004);
and U39659 (N_39659,N_39051,N_39301);
xnor U39660 (N_39660,N_39079,N_39381);
nand U39661 (N_39661,N_39314,N_39017);
nor U39662 (N_39662,N_39402,N_39433);
nor U39663 (N_39663,N_39047,N_39436);
xnor U39664 (N_39664,N_39019,N_39243);
nor U39665 (N_39665,N_39124,N_39415);
nand U39666 (N_39666,N_39231,N_39158);
and U39667 (N_39667,N_39493,N_39144);
xnor U39668 (N_39668,N_39099,N_39063);
and U39669 (N_39669,N_39228,N_39344);
nor U39670 (N_39670,N_39216,N_39434);
xor U39671 (N_39671,N_39035,N_39442);
or U39672 (N_39672,N_39378,N_39189);
xnor U39673 (N_39673,N_39361,N_39088);
xnor U39674 (N_39674,N_39392,N_39458);
nand U39675 (N_39675,N_39400,N_39397);
xor U39676 (N_39676,N_39055,N_39337);
nor U39677 (N_39677,N_39488,N_39166);
nor U39678 (N_39678,N_39348,N_39174);
nor U39679 (N_39679,N_39209,N_39330);
nand U39680 (N_39680,N_39040,N_39448);
and U39681 (N_39681,N_39367,N_39107);
or U39682 (N_39682,N_39137,N_39322);
nor U39683 (N_39683,N_39355,N_39376);
or U39684 (N_39684,N_39129,N_39087);
or U39685 (N_39685,N_39236,N_39098);
nand U39686 (N_39686,N_39247,N_39286);
and U39687 (N_39687,N_39066,N_39042);
xnor U39688 (N_39688,N_39185,N_39288);
nand U39689 (N_39689,N_39154,N_39423);
nor U39690 (N_39690,N_39299,N_39230);
and U39691 (N_39691,N_39156,N_39277);
and U39692 (N_39692,N_39451,N_39307);
xnor U39693 (N_39693,N_39273,N_39352);
or U39694 (N_39694,N_39497,N_39343);
nor U39695 (N_39695,N_39287,N_39371);
nor U39696 (N_39696,N_39200,N_39422);
nand U39697 (N_39697,N_39084,N_39317);
nand U39698 (N_39698,N_39490,N_39312);
and U39699 (N_39699,N_39083,N_39226);
nand U39700 (N_39700,N_39196,N_39300);
nor U39701 (N_39701,N_39270,N_39276);
nor U39702 (N_39702,N_39151,N_39421);
nor U39703 (N_39703,N_39284,N_39177);
and U39704 (N_39704,N_39136,N_39306);
nor U39705 (N_39705,N_39401,N_39334);
or U39706 (N_39706,N_39399,N_39032);
or U39707 (N_39707,N_39305,N_39427);
xnor U39708 (N_39708,N_39428,N_39112);
xnor U39709 (N_39709,N_39435,N_39052);
and U39710 (N_39710,N_39149,N_39468);
xnor U39711 (N_39711,N_39258,N_39463);
nand U39712 (N_39712,N_39496,N_39475);
or U39713 (N_39713,N_39424,N_39308);
nand U39714 (N_39714,N_39366,N_39018);
xnor U39715 (N_39715,N_39290,N_39096);
nor U39716 (N_39716,N_39027,N_39097);
nand U39717 (N_39717,N_39140,N_39498);
nand U39718 (N_39718,N_39482,N_39152);
and U39719 (N_39719,N_39444,N_39116);
nor U39720 (N_39720,N_39013,N_39411);
or U39721 (N_39721,N_39407,N_39333);
xnor U39722 (N_39722,N_39167,N_39404);
and U39723 (N_39723,N_39118,N_39257);
xnor U39724 (N_39724,N_39321,N_39242);
xor U39725 (N_39725,N_39131,N_39095);
or U39726 (N_39726,N_39319,N_39220);
and U39727 (N_39727,N_39480,N_39359);
or U39728 (N_39728,N_39159,N_39362);
xnor U39729 (N_39729,N_39269,N_39011);
or U39730 (N_39730,N_39049,N_39420);
and U39731 (N_39731,N_39335,N_39041);
or U39732 (N_39732,N_39271,N_39261);
nand U39733 (N_39733,N_39263,N_39479);
nand U39734 (N_39734,N_39023,N_39117);
nor U39735 (N_39735,N_39071,N_39363);
xnor U39736 (N_39736,N_39198,N_39130);
nor U39737 (N_39737,N_39123,N_39295);
nand U39738 (N_39738,N_39207,N_39259);
nor U39739 (N_39739,N_39109,N_39057);
nand U39740 (N_39740,N_39298,N_39382);
or U39741 (N_39741,N_39351,N_39364);
nand U39742 (N_39742,N_39477,N_39418);
nand U39743 (N_39743,N_39184,N_39204);
and U39744 (N_39744,N_39197,N_39467);
nor U39745 (N_39745,N_39275,N_39021);
nor U39746 (N_39746,N_39093,N_39060);
nor U39747 (N_39747,N_39029,N_39406);
or U39748 (N_39748,N_39292,N_39106);
nand U39749 (N_39749,N_39370,N_39046);
or U39750 (N_39750,N_39339,N_39143);
xnor U39751 (N_39751,N_39459,N_39367);
nor U39752 (N_39752,N_39297,N_39065);
xnor U39753 (N_39753,N_39157,N_39416);
xor U39754 (N_39754,N_39310,N_39083);
nor U39755 (N_39755,N_39406,N_39395);
nand U39756 (N_39756,N_39390,N_39283);
xor U39757 (N_39757,N_39469,N_39314);
or U39758 (N_39758,N_39430,N_39203);
or U39759 (N_39759,N_39079,N_39277);
and U39760 (N_39760,N_39321,N_39241);
xnor U39761 (N_39761,N_39342,N_39366);
xnor U39762 (N_39762,N_39276,N_39499);
and U39763 (N_39763,N_39055,N_39053);
nor U39764 (N_39764,N_39423,N_39100);
xor U39765 (N_39765,N_39293,N_39042);
or U39766 (N_39766,N_39341,N_39498);
or U39767 (N_39767,N_39433,N_39308);
nor U39768 (N_39768,N_39004,N_39330);
and U39769 (N_39769,N_39099,N_39339);
or U39770 (N_39770,N_39151,N_39316);
nor U39771 (N_39771,N_39304,N_39135);
nor U39772 (N_39772,N_39142,N_39108);
and U39773 (N_39773,N_39342,N_39221);
and U39774 (N_39774,N_39446,N_39105);
nand U39775 (N_39775,N_39179,N_39067);
nand U39776 (N_39776,N_39392,N_39188);
or U39777 (N_39777,N_39325,N_39357);
xor U39778 (N_39778,N_39137,N_39453);
xor U39779 (N_39779,N_39467,N_39407);
xnor U39780 (N_39780,N_39044,N_39172);
nand U39781 (N_39781,N_39185,N_39010);
nand U39782 (N_39782,N_39168,N_39009);
and U39783 (N_39783,N_39227,N_39258);
or U39784 (N_39784,N_39071,N_39139);
nand U39785 (N_39785,N_39448,N_39211);
nand U39786 (N_39786,N_39244,N_39424);
nor U39787 (N_39787,N_39373,N_39237);
nor U39788 (N_39788,N_39116,N_39382);
and U39789 (N_39789,N_39069,N_39268);
nor U39790 (N_39790,N_39305,N_39128);
nand U39791 (N_39791,N_39127,N_39438);
or U39792 (N_39792,N_39480,N_39167);
nand U39793 (N_39793,N_39229,N_39207);
or U39794 (N_39794,N_39461,N_39230);
nor U39795 (N_39795,N_39461,N_39217);
and U39796 (N_39796,N_39133,N_39066);
nand U39797 (N_39797,N_39095,N_39430);
xnor U39798 (N_39798,N_39091,N_39425);
and U39799 (N_39799,N_39456,N_39201);
nand U39800 (N_39800,N_39390,N_39322);
xor U39801 (N_39801,N_39294,N_39027);
xor U39802 (N_39802,N_39294,N_39295);
nand U39803 (N_39803,N_39321,N_39499);
xor U39804 (N_39804,N_39047,N_39140);
nor U39805 (N_39805,N_39071,N_39276);
or U39806 (N_39806,N_39088,N_39357);
and U39807 (N_39807,N_39456,N_39052);
xnor U39808 (N_39808,N_39130,N_39025);
nor U39809 (N_39809,N_39445,N_39495);
nor U39810 (N_39810,N_39240,N_39303);
nor U39811 (N_39811,N_39152,N_39381);
nand U39812 (N_39812,N_39150,N_39187);
nand U39813 (N_39813,N_39161,N_39121);
xnor U39814 (N_39814,N_39133,N_39328);
and U39815 (N_39815,N_39420,N_39143);
nor U39816 (N_39816,N_39074,N_39076);
xor U39817 (N_39817,N_39038,N_39396);
xor U39818 (N_39818,N_39128,N_39078);
nand U39819 (N_39819,N_39181,N_39351);
and U39820 (N_39820,N_39110,N_39331);
or U39821 (N_39821,N_39001,N_39094);
nand U39822 (N_39822,N_39326,N_39048);
xor U39823 (N_39823,N_39018,N_39066);
and U39824 (N_39824,N_39097,N_39044);
nor U39825 (N_39825,N_39091,N_39272);
and U39826 (N_39826,N_39122,N_39207);
and U39827 (N_39827,N_39061,N_39049);
nor U39828 (N_39828,N_39276,N_39430);
or U39829 (N_39829,N_39215,N_39062);
nand U39830 (N_39830,N_39055,N_39227);
and U39831 (N_39831,N_39161,N_39077);
and U39832 (N_39832,N_39393,N_39013);
and U39833 (N_39833,N_39409,N_39495);
nand U39834 (N_39834,N_39486,N_39102);
and U39835 (N_39835,N_39317,N_39215);
xor U39836 (N_39836,N_39490,N_39111);
nor U39837 (N_39837,N_39471,N_39092);
xnor U39838 (N_39838,N_39497,N_39429);
nor U39839 (N_39839,N_39266,N_39371);
and U39840 (N_39840,N_39011,N_39359);
and U39841 (N_39841,N_39446,N_39234);
nor U39842 (N_39842,N_39492,N_39303);
nand U39843 (N_39843,N_39142,N_39060);
and U39844 (N_39844,N_39382,N_39195);
or U39845 (N_39845,N_39088,N_39180);
or U39846 (N_39846,N_39115,N_39026);
xor U39847 (N_39847,N_39473,N_39255);
nor U39848 (N_39848,N_39005,N_39253);
xor U39849 (N_39849,N_39255,N_39182);
nor U39850 (N_39850,N_39349,N_39108);
nand U39851 (N_39851,N_39058,N_39051);
and U39852 (N_39852,N_39153,N_39459);
nand U39853 (N_39853,N_39278,N_39267);
nand U39854 (N_39854,N_39135,N_39258);
nand U39855 (N_39855,N_39040,N_39303);
nor U39856 (N_39856,N_39096,N_39110);
nor U39857 (N_39857,N_39187,N_39406);
or U39858 (N_39858,N_39256,N_39091);
or U39859 (N_39859,N_39292,N_39259);
or U39860 (N_39860,N_39006,N_39275);
and U39861 (N_39861,N_39483,N_39034);
nor U39862 (N_39862,N_39319,N_39217);
and U39863 (N_39863,N_39001,N_39260);
and U39864 (N_39864,N_39369,N_39463);
or U39865 (N_39865,N_39295,N_39458);
nand U39866 (N_39866,N_39173,N_39371);
and U39867 (N_39867,N_39121,N_39454);
xnor U39868 (N_39868,N_39475,N_39186);
xor U39869 (N_39869,N_39072,N_39188);
nand U39870 (N_39870,N_39315,N_39016);
xor U39871 (N_39871,N_39155,N_39377);
nor U39872 (N_39872,N_39164,N_39204);
xnor U39873 (N_39873,N_39028,N_39301);
xnor U39874 (N_39874,N_39251,N_39180);
xnor U39875 (N_39875,N_39200,N_39447);
nor U39876 (N_39876,N_39062,N_39069);
nand U39877 (N_39877,N_39126,N_39137);
xor U39878 (N_39878,N_39238,N_39345);
and U39879 (N_39879,N_39365,N_39033);
and U39880 (N_39880,N_39105,N_39186);
or U39881 (N_39881,N_39224,N_39337);
or U39882 (N_39882,N_39226,N_39229);
nand U39883 (N_39883,N_39442,N_39436);
or U39884 (N_39884,N_39279,N_39218);
xnor U39885 (N_39885,N_39026,N_39092);
nor U39886 (N_39886,N_39045,N_39230);
or U39887 (N_39887,N_39261,N_39027);
xor U39888 (N_39888,N_39445,N_39163);
nand U39889 (N_39889,N_39122,N_39195);
or U39890 (N_39890,N_39033,N_39353);
nor U39891 (N_39891,N_39328,N_39315);
xor U39892 (N_39892,N_39461,N_39394);
or U39893 (N_39893,N_39299,N_39371);
xor U39894 (N_39894,N_39462,N_39340);
and U39895 (N_39895,N_39386,N_39411);
nand U39896 (N_39896,N_39088,N_39339);
xor U39897 (N_39897,N_39032,N_39022);
xor U39898 (N_39898,N_39185,N_39032);
xnor U39899 (N_39899,N_39144,N_39171);
nand U39900 (N_39900,N_39185,N_39127);
and U39901 (N_39901,N_39023,N_39150);
nand U39902 (N_39902,N_39074,N_39113);
or U39903 (N_39903,N_39333,N_39450);
xor U39904 (N_39904,N_39188,N_39423);
nand U39905 (N_39905,N_39084,N_39135);
nand U39906 (N_39906,N_39393,N_39330);
nand U39907 (N_39907,N_39461,N_39119);
and U39908 (N_39908,N_39223,N_39368);
nor U39909 (N_39909,N_39068,N_39129);
nand U39910 (N_39910,N_39010,N_39023);
xnor U39911 (N_39911,N_39317,N_39001);
xnor U39912 (N_39912,N_39422,N_39291);
nand U39913 (N_39913,N_39171,N_39157);
xor U39914 (N_39914,N_39089,N_39048);
or U39915 (N_39915,N_39222,N_39479);
nor U39916 (N_39916,N_39268,N_39015);
nand U39917 (N_39917,N_39488,N_39268);
and U39918 (N_39918,N_39448,N_39280);
nor U39919 (N_39919,N_39489,N_39046);
nand U39920 (N_39920,N_39217,N_39029);
nand U39921 (N_39921,N_39266,N_39100);
nor U39922 (N_39922,N_39274,N_39095);
nand U39923 (N_39923,N_39100,N_39180);
and U39924 (N_39924,N_39025,N_39419);
and U39925 (N_39925,N_39290,N_39389);
xor U39926 (N_39926,N_39371,N_39435);
or U39927 (N_39927,N_39499,N_39272);
and U39928 (N_39928,N_39446,N_39223);
or U39929 (N_39929,N_39136,N_39409);
and U39930 (N_39930,N_39219,N_39037);
nor U39931 (N_39931,N_39255,N_39262);
or U39932 (N_39932,N_39407,N_39038);
nand U39933 (N_39933,N_39136,N_39440);
and U39934 (N_39934,N_39319,N_39083);
or U39935 (N_39935,N_39195,N_39219);
nand U39936 (N_39936,N_39203,N_39282);
or U39937 (N_39937,N_39421,N_39417);
xnor U39938 (N_39938,N_39180,N_39073);
nand U39939 (N_39939,N_39227,N_39174);
or U39940 (N_39940,N_39028,N_39109);
nand U39941 (N_39941,N_39192,N_39055);
nand U39942 (N_39942,N_39022,N_39468);
nand U39943 (N_39943,N_39301,N_39365);
xor U39944 (N_39944,N_39262,N_39026);
nor U39945 (N_39945,N_39106,N_39126);
xor U39946 (N_39946,N_39147,N_39379);
or U39947 (N_39947,N_39200,N_39255);
nor U39948 (N_39948,N_39061,N_39079);
xor U39949 (N_39949,N_39225,N_39107);
or U39950 (N_39950,N_39313,N_39040);
and U39951 (N_39951,N_39096,N_39363);
nor U39952 (N_39952,N_39381,N_39380);
nor U39953 (N_39953,N_39348,N_39116);
xor U39954 (N_39954,N_39396,N_39324);
nand U39955 (N_39955,N_39456,N_39444);
and U39956 (N_39956,N_39247,N_39191);
and U39957 (N_39957,N_39201,N_39285);
nand U39958 (N_39958,N_39118,N_39281);
or U39959 (N_39959,N_39459,N_39058);
xnor U39960 (N_39960,N_39199,N_39033);
nor U39961 (N_39961,N_39304,N_39263);
nor U39962 (N_39962,N_39128,N_39472);
nand U39963 (N_39963,N_39043,N_39115);
nand U39964 (N_39964,N_39139,N_39372);
nand U39965 (N_39965,N_39382,N_39371);
nor U39966 (N_39966,N_39216,N_39214);
and U39967 (N_39967,N_39217,N_39033);
nand U39968 (N_39968,N_39126,N_39120);
nor U39969 (N_39969,N_39408,N_39048);
nor U39970 (N_39970,N_39431,N_39125);
or U39971 (N_39971,N_39385,N_39117);
xnor U39972 (N_39972,N_39460,N_39034);
nand U39973 (N_39973,N_39211,N_39355);
or U39974 (N_39974,N_39478,N_39493);
nor U39975 (N_39975,N_39067,N_39292);
and U39976 (N_39976,N_39059,N_39141);
nor U39977 (N_39977,N_39351,N_39129);
or U39978 (N_39978,N_39414,N_39152);
nor U39979 (N_39979,N_39248,N_39283);
and U39980 (N_39980,N_39012,N_39089);
nor U39981 (N_39981,N_39323,N_39397);
nand U39982 (N_39982,N_39144,N_39176);
and U39983 (N_39983,N_39336,N_39227);
and U39984 (N_39984,N_39197,N_39108);
nand U39985 (N_39985,N_39023,N_39206);
or U39986 (N_39986,N_39302,N_39113);
and U39987 (N_39987,N_39384,N_39029);
or U39988 (N_39988,N_39041,N_39444);
nor U39989 (N_39989,N_39096,N_39464);
or U39990 (N_39990,N_39412,N_39449);
or U39991 (N_39991,N_39324,N_39033);
nor U39992 (N_39992,N_39398,N_39187);
nand U39993 (N_39993,N_39175,N_39116);
nand U39994 (N_39994,N_39016,N_39342);
and U39995 (N_39995,N_39178,N_39244);
xnor U39996 (N_39996,N_39085,N_39110);
or U39997 (N_39997,N_39161,N_39071);
or U39998 (N_39998,N_39179,N_39152);
or U39999 (N_39999,N_39255,N_39269);
and U40000 (N_40000,N_39855,N_39812);
nand U40001 (N_40001,N_39981,N_39880);
nor U40002 (N_40002,N_39518,N_39945);
nand U40003 (N_40003,N_39608,N_39811);
nand U40004 (N_40004,N_39602,N_39976);
nor U40005 (N_40005,N_39515,N_39962);
nand U40006 (N_40006,N_39785,N_39511);
and U40007 (N_40007,N_39825,N_39618);
or U40008 (N_40008,N_39826,N_39556);
or U40009 (N_40009,N_39600,N_39992);
nand U40010 (N_40010,N_39781,N_39660);
nand U40011 (N_40011,N_39776,N_39978);
nand U40012 (N_40012,N_39847,N_39928);
or U40013 (N_40013,N_39589,N_39920);
and U40014 (N_40014,N_39873,N_39703);
nand U40015 (N_40015,N_39995,N_39576);
or U40016 (N_40016,N_39539,N_39744);
or U40017 (N_40017,N_39846,N_39930);
or U40018 (N_40018,N_39712,N_39590);
and U40019 (N_40019,N_39698,N_39527);
or U40020 (N_40020,N_39676,N_39742);
nand U40021 (N_40021,N_39876,N_39998);
nand U40022 (N_40022,N_39691,N_39609);
nor U40023 (N_40023,N_39782,N_39655);
and U40024 (N_40024,N_39854,N_39759);
and U40025 (N_40025,N_39637,N_39516);
nor U40026 (N_40026,N_39977,N_39874);
nor U40027 (N_40027,N_39708,N_39794);
or U40028 (N_40028,N_39633,N_39500);
xnor U40029 (N_40029,N_39842,N_39840);
nand U40030 (N_40030,N_39533,N_39619);
nand U40031 (N_40031,N_39634,N_39766);
nand U40032 (N_40032,N_39603,N_39592);
nor U40033 (N_40033,N_39764,N_39886);
and U40034 (N_40034,N_39683,N_39700);
nand U40035 (N_40035,N_39587,N_39643);
xnor U40036 (N_40036,N_39843,N_39582);
and U40037 (N_40037,N_39925,N_39865);
nor U40038 (N_40038,N_39557,N_39724);
nor U40039 (N_40039,N_39638,N_39627);
xor U40040 (N_40040,N_39620,N_39960);
and U40041 (N_40041,N_39508,N_39635);
nor U40042 (N_40042,N_39631,N_39917);
or U40043 (N_40043,N_39974,N_39561);
nor U40044 (N_40044,N_39733,N_39520);
and U40045 (N_40045,N_39999,N_39911);
and U40046 (N_40046,N_39957,N_39816);
and U40047 (N_40047,N_39517,N_39975);
nand U40048 (N_40048,N_39571,N_39991);
nor U40049 (N_40049,N_39778,N_39612);
nand U40050 (N_40050,N_39573,N_39552);
xnor U40051 (N_40051,N_39659,N_39726);
nand U40052 (N_40052,N_39509,N_39697);
nor U40053 (N_40053,N_39687,N_39615);
xnor U40054 (N_40054,N_39820,N_39929);
or U40055 (N_40055,N_39786,N_39554);
or U40056 (N_40056,N_39530,N_39649);
and U40057 (N_40057,N_39809,N_39597);
xnor U40058 (N_40058,N_39662,N_39829);
nand U40059 (N_40059,N_39896,N_39982);
nand U40060 (N_40060,N_39755,N_39535);
nor U40061 (N_40061,N_39803,N_39885);
or U40062 (N_40062,N_39679,N_39965);
xor U40063 (N_40063,N_39636,N_39952);
or U40064 (N_40064,N_39707,N_39891);
and U40065 (N_40065,N_39625,N_39828);
nand U40066 (N_40066,N_39948,N_39719);
xor U40067 (N_40067,N_39705,N_39756);
xor U40068 (N_40068,N_39601,N_39706);
or U40069 (N_40069,N_39946,N_39875);
or U40070 (N_40070,N_39933,N_39950);
or U40071 (N_40071,N_39585,N_39939);
and U40072 (N_40072,N_39598,N_39839);
xor U40073 (N_40073,N_39848,N_39758);
and U40074 (N_40074,N_39654,N_39806);
nor U40075 (N_40075,N_39797,N_39640);
nor U40076 (N_40076,N_39593,N_39963);
and U40077 (N_40077,N_39834,N_39578);
and U40078 (N_40078,N_39793,N_39727);
xor U40079 (N_40079,N_39969,N_39681);
nor U40080 (N_40080,N_39558,N_39837);
nand U40081 (N_40081,N_39941,N_39728);
nand U40082 (N_40082,N_39947,N_39575);
nand U40083 (N_40083,N_39753,N_39818);
nor U40084 (N_40084,N_39872,N_39729);
nand U40085 (N_40085,N_39967,N_39888);
nand U40086 (N_40086,N_39532,N_39606);
nor U40087 (N_40087,N_39616,N_39682);
nand U40088 (N_40088,N_39833,N_39749);
nand U40089 (N_40089,N_39802,N_39762);
and U40090 (N_40090,N_39718,N_39892);
nand U40091 (N_40091,N_39584,N_39746);
nor U40092 (N_40092,N_39966,N_39912);
and U40093 (N_40093,N_39689,N_39628);
nor U40094 (N_40094,N_39990,N_39979);
xnor U40095 (N_40095,N_39559,N_39717);
nand U40096 (N_40096,N_39835,N_39993);
nand U40097 (N_40097,N_39611,N_39823);
xnor U40098 (N_40098,N_39548,N_39672);
and U40099 (N_40099,N_39959,N_39522);
and U40100 (N_40100,N_39506,N_39798);
nor U40101 (N_40101,N_39866,N_39827);
and U40102 (N_40102,N_39629,N_39537);
xor U40103 (N_40103,N_39821,N_39883);
and U40104 (N_40104,N_39736,N_39772);
and U40105 (N_40105,N_39968,N_39581);
nor U40106 (N_40106,N_39543,N_39890);
nand U40107 (N_40107,N_39622,N_39881);
nor U40108 (N_40108,N_39723,N_39800);
and U40109 (N_40109,N_39791,N_39650);
xnor U40110 (N_40110,N_39770,N_39735);
nand U40111 (N_40111,N_39599,N_39651);
nand U40112 (N_40112,N_39645,N_39997);
xnor U40113 (N_40113,N_39961,N_39653);
and U40114 (N_40114,N_39531,N_39524);
xnor U40115 (N_40115,N_39862,N_39754);
xor U40116 (N_40116,N_39505,N_39594);
xor U40117 (N_40117,N_39512,N_39956);
nor U40118 (N_40118,N_39663,N_39868);
nand U40119 (N_40119,N_39910,N_39652);
and U40120 (N_40120,N_39757,N_39893);
nand U40121 (N_40121,N_39536,N_39796);
and U40122 (N_40122,N_39894,N_39869);
and U40123 (N_40123,N_39924,N_39503);
and U40124 (N_40124,N_39824,N_39591);
xnor U40125 (N_40125,N_39788,N_39739);
nor U40126 (N_40126,N_39692,N_39669);
or U40127 (N_40127,N_39784,N_39607);
xor U40128 (N_40128,N_39921,N_39546);
and U40129 (N_40129,N_39942,N_39605);
nor U40130 (N_40130,N_39570,N_39549);
and U40131 (N_40131,N_39748,N_39579);
or U40132 (N_40132,N_39765,N_39918);
or U40133 (N_40133,N_39678,N_39715);
and U40134 (N_40134,N_39519,N_39617);
or U40135 (N_40135,N_39937,N_39808);
xnor U40136 (N_40136,N_39819,N_39673);
nand U40137 (N_40137,N_39664,N_39630);
xnor U40138 (N_40138,N_39523,N_39560);
and U40139 (N_40139,N_39752,N_39830);
nor U40140 (N_40140,N_39882,N_39804);
xnor U40141 (N_40141,N_39879,N_39773);
xnor U40142 (N_40142,N_39667,N_39714);
or U40143 (N_40143,N_39538,N_39988);
nand U40144 (N_40144,N_39996,N_39904);
and U40145 (N_40145,N_39905,N_39934);
xor U40146 (N_40146,N_39908,N_39780);
nor U40147 (N_40147,N_39926,N_39774);
nor U40148 (N_40148,N_39731,N_39913);
and U40149 (N_40149,N_39940,N_39850);
and U40150 (N_40150,N_39747,N_39973);
xnor U40151 (N_40151,N_39701,N_39613);
and U40152 (N_40152,N_39761,N_39877);
or U40153 (N_40153,N_39565,N_39716);
and U40154 (N_40154,N_39648,N_39887);
or U40155 (N_40155,N_39684,N_39895);
nand U40156 (N_40156,N_39938,N_39971);
and U40157 (N_40157,N_39621,N_39562);
nor U40158 (N_40158,N_39871,N_39639);
and U40159 (N_40159,N_39657,N_39771);
nand U40160 (N_40160,N_39721,N_39529);
xor U40161 (N_40161,N_39553,N_39685);
and U40162 (N_40162,N_39641,N_39951);
nand U40163 (N_40163,N_39709,N_39884);
and U40164 (N_40164,N_39586,N_39743);
xnor U40165 (N_40165,N_39914,N_39859);
nor U40166 (N_40166,N_39994,N_39935);
nand U40167 (N_40167,N_39710,N_39722);
and U40168 (N_40168,N_39514,N_39738);
nand U40169 (N_40169,N_39547,N_39838);
nor U40170 (N_40170,N_39661,N_39943);
nor U40171 (N_40171,N_39916,N_39769);
and U40172 (N_40172,N_39900,N_39521);
and U40173 (N_40173,N_39949,N_39856);
xor U40174 (N_40174,N_39550,N_39671);
and U40175 (N_40175,N_39695,N_39642);
and U40176 (N_40176,N_39541,N_39668);
nand U40177 (N_40177,N_39767,N_39675);
or U40178 (N_40178,N_39899,N_39566);
or U40179 (N_40179,N_39987,N_39870);
nand U40180 (N_40180,N_39725,N_39790);
nand U40181 (N_40181,N_39944,N_39763);
nor U40182 (N_40182,N_39544,N_39775);
nor U40183 (N_40183,N_39955,N_39588);
and U40184 (N_40184,N_39972,N_39779);
or U40185 (N_40185,N_39568,N_39953);
nand U40186 (N_40186,N_39693,N_39583);
nor U40187 (N_40187,N_39732,N_39632);
nand U40188 (N_40188,N_39989,N_39958);
xor U40189 (N_40189,N_39907,N_39898);
xor U40190 (N_40190,N_39574,N_39670);
nand U40191 (N_40191,N_39909,N_39572);
and U40192 (N_40192,N_39787,N_39936);
xnor U40193 (N_40193,N_39624,N_39688);
xor U40194 (N_40194,N_39915,N_39551);
nand U40195 (N_40195,N_39507,N_39813);
nor U40196 (N_40196,N_39555,N_39919);
xnor U40197 (N_40197,N_39677,N_39832);
nand U40198 (N_40198,N_39903,N_39923);
xor U40199 (N_40199,N_39985,N_39751);
or U40200 (N_40200,N_39858,N_39694);
and U40201 (N_40201,N_39504,N_39542);
and U40202 (N_40202,N_39852,N_39502);
nand U40203 (N_40203,N_39932,N_39696);
nand U40204 (N_40204,N_39704,N_39792);
xnor U40205 (N_40205,N_39831,N_39970);
nand U40206 (N_40206,N_39906,N_39902);
or U40207 (N_40207,N_39801,N_39604);
or U40208 (N_40208,N_39844,N_39931);
nor U40209 (N_40209,N_39730,N_39577);
and U40210 (N_40210,N_39836,N_39863);
or U40211 (N_40211,N_39644,N_39646);
and U40212 (N_40212,N_39534,N_39674);
or U40213 (N_40213,N_39861,N_39889);
nor U40214 (N_40214,N_39680,N_39986);
nand U40215 (N_40215,N_39768,N_39815);
and U40216 (N_40216,N_39851,N_39822);
nand U40217 (N_40217,N_39927,N_39737);
and U40218 (N_40218,N_39658,N_39745);
or U40219 (N_40219,N_39878,N_39528);
xnor U40220 (N_40220,N_39720,N_39795);
or U40221 (N_40221,N_39596,N_39510);
xor U40222 (N_40222,N_39741,N_39540);
and U40223 (N_40223,N_39580,N_39841);
nand U40224 (N_40224,N_39760,N_39980);
xnor U40225 (N_40225,N_39814,N_39713);
and U40226 (N_40226,N_39545,N_39799);
xnor U40227 (N_40227,N_39860,N_39805);
and U40228 (N_40228,N_39563,N_39954);
nand U40229 (N_40229,N_39789,N_39783);
and U40230 (N_40230,N_39853,N_39922);
xnor U40231 (N_40231,N_39983,N_39626);
or U40232 (N_40232,N_39513,N_39807);
or U40233 (N_40233,N_39690,N_39564);
nor U40234 (N_40234,N_39817,N_39845);
or U40235 (N_40235,N_39699,N_39864);
and U40236 (N_40236,N_39964,N_39623);
nand U40237 (N_40237,N_39686,N_39867);
xor U40238 (N_40238,N_39525,N_39897);
and U40239 (N_40239,N_39702,N_39610);
or U40240 (N_40240,N_39656,N_39734);
nand U40241 (N_40241,N_39595,N_39666);
or U40242 (N_40242,N_39567,N_39849);
nand U40243 (N_40243,N_39526,N_39711);
and U40244 (N_40244,N_39569,N_39647);
and U40245 (N_40245,N_39740,N_39750);
or U40246 (N_40246,N_39857,N_39777);
nand U40247 (N_40247,N_39614,N_39665);
or U40248 (N_40248,N_39984,N_39901);
xor U40249 (N_40249,N_39810,N_39501);
nor U40250 (N_40250,N_39941,N_39666);
nand U40251 (N_40251,N_39907,N_39771);
xnor U40252 (N_40252,N_39543,N_39760);
nand U40253 (N_40253,N_39620,N_39775);
and U40254 (N_40254,N_39711,N_39730);
nand U40255 (N_40255,N_39502,N_39607);
and U40256 (N_40256,N_39903,N_39691);
xnor U40257 (N_40257,N_39936,N_39946);
or U40258 (N_40258,N_39803,N_39892);
and U40259 (N_40259,N_39598,N_39508);
nor U40260 (N_40260,N_39843,N_39891);
and U40261 (N_40261,N_39633,N_39725);
xnor U40262 (N_40262,N_39710,N_39956);
nor U40263 (N_40263,N_39879,N_39828);
nand U40264 (N_40264,N_39551,N_39503);
and U40265 (N_40265,N_39518,N_39556);
xor U40266 (N_40266,N_39817,N_39508);
or U40267 (N_40267,N_39974,N_39746);
and U40268 (N_40268,N_39813,N_39831);
and U40269 (N_40269,N_39962,N_39756);
or U40270 (N_40270,N_39507,N_39632);
nand U40271 (N_40271,N_39725,N_39537);
nor U40272 (N_40272,N_39862,N_39829);
xnor U40273 (N_40273,N_39538,N_39717);
xnor U40274 (N_40274,N_39593,N_39607);
nand U40275 (N_40275,N_39677,N_39986);
nor U40276 (N_40276,N_39910,N_39684);
or U40277 (N_40277,N_39840,N_39985);
xor U40278 (N_40278,N_39528,N_39509);
xnor U40279 (N_40279,N_39700,N_39592);
nor U40280 (N_40280,N_39577,N_39742);
or U40281 (N_40281,N_39753,N_39950);
nor U40282 (N_40282,N_39545,N_39709);
nand U40283 (N_40283,N_39696,N_39955);
or U40284 (N_40284,N_39903,N_39801);
and U40285 (N_40285,N_39984,N_39576);
nor U40286 (N_40286,N_39852,N_39860);
nand U40287 (N_40287,N_39979,N_39501);
and U40288 (N_40288,N_39685,N_39793);
xnor U40289 (N_40289,N_39942,N_39764);
xor U40290 (N_40290,N_39912,N_39908);
nor U40291 (N_40291,N_39749,N_39511);
nor U40292 (N_40292,N_39910,N_39560);
and U40293 (N_40293,N_39557,N_39824);
nand U40294 (N_40294,N_39736,N_39954);
nand U40295 (N_40295,N_39975,N_39630);
and U40296 (N_40296,N_39508,N_39892);
nor U40297 (N_40297,N_39582,N_39661);
nor U40298 (N_40298,N_39715,N_39531);
nor U40299 (N_40299,N_39889,N_39746);
and U40300 (N_40300,N_39561,N_39609);
nand U40301 (N_40301,N_39830,N_39834);
and U40302 (N_40302,N_39716,N_39888);
xnor U40303 (N_40303,N_39964,N_39822);
nor U40304 (N_40304,N_39713,N_39890);
or U40305 (N_40305,N_39731,N_39820);
nor U40306 (N_40306,N_39770,N_39920);
or U40307 (N_40307,N_39505,N_39882);
nor U40308 (N_40308,N_39986,N_39918);
nor U40309 (N_40309,N_39636,N_39889);
and U40310 (N_40310,N_39829,N_39905);
or U40311 (N_40311,N_39899,N_39731);
nor U40312 (N_40312,N_39574,N_39745);
nor U40313 (N_40313,N_39983,N_39529);
or U40314 (N_40314,N_39975,N_39670);
and U40315 (N_40315,N_39513,N_39733);
nor U40316 (N_40316,N_39921,N_39804);
nand U40317 (N_40317,N_39627,N_39753);
nand U40318 (N_40318,N_39855,N_39785);
or U40319 (N_40319,N_39621,N_39767);
nor U40320 (N_40320,N_39518,N_39740);
nand U40321 (N_40321,N_39557,N_39889);
or U40322 (N_40322,N_39528,N_39653);
nor U40323 (N_40323,N_39791,N_39665);
nand U40324 (N_40324,N_39875,N_39786);
nor U40325 (N_40325,N_39749,N_39577);
xnor U40326 (N_40326,N_39970,N_39721);
nor U40327 (N_40327,N_39806,N_39968);
or U40328 (N_40328,N_39639,N_39957);
nor U40329 (N_40329,N_39550,N_39548);
xor U40330 (N_40330,N_39563,N_39920);
xor U40331 (N_40331,N_39548,N_39539);
xor U40332 (N_40332,N_39892,N_39514);
and U40333 (N_40333,N_39980,N_39755);
nand U40334 (N_40334,N_39560,N_39921);
xnor U40335 (N_40335,N_39892,N_39532);
nor U40336 (N_40336,N_39538,N_39591);
nor U40337 (N_40337,N_39960,N_39593);
nand U40338 (N_40338,N_39722,N_39925);
and U40339 (N_40339,N_39584,N_39878);
or U40340 (N_40340,N_39603,N_39892);
nand U40341 (N_40341,N_39727,N_39879);
xnor U40342 (N_40342,N_39916,N_39823);
and U40343 (N_40343,N_39639,N_39733);
xnor U40344 (N_40344,N_39511,N_39737);
or U40345 (N_40345,N_39953,N_39582);
or U40346 (N_40346,N_39872,N_39752);
and U40347 (N_40347,N_39708,N_39756);
xnor U40348 (N_40348,N_39911,N_39592);
nor U40349 (N_40349,N_39834,N_39533);
and U40350 (N_40350,N_39616,N_39760);
nand U40351 (N_40351,N_39549,N_39943);
nor U40352 (N_40352,N_39948,N_39914);
or U40353 (N_40353,N_39543,N_39910);
nor U40354 (N_40354,N_39690,N_39718);
nand U40355 (N_40355,N_39623,N_39694);
nor U40356 (N_40356,N_39684,N_39699);
xnor U40357 (N_40357,N_39551,N_39959);
and U40358 (N_40358,N_39923,N_39754);
or U40359 (N_40359,N_39748,N_39845);
nand U40360 (N_40360,N_39996,N_39565);
and U40361 (N_40361,N_39880,N_39863);
and U40362 (N_40362,N_39992,N_39888);
nand U40363 (N_40363,N_39567,N_39503);
or U40364 (N_40364,N_39568,N_39535);
nor U40365 (N_40365,N_39520,N_39822);
or U40366 (N_40366,N_39511,N_39950);
nor U40367 (N_40367,N_39937,N_39719);
xor U40368 (N_40368,N_39924,N_39956);
or U40369 (N_40369,N_39654,N_39904);
xnor U40370 (N_40370,N_39763,N_39997);
and U40371 (N_40371,N_39566,N_39980);
nor U40372 (N_40372,N_39986,N_39600);
and U40373 (N_40373,N_39592,N_39957);
nand U40374 (N_40374,N_39529,N_39972);
nand U40375 (N_40375,N_39980,N_39875);
nand U40376 (N_40376,N_39552,N_39989);
nor U40377 (N_40377,N_39824,N_39634);
and U40378 (N_40378,N_39966,N_39725);
xor U40379 (N_40379,N_39996,N_39827);
nand U40380 (N_40380,N_39557,N_39926);
xnor U40381 (N_40381,N_39609,N_39725);
nand U40382 (N_40382,N_39743,N_39730);
nand U40383 (N_40383,N_39847,N_39792);
nor U40384 (N_40384,N_39654,N_39651);
nor U40385 (N_40385,N_39548,N_39937);
or U40386 (N_40386,N_39655,N_39558);
nor U40387 (N_40387,N_39683,N_39582);
nand U40388 (N_40388,N_39964,N_39647);
nand U40389 (N_40389,N_39505,N_39620);
nand U40390 (N_40390,N_39521,N_39941);
xnor U40391 (N_40391,N_39582,N_39949);
nand U40392 (N_40392,N_39580,N_39582);
nand U40393 (N_40393,N_39839,N_39801);
xor U40394 (N_40394,N_39567,N_39937);
xor U40395 (N_40395,N_39627,N_39876);
xor U40396 (N_40396,N_39863,N_39937);
or U40397 (N_40397,N_39776,N_39802);
and U40398 (N_40398,N_39922,N_39803);
xor U40399 (N_40399,N_39690,N_39796);
nand U40400 (N_40400,N_39735,N_39976);
nor U40401 (N_40401,N_39843,N_39868);
xnor U40402 (N_40402,N_39713,N_39505);
nor U40403 (N_40403,N_39586,N_39527);
nor U40404 (N_40404,N_39678,N_39611);
nor U40405 (N_40405,N_39816,N_39510);
or U40406 (N_40406,N_39603,N_39625);
or U40407 (N_40407,N_39684,N_39601);
nor U40408 (N_40408,N_39753,N_39709);
nand U40409 (N_40409,N_39737,N_39972);
and U40410 (N_40410,N_39614,N_39679);
and U40411 (N_40411,N_39505,N_39888);
nand U40412 (N_40412,N_39581,N_39634);
or U40413 (N_40413,N_39685,N_39822);
nand U40414 (N_40414,N_39550,N_39801);
nand U40415 (N_40415,N_39991,N_39563);
nor U40416 (N_40416,N_39948,N_39814);
nor U40417 (N_40417,N_39541,N_39532);
or U40418 (N_40418,N_39919,N_39979);
nor U40419 (N_40419,N_39974,N_39999);
nand U40420 (N_40420,N_39976,N_39801);
or U40421 (N_40421,N_39533,N_39876);
nand U40422 (N_40422,N_39703,N_39568);
nand U40423 (N_40423,N_39618,N_39688);
xnor U40424 (N_40424,N_39673,N_39514);
nand U40425 (N_40425,N_39848,N_39992);
nand U40426 (N_40426,N_39842,N_39779);
or U40427 (N_40427,N_39680,N_39866);
nand U40428 (N_40428,N_39821,N_39699);
xor U40429 (N_40429,N_39890,N_39714);
nand U40430 (N_40430,N_39577,N_39752);
nand U40431 (N_40431,N_39699,N_39651);
nor U40432 (N_40432,N_39925,N_39679);
nor U40433 (N_40433,N_39524,N_39758);
nand U40434 (N_40434,N_39642,N_39843);
xor U40435 (N_40435,N_39749,N_39625);
xnor U40436 (N_40436,N_39721,N_39611);
xor U40437 (N_40437,N_39929,N_39623);
and U40438 (N_40438,N_39991,N_39548);
and U40439 (N_40439,N_39585,N_39691);
xnor U40440 (N_40440,N_39625,N_39501);
xor U40441 (N_40441,N_39906,N_39969);
or U40442 (N_40442,N_39979,N_39997);
xor U40443 (N_40443,N_39592,N_39609);
and U40444 (N_40444,N_39818,N_39585);
xnor U40445 (N_40445,N_39715,N_39961);
or U40446 (N_40446,N_39807,N_39838);
and U40447 (N_40447,N_39884,N_39804);
xor U40448 (N_40448,N_39974,N_39868);
nor U40449 (N_40449,N_39820,N_39610);
xor U40450 (N_40450,N_39925,N_39520);
xor U40451 (N_40451,N_39890,N_39886);
or U40452 (N_40452,N_39761,N_39729);
and U40453 (N_40453,N_39861,N_39749);
nor U40454 (N_40454,N_39705,N_39872);
and U40455 (N_40455,N_39844,N_39801);
nor U40456 (N_40456,N_39516,N_39963);
and U40457 (N_40457,N_39984,N_39701);
nor U40458 (N_40458,N_39620,N_39752);
xor U40459 (N_40459,N_39528,N_39968);
nand U40460 (N_40460,N_39522,N_39678);
or U40461 (N_40461,N_39602,N_39988);
xor U40462 (N_40462,N_39803,N_39535);
nand U40463 (N_40463,N_39840,N_39785);
xnor U40464 (N_40464,N_39644,N_39696);
nand U40465 (N_40465,N_39703,N_39569);
or U40466 (N_40466,N_39883,N_39871);
nor U40467 (N_40467,N_39760,N_39598);
nand U40468 (N_40468,N_39816,N_39929);
and U40469 (N_40469,N_39531,N_39870);
xor U40470 (N_40470,N_39999,N_39843);
nor U40471 (N_40471,N_39850,N_39973);
or U40472 (N_40472,N_39733,N_39666);
nor U40473 (N_40473,N_39665,N_39913);
nand U40474 (N_40474,N_39695,N_39821);
nand U40475 (N_40475,N_39715,N_39914);
xor U40476 (N_40476,N_39522,N_39535);
nor U40477 (N_40477,N_39785,N_39775);
and U40478 (N_40478,N_39871,N_39535);
and U40479 (N_40479,N_39646,N_39893);
nor U40480 (N_40480,N_39987,N_39931);
nor U40481 (N_40481,N_39957,N_39682);
nand U40482 (N_40482,N_39657,N_39849);
and U40483 (N_40483,N_39709,N_39636);
xor U40484 (N_40484,N_39927,N_39719);
and U40485 (N_40485,N_39581,N_39944);
or U40486 (N_40486,N_39771,N_39631);
or U40487 (N_40487,N_39989,N_39561);
xnor U40488 (N_40488,N_39810,N_39870);
and U40489 (N_40489,N_39603,N_39917);
and U40490 (N_40490,N_39923,N_39936);
and U40491 (N_40491,N_39984,N_39822);
xnor U40492 (N_40492,N_39955,N_39737);
xor U40493 (N_40493,N_39806,N_39843);
nand U40494 (N_40494,N_39909,N_39599);
xor U40495 (N_40495,N_39949,N_39779);
nor U40496 (N_40496,N_39517,N_39952);
or U40497 (N_40497,N_39731,N_39586);
nand U40498 (N_40498,N_39506,N_39737);
or U40499 (N_40499,N_39692,N_39993);
and U40500 (N_40500,N_40164,N_40180);
or U40501 (N_40501,N_40388,N_40458);
xor U40502 (N_40502,N_40283,N_40234);
nand U40503 (N_40503,N_40034,N_40364);
nand U40504 (N_40504,N_40319,N_40462);
nand U40505 (N_40505,N_40113,N_40246);
nor U40506 (N_40506,N_40482,N_40201);
nand U40507 (N_40507,N_40263,N_40274);
nand U40508 (N_40508,N_40367,N_40424);
nor U40509 (N_40509,N_40259,N_40317);
nand U40510 (N_40510,N_40225,N_40257);
nand U40511 (N_40511,N_40476,N_40243);
xnor U40512 (N_40512,N_40249,N_40146);
nor U40513 (N_40513,N_40419,N_40278);
xnor U40514 (N_40514,N_40035,N_40298);
or U40515 (N_40515,N_40383,N_40357);
nand U40516 (N_40516,N_40245,N_40079);
or U40517 (N_40517,N_40374,N_40229);
and U40518 (N_40518,N_40491,N_40067);
nor U40519 (N_40519,N_40227,N_40108);
and U40520 (N_40520,N_40276,N_40461);
or U40521 (N_40521,N_40255,N_40161);
and U40522 (N_40522,N_40405,N_40314);
and U40523 (N_40523,N_40203,N_40185);
or U40524 (N_40524,N_40187,N_40421);
and U40525 (N_40525,N_40474,N_40100);
and U40526 (N_40526,N_40358,N_40495);
and U40527 (N_40527,N_40432,N_40214);
nand U40528 (N_40528,N_40007,N_40463);
or U40529 (N_40529,N_40157,N_40247);
nand U40530 (N_40530,N_40331,N_40332);
nand U40531 (N_40531,N_40305,N_40075);
or U40532 (N_40532,N_40097,N_40215);
or U40533 (N_40533,N_40196,N_40231);
nand U40534 (N_40534,N_40111,N_40488);
xor U40535 (N_40535,N_40415,N_40397);
nand U40536 (N_40536,N_40381,N_40320);
xnor U40537 (N_40537,N_40178,N_40375);
xor U40538 (N_40538,N_40147,N_40114);
or U40539 (N_40539,N_40135,N_40430);
nor U40540 (N_40540,N_40412,N_40418);
nand U40541 (N_40541,N_40233,N_40059);
nand U40542 (N_40542,N_40083,N_40384);
nor U40543 (N_40543,N_40359,N_40428);
and U40544 (N_40544,N_40264,N_40173);
and U40545 (N_40545,N_40466,N_40343);
nor U40546 (N_40546,N_40094,N_40478);
nor U40547 (N_40547,N_40315,N_40254);
nor U40548 (N_40548,N_40148,N_40139);
nor U40549 (N_40549,N_40363,N_40289);
or U40550 (N_40550,N_40177,N_40217);
or U40551 (N_40551,N_40029,N_40369);
nand U40552 (N_40552,N_40209,N_40226);
nand U40553 (N_40553,N_40301,N_40268);
xor U40554 (N_40554,N_40133,N_40292);
nand U40555 (N_40555,N_40069,N_40248);
xnor U40556 (N_40556,N_40390,N_40436);
xor U40557 (N_40557,N_40077,N_40013);
nand U40558 (N_40558,N_40055,N_40475);
and U40559 (N_40559,N_40408,N_40334);
nor U40560 (N_40560,N_40160,N_40449);
nand U40561 (N_40561,N_40356,N_40239);
nor U40562 (N_40562,N_40081,N_40186);
nor U40563 (N_40563,N_40130,N_40445);
or U40564 (N_40564,N_40211,N_40000);
nand U40565 (N_40565,N_40306,N_40310);
xor U40566 (N_40566,N_40071,N_40240);
and U40567 (N_40567,N_40096,N_40103);
or U40568 (N_40568,N_40342,N_40095);
nor U40569 (N_40569,N_40413,N_40460);
xnor U40570 (N_40570,N_40321,N_40167);
xnor U40571 (N_40571,N_40107,N_40435);
or U40572 (N_40572,N_40145,N_40382);
nor U40573 (N_40573,N_40191,N_40399);
and U40574 (N_40574,N_40499,N_40008);
nand U40575 (N_40575,N_40417,N_40426);
or U40576 (N_40576,N_40250,N_40377);
xnor U40577 (N_40577,N_40032,N_40026);
xor U40578 (N_40578,N_40308,N_40414);
xor U40579 (N_40579,N_40294,N_40004);
nor U40580 (N_40580,N_40024,N_40093);
and U40581 (N_40581,N_40447,N_40483);
or U40582 (N_40582,N_40101,N_40425);
and U40583 (N_40583,N_40181,N_40057);
or U40584 (N_40584,N_40464,N_40080);
and U40585 (N_40585,N_40400,N_40339);
and U40586 (N_40586,N_40385,N_40162);
nand U40587 (N_40587,N_40170,N_40354);
nor U40588 (N_40588,N_40090,N_40485);
and U40589 (N_40589,N_40442,N_40043);
nand U40590 (N_40590,N_40338,N_40070);
xor U40591 (N_40591,N_40251,N_40403);
or U40592 (N_40592,N_40282,N_40056);
and U40593 (N_40593,N_40228,N_40312);
or U40594 (N_40594,N_40378,N_40365);
or U40595 (N_40595,N_40453,N_40015);
or U40596 (N_40596,N_40150,N_40344);
nand U40597 (N_40597,N_40110,N_40340);
xor U40598 (N_40598,N_40052,N_40376);
nor U40599 (N_40599,N_40126,N_40038);
nor U40600 (N_40600,N_40444,N_40119);
nor U40601 (N_40601,N_40309,N_40362);
or U40602 (N_40602,N_40207,N_40153);
nor U40603 (N_40603,N_40063,N_40115);
xor U40604 (N_40604,N_40188,N_40109);
xnor U40605 (N_40605,N_40204,N_40280);
or U40606 (N_40606,N_40102,N_40064);
xnor U40607 (N_40607,N_40333,N_40218);
or U40608 (N_40608,N_40323,N_40456);
and U40609 (N_40609,N_40129,N_40267);
or U40610 (N_40610,N_40244,N_40302);
and U40611 (N_40611,N_40222,N_40434);
and U40612 (N_40612,N_40065,N_40172);
and U40613 (N_40613,N_40144,N_40237);
nor U40614 (N_40614,N_40446,N_40346);
and U40615 (N_40615,N_40001,N_40492);
and U40616 (N_40616,N_40422,N_40078);
nor U40617 (N_40617,N_40465,N_40051);
nor U40618 (N_40618,N_40467,N_40060);
or U40619 (N_40619,N_40036,N_40118);
and U40620 (N_40620,N_40195,N_40206);
nand U40621 (N_40621,N_40355,N_40149);
xor U40622 (N_40622,N_40014,N_40041);
and U40623 (N_40623,N_40290,N_40262);
and U40624 (N_40624,N_40140,N_40406);
nor U40625 (N_40625,N_40299,N_40479);
xor U40626 (N_40626,N_40137,N_40128);
xor U40627 (N_40627,N_40353,N_40285);
nor U40628 (N_40628,N_40493,N_40045);
or U40629 (N_40629,N_40325,N_40189);
xnor U40630 (N_40630,N_40404,N_40028);
nand U40631 (N_40631,N_40471,N_40288);
nand U40632 (N_40632,N_40303,N_40120);
and U40633 (N_40633,N_40368,N_40392);
and U40634 (N_40634,N_40098,N_40345);
and U40635 (N_40635,N_40198,N_40125);
or U40636 (N_40636,N_40387,N_40341);
and U40637 (N_40637,N_40272,N_40054);
or U40638 (N_40638,N_40158,N_40131);
and U40639 (N_40639,N_40494,N_40042);
xnor U40640 (N_40640,N_40061,N_40469);
nand U40641 (N_40641,N_40104,N_40473);
or U40642 (N_40642,N_40123,N_40027);
and U40643 (N_40643,N_40087,N_40010);
or U40644 (N_40644,N_40261,N_40448);
nand U40645 (N_40645,N_40210,N_40112);
and U40646 (N_40646,N_40219,N_40452);
nor U40647 (N_40647,N_40124,N_40277);
or U40648 (N_40648,N_40266,N_40171);
xor U40649 (N_40649,N_40213,N_40242);
nand U40650 (N_40650,N_40197,N_40295);
nand U40651 (N_40651,N_40260,N_40351);
or U40652 (N_40652,N_40361,N_40179);
nor U40653 (N_40653,N_40006,N_40440);
and U40654 (N_40654,N_40327,N_40286);
and U40655 (N_40655,N_40450,N_40402);
nand U40656 (N_40656,N_40304,N_40481);
xor U40657 (N_40657,N_40088,N_40205);
nor U40658 (N_40658,N_40194,N_40165);
and U40659 (N_40659,N_40349,N_40062);
xor U40660 (N_40660,N_40132,N_40127);
nor U40661 (N_40661,N_40105,N_40275);
or U40662 (N_40662,N_40287,N_40050);
nand U40663 (N_40663,N_40151,N_40166);
and U40664 (N_40664,N_40053,N_40011);
and U40665 (N_40665,N_40241,N_40136);
xor U40666 (N_40666,N_40037,N_40238);
and U40667 (N_40667,N_40313,N_40373);
nor U40668 (N_40668,N_40371,N_40138);
nor U40669 (N_40669,N_40152,N_40370);
or U40670 (N_40670,N_40270,N_40386);
nor U40671 (N_40671,N_40086,N_40183);
or U40672 (N_40672,N_40352,N_40085);
xor U40673 (N_40673,N_40389,N_40427);
nor U40674 (N_40674,N_40416,N_40159);
xor U40675 (N_40675,N_40017,N_40141);
xnor U40676 (N_40676,N_40033,N_40269);
and U40677 (N_40677,N_40019,N_40429);
and U40678 (N_40678,N_40143,N_40433);
nor U40679 (N_40679,N_40468,N_40438);
or U40680 (N_40680,N_40224,N_40092);
xor U40681 (N_40681,N_40220,N_40184);
nand U40682 (N_40682,N_40082,N_40208);
nor U40683 (N_40683,N_40066,N_40284);
nor U40684 (N_40684,N_40300,N_40047);
or U40685 (N_40685,N_40044,N_40009);
and U40686 (N_40686,N_40169,N_40230);
nor U40687 (N_40687,N_40122,N_40484);
and U40688 (N_40688,N_40336,N_40048);
or U40689 (N_40689,N_40003,N_40279);
or U40690 (N_40690,N_40020,N_40423);
xor U40691 (N_40691,N_40040,N_40350);
or U40692 (N_40692,N_40487,N_40311);
nor U40693 (N_40693,N_40497,N_40223);
or U40694 (N_40694,N_40410,N_40407);
and U40695 (N_40695,N_40023,N_40457);
nor U40696 (N_40696,N_40271,N_40089);
nand U40697 (N_40697,N_40182,N_40021);
nor U40698 (N_40698,N_40372,N_40074);
xnor U40699 (N_40699,N_40200,N_40121);
nand U40700 (N_40700,N_40437,N_40459);
nand U40701 (N_40701,N_40393,N_40199);
nand U40702 (N_40702,N_40411,N_40221);
or U40703 (N_40703,N_40176,N_40324);
nor U40704 (N_40704,N_40046,N_40072);
or U40705 (N_40705,N_40163,N_40232);
nand U40706 (N_40706,N_40281,N_40273);
or U40707 (N_40707,N_40409,N_40058);
and U40708 (N_40708,N_40498,N_40455);
xor U40709 (N_40709,N_40431,N_40134);
xor U40710 (N_40710,N_40016,N_40477);
or U40711 (N_40711,N_40451,N_40439);
or U40712 (N_40712,N_40252,N_40192);
or U40713 (N_40713,N_40293,N_40401);
or U40714 (N_40714,N_40335,N_40005);
nor U40715 (N_40715,N_40307,N_40031);
nand U40716 (N_40716,N_40049,N_40175);
nand U40717 (N_40717,N_40099,N_40391);
xor U40718 (N_40718,N_40329,N_40454);
nand U40719 (N_40719,N_40420,N_40330);
and U40720 (N_40720,N_40348,N_40360);
xor U40721 (N_40721,N_40084,N_40328);
or U40722 (N_40722,N_40470,N_40398);
or U40723 (N_40723,N_40396,N_40174);
nand U40724 (N_40724,N_40337,N_40472);
xnor U40725 (N_40725,N_40030,N_40366);
nor U40726 (N_40726,N_40073,N_40297);
nand U40727 (N_40727,N_40216,N_40106);
xnor U40728 (N_40728,N_40116,N_40142);
or U40729 (N_40729,N_40236,N_40394);
nor U40730 (N_40730,N_40265,N_40022);
xor U40731 (N_40731,N_40322,N_40316);
and U40732 (N_40732,N_40202,N_40291);
nor U40733 (N_40733,N_40318,N_40490);
nor U40734 (N_40734,N_40091,N_40155);
nor U40735 (N_40735,N_40486,N_40256);
and U40736 (N_40736,N_40156,N_40039);
nand U40737 (N_40737,N_40395,N_40296);
xnor U40738 (N_40738,N_40018,N_40380);
nor U40739 (N_40739,N_40258,N_40443);
xnor U40740 (N_40740,N_40193,N_40489);
and U40741 (N_40741,N_40347,N_40496);
nand U40742 (N_40742,N_40154,N_40212);
and U40743 (N_40743,N_40012,N_40117);
or U40744 (N_40744,N_40168,N_40326);
nor U40745 (N_40745,N_40235,N_40480);
xnor U40746 (N_40746,N_40076,N_40441);
or U40747 (N_40747,N_40190,N_40002);
nor U40748 (N_40748,N_40253,N_40068);
nand U40749 (N_40749,N_40025,N_40379);
nor U40750 (N_40750,N_40001,N_40004);
or U40751 (N_40751,N_40064,N_40186);
or U40752 (N_40752,N_40300,N_40350);
nand U40753 (N_40753,N_40049,N_40358);
nor U40754 (N_40754,N_40127,N_40487);
or U40755 (N_40755,N_40465,N_40449);
and U40756 (N_40756,N_40495,N_40424);
or U40757 (N_40757,N_40094,N_40112);
nand U40758 (N_40758,N_40319,N_40047);
nand U40759 (N_40759,N_40105,N_40407);
and U40760 (N_40760,N_40316,N_40418);
or U40761 (N_40761,N_40036,N_40130);
or U40762 (N_40762,N_40044,N_40373);
or U40763 (N_40763,N_40131,N_40437);
and U40764 (N_40764,N_40221,N_40382);
xnor U40765 (N_40765,N_40129,N_40497);
nor U40766 (N_40766,N_40340,N_40128);
nor U40767 (N_40767,N_40486,N_40469);
nand U40768 (N_40768,N_40175,N_40230);
nand U40769 (N_40769,N_40336,N_40404);
or U40770 (N_40770,N_40185,N_40451);
nand U40771 (N_40771,N_40130,N_40408);
or U40772 (N_40772,N_40468,N_40339);
nor U40773 (N_40773,N_40026,N_40441);
nor U40774 (N_40774,N_40450,N_40235);
nand U40775 (N_40775,N_40365,N_40472);
nand U40776 (N_40776,N_40197,N_40216);
and U40777 (N_40777,N_40489,N_40032);
nand U40778 (N_40778,N_40404,N_40389);
nand U40779 (N_40779,N_40172,N_40099);
nand U40780 (N_40780,N_40220,N_40012);
nor U40781 (N_40781,N_40280,N_40455);
nand U40782 (N_40782,N_40322,N_40054);
and U40783 (N_40783,N_40309,N_40423);
nor U40784 (N_40784,N_40185,N_40285);
and U40785 (N_40785,N_40110,N_40215);
nor U40786 (N_40786,N_40176,N_40051);
xnor U40787 (N_40787,N_40190,N_40487);
nand U40788 (N_40788,N_40256,N_40293);
nand U40789 (N_40789,N_40264,N_40405);
or U40790 (N_40790,N_40280,N_40103);
xor U40791 (N_40791,N_40222,N_40295);
xnor U40792 (N_40792,N_40174,N_40093);
and U40793 (N_40793,N_40175,N_40412);
or U40794 (N_40794,N_40054,N_40318);
xnor U40795 (N_40795,N_40466,N_40186);
xor U40796 (N_40796,N_40219,N_40497);
nor U40797 (N_40797,N_40131,N_40482);
and U40798 (N_40798,N_40311,N_40086);
and U40799 (N_40799,N_40300,N_40159);
xor U40800 (N_40800,N_40066,N_40418);
and U40801 (N_40801,N_40389,N_40003);
or U40802 (N_40802,N_40118,N_40424);
nor U40803 (N_40803,N_40288,N_40180);
nor U40804 (N_40804,N_40023,N_40427);
xor U40805 (N_40805,N_40097,N_40028);
nand U40806 (N_40806,N_40474,N_40112);
nand U40807 (N_40807,N_40384,N_40241);
and U40808 (N_40808,N_40151,N_40318);
nand U40809 (N_40809,N_40146,N_40394);
nor U40810 (N_40810,N_40348,N_40147);
nor U40811 (N_40811,N_40032,N_40344);
xnor U40812 (N_40812,N_40143,N_40153);
or U40813 (N_40813,N_40345,N_40473);
nor U40814 (N_40814,N_40339,N_40304);
xor U40815 (N_40815,N_40188,N_40098);
nand U40816 (N_40816,N_40298,N_40394);
nand U40817 (N_40817,N_40140,N_40340);
or U40818 (N_40818,N_40189,N_40179);
and U40819 (N_40819,N_40483,N_40143);
nand U40820 (N_40820,N_40440,N_40400);
nor U40821 (N_40821,N_40069,N_40410);
xor U40822 (N_40822,N_40327,N_40153);
and U40823 (N_40823,N_40393,N_40356);
xnor U40824 (N_40824,N_40014,N_40420);
and U40825 (N_40825,N_40404,N_40094);
or U40826 (N_40826,N_40481,N_40058);
nand U40827 (N_40827,N_40387,N_40486);
or U40828 (N_40828,N_40055,N_40168);
or U40829 (N_40829,N_40033,N_40454);
and U40830 (N_40830,N_40232,N_40454);
and U40831 (N_40831,N_40176,N_40199);
nand U40832 (N_40832,N_40472,N_40288);
xnor U40833 (N_40833,N_40276,N_40492);
or U40834 (N_40834,N_40474,N_40111);
and U40835 (N_40835,N_40168,N_40020);
and U40836 (N_40836,N_40466,N_40486);
nor U40837 (N_40837,N_40175,N_40300);
nand U40838 (N_40838,N_40352,N_40410);
nor U40839 (N_40839,N_40185,N_40435);
or U40840 (N_40840,N_40383,N_40100);
and U40841 (N_40841,N_40462,N_40252);
nor U40842 (N_40842,N_40394,N_40014);
nand U40843 (N_40843,N_40085,N_40325);
or U40844 (N_40844,N_40204,N_40119);
nand U40845 (N_40845,N_40337,N_40041);
nand U40846 (N_40846,N_40060,N_40217);
xor U40847 (N_40847,N_40003,N_40190);
nand U40848 (N_40848,N_40387,N_40050);
nor U40849 (N_40849,N_40152,N_40047);
and U40850 (N_40850,N_40328,N_40163);
or U40851 (N_40851,N_40479,N_40418);
xnor U40852 (N_40852,N_40349,N_40223);
and U40853 (N_40853,N_40330,N_40474);
or U40854 (N_40854,N_40433,N_40206);
xnor U40855 (N_40855,N_40457,N_40206);
xor U40856 (N_40856,N_40216,N_40380);
or U40857 (N_40857,N_40135,N_40366);
xor U40858 (N_40858,N_40018,N_40460);
nor U40859 (N_40859,N_40286,N_40120);
or U40860 (N_40860,N_40042,N_40222);
nor U40861 (N_40861,N_40338,N_40292);
nor U40862 (N_40862,N_40021,N_40422);
nor U40863 (N_40863,N_40176,N_40134);
nand U40864 (N_40864,N_40423,N_40016);
nand U40865 (N_40865,N_40132,N_40031);
and U40866 (N_40866,N_40430,N_40403);
xnor U40867 (N_40867,N_40063,N_40485);
or U40868 (N_40868,N_40045,N_40481);
xnor U40869 (N_40869,N_40289,N_40291);
nor U40870 (N_40870,N_40020,N_40180);
xor U40871 (N_40871,N_40149,N_40412);
or U40872 (N_40872,N_40051,N_40398);
nor U40873 (N_40873,N_40318,N_40210);
xnor U40874 (N_40874,N_40199,N_40029);
and U40875 (N_40875,N_40419,N_40104);
and U40876 (N_40876,N_40114,N_40425);
and U40877 (N_40877,N_40222,N_40256);
nor U40878 (N_40878,N_40123,N_40186);
nand U40879 (N_40879,N_40264,N_40207);
nor U40880 (N_40880,N_40477,N_40032);
nand U40881 (N_40881,N_40344,N_40380);
and U40882 (N_40882,N_40112,N_40067);
xnor U40883 (N_40883,N_40184,N_40060);
nand U40884 (N_40884,N_40454,N_40316);
xor U40885 (N_40885,N_40404,N_40098);
xnor U40886 (N_40886,N_40465,N_40071);
or U40887 (N_40887,N_40336,N_40147);
nand U40888 (N_40888,N_40449,N_40351);
nand U40889 (N_40889,N_40158,N_40005);
or U40890 (N_40890,N_40366,N_40041);
and U40891 (N_40891,N_40118,N_40230);
nor U40892 (N_40892,N_40051,N_40356);
nand U40893 (N_40893,N_40419,N_40171);
and U40894 (N_40894,N_40410,N_40291);
nand U40895 (N_40895,N_40413,N_40305);
nor U40896 (N_40896,N_40312,N_40319);
xnor U40897 (N_40897,N_40397,N_40447);
and U40898 (N_40898,N_40374,N_40473);
xnor U40899 (N_40899,N_40456,N_40015);
nand U40900 (N_40900,N_40225,N_40404);
xnor U40901 (N_40901,N_40493,N_40339);
nand U40902 (N_40902,N_40278,N_40156);
nor U40903 (N_40903,N_40033,N_40261);
xor U40904 (N_40904,N_40236,N_40492);
or U40905 (N_40905,N_40222,N_40086);
nor U40906 (N_40906,N_40117,N_40133);
and U40907 (N_40907,N_40387,N_40105);
or U40908 (N_40908,N_40355,N_40018);
and U40909 (N_40909,N_40070,N_40150);
nor U40910 (N_40910,N_40491,N_40458);
or U40911 (N_40911,N_40496,N_40197);
xnor U40912 (N_40912,N_40488,N_40222);
and U40913 (N_40913,N_40325,N_40166);
or U40914 (N_40914,N_40140,N_40175);
or U40915 (N_40915,N_40060,N_40007);
nand U40916 (N_40916,N_40205,N_40249);
xnor U40917 (N_40917,N_40254,N_40320);
nor U40918 (N_40918,N_40390,N_40126);
or U40919 (N_40919,N_40298,N_40181);
nand U40920 (N_40920,N_40237,N_40398);
or U40921 (N_40921,N_40271,N_40132);
nor U40922 (N_40922,N_40185,N_40369);
xor U40923 (N_40923,N_40472,N_40221);
and U40924 (N_40924,N_40143,N_40348);
and U40925 (N_40925,N_40445,N_40187);
or U40926 (N_40926,N_40009,N_40477);
nor U40927 (N_40927,N_40021,N_40303);
xor U40928 (N_40928,N_40255,N_40187);
nor U40929 (N_40929,N_40262,N_40123);
nand U40930 (N_40930,N_40183,N_40242);
nand U40931 (N_40931,N_40122,N_40295);
xnor U40932 (N_40932,N_40109,N_40110);
nand U40933 (N_40933,N_40141,N_40399);
and U40934 (N_40934,N_40135,N_40492);
and U40935 (N_40935,N_40218,N_40105);
or U40936 (N_40936,N_40062,N_40166);
xnor U40937 (N_40937,N_40087,N_40498);
nor U40938 (N_40938,N_40304,N_40468);
nand U40939 (N_40939,N_40264,N_40382);
xnor U40940 (N_40940,N_40288,N_40164);
nor U40941 (N_40941,N_40175,N_40399);
nand U40942 (N_40942,N_40092,N_40048);
nor U40943 (N_40943,N_40057,N_40395);
and U40944 (N_40944,N_40489,N_40455);
nand U40945 (N_40945,N_40173,N_40492);
xnor U40946 (N_40946,N_40163,N_40156);
nor U40947 (N_40947,N_40060,N_40113);
nor U40948 (N_40948,N_40011,N_40216);
nor U40949 (N_40949,N_40398,N_40423);
xnor U40950 (N_40950,N_40013,N_40433);
nand U40951 (N_40951,N_40113,N_40025);
nor U40952 (N_40952,N_40453,N_40417);
and U40953 (N_40953,N_40006,N_40310);
nor U40954 (N_40954,N_40246,N_40344);
or U40955 (N_40955,N_40485,N_40141);
nor U40956 (N_40956,N_40057,N_40278);
and U40957 (N_40957,N_40202,N_40072);
xor U40958 (N_40958,N_40151,N_40398);
nor U40959 (N_40959,N_40457,N_40008);
and U40960 (N_40960,N_40019,N_40402);
xnor U40961 (N_40961,N_40432,N_40498);
and U40962 (N_40962,N_40023,N_40029);
or U40963 (N_40963,N_40293,N_40344);
xnor U40964 (N_40964,N_40424,N_40239);
nor U40965 (N_40965,N_40086,N_40450);
nand U40966 (N_40966,N_40142,N_40197);
nand U40967 (N_40967,N_40321,N_40093);
nand U40968 (N_40968,N_40264,N_40093);
nand U40969 (N_40969,N_40190,N_40371);
nor U40970 (N_40970,N_40406,N_40318);
and U40971 (N_40971,N_40426,N_40258);
and U40972 (N_40972,N_40492,N_40084);
or U40973 (N_40973,N_40412,N_40411);
nor U40974 (N_40974,N_40111,N_40193);
or U40975 (N_40975,N_40270,N_40196);
or U40976 (N_40976,N_40303,N_40032);
nor U40977 (N_40977,N_40002,N_40194);
or U40978 (N_40978,N_40470,N_40206);
and U40979 (N_40979,N_40436,N_40121);
nor U40980 (N_40980,N_40373,N_40171);
nand U40981 (N_40981,N_40348,N_40032);
and U40982 (N_40982,N_40258,N_40034);
and U40983 (N_40983,N_40033,N_40490);
xor U40984 (N_40984,N_40058,N_40304);
and U40985 (N_40985,N_40014,N_40211);
xor U40986 (N_40986,N_40334,N_40477);
nor U40987 (N_40987,N_40124,N_40092);
nand U40988 (N_40988,N_40024,N_40360);
nor U40989 (N_40989,N_40070,N_40120);
xor U40990 (N_40990,N_40315,N_40186);
or U40991 (N_40991,N_40485,N_40377);
nor U40992 (N_40992,N_40037,N_40213);
nor U40993 (N_40993,N_40282,N_40297);
and U40994 (N_40994,N_40055,N_40099);
nand U40995 (N_40995,N_40395,N_40456);
nand U40996 (N_40996,N_40329,N_40016);
or U40997 (N_40997,N_40422,N_40265);
nor U40998 (N_40998,N_40106,N_40246);
or U40999 (N_40999,N_40456,N_40063);
nand U41000 (N_41000,N_40663,N_40696);
and U41001 (N_41001,N_40731,N_40613);
xor U41002 (N_41002,N_40713,N_40777);
or U41003 (N_41003,N_40709,N_40590);
nor U41004 (N_41004,N_40843,N_40558);
nand U41005 (N_41005,N_40623,N_40618);
xnor U41006 (N_41006,N_40534,N_40783);
xnor U41007 (N_41007,N_40738,N_40900);
and U41008 (N_41008,N_40625,N_40581);
nand U41009 (N_41009,N_40881,N_40782);
xnor U41010 (N_41010,N_40809,N_40703);
xnor U41011 (N_41011,N_40903,N_40682);
nor U41012 (N_41012,N_40688,N_40943);
and U41013 (N_41013,N_40659,N_40811);
nand U41014 (N_41014,N_40819,N_40914);
nand U41015 (N_41015,N_40949,N_40998);
nor U41016 (N_41016,N_40673,N_40630);
xor U41017 (N_41017,N_40946,N_40816);
nand U41018 (N_41018,N_40970,N_40854);
and U41019 (N_41019,N_40707,N_40667);
xor U41020 (N_41020,N_40990,N_40825);
nor U41021 (N_41021,N_40901,N_40519);
nor U41022 (N_41022,N_40657,N_40884);
xnor U41023 (N_41023,N_40873,N_40741);
and U41024 (N_41024,N_40617,N_40547);
and U41025 (N_41025,N_40789,N_40818);
or U41026 (N_41026,N_40660,N_40747);
nand U41027 (N_41027,N_40714,N_40891);
nor U41028 (N_41028,N_40542,N_40523);
nor U41029 (N_41029,N_40629,N_40728);
nor U41030 (N_41030,N_40948,N_40537);
xnor U41031 (N_41031,N_40940,N_40722);
nand U41032 (N_41032,N_40958,N_40744);
and U41033 (N_41033,N_40762,N_40679);
xnor U41034 (N_41034,N_40608,N_40504);
nor U41035 (N_41035,N_40899,N_40692);
nor U41036 (N_41036,N_40592,N_40665);
or U41037 (N_41037,N_40971,N_40862);
and U41038 (N_41038,N_40840,N_40969);
nor U41039 (N_41039,N_40829,N_40616);
or U41040 (N_41040,N_40520,N_40574);
nand U41041 (N_41041,N_40935,N_40975);
or U41042 (N_41042,N_40906,N_40742);
nor U41043 (N_41043,N_40869,N_40951);
nor U41044 (N_41044,N_40996,N_40539);
xor U41045 (N_41045,N_40973,N_40536);
nand U41046 (N_41046,N_40565,N_40955);
and U41047 (N_41047,N_40761,N_40868);
xor U41048 (N_41048,N_40930,N_40720);
xnor U41049 (N_41049,N_40705,N_40904);
xor U41050 (N_41050,N_40965,N_40598);
and U41051 (N_41051,N_40745,N_40715);
and U41052 (N_41052,N_40963,N_40995);
xor U41053 (N_41053,N_40781,N_40509);
xnor U41054 (N_41054,N_40966,N_40627);
or U41055 (N_41055,N_40878,N_40922);
or U41056 (N_41056,N_40837,N_40985);
and U41057 (N_41057,N_40620,N_40847);
xnor U41058 (N_41058,N_40656,N_40924);
xnor U41059 (N_41059,N_40954,N_40987);
xnor U41060 (N_41060,N_40612,N_40810);
and U41061 (N_41061,N_40826,N_40572);
nand U41062 (N_41062,N_40957,N_40889);
and U41063 (N_41063,N_40516,N_40893);
and U41064 (N_41064,N_40575,N_40902);
nand U41065 (N_41065,N_40897,N_40806);
xor U41066 (N_41066,N_40723,N_40799);
and U41067 (N_41067,N_40875,N_40942);
xnor U41068 (N_41068,N_40931,N_40538);
or U41069 (N_41069,N_40918,N_40756);
or U41070 (N_41070,N_40726,N_40595);
xnor U41071 (N_41071,N_40680,N_40774);
and U41072 (N_41072,N_40813,N_40877);
and U41073 (N_41073,N_40508,N_40736);
xnor U41074 (N_41074,N_40796,N_40882);
or U41075 (N_41075,N_40808,N_40588);
xnor U41076 (N_41076,N_40765,N_40863);
nor U41077 (N_41077,N_40671,N_40716);
nand U41078 (N_41078,N_40820,N_40913);
nand U41079 (N_41079,N_40658,N_40921);
or U41080 (N_41080,N_40593,N_40981);
and U41081 (N_41081,N_40936,N_40859);
or U41082 (N_41082,N_40685,N_40621);
or U41083 (N_41083,N_40732,N_40670);
xor U41084 (N_41084,N_40886,N_40832);
and U41085 (N_41085,N_40580,N_40769);
nor U41086 (N_41086,N_40999,N_40645);
nand U41087 (N_41087,N_40833,N_40545);
nand U41088 (N_41088,N_40532,N_40885);
nor U41089 (N_41089,N_40635,N_40586);
nor U41090 (N_41090,N_40944,N_40896);
or U41091 (N_41091,N_40546,N_40561);
or U41092 (N_41092,N_40780,N_40968);
or U41093 (N_41093,N_40980,N_40651);
or U41094 (N_41094,N_40648,N_40779);
nor U41095 (N_41095,N_40945,N_40652);
or U41096 (N_41096,N_40555,N_40915);
nor U41097 (N_41097,N_40950,N_40690);
xnor U41098 (N_41098,N_40522,N_40937);
and U41099 (N_41099,N_40784,N_40661);
nand U41100 (N_41100,N_40846,N_40636);
nor U41101 (N_41101,N_40753,N_40543);
or U41102 (N_41102,N_40755,N_40735);
nor U41103 (N_41103,N_40668,N_40835);
xnor U41104 (N_41104,N_40876,N_40763);
nor U41105 (N_41105,N_40737,N_40601);
or U41106 (N_41106,N_40619,N_40802);
and U41107 (N_41107,N_40631,N_40710);
nand U41108 (N_41108,N_40834,N_40997);
xor U41109 (N_41109,N_40634,N_40920);
xnor U41110 (N_41110,N_40719,N_40739);
xor U41111 (N_41111,N_40778,N_40655);
xor U41112 (N_41112,N_40677,N_40867);
and U41113 (N_41113,N_40866,N_40684);
nand U41114 (N_41114,N_40919,N_40979);
xor U41115 (N_41115,N_40573,N_40552);
xnor U41116 (N_41116,N_40959,N_40910);
nor U41117 (N_41117,N_40697,N_40579);
nor U41118 (N_41118,N_40515,N_40939);
and U41119 (N_41119,N_40853,N_40842);
xnor U41120 (N_41120,N_40960,N_40767);
nor U41121 (N_41121,N_40609,N_40535);
nor U41122 (N_41122,N_40928,N_40503);
nand U41123 (N_41123,N_40938,N_40956);
nand U41124 (N_41124,N_40585,N_40838);
xnor U41125 (N_41125,N_40757,N_40754);
nand U41126 (N_41126,N_40982,N_40553);
xnor U41127 (N_41127,N_40871,N_40698);
or U41128 (N_41128,N_40798,N_40894);
or U41129 (N_41129,N_40992,N_40725);
nor U41130 (N_41130,N_40740,N_40927);
nor U41131 (N_41131,N_40977,N_40815);
nand U41132 (N_41132,N_40734,N_40908);
nor U41133 (N_41133,N_40702,N_40510);
or U41134 (N_41134,N_40639,N_40786);
and U41135 (N_41135,N_40770,N_40706);
nor U41136 (N_41136,N_40701,N_40972);
nand U41137 (N_41137,N_40895,N_40967);
and U41138 (N_41138,N_40856,N_40604);
nand U41139 (N_41139,N_40898,N_40917);
nor U41140 (N_41140,N_40772,N_40501);
xnor U41141 (N_41141,N_40564,N_40531);
nand U41142 (N_41142,N_40525,N_40794);
nor U41143 (N_41143,N_40708,N_40812);
nand U41144 (N_41144,N_40600,N_40821);
xor U41145 (N_41145,N_40978,N_40879);
nand U41146 (N_41146,N_40724,N_40548);
or U41147 (N_41147,N_40888,N_40584);
xor U41148 (N_41148,N_40610,N_40599);
and U41149 (N_41149,N_40807,N_40817);
xnor U41150 (N_41150,N_40865,N_40790);
and U41151 (N_41151,N_40567,N_40589);
xor U41152 (N_41152,N_40549,N_40550);
xnor U41153 (N_41153,N_40828,N_40594);
xnor U41154 (N_41154,N_40596,N_40932);
nand U41155 (N_41155,N_40526,N_40562);
and U41156 (N_41156,N_40524,N_40729);
nand U41157 (N_41157,N_40974,N_40801);
xor U41158 (N_41158,N_40712,N_40760);
xor U41159 (N_41159,N_40788,N_40864);
or U41160 (N_41160,N_40986,N_40803);
or U41161 (N_41161,N_40576,N_40674);
nand U41162 (N_41162,N_40764,N_40749);
xor U41163 (N_41163,N_40676,N_40583);
xor U41164 (N_41164,N_40672,N_40560);
xor U41165 (N_41165,N_40923,N_40822);
and U41166 (N_41166,N_40533,N_40528);
and U41167 (N_41167,N_40664,N_40711);
xor U41168 (N_41168,N_40892,N_40855);
or U41169 (N_41169,N_40751,N_40653);
nor U41170 (N_41170,N_40839,N_40683);
xnor U41171 (N_41171,N_40797,N_40953);
nand U41172 (N_41172,N_40880,N_40785);
nand U41173 (N_41173,N_40861,N_40527);
and U41174 (N_41174,N_40993,N_40603);
nand U41175 (N_41175,N_40795,N_40976);
or U41176 (N_41176,N_40518,N_40607);
xnor U41177 (N_41177,N_40872,N_40556);
nor U41178 (N_41178,N_40551,N_40626);
nand U41179 (N_41179,N_40768,N_40718);
nor U41180 (N_41180,N_40606,N_40704);
nor U41181 (N_41181,N_40500,N_40849);
nor U41182 (N_41182,N_40644,N_40746);
xnor U41183 (N_41183,N_40577,N_40650);
xnor U41184 (N_41184,N_40571,N_40773);
xnor U41185 (N_41185,N_40907,N_40568);
or U41186 (N_41186,N_40654,N_40637);
nor U41187 (N_41187,N_40814,N_40721);
nor U41188 (N_41188,N_40752,N_40994);
xnor U41189 (N_41189,N_40952,N_40544);
nand U41190 (N_41190,N_40929,N_40597);
nor U41191 (N_41191,N_40681,N_40771);
xnor U41192 (N_41192,N_40694,N_40850);
xor U41193 (N_41193,N_40727,N_40529);
nor U41194 (N_41194,N_40874,N_40750);
and U41195 (N_41195,N_40824,N_40554);
or U41196 (N_41196,N_40941,N_40649);
xor U41197 (N_41197,N_40633,N_40800);
xnor U41198 (N_41198,N_40883,N_40860);
or U41199 (N_41199,N_40557,N_40909);
and U41200 (N_41200,N_40689,N_40514);
xnor U41201 (N_41201,N_40793,N_40691);
nor U41202 (N_41202,N_40759,N_40787);
nor U41203 (N_41203,N_40890,N_40628);
or U41204 (N_41204,N_40743,N_40934);
or U41205 (N_41205,N_40662,N_40506);
and U41206 (N_41206,N_40717,N_40611);
or U41207 (N_41207,N_40541,N_40730);
and U41208 (N_41208,N_40669,N_40587);
nor U41209 (N_41209,N_40858,N_40733);
nand U41210 (N_41210,N_40766,N_40693);
and U41211 (N_41211,N_40686,N_40517);
xor U41212 (N_41212,N_40845,N_40513);
and U41213 (N_41213,N_40988,N_40640);
or U41214 (N_41214,N_40638,N_40823);
nand U41215 (N_41215,N_40905,N_40605);
nand U41216 (N_41216,N_40887,N_40502);
nor U41217 (N_41217,N_40852,N_40622);
nand U41218 (N_41218,N_40505,N_40624);
nor U41219 (N_41219,N_40962,N_40848);
or U41220 (N_41220,N_40804,N_40827);
and U41221 (N_41221,N_40559,N_40646);
nor U41222 (N_41222,N_40916,N_40570);
and U41223 (N_41223,N_40540,N_40925);
xor U41224 (N_41224,N_40511,N_40602);
nor U41225 (N_41225,N_40700,N_40911);
nand U41226 (N_41226,N_40566,N_40912);
or U41227 (N_41227,N_40964,N_40530);
or U41228 (N_41228,N_40591,N_40699);
nand U41229 (N_41229,N_40851,N_40512);
and U41230 (N_41230,N_40641,N_40748);
xnor U41231 (N_41231,N_40675,N_40830);
and U41232 (N_41232,N_40961,N_40831);
nor U41233 (N_41233,N_40857,N_40632);
nor U41234 (N_41234,N_40678,N_40507);
and U41235 (N_41235,N_40643,N_40578);
xor U41236 (N_41236,N_40687,N_40947);
nand U41237 (N_41237,N_40989,N_40933);
or U41238 (N_41238,N_40792,N_40836);
and U41239 (N_41239,N_40642,N_40614);
or U41240 (N_41240,N_40805,N_40615);
or U41241 (N_41241,N_40776,N_40984);
nand U41242 (N_41242,N_40775,N_40841);
xor U41243 (N_41243,N_40647,N_40844);
xor U41244 (N_41244,N_40582,N_40870);
xnor U41245 (N_41245,N_40569,N_40926);
and U41246 (N_41246,N_40991,N_40758);
xnor U41247 (N_41247,N_40563,N_40983);
xnor U41248 (N_41248,N_40666,N_40791);
or U41249 (N_41249,N_40521,N_40695);
nor U41250 (N_41250,N_40609,N_40951);
xnor U41251 (N_41251,N_40872,N_40864);
and U41252 (N_41252,N_40583,N_40945);
nor U41253 (N_41253,N_40985,N_40542);
or U41254 (N_41254,N_40510,N_40901);
nand U41255 (N_41255,N_40828,N_40735);
nor U41256 (N_41256,N_40656,N_40822);
xnor U41257 (N_41257,N_40817,N_40996);
nand U41258 (N_41258,N_40892,N_40560);
and U41259 (N_41259,N_40887,N_40741);
and U41260 (N_41260,N_40973,N_40951);
or U41261 (N_41261,N_40732,N_40709);
nand U41262 (N_41262,N_40642,N_40620);
and U41263 (N_41263,N_40898,N_40873);
nand U41264 (N_41264,N_40882,N_40902);
and U41265 (N_41265,N_40700,N_40995);
xnor U41266 (N_41266,N_40605,N_40778);
nor U41267 (N_41267,N_40710,N_40585);
nor U41268 (N_41268,N_40990,N_40888);
nand U41269 (N_41269,N_40902,N_40530);
and U41270 (N_41270,N_40509,N_40693);
nor U41271 (N_41271,N_40510,N_40500);
or U41272 (N_41272,N_40923,N_40551);
nor U41273 (N_41273,N_40551,N_40521);
or U41274 (N_41274,N_40515,N_40820);
and U41275 (N_41275,N_40635,N_40660);
and U41276 (N_41276,N_40823,N_40841);
or U41277 (N_41277,N_40566,N_40857);
and U41278 (N_41278,N_40852,N_40975);
nand U41279 (N_41279,N_40598,N_40670);
nor U41280 (N_41280,N_40713,N_40696);
and U41281 (N_41281,N_40506,N_40577);
nor U41282 (N_41282,N_40594,N_40617);
nand U41283 (N_41283,N_40552,N_40590);
xnor U41284 (N_41284,N_40611,N_40724);
and U41285 (N_41285,N_40960,N_40785);
or U41286 (N_41286,N_40746,N_40673);
nand U41287 (N_41287,N_40755,N_40531);
or U41288 (N_41288,N_40529,N_40856);
and U41289 (N_41289,N_40902,N_40984);
nand U41290 (N_41290,N_40992,N_40504);
nand U41291 (N_41291,N_40716,N_40786);
xor U41292 (N_41292,N_40867,N_40693);
or U41293 (N_41293,N_40862,N_40827);
xor U41294 (N_41294,N_40590,N_40934);
or U41295 (N_41295,N_40538,N_40810);
or U41296 (N_41296,N_40900,N_40913);
xor U41297 (N_41297,N_40658,N_40759);
and U41298 (N_41298,N_40759,N_40686);
and U41299 (N_41299,N_40765,N_40716);
xnor U41300 (N_41300,N_40964,N_40989);
or U41301 (N_41301,N_40529,N_40847);
nand U41302 (N_41302,N_40516,N_40721);
and U41303 (N_41303,N_40829,N_40972);
xor U41304 (N_41304,N_40692,N_40941);
xor U41305 (N_41305,N_40946,N_40549);
and U41306 (N_41306,N_40907,N_40623);
xnor U41307 (N_41307,N_40687,N_40622);
or U41308 (N_41308,N_40508,N_40640);
xnor U41309 (N_41309,N_40782,N_40554);
nor U41310 (N_41310,N_40602,N_40896);
nor U41311 (N_41311,N_40606,N_40675);
xnor U41312 (N_41312,N_40609,N_40512);
nor U41313 (N_41313,N_40768,N_40807);
and U41314 (N_41314,N_40689,N_40972);
xnor U41315 (N_41315,N_40798,N_40595);
nand U41316 (N_41316,N_40649,N_40710);
xnor U41317 (N_41317,N_40836,N_40625);
or U41318 (N_41318,N_40827,N_40669);
xor U41319 (N_41319,N_40500,N_40876);
nor U41320 (N_41320,N_40602,N_40743);
nand U41321 (N_41321,N_40505,N_40693);
nor U41322 (N_41322,N_40813,N_40705);
and U41323 (N_41323,N_40690,N_40976);
nor U41324 (N_41324,N_40546,N_40669);
nand U41325 (N_41325,N_40668,N_40974);
xor U41326 (N_41326,N_40815,N_40707);
or U41327 (N_41327,N_40927,N_40633);
or U41328 (N_41328,N_40922,N_40674);
and U41329 (N_41329,N_40572,N_40671);
or U41330 (N_41330,N_40688,N_40597);
or U41331 (N_41331,N_40878,N_40526);
and U41332 (N_41332,N_40598,N_40665);
or U41333 (N_41333,N_40851,N_40924);
and U41334 (N_41334,N_40525,N_40580);
or U41335 (N_41335,N_40588,N_40716);
xor U41336 (N_41336,N_40856,N_40981);
nand U41337 (N_41337,N_40888,N_40794);
and U41338 (N_41338,N_40569,N_40933);
xnor U41339 (N_41339,N_40883,N_40562);
or U41340 (N_41340,N_40601,N_40693);
or U41341 (N_41341,N_40684,N_40725);
xor U41342 (N_41342,N_40995,N_40744);
nor U41343 (N_41343,N_40840,N_40853);
and U41344 (N_41344,N_40529,N_40546);
nor U41345 (N_41345,N_40831,N_40980);
nand U41346 (N_41346,N_40913,N_40658);
xnor U41347 (N_41347,N_40520,N_40898);
and U41348 (N_41348,N_40976,N_40925);
nor U41349 (N_41349,N_40614,N_40581);
xor U41350 (N_41350,N_40994,N_40899);
or U41351 (N_41351,N_40553,N_40543);
or U41352 (N_41352,N_40973,N_40932);
xor U41353 (N_41353,N_40879,N_40573);
and U41354 (N_41354,N_40536,N_40857);
nand U41355 (N_41355,N_40928,N_40835);
nand U41356 (N_41356,N_40542,N_40662);
nor U41357 (N_41357,N_40830,N_40768);
xnor U41358 (N_41358,N_40641,N_40598);
nor U41359 (N_41359,N_40551,N_40781);
nor U41360 (N_41360,N_40547,N_40981);
xnor U41361 (N_41361,N_40588,N_40681);
nor U41362 (N_41362,N_40872,N_40926);
nand U41363 (N_41363,N_40521,N_40601);
or U41364 (N_41364,N_40529,N_40621);
and U41365 (N_41365,N_40895,N_40698);
nand U41366 (N_41366,N_40994,N_40551);
nor U41367 (N_41367,N_40636,N_40825);
xor U41368 (N_41368,N_40578,N_40949);
xor U41369 (N_41369,N_40902,N_40689);
and U41370 (N_41370,N_40998,N_40627);
xor U41371 (N_41371,N_40776,N_40780);
or U41372 (N_41372,N_40707,N_40734);
and U41373 (N_41373,N_40691,N_40765);
or U41374 (N_41374,N_40783,N_40883);
nand U41375 (N_41375,N_40759,N_40610);
nor U41376 (N_41376,N_40763,N_40922);
nor U41377 (N_41377,N_40753,N_40768);
or U41378 (N_41378,N_40959,N_40690);
nand U41379 (N_41379,N_40916,N_40850);
nand U41380 (N_41380,N_40513,N_40777);
nand U41381 (N_41381,N_40677,N_40640);
or U41382 (N_41382,N_40940,N_40921);
and U41383 (N_41383,N_40876,N_40694);
xnor U41384 (N_41384,N_40930,N_40971);
nand U41385 (N_41385,N_40532,N_40500);
xnor U41386 (N_41386,N_40996,N_40980);
and U41387 (N_41387,N_40678,N_40555);
and U41388 (N_41388,N_40747,N_40885);
nand U41389 (N_41389,N_40978,N_40621);
or U41390 (N_41390,N_40989,N_40619);
and U41391 (N_41391,N_40804,N_40608);
or U41392 (N_41392,N_40893,N_40530);
nor U41393 (N_41393,N_40980,N_40909);
or U41394 (N_41394,N_40912,N_40780);
and U41395 (N_41395,N_40669,N_40892);
or U41396 (N_41396,N_40664,N_40749);
nand U41397 (N_41397,N_40540,N_40612);
and U41398 (N_41398,N_40806,N_40559);
nand U41399 (N_41399,N_40651,N_40658);
and U41400 (N_41400,N_40689,N_40988);
nor U41401 (N_41401,N_40787,N_40707);
or U41402 (N_41402,N_40634,N_40723);
nor U41403 (N_41403,N_40744,N_40554);
or U41404 (N_41404,N_40629,N_40731);
or U41405 (N_41405,N_40968,N_40813);
and U41406 (N_41406,N_40732,N_40876);
xnor U41407 (N_41407,N_40915,N_40765);
nand U41408 (N_41408,N_40884,N_40621);
nand U41409 (N_41409,N_40918,N_40801);
nor U41410 (N_41410,N_40507,N_40550);
nor U41411 (N_41411,N_40539,N_40517);
and U41412 (N_41412,N_40577,N_40565);
or U41413 (N_41413,N_40721,N_40936);
and U41414 (N_41414,N_40898,N_40566);
nor U41415 (N_41415,N_40875,N_40888);
nor U41416 (N_41416,N_40627,N_40883);
or U41417 (N_41417,N_40576,N_40607);
and U41418 (N_41418,N_40994,N_40851);
nor U41419 (N_41419,N_40917,N_40850);
and U41420 (N_41420,N_40583,N_40550);
and U41421 (N_41421,N_40998,N_40885);
xor U41422 (N_41422,N_40758,N_40870);
nand U41423 (N_41423,N_40922,N_40952);
or U41424 (N_41424,N_40635,N_40838);
xor U41425 (N_41425,N_40646,N_40678);
or U41426 (N_41426,N_40882,N_40769);
xnor U41427 (N_41427,N_40844,N_40814);
nand U41428 (N_41428,N_40624,N_40854);
nor U41429 (N_41429,N_40581,N_40867);
and U41430 (N_41430,N_40700,N_40752);
nand U41431 (N_41431,N_40927,N_40971);
nor U41432 (N_41432,N_40674,N_40916);
nand U41433 (N_41433,N_40995,N_40566);
or U41434 (N_41434,N_40750,N_40676);
and U41435 (N_41435,N_40778,N_40685);
or U41436 (N_41436,N_40984,N_40699);
xor U41437 (N_41437,N_40739,N_40787);
or U41438 (N_41438,N_40827,N_40585);
nor U41439 (N_41439,N_40990,N_40697);
nand U41440 (N_41440,N_40542,N_40711);
nand U41441 (N_41441,N_40650,N_40718);
nor U41442 (N_41442,N_40685,N_40937);
nor U41443 (N_41443,N_40637,N_40869);
nor U41444 (N_41444,N_40637,N_40605);
and U41445 (N_41445,N_40924,N_40520);
and U41446 (N_41446,N_40621,N_40829);
nor U41447 (N_41447,N_40914,N_40956);
nor U41448 (N_41448,N_40871,N_40510);
or U41449 (N_41449,N_40748,N_40735);
and U41450 (N_41450,N_40821,N_40702);
or U41451 (N_41451,N_40794,N_40801);
nor U41452 (N_41452,N_40593,N_40752);
nand U41453 (N_41453,N_40905,N_40869);
xor U41454 (N_41454,N_40524,N_40802);
or U41455 (N_41455,N_40935,N_40637);
nor U41456 (N_41456,N_40732,N_40696);
nand U41457 (N_41457,N_40903,N_40724);
xnor U41458 (N_41458,N_40925,N_40572);
and U41459 (N_41459,N_40856,N_40603);
xor U41460 (N_41460,N_40653,N_40603);
or U41461 (N_41461,N_40677,N_40795);
nor U41462 (N_41462,N_40640,N_40933);
nor U41463 (N_41463,N_40589,N_40707);
nor U41464 (N_41464,N_40657,N_40507);
or U41465 (N_41465,N_40866,N_40556);
and U41466 (N_41466,N_40859,N_40856);
xnor U41467 (N_41467,N_40946,N_40602);
xnor U41468 (N_41468,N_40723,N_40604);
nor U41469 (N_41469,N_40900,N_40887);
xnor U41470 (N_41470,N_40991,N_40573);
xor U41471 (N_41471,N_40854,N_40882);
xnor U41472 (N_41472,N_40698,N_40604);
nand U41473 (N_41473,N_40524,N_40940);
nand U41474 (N_41474,N_40927,N_40701);
nor U41475 (N_41475,N_40699,N_40917);
or U41476 (N_41476,N_40820,N_40765);
nor U41477 (N_41477,N_40964,N_40544);
or U41478 (N_41478,N_40822,N_40574);
nor U41479 (N_41479,N_40915,N_40582);
and U41480 (N_41480,N_40755,N_40747);
xnor U41481 (N_41481,N_40713,N_40879);
nor U41482 (N_41482,N_40931,N_40972);
nor U41483 (N_41483,N_40963,N_40978);
nor U41484 (N_41484,N_40594,N_40563);
xnor U41485 (N_41485,N_40792,N_40634);
nor U41486 (N_41486,N_40679,N_40809);
nand U41487 (N_41487,N_40894,N_40697);
xnor U41488 (N_41488,N_40556,N_40945);
nand U41489 (N_41489,N_40796,N_40566);
or U41490 (N_41490,N_40606,N_40919);
and U41491 (N_41491,N_40618,N_40792);
or U41492 (N_41492,N_40865,N_40659);
xnor U41493 (N_41493,N_40792,N_40947);
and U41494 (N_41494,N_40774,N_40809);
xnor U41495 (N_41495,N_40895,N_40556);
xnor U41496 (N_41496,N_40667,N_40501);
and U41497 (N_41497,N_40776,N_40870);
nor U41498 (N_41498,N_40910,N_40832);
or U41499 (N_41499,N_40912,N_40741);
or U41500 (N_41500,N_41126,N_41474);
nand U41501 (N_41501,N_41499,N_41356);
nand U41502 (N_41502,N_41434,N_41419);
nor U41503 (N_41503,N_41128,N_41002);
xnor U41504 (N_41504,N_41498,N_41164);
nand U41505 (N_41505,N_41078,N_41281);
and U41506 (N_41506,N_41459,N_41248);
nor U41507 (N_41507,N_41127,N_41407);
and U41508 (N_41508,N_41008,N_41272);
and U41509 (N_41509,N_41184,N_41314);
nor U41510 (N_41510,N_41436,N_41261);
and U41511 (N_41511,N_41321,N_41453);
xnor U41512 (N_41512,N_41188,N_41312);
or U41513 (N_41513,N_41339,N_41165);
and U41514 (N_41514,N_41101,N_41420);
nor U41515 (N_41515,N_41107,N_41087);
nor U41516 (N_41516,N_41462,N_41088);
or U41517 (N_41517,N_41149,N_41297);
or U41518 (N_41518,N_41387,N_41362);
nor U41519 (N_41519,N_41176,N_41284);
nor U41520 (N_41520,N_41195,N_41080);
and U41521 (N_41521,N_41031,N_41024);
or U41522 (N_41522,N_41059,N_41342);
nand U41523 (N_41523,N_41202,N_41097);
and U41524 (N_41524,N_41317,N_41051);
or U41525 (N_41525,N_41390,N_41114);
nand U41526 (N_41526,N_41057,N_41204);
nand U41527 (N_41527,N_41346,N_41327);
xnor U41528 (N_41528,N_41058,N_41095);
and U41529 (N_41529,N_41098,N_41357);
or U41530 (N_41530,N_41181,N_41467);
and U41531 (N_41531,N_41105,N_41163);
or U41532 (N_41532,N_41466,N_41247);
xnor U41533 (N_41533,N_41300,N_41289);
nand U41534 (N_41534,N_41444,N_41416);
or U41535 (N_41535,N_41151,N_41066);
nor U41536 (N_41536,N_41489,N_41380);
xor U41537 (N_41537,N_41180,N_41410);
nor U41538 (N_41538,N_41000,N_41295);
and U41539 (N_41539,N_41381,N_41372);
and U41540 (N_41540,N_41255,N_41085);
nor U41541 (N_41541,N_41082,N_41166);
xnor U41542 (N_41542,N_41113,N_41325);
xnor U41543 (N_41543,N_41009,N_41413);
xor U41544 (N_41544,N_41409,N_41012);
and U41545 (N_41545,N_41182,N_41316);
xor U41546 (N_41546,N_41318,N_41207);
xor U41547 (N_41547,N_41071,N_41227);
or U41548 (N_41548,N_41435,N_41240);
xnor U41549 (N_41549,N_41292,N_41286);
and U41550 (N_41550,N_41469,N_41179);
or U41551 (N_41551,N_41236,N_41385);
xor U41552 (N_41552,N_41359,N_41368);
xor U41553 (N_41553,N_41015,N_41138);
nand U41554 (N_41554,N_41347,N_41104);
xnor U41555 (N_41555,N_41460,N_41230);
or U41556 (N_41556,N_41322,N_41193);
and U41557 (N_41557,N_41427,N_41476);
nor U41558 (N_41558,N_41003,N_41019);
nand U41559 (N_41559,N_41121,N_41177);
nor U41560 (N_41560,N_41254,N_41415);
nand U41561 (N_41561,N_41364,N_41054);
and U41562 (N_41562,N_41200,N_41111);
or U41563 (N_41563,N_41482,N_41344);
nand U41564 (N_41564,N_41172,N_41360);
and U41565 (N_41565,N_41146,N_41171);
xor U41566 (N_41566,N_41418,N_41053);
nand U41567 (N_41567,N_41405,N_41139);
xnor U41568 (N_41568,N_41142,N_41417);
or U41569 (N_41569,N_41096,N_41298);
xor U41570 (N_41570,N_41304,N_41369);
nor U41571 (N_41571,N_41376,N_41170);
or U41572 (N_41572,N_41447,N_41355);
and U41573 (N_41573,N_41190,N_41153);
or U41574 (N_41574,N_41253,N_41186);
and U41575 (N_41575,N_41335,N_41131);
and U41576 (N_41576,N_41354,N_41358);
nor U41577 (N_41577,N_41154,N_41307);
and U41578 (N_41578,N_41198,N_41404);
or U41579 (N_41579,N_41264,N_41068);
and U41580 (N_41580,N_41205,N_41201);
nor U41581 (N_41581,N_41061,N_41238);
xnor U41582 (N_41582,N_41123,N_41218);
and U41583 (N_41583,N_41442,N_41388);
or U41584 (N_41584,N_41135,N_41320);
nor U41585 (N_41585,N_41167,N_41137);
nand U41586 (N_41586,N_41394,N_41004);
and U41587 (N_41587,N_41348,N_41456);
or U41588 (N_41588,N_41283,N_41382);
or U41589 (N_41589,N_41268,N_41219);
xnor U41590 (N_41590,N_41326,N_41036);
nor U41591 (N_41591,N_41150,N_41299);
and U41592 (N_41592,N_41400,N_41412);
xnor U41593 (N_41593,N_41408,N_41373);
xor U41594 (N_41594,N_41161,N_41371);
or U41595 (N_41595,N_41393,N_41311);
and U41596 (N_41596,N_41148,N_41293);
nand U41597 (N_41597,N_41367,N_41158);
and U41598 (N_41598,N_41069,N_41398);
or U41599 (N_41599,N_41162,N_41155);
xor U41600 (N_41600,N_41374,N_41099);
or U41601 (N_41601,N_41199,N_41210);
nor U41602 (N_41602,N_41232,N_41370);
or U41603 (N_41603,N_41256,N_41022);
and U41604 (N_41604,N_41032,N_41076);
or U41605 (N_41605,N_41430,N_41052);
nor U41606 (N_41606,N_41140,N_41470);
nor U41607 (N_41607,N_41334,N_41132);
nor U41608 (N_41608,N_41115,N_41214);
nor U41609 (N_41609,N_41239,N_41090);
nor U41610 (N_41610,N_41483,N_41129);
nor U41611 (N_41611,N_41110,N_41465);
or U41612 (N_41612,N_41014,N_41443);
and U41613 (N_41613,N_41067,N_41455);
nor U41614 (N_41614,N_41157,N_41102);
nor U41615 (N_41615,N_41433,N_41475);
and U41616 (N_41616,N_41363,N_41220);
or U41617 (N_41617,N_41309,N_41136);
nor U41618 (N_41618,N_41235,N_41147);
or U41619 (N_41619,N_41037,N_41496);
and U41620 (N_41620,N_41143,N_41077);
nand U41621 (N_41621,N_41118,N_41464);
nor U41622 (N_41622,N_41124,N_41481);
nor U41623 (N_41623,N_41056,N_41340);
nor U41624 (N_41624,N_41454,N_41492);
xnor U41625 (N_41625,N_41478,N_41332);
xor U41626 (N_41626,N_41221,N_41485);
and U41627 (N_41627,N_41391,N_41323);
nor U41628 (N_41628,N_41040,N_41079);
nand U41629 (N_41629,N_41401,N_41366);
nor U41630 (N_41630,N_41493,N_41187);
and U41631 (N_41631,N_41074,N_41395);
nor U41632 (N_41632,N_41487,N_41065);
xnor U41633 (N_41633,N_41345,N_41389);
and U41634 (N_41634,N_41275,N_41144);
and U41635 (N_41635,N_41249,N_41237);
xor U41636 (N_41636,N_41439,N_41451);
and U41637 (N_41637,N_41486,N_41431);
or U41638 (N_41638,N_41440,N_41156);
nand U41639 (N_41639,N_41263,N_41026);
nor U41640 (N_41640,N_41423,N_41437);
nand U41641 (N_41641,N_41016,N_41203);
xnor U41642 (N_41642,N_41134,N_41365);
nand U41643 (N_41643,N_41461,N_41178);
or U41644 (N_41644,N_41062,N_41086);
nor U41645 (N_41645,N_41288,N_41120);
xnor U41646 (N_41646,N_41396,N_41445);
nor U41647 (N_41647,N_41045,N_41411);
or U41648 (N_41648,N_41215,N_41006);
nand U41649 (N_41649,N_41336,N_41035);
and U41650 (N_41650,N_41094,N_41290);
or U41651 (N_41651,N_41426,N_41243);
nor U41652 (N_41652,N_41241,N_41029);
nand U41653 (N_41653,N_41007,N_41497);
nand U41654 (N_41654,N_41479,N_41250);
nor U41655 (N_41655,N_41046,N_41038);
xor U41656 (N_41656,N_41276,N_41055);
nand U41657 (N_41657,N_41183,N_41048);
and U41658 (N_41658,N_41018,N_41225);
xnor U41659 (N_41659,N_41027,N_41194);
xnor U41660 (N_41660,N_41377,N_41216);
or U41661 (N_41661,N_41108,N_41343);
nand U41662 (N_41662,N_41224,N_41125);
nor U41663 (N_41663,N_41429,N_41477);
xor U41664 (N_41664,N_41173,N_41285);
nor U41665 (N_41665,N_41021,N_41428);
or U41666 (N_41666,N_41025,N_41331);
nor U41667 (N_41667,N_41130,N_41452);
and U41668 (N_41668,N_41338,N_41260);
xnor U41669 (N_41669,N_41034,N_41033);
nand U41670 (N_41670,N_41185,N_41231);
nor U41671 (N_41671,N_41266,N_41217);
or U41672 (N_41672,N_41257,N_41072);
xnor U41673 (N_41673,N_41228,N_41206);
nor U41674 (N_41674,N_41100,N_41277);
and U41675 (N_41675,N_41064,N_41208);
or U41676 (N_41676,N_41406,N_41226);
xnor U41677 (N_41677,N_41092,N_41005);
nand U41678 (N_41678,N_41490,N_41116);
nand U41679 (N_41679,N_41267,N_41378);
or U41680 (N_41680,N_41273,N_41028);
xnor U41681 (N_41681,N_41287,N_41313);
nand U41682 (N_41682,N_41013,N_41352);
nor U41683 (N_41683,N_41303,N_41073);
xnor U41684 (N_41684,N_41089,N_41446);
xor U41685 (N_41685,N_41211,N_41106);
xor U41686 (N_41686,N_41457,N_41122);
nand U41687 (N_41687,N_41229,N_41084);
or U41688 (N_41688,N_41246,N_41463);
or U41689 (N_41689,N_41341,N_41432);
xor U41690 (N_41690,N_41112,N_41421);
and U41691 (N_41691,N_41424,N_41392);
nor U41692 (N_41692,N_41049,N_41450);
and U41693 (N_41693,N_41197,N_41222);
or U41694 (N_41694,N_41480,N_41196);
or U41695 (N_41695,N_41133,N_41001);
and U41696 (N_41696,N_41044,N_41258);
nand U41697 (N_41697,N_41383,N_41192);
or U41698 (N_41698,N_41386,N_41361);
nor U41699 (N_41699,N_41422,N_41353);
nand U41700 (N_41700,N_41093,N_41117);
and U41701 (N_41701,N_41103,N_41043);
and U41702 (N_41702,N_41109,N_41175);
and U41703 (N_41703,N_41050,N_41168);
and U41704 (N_41704,N_41213,N_41242);
and U41705 (N_41705,N_41269,N_41119);
xor U41706 (N_41706,N_41351,N_41244);
or U41707 (N_41707,N_41330,N_41402);
xor U41708 (N_41708,N_41020,N_41223);
nand U41709 (N_41709,N_41145,N_41251);
and U41710 (N_41710,N_41152,N_41472);
or U41711 (N_41711,N_41491,N_41141);
xor U41712 (N_41712,N_41425,N_41234);
and U41713 (N_41713,N_41337,N_41047);
and U41714 (N_41714,N_41379,N_41209);
xor U41715 (N_41715,N_41301,N_41495);
or U41716 (N_41716,N_41274,N_41449);
and U41717 (N_41717,N_41245,N_41011);
nor U41718 (N_41718,N_41329,N_41319);
xor U41719 (N_41719,N_41262,N_41296);
nand U41720 (N_41720,N_41174,N_41441);
xor U41721 (N_41721,N_41397,N_41042);
and U41722 (N_41722,N_41471,N_41160);
nand U41723 (N_41723,N_41399,N_41280);
nand U41724 (N_41724,N_41333,N_41484);
nand U41725 (N_41725,N_41310,N_41233);
xnor U41726 (N_41726,N_41010,N_41030);
xor U41727 (N_41727,N_41291,N_41328);
nor U41728 (N_41728,N_41375,N_41083);
xnor U41729 (N_41729,N_41023,N_41403);
nor U41730 (N_41730,N_41350,N_41282);
and U41731 (N_41731,N_41270,N_41189);
or U41732 (N_41732,N_41265,N_41494);
xor U41733 (N_41733,N_41091,N_41448);
xor U41734 (N_41734,N_41212,N_41039);
or U41735 (N_41735,N_41414,N_41308);
nand U41736 (N_41736,N_41324,N_41438);
nand U41737 (N_41737,N_41271,N_41473);
xor U41738 (N_41738,N_41315,N_41041);
xnor U41739 (N_41739,N_41169,N_41060);
nand U41740 (N_41740,N_41458,N_41488);
nor U41741 (N_41741,N_41259,N_41302);
xnor U41742 (N_41742,N_41017,N_41063);
xnor U41743 (N_41743,N_41349,N_41384);
and U41744 (N_41744,N_41252,N_41159);
nor U41745 (N_41745,N_41191,N_41081);
and U41746 (N_41746,N_41279,N_41278);
and U41747 (N_41747,N_41468,N_41306);
or U41748 (N_41748,N_41075,N_41070);
and U41749 (N_41749,N_41294,N_41305);
xor U41750 (N_41750,N_41307,N_41454);
nand U41751 (N_41751,N_41152,N_41305);
or U41752 (N_41752,N_41135,N_41061);
and U41753 (N_41753,N_41186,N_41361);
or U41754 (N_41754,N_41161,N_41023);
and U41755 (N_41755,N_41254,N_41188);
xnor U41756 (N_41756,N_41384,N_41264);
or U41757 (N_41757,N_41090,N_41360);
nor U41758 (N_41758,N_41192,N_41356);
nor U41759 (N_41759,N_41444,N_41072);
or U41760 (N_41760,N_41033,N_41411);
nand U41761 (N_41761,N_41066,N_41324);
xor U41762 (N_41762,N_41450,N_41322);
or U41763 (N_41763,N_41366,N_41293);
or U41764 (N_41764,N_41233,N_41026);
or U41765 (N_41765,N_41059,N_41058);
or U41766 (N_41766,N_41306,N_41351);
and U41767 (N_41767,N_41135,N_41143);
or U41768 (N_41768,N_41494,N_41133);
and U41769 (N_41769,N_41229,N_41354);
or U41770 (N_41770,N_41451,N_41049);
xnor U41771 (N_41771,N_41062,N_41401);
and U41772 (N_41772,N_41121,N_41045);
nor U41773 (N_41773,N_41272,N_41452);
and U41774 (N_41774,N_41123,N_41101);
nand U41775 (N_41775,N_41131,N_41005);
xor U41776 (N_41776,N_41262,N_41125);
and U41777 (N_41777,N_41494,N_41315);
nand U41778 (N_41778,N_41287,N_41052);
or U41779 (N_41779,N_41423,N_41056);
and U41780 (N_41780,N_41491,N_41188);
and U41781 (N_41781,N_41203,N_41108);
xnor U41782 (N_41782,N_41040,N_41059);
xnor U41783 (N_41783,N_41072,N_41362);
nand U41784 (N_41784,N_41055,N_41195);
nor U41785 (N_41785,N_41095,N_41457);
and U41786 (N_41786,N_41273,N_41148);
and U41787 (N_41787,N_41074,N_41077);
xnor U41788 (N_41788,N_41138,N_41426);
nor U41789 (N_41789,N_41297,N_41103);
nand U41790 (N_41790,N_41245,N_41083);
or U41791 (N_41791,N_41469,N_41005);
xor U41792 (N_41792,N_41340,N_41347);
nor U41793 (N_41793,N_41458,N_41499);
or U41794 (N_41794,N_41353,N_41046);
nor U41795 (N_41795,N_41461,N_41010);
xor U41796 (N_41796,N_41262,N_41448);
or U41797 (N_41797,N_41355,N_41082);
xnor U41798 (N_41798,N_41000,N_41005);
and U41799 (N_41799,N_41409,N_41182);
xnor U41800 (N_41800,N_41397,N_41371);
or U41801 (N_41801,N_41136,N_41343);
xor U41802 (N_41802,N_41393,N_41238);
nand U41803 (N_41803,N_41232,N_41284);
nor U41804 (N_41804,N_41097,N_41179);
xor U41805 (N_41805,N_41165,N_41047);
xor U41806 (N_41806,N_41177,N_41189);
nor U41807 (N_41807,N_41473,N_41453);
and U41808 (N_41808,N_41042,N_41017);
nor U41809 (N_41809,N_41223,N_41130);
and U41810 (N_41810,N_41123,N_41344);
nor U41811 (N_41811,N_41486,N_41473);
nand U41812 (N_41812,N_41319,N_41152);
xnor U41813 (N_41813,N_41044,N_41480);
and U41814 (N_41814,N_41010,N_41232);
and U41815 (N_41815,N_41458,N_41325);
xor U41816 (N_41816,N_41177,N_41457);
xor U41817 (N_41817,N_41015,N_41022);
xor U41818 (N_41818,N_41254,N_41004);
nor U41819 (N_41819,N_41338,N_41346);
nand U41820 (N_41820,N_41113,N_41319);
or U41821 (N_41821,N_41156,N_41399);
nand U41822 (N_41822,N_41082,N_41499);
and U41823 (N_41823,N_41122,N_41327);
xnor U41824 (N_41824,N_41474,N_41362);
nor U41825 (N_41825,N_41317,N_41181);
nand U41826 (N_41826,N_41374,N_41121);
xnor U41827 (N_41827,N_41097,N_41346);
nand U41828 (N_41828,N_41334,N_41177);
or U41829 (N_41829,N_41012,N_41258);
xnor U41830 (N_41830,N_41269,N_41371);
or U41831 (N_41831,N_41437,N_41330);
nand U41832 (N_41832,N_41411,N_41367);
and U41833 (N_41833,N_41014,N_41121);
or U41834 (N_41834,N_41311,N_41081);
or U41835 (N_41835,N_41386,N_41342);
or U41836 (N_41836,N_41029,N_41368);
or U41837 (N_41837,N_41027,N_41008);
and U41838 (N_41838,N_41304,N_41268);
nand U41839 (N_41839,N_41497,N_41499);
nand U41840 (N_41840,N_41201,N_41132);
or U41841 (N_41841,N_41349,N_41095);
nand U41842 (N_41842,N_41285,N_41017);
nand U41843 (N_41843,N_41347,N_41366);
nand U41844 (N_41844,N_41220,N_41223);
and U41845 (N_41845,N_41405,N_41113);
nand U41846 (N_41846,N_41084,N_41123);
and U41847 (N_41847,N_41129,N_41109);
and U41848 (N_41848,N_41156,N_41224);
nor U41849 (N_41849,N_41066,N_41264);
nor U41850 (N_41850,N_41472,N_41334);
and U41851 (N_41851,N_41030,N_41126);
nor U41852 (N_41852,N_41313,N_41401);
nor U41853 (N_41853,N_41395,N_41266);
nor U41854 (N_41854,N_41359,N_41130);
nor U41855 (N_41855,N_41498,N_41418);
nand U41856 (N_41856,N_41442,N_41002);
nand U41857 (N_41857,N_41428,N_41145);
xor U41858 (N_41858,N_41393,N_41216);
and U41859 (N_41859,N_41280,N_41103);
nor U41860 (N_41860,N_41122,N_41023);
nand U41861 (N_41861,N_41104,N_41013);
xnor U41862 (N_41862,N_41062,N_41183);
xor U41863 (N_41863,N_41425,N_41075);
and U41864 (N_41864,N_41258,N_41036);
xor U41865 (N_41865,N_41058,N_41008);
and U41866 (N_41866,N_41013,N_41247);
nand U41867 (N_41867,N_41377,N_41433);
and U41868 (N_41868,N_41313,N_41069);
and U41869 (N_41869,N_41339,N_41341);
xor U41870 (N_41870,N_41184,N_41037);
or U41871 (N_41871,N_41168,N_41052);
and U41872 (N_41872,N_41492,N_41238);
xnor U41873 (N_41873,N_41298,N_41478);
and U41874 (N_41874,N_41134,N_41209);
nor U41875 (N_41875,N_41425,N_41008);
nand U41876 (N_41876,N_41304,N_41028);
xor U41877 (N_41877,N_41198,N_41080);
or U41878 (N_41878,N_41419,N_41049);
and U41879 (N_41879,N_41390,N_41017);
and U41880 (N_41880,N_41347,N_41327);
nand U41881 (N_41881,N_41376,N_41484);
nand U41882 (N_41882,N_41385,N_41211);
nand U41883 (N_41883,N_41200,N_41306);
or U41884 (N_41884,N_41188,N_41335);
nor U41885 (N_41885,N_41150,N_41444);
nor U41886 (N_41886,N_41376,N_41172);
or U41887 (N_41887,N_41470,N_41286);
nand U41888 (N_41888,N_41056,N_41219);
xnor U41889 (N_41889,N_41172,N_41355);
xor U41890 (N_41890,N_41109,N_41063);
and U41891 (N_41891,N_41192,N_41286);
nand U41892 (N_41892,N_41266,N_41462);
xor U41893 (N_41893,N_41468,N_41373);
and U41894 (N_41894,N_41105,N_41221);
or U41895 (N_41895,N_41485,N_41037);
or U41896 (N_41896,N_41043,N_41160);
nor U41897 (N_41897,N_41017,N_41290);
nand U41898 (N_41898,N_41231,N_41326);
nand U41899 (N_41899,N_41207,N_41454);
and U41900 (N_41900,N_41141,N_41262);
nand U41901 (N_41901,N_41010,N_41065);
and U41902 (N_41902,N_41107,N_41414);
nor U41903 (N_41903,N_41376,N_41301);
or U41904 (N_41904,N_41362,N_41060);
and U41905 (N_41905,N_41340,N_41018);
or U41906 (N_41906,N_41111,N_41280);
or U41907 (N_41907,N_41492,N_41108);
xnor U41908 (N_41908,N_41499,N_41443);
nand U41909 (N_41909,N_41428,N_41284);
and U41910 (N_41910,N_41492,N_41345);
nor U41911 (N_41911,N_41469,N_41435);
xnor U41912 (N_41912,N_41472,N_41139);
or U41913 (N_41913,N_41423,N_41079);
xnor U41914 (N_41914,N_41331,N_41078);
nand U41915 (N_41915,N_41481,N_41039);
nand U41916 (N_41916,N_41160,N_41165);
xnor U41917 (N_41917,N_41013,N_41246);
nand U41918 (N_41918,N_41472,N_41229);
nor U41919 (N_41919,N_41012,N_41436);
or U41920 (N_41920,N_41265,N_41010);
xnor U41921 (N_41921,N_41207,N_41182);
nand U41922 (N_41922,N_41228,N_41084);
nor U41923 (N_41923,N_41324,N_41418);
nor U41924 (N_41924,N_41218,N_41461);
nand U41925 (N_41925,N_41267,N_41124);
or U41926 (N_41926,N_41111,N_41024);
or U41927 (N_41927,N_41433,N_41455);
xor U41928 (N_41928,N_41217,N_41260);
xnor U41929 (N_41929,N_41134,N_41380);
nor U41930 (N_41930,N_41421,N_41338);
or U41931 (N_41931,N_41236,N_41345);
xor U41932 (N_41932,N_41173,N_41236);
xnor U41933 (N_41933,N_41222,N_41014);
and U41934 (N_41934,N_41294,N_41193);
nor U41935 (N_41935,N_41326,N_41265);
nor U41936 (N_41936,N_41139,N_41487);
and U41937 (N_41937,N_41254,N_41147);
xnor U41938 (N_41938,N_41167,N_41407);
nand U41939 (N_41939,N_41494,N_41466);
xnor U41940 (N_41940,N_41179,N_41413);
xnor U41941 (N_41941,N_41239,N_41188);
nand U41942 (N_41942,N_41140,N_41368);
xor U41943 (N_41943,N_41348,N_41491);
nor U41944 (N_41944,N_41132,N_41183);
and U41945 (N_41945,N_41102,N_41072);
xnor U41946 (N_41946,N_41355,N_41350);
and U41947 (N_41947,N_41125,N_41244);
nor U41948 (N_41948,N_41069,N_41273);
nor U41949 (N_41949,N_41026,N_41430);
or U41950 (N_41950,N_41341,N_41370);
nand U41951 (N_41951,N_41217,N_41037);
and U41952 (N_41952,N_41408,N_41394);
and U41953 (N_41953,N_41097,N_41343);
nor U41954 (N_41954,N_41233,N_41053);
and U41955 (N_41955,N_41073,N_41477);
and U41956 (N_41956,N_41325,N_41198);
and U41957 (N_41957,N_41032,N_41430);
and U41958 (N_41958,N_41214,N_41032);
and U41959 (N_41959,N_41163,N_41420);
xor U41960 (N_41960,N_41285,N_41071);
and U41961 (N_41961,N_41374,N_41077);
nor U41962 (N_41962,N_41246,N_41308);
nor U41963 (N_41963,N_41001,N_41033);
and U41964 (N_41964,N_41370,N_41337);
nand U41965 (N_41965,N_41474,N_41023);
and U41966 (N_41966,N_41135,N_41469);
or U41967 (N_41967,N_41284,N_41249);
or U41968 (N_41968,N_41187,N_41408);
and U41969 (N_41969,N_41023,N_41316);
or U41970 (N_41970,N_41416,N_41403);
nand U41971 (N_41971,N_41200,N_41484);
nor U41972 (N_41972,N_41179,N_41492);
xnor U41973 (N_41973,N_41372,N_41004);
nor U41974 (N_41974,N_41460,N_41171);
nand U41975 (N_41975,N_41442,N_41280);
nor U41976 (N_41976,N_41152,N_41200);
or U41977 (N_41977,N_41487,N_41176);
or U41978 (N_41978,N_41221,N_41204);
and U41979 (N_41979,N_41225,N_41135);
xnor U41980 (N_41980,N_41330,N_41472);
and U41981 (N_41981,N_41408,N_41170);
nand U41982 (N_41982,N_41295,N_41155);
xor U41983 (N_41983,N_41434,N_41166);
or U41984 (N_41984,N_41362,N_41304);
xor U41985 (N_41985,N_41472,N_41207);
xor U41986 (N_41986,N_41317,N_41498);
nor U41987 (N_41987,N_41336,N_41427);
nor U41988 (N_41988,N_41349,N_41445);
and U41989 (N_41989,N_41474,N_41244);
and U41990 (N_41990,N_41387,N_41494);
xnor U41991 (N_41991,N_41111,N_41281);
nor U41992 (N_41992,N_41268,N_41247);
or U41993 (N_41993,N_41330,N_41449);
xnor U41994 (N_41994,N_41319,N_41421);
nor U41995 (N_41995,N_41497,N_41204);
and U41996 (N_41996,N_41485,N_41002);
nand U41997 (N_41997,N_41034,N_41159);
or U41998 (N_41998,N_41046,N_41371);
xor U41999 (N_41999,N_41323,N_41121);
nor U42000 (N_42000,N_41614,N_41805);
and U42001 (N_42001,N_41511,N_41735);
nand U42002 (N_42002,N_41709,N_41727);
nand U42003 (N_42003,N_41571,N_41757);
xor U42004 (N_42004,N_41711,N_41885);
xor U42005 (N_42005,N_41586,N_41626);
and U42006 (N_42006,N_41965,N_41654);
nor U42007 (N_42007,N_41613,N_41978);
and U42008 (N_42008,N_41646,N_41559);
and U42009 (N_42009,N_41828,N_41523);
xnor U42010 (N_42010,N_41503,N_41685);
nor U42011 (N_42011,N_41909,N_41898);
and U42012 (N_42012,N_41619,N_41667);
xnor U42013 (N_42013,N_41836,N_41684);
xnor U42014 (N_42014,N_41821,N_41532);
nand U42015 (N_42015,N_41873,N_41699);
or U42016 (N_42016,N_41793,N_41715);
and U42017 (N_42017,N_41723,N_41950);
or U42018 (N_42018,N_41913,N_41714);
and U42019 (N_42019,N_41765,N_41809);
or U42020 (N_42020,N_41760,N_41674);
and U42021 (N_42021,N_41956,N_41948);
xnor U42022 (N_42022,N_41936,N_41697);
xor U42023 (N_42023,N_41591,N_41678);
nand U42024 (N_42024,N_41533,N_41624);
xnor U42025 (N_42025,N_41790,N_41534);
nand U42026 (N_42026,N_41638,N_41955);
or U42027 (N_42027,N_41739,N_41866);
nor U42028 (N_42028,N_41995,N_41600);
or U42029 (N_42029,N_41680,N_41817);
and U42030 (N_42030,N_41939,N_41721);
nor U42031 (N_42031,N_41779,N_41850);
xor U42032 (N_42032,N_41629,N_41831);
nor U42033 (N_42033,N_41710,N_41700);
xor U42034 (N_42034,N_41754,N_41857);
or U42035 (N_42035,N_41780,N_41887);
and U42036 (N_42036,N_41751,N_41753);
nor U42037 (N_42037,N_41900,N_41545);
nor U42038 (N_42038,N_41968,N_41679);
and U42039 (N_42039,N_41612,N_41557);
or U42040 (N_42040,N_41564,N_41724);
xnor U42041 (N_42041,N_41840,N_41568);
nand U42042 (N_42042,N_41962,N_41693);
and U42043 (N_42043,N_41588,N_41556);
and U42044 (N_42044,N_41830,N_41759);
xnor U42045 (N_42045,N_41903,N_41905);
nor U42046 (N_42046,N_41774,N_41964);
nor U42047 (N_42047,N_41932,N_41746);
nor U42048 (N_42048,N_41620,N_41871);
and U42049 (N_42049,N_41637,N_41756);
nor U42050 (N_42050,N_41931,N_41703);
nand U42051 (N_42051,N_41917,N_41601);
nor U42052 (N_42052,N_41843,N_41888);
and U42053 (N_42053,N_41642,N_41550);
xor U42054 (N_42054,N_41512,N_41648);
xnor U42055 (N_42055,N_41846,N_41582);
nand U42056 (N_42056,N_41940,N_41918);
nand U42057 (N_42057,N_41824,N_41854);
nor U42058 (N_42058,N_41785,N_41596);
nand U42059 (N_42059,N_41827,N_41838);
and U42060 (N_42060,N_41635,N_41676);
or U42061 (N_42061,N_41848,N_41755);
and U42062 (N_42062,N_41945,N_41907);
or U42063 (N_42063,N_41623,N_41897);
nand U42064 (N_42064,N_41593,N_41603);
nor U42065 (N_42065,N_41504,N_41875);
nand U42066 (N_42066,N_41772,N_41664);
and U42067 (N_42067,N_41926,N_41781);
nand U42068 (N_42068,N_41577,N_41608);
or U42069 (N_42069,N_41858,N_41740);
xnor U42070 (N_42070,N_41972,N_41585);
xor U42071 (N_42071,N_41802,N_41743);
nor U42072 (N_42072,N_41561,N_41544);
and U42073 (N_42073,N_41555,N_41868);
nor U42074 (N_42074,N_41653,N_41528);
or U42075 (N_42075,N_41876,N_41801);
or U42076 (N_42076,N_41563,N_41869);
nor U42077 (N_42077,N_41922,N_41736);
and U42078 (N_42078,N_41598,N_41645);
and U42079 (N_42079,N_41804,N_41763);
nor U42080 (N_42080,N_41764,N_41670);
nor U42081 (N_42081,N_41811,N_41967);
nand U42082 (N_42082,N_41716,N_41651);
and U42083 (N_42083,N_41722,N_41702);
xnor U42084 (N_42084,N_41852,N_41777);
nor U42085 (N_42085,N_41853,N_41656);
and U42086 (N_42086,N_41971,N_41986);
xor U42087 (N_42087,N_41649,N_41881);
xnor U42088 (N_42088,N_41732,N_41813);
nand U42089 (N_42089,N_41610,N_41961);
nand U42090 (N_42090,N_41604,N_41923);
nor U42091 (N_42091,N_41818,N_41566);
or U42092 (N_42092,N_41867,N_41558);
nand U42093 (N_42093,N_41959,N_41856);
xnor U42094 (N_42094,N_41597,N_41643);
and U42095 (N_42095,N_41944,N_41847);
nand U42096 (N_42096,N_41509,N_41865);
xnor U42097 (N_42097,N_41560,N_41992);
and U42098 (N_42098,N_41542,N_41578);
xnor U42099 (N_42099,N_41834,N_41652);
xor U42100 (N_42100,N_41730,N_41541);
nand U42101 (N_42101,N_41718,N_41663);
nor U42102 (N_42102,N_41641,N_41636);
nor U42103 (N_42103,N_41567,N_41919);
xor U42104 (N_42104,N_41605,N_41606);
xnor U42105 (N_42105,N_41647,N_41627);
nand U42106 (N_42106,N_41969,N_41799);
nand U42107 (N_42107,N_41726,N_41698);
or U42108 (N_42108,N_41675,N_41942);
nand U42109 (N_42109,N_41958,N_41729);
or U42110 (N_42110,N_41569,N_41974);
or U42111 (N_42111,N_41806,N_41659);
nand U42112 (N_42112,N_41607,N_41531);
xnor U42113 (N_42113,N_41796,N_41516);
xnor U42114 (N_42114,N_41937,N_41951);
nor U42115 (N_42115,N_41895,N_41547);
nor U42116 (N_42116,N_41631,N_41935);
nor U42117 (N_42117,N_41855,N_41553);
xor U42118 (N_42118,N_41946,N_41771);
nand U42119 (N_42119,N_41690,N_41508);
and U42120 (N_42120,N_41835,N_41632);
or U42121 (N_42121,N_41924,N_41930);
xnor U42122 (N_42122,N_41878,N_41841);
nand U42123 (N_42123,N_41860,N_41506);
xnor U42124 (N_42124,N_41904,N_41691);
nand U42125 (N_42125,N_41800,N_41581);
xnor U42126 (N_42126,N_41928,N_41524);
and U42127 (N_42127,N_41826,N_41748);
xnor U42128 (N_42128,N_41915,N_41775);
or U42129 (N_42129,N_41769,N_41982);
or U42130 (N_42130,N_41773,N_41546);
or U42131 (N_42131,N_41551,N_41692);
and U42132 (N_42132,N_41750,N_41980);
nand U42133 (N_42133,N_41701,N_41807);
and U42134 (N_42134,N_41966,N_41872);
or U42135 (N_42135,N_41639,N_41910);
xnor U42136 (N_42136,N_41745,N_41877);
or U42137 (N_42137,N_41576,N_41505);
xnor U42138 (N_42138,N_41665,N_41975);
or U42139 (N_42139,N_41921,N_41795);
and U42140 (N_42140,N_41517,N_41993);
and U42141 (N_42141,N_41687,N_41666);
nand U42142 (N_42142,N_41814,N_41999);
xor U42143 (N_42143,N_41574,N_41625);
nand U42144 (N_42144,N_41941,N_41733);
xor U42145 (N_42145,N_41671,N_41812);
xor U42146 (N_42146,N_41741,N_41529);
xnor U42147 (N_42147,N_41535,N_41514);
nor U42148 (N_42148,N_41552,N_41633);
nor U42149 (N_42149,N_41902,N_41719);
nor U42150 (N_42150,N_41851,N_41880);
xor U42151 (N_42151,N_41996,N_41766);
nand U42152 (N_42152,N_41893,N_41889);
or U42153 (N_42153,N_41500,N_41984);
nor U42154 (N_42154,N_41983,N_41960);
or U42155 (N_42155,N_41820,N_41837);
nand U42156 (N_42156,N_41655,N_41554);
xnor U42157 (N_42157,N_41762,N_41594);
and U42158 (N_42158,N_41879,N_41658);
xor U42159 (N_42159,N_41768,N_41536);
nor U42160 (N_42160,N_41518,N_41938);
and U42161 (N_42161,N_41522,N_41704);
and U42162 (N_42162,N_41862,N_41849);
xnor U42163 (N_42163,N_41525,N_41979);
xor U42164 (N_42164,N_41815,N_41792);
xor U42165 (N_42165,N_41891,N_41839);
or U42166 (N_42166,N_41808,N_41803);
nand U42167 (N_42167,N_41816,N_41713);
nand U42168 (N_42168,N_41537,N_41989);
xnor U42169 (N_42169,N_41747,N_41530);
nor U42170 (N_42170,N_41997,N_41844);
and U42171 (N_42171,N_41543,N_41916);
nor U42172 (N_42172,N_41681,N_41778);
or U42173 (N_42173,N_41595,N_41977);
or U42174 (N_42174,N_41527,N_41616);
nor U42175 (N_42175,N_41819,N_41519);
xor U42176 (N_42176,N_41584,N_41521);
and U42177 (N_42177,N_41720,N_41987);
nor U42178 (N_42178,N_41717,N_41611);
or U42179 (N_42179,N_41782,N_41863);
or U42180 (N_42180,N_41575,N_41660);
or U42181 (N_42181,N_41954,N_41731);
xnor U42182 (N_42182,N_41749,N_41973);
and U42183 (N_42183,N_41617,N_41609);
xnor U42184 (N_42184,N_41657,N_41630);
and U42185 (N_42185,N_41672,N_41833);
nand U42186 (N_42186,N_41640,N_41510);
or U42187 (N_42187,N_41602,N_41583);
xor U42188 (N_42188,N_41507,N_41894);
and U42189 (N_42189,N_41914,N_41562);
and U42190 (N_42190,N_41538,N_41580);
nand U42191 (N_42191,N_41688,N_41761);
xor U42192 (N_42192,N_41682,N_41952);
and U42193 (N_42193,N_41695,N_41892);
nand U42194 (N_42194,N_41883,N_41920);
nor U42195 (N_42195,N_41644,N_41970);
or U42196 (N_42196,N_41789,N_41994);
xor U42197 (N_42197,N_41615,N_41696);
and U42198 (N_42198,N_41985,N_41686);
nor U42199 (N_42199,N_41549,N_41845);
xnor U42200 (N_42200,N_41791,N_41988);
xor U42201 (N_42201,N_41502,N_41798);
or U42202 (N_42202,N_41933,N_41998);
and U42203 (N_42203,N_41829,N_41823);
or U42204 (N_42204,N_41662,N_41925);
or U42205 (N_42205,N_41783,N_41573);
nor U42206 (N_42206,N_41787,N_41899);
xor U42207 (N_42207,N_41874,N_41784);
nor U42208 (N_42208,N_41981,N_41515);
nor U42209 (N_42209,N_41650,N_41842);
and U42210 (N_42210,N_41520,N_41929);
xor U42211 (N_42211,N_41683,N_41884);
xor U42212 (N_42212,N_41943,N_41694);
nand U42213 (N_42213,N_41908,N_41599);
and U42214 (N_42214,N_41728,N_41707);
and U42215 (N_42215,N_41708,N_41861);
nand U42216 (N_42216,N_41734,N_41621);
nand U42217 (N_42217,N_41870,N_41770);
and U42218 (N_42218,N_41767,N_41579);
and U42219 (N_42219,N_41668,N_41526);
or U42220 (N_42220,N_41622,N_41991);
xnor U42221 (N_42221,N_41587,N_41976);
or U42222 (N_42222,N_41912,N_41797);
nand U42223 (N_42223,N_41661,N_41669);
and U42224 (N_42224,N_41513,N_41825);
nand U42225 (N_42225,N_41628,N_41786);
xnor U42226 (N_42226,N_41752,N_41957);
nor U42227 (N_42227,N_41953,N_41927);
nor U42228 (N_42228,N_41744,N_41832);
nor U42229 (N_42229,N_41934,N_41572);
or U42230 (N_42230,N_41864,N_41990);
and U42231 (N_42231,N_41589,N_41570);
nor U42232 (N_42232,N_41859,N_41592);
and U42233 (N_42233,N_41822,N_41882);
nand U42234 (N_42234,N_41548,N_41886);
nor U42235 (N_42235,N_41712,N_41738);
nor U42236 (N_42236,N_41949,N_41947);
or U42237 (N_42237,N_41742,N_41963);
or U42238 (N_42238,N_41776,N_41794);
xnor U42239 (N_42239,N_41677,N_41689);
xor U42240 (N_42240,N_41705,N_41890);
and U42241 (N_42241,N_41590,N_41618);
nand U42242 (N_42242,N_41706,N_41565);
nor U42243 (N_42243,N_41901,N_41810);
nor U42244 (N_42244,N_41737,N_41758);
nor U42245 (N_42245,N_41673,N_41634);
or U42246 (N_42246,N_41725,N_41788);
xnor U42247 (N_42247,N_41501,N_41906);
nand U42248 (N_42248,N_41540,N_41896);
xor U42249 (N_42249,N_41911,N_41539);
or U42250 (N_42250,N_41689,N_41729);
xnor U42251 (N_42251,N_41927,N_41618);
xor U42252 (N_42252,N_41575,N_41970);
xor U42253 (N_42253,N_41765,N_41577);
or U42254 (N_42254,N_41613,N_41965);
or U42255 (N_42255,N_41904,N_41709);
or U42256 (N_42256,N_41773,N_41611);
and U42257 (N_42257,N_41646,N_41594);
or U42258 (N_42258,N_41608,N_41967);
nand U42259 (N_42259,N_41571,N_41610);
nand U42260 (N_42260,N_41766,N_41586);
nor U42261 (N_42261,N_41559,N_41653);
or U42262 (N_42262,N_41658,N_41765);
or U42263 (N_42263,N_41829,N_41950);
nor U42264 (N_42264,N_41575,N_41975);
nand U42265 (N_42265,N_41933,N_41542);
or U42266 (N_42266,N_41764,N_41805);
or U42267 (N_42267,N_41703,N_41746);
nand U42268 (N_42268,N_41524,N_41812);
nor U42269 (N_42269,N_41701,N_41772);
nor U42270 (N_42270,N_41622,N_41705);
nand U42271 (N_42271,N_41960,N_41922);
and U42272 (N_42272,N_41660,N_41692);
and U42273 (N_42273,N_41644,N_41572);
and U42274 (N_42274,N_41610,N_41614);
nor U42275 (N_42275,N_41874,N_41514);
and U42276 (N_42276,N_41807,N_41536);
nor U42277 (N_42277,N_41687,N_41842);
xor U42278 (N_42278,N_41569,N_41730);
nor U42279 (N_42279,N_41948,N_41599);
or U42280 (N_42280,N_41846,N_41701);
or U42281 (N_42281,N_41759,N_41695);
and U42282 (N_42282,N_41968,N_41619);
nor U42283 (N_42283,N_41825,N_41551);
or U42284 (N_42284,N_41740,N_41549);
xnor U42285 (N_42285,N_41881,N_41755);
or U42286 (N_42286,N_41929,N_41763);
xor U42287 (N_42287,N_41840,N_41900);
and U42288 (N_42288,N_41677,N_41923);
or U42289 (N_42289,N_41634,N_41730);
and U42290 (N_42290,N_41666,N_41721);
and U42291 (N_42291,N_41598,N_41676);
xnor U42292 (N_42292,N_41641,N_41724);
nand U42293 (N_42293,N_41532,N_41550);
xnor U42294 (N_42294,N_41635,N_41941);
nor U42295 (N_42295,N_41702,N_41864);
nand U42296 (N_42296,N_41829,N_41558);
xor U42297 (N_42297,N_41636,N_41749);
nand U42298 (N_42298,N_41641,N_41596);
or U42299 (N_42299,N_41955,N_41637);
nor U42300 (N_42300,N_41655,N_41914);
nor U42301 (N_42301,N_41702,N_41536);
xor U42302 (N_42302,N_41616,N_41994);
nor U42303 (N_42303,N_41882,N_41759);
and U42304 (N_42304,N_41828,N_41991);
or U42305 (N_42305,N_41834,N_41999);
xor U42306 (N_42306,N_41505,N_41513);
nor U42307 (N_42307,N_41571,N_41659);
and U42308 (N_42308,N_41752,N_41602);
nor U42309 (N_42309,N_41622,N_41751);
and U42310 (N_42310,N_41999,N_41827);
nand U42311 (N_42311,N_41844,N_41588);
nor U42312 (N_42312,N_41919,N_41624);
nor U42313 (N_42313,N_41538,N_41996);
and U42314 (N_42314,N_41714,N_41632);
and U42315 (N_42315,N_41693,N_41957);
nor U42316 (N_42316,N_41683,N_41718);
nor U42317 (N_42317,N_41927,N_41776);
and U42318 (N_42318,N_41752,N_41748);
xor U42319 (N_42319,N_41657,N_41517);
nand U42320 (N_42320,N_41799,N_41782);
nor U42321 (N_42321,N_41704,N_41922);
and U42322 (N_42322,N_41521,N_41908);
or U42323 (N_42323,N_41729,N_41979);
nor U42324 (N_42324,N_41804,N_41752);
and U42325 (N_42325,N_41653,N_41598);
nand U42326 (N_42326,N_41819,N_41654);
xnor U42327 (N_42327,N_41769,N_41721);
nor U42328 (N_42328,N_41533,N_41586);
nor U42329 (N_42329,N_41715,N_41814);
and U42330 (N_42330,N_41992,N_41910);
or U42331 (N_42331,N_41670,N_41860);
nand U42332 (N_42332,N_41730,N_41705);
or U42333 (N_42333,N_41901,N_41862);
nand U42334 (N_42334,N_41657,N_41690);
nand U42335 (N_42335,N_41681,N_41932);
and U42336 (N_42336,N_41704,N_41557);
or U42337 (N_42337,N_41614,N_41532);
nand U42338 (N_42338,N_41503,N_41885);
or U42339 (N_42339,N_41870,N_41905);
or U42340 (N_42340,N_41856,N_41613);
nand U42341 (N_42341,N_41792,N_41996);
nor U42342 (N_42342,N_41802,N_41523);
nand U42343 (N_42343,N_41765,N_41791);
or U42344 (N_42344,N_41698,N_41759);
and U42345 (N_42345,N_41513,N_41618);
nand U42346 (N_42346,N_41882,N_41903);
or U42347 (N_42347,N_41988,N_41998);
nor U42348 (N_42348,N_41759,N_41995);
xor U42349 (N_42349,N_41801,N_41992);
nand U42350 (N_42350,N_41826,N_41792);
xnor U42351 (N_42351,N_41669,N_41619);
and U42352 (N_42352,N_41779,N_41570);
or U42353 (N_42353,N_41717,N_41671);
nand U42354 (N_42354,N_41619,N_41783);
xnor U42355 (N_42355,N_41924,N_41941);
nand U42356 (N_42356,N_41901,N_41779);
xnor U42357 (N_42357,N_41859,N_41836);
or U42358 (N_42358,N_41528,N_41996);
and U42359 (N_42359,N_41924,N_41611);
or U42360 (N_42360,N_41605,N_41826);
and U42361 (N_42361,N_41753,N_41514);
nor U42362 (N_42362,N_41982,N_41711);
nand U42363 (N_42363,N_41884,N_41593);
or U42364 (N_42364,N_41557,N_41850);
nand U42365 (N_42365,N_41948,N_41708);
or U42366 (N_42366,N_41801,N_41878);
or U42367 (N_42367,N_41886,N_41539);
or U42368 (N_42368,N_41817,N_41832);
xnor U42369 (N_42369,N_41807,N_41720);
nand U42370 (N_42370,N_41668,N_41958);
and U42371 (N_42371,N_41648,N_41767);
and U42372 (N_42372,N_41949,N_41614);
or U42373 (N_42373,N_41864,N_41758);
xnor U42374 (N_42374,N_41906,N_41523);
nand U42375 (N_42375,N_41715,N_41666);
nor U42376 (N_42376,N_41848,N_41983);
xnor U42377 (N_42377,N_41777,N_41627);
nor U42378 (N_42378,N_41586,N_41786);
or U42379 (N_42379,N_41706,N_41801);
xnor U42380 (N_42380,N_41531,N_41589);
or U42381 (N_42381,N_41563,N_41816);
and U42382 (N_42382,N_41881,N_41626);
nand U42383 (N_42383,N_41660,N_41714);
nor U42384 (N_42384,N_41724,N_41791);
nor U42385 (N_42385,N_41977,N_41640);
and U42386 (N_42386,N_41862,N_41507);
and U42387 (N_42387,N_41571,N_41792);
and U42388 (N_42388,N_41629,N_41741);
or U42389 (N_42389,N_41648,N_41735);
and U42390 (N_42390,N_41727,N_41968);
or U42391 (N_42391,N_41703,N_41573);
nand U42392 (N_42392,N_41813,N_41712);
nand U42393 (N_42393,N_41750,N_41792);
nor U42394 (N_42394,N_41765,N_41959);
and U42395 (N_42395,N_41624,N_41732);
or U42396 (N_42396,N_41631,N_41595);
and U42397 (N_42397,N_41631,N_41977);
or U42398 (N_42398,N_41869,N_41999);
and U42399 (N_42399,N_41857,N_41863);
xor U42400 (N_42400,N_41785,N_41770);
or U42401 (N_42401,N_41775,N_41900);
nand U42402 (N_42402,N_41754,N_41625);
nand U42403 (N_42403,N_41677,N_41566);
or U42404 (N_42404,N_41744,N_41917);
and U42405 (N_42405,N_41668,N_41790);
xnor U42406 (N_42406,N_41687,N_41553);
nor U42407 (N_42407,N_41711,N_41802);
nor U42408 (N_42408,N_41683,N_41971);
nand U42409 (N_42409,N_41658,N_41988);
or U42410 (N_42410,N_41696,N_41588);
nand U42411 (N_42411,N_41918,N_41658);
xnor U42412 (N_42412,N_41571,N_41630);
and U42413 (N_42413,N_41512,N_41802);
nor U42414 (N_42414,N_41590,N_41808);
nand U42415 (N_42415,N_41565,N_41616);
or U42416 (N_42416,N_41649,N_41808);
and U42417 (N_42417,N_41697,N_41545);
nor U42418 (N_42418,N_41980,N_41805);
nor U42419 (N_42419,N_41523,N_41946);
nor U42420 (N_42420,N_41908,N_41744);
or U42421 (N_42421,N_41513,N_41511);
nand U42422 (N_42422,N_41982,N_41617);
or U42423 (N_42423,N_41824,N_41715);
xor U42424 (N_42424,N_41940,N_41873);
or U42425 (N_42425,N_41751,N_41565);
and U42426 (N_42426,N_41790,N_41526);
xor U42427 (N_42427,N_41770,N_41934);
nor U42428 (N_42428,N_41583,N_41920);
or U42429 (N_42429,N_41869,N_41862);
or U42430 (N_42430,N_41884,N_41774);
nor U42431 (N_42431,N_41597,N_41836);
xnor U42432 (N_42432,N_41503,N_41521);
and U42433 (N_42433,N_41970,N_41726);
or U42434 (N_42434,N_41604,N_41834);
and U42435 (N_42435,N_41964,N_41550);
nand U42436 (N_42436,N_41792,N_41963);
xnor U42437 (N_42437,N_41899,N_41718);
or U42438 (N_42438,N_41949,N_41504);
xnor U42439 (N_42439,N_41695,N_41596);
xor U42440 (N_42440,N_41686,N_41695);
nor U42441 (N_42441,N_41732,N_41582);
and U42442 (N_42442,N_41819,N_41875);
nor U42443 (N_42443,N_41673,N_41642);
or U42444 (N_42444,N_41511,N_41939);
and U42445 (N_42445,N_41569,N_41589);
nor U42446 (N_42446,N_41639,N_41567);
and U42447 (N_42447,N_41653,N_41734);
nand U42448 (N_42448,N_41678,N_41802);
or U42449 (N_42449,N_41818,N_41809);
and U42450 (N_42450,N_41975,N_41724);
xnor U42451 (N_42451,N_41740,N_41916);
or U42452 (N_42452,N_41597,N_41563);
or U42453 (N_42453,N_41543,N_41767);
and U42454 (N_42454,N_41822,N_41896);
nor U42455 (N_42455,N_41734,N_41529);
and U42456 (N_42456,N_41718,N_41706);
xnor U42457 (N_42457,N_41775,N_41796);
or U42458 (N_42458,N_41842,N_41691);
nand U42459 (N_42459,N_41781,N_41862);
nand U42460 (N_42460,N_41676,N_41677);
nand U42461 (N_42461,N_41944,N_41526);
and U42462 (N_42462,N_41805,N_41662);
nor U42463 (N_42463,N_41849,N_41856);
and U42464 (N_42464,N_41662,N_41940);
nor U42465 (N_42465,N_41708,N_41821);
xnor U42466 (N_42466,N_41940,N_41903);
and U42467 (N_42467,N_41723,N_41656);
nor U42468 (N_42468,N_41781,N_41571);
and U42469 (N_42469,N_41573,N_41730);
and U42470 (N_42470,N_41583,N_41703);
or U42471 (N_42471,N_41813,N_41623);
xnor U42472 (N_42472,N_41597,N_41997);
or U42473 (N_42473,N_41613,N_41966);
nor U42474 (N_42474,N_41595,N_41810);
xor U42475 (N_42475,N_41844,N_41861);
xnor U42476 (N_42476,N_41733,N_41538);
or U42477 (N_42477,N_41540,N_41956);
and U42478 (N_42478,N_41751,N_41791);
nand U42479 (N_42479,N_41909,N_41920);
or U42480 (N_42480,N_41802,N_41776);
and U42481 (N_42481,N_41910,N_41930);
nor U42482 (N_42482,N_41848,N_41571);
nor U42483 (N_42483,N_41516,N_41692);
and U42484 (N_42484,N_41602,N_41963);
nand U42485 (N_42485,N_41742,N_41745);
and U42486 (N_42486,N_41756,N_41523);
and U42487 (N_42487,N_41584,N_41531);
nand U42488 (N_42488,N_41723,N_41501);
or U42489 (N_42489,N_41739,N_41775);
or U42490 (N_42490,N_41947,N_41733);
nand U42491 (N_42491,N_41649,N_41930);
or U42492 (N_42492,N_41675,N_41596);
nor U42493 (N_42493,N_41689,N_41742);
and U42494 (N_42494,N_41504,N_41518);
nand U42495 (N_42495,N_41701,N_41965);
or U42496 (N_42496,N_41969,N_41922);
nand U42497 (N_42497,N_41581,N_41553);
nor U42498 (N_42498,N_41680,N_41913);
and U42499 (N_42499,N_41581,N_41692);
and U42500 (N_42500,N_42048,N_42088);
and U42501 (N_42501,N_42191,N_42238);
xnor U42502 (N_42502,N_42265,N_42372);
nor U42503 (N_42503,N_42051,N_42195);
nand U42504 (N_42504,N_42405,N_42093);
nor U42505 (N_42505,N_42327,N_42024);
nand U42506 (N_42506,N_42062,N_42146);
nand U42507 (N_42507,N_42494,N_42425);
or U42508 (N_42508,N_42483,N_42039);
or U42509 (N_42509,N_42326,N_42204);
nand U42510 (N_42510,N_42015,N_42286);
nand U42511 (N_42511,N_42356,N_42205);
or U42512 (N_42512,N_42177,N_42236);
xnor U42513 (N_42513,N_42192,N_42431);
xor U42514 (N_42514,N_42404,N_42147);
xor U42515 (N_42515,N_42008,N_42428);
nand U42516 (N_42516,N_42346,N_42374);
nor U42517 (N_42517,N_42475,N_42268);
or U42518 (N_42518,N_42432,N_42173);
and U42519 (N_42519,N_42190,N_42114);
or U42520 (N_42520,N_42399,N_42160);
and U42521 (N_42521,N_42193,N_42186);
nor U42522 (N_42522,N_42396,N_42227);
nand U42523 (N_42523,N_42184,N_42077);
xnor U42524 (N_42524,N_42253,N_42031);
and U42525 (N_42525,N_42115,N_42306);
nor U42526 (N_42526,N_42493,N_42068);
or U42527 (N_42527,N_42437,N_42163);
and U42528 (N_42528,N_42004,N_42162);
nor U42529 (N_42529,N_42267,N_42311);
xnor U42530 (N_42530,N_42188,N_42079);
or U42531 (N_42531,N_42148,N_42445);
nand U42532 (N_42532,N_42002,N_42156);
or U42533 (N_42533,N_42413,N_42053);
nand U42534 (N_42534,N_42187,N_42000);
nand U42535 (N_42535,N_42451,N_42076);
xor U42536 (N_42536,N_42397,N_42219);
xor U42537 (N_42537,N_42270,N_42119);
and U42538 (N_42538,N_42474,N_42018);
nor U42539 (N_42539,N_42304,N_42027);
nand U42540 (N_42540,N_42151,N_42030);
or U42541 (N_42541,N_42172,N_42106);
nor U42542 (N_42542,N_42370,N_42387);
or U42543 (N_42543,N_42298,N_42411);
and U42544 (N_42544,N_42368,N_42080);
xnor U42545 (N_42545,N_42276,N_42386);
or U42546 (N_42546,N_42479,N_42121);
xnor U42547 (N_42547,N_42029,N_42330);
or U42548 (N_42548,N_42460,N_42241);
nand U42549 (N_42549,N_42215,N_42013);
nand U42550 (N_42550,N_42033,N_42367);
xor U42551 (N_42551,N_42357,N_42258);
and U42552 (N_42552,N_42273,N_42005);
nand U42553 (N_42553,N_42045,N_42351);
xor U42554 (N_42554,N_42251,N_42320);
xor U42555 (N_42555,N_42266,N_42426);
nand U42556 (N_42556,N_42061,N_42429);
and U42557 (N_42557,N_42279,N_42323);
or U42558 (N_42558,N_42171,N_42491);
nor U42559 (N_42559,N_42457,N_42492);
nor U42560 (N_42560,N_42255,N_42481);
xnor U42561 (N_42561,N_42262,N_42398);
xnor U42562 (N_42562,N_42317,N_42244);
and U42563 (N_42563,N_42469,N_42319);
nand U42564 (N_42564,N_42249,N_42185);
xnor U42565 (N_42565,N_42455,N_42235);
or U42566 (N_42566,N_42449,N_42225);
nand U42567 (N_42567,N_42250,N_42022);
nor U42568 (N_42568,N_42452,N_42091);
or U42569 (N_42569,N_42289,N_42296);
nor U42570 (N_42570,N_42316,N_42158);
and U42571 (N_42571,N_42047,N_42167);
xnor U42572 (N_42572,N_42059,N_42189);
nand U42573 (N_42573,N_42216,N_42028);
nor U42574 (N_42574,N_42389,N_42159);
nand U42575 (N_42575,N_42136,N_42463);
and U42576 (N_42576,N_42078,N_42166);
or U42577 (N_42577,N_42450,N_42335);
or U42578 (N_42578,N_42318,N_42019);
xnor U42579 (N_42579,N_42035,N_42081);
nor U42580 (N_42580,N_42294,N_42430);
nand U42581 (N_42581,N_42054,N_42170);
or U42582 (N_42582,N_42340,N_42380);
xnor U42583 (N_42583,N_42496,N_42211);
nand U42584 (N_42584,N_42199,N_42108);
or U42585 (N_42585,N_42362,N_42456);
or U42586 (N_42586,N_42461,N_42245);
xor U42587 (N_42587,N_42407,N_42152);
nor U42588 (N_42588,N_42111,N_42495);
nand U42589 (N_42589,N_42467,N_42365);
nand U42590 (N_42590,N_42223,N_42472);
xor U42591 (N_42591,N_42126,N_42098);
or U42592 (N_42592,N_42096,N_42196);
and U42593 (N_42593,N_42021,N_42395);
and U42594 (N_42594,N_42478,N_42313);
nand U42595 (N_42595,N_42110,N_42150);
nand U42596 (N_42596,N_42157,N_42116);
or U42597 (N_42597,N_42269,N_42310);
and U42598 (N_42598,N_42003,N_42322);
or U42599 (N_42599,N_42099,N_42036);
nor U42600 (N_42600,N_42181,N_42207);
or U42601 (N_42601,N_42400,N_42014);
nor U42602 (N_42602,N_42339,N_42288);
and U42603 (N_42603,N_42485,N_42070);
and U42604 (N_42604,N_42131,N_42448);
nand U42605 (N_42605,N_42497,N_42376);
nor U42606 (N_42606,N_42153,N_42214);
or U42607 (N_42607,N_42044,N_42302);
nand U42608 (N_42608,N_42348,N_42125);
nand U42609 (N_42609,N_42210,N_42402);
nor U42610 (N_42610,N_42272,N_42353);
or U42611 (N_42611,N_42174,N_42071);
or U42612 (N_42612,N_42050,N_42275);
and U42613 (N_42613,N_42490,N_42086);
or U42614 (N_42614,N_42038,N_42458);
nor U42615 (N_42615,N_42222,N_42109);
nand U42616 (N_42616,N_42419,N_42127);
or U42617 (N_42617,N_42464,N_42041);
or U42618 (N_42618,N_42325,N_42100);
xnor U42619 (N_42619,N_42355,N_42454);
nor U42620 (N_42620,N_42239,N_42482);
xor U42621 (N_42621,N_42349,N_42314);
or U42622 (N_42622,N_42040,N_42331);
or U42623 (N_42623,N_42139,N_42352);
nand U42624 (N_42624,N_42228,N_42486);
nand U42625 (N_42625,N_42281,N_42058);
nor U42626 (N_42626,N_42137,N_42334);
nand U42627 (N_42627,N_42459,N_42421);
xnor U42628 (N_42628,N_42256,N_42084);
xor U42629 (N_42629,N_42447,N_42175);
nand U42630 (N_42630,N_42082,N_42438);
nand U42631 (N_42631,N_42203,N_42252);
and U42632 (N_42632,N_42422,N_42297);
and U42633 (N_42633,N_42043,N_42287);
xor U42634 (N_42634,N_42394,N_42333);
xor U42635 (N_42635,N_42149,N_42446);
and U42636 (N_42636,N_42409,N_42290);
nor U42637 (N_42637,N_42328,N_42064);
nand U42638 (N_42638,N_42130,N_42308);
nor U42639 (N_42639,N_42006,N_42083);
nand U42640 (N_42640,N_42011,N_42092);
nand U42641 (N_42641,N_42301,N_42133);
nor U42642 (N_42642,N_42418,N_42435);
nand U42643 (N_42643,N_42344,N_42471);
or U42644 (N_42644,N_42345,N_42439);
xnor U42645 (N_42645,N_42012,N_42385);
nand U42646 (N_42646,N_42120,N_42423);
or U42647 (N_42647,N_42414,N_42390);
xor U42648 (N_42648,N_42300,N_42201);
or U42649 (N_42649,N_42178,N_42055);
and U42650 (N_42650,N_42180,N_42221);
nor U42651 (N_42651,N_42140,N_42072);
xnor U42652 (N_42652,N_42208,N_42154);
or U42653 (N_42653,N_42263,N_42442);
or U42654 (N_42654,N_42232,N_42212);
or U42655 (N_42655,N_42336,N_42155);
or U42656 (N_42656,N_42498,N_42046);
and U42657 (N_42657,N_42261,N_42373);
and U42658 (N_42658,N_42220,N_42129);
or U42659 (N_42659,N_42324,N_42388);
xnor U42660 (N_42660,N_42128,N_42284);
nand U42661 (N_42661,N_42283,N_42309);
and U42662 (N_42662,N_42259,N_42246);
xor U42663 (N_42663,N_42307,N_42097);
xnor U42664 (N_42664,N_42441,N_42254);
xor U42665 (N_42665,N_42278,N_42257);
or U42666 (N_42666,N_42364,N_42434);
nand U42667 (N_42667,N_42465,N_42264);
xnor U42668 (N_42668,N_42104,N_42017);
nor U42669 (N_42669,N_42379,N_42360);
or U42670 (N_42670,N_42384,N_42391);
nand U42671 (N_42671,N_42293,N_42295);
nand U42672 (N_42672,N_42176,N_42124);
and U42673 (N_42673,N_42102,N_42007);
or U42674 (N_42674,N_42417,N_42277);
and U42675 (N_42675,N_42424,N_42470);
nand U42676 (N_42676,N_42489,N_42393);
and U42677 (N_42677,N_42342,N_42443);
and U42678 (N_42678,N_42226,N_42066);
or U42679 (N_42679,N_42023,N_42020);
and U42680 (N_42680,N_42206,N_42063);
or U42681 (N_42681,N_42484,N_42406);
nand U42682 (N_42682,N_42444,N_42240);
and U42683 (N_42683,N_42305,N_42144);
nand U42684 (N_42684,N_42009,N_42381);
nand U42685 (N_42685,N_42366,N_42477);
or U42686 (N_42686,N_42359,N_42052);
nor U42687 (N_42687,N_42291,N_42087);
nor U42688 (N_42688,N_42230,N_42090);
and U42689 (N_42689,N_42138,N_42476);
or U42690 (N_42690,N_42285,N_42034);
and U42691 (N_42691,N_42303,N_42117);
and U42692 (N_42692,N_42089,N_42383);
and U42693 (N_42693,N_42361,N_42488);
xor U42694 (N_42694,N_42274,N_42231);
or U42695 (N_42695,N_42321,N_42412);
nor U42696 (N_42696,N_42161,N_42198);
or U42697 (N_42697,N_42341,N_42466);
and U42698 (N_42698,N_42143,N_42113);
nand U42699 (N_42699,N_42408,N_42480);
xnor U42700 (N_42700,N_42315,N_42415);
and U42701 (N_42701,N_42242,N_42032);
or U42702 (N_42702,N_42358,N_42142);
xnor U42703 (N_42703,N_42141,N_42347);
nand U42704 (N_42704,N_42343,N_42234);
or U42705 (N_42705,N_42280,N_42179);
and U42706 (N_42706,N_42122,N_42299);
nand U42707 (N_42707,N_42350,N_42473);
or U42708 (N_42708,N_42112,N_42168);
nor U42709 (N_42709,N_42427,N_42069);
nand U42710 (N_42710,N_42229,N_42487);
xor U42711 (N_42711,N_42499,N_42169);
nor U42712 (N_42712,N_42378,N_42243);
xor U42713 (N_42713,N_42182,N_42332);
nand U42714 (N_42714,N_42042,N_42165);
xnor U42715 (N_42715,N_42468,N_42073);
xnor U42716 (N_42716,N_42085,N_42025);
and U42717 (N_42717,N_42375,N_42194);
or U42718 (N_42718,N_42354,N_42209);
xor U42719 (N_42719,N_42016,N_42202);
nand U42720 (N_42720,N_42237,N_42453);
xnor U42721 (N_42721,N_42392,N_42095);
nor U42722 (N_42722,N_42224,N_42001);
xor U42723 (N_42723,N_42369,N_42371);
and U42724 (N_42724,N_42363,N_42401);
and U42725 (N_42725,N_42247,N_42134);
xnor U42726 (N_42726,N_42197,N_42329);
nor U42727 (N_42727,N_42462,N_42403);
or U42728 (N_42728,N_42233,N_42145);
xnor U42729 (N_42729,N_42292,N_42420);
nor U42730 (N_42730,N_42132,N_42049);
nand U42731 (N_42731,N_42436,N_42123);
or U42732 (N_42732,N_42183,N_42105);
or U42733 (N_42733,N_42107,N_42416);
nor U42734 (N_42734,N_42074,N_42200);
xnor U42735 (N_42735,N_42440,N_42213);
or U42736 (N_42736,N_42067,N_42382);
xnor U42737 (N_42737,N_42218,N_42057);
or U42738 (N_42738,N_42103,N_42010);
nand U42739 (N_42739,N_42433,N_42135);
and U42740 (N_42740,N_42377,N_42094);
nor U42741 (N_42741,N_42338,N_42065);
nand U42742 (N_42742,N_42248,N_42217);
or U42743 (N_42743,N_42026,N_42271);
xnor U42744 (N_42744,N_42101,N_42056);
xor U42745 (N_42745,N_42260,N_42164);
nand U42746 (N_42746,N_42037,N_42060);
nand U42747 (N_42747,N_42312,N_42410);
xor U42748 (N_42748,N_42075,N_42118);
or U42749 (N_42749,N_42282,N_42337);
nor U42750 (N_42750,N_42246,N_42097);
or U42751 (N_42751,N_42298,N_42054);
and U42752 (N_42752,N_42039,N_42123);
or U42753 (N_42753,N_42295,N_42363);
nor U42754 (N_42754,N_42447,N_42232);
and U42755 (N_42755,N_42273,N_42432);
nor U42756 (N_42756,N_42407,N_42424);
or U42757 (N_42757,N_42448,N_42165);
nor U42758 (N_42758,N_42042,N_42431);
nand U42759 (N_42759,N_42497,N_42209);
nor U42760 (N_42760,N_42173,N_42006);
or U42761 (N_42761,N_42341,N_42101);
nand U42762 (N_42762,N_42252,N_42364);
or U42763 (N_42763,N_42326,N_42095);
xnor U42764 (N_42764,N_42475,N_42330);
xnor U42765 (N_42765,N_42126,N_42214);
nor U42766 (N_42766,N_42372,N_42460);
xnor U42767 (N_42767,N_42459,N_42371);
nor U42768 (N_42768,N_42318,N_42478);
or U42769 (N_42769,N_42124,N_42097);
nand U42770 (N_42770,N_42124,N_42467);
or U42771 (N_42771,N_42257,N_42403);
nor U42772 (N_42772,N_42309,N_42033);
xnor U42773 (N_42773,N_42046,N_42397);
xnor U42774 (N_42774,N_42109,N_42121);
xnor U42775 (N_42775,N_42288,N_42156);
or U42776 (N_42776,N_42348,N_42201);
and U42777 (N_42777,N_42087,N_42424);
nand U42778 (N_42778,N_42475,N_42470);
and U42779 (N_42779,N_42330,N_42123);
nor U42780 (N_42780,N_42351,N_42177);
nor U42781 (N_42781,N_42416,N_42315);
nor U42782 (N_42782,N_42279,N_42286);
and U42783 (N_42783,N_42328,N_42454);
xnor U42784 (N_42784,N_42137,N_42131);
xnor U42785 (N_42785,N_42022,N_42002);
xnor U42786 (N_42786,N_42194,N_42043);
or U42787 (N_42787,N_42455,N_42311);
xor U42788 (N_42788,N_42232,N_42193);
or U42789 (N_42789,N_42451,N_42046);
nor U42790 (N_42790,N_42202,N_42326);
and U42791 (N_42791,N_42140,N_42318);
and U42792 (N_42792,N_42318,N_42291);
xnor U42793 (N_42793,N_42392,N_42135);
nand U42794 (N_42794,N_42229,N_42417);
nand U42795 (N_42795,N_42223,N_42300);
nand U42796 (N_42796,N_42005,N_42457);
and U42797 (N_42797,N_42059,N_42474);
or U42798 (N_42798,N_42085,N_42158);
and U42799 (N_42799,N_42420,N_42370);
xnor U42800 (N_42800,N_42140,N_42317);
xor U42801 (N_42801,N_42489,N_42037);
nor U42802 (N_42802,N_42374,N_42244);
and U42803 (N_42803,N_42302,N_42154);
or U42804 (N_42804,N_42195,N_42121);
and U42805 (N_42805,N_42283,N_42347);
nand U42806 (N_42806,N_42031,N_42257);
nor U42807 (N_42807,N_42322,N_42295);
nor U42808 (N_42808,N_42352,N_42413);
nor U42809 (N_42809,N_42467,N_42324);
nor U42810 (N_42810,N_42336,N_42107);
nand U42811 (N_42811,N_42255,N_42320);
nand U42812 (N_42812,N_42358,N_42177);
nor U42813 (N_42813,N_42302,N_42174);
and U42814 (N_42814,N_42328,N_42447);
or U42815 (N_42815,N_42456,N_42214);
and U42816 (N_42816,N_42487,N_42422);
and U42817 (N_42817,N_42387,N_42205);
or U42818 (N_42818,N_42115,N_42236);
nand U42819 (N_42819,N_42481,N_42217);
nand U42820 (N_42820,N_42237,N_42382);
nand U42821 (N_42821,N_42220,N_42243);
or U42822 (N_42822,N_42196,N_42108);
or U42823 (N_42823,N_42190,N_42314);
xnor U42824 (N_42824,N_42047,N_42100);
or U42825 (N_42825,N_42368,N_42361);
xnor U42826 (N_42826,N_42244,N_42044);
nand U42827 (N_42827,N_42458,N_42048);
xnor U42828 (N_42828,N_42135,N_42387);
or U42829 (N_42829,N_42495,N_42181);
or U42830 (N_42830,N_42429,N_42055);
and U42831 (N_42831,N_42164,N_42177);
and U42832 (N_42832,N_42179,N_42246);
nor U42833 (N_42833,N_42438,N_42036);
and U42834 (N_42834,N_42496,N_42241);
nor U42835 (N_42835,N_42499,N_42313);
or U42836 (N_42836,N_42134,N_42266);
and U42837 (N_42837,N_42489,N_42168);
nor U42838 (N_42838,N_42088,N_42416);
or U42839 (N_42839,N_42307,N_42323);
and U42840 (N_42840,N_42194,N_42462);
nand U42841 (N_42841,N_42328,N_42489);
or U42842 (N_42842,N_42367,N_42403);
nor U42843 (N_42843,N_42275,N_42323);
nand U42844 (N_42844,N_42450,N_42320);
nor U42845 (N_42845,N_42346,N_42318);
or U42846 (N_42846,N_42214,N_42131);
nor U42847 (N_42847,N_42067,N_42372);
nand U42848 (N_42848,N_42107,N_42344);
xor U42849 (N_42849,N_42390,N_42307);
nand U42850 (N_42850,N_42061,N_42013);
nand U42851 (N_42851,N_42256,N_42487);
nand U42852 (N_42852,N_42072,N_42161);
or U42853 (N_42853,N_42173,N_42279);
and U42854 (N_42854,N_42139,N_42149);
nor U42855 (N_42855,N_42345,N_42348);
xnor U42856 (N_42856,N_42499,N_42368);
or U42857 (N_42857,N_42187,N_42186);
or U42858 (N_42858,N_42296,N_42037);
nand U42859 (N_42859,N_42216,N_42323);
and U42860 (N_42860,N_42205,N_42227);
or U42861 (N_42861,N_42399,N_42452);
nand U42862 (N_42862,N_42094,N_42206);
nor U42863 (N_42863,N_42297,N_42333);
nand U42864 (N_42864,N_42079,N_42012);
nand U42865 (N_42865,N_42325,N_42011);
nor U42866 (N_42866,N_42007,N_42447);
nor U42867 (N_42867,N_42008,N_42249);
nand U42868 (N_42868,N_42012,N_42227);
and U42869 (N_42869,N_42469,N_42168);
and U42870 (N_42870,N_42171,N_42351);
nand U42871 (N_42871,N_42069,N_42475);
nor U42872 (N_42872,N_42142,N_42317);
xnor U42873 (N_42873,N_42162,N_42052);
nor U42874 (N_42874,N_42027,N_42447);
nand U42875 (N_42875,N_42338,N_42231);
or U42876 (N_42876,N_42025,N_42280);
or U42877 (N_42877,N_42267,N_42476);
and U42878 (N_42878,N_42428,N_42415);
xor U42879 (N_42879,N_42013,N_42288);
nand U42880 (N_42880,N_42442,N_42381);
nand U42881 (N_42881,N_42364,N_42054);
nand U42882 (N_42882,N_42484,N_42474);
and U42883 (N_42883,N_42027,N_42043);
or U42884 (N_42884,N_42075,N_42161);
nor U42885 (N_42885,N_42207,N_42424);
xnor U42886 (N_42886,N_42367,N_42398);
xor U42887 (N_42887,N_42174,N_42486);
or U42888 (N_42888,N_42105,N_42034);
nand U42889 (N_42889,N_42248,N_42427);
xor U42890 (N_42890,N_42137,N_42301);
nand U42891 (N_42891,N_42236,N_42230);
nand U42892 (N_42892,N_42437,N_42290);
xor U42893 (N_42893,N_42275,N_42322);
xor U42894 (N_42894,N_42318,N_42217);
nor U42895 (N_42895,N_42464,N_42094);
nor U42896 (N_42896,N_42345,N_42138);
or U42897 (N_42897,N_42469,N_42121);
nor U42898 (N_42898,N_42458,N_42389);
nand U42899 (N_42899,N_42374,N_42349);
nor U42900 (N_42900,N_42177,N_42134);
or U42901 (N_42901,N_42024,N_42453);
xnor U42902 (N_42902,N_42255,N_42073);
or U42903 (N_42903,N_42024,N_42206);
xor U42904 (N_42904,N_42248,N_42176);
xnor U42905 (N_42905,N_42081,N_42042);
nand U42906 (N_42906,N_42291,N_42389);
or U42907 (N_42907,N_42030,N_42454);
nand U42908 (N_42908,N_42069,N_42259);
and U42909 (N_42909,N_42483,N_42432);
xor U42910 (N_42910,N_42272,N_42075);
nand U42911 (N_42911,N_42150,N_42139);
or U42912 (N_42912,N_42269,N_42330);
and U42913 (N_42913,N_42135,N_42037);
xnor U42914 (N_42914,N_42087,N_42308);
and U42915 (N_42915,N_42268,N_42289);
or U42916 (N_42916,N_42314,N_42495);
and U42917 (N_42917,N_42227,N_42377);
and U42918 (N_42918,N_42420,N_42269);
and U42919 (N_42919,N_42286,N_42141);
nor U42920 (N_42920,N_42499,N_42179);
or U42921 (N_42921,N_42471,N_42450);
and U42922 (N_42922,N_42461,N_42411);
and U42923 (N_42923,N_42202,N_42376);
or U42924 (N_42924,N_42214,N_42475);
and U42925 (N_42925,N_42049,N_42321);
and U42926 (N_42926,N_42238,N_42297);
and U42927 (N_42927,N_42279,N_42040);
and U42928 (N_42928,N_42236,N_42005);
or U42929 (N_42929,N_42495,N_42003);
and U42930 (N_42930,N_42227,N_42371);
nor U42931 (N_42931,N_42153,N_42377);
xor U42932 (N_42932,N_42166,N_42169);
nand U42933 (N_42933,N_42438,N_42475);
nor U42934 (N_42934,N_42185,N_42027);
xnor U42935 (N_42935,N_42234,N_42339);
or U42936 (N_42936,N_42478,N_42048);
or U42937 (N_42937,N_42474,N_42128);
and U42938 (N_42938,N_42305,N_42497);
or U42939 (N_42939,N_42319,N_42295);
or U42940 (N_42940,N_42045,N_42393);
nor U42941 (N_42941,N_42281,N_42248);
nand U42942 (N_42942,N_42439,N_42476);
nor U42943 (N_42943,N_42261,N_42429);
or U42944 (N_42944,N_42039,N_42251);
nor U42945 (N_42945,N_42389,N_42358);
or U42946 (N_42946,N_42481,N_42473);
and U42947 (N_42947,N_42079,N_42454);
nand U42948 (N_42948,N_42499,N_42004);
nor U42949 (N_42949,N_42327,N_42057);
nor U42950 (N_42950,N_42163,N_42132);
or U42951 (N_42951,N_42177,N_42303);
nor U42952 (N_42952,N_42303,N_42124);
nand U42953 (N_42953,N_42301,N_42259);
xnor U42954 (N_42954,N_42429,N_42023);
or U42955 (N_42955,N_42141,N_42358);
nand U42956 (N_42956,N_42490,N_42242);
xor U42957 (N_42957,N_42093,N_42396);
nand U42958 (N_42958,N_42477,N_42423);
xnor U42959 (N_42959,N_42424,N_42093);
nor U42960 (N_42960,N_42478,N_42480);
nor U42961 (N_42961,N_42133,N_42434);
or U42962 (N_42962,N_42246,N_42015);
xor U42963 (N_42963,N_42134,N_42425);
and U42964 (N_42964,N_42241,N_42464);
nor U42965 (N_42965,N_42057,N_42434);
nand U42966 (N_42966,N_42478,N_42153);
nor U42967 (N_42967,N_42231,N_42495);
and U42968 (N_42968,N_42238,N_42439);
and U42969 (N_42969,N_42128,N_42134);
nand U42970 (N_42970,N_42375,N_42431);
and U42971 (N_42971,N_42323,N_42249);
xnor U42972 (N_42972,N_42450,N_42270);
or U42973 (N_42973,N_42095,N_42231);
or U42974 (N_42974,N_42252,N_42432);
xnor U42975 (N_42975,N_42226,N_42035);
nand U42976 (N_42976,N_42369,N_42012);
and U42977 (N_42977,N_42216,N_42432);
nor U42978 (N_42978,N_42489,N_42242);
or U42979 (N_42979,N_42004,N_42337);
or U42980 (N_42980,N_42082,N_42475);
nand U42981 (N_42981,N_42328,N_42371);
xnor U42982 (N_42982,N_42201,N_42301);
or U42983 (N_42983,N_42442,N_42131);
nand U42984 (N_42984,N_42151,N_42109);
nor U42985 (N_42985,N_42001,N_42195);
nor U42986 (N_42986,N_42007,N_42266);
and U42987 (N_42987,N_42370,N_42162);
nand U42988 (N_42988,N_42014,N_42182);
or U42989 (N_42989,N_42130,N_42387);
xnor U42990 (N_42990,N_42436,N_42131);
nor U42991 (N_42991,N_42353,N_42202);
nor U42992 (N_42992,N_42381,N_42057);
and U42993 (N_42993,N_42093,N_42060);
xnor U42994 (N_42994,N_42314,N_42042);
nand U42995 (N_42995,N_42214,N_42300);
nor U42996 (N_42996,N_42152,N_42352);
xor U42997 (N_42997,N_42008,N_42061);
or U42998 (N_42998,N_42223,N_42438);
nand U42999 (N_42999,N_42111,N_42359);
or U43000 (N_43000,N_42978,N_42609);
and U43001 (N_43001,N_42667,N_42975);
nor U43002 (N_43002,N_42962,N_42508);
nor U43003 (N_43003,N_42695,N_42993);
nor U43004 (N_43004,N_42929,N_42703);
or U43005 (N_43005,N_42640,N_42729);
and U43006 (N_43006,N_42678,N_42600);
nor U43007 (N_43007,N_42854,N_42803);
and U43008 (N_43008,N_42802,N_42608);
and U43009 (N_43009,N_42817,N_42941);
or U43010 (N_43010,N_42659,N_42859);
or U43011 (N_43011,N_42568,N_42708);
nor U43012 (N_43012,N_42663,N_42737);
xor U43013 (N_43013,N_42931,N_42951);
nor U43014 (N_43014,N_42810,N_42945);
nand U43015 (N_43015,N_42831,N_42572);
nand U43016 (N_43016,N_42840,N_42629);
nor U43017 (N_43017,N_42584,N_42687);
and U43018 (N_43018,N_42519,N_42949);
or U43019 (N_43019,N_42719,N_42655);
xor U43020 (N_43020,N_42551,N_42815);
and U43021 (N_43021,N_42633,N_42755);
or U43022 (N_43022,N_42943,N_42807);
nand U43023 (N_43023,N_42959,N_42707);
or U43024 (N_43024,N_42699,N_42919);
nor U43025 (N_43025,N_42739,N_42862);
nor U43026 (N_43026,N_42961,N_42611);
or U43027 (N_43027,N_42642,N_42774);
nor U43028 (N_43028,N_42883,N_42786);
xnor U43029 (N_43029,N_42821,N_42999);
or U43030 (N_43030,N_42776,N_42620);
nor U43031 (N_43031,N_42882,N_42857);
xor U43032 (N_43032,N_42670,N_42845);
or U43033 (N_43033,N_42747,N_42886);
nor U43034 (N_43034,N_42903,N_42805);
nand U43035 (N_43035,N_42897,N_42875);
nand U43036 (N_43036,N_42734,N_42916);
or U43037 (N_43037,N_42935,N_42933);
or U43038 (N_43038,N_42520,N_42760);
or U43039 (N_43039,N_42689,N_42824);
and U43040 (N_43040,N_42826,N_42592);
nor U43041 (N_43041,N_42740,N_42991);
and U43042 (N_43042,N_42795,N_42730);
and U43043 (N_43043,N_42523,N_42578);
and U43044 (N_43044,N_42535,N_42717);
xnor U43045 (N_43045,N_42938,N_42696);
or U43046 (N_43046,N_42868,N_42727);
xor U43047 (N_43047,N_42843,N_42563);
nand U43048 (N_43048,N_42521,N_42722);
or U43049 (N_43049,N_42529,N_42564);
nand U43050 (N_43050,N_42861,N_42559);
and U43051 (N_43051,N_42829,N_42796);
or U43052 (N_43052,N_42507,N_42928);
or U43053 (N_43053,N_42567,N_42997);
or U43054 (N_43054,N_42579,N_42725);
and U43055 (N_43055,N_42517,N_42968);
or U43056 (N_43056,N_42524,N_42974);
and U43057 (N_43057,N_42501,N_42867);
nor U43058 (N_43058,N_42809,N_42621);
and U43059 (N_43059,N_42674,N_42615);
nand U43060 (N_43060,N_42606,N_42542);
nand U43061 (N_43061,N_42808,N_42917);
nor U43062 (N_43062,N_42622,N_42522);
and U43063 (N_43063,N_42632,N_42716);
nor U43064 (N_43064,N_42847,N_42896);
nor U43065 (N_43065,N_42823,N_42749);
nor U43066 (N_43066,N_42661,N_42753);
nand U43067 (N_43067,N_42791,N_42799);
xor U43068 (N_43068,N_42971,N_42890);
xor U43069 (N_43069,N_42595,N_42530);
and U43070 (N_43070,N_42713,N_42969);
nand U43071 (N_43071,N_42976,N_42569);
xnor U43072 (N_43072,N_42770,N_42988);
nor U43073 (N_43073,N_42972,N_42733);
xor U43074 (N_43074,N_42736,N_42677);
nor U43075 (N_43075,N_42798,N_42647);
nor U43076 (N_43076,N_42757,N_42652);
nor U43077 (N_43077,N_42554,N_42947);
nor U43078 (N_43078,N_42830,N_42833);
nand U43079 (N_43079,N_42514,N_42926);
or U43080 (N_43080,N_42819,N_42536);
nand U43081 (N_43081,N_42697,N_42921);
xor U43082 (N_43082,N_42956,N_42671);
xor U43083 (N_43083,N_42894,N_42626);
and U43084 (N_43084,N_42700,N_42992);
nor U43085 (N_43085,N_42793,N_42714);
xor U43086 (N_43086,N_42533,N_42984);
nand U43087 (N_43087,N_42724,N_42765);
and U43088 (N_43088,N_42915,N_42658);
nand U43089 (N_43089,N_42906,N_42601);
and U43090 (N_43090,N_42756,N_42726);
or U43091 (N_43091,N_42966,N_42851);
and U43092 (N_43092,N_42635,N_42591);
or U43093 (N_43093,N_42630,N_42813);
nand U43094 (N_43094,N_42675,N_42781);
xor U43095 (N_43095,N_42923,N_42534);
nand U43096 (N_43096,N_42679,N_42594);
nor U43097 (N_43097,N_42922,N_42586);
or U43098 (N_43098,N_42780,N_42925);
or U43099 (N_43099,N_42684,N_42761);
nand U43100 (N_43100,N_42650,N_42806);
nand U43101 (N_43101,N_42599,N_42500);
or U43102 (N_43102,N_42914,N_42668);
and U43103 (N_43103,N_42553,N_42986);
nor U43104 (N_43104,N_42548,N_42930);
nor U43105 (N_43105,N_42979,N_42628);
xnor U43106 (N_43106,N_42881,N_42814);
nand U43107 (N_43107,N_42698,N_42528);
and U43108 (N_43108,N_42918,N_42602);
nand U43109 (N_43109,N_42623,N_42904);
xnor U43110 (N_43110,N_42526,N_42811);
nand U43111 (N_43111,N_42583,N_42792);
nand U43112 (N_43112,N_42646,N_42638);
nor U43113 (N_43113,N_42898,N_42634);
nand U43114 (N_43114,N_42872,N_42587);
nor U43115 (N_43115,N_42664,N_42718);
and U43116 (N_43116,N_42871,N_42607);
or U43117 (N_43117,N_42510,N_42772);
xor U43118 (N_43118,N_42768,N_42955);
or U43119 (N_43119,N_42527,N_42525);
and U43120 (N_43120,N_42574,N_42552);
nand U43121 (N_43121,N_42758,N_42750);
or U43122 (N_43122,N_42751,N_42538);
nand U43123 (N_43123,N_42785,N_42545);
and U43124 (N_43124,N_42920,N_42989);
nor U43125 (N_43125,N_42560,N_42651);
or U43126 (N_43126,N_42889,N_42649);
and U43127 (N_43127,N_42644,N_42627);
nor U43128 (N_43128,N_42596,N_42790);
or U43129 (N_43129,N_42812,N_42543);
or U43130 (N_43130,N_42878,N_42777);
xor U43131 (N_43131,N_42709,N_42769);
and U43132 (N_43132,N_42963,N_42953);
nor U43133 (N_43133,N_42597,N_42575);
or U43134 (N_43134,N_42539,N_42705);
nor U43135 (N_43135,N_42994,N_42616);
and U43136 (N_43136,N_42998,N_42869);
and U43137 (N_43137,N_42879,N_42827);
and U43138 (N_43138,N_42852,N_42762);
or U43139 (N_43139,N_42641,N_42673);
xnor U43140 (N_43140,N_42832,N_42745);
xor U43141 (N_43141,N_42907,N_42771);
nand U43142 (N_43142,N_42549,N_42842);
xor U43143 (N_43143,N_42556,N_42888);
or U43144 (N_43144,N_42764,N_42816);
nor U43145 (N_43145,N_42980,N_42853);
and U43146 (N_43146,N_42789,N_42746);
and U43147 (N_43147,N_42558,N_42656);
xor U43148 (N_43148,N_42688,N_42728);
or U43149 (N_43149,N_42910,N_42504);
and U43150 (N_43150,N_42932,N_42721);
nand U43151 (N_43151,N_42794,N_42619);
or U43152 (N_43152,N_42912,N_42565);
nor U43153 (N_43153,N_42748,N_42895);
xnor U43154 (N_43154,N_42893,N_42874);
nand U43155 (N_43155,N_42909,N_42715);
xor U43156 (N_43156,N_42518,N_42835);
nor U43157 (N_43157,N_42509,N_42577);
nand U43158 (N_43158,N_42787,N_42754);
and U43159 (N_43159,N_42511,N_42547);
nor U43160 (N_43160,N_42686,N_42503);
or U43161 (N_43161,N_42983,N_42982);
xnor U43162 (N_43162,N_42855,N_42701);
and U43163 (N_43163,N_42981,N_42576);
nand U43164 (N_43164,N_42990,N_42515);
nor U43165 (N_43165,N_42561,N_42741);
xor U43166 (N_43166,N_42838,N_42804);
xor U43167 (N_43167,N_42582,N_42850);
and U43168 (N_43168,N_42939,N_42537);
xor U43169 (N_43169,N_42544,N_42512);
and U43170 (N_43170,N_42797,N_42704);
nand U43171 (N_43171,N_42566,N_42513);
xor U43172 (N_43172,N_42706,N_42901);
or U43173 (N_43173,N_42657,N_42618);
and U43174 (N_43174,N_42766,N_42885);
xnor U43175 (N_43175,N_42767,N_42987);
and U43176 (N_43176,N_42887,N_42944);
and U43177 (N_43177,N_42660,N_42864);
nand U43178 (N_43178,N_42877,N_42532);
and U43179 (N_43179,N_42702,N_42555);
nand U43180 (N_43180,N_42763,N_42589);
xnor U43181 (N_43181,N_42645,N_42977);
or U43182 (N_43182,N_42680,N_42849);
and U43183 (N_43183,N_42884,N_42665);
or U43184 (N_43184,N_42800,N_42957);
nor U43185 (N_43185,N_42581,N_42822);
nand U43186 (N_43186,N_42669,N_42752);
and U43187 (N_43187,N_42940,N_42643);
nor U43188 (N_43188,N_42676,N_42580);
xnor U43189 (N_43189,N_42783,N_42735);
or U43190 (N_43190,N_42778,N_42996);
xnor U43191 (N_43191,N_42846,N_42967);
or U43192 (N_43192,N_42856,N_42900);
and U43193 (N_43193,N_42905,N_42891);
and U43194 (N_43194,N_42653,N_42631);
xnor U43195 (N_43195,N_42531,N_42557);
and U43196 (N_43196,N_42876,N_42694);
nand U43197 (N_43197,N_42573,N_42712);
nand U43198 (N_43198,N_42637,N_42541);
and U43199 (N_43199,N_42958,N_42720);
or U43200 (N_43200,N_42870,N_42866);
and U43201 (N_43201,N_42731,N_42784);
and U43202 (N_43202,N_42950,N_42865);
and U43203 (N_43203,N_42711,N_42672);
nor U43204 (N_43204,N_42742,N_42710);
nor U43205 (N_43205,N_42934,N_42965);
and U43206 (N_43206,N_42863,N_42562);
and U43207 (N_43207,N_42505,N_42683);
xnor U43208 (N_43208,N_42942,N_42848);
or U43209 (N_43209,N_42964,N_42828);
and U43210 (N_43210,N_42902,N_42612);
xnor U43211 (N_43211,N_42662,N_42502);
or U43212 (N_43212,N_42546,N_42570);
xor U43213 (N_43213,N_42985,N_42839);
and U43214 (N_43214,N_42639,N_42648);
nand U43215 (N_43215,N_42506,N_42681);
nor U43216 (N_43216,N_42995,N_42801);
or U43217 (N_43217,N_42952,N_42820);
nand U43218 (N_43218,N_42625,N_42841);
and U43219 (N_43219,N_42604,N_42614);
nor U43220 (N_43220,N_42908,N_42936);
and U43221 (N_43221,N_42899,N_42693);
nand U43222 (N_43222,N_42892,N_42744);
nand U43223 (N_43223,N_42973,N_42682);
or U43224 (N_43224,N_42690,N_42743);
nor U43225 (N_43225,N_42588,N_42516);
nand U43226 (N_43226,N_42818,N_42773);
xor U43227 (N_43227,N_42685,N_42666);
xnor U43228 (N_43228,N_42691,N_42924);
or U43229 (N_43229,N_42825,N_42540);
xnor U43230 (N_43230,N_42550,N_42927);
and U43231 (N_43231,N_42585,N_42617);
xor U43232 (N_43232,N_42911,N_42782);
or U43233 (N_43233,N_42723,N_42970);
or U43234 (N_43234,N_42738,N_42590);
nand U43235 (N_43235,N_42960,N_42571);
xor U43236 (N_43236,N_42937,N_42913);
xnor U43237 (N_43237,N_42654,N_42880);
xnor U43238 (N_43238,N_42732,N_42788);
xnor U43239 (N_43239,N_42954,N_42605);
or U43240 (N_43240,N_42873,N_42759);
or U43241 (N_43241,N_42613,N_42844);
and U43242 (N_43242,N_42598,N_42603);
nor U43243 (N_43243,N_42858,N_42948);
or U43244 (N_43244,N_42692,N_42624);
nor U43245 (N_43245,N_42837,N_42860);
nor U43246 (N_43246,N_42946,N_42836);
or U43247 (N_43247,N_42636,N_42779);
or U43248 (N_43248,N_42593,N_42610);
or U43249 (N_43249,N_42834,N_42775);
and U43250 (N_43250,N_42880,N_42714);
xor U43251 (N_43251,N_42580,N_42864);
and U43252 (N_43252,N_42842,N_42938);
xor U43253 (N_43253,N_42913,N_42943);
nor U43254 (N_43254,N_42661,N_42994);
nor U43255 (N_43255,N_42553,N_42776);
nand U43256 (N_43256,N_42822,N_42558);
xor U43257 (N_43257,N_42571,N_42809);
nor U43258 (N_43258,N_42849,N_42971);
and U43259 (N_43259,N_42747,N_42647);
xnor U43260 (N_43260,N_42556,N_42608);
and U43261 (N_43261,N_42579,N_42578);
xor U43262 (N_43262,N_42653,N_42796);
xor U43263 (N_43263,N_42537,N_42618);
xnor U43264 (N_43264,N_42544,N_42797);
nor U43265 (N_43265,N_42883,N_42523);
and U43266 (N_43266,N_42710,N_42928);
nand U43267 (N_43267,N_42798,N_42595);
xor U43268 (N_43268,N_42948,N_42754);
and U43269 (N_43269,N_42815,N_42722);
or U43270 (N_43270,N_42725,N_42974);
xnor U43271 (N_43271,N_42883,N_42876);
xnor U43272 (N_43272,N_42966,N_42598);
or U43273 (N_43273,N_42573,N_42974);
or U43274 (N_43274,N_42640,N_42906);
nand U43275 (N_43275,N_42824,N_42927);
nand U43276 (N_43276,N_42944,N_42963);
xor U43277 (N_43277,N_42782,N_42546);
nor U43278 (N_43278,N_42685,N_42965);
xor U43279 (N_43279,N_42755,N_42811);
and U43280 (N_43280,N_42796,N_42608);
xor U43281 (N_43281,N_42935,N_42768);
xor U43282 (N_43282,N_42835,N_42938);
xor U43283 (N_43283,N_42934,N_42819);
nand U43284 (N_43284,N_42996,N_42826);
nor U43285 (N_43285,N_42816,N_42901);
nor U43286 (N_43286,N_42581,N_42563);
nor U43287 (N_43287,N_42751,N_42879);
nand U43288 (N_43288,N_42596,N_42728);
or U43289 (N_43289,N_42984,N_42685);
nor U43290 (N_43290,N_42827,N_42698);
and U43291 (N_43291,N_42973,N_42610);
xor U43292 (N_43292,N_42946,N_42579);
xor U43293 (N_43293,N_42728,N_42833);
xnor U43294 (N_43294,N_42513,N_42720);
nor U43295 (N_43295,N_42951,N_42624);
and U43296 (N_43296,N_42535,N_42580);
xnor U43297 (N_43297,N_42986,N_42508);
or U43298 (N_43298,N_42579,N_42615);
or U43299 (N_43299,N_42802,N_42926);
nand U43300 (N_43300,N_42859,N_42982);
nand U43301 (N_43301,N_42842,N_42699);
nor U43302 (N_43302,N_42624,N_42709);
or U43303 (N_43303,N_42808,N_42703);
or U43304 (N_43304,N_42896,N_42825);
nor U43305 (N_43305,N_42868,N_42813);
or U43306 (N_43306,N_42719,N_42990);
nand U43307 (N_43307,N_42901,N_42521);
or U43308 (N_43308,N_42569,N_42549);
or U43309 (N_43309,N_42896,N_42586);
nor U43310 (N_43310,N_42694,N_42935);
nor U43311 (N_43311,N_42825,N_42549);
nand U43312 (N_43312,N_42801,N_42813);
xnor U43313 (N_43313,N_42534,N_42614);
nor U43314 (N_43314,N_42619,N_42578);
or U43315 (N_43315,N_42517,N_42613);
and U43316 (N_43316,N_42807,N_42855);
nand U43317 (N_43317,N_42532,N_42682);
and U43318 (N_43318,N_42631,N_42796);
xnor U43319 (N_43319,N_42595,N_42887);
nand U43320 (N_43320,N_42962,N_42553);
nor U43321 (N_43321,N_42546,N_42733);
or U43322 (N_43322,N_42899,N_42957);
or U43323 (N_43323,N_42774,N_42925);
and U43324 (N_43324,N_42948,N_42677);
nand U43325 (N_43325,N_42721,N_42854);
nor U43326 (N_43326,N_42558,N_42979);
nor U43327 (N_43327,N_42631,N_42608);
nand U43328 (N_43328,N_42545,N_42613);
and U43329 (N_43329,N_42706,N_42665);
or U43330 (N_43330,N_42585,N_42541);
or U43331 (N_43331,N_42844,N_42683);
xor U43332 (N_43332,N_42886,N_42770);
and U43333 (N_43333,N_42826,N_42924);
xnor U43334 (N_43334,N_42633,N_42685);
xor U43335 (N_43335,N_42553,N_42788);
nand U43336 (N_43336,N_42839,N_42910);
or U43337 (N_43337,N_42851,N_42771);
and U43338 (N_43338,N_42794,N_42901);
nand U43339 (N_43339,N_42854,N_42961);
nor U43340 (N_43340,N_42665,N_42604);
nand U43341 (N_43341,N_42848,N_42736);
and U43342 (N_43342,N_42661,N_42779);
nand U43343 (N_43343,N_42710,N_42646);
and U43344 (N_43344,N_42599,N_42630);
and U43345 (N_43345,N_42630,N_42728);
xor U43346 (N_43346,N_42967,N_42937);
and U43347 (N_43347,N_42710,N_42994);
nand U43348 (N_43348,N_42805,N_42813);
nor U43349 (N_43349,N_42671,N_42764);
nand U43350 (N_43350,N_42891,N_42881);
or U43351 (N_43351,N_42531,N_42682);
or U43352 (N_43352,N_42581,N_42865);
and U43353 (N_43353,N_42533,N_42837);
or U43354 (N_43354,N_42597,N_42800);
and U43355 (N_43355,N_42662,N_42530);
and U43356 (N_43356,N_42617,N_42666);
and U43357 (N_43357,N_42503,N_42630);
or U43358 (N_43358,N_42928,N_42916);
or U43359 (N_43359,N_42769,N_42555);
nor U43360 (N_43360,N_42844,N_42930);
and U43361 (N_43361,N_42554,N_42922);
and U43362 (N_43362,N_42602,N_42912);
xor U43363 (N_43363,N_42705,N_42513);
nand U43364 (N_43364,N_42852,N_42760);
xnor U43365 (N_43365,N_42520,N_42966);
and U43366 (N_43366,N_42512,N_42853);
or U43367 (N_43367,N_42740,N_42932);
nand U43368 (N_43368,N_42523,N_42823);
and U43369 (N_43369,N_42754,N_42758);
or U43370 (N_43370,N_42916,N_42925);
nor U43371 (N_43371,N_42584,N_42659);
and U43372 (N_43372,N_42691,N_42656);
xnor U43373 (N_43373,N_42786,N_42754);
or U43374 (N_43374,N_42938,N_42569);
or U43375 (N_43375,N_42736,N_42501);
or U43376 (N_43376,N_42758,N_42546);
nor U43377 (N_43377,N_42780,N_42764);
and U43378 (N_43378,N_42575,N_42734);
and U43379 (N_43379,N_42906,N_42600);
or U43380 (N_43380,N_42545,N_42970);
xnor U43381 (N_43381,N_42755,N_42821);
or U43382 (N_43382,N_42929,N_42576);
or U43383 (N_43383,N_42728,N_42846);
xnor U43384 (N_43384,N_42852,N_42954);
nand U43385 (N_43385,N_42864,N_42769);
nor U43386 (N_43386,N_42978,N_42965);
or U43387 (N_43387,N_42861,N_42893);
or U43388 (N_43388,N_42642,N_42707);
nand U43389 (N_43389,N_42712,N_42899);
and U43390 (N_43390,N_42503,N_42502);
or U43391 (N_43391,N_42823,N_42826);
or U43392 (N_43392,N_42801,N_42569);
nor U43393 (N_43393,N_42907,N_42879);
and U43394 (N_43394,N_42849,N_42695);
nand U43395 (N_43395,N_42527,N_42710);
nand U43396 (N_43396,N_42912,N_42995);
and U43397 (N_43397,N_42593,N_42547);
nand U43398 (N_43398,N_42728,N_42839);
nor U43399 (N_43399,N_42716,N_42642);
xnor U43400 (N_43400,N_42884,N_42821);
or U43401 (N_43401,N_42925,N_42579);
nand U43402 (N_43402,N_42598,N_42986);
or U43403 (N_43403,N_42650,N_42683);
xor U43404 (N_43404,N_42880,N_42607);
nand U43405 (N_43405,N_42596,N_42817);
nor U43406 (N_43406,N_42604,N_42631);
nor U43407 (N_43407,N_42888,N_42752);
nand U43408 (N_43408,N_42666,N_42814);
nor U43409 (N_43409,N_42724,N_42504);
xnor U43410 (N_43410,N_42917,N_42984);
nand U43411 (N_43411,N_42629,N_42697);
nand U43412 (N_43412,N_42828,N_42907);
nor U43413 (N_43413,N_42743,N_42598);
nor U43414 (N_43414,N_42848,N_42619);
xor U43415 (N_43415,N_42962,N_42904);
nand U43416 (N_43416,N_42680,N_42650);
xnor U43417 (N_43417,N_42919,N_42843);
nor U43418 (N_43418,N_42517,N_42698);
or U43419 (N_43419,N_42986,N_42966);
xor U43420 (N_43420,N_42565,N_42921);
nand U43421 (N_43421,N_42675,N_42509);
nor U43422 (N_43422,N_42734,N_42719);
or U43423 (N_43423,N_42633,N_42540);
nand U43424 (N_43424,N_42769,N_42868);
or U43425 (N_43425,N_42935,N_42750);
nand U43426 (N_43426,N_42959,N_42996);
nor U43427 (N_43427,N_42959,N_42863);
nor U43428 (N_43428,N_42844,N_42724);
or U43429 (N_43429,N_42829,N_42710);
and U43430 (N_43430,N_42917,N_42561);
xor U43431 (N_43431,N_42627,N_42641);
nand U43432 (N_43432,N_42942,N_42520);
or U43433 (N_43433,N_42717,N_42819);
or U43434 (N_43434,N_42782,N_42506);
xor U43435 (N_43435,N_42856,N_42812);
nand U43436 (N_43436,N_42830,N_42578);
xnor U43437 (N_43437,N_42979,N_42647);
and U43438 (N_43438,N_42729,N_42691);
nand U43439 (N_43439,N_42618,N_42561);
or U43440 (N_43440,N_42817,N_42615);
xor U43441 (N_43441,N_42600,N_42992);
or U43442 (N_43442,N_42574,N_42528);
nor U43443 (N_43443,N_42933,N_42765);
nor U43444 (N_43444,N_42648,N_42689);
and U43445 (N_43445,N_42667,N_42967);
xnor U43446 (N_43446,N_42546,N_42892);
or U43447 (N_43447,N_42625,N_42716);
nand U43448 (N_43448,N_42516,N_42714);
and U43449 (N_43449,N_42960,N_42910);
and U43450 (N_43450,N_42988,N_42696);
nand U43451 (N_43451,N_42677,N_42528);
nand U43452 (N_43452,N_42541,N_42678);
and U43453 (N_43453,N_42967,N_42958);
nor U43454 (N_43454,N_42848,N_42742);
or U43455 (N_43455,N_42874,N_42626);
nand U43456 (N_43456,N_42965,N_42794);
nor U43457 (N_43457,N_42744,N_42774);
nand U43458 (N_43458,N_42964,N_42946);
and U43459 (N_43459,N_42574,N_42687);
nor U43460 (N_43460,N_42867,N_42880);
nand U43461 (N_43461,N_42657,N_42687);
or U43462 (N_43462,N_42938,N_42931);
nand U43463 (N_43463,N_42889,N_42573);
or U43464 (N_43464,N_42804,N_42896);
xor U43465 (N_43465,N_42804,N_42666);
xor U43466 (N_43466,N_42726,N_42736);
xnor U43467 (N_43467,N_42778,N_42616);
nor U43468 (N_43468,N_42865,N_42757);
nand U43469 (N_43469,N_42636,N_42514);
nor U43470 (N_43470,N_42696,N_42898);
and U43471 (N_43471,N_42994,N_42507);
nor U43472 (N_43472,N_42977,N_42537);
xor U43473 (N_43473,N_42601,N_42839);
or U43474 (N_43474,N_42877,N_42808);
nand U43475 (N_43475,N_42653,N_42970);
xnor U43476 (N_43476,N_42542,N_42524);
and U43477 (N_43477,N_42940,N_42987);
xnor U43478 (N_43478,N_42807,N_42664);
and U43479 (N_43479,N_42770,N_42720);
or U43480 (N_43480,N_42753,N_42780);
and U43481 (N_43481,N_42584,N_42974);
nand U43482 (N_43482,N_42831,N_42624);
nand U43483 (N_43483,N_42766,N_42768);
nor U43484 (N_43484,N_42676,N_42779);
nand U43485 (N_43485,N_42666,N_42922);
xor U43486 (N_43486,N_42547,N_42839);
nor U43487 (N_43487,N_42947,N_42588);
and U43488 (N_43488,N_42766,N_42690);
nand U43489 (N_43489,N_42819,N_42666);
nor U43490 (N_43490,N_42920,N_42549);
or U43491 (N_43491,N_42538,N_42961);
or U43492 (N_43492,N_42745,N_42638);
xor U43493 (N_43493,N_42818,N_42861);
nor U43494 (N_43494,N_42653,N_42786);
or U43495 (N_43495,N_42666,N_42859);
and U43496 (N_43496,N_42987,N_42543);
or U43497 (N_43497,N_42795,N_42948);
and U43498 (N_43498,N_42895,N_42801);
nand U43499 (N_43499,N_42738,N_42972);
xor U43500 (N_43500,N_43091,N_43145);
and U43501 (N_43501,N_43395,N_43082);
nand U43502 (N_43502,N_43223,N_43457);
xor U43503 (N_43503,N_43024,N_43479);
xnor U43504 (N_43504,N_43261,N_43341);
and U43505 (N_43505,N_43268,N_43121);
nor U43506 (N_43506,N_43230,N_43054);
nand U43507 (N_43507,N_43345,N_43129);
and U43508 (N_43508,N_43052,N_43119);
nor U43509 (N_43509,N_43250,N_43017);
nand U43510 (N_43510,N_43254,N_43374);
xor U43511 (N_43511,N_43390,N_43138);
nand U43512 (N_43512,N_43367,N_43309);
nand U43513 (N_43513,N_43484,N_43072);
nor U43514 (N_43514,N_43216,N_43325);
or U43515 (N_43515,N_43346,N_43385);
nand U43516 (N_43516,N_43061,N_43260);
and U43517 (N_43517,N_43299,N_43146);
xor U43518 (N_43518,N_43469,N_43437);
xor U43519 (N_43519,N_43222,N_43173);
xnor U43520 (N_43520,N_43131,N_43047);
nor U43521 (N_43521,N_43422,N_43004);
or U43522 (N_43522,N_43231,N_43485);
and U43523 (N_43523,N_43062,N_43275);
or U43524 (N_43524,N_43156,N_43025);
nand U43525 (N_43525,N_43339,N_43132);
nand U43526 (N_43526,N_43413,N_43000);
nor U43527 (N_43527,N_43199,N_43241);
xor U43528 (N_43528,N_43314,N_43125);
xnor U43529 (N_43529,N_43462,N_43111);
or U43530 (N_43530,N_43371,N_43201);
and U43531 (N_43531,N_43320,N_43414);
nand U43532 (N_43532,N_43059,N_43391);
xor U43533 (N_43533,N_43240,N_43468);
and U43534 (N_43534,N_43203,N_43397);
and U43535 (N_43535,N_43116,N_43445);
and U43536 (N_43536,N_43482,N_43476);
nand U43537 (N_43537,N_43432,N_43381);
and U43538 (N_43538,N_43069,N_43166);
xor U43539 (N_43539,N_43327,N_43343);
nor U43540 (N_43540,N_43196,N_43194);
xnor U43541 (N_43541,N_43271,N_43489);
xnor U43542 (N_43542,N_43434,N_43493);
nand U43543 (N_43543,N_43488,N_43283);
nand U43544 (N_43544,N_43060,N_43234);
xor U43545 (N_43545,N_43093,N_43405);
xnor U43546 (N_43546,N_43195,N_43294);
nor U43547 (N_43547,N_43255,N_43155);
and U43548 (N_43548,N_43435,N_43092);
or U43549 (N_43549,N_43208,N_43356);
nand U43550 (N_43550,N_43454,N_43179);
nand U43551 (N_43551,N_43086,N_43105);
xnor U43552 (N_43552,N_43399,N_43313);
xor U43553 (N_43553,N_43012,N_43311);
and U43554 (N_43554,N_43494,N_43340);
or U43555 (N_43555,N_43338,N_43152);
nand U43556 (N_43556,N_43035,N_43363);
and U43557 (N_43557,N_43163,N_43274);
nor U43558 (N_43558,N_43321,N_43158);
xor U43559 (N_43559,N_43408,N_43384);
or U43560 (N_43560,N_43229,N_43227);
and U43561 (N_43561,N_43134,N_43070);
and U43562 (N_43562,N_43067,N_43026);
or U43563 (N_43563,N_43213,N_43358);
and U43564 (N_43564,N_43104,N_43188);
nor U43565 (N_43565,N_43492,N_43211);
xnor U43566 (N_43566,N_43330,N_43406);
and U43567 (N_43567,N_43467,N_43252);
nand U43568 (N_43568,N_43300,N_43370);
and U43569 (N_43569,N_43392,N_43162);
nor U43570 (N_43570,N_43065,N_43329);
nor U43571 (N_43571,N_43135,N_43427);
and U43572 (N_43572,N_43324,N_43192);
nand U43573 (N_43573,N_43307,N_43349);
and U43574 (N_43574,N_43386,N_43176);
xnor U43575 (N_43575,N_43142,N_43248);
and U43576 (N_43576,N_43396,N_43287);
nand U43577 (N_43577,N_43001,N_43027);
nand U43578 (N_43578,N_43455,N_43441);
nor U43579 (N_43579,N_43433,N_43029);
and U43580 (N_43580,N_43041,N_43398);
nand U43581 (N_43581,N_43184,N_43465);
nand U43582 (N_43582,N_43013,N_43015);
xnor U43583 (N_43583,N_43273,N_43483);
nand U43584 (N_43584,N_43318,N_43481);
nor U43585 (N_43585,N_43157,N_43154);
nor U43586 (N_43586,N_43471,N_43310);
nand U43587 (N_43587,N_43301,N_43197);
or U43588 (N_43588,N_43394,N_43127);
xnor U43589 (N_43589,N_43021,N_43113);
or U43590 (N_43590,N_43190,N_43045);
xnor U43591 (N_43591,N_43264,N_43030);
nor U43592 (N_43592,N_43217,N_43344);
or U43593 (N_43593,N_43186,N_43083);
nor U43594 (N_43594,N_43172,N_43251);
or U43595 (N_43595,N_43259,N_43456);
nand U43596 (N_43596,N_43218,N_43221);
nand U43597 (N_43597,N_43238,N_43031);
xor U43598 (N_43598,N_43315,N_43464);
and U43599 (N_43599,N_43044,N_43170);
nand U43600 (N_43600,N_43244,N_43232);
or U43601 (N_43601,N_43326,N_43486);
or U43602 (N_43602,N_43088,N_43480);
xnor U43603 (N_43603,N_43149,N_43191);
nor U43604 (N_43604,N_43245,N_43051);
nand U43605 (N_43605,N_43057,N_43016);
nor U43606 (N_43606,N_43110,N_43354);
nor U43607 (N_43607,N_43277,N_43351);
and U43608 (N_43608,N_43303,N_43499);
nand U43609 (N_43609,N_43348,N_43377);
and U43610 (N_43610,N_43498,N_43099);
and U43611 (N_43611,N_43302,N_43402);
or U43612 (N_43612,N_43079,N_43281);
or U43613 (N_43613,N_43153,N_43436);
and U43614 (N_43614,N_43247,N_43005);
and U43615 (N_43615,N_43382,N_43106);
nor U43616 (N_43616,N_43175,N_43228);
or U43617 (N_43617,N_43198,N_43298);
xor U43618 (N_43618,N_43018,N_43074);
and U43619 (N_43619,N_43447,N_43151);
and U43620 (N_43620,N_43084,N_43028);
nor U43621 (N_43621,N_43064,N_43076);
nor U43622 (N_43622,N_43056,N_43442);
or U43623 (N_43623,N_43187,N_43128);
nand U43624 (N_43624,N_43425,N_43270);
nor U43625 (N_43625,N_43478,N_43117);
nand U43626 (N_43626,N_43350,N_43058);
nor U43627 (N_43627,N_43081,N_43183);
nand U43628 (N_43628,N_43331,N_43265);
nand U43629 (N_43629,N_43055,N_43421);
nand U43630 (N_43630,N_43272,N_43235);
nor U43631 (N_43631,N_43256,N_43050);
or U43632 (N_43632,N_43066,N_43316);
xnor U43633 (N_43633,N_43169,N_43410);
nor U43634 (N_43634,N_43160,N_43010);
and U43635 (N_43635,N_43209,N_43077);
xnor U43636 (N_43636,N_43378,N_43267);
and U43637 (N_43637,N_43144,N_43034);
and U43638 (N_43638,N_43461,N_43164);
or U43639 (N_43639,N_43049,N_43008);
or U43640 (N_43640,N_43185,N_43114);
xor U43641 (N_43641,N_43141,N_43417);
nor U43642 (N_43642,N_43071,N_43204);
nor U43643 (N_43643,N_43328,N_43150);
nor U43644 (N_43644,N_43389,N_43475);
nor U43645 (N_43645,N_43249,N_43167);
or U43646 (N_43646,N_43007,N_43323);
xnor U43647 (N_43647,N_43096,N_43292);
nand U43648 (N_43648,N_43118,N_43237);
nor U43649 (N_43649,N_43403,N_43120);
and U43650 (N_43650,N_43379,N_43233);
xor U43651 (N_43651,N_43419,N_43446);
or U43652 (N_43652,N_43189,N_43112);
nand U43653 (N_43653,N_43383,N_43495);
xor U43654 (N_43654,N_43263,N_43450);
and U43655 (N_43655,N_43282,N_43243);
nor U43656 (N_43656,N_43449,N_43366);
xnor U43657 (N_43657,N_43246,N_43278);
xor U43658 (N_43658,N_43168,N_43124);
nand U43659 (N_43659,N_43451,N_43095);
or U43660 (N_43660,N_43126,N_43053);
nor U43661 (N_43661,N_43333,N_43337);
and U43662 (N_43662,N_43257,N_43137);
or U43663 (N_43663,N_43214,N_43317);
nor U43664 (N_43664,N_43215,N_43290);
and U43665 (N_43665,N_43411,N_43429);
and U43666 (N_43666,N_43087,N_43140);
nor U43667 (N_43667,N_43400,N_43133);
nor U43668 (N_43668,N_43409,N_43068);
nor U43669 (N_43669,N_43342,N_43103);
or U43670 (N_43670,N_43143,N_43332);
nor U43671 (N_43671,N_43048,N_43431);
nand U43672 (N_43672,N_43473,N_43098);
xnor U43673 (N_43673,N_43100,N_43297);
and U43674 (N_43674,N_43293,N_43401);
or U43675 (N_43675,N_43423,N_43239);
and U43676 (N_43676,N_43033,N_43448);
nor U43677 (N_43677,N_43123,N_43090);
nand U43678 (N_43678,N_43080,N_43219);
xnor U43679 (N_43679,N_43279,N_43296);
xor U43680 (N_43680,N_43205,N_43491);
or U43681 (N_43681,N_43075,N_43415);
xnor U43682 (N_43682,N_43412,N_43497);
nand U43683 (N_43683,N_43202,N_43352);
or U43684 (N_43684,N_43085,N_43380);
nand U43685 (N_43685,N_43078,N_43159);
nor U43686 (N_43686,N_43107,N_43336);
and U43687 (N_43687,N_43472,N_43207);
xnor U43688 (N_43688,N_43470,N_43477);
nand U43689 (N_43689,N_43073,N_43387);
nor U43690 (N_43690,N_43319,N_43101);
nand U43691 (N_43691,N_43286,N_43460);
and U43692 (N_43692,N_43291,N_43182);
or U43693 (N_43693,N_43474,N_43368);
or U43694 (N_43694,N_43014,N_43200);
or U43695 (N_43695,N_43020,N_43308);
nor U43696 (N_43696,N_43373,N_43011);
or U43697 (N_43697,N_43306,N_43006);
xor U43698 (N_43698,N_43042,N_43407);
and U43699 (N_43699,N_43426,N_43452);
and U43700 (N_43700,N_43335,N_43210);
nor U43701 (N_43701,N_43063,N_43416);
and U43702 (N_43702,N_43174,N_43404);
nor U43703 (N_43703,N_43220,N_43139);
or U43704 (N_43704,N_43388,N_43360);
and U43705 (N_43705,N_43347,N_43276);
nor U43706 (N_43706,N_43376,N_43459);
nor U43707 (N_43707,N_43487,N_43039);
nor U43708 (N_43708,N_43284,N_43369);
or U43709 (N_43709,N_43165,N_43364);
and U43710 (N_43710,N_43180,N_43453);
xnor U43711 (N_43711,N_43178,N_43463);
or U43712 (N_43712,N_43295,N_43148);
and U43713 (N_43713,N_43040,N_43102);
or U43714 (N_43714,N_43362,N_43253);
or U43715 (N_43715,N_43322,N_43258);
nand U43716 (N_43716,N_43440,N_43430);
xnor U43717 (N_43717,N_43365,N_43444);
nand U43718 (N_43718,N_43289,N_43266);
xor U43719 (N_43719,N_43375,N_43359);
and U43720 (N_43720,N_43458,N_43280);
nand U43721 (N_43721,N_43108,N_43089);
and U43722 (N_43722,N_43334,N_43372);
or U43723 (N_43723,N_43424,N_43003);
and U43724 (N_43724,N_43002,N_43269);
and U43725 (N_43725,N_43262,N_43353);
xnor U43726 (N_43726,N_43438,N_43181);
or U43727 (N_43727,N_43428,N_43357);
xor U43728 (N_43728,N_43036,N_43225);
or U43729 (N_43729,N_43206,N_43226);
or U43730 (N_43730,N_43193,N_43171);
and U43731 (N_43731,N_43023,N_43288);
xor U43732 (N_43732,N_43312,N_43236);
or U43733 (N_43733,N_43094,N_43224);
and U43734 (N_43734,N_43046,N_43161);
or U43735 (N_43735,N_43305,N_43009);
or U43736 (N_43736,N_43022,N_43285);
nand U43737 (N_43737,N_43466,N_43304);
nor U43738 (N_43738,N_43439,N_43038);
nand U43739 (N_43739,N_43361,N_43043);
nor U43740 (N_43740,N_43115,N_43242);
nor U43741 (N_43741,N_43147,N_43032);
or U43742 (N_43742,N_43177,N_43355);
or U43743 (N_43743,N_43496,N_43490);
or U43744 (N_43744,N_43418,N_43109);
nand U43745 (N_43745,N_43420,N_43393);
nor U43746 (N_43746,N_43130,N_43136);
nor U43747 (N_43747,N_43212,N_43122);
nor U43748 (N_43748,N_43037,N_43097);
or U43749 (N_43749,N_43019,N_43443);
and U43750 (N_43750,N_43141,N_43004);
nand U43751 (N_43751,N_43049,N_43052);
nor U43752 (N_43752,N_43044,N_43166);
and U43753 (N_43753,N_43351,N_43415);
or U43754 (N_43754,N_43240,N_43015);
or U43755 (N_43755,N_43014,N_43073);
xnor U43756 (N_43756,N_43070,N_43353);
nand U43757 (N_43757,N_43355,N_43175);
and U43758 (N_43758,N_43226,N_43176);
nor U43759 (N_43759,N_43435,N_43238);
nand U43760 (N_43760,N_43082,N_43246);
and U43761 (N_43761,N_43057,N_43302);
xor U43762 (N_43762,N_43406,N_43014);
nor U43763 (N_43763,N_43241,N_43364);
nand U43764 (N_43764,N_43124,N_43111);
xnor U43765 (N_43765,N_43158,N_43485);
nor U43766 (N_43766,N_43091,N_43065);
or U43767 (N_43767,N_43247,N_43357);
or U43768 (N_43768,N_43452,N_43359);
and U43769 (N_43769,N_43035,N_43247);
nand U43770 (N_43770,N_43306,N_43343);
and U43771 (N_43771,N_43472,N_43334);
and U43772 (N_43772,N_43367,N_43105);
and U43773 (N_43773,N_43465,N_43134);
nor U43774 (N_43774,N_43173,N_43241);
xnor U43775 (N_43775,N_43112,N_43163);
and U43776 (N_43776,N_43447,N_43233);
nand U43777 (N_43777,N_43489,N_43059);
and U43778 (N_43778,N_43343,N_43097);
nor U43779 (N_43779,N_43476,N_43227);
or U43780 (N_43780,N_43251,N_43237);
nor U43781 (N_43781,N_43087,N_43002);
nand U43782 (N_43782,N_43414,N_43161);
or U43783 (N_43783,N_43340,N_43462);
nand U43784 (N_43784,N_43063,N_43051);
and U43785 (N_43785,N_43069,N_43367);
or U43786 (N_43786,N_43299,N_43402);
or U43787 (N_43787,N_43003,N_43418);
nand U43788 (N_43788,N_43418,N_43379);
xor U43789 (N_43789,N_43477,N_43064);
nand U43790 (N_43790,N_43348,N_43021);
and U43791 (N_43791,N_43179,N_43204);
nor U43792 (N_43792,N_43194,N_43025);
nand U43793 (N_43793,N_43404,N_43221);
nand U43794 (N_43794,N_43215,N_43401);
xnor U43795 (N_43795,N_43153,N_43243);
nor U43796 (N_43796,N_43390,N_43052);
nand U43797 (N_43797,N_43176,N_43070);
nand U43798 (N_43798,N_43042,N_43232);
nand U43799 (N_43799,N_43258,N_43327);
nand U43800 (N_43800,N_43130,N_43339);
nand U43801 (N_43801,N_43111,N_43156);
nor U43802 (N_43802,N_43297,N_43181);
and U43803 (N_43803,N_43244,N_43438);
nand U43804 (N_43804,N_43483,N_43154);
or U43805 (N_43805,N_43320,N_43110);
nor U43806 (N_43806,N_43021,N_43339);
nand U43807 (N_43807,N_43168,N_43392);
nand U43808 (N_43808,N_43244,N_43186);
xor U43809 (N_43809,N_43428,N_43003);
or U43810 (N_43810,N_43325,N_43357);
xor U43811 (N_43811,N_43155,N_43338);
xor U43812 (N_43812,N_43072,N_43410);
nor U43813 (N_43813,N_43362,N_43283);
nor U43814 (N_43814,N_43468,N_43413);
nand U43815 (N_43815,N_43201,N_43215);
and U43816 (N_43816,N_43431,N_43401);
and U43817 (N_43817,N_43499,N_43456);
nor U43818 (N_43818,N_43117,N_43435);
xnor U43819 (N_43819,N_43303,N_43151);
nor U43820 (N_43820,N_43488,N_43306);
xor U43821 (N_43821,N_43382,N_43348);
nand U43822 (N_43822,N_43429,N_43200);
nand U43823 (N_43823,N_43396,N_43405);
nor U43824 (N_43824,N_43164,N_43487);
xnor U43825 (N_43825,N_43470,N_43280);
nand U43826 (N_43826,N_43376,N_43396);
nor U43827 (N_43827,N_43145,N_43354);
and U43828 (N_43828,N_43193,N_43465);
and U43829 (N_43829,N_43011,N_43046);
nor U43830 (N_43830,N_43193,N_43475);
xnor U43831 (N_43831,N_43151,N_43333);
nand U43832 (N_43832,N_43218,N_43337);
nand U43833 (N_43833,N_43371,N_43243);
and U43834 (N_43834,N_43277,N_43079);
and U43835 (N_43835,N_43007,N_43094);
nand U43836 (N_43836,N_43222,N_43275);
and U43837 (N_43837,N_43030,N_43194);
and U43838 (N_43838,N_43297,N_43046);
xnor U43839 (N_43839,N_43091,N_43054);
nand U43840 (N_43840,N_43142,N_43347);
and U43841 (N_43841,N_43490,N_43259);
nor U43842 (N_43842,N_43002,N_43108);
or U43843 (N_43843,N_43450,N_43281);
nor U43844 (N_43844,N_43017,N_43203);
nor U43845 (N_43845,N_43066,N_43175);
or U43846 (N_43846,N_43412,N_43193);
or U43847 (N_43847,N_43412,N_43241);
and U43848 (N_43848,N_43252,N_43165);
xor U43849 (N_43849,N_43365,N_43013);
or U43850 (N_43850,N_43497,N_43291);
xor U43851 (N_43851,N_43188,N_43438);
xor U43852 (N_43852,N_43423,N_43181);
nor U43853 (N_43853,N_43472,N_43141);
nor U43854 (N_43854,N_43496,N_43023);
or U43855 (N_43855,N_43420,N_43484);
xnor U43856 (N_43856,N_43233,N_43167);
nor U43857 (N_43857,N_43014,N_43215);
nor U43858 (N_43858,N_43294,N_43494);
xnor U43859 (N_43859,N_43005,N_43415);
and U43860 (N_43860,N_43434,N_43018);
and U43861 (N_43861,N_43223,N_43226);
nor U43862 (N_43862,N_43425,N_43447);
or U43863 (N_43863,N_43334,N_43083);
nand U43864 (N_43864,N_43488,N_43229);
or U43865 (N_43865,N_43390,N_43302);
and U43866 (N_43866,N_43085,N_43442);
and U43867 (N_43867,N_43321,N_43493);
nor U43868 (N_43868,N_43361,N_43291);
and U43869 (N_43869,N_43369,N_43059);
nand U43870 (N_43870,N_43088,N_43459);
nor U43871 (N_43871,N_43437,N_43369);
nor U43872 (N_43872,N_43082,N_43216);
nor U43873 (N_43873,N_43098,N_43234);
nand U43874 (N_43874,N_43434,N_43421);
nor U43875 (N_43875,N_43091,N_43152);
and U43876 (N_43876,N_43025,N_43480);
xnor U43877 (N_43877,N_43435,N_43197);
xnor U43878 (N_43878,N_43326,N_43034);
xnor U43879 (N_43879,N_43460,N_43040);
nor U43880 (N_43880,N_43084,N_43271);
xnor U43881 (N_43881,N_43040,N_43098);
nor U43882 (N_43882,N_43255,N_43091);
nor U43883 (N_43883,N_43402,N_43160);
or U43884 (N_43884,N_43010,N_43081);
nor U43885 (N_43885,N_43199,N_43425);
xnor U43886 (N_43886,N_43231,N_43143);
or U43887 (N_43887,N_43440,N_43174);
nor U43888 (N_43888,N_43089,N_43316);
or U43889 (N_43889,N_43411,N_43469);
or U43890 (N_43890,N_43370,N_43419);
nand U43891 (N_43891,N_43222,N_43318);
xnor U43892 (N_43892,N_43324,N_43429);
nor U43893 (N_43893,N_43329,N_43369);
or U43894 (N_43894,N_43117,N_43056);
and U43895 (N_43895,N_43349,N_43282);
nand U43896 (N_43896,N_43459,N_43260);
and U43897 (N_43897,N_43082,N_43489);
xor U43898 (N_43898,N_43193,N_43253);
nor U43899 (N_43899,N_43350,N_43471);
and U43900 (N_43900,N_43241,N_43181);
or U43901 (N_43901,N_43498,N_43102);
and U43902 (N_43902,N_43489,N_43166);
and U43903 (N_43903,N_43041,N_43271);
xnor U43904 (N_43904,N_43069,N_43476);
nor U43905 (N_43905,N_43160,N_43156);
and U43906 (N_43906,N_43334,N_43001);
or U43907 (N_43907,N_43453,N_43125);
xnor U43908 (N_43908,N_43071,N_43331);
xor U43909 (N_43909,N_43312,N_43265);
xor U43910 (N_43910,N_43317,N_43245);
or U43911 (N_43911,N_43233,N_43329);
or U43912 (N_43912,N_43399,N_43165);
nand U43913 (N_43913,N_43138,N_43256);
nor U43914 (N_43914,N_43454,N_43415);
or U43915 (N_43915,N_43421,N_43197);
or U43916 (N_43916,N_43488,N_43175);
xnor U43917 (N_43917,N_43315,N_43034);
xnor U43918 (N_43918,N_43035,N_43272);
xor U43919 (N_43919,N_43174,N_43045);
nor U43920 (N_43920,N_43029,N_43261);
and U43921 (N_43921,N_43266,N_43214);
xnor U43922 (N_43922,N_43463,N_43482);
nand U43923 (N_43923,N_43322,N_43224);
nor U43924 (N_43924,N_43464,N_43327);
nand U43925 (N_43925,N_43123,N_43159);
or U43926 (N_43926,N_43274,N_43405);
or U43927 (N_43927,N_43048,N_43488);
nor U43928 (N_43928,N_43102,N_43375);
xnor U43929 (N_43929,N_43105,N_43125);
or U43930 (N_43930,N_43180,N_43054);
or U43931 (N_43931,N_43027,N_43359);
or U43932 (N_43932,N_43374,N_43491);
xnor U43933 (N_43933,N_43179,N_43330);
and U43934 (N_43934,N_43121,N_43349);
xor U43935 (N_43935,N_43349,N_43331);
and U43936 (N_43936,N_43090,N_43004);
or U43937 (N_43937,N_43464,N_43186);
nand U43938 (N_43938,N_43497,N_43360);
and U43939 (N_43939,N_43213,N_43026);
nor U43940 (N_43940,N_43481,N_43208);
nor U43941 (N_43941,N_43381,N_43383);
nor U43942 (N_43942,N_43158,N_43017);
xor U43943 (N_43943,N_43195,N_43158);
and U43944 (N_43944,N_43422,N_43118);
xnor U43945 (N_43945,N_43176,N_43496);
and U43946 (N_43946,N_43338,N_43116);
xnor U43947 (N_43947,N_43217,N_43174);
xnor U43948 (N_43948,N_43265,N_43229);
nand U43949 (N_43949,N_43385,N_43374);
and U43950 (N_43950,N_43273,N_43183);
xnor U43951 (N_43951,N_43093,N_43075);
or U43952 (N_43952,N_43112,N_43108);
xnor U43953 (N_43953,N_43004,N_43111);
nand U43954 (N_43954,N_43466,N_43438);
nor U43955 (N_43955,N_43157,N_43485);
xnor U43956 (N_43956,N_43008,N_43005);
and U43957 (N_43957,N_43250,N_43016);
xnor U43958 (N_43958,N_43072,N_43235);
and U43959 (N_43959,N_43360,N_43008);
nand U43960 (N_43960,N_43477,N_43222);
and U43961 (N_43961,N_43484,N_43324);
nor U43962 (N_43962,N_43154,N_43047);
or U43963 (N_43963,N_43234,N_43374);
xor U43964 (N_43964,N_43346,N_43109);
nand U43965 (N_43965,N_43252,N_43462);
xnor U43966 (N_43966,N_43092,N_43476);
xnor U43967 (N_43967,N_43179,N_43281);
xnor U43968 (N_43968,N_43227,N_43015);
nor U43969 (N_43969,N_43264,N_43384);
or U43970 (N_43970,N_43429,N_43081);
nor U43971 (N_43971,N_43120,N_43445);
or U43972 (N_43972,N_43276,N_43162);
and U43973 (N_43973,N_43104,N_43039);
and U43974 (N_43974,N_43127,N_43158);
and U43975 (N_43975,N_43437,N_43338);
xor U43976 (N_43976,N_43154,N_43161);
nand U43977 (N_43977,N_43451,N_43002);
xnor U43978 (N_43978,N_43487,N_43054);
or U43979 (N_43979,N_43058,N_43190);
xor U43980 (N_43980,N_43082,N_43305);
xor U43981 (N_43981,N_43126,N_43085);
nand U43982 (N_43982,N_43245,N_43286);
or U43983 (N_43983,N_43289,N_43010);
or U43984 (N_43984,N_43479,N_43061);
nand U43985 (N_43985,N_43285,N_43023);
nor U43986 (N_43986,N_43439,N_43155);
and U43987 (N_43987,N_43196,N_43042);
nand U43988 (N_43988,N_43442,N_43287);
nand U43989 (N_43989,N_43234,N_43115);
and U43990 (N_43990,N_43184,N_43182);
and U43991 (N_43991,N_43069,N_43479);
nor U43992 (N_43992,N_43093,N_43111);
xnor U43993 (N_43993,N_43211,N_43030);
or U43994 (N_43994,N_43332,N_43103);
nor U43995 (N_43995,N_43474,N_43009);
xor U43996 (N_43996,N_43221,N_43356);
and U43997 (N_43997,N_43346,N_43471);
nor U43998 (N_43998,N_43172,N_43412);
xor U43999 (N_43999,N_43410,N_43317);
and U44000 (N_44000,N_43809,N_43552);
xor U44001 (N_44001,N_43556,N_43919);
nand U44002 (N_44002,N_43584,N_43637);
or U44003 (N_44003,N_43751,N_43537);
or U44004 (N_44004,N_43957,N_43638);
or U44005 (N_44005,N_43850,N_43807);
or U44006 (N_44006,N_43626,N_43539);
and U44007 (N_44007,N_43906,N_43649);
nor U44008 (N_44008,N_43814,N_43632);
or U44009 (N_44009,N_43826,N_43565);
nor U44010 (N_44010,N_43846,N_43530);
nand U44011 (N_44011,N_43593,N_43643);
nor U44012 (N_44012,N_43761,N_43998);
or U44013 (N_44013,N_43728,N_43679);
nand U44014 (N_44014,N_43705,N_43877);
xor U44015 (N_44015,N_43922,N_43940);
nor U44016 (N_44016,N_43516,N_43839);
or U44017 (N_44017,N_43609,N_43722);
nand U44018 (N_44018,N_43640,N_43520);
xor U44019 (N_44019,N_43712,N_43695);
or U44020 (N_44020,N_43575,N_43574);
or U44021 (N_44021,N_43996,N_43929);
nor U44022 (N_44022,N_43675,N_43543);
xor U44023 (N_44023,N_43691,N_43799);
xor U44024 (N_44024,N_43931,N_43732);
xnor U44025 (N_44025,N_43849,N_43604);
xor U44026 (N_44026,N_43865,N_43914);
nand U44027 (N_44027,N_43968,N_43887);
or U44028 (N_44028,N_43829,N_43548);
or U44029 (N_44029,N_43650,N_43591);
and U44030 (N_44030,N_43708,N_43738);
nand U44031 (N_44031,N_43923,N_43731);
xnor U44032 (N_44032,N_43802,N_43724);
nor U44033 (N_44033,N_43874,N_43557);
nand U44034 (N_44034,N_43803,N_43966);
nand U44035 (N_44035,N_43958,N_43563);
or U44036 (N_44036,N_43955,N_43676);
or U44037 (N_44037,N_43735,N_43525);
or U44038 (N_44038,N_43586,N_43875);
or U44039 (N_44039,N_43930,N_43827);
nor U44040 (N_44040,N_43583,N_43717);
nor U44041 (N_44041,N_43685,N_43746);
nand U44042 (N_44042,N_43531,N_43805);
xnor U44043 (N_44043,N_43924,N_43707);
and U44044 (N_44044,N_43630,N_43793);
and U44045 (N_44045,N_43851,N_43665);
and U44046 (N_44046,N_43784,N_43641);
and U44047 (N_44047,N_43519,N_43551);
or U44048 (N_44048,N_43673,N_43892);
xor U44049 (N_44049,N_43739,N_43939);
or U44050 (N_44050,N_43750,N_43536);
nor U44051 (N_44051,N_43507,N_43611);
or U44052 (N_44052,N_43830,N_43541);
and U44053 (N_44053,N_43606,N_43843);
nand U44054 (N_44054,N_43510,N_43704);
nand U44055 (N_44055,N_43748,N_43734);
nand U44056 (N_44056,N_43896,N_43585);
nand U44057 (N_44057,N_43813,N_43866);
nand U44058 (N_44058,N_43771,N_43975);
and U44059 (N_44059,N_43797,N_43812);
xor U44060 (N_44060,N_43648,N_43895);
xor U44061 (N_44061,N_43686,N_43835);
nor U44062 (N_44062,N_43757,N_43971);
nor U44063 (N_44063,N_43762,N_43512);
or U44064 (N_44064,N_43654,N_43969);
and U44065 (N_44065,N_43566,N_43780);
xor U44066 (N_44066,N_43999,N_43607);
and U44067 (N_44067,N_43727,N_43703);
nor U44068 (N_44068,N_43942,N_43657);
nand U44069 (N_44069,N_43687,N_43639);
nand U44070 (N_44070,N_43845,N_43909);
and U44071 (N_44071,N_43621,N_43786);
nand U44072 (N_44072,N_43625,N_43898);
or U44073 (N_44073,N_43964,N_43573);
xnor U44074 (N_44074,N_43822,N_43936);
nor U44075 (N_44075,N_43821,N_43555);
nor U44076 (N_44076,N_43804,N_43989);
nor U44077 (N_44077,N_43546,N_43571);
and U44078 (N_44078,N_43943,N_43538);
nor U44079 (N_44079,N_43925,N_43860);
xnor U44080 (N_44080,N_43505,N_43858);
or U44081 (N_44081,N_43733,N_43913);
and U44082 (N_44082,N_43580,N_43721);
nand U44083 (N_44083,N_43915,N_43535);
and U44084 (N_44084,N_43970,N_43868);
or U44085 (N_44085,N_43698,N_43579);
or U44086 (N_44086,N_43619,N_43545);
nor U44087 (N_44087,N_43715,N_43774);
nand U44088 (N_44088,N_43997,N_43542);
xor U44089 (N_44089,N_43979,N_43980);
or U44090 (N_44090,N_43963,N_43859);
xor U44091 (N_44091,N_43590,N_43529);
nor U44092 (N_44092,N_43718,N_43599);
xnor U44093 (N_44093,N_43720,N_43681);
nand U44094 (N_44094,N_43932,N_43689);
xnor U44095 (N_44095,N_43948,N_43974);
and U44096 (N_44096,N_43792,N_43743);
nor U44097 (N_44097,N_43862,N_43987);
or U44098 (N_44098,N_43820,N_43674);
xor U44099 (N_44099,N_43816,N_43570);
nand U44100 (N_44100,N_43918,N_43944);
xor U44101 (N_44101,N_43785,N_43569);
nor U44102 (N_44102,N_43842,N_43897);
xor U44103 (N_44103,N_43811,N_43636);
nand U44104 (N_44104,N_43995,N_43564);
or U44105 (N_44105,N_43962,N_43700);
and U44106 (N_44106,N_43628,N_43755);
nand U44107 (N_44107,N_43992,N_43946);
nand U44108 (N_44108,N_43870,N_43624);
nor U44109 (N_44109,N_43938,N_43941);
xor U44110 (N_44110,N_43978,N_43553);
and U44111 (N_44111,N_43560,N_43869);
nor U44112 (N_44112,N_43756,N_43795);
nand U44113 (N_44113,N_43965,N_43776);
nor U44114 (N_44114,N_43711,N_43781);
xor U44115 (N_44115,N_43582,N_43916);
or U44116 (N_44116,N_43982,N_43894);
and U44117 (N_44117,N_43810,N_43884);
nor U44118 (N_44118,N_43881,N_43608);
nand U44119 (N_44119,N_43752,N_43680);
or U44120 (N_44120,N_43701,N_43514);
nand U44121 (N_44121,N_43764,N_43873);
xnor U44122 (N_44122,N_43672,N_43986);
xor U44123 (N_44123,N_43838,N_43824);
nor U44124 (N_44124,N_43544,N_43620);
and U44125 (N_44125,N_43782,N_43837);
nand U44126 (N_44126,N_43614,N_43900);
nand U44127 (N_44127,N_43719,N_43652);
or U44128 (N_44128,N_43840,N_43935);
nor U44129 (N_44129,N_43864,N_43693);
or U44130 (N_44130,N_43800,N_43984);
nor U44131 (N_44131,N_43947,N_43567);
xor U44132 (N_44132,N_43902,N_43668);
or U44133 (N_44133,N_43778,N_43753);
xnor U44134 (N_44134,N_43857,N_43832);
xor U44135 (N_44135,N_43907,N_43716);
and U44136 (N_44136,N_43549,N_43889);
or U44137 (N_44137,N_43759,N_43767);
nor U44138 (N_44138,N_43796,N_43863);
nor U44139 (N_44139,N_43928,N_43819);
nor U44140 (N_44140,N_43888,N_43741);
and U44141 (N_44141,N_43742,N_43550);
nand U44142 (N_44142,N_43522,N_43815);
nor U44143 (N_44143,N_43736,N_43595);
nor U44144 (N_44144,N_43794,N_43667);
or U44145 (N_44145,N_43508,N_43952);
and U44146 (N_44146,N_43683,N_43901);
nor U44147 (N_44147,N_43616,N_43500);
nand U44148 (N_44148,N_43749,N_43745);
xnor U44149 (N_44149,N_43853,N_43951);
nor U44150 (N_44150,N_43910,N_43502);
or U44151 (N_44151,N_43589,N_43880);
nor U44152 (N_44152,N_43765,N_43920);
and U44153 (N_44153,N_43893,N_43867);
and U44154 (N_44154,N_43671,N_43828);
and U44155 (N_44155,N_43713,N_43823);
or U44156 (N_44156,N_43769,N_43655);
nand U44157 (N_44157,N_43788,N_43981);
or U44158 (N_44158,N_43528,N_43953);
nand U44159 (N_44159,N_43592,N_43760);
nor U44160 (N_44160,N_43532,N_43959);
nor U44161 (N_44161,N_43527,N_43891);
xnor U44162 (N_44162,N_43740,N_43775);
nand U44163 (N_44163,N_43598,N_43678);
xnor U44164 (N_44164,N_43988,N_43706);
or U44165 (N_44165,N_43945,N_43991);
xnor U44166 (N_44166,N_43696,N_43967);
xor U44167 (N_44167,N_43730,N_43770);
xor U44168 (N_44168,N_43661,N_43601);
nand U44169 (N_44169,N_43596,N_43533);
and U44170 (N_44170,N_43600,N_43977);
nand U44171 (N_44171,N_43871,N_43677);
or U44172 (N_44172,N_43956,N_43976);
nor U44173 (N_44173,N_43882,N_43856);
nor U44174 (N_44174,N_43872,N_43806);
nand U44175 (N_44175,N_43526,N_43576);
or U44176 (N_44176,N_43656,N_43773);
nand U44177 (N_44177,N_43983,N_43670);
nand U44178 (N_44178,N_43825,N_43990);
nor U44179 (N_44179,N_43899,N_43682);
xnor U44180 (N_44180,N_43554,N_43768);
nor U44181 (N_44181,N_43578,N_43833);
nor U44182 (N_44182,N_43623,N_43503);
nand U44183 (N_44183,N_43699,N_43848);
and U44184 (N_44184,N_43783,N_43801);
xor U44185 (N_44185,N_43808,N_43697);
nor U44186 (N_44186,N_43613,N_43917);
nor U44187 (N_44187,N_43985,N_43644);
xnor U44188 (N_44188,N_43534,N_43993);
nand U44189 (N_44189,N_43660,N_43777);
or U44190 (N_44190,N_43927,N_43635);
nor U44191 (N_44191,N_43577,N_43836);
xnor U44192 (N_44192,N_43523,N_43663);
or U44193 (N_44193,N_43562,N_43587);
and U44194 (N_44194,N_43876,N_43540);
nand U44195 (N_44195,N_43588,N_43921);
nand U44196 (N_44196,N_43518,N_43949);
and U44197 (N_44197,N_43817,N_43688);
nor U44198 (N_44198,N_43912,N_43852);
or U44199 (N_44199,N_43911,N_43798);
and U44200 (N_44200,N_43779,N_43818);
nand U44201 (N_44201,N_43631,N_43766);
nor U44202 (N_44202,N_43506,N_43615);
or U44203 (N_44203,N_43702,N_43511);
and U44204 (N_44204,N_43885,N_43725);
xnor U44205 (N_44205,N_43581,N_43847);
or U44206 (N_44206,N_43610,N_43513);
nand U44207 (N_44207,N_43690,N_43934);
nor U44208 (N_44208,N_43950,N_43629);
or U44209 (N_44209,N_43612,N_43758);
nor U44210 (N_44210,N_43855,N_43890);
nand U44211 (N_44211,N_43694,N_43961);
and U44212 (N_44212,N_43926,N_43617);
nor U44213 (N_44213,N_43933,N_43572);
nand U44214 (N_44214,N_43954,N_43729);
nand U44215 (N_44215,N_43501,N_43905);
or U44216 (N_44216,N_43664,N_43618);
nand U44217 (N_44217,N_43658,N_43646);
or U44218 (N_44218,N_43504,N_43878);
nand U44219 (N_44219,N_43561,N_43831);
and U44220 (N_44220,N_43960,N_43714);
nand U44221 (N_44221,N_43559,N_43515);
nand U44222 (N_44222,N_43622,N_43627);
or U44223 (N_44223,N_43904,N_43908);
nand U44224 (N_44224,N_43603,N_43633);
or U44225 (N_44225,N_43747,N_43547);
nand U44226 (N_44226,N_43726,N_43709);
xor U44227 (N_44227,N_43597,N_43854);
xnor U44228 (N_44228,N_43509,N_43642);
or U44229 (N_44229,N_43653,N_43651);
or U44230 (N_44230,N_43789,N_43879);
nor U44231 (N_44231,N_43973,N_43841);
or U44232 (N_44232,N_43659,N_43861);
or U44233 (N_44233,N_43568,N_43744);
nor U44234 (N_44234,N_43790,N_43517);
or U44235 (N_44235,N_43937,N_43723);
and U44236 (N_44236,N_43524,N_43692);
or U44237 (N_44237,N_43710,N_43594);
and U44238 (N_44238,N_43684,N_43886);
or U44239 (N_44239,N_43754,N_43662);
or U44240 (N_44240,N_43903,N_43834);
nand U44241 (N_44241,N_43647,N_43791);
nor U44242 (N_44242,N_43521,N_43763);
nor U44243 (N_44243,N_43605,N_43669);
and U44244 (N_44244,N_43634,N_43994);
nor U44245 (N_44245,N_43737,N_43787);
xnor U44246 (N_44246,N_43602,N_43645);
and U44247 (N_44247,N_43558,N_43844);
and U44248 (N_44248,N_43972,N_43772);
xnor U44249 (N_44249,N_43883,N_43666);
and U44250 (N_44250,N_43633,N_43711);
xor U44251 (N_44251,N_43607,N_43761);
nand U44252 (N_44252,N_43646,N_43978);
xor U44253 (N_44253,N_43949,N_43797);
and U44254 (N_44254,N_43548,N_43782);
and U44255 (N_44255,N_43978,N_43548);
or U44256 (N_44256,N_43777,N_43696);
xnor U44257 (N_44257,N_43607,N_43963);
and U44258 (N_44258,N_43722,N_43851);
nor U44259 (N_44259,N_43835,N_43895);
and U44260 (N_44260,N_43576,N_43821);
nand U44261 (N_44261,N_43846,N_43645);
nor U44262 (N_44262,N_43765,N_43526);
nand U44263 (N_44263,N_43628,N_43954);
and U44264 (N_44264,N_43690,N_43919);
nand U44265 (N_44265,N_43707,N_43733);
xor U44266 (N_44266,N_43678,N_43758);
xor U44267 (N_44267,N_43951,N_43646);
nor U44268 (N_44268,N_43827,N_43781);
or U44269 (N_44269,N_43667,N_43798);
nand U44270 (N_44270,N_43954,N_43505);
nand U44271 (N_44271,N_43568,N_43588);
nor U44272 (N_44272,N_43865,N_43877);
nor U44273 (N_44273,N_43845,N_43535);
or U44274 (N_44274,N_43546,N_43728);
and U44275 (N_44275,N_43660,N_43900);
or U44276 (N_44276,N_43965,N_43583);
and U44277 (N_44277,N_43980,N_43716);
and U44278 (N_44278,N_43647,N_43924);
xnor U44279 (N_44279,N_43660,N_43969);
or U44280 (N_44280,N_43759,N_43905);
and U44281 (N_44281,N_43501,N_43890);
xor U44282 (N_44282,N_43505,N_43658);
or U44283 (N_44283,N_43955,N_43537);
nor U44284 (N_44284,N_43773,N_43704);
nand U44285 (N_44285,N_43606,N_43737);
xor U44286 (N_44286,N_43578,N_43516);
and U44287 (N_44287,N_43923,N_43500);
or U44288 (N_44288,N_43652,N_43546);
nand U44289 (N_44289,N_43944,N_43657);
and U44290 (N_44290,N_43523,N_43759);
or U44291 (N_44291,N_43503,N_43556);
xnor U44292 (N_44292,N_43924,N_43880);
nand U44293 (N_44293,N_43900,N_43743);
or U44294 (N_44294,N_43920,N_43833);
nor U44295 (N_44295,N_43604,N_43721);
or U44296 (N_44296,N_43931,N_43809);
nand U44297 (N_44297,N_43569,N_43523);
or U44298 (N_44298,N_43913,N_43730);
and U44299 (N_44299,N_43801,N_43907);
nor U44300 (N_44300,N_43894,N_43617);
or U44301 (N_44301,N_43567,N_43869);
or U44302 (N_44302,N_43649,N_43959);
and U44303 (N_44303,N_43782,N_43527);
nor U44304 (N_44304,N_43642,N_43976);
nor U44305 (N_44305,N_43835,N_43940);
nand U44306 (N_44306,N_43601,N_43752);
or U44307 (N_44307,N_43881,N_43706);
xor U44308 (N_44308,N_43853,N_43988);
and U44309 (N_44309,N_43503,N_43847);
or U44310 (N_44310,N_43647,N_43874);
or U44311 (N_44311,N_43876,N_43546);
nand U44312 (N_44312,N_43966,N_43683);
nor U44313 (N_44313,N_43593,N_43885);
nand U44314 (N_44314,N_43907,N_43736);
nor U44315 (N_44315,N_43630,N_43700);
nand U44316 (N_44316,N_43851,N_43684);
or U44317 (N_44317,N_43718,N_43993);
or U44318 (N_44318,N_43723,N_43769);
nor U44319 (N_44319,N_43737,N_43768);
xnor U44320 (N_44320,N_43937,N_43965);
or U44321 (N_44321,N_43542,N_43944);
or U44322 (N_44322,N_43600,N_43533);
xor U44323 (N_44323,N_43718,N_43866);
nand U44324 (N_44324,N_43604,N_43638);
nand U44325 (N_44325,N_43557,N_43971);
nor U44326 (N_44326,N_43754,N_43747);
nand U44327 (N_44327,N_43581,N_43983);
nor U44328 (N_44328,N_43784,N_43982);
and U44329 (N_44329,N_43641,N_43894);
nand U44330 (N_44330,N_43614,N_43622);
nor U44331 (N_44331,N_43967,N_43507);
nor U44332 (N_44332,N_43678,N_43847);
nand U44333 (N_44333,N_43998,N_43611);
or U44334 (N_44334,N_43880,N_43500);
xor U44335 (N_44335,N_43848,N_43608);
nor U44336 (N_44336,N_43579,N_43782);
and U44337 (N_44337,N_43693,N_43836);
nor U44338 (N_44338,N_43629,N_43579);
nor U44339 (N_44339,N_43760,N_43516);
nor U44340 (N_44340,N_43508,N_43674);
or U44341 (N_44341,N_43642,N_43736);
xnor U44342 (N_44342,N_43767,N_43867);
nor U44343 (N_44343,N_43781,N_43806);
or U44344 (N_44344,N_43994,N_43643);
or U44345 (N_44345,N_43859,N_43662);
xnor U44346 (N_44346,N_43950,N_43535);
and U44347 (N_44347,N_43716,N_43645);
or U44348 (N_44348,N_43519,N_43991);
xnor U44349 (N_44349,N_43750,N_43609);
xnor U44350 (N_44350,N_43689,N_43551);
or U44351 (N_44351,N_43549,N_43698);
nor U44352 (N_44352,N_43976,N_43622);
nor U44353 (N_44353,N_43664,N_43669);
nor U44354 (N_44354,N_43845,N_43780);
or U44355 (N_44355,N_43604,N_43685);
nor U44356 (N_44356,N_43814,N_43969);
nand U44357 (N_44357,N_43642,N_43658);
xnor U44358 (N_44358,N_43862,N_43928);
nor U44359 (N_44359,N_43573,N_43791);
and U44360 (N_44360,N_43832,N_43881);
or U44361 (N_44361,N_43703,N_43888);
and U44362 (N_44362,N_43661,N_43967);
nor U44363 (N_44363,N_43746,N_43970);
nor U44364 (N_44364,N_43555,N_43810);
xor U44365 (N_44365,N_43720,N_43827);
or U44366 (N_44366,N_43983,N_43590);
nand U44367 (N_44367,N_43849,N_43774);
xnor U44368 (N_44368,N_43510,N_43889);
xnor U44369 (N_44369,N_43788,N_43920);
and U44370 (N_44370,N_43690,N_43967);
and U44371 (N_44371,N_43873,N_43541);
or U44372 (N_44372,N_43939,N_43502);
xnor U44373 (N_44373,N_43929,N_43535);
nand U44374 (N_44374,N_43655,N_43658);
nand U44375 (N_44375,N_43864,N_43960);
nor U44376 (N_44376,N_43597,N_43893);
nor U44377 (N_44377,N_43834,N_43942);
nand U44378 (N_44378,N_43816,N_43878);
nand U44379 (N_44379,N_43733,N_43979);
and U44380 (N_44380,N_43501,N_43885);
and U44381 (N_44381,N_43556,N_43595);
nand U44382 (N_44382,N_43908,N_43582);
and U44383 (N_44383,N_43716,N_43622);
and U44384 (N_44384,N_43968,N_43690);
nand U44385 (N_44385,N_43728,N_43700);
nor U44386 (N_44386,N_43590,N_43719);
nand U44387 (N_44387,N_43808,N_43978);
xnor U44388 (N_44388,N_43976,N_43523);
nand U44389 (N_44389,N_43786,N_43766);
or U44390 (N_44390,N_43798,N_43535);
xor U44391 (N_44391,N_43576,N_43842);
and U44392 (N_44392,N_43620,N_43958);
nand U44393 (N_44393,N_43602,N_43516);
and U44394 (N_44394,N_43880,N_43911);
xor U44395 (N_44395,N_43615,N_43917);
or U44396 (N_44396,N_43537,N_43534);
xor U44397 (N_44397,N_43550,N_43764);
or U44398 (N_44398,N_43835,N_43682);
nand U44399 (N_44399,N_43740,N_43712);
nand U44400 (N_44400,N_43584,N_43531);
and U44401 (N_44401,N_43525,N_43798);
or U44402 (N_44402,N_43682,N_43555);
and U44403 (N_44403,N_43867,N_43630);
nor U44404 (N_44404,N_43980,N_43718);
xor U44405 (N_44405,N_43533,N_43781);
nor U44406 (N_44406,N_43672,N_43532);
nor U44407 (N_44407,N_43789,N_43744);
nand U44408 (N_44408,N_43553,N_43828);
nor U44409 (N_44409,N_43966,N_43935);
xnor U44410 (N_44410,N_43793,N_43651);
nor U44411 (N_44411,N_43887,N_43697);
nand U44412 (N_44412,N_43969,N_43738);
xnor U44413 (N_44413,N_43980,N_43652);
and U44414 (N_44414,N_43634,N_43726);
nand U44415 (N_44415,N_43961,N_43897);
nor U44416 (N_44416,N_43996,N_43812);
and U44417 (N_44417,N_43667,N_43698);
nor U44418 (N_44418,N_43625,N_43520);
nor U44419 (N_44419,N_43869,N_43999);
nand U44420 (N_44420,N_43818,N_43771);
and U44421 (N_44421,N_43726,N_43628);
nand U44422 (N_44422,N_43688,N_43788);
or U44423 (N_44423,N_43523,N_43556);
nor U44424 (N_44424,N_43652,N_43735);
nor U44425 (N_44425,N_43604,N_43689);
nand U44426 (N_44426,N_43763,N_43586);
or U44427 (N_44427,N_43560,N_43851);
xor U44428 (N_44428,N_43691,N_43738);
nand U44429 (N_44429,N_43910,N_43735);
nand U44430 (N_44430,N_43585,N_43862);
xnor U44431 (N_44431,N_43520,N_43865);
or U44432 (N_44432,N_43910,N_43659);
and U44433 (N_44433,N_43844,N_43876);
nand U44434 (N_44434,N_43908,N_43882);
and U44435 (N_44435,N_43948,N_43795);
and U44436 (N_44436,N_43861,N_43802);
and U44437 (N_44437,N_43549,N_43722);
and U44438 (N_44438,N_43801,N_43975);
or U44439 (N_44439,N_43702,N_43911);
or U44440 (N_44440,N_43898,N_43605);
nand U44441 (N_44441,N_43626,N_43834);
nor U44442 (N_44442,N_43800,N_43862);
and U44443 (N_44443,N_43760,N_43786);
or U44444 (N_44444,N_43722,N_43905);
nand U44445 (N_44445,N_43921,N_43739);
nor U44446 (N_44446,N_43874,N_43697);
nor U44447 (N_44447,N_43667,N_43937);
nor U44448 (N_44448,N_43789,N_43540);
nand U44449 (N_44449,N_43930,N_43507);
and U44450 (N_44450,N_43508,N_43732);
xor U44451 (N_44451,N_43785,N_43518);
xor U44452 (N_44452,N_43884,N_43518);
nor U44453 (N_44453,N_43917,N_43897);
and U44454 (N_44454,N_43882,N_43903);
or U44455 (N_44455,N_43801,N_43838);
nand U44456 (N_44456,N_43748,N_43638);
nor U44457 (N_44457,N_43662,N_43653);
xnor U44458 (N_44458,N_43947,N_43664);
or U44459 (N_44459,N_43534,N_43516);
and U44460 (N_44460,N_43876,N_43809);
xor U44461 (N_44461,N_43620,N_43520);
and U44462 (N_44462,N_43769,N_43540);
or U44463 (N_44463,N_43870,N_43862);
nand U44464 (N_44464,N_43915,N_43779);
xnor U44465 (N_44465,N_43745,N_43544);
or U44466 (N_44466,N_43834,N_43845);
nor U44467 (N_44467,N_43988,N_43507);
nor U44468 (N_44468,N_43887,N_43992);
and U44469 (N_44469,N_43526,N_43848);
xor U44470 (N_44470,N_43671,N_43952);
xnor U44471 (N_44471,N_43599,N_43874);
nand U44472 (N_44472,N_43909,N_43751);
nand U44473 (N_44473,N_43738,N_43880);
and U44474 (N_44474,N_43682,N_43891);
or U44475 (N_44475,N_43521,N_43860);
nand U44476 (N_44476,N_43857,N_43844);
or U44477 (N_44477,N_43938,N_43786);
nand U44478 (N_44478,N_43520,N_43947);
and U44479 (N_44479,N_43678,N_43514);
xnor U44480 (N_44480,N_43953,N_43825);
nand U44481 (N_44481,N_43794,N_43777);
and U44482 (N_44482,N_43728,N_43842);
xnor U44483 (N_44483,N_43680,N_43865);
xnor U44484 (N_44484,N_43869,N_43696);
nand U44485 (N_44485,N_43978,N_43814);
or U44486 (N_44486,N_43700,N_43885);
and U44487 (N_44487,N_43841,N_43830);
xor U44488 (N_44488,N_43573,N_43899);
nor U44489 (N_44489,N_43928,N_43501);
nor U44490 (N_44490,N_43614,N_43628);
or U44491 (N_44491,N_43975,N_43822);
nor U44492 (N_44492,N_43657,N_43811);
or U44493 (N_44493,N_43946,N_43688);
nand U44494 (N_44494,N_43531,N_43735);
and U44495 (N_44495,N_43520,N_43944);
and U44496 (N_44496,N_43769,N_43770);
xor U44497 (N_44497,N_43873,N_43550);
or U44498 (N_44498,N_43811,N_43553);
nand U44499 (N_44499,N_43660,N_43894);
xor U44500 (N_44500,N_44355,N_44285);
nand U44501 (N_44501,N_44254,N_44033);
nor U44502 (N_44502,N_44329,N_44128);
or U44503 (N_44503,N_44093,N_44434);
xnor U44504 (N_44504,N_44428,N_44118);
xnor U44505 (N_44505,N_44133,N_44002);
xor U44506 (N_44506,N_44491,N_44039);
nand U44507 (N_44507,N_44288,N_44143);
xor U44508 (N_44508,N_44424,N_44494);
nor U44509 (N_44509,N_44216,N_44295);
nor U44510 (N_44510,N_44433,N_44200);
nor U44511 (N_44511,N_44098,N_44001);
and U44512 (N_44512,N_44299,N_44136);
nor U44513 (N_44513,N_44168,N_44248);
or U44514 (N_44514,N_44078,N_44201);
nor U44515 (N_44515,N_44478,N_44479);
nor U44516 (N_44516,N_44330,N_44403);
or U44517 (N_44517,N_44496,N_44090);
and U44518 (N_44518,N_44409,N_44317);
and U44519 (N_44519,N_44177,N_44184);
and U44520 (N_44520,N_44392,N_44206);
or U44521 (N_44521,N_44144,N_44182);
nand U44522 (N_44522,N_44237,N_44176);
or U44523 (N_44523,N_44436,N_44296);
nand U44524 (N_44524,N_44287,N_44187);
nor U44525 (N_44525,N_44195,N_44351);
xnor U44526 (N_44526,N_44360,N_44461);
nor U44527 (N_44527,N_44464,N_44228);
nand U44528 (N_44528,N_44339,N_44394);
nand U44529 (N_44529,N_44475,N_44198);
nand U44530 (N_44530,N_44453,N_44476);
nand U44531 (N_44531,N_44325,N_44473);
xor U44532 (N_44532,N_44253,N_44042);
xnor U44533 (N_44533,N_44105,N_44352);
xor U44534 (N_44534,N_44115,N_44036);
and U44535 (N_44535,N_44192,N_44247);
and U44536 (N_44536,N_44114,N_44196);
nor U44537 (N_44537,N_44481,N_44463);
nand U44538 (N_44538,N_44414,N_44180);
xor U44539 (N_44539,N_44310,N_44175);
xor U44540 (N_44540,N_44334,N_44395);
and U44541 (N_44541,N_44112,N_44365);
xor U44542 (N_44542,N_44440,N_44493);
and U44543 (N_44543,N_44265,N_44448);
nor U44544 (N_44544,N_44354,N_44017);
nand U44545 (N_44545,N_44408,N_44263);
or U44546 (N_44546,N_44186,N_44495);
nor U44547 (N_44547,N_44024,N_44306);
nor U44548 (N_44548,N_44333,N_44243);
xor U44549 (N_44549,N_44122,N_44003);
or U44550 (N_44550,N_44223,N_44413);
or U44551 (N_44551,N_44350,N_44154);
nand U44552 (N_44552,N_44373,N_44009);
or U44553 (N_44553,N_44139,N_44239);
and U44554 (N_44554,N_44018,N_44362);
xnor U44555 (N_44555,N_44107,N_44415);
xnor U44556 (N_44556,N_44034,N_44435);
or U44557 (N_44557,N_44193,N_44369);
and U44558 (N_44558,N_44467,N_44474);
nor U44559 (N_44559,N_44205,N_44104);
or U44560 (N_44560,N_44393,N_44209);
nor U44561 (N_44561,N_44217,N_44286);
nor U44562 (N_44562,N_44095,N_44088);
xor U44563 (N_44563,N_44447,N_44173);
nand U44564 (N_44564,N_44137,N_44199);
and U44565 (N_44565,N_44170,N_44047);
and U44566 (N_44566,N_44082,N_44208);
xor U44567 (N_44567,N_44148,N_44004);
nor U44568 (N_44568,N_44059,N_44230);
nor U44569 (N_44569,N_44272,N_44138);
or U44570 (N_44570,N_44134,N_44449);
and U44571 (N_44571,N_44419,N_44101);
nand U44572 (N_44572,N_44212,N_44099);
nand U44573 (N_44573,N_44378,N_44280);
or U44574 (N_44574,N_44037,N_44404);
or U44575 (N_44575,N_44313,N_44353);
or U44576 (N_44576,N_44211,N_44357);
nand U44577 (N_44577,N_44091,N_44356);
or U44578 (N_44578,N_44062,N_44061);
or U44579 (N_44579,N_44087,N_44497);
nand U44580 (N_44580,N_44292,N_44163);
xor U44581 (N_44581,N_44048,N_44063);
or U44582 (N_44582,N_44049,N_44227);
or U44583 (N_44583,N_44194,N_44382);
xnor U44584 (N_44584,N_44197,N_44147);
or U44585 (N_44585,N_44152,N_44468);
nor U44586 (N_44586,N_44318,N_44273);
xnor U44587 (N_44587,N_44210,N_44301);
nand U44588 (N_44588,N_44086,N_44241);
nor U44589 (N_44589,N_44375,N_44162);
or U44590 (N_44590,N_44027,N_44387);
and U44591 (N_44591,N_44376,N_44271);
and U44592 (N_44592,N_44315,N_44055);
nand U44593 (N_44593,N_44056,N_44261);
xnor U44594 (N_44594,N_44269,N_44160);
nand U44595 (N_44595,N_44094,N_44251);
nand U44596 (N_44596,N_44486,N_44010);
xnor U44597 (N_44597,N_44281,N_44454);
or U44598 (N_44598,N_44399,N_44383);
or U44599 (N_44599,N_44283,N_44293);
nor U44600 (N_44600,N_44384,N_44172);
and U44601 (N_44601,N_44492,N_44322);
or U44602 (N_44602,N_44343,N_44290);
or U44603 (N_44603,N_44312,N_44423);
or U44604 (N_44604,N_44266,N_44060);
or U44605 (N_44605,N_44014,N_44308);
nand U44606 (N_44606,N_44234,N_44328);
nor U44607 (N_44607,N_44158,N_44368);
or U44608 (N_44608,N_44364,N_44074);
nor U44609 (N_44609,N_44401,N_44022);
nor U44610 (N_44610,N_44142,N_44275);
xnor U44611 (N_44611,N_44420,N_44080);
or U44612 (N_44612,N_44425,N_44096);
nand U44613 (N_44613,N_44097,N_44165);
nor U44614 (N_44614,N_44075,N_44013);
xnor U44615 (N_44615,N_44307,N_44438);
nor U44616 (N_44616,N_44057,N_44426);
xnor U44617 (N_44617,N_44381,N_44044);
nand U44618 (N_44618,N_44462,N_44072);
nand U44619 (N_44619,N_44242,N_44498);
nand U44620 (N_44620,N_44233,N_44316);
and U44621 (N_44621,N_44278,N_44410);
or U44622 (N_44622,N_44256,N_44458);
and U44623 (N_44623,N_44341,N_44077);
xor U44624 (N_44624,N_44366,N_44011);
and U44625 (N_44625,N_44260,N_44043);
nand U44626 (N_44626,N_44471,N_44477);
xnor U44627 (N_44627,N_44385,N_44250);
xnor U44628 (N_44628,N_44411,N_44314);
nand U44629 (N_44629,N_44178,N_44231);
and U44630 (N_44630,N_44167,N_44150);
xor U44631 (N_44631,N_44064,N_44370);
xor U44632 (N_44632,N_44084,N_44465);
and U44633 (N_44633,N_44116,N_44297);
nor U44634 (N_44634,N_44300,N_44050);
nor U44635 (N_44635,N_44085,N_44396);
xor U44636 (N_44636,N_44023,N_44021);
nor U44637 (N_44637,N_44008,N_44181);
nand U44638 (N_44638,N_44188,N_44157);
nand U44639 (N_44639,N_44470,N_44207);
and U44640 (N_44640,N_44252,N_44402);
nand U44641 (N_44641,N_44282,N_44026);
xor U44642 (N_44642,N_44397,N_44111);
nand U44643 (N_44643,N_44141,N_44416);
xnor U44644 (N_44644,N_44482,N_44390);
and U44645 (N_44645,N_44340,N_44145);
or U44646 (N_44646,N_44218,N_44102);
and U44647 (N_44647,N_44421,N_44274);
or U44648 (N_44648,N_44249,N_44345);
nand U44649 (N_44649,N_44130,N_44380);
nand U44650 (N_44650,N_44065,N_44069);
or U44651 (N_44651,N_44441,N_44444);
xnor U44652 (N_44652,N_44466,N_44119);
or U44653 (N_44653,N_44040,N_44156);
or U44654 (N_44654,N_44389,N_44359);
or U44655 (N_44655,N_44487,N_44391);
and U44656 (N_44656,N_44245,N_44452);
xnor U44657 (N_44657,N_44222,N_44108);
or U44658 (N_44658,N_44161,N_44131);
and U44659 (N_44659,N_44149,N_44405);
xnor U44660 (N_44660,N_44092,N_44321);
nor U44661 (N_44661,N_44164,N_44304);
or U44662 (N_44662,N_44073,N_44109);
or U44663 (N_44663,N_44371,N_44103);
and U44664 (N_44664,N_44019,N_44335);
and U44665 (N_44665,N_44146,N_44309);
nand U44666 (N_44666,N_44469,N_44202);
and U44667 (N_44667,N_44244,N_44015);
nor U44668 (N_44668,N_44025,N_44336);
and U44669 (N_44669,N_44456,N_44174);
xor U44670 (N_44670,N_44123,N_44153);
nand U44671 (N_44671,N_44262,N_44398);
or U44672 (N_44672,N_44289,N_44264);
and U44673 (N_44673,N_44132,N_44344);
nand U44674 (N_44674,N_44358,N_44298);
nor U44675 (N_44675,N_44220,N_44030);
nor U44676 (N_44676,N_44191,N_44028);
and U44677 (N_44677,N_44159,N_44459);
and U44678 (N_44678,N_44219,N_44437);
nor U44679 (N_44679,N_44291,N_44016);
or U44680 (N_44680,N_44430,N_44240);
xnor U44681 (N_44681,N_44327,N_44089);
or U44682 (N_44682,N_44054,N_44361);
nand U44683 (N_44683,N_44258,N_44499);
or U44684 (N_44684,N_44267,N_44007);
or U44685 (N_44685,N_44337,N_44113);
nand U44686 (N_44686,N_44045,N_44035);
or U44687 (N_44687,N_44129,N_44483);
and U44688 (N_44688,N_44100,N_44204);
and U44689 (N_44689,N_44412,N_44229);
or U44690 (N_44690,N_44224,N_44480);
xnor U44691 (N_44691,N_44140,N_44439);
xor U44692 (N_44692,N_44377,N_44268);
xor U44693 (N_44693,N_44257,N_44347);
nand U44694 (N_44694,N_44221,N_44071);
nand U44695 (N_44695,N_44422,N_44179);
xor U44696 (N_44696,N_44053,N_44490);
nor U44697 (N_44697,N_44276,N_44386);
xor U44698 (N_44698,N_44126,N_44000);
nand U44699 (N_44699,N_44379,N_44374);
or U44700 (N_44700,N_44155,N_44284);
xor U44701 (N_44701,N_44303,N_44319);
and U44702 (N_44702,N_44406,N_44135);
or U44703 (N_44703,N_44067,N_44151);
nor U44704 (N_44704,N_44431,N_44443);
or U44705 (N_44705,N_44326,N_44110);
nand U44706 (N_44706,N_44445,N_44255);
or U44707 (N_44707,N_44332,N_44079);
or U44708 (N_44708,N_44294,N_44225);
xor U44709 (N_44709,N_44070,N_44418);
xnor U44710 (N_44710,N_44277,N_44432);
or U44711 (N_44711,N_44203,N_44076);
and U44712 (N_44712,N_44214,N_44081);
and U44713 (N_44713,N_44323,N_44320);
or U44714 (N_44714,N_44171,N_44388);
and U44715 (N_44715,N_44120,N_44457);
nand U44716 (N_44716,N_44213,N_44046);
nor U44717 (N_44717,N_44215,N_44442);
nor U44718 (N_44718,N_44185,N_44006);
nand U44719 (N_44719,N_44429,N_44183);
and U44720 (N_44720,N_44417,N_44189);
xnor U44721 (N_44721,N_44012,N_44029);
xor U44722 (N_44722,N_44489,N_44020);
xor U44723 (N_44723,N_44246,N_44031);
or U44724 (N_44724,N_44083,N_44331);
xnor U44725 (N_44725,N_44484,N_44117);
nand U44726 (N_44726,N_44451,N_44349);
xor U44727 (N_44727,N_44346,N_44259);
nor U44728 (N_44728,N_44342,N_44348);
xor U44729 (N_44729,N_44450,N_44311);
and U44730 (N_44730,N_44485,N_44032);
nand U44731 (N_44731,N_44235,N_44236);
xnor U44732 (N_44732,N_44446,N_44367);
or U44733 (N_44733,N_44125,N_44302);
or U44734 (N_44734,N_44270,N_44279);
xnor U44735 (N_44735,N_44041,N_44324);
xor U44736 (N_44736,N_44106,N_44005);
and U44737 (N_44737,N_44305,N_44127);
or U44738 (N_44738,N_44226,N_44124);
nor U44739 (N_44739,N_44169,N_44052);
nand U44740 (N_44740,N_44363,N_44051);
nor U44741 (N_44741,N_44121,N_44066);
and U44742 (N_44742,N_44427,N_44472);
xor U44743 (N_44743,N_44400,N_44460);
xnor U44744 (N_44744,N_44190,N_44488);
and U44745 (N_44745,N_44068,N_44238);
xnor U44746 (N_44746,N_44166,N_44338);
nor U44747 (N_44747,N_44455,N_44407);
and U44748 (N_44748,N_44372,N_44232);
nor U44749 (N_44749,N_44058,N_44038);
or U44750 (N_44750,N_44250,N_44409);
and U44751 (N_44751,N_44074,N_44045);
or U44752 (N_44752,N_44301,N_44208);
xnor U44753 (N_44753,N_44142,N_44163);
and U44754 (N_44754,N_44492,N_44302);
and U44755 (N_44755,N_44003,N_44441);
nand U44756 (N_44756,N_44355,N_44346);
or U44757 (N_44757,N_44456,N_44250);
xor U44758 (N_44758,N_44329,N_44315);
and U44759 (N_44759,N_44398,N_44414);
nand U44760 (N_44760,N_44180,N_44151);
xor U44761 (N_44761,N_44133,N_44299);
or U44762 (N_44762,N_44420,N_44047);
nand U44763 (N_44763,N_44450,N_44178);
and U44764 (N_44764,N_44313,N_44379);
nor U44765 (N_44765,N_44014,N_44106);
and U44766 (N_44766,N_44073,N_44244);
and U44767 (N_44767,N_44462,N_44067);
and U44768 (N_44768,N_44386,N_44405);
and U44769 (N_44769,N_44174,N_44055);
and U44770 (N_44770,N_44484,N_44287);
nand U44771 (N_44771,N_44426,N_44249);
or U44772 (N_44772,N_44026,N_44475);
and U44773 (N_44773,N_44434,N_44124);
and U44774 (N_44774,N_44219,N_44178);
nor U44775 (N_44775,N_44462,N_44053);
or U44776 (N_44776,N_44043,N_44385);
nand U44777 (N_44777,N_44177,N_44269);
nand U44778 (N_44778,N_44423,N_44141);
nor U44779 (N_44779,N_44493,N_44433);
nor U44780 (N_44780,N_44331,N_44260);
nand U44781 (N_44781,N_44048,N_44234);
and U44782 (N_44782,N_44274,N_44192);
nand U44783 (N_44783,N_44089,N_44337);
xnor U44784 (N_44784,N_44031,N_44111);
or U44785 (N_44785,N_44303,N_44156);
and U44786 (N_44786,N_44367,N_44313);
nor U44787 (N_44787,N_44469,N_44362);
and U44788 (N_44788,N_44410,N_44163);
xor U44789 (N_44789,N_44352,N_44342);
or U44790 (N_44790,N_44033,N_44213);
nor U44791 (N_44791,N_44207,N_44322);
nor U44792 (N_44792,N_44321,N_44174);
nand U44793 (N_44793,N_44076,N_44349);
nand U44794 (N_44794,N_44007,N_44057);
nor U44795 (N_44795,N_44243,N_44107);
or U44796 (N_44796,N_44152,N_44153);
nand U44797 (N_44797,N_44294,N_44244);
xor U44798 (N_44798,N_44194,N_44417);
and U44799 (N_44799,N_44421,N_44303);
and U44800 (N_44800,N_44103,N_44064);
or U44801 (N_44801,N_44362,N_44196);
and U44802 (N_44802,N_44224,N_44434);
or U44803 (N_44803,N_44392,N_44373);
or U44804 (N_44804,N_44223,N_44066);
and U44805 (N_44805,N_44342,N_44129);
or U44806 (N_44806,N_44011,N_44457);
or U44807 (N_44807,N_44056,N_44140);
nor U44808 (N_44808,N_44170,N_44094);
nand U44809 (N_44809,N_44412,N_44164);
nor U44810 (N_44810,N_44159,N_44129);
and U44811 (N_44811,N_44270,N_44376);
or U44812 (N_44812,N_44457,N_44445);
and U44813 (N_44813,N_44245,N_44124);
and U44814 (N_44814,N_44155,N_44403);
and U44815 (N_44815,N_44262,N_44272);
nand U44816 (N_44816,N_44258,N_44313);
and U44817 (N_44817,N_44083,N_44082);
nor U44818 (N_44818,N_44161,N_44462);
or U44819 (N_44819,N_44042,N_44429);
or U44820 (N_44820,N_44341,N_44034);
xor U44821 (N_44821,N_44231,N_44445);
nor U44822 (N_44822,N_44269,N_44333);
and U44823 (N_44823,N_44006,N_44111);
or U44824 (N_44824,N_44055,N_44203);
nand U44825 (N_44825,N_44112,N_44231);
xnor U44826 (N_44826,N_44082,N_44296);
and U44827 (N_44827,N_44153,N_44365);
or U44828 (N_44828,N_44111,N_44049);
nor U44829 (N_44829,N_44495,N_44466);
nor U44830 (N_44830,N_44402,N_44315);
xor U44831 (N_44831,N_44017,N_44461);
nor U44832 (N_44832,N_44442,N_44269);
or U44833 (N_44833,N_44245,N_44165);
and U44834 (N_44834,N_44039,N_44465);
xor U44835 (N_44835,N_44300,N_44378);
xor U44836 (N_44836,N_44056,N_44237);
xnor U44837 (N_44837,N_44175,N_44015);
and U44838 (N_44838,N_44201,N_44398);
xnor U44839 (N_44839,N_44450,N_44258);
nor U44840 (N_44840,N_44171,N_44000);
xor U44841 (N_44841,N_44307,N_44202);
and U44842 (N_44842,N_44017,N_44023);
nand U44843 (N_44843,N_44146,N_44001);
and U44844 (N_44844,N_44296,N_44096);
nor U44845 (N_44845,N_44364,N_44325);
xor U44846 (N_44846,N_44304,N_44490);
xnor U44847 (N_44847,N_44428,N_44327);
nor U44848 (N_44848,N_44128,N_44278);
xor U44849 (N_44849,N_44485,N_44025);
or U44850 (N_44850,N_44420,N_44022);
nor U44851 (N_44851,N_44153,N_44282);
xnor U44852 (N_44852,N_44053,N_44378);
xnor U44853 (N_44853,N_44314,N_44170);
or U44854 (N_44854,N_44087,N_44163);
nor U44855 (N_44855,N_44317,N_44374);
xor U44856 (N_44856,N_44232,N_44248);
and U44857 (N_44857,N_44280,N_44101);
and U44858 (N_44858,N_44261,N_44011);
xnor U44859 (N_44859,N_44049,N_44420);
xor U44860 (N_44860,N_44142,N_44268);
nor U44861 (N_44861,N_44072,N_44190);
and U44862 (N_44862,N_44119,N_44266);
or U44863 (N_44863,N_44493,N_44307);
nand U44864 (N_44864,N_44050,N_44302);
and U44865 (N_44865,N_44472,N_44268);
xor U44866 (N_44866,N_44039,N_44239);
and U44867 (N_44867,N_44360,N_44029);
nor U44868 (N_44868,N_44080,N_44123);
and U44869 (N_44869,N_44488,N_44487);
nor U44870 (N_44870,N_44134,N_44460);
or U44871 (N_44871,N_44214,N_44037);
and U44872 (N_44872,N_44007,N_44047);
or U44873 (N_44873,N_44381,N_44213);
and U44874 (N_44874,N_44179,N_44384);
xor U44875 (N_44875,N_44348,N_44433);
and U44876 (N_44876,N_44344,N_44172);
or U44877 (N_44877,N_44429,N_44174);
and U44878 (N_44878,N_44263,N_44061);
nor U44879 (N_44879,N_44068,N_44203);
xnor U44880 (N_44880,N_44363,N_44182);
nand U44881 (N_44881,N_44223,N_44157);
nand U44882 (N_44882,N_44473,N_44209);
nand U44883 (N_44883,N_44398,N_44193);
nand U44884 (N_44884,N_44360,N_44355);
nor U44885 (N_44885,N_44366,N_44341);
xor U44886 (N_44886,N_44439,N_44289);
or U44887 (N_44887,N_44169,N_44249);
xor U44888 (N_44888,N_44068,N_44429);
and U44889 (N_44889,N_44144,N_44088);
nor U44890 (N_44890,N_44110,N_44426);
nand U44891 (N_44891,N_44118,N_44247);
or U44892 (N_44892,N_44491,N_44442);
nor U44893 (N_44893,N_44291,N_44312);
xor U44894 (N_44894,N_44175,N_44211);
nor U44895 (N_44895,N_44052,N_44291);
nor U44896 (N_44896,N_44113,N_44037);
or U44897 (N_44897,N_44492,N_44420);
or U44898 (N_44898,N_44415,N_44039);
xor U44899 (N_44899,N_44296,N_44269);
or U44900 (N_44900,N_44323,N_44406);
xor U44901 (N_44901,N_44230,N_44371);
or U44902 (N_44902,N_44086,N_44167);
nor U44903 (N_44903,N_44107,N_44411);
nand U44904 (N_44904,N_44198,N_44002);
nand U44905 (N_44905,N_44440,N_44054);
or U44906 (N_44906,N_44211,N_44361);
and U44907 (N_44907,N_44457,N_44340);
nor U44908 (N_44908,N_44211,N_44024);
xor U44909 (N_44909,N_44355,N_44332);
xnor U44910 (N_44910,N_44238,N_44428);
and U44911 (N_44911,N_44008,N_44493);
xor U44912 (N_44912,N_44439,N_44181);
nor U44913 (N_44913,N_44008,N_44362);
and U44914 (N_44914,N_44124,N_44407);
and U44915 (N_44915,N_44040,N_44342);
nand U44916 (N_44916,N_44368,N_44460);
xor U44917 (N_44917,N_44219,N_44284);
nand U44918 (N_44918,N_44320,N_44070);
and U44919 (N_44919,N_44410,N_44011);
nand U44920 (N_44920,N_44186,N_44031);
xnor U44921 (N_44921,N_44455,N_44418);
nor U44922 (N_44922,N_44073,N_44001);
or U44923 (N_44923,N_44249,N_44168);
nand U44924 (N_44924,N_44191,N_44261);
xnor U44925 (N_44925,N_44036,N_44249);
and U44926 (N_44926,N_44232,N_44027);
nor U44927 (N_44927,N_44322,N_44434);
xor U44928 (N_44928,N_44090,N_44245);
and U44929 (N_44929,N_44419,N_44385);
nor U44930 (N_44930,N_44456,N_44227);
and U44931 (N_44931,N_44189,N_44161);
nor U44932 (N_44932,N_44346,N_44225);
or U44933 (N_44933,N_44211,N_44213);
nor U44934 (N_44934,N_44374,N_44088);
xnor U44935 (N_44935,N_44088,N_44196);
nor U44936 (N_44936,N_44229,N_44114);
xor U44937 (N_44937,N_44180,N_44345);
or U44938 (N_44938,N_44473,N_44249);
or U44939 (N_44939,N_44324,N_44132);
or U44940 (N_44940,N_44235,N_44420);
nor U44941 (N_44941,N_44307,N_44061);
nor U44942 (N_44942,N_44113,N_44447);
or U44943 (N_44943,N_44106,N_44329);
and U44944 (N_44944,N_44214,N_44134);
or U44945 (N_44945,N_44407,N_44377);
nor U44946 (N_44946,N_44203,N_44119);
xor U44947 (N_44947,N_44128,N_44150);
nand U44948 (N_44948,N_44349,N_44334);
nand U44949 (N_44949,N_44388,N_44284);
and U44950 (N_44950,N_44302,N_44087);
and U44951 (N_44951,N_44121,N_44141);
or U44952 (N_44952,N_44423,N_44013);
or U44953 (N_44953,N_44130,N_44338);
nand U44954 (N_44954,N_44423,N_44384);
nand U44955 (N_44955,N_44345,N_44375);
or U44956 (N_44956,N_44168,N_44354);
or U44957 (N_44957,N_44401,N_44478);
xor U44958 (N_44958,N_44021,N_44047);
nor U44959 (N_44959,N_44427,N_44460);
nor U44960 (N_44960,N_44240,N_44043);
nor U44961 (N_44961,N_44241,N_44129);
and U44962 (N_44962,N_44421,N_44210);
and U44963 (N_44963,N_44352,N_44461);
or U44964 (N_44964,N_44303,N_44121);
nand U44965 (N_44965,N_44404,N_44152);
nand U44966 (N_44966,N_44275,N_44107);
and U44967 (N_44967,N_44003,N_44079);
or U44968 (N_44968,N_44329,N_44031);
xnor U44969 (N_44969,N_44015,N_44062);
nand U44970 (N_44970,N_44436,N_44059);
and U44971 (N_44971,N_44216,N_44397);
nor U44972 (N_44972,N_44480,N_44459);
nor U44973 (N_44973,N_44045,N_44368);
nor U44974 (N_44974,N_44172,N_44389);
nand U44975 (N_44975,N_44394,N_44038);
nand U44976 (N_44976,N_44125,N_44299);
nand U44977 (N_44977,N_44297,N_44455);
or U44978 (N_44978,N_44227,N_44053);
and U44979 (N_44979,N_44278,N_44184);
nor U44980 (N_44980,N_44146,N_44088);
nand U44981 (N_44981,N_44052,N_44084);
xnor U44982 (N_44982,N_44283,N_44086);
nor U44983 (N_44983,N_44099,N_44342);
and U44984 (N_44984,N_44210,N_44063);
and U44985 (N_44985,N_44488,N_44325);
and U44986 (N_44986,N_44039,N_44261);
xor U44987 (N_44987,N_44243,N_44486);
xnor U44988 (N_44988,N_44210,N_44285);
xor U44989 (N_44989,N_44235,N_44034);
and U44990 (N_44990,N_44316,N_44322);
or U44991 (N_44991,N_44250,N_44147);
nand U44992 (N_44992,N_44093,N_44475);
or U44993 (N_44993,N_44436,N_44427);
nor U44994 (N_44994,N_44006,N_44329);
and U44995 (N_44995,N_44205,N_44079);
or U44996 (N_44996,N_44221,N_44199);
nand U44997 (N_44997,N_44101,N_44138);
and U44998 (N_44998,N_44303,N_44104);
xnor U44999 (N_44999,N_44165,N_44054);
nand U45000 (N_45000,N_44929,N_44669);
or U45001 (N_45001,N_44838,N_44877);
and U45002 (N_45002,N_44664,N_44813);
nor U45003 (N_45003,N_44662,N_44953);
nand U45004 (N_45004,N_44733,N_44609);
or U45005 (N_45005,N_44831,N_44699);
or U45006 (N_45006,N_44907,N_44864);
and U45007 (N_45007,N_44668,N_44741);
nand U45008 (N_45008,N_44819,N_44671);
and U45009 (N_45009,N_44695,N_44684);
and U45010 (N_45010,N_44646,N_44795);
and U45011 (N_45011,N_44944,N_44634);
and U45012 (N_45012,N_44899,N_44557);
or U45013 (N_45013,N_44886,N_44502);
and U45014 (N_45014,N_44517,N_44859);
xor U45015 (N_45015,N_44670,N_44627);
or U45016 (N_45016,N_44617,N_44694);
nor U45017 (N_45017,N_44587,N_44564);
and U45018 (N_45018,N_44576,N_44784);
or U45019 (N_45019,N_44853,N_44606);
and U45020 (N_45020,N_44769,N_44940);
or U45021 (N_45021,N_44704,N_44541);
nor U45022 (N_45022,N_44901,N_44780);
or U45023 (N_45023,N_44559,N_44661);
nand U45024 (N_45024,N_44975,N_44807);
or U45025 (N_45025,N_44536,N_44880);
and U45026 (N_45026,N_44928,N_44696);
nand U45027 (N_45027,N_44991,N_44958);
xnor U45028 (N_45028,N_44895,N_44526);
or U45029 (N_45029,N_44650,N_44777);
or U45030 (N_45030,N_44628,N_44547);
nand U45031 (N_45031,N_44837,N_44791);
nor U45032 (N_45032,N_44803,N_44505);
xnor U45033 (N_45033,N_44774,N_44535);
or U45034 (N_45034,N_44866,N_44654);
and U45035 (N_45035,N_44821,N_44832);
or U45036 (N_45036,N_44910,N_44569);
xnor U45037 (N_45037,N_44677,N_44989);
and U45038 (N_45038,N_44960,N_44705);
nor U45039 (N_45039,N_44739,N_44501);
xnor U45040 (N_45040,N_44922,N_44625);
and U45041 (N_45041,N_44720,N_44924);
and U45042 (N_45042,N_44916,N_44714);
nand U45043 (N_45043,N_44852,N_44596);
nor U45044 (N_45044,N_44726,N_44568);
and U45045 (N_45045,N_44851,N_44939);
xor U45046 (N_45046,N_44787,N_44630);
or U45047 (N_45047,N_44912,N_44512);
xnor U45048 (N_45048,N_44950,N_44845);
or U45049 (N_45049,N_44996,N_44843);
and U45050 (N_45050,N_44841,N_44760);
nand U45051 (N_45051,N_44583,N_44666);
or U45052 (N_45052,N_44629,N_44794);
nor U45053 (N_45053,N_44834,N_44827);
nor U45054 (N_45054,N_44632,N_44826);
nand U45055 (N_45055,N_44767,N_44667);
or U45056 (N_45056,N_44915,N_44936);
or U45057 (N_45057,N_44847,N_44633);
xnor U45058 (N_45058,N_44624,N_44812);
nand U45059 (N_45059,N_44799,N_44875);
nor U45060 (N_45060,N_44570,N_44572);
nand U45061 (N_45061,N_44607,N_44722);
and U45062 (N_45062,N_44678,N_44893);
nor U45063 (N_45063,N_44676,N_44649);
xnor U45064 (N_45064,N_44923,N_44555);
nor U45065 (N_45065,N_44801,N_44959);
or U45066 (N_45066,N_44525,N_44833);
or U45067 (N_45067,N_44779,N_44626);
nor U45068 (N_45068,N_44729,N_44565);
nor U45069 (N_45069,N_44605,N_44946);
and U45070 (N_45070,N_44721,N_44644);
xor U45071 (N_45071,N_44882,N_44603);
and U45072 (N_45072,N_44898,N_44824);
nor U45073 (N_45073,N_44942,N_44804);
nor U45074 (N_45074,N_44746,N_44692);
nor U45075 (N_45075,N_44917,N_44580);
nor U45076 (N_45076,N_44796,N_44690);
nand U45077 (N_45077,N_44905,N_44506);
and U45078 (N_45078,N_44839,N_44658);
nor U45079 (N_45079,N_44691,N_44884);
nand U45080 (N_45080,N_44542,N_44885);
nand U45081 (N_45081,N_44503,N_44793);
and U45082 (N_45082,N_44823,N_44814);
nand U45083 (N_45083,N_44653,N_44969);
nand U45084 (N_45084,N_44848,N_44518);
nand U45085 (N_45085,N_44749,N_44703);
nor U45086 (N_45086,N_44934,N_44665);
nor U45087 (N_45087,N_44992,N_44577);
and U45088 (N_45088,N_44556,N_44763);
or U45089 (N_45089,N_44752,N_44595);
and U45090 (N_45090,N_44655,N_44520);
and U45091 (N_45091,N_44900,N_44904);
or U45092 (N_45092,N_44613,N_44510);
nor U45093 (N_45093,N_44938,N_44598);
or U45094 (N_45094,N_44717,N_44636);
xnor U45095 (N_45095,N_44840,N_44945);
nand U45096 (N_45096,N_44710,N_44527);
nand U45097 (N_45097,N_44957,N_44941);
or U45098 (N_45098,N_44964,N_44600);
xor U45099 (N_45099,N_44623,N_44849);
nor U45100 (N_45100,N_44894,N_44718);
xor U45101 (N_45101,N_44802,N_44775);
nor U45102 (N_45102,N_44528,N_44659);
xnor U45103 (N_45103,N_44750,N_44782);
and U45104 (N_45104,N_44903,N_44687);
or U45105 (N_45105,N_44748,N_44762);
nor U45106 (N_45106,N_44619,N_44810);
nand U45107 (N_45107,N_44640,N_44601);
nand U45108 (N_45108,N_44701,N_44708);
xnor U45109 (N_45109,N_44973,N_44551);
nand U45110 (N_45110,N_44645,N_44867);
nand U45111 (N_45111,N_44735,N_44514);
or U45112 (N_45112,N_44642,N_44567);
and U45113 (N_45113,N_44571,N_44612);
nor U45114 (N_45114,N_44835,N_44713);
nand U45115 (N_45115,N_44682,N_44737);
nor U45116 (N_45116,N_44967,N_44756);
xnor U45117 (N_45117,N_44611,N_44906);
xor U45118 (N_45118,N_44971,N_44783);
or U45119 (N_45119,N_44686,N_44995);
nand U45120 (N_45120,N_44742,N_44816);
nor U45121 (N_45121,N_44730,N_44956);
nor U45122 (N_45122,N_44672,N_44902);
nand U45123 (N_45123,N_44546,N_44772);
nand U45124 (N_45124,N_44549,N_44727);
nand U45125 (N_45125,N_44778,N_44872);
and U45126 (N_45126,N_44863,N_44978);
or U45127 (N_45127,N_44738,N_44757);
or U45128 (N_45128,N_44681,N_44652);
or U45129 (N_45129,N_44519,N_44736);
and U45130 (N_45130,N_44862,N_44543);
and U45131 (N_45131,N_44637,N_44508);
or U45132 (N_45132,N_44651,N_44643);
or U45133 (N_45133,N_44965,N_44604);
or U45134 (N_45134,N_44954,N_44981);
nor U45135 (N_45135,N_44798,N_44500);
nor U45136 (N_45136,N_44822,N_44610);
xnor U45137 (N_45137,N_44999,N_44548);
nor U45138 (N_45138,N_44788,N_44707);
or U45139 (N_45139,N_44639,N_44581);
nand U45140 (N_45140,N_44908,N_44800);
or U45141 (N_45141,N_44562,N_44868);
nor U45142 (N_45142,N_44589,N_44920);
nand U45143 (N_45143,N_44766,N_44693);
nand U45144 (N_45144,N_44573,N_44952);
xor U45145 (N_45145,N_44702,N_44584);
and U45146 (N_45146,N_44968,N_44776);
and U45147 (N_45147,N_44511,N_44516);
and U45148 (N_45148,N_44734,N_44685);
or U45149 (N_45149,N_44984,N_44926);
nand U45150 (N_45150,N_44558,N_44860);
and U45151 (N_45151,N_44948,N_44574);
nand U45152 (N_45152,N_44594,N_44770);
or U45153 (N_45153,N_44909,N_44648);
nor U45154 (N_45154,N_44871,N_44919);
and U45155 (N_45155,N_44550,N_44997);
nor U45156 (N_45156,N_44879,N_44876);
xnor U45157 (N_45157,N_44986,N_44943);
xnor U45158 (N_45158,N_44870,N_44855);
xor U45159 (N_45159,N_44622,N_44673);
or U45160 (N_45160,N_44680,N_44933);
or U45161 (N_45161,N_44888,N_44951);
nand U45162 (N_45162,N_44647,N_44590);
or U45163 (N_45163,N_44635,N_44828);
nor U45164 (N_45164,N_44615,N_44931);
nor U45165 (N_45165,N_44723,N_44990);
xor U45166 (N_45166,N_44771,N_44533);
nand U45167 (N_45167,N_44744,N_44523);
xnor U45168 (N_45168,N_44621,N_44854);
nor U45169 (N_45169,N_44585,N_44544);
nor U45170 (N_45170,N_44540,N_44842);
nand U45171 (N_45171,N_44972,N_44679);
nor U45172 (N_45172,N_44809,N_44728);
or U45173 (N_45173,N_44789,N_44918);
xor U45174 (N_45174,N_44874,N_44856);
nor U45175 (N_45175,N_44561,N_44731);
and U45176 (N_45176,N_44808,N_44980);
or U45177 (N_45177,N_44698,N_44553);
nand U45178 (N_45178,N_44790,N_44993);
nand U45179 (N_45179,N_44873,N_44925);
and U45180 (N_45180,N_44732,N_44579);
and U45181 (N_45181,N_44921,N_44883);
xnor U45182 (N_45182,N_44712,N_44785);
or U45183 (N_45183,N_44881,N_44534);
or U45184 (N_45184,N_44554,N_44560);
nand U45185 (N_45185,N_44811,N_44599);
nor U45186 (N_45186,N_44751,N_44985);
and U45187 (N_45187,N_44675,N_44753);
nand U45188 (N_45188,N_44608,N_44869);
nand U45189 (N_45189,N_44586,N_44724);
and U45190 (N_45190,N_44697,N_44932);
and U45191 (N_45191,N_44578,N_44937);
or U45192 (N_45192,N_44522,N_44955);
nand U45193 (N_45193,N_44805,N_44660);
nand U45194 (N_45194,N_44592,N_44935);
nand U45195 (N_45195,N_44552,N_44844);
xnor U45196 (N_45196,N_44575,N_44988);
nor U45197 (N_45197,N_44887,N_44889);
nor U45198 (N_45198,N_44689,N_44892);
xnor U45199 (N_45199,N_44982,N_44979);
nor U45200 (N_45200,N_44850,N_44591);
xnor U45201 (N_45201,N_44878,N_44758);
xnor U45202 (N_45202,N_44706,N_44754);
or U45203 (N_45203,N_44861,N_44961);
xor U45204 (N_45204,N_44588,N_44768);
xnor U45205 (N_45205,N_44836,N_44820);
and U45206 (N_45206,N_44829,N_44566);
and U45207 (N_45207,N_44891,N_44846);
nor U45208 (N_45208,N_44970,N_44530);
xor U45209 (N_45209,N_44927,N_44759);
xor U45210 (N_45210,N_44674,N_44515);
xor U45211 (N_45211,N_44817,N_44781);
or U45212 (N_45212,N_44582,N_44509);
and U45213 (N_45213,N_44529,N_44911);
or U45214 (N_45214,N_44865,N_44597);
xnor U45215 (N_45215,N_44593,N_44896);
nor U45216 (N_45216,N_44963,N_44761);
nor U45217 (N_45217,N_44620,N_44715);
or U45218 (N_45218,N_44815,N_44743);
and U45219 (N_45219,N_44719,N_44531);
or U45220 (N_45220,N_44857,N_44657);
nand U45221 (N_45221,N_44792,N_44976);
and U45222 (N_45222,N_44858,N_44700);
and U45223 (N_45223,N_44641,N_44998);
and U45224 (N_45224,N_44962,N_44797);
or U45225 (N_45225,N_44618,N_44524);
nand U45226 (N_45226,N_44983,N_44537);
or U45227 (N_45227,N_44773,N_44977);
xnor U45228 (N_45228,N_44974,N_44538);
or U45229 (N_45229,N_44806,N_44890);
nor U45230 (N_45230,N_44521,N_44616);
nor U45231 (N_45231,N_44947,N_44545);
and U45232 (N_45232,N_44914,N_44764);
xnor U45233 (N_45233,N_44507,N_44539);
nand U45234 (N_45234,N_44716,N_44949);
or U45235 (N_45235,N_44725,N_44755);
or U45236 (N_45236,N_44966,N_44663);
xor U45237 (N_45237,N_44638,N_44818);
and U45238 (N_45238,N_44504,N_44747);
xor U45239 (N_45239,N_44745,N_44897);
nor U45240 (N_45240,N_44765,N_44709);
or U45241 (N_45241,N_44830,N_44688);
nand U45242 (N_45242,N_44740,N_44532);
nor U45243 (N_45243,N_44994,N_44930);
nand U45244 (N_45244,N_44656,N_44683);
nand U45245 (N_45245,N_44614,N_44602);
nand U45246 (N_45246,N_44987,N_44563);
xor U45247 (N_45247,N_44786,N_44631);
and U45248 (N_45248,N_44513,N_44711);
nor U45249 (N_45249,N_44913,N_44825);
or U45250 (N_45250,N_44572,N_44745);
and U45251 (N_45251,N_44560,N_44711);
or U45252 (N_45252,N_44850,N_44578);
xnor U45253 (N_45253,N_44503,N_44507);
xor U45254 (N_45254,N_44814,N_44903);
nor U45255 (N_45255,N_44903,N_44690);
nor U45256 (N_45256,N_44601,N_44756);
and U45257 (N_45257,N_44792,N_44577);
nand U45258 (N_45258,N_44736,N_44506);
or U45259 (N_45259,N_44956,N_44862);
nor U45260 (N_45260,N_44840,N_44768);
and U45261 (N_45261,N_44778,N_44902);
or U45262 (N_45262,N_44517,N_44950);
nand U45263 (N_45263,N_44537,N_44743);
and U45264 (N_45264,N_44780,N_44783);
or U45265 (N_45265,N_44635,N_44917);
nor U45266 (N_45266,N_44713,N_44730);
xor U45267 (N_45267,N_44980,N_44554);
nor U45268 (N_45268,N_44578,N_44965);
nand U45269 (N_45269,N_44504,N_44764);
xnor U45270 (N_45270,N_44902,N_44770);
nor U45271 (N_45271,N_44650,N_44960);
and U45272 (N_45272,N_44552,N_44656);
and U45273 (N_45273,N_44671,N_44977);
nor U45274 (N_45274,N_44998,N_44937);
or U45275 (N_45275,N_44604,N_44513);
nor U45276 (N_45276,N_44810,N_44610);
nor U45277 (N_45277,N_44668,N_44832);
nand U45278 (N_45278,N_44726,N_44640);
or U45279 (N_45279,N_44558,N_44544);
and U45280 (N_45280,N_44854,N_44997);
xor U45281 (N_45281,N_44552,N_44503);
nand U45282 (N_45282,N_44952,N_44690);
nand U45283 (N_45283,N_44758,N_44679);
or U45284 (N_45284,N_44603,N_44881);
nor U45285 (N_45285,N_44671,N_44603);
nor U45286 (N_45286,N_44869,N_44635);
xor U45287 (N_45287,N_44876,N_44595);
nand U45288 (N_45288,N_44529,N_44890);
nand U45289 (N_45289,N_44549,N_44818);
nand U45290 (N_45290,N_44652,N_44573);
nand U45291 (N_45291,N_44698,N_44569);
xor U45292 (N_45292,N_44778,N_44866);
nand U45293 (N_45293,N_44893,N_44510);
nand U45294 (N_45294,N_44711,N_44585);
nor U45295 (N_45295,N_44853,N_44558);
nand U45296 (N_45296,N_44636,N_44978);
nor U45297 (N_45297,N_44886,N_44597);
nor U45298 (N_45298,N_44627,N_44973);
nand U45299 (N_45299,N_44759,N_44982);
nand U45300 (N_45300,N_44614,N_44587);
or U45301 (N_45301,N_44783,N_44837);
nor U45302 (N_45302,N_44911,N_44746);
nand U45303 (N_45303,N_44962,N_44710);
xnor U45304 (N_45304,N_44779,N_44826);
xnor U45305 (N_45305,N_44821,N_44535);
xnor U45306 (N_45306,N_44504,N_44925);
xnor U45307 (N_45307,N_44622,N_44631);
xnor U45308 (N_45308,N_44804,N_44654);
nor U45309 (N_45309,N_44505,N_44677);
or U45310 (N_45310,N_44584,N_44540);
xor U45311 (N_45311,N_44755,N_44685);
nor U45312 (N_45312,N_44862,N_44975);
or U45313 (N_45313,N_44896,N_44903);
nor U45314 (N_45314,N_44958,N_44581);
xor U45315 (N_45315,N_44502,N_44827);
and U45316 (N_45316,N_44529,N_44917);
nor U45317 (N_45317,N_44915,N_44798);
and U45318 (N_45318,N_44804,N_44985);
xnor U45319 (N_45319,N_44829,N_44738);
nand U45320 (N_45320,N_44781,N_44664);
or U45321 (N_45321,N_44554,N_44753);
nand U45322 (N_45322,N_44625,N_44717);
xnor U45323 (N_45323,N_44610,N_44930);
nor U45324 (N_45324,N_44516,N_44509);
xnor U45325 (N_45325,N_44879,N_44662);
nand U45326 (N_45326,N_44988,N_44952);
or U45327 (N_45327,N_44902,N_44877);
xor U45328 (N_45328,N_44556,N_44735);
xnor U45329 (N_45329,N_44983,N_44538);
and U45330 (N_45330,N_44517,N_44708);
nor U45331 (N_45331,N_44985,N_44508);
or U45332 (N_45332,N_44938,N_44567);
nand U45333 (N_45333,N_44865,N_44788);
nor U45334 (N_45334,N_44727,N_44562);
xor U45335 (N_45335,N_44633,N_44845);
and U45336 (N_45336,N_44844,N_44514);
or U45337 (N_45337,N_44688,N_44554);
or U45338 (N_45338,N_44557,N_44513);
nor U45339 (N_45339,N_44779,N_44646);
and U45340 (N_45340,N_44567,N_44840);
or U45341 (N_45341,N_44529,N_44703);
and U45342 (N_45342,N_44667,N_44974);
and U45343 (N_45343,N_44664,N_44828);
and U45344 (N_45344,N_44766,N_44653);
nand U45345 (N_45345,N_44809,N_44665);
nor U45346 (N_45346,N_44963,N_44740);
nor U45347 (N_45347,N_44784,N_44582);
xnor U45348 (N_45348,N_44857,N_44692);
nand U45349 (N_45349,N_44691,N_44852);
and U45350 (N_45350,N_44561,N_44581);
nand U45351 (N_45351,N_44892,N_44935);
or U45352 (N_45352,N_44538,N_44805);
xnor U45353 (N_45353,N_44506,N_44876);
xnor U45354 (N_45354,N_44771,N_44552);
xnor U45355 (N_45355,N_44563,N_44615);
and U45356 (N_45356,N_44586,N_44756);
xnor U45357 (N_45357,N_44681,N_44710);
nor U45358 (N_45358,N_44909,N_44893);
nor U45359 (N_45359,N_44822,N_44729);
and U45360 (N_45360,N_44876,N_44808);
nor U45361 (N_45361,N_44861,N_44658);
or U45362 (N_45362,N_44978,N_44869);
xor U45363 (N_45363,N_44854,N_44610);
nor U45364 (N_45364,N_44994,N_44700);
nor U45365 (N_45365,N_44634,N_44777);
xnor U45366 (N_45366,N_44511,N_44681);
and U45367 (N_45367,N_44616,N_44856);
nor U45368 (N_45368,N_44828,N_44578);
nor U45369 (N_45369,N_44696,N_44823);
or U45370 (N_45370,N_44615,N_44718);
xor U45371 (N_45371,N_44676,N_44885);
xor U45372 (N_45372,N_44890,N_44834);
and U45373 (N_45373,N_44850,N_44663);
nand U45374 (N_45374,N_44689,N_44886);
and U45375 (N_45375,N_44617,N_44854);
nor U45376 (N_45376,N_44732,N_44823);
nor U45377 (N_45377,N_44711,N_44881);
xor U45378 (N_45378,N_44737,N_44825);
nand U45379 (N_45379,N_44579,N_44934);
nor U45380 (N_45380,N_44569,N_44718);
xnor U45381 (N_45381,N_44777,N_44615);
and U45382 (N_45382,N_44688,N_44952);
and U45383 (N_45383,N_44717,N_44899);
xnor U45384 (N_45384,N_44610,N_44540);
xnor U45385 (N_45385,N_44619,N_44597);
and U45386 (N_45386,N_44872,N_44612);
or U45387 (N_45387,N_44645,N_44707);
nand U45388 (N_45388,N_44935,N_44635);
nand U45389 (N_45389,N_44810,N_44711);
nor U45390 (N_45390,N_44925,N_44577);
nand U45391 (N_45391,N_44542,N_44944);
and U45392 (N_45392,N_44670,N_44927);
xor U45393 (N_45393,N_44912,N_44682);
and U45394 (N_45394,N_44573,N_44963);
xor U45395 (N_45395,N_44539,N_44709);
and U45396 (N_45396,N_44761,N_44648);
nand U45397 (N_45397,N_44763,N_44574);
nor U45398 (N_45398,N_44651,N_44831);
nand U45399 (N_45399,N_44927,N_44900);
and U45400 (N_45400,N_44837,N_44931);
or U45401 (N_45401,N_44842,N_44655);
and U45402 (N_45402,N_44567,N_44524);
or U45403 (N_45403,N_44680,N_44799);
and U45404 (N_45404,N_44632,N_44886);
nor U45405 (N_45405,N_44593,N_44968);
and U45406 (N_45406,N_44902,N_44889);
or U45407 (N_45407,N_44631,N_44726);
nand U45408 (N_45408,N_44686,N_44727);
nand U45409 (N_45409,N_44818,N_44946);
and U45410 (N_45410,N_44569,N_44581);
and U45411 (N_45411,N_44717,N_44712);
or U45412 (N_45412,N_44695,N_44508);
nand U45413 (N_45413,N_44783,N_44863);
xnor U45414 (N_45414,N_44957,N_44765);
nand U45415 (N_45415,N_44819,N_44512);
xnor U45416 (N_45416,N_44661,N_44755);
xor U45417 (N_45417,N_44955,N_44789);
or U45418 (N_45418,N_44619,N_44514);
nand U45419 (N_45419,N_44950,N_44941);
xor U45420 (N_45420,N_44802,N_44647);
and U45421 (N_45421,N_44954,N_44600);
and U45422 (N_45422,N_44929,N_44673);
nand U45423 (N_45423,N_44907,N_44780);
and U45424 (N_45424,N_44950,N_44634);
xnor U45425 (N_45425,N_44758,N_44853);
nor U45426 (N_45426,N_44963,N_44879);
nand U45427 (N_45427,N_44634,N_44545);
nand U45428 (N_45428,N_44690,N_44897);
and U45429 (N_45429,N_44996,N_44915);
and U45430 (N_45430,N_44856,N_44511);
and U45431 (N_45431,N_44878,N_44640);
xnor U45432 (N_45432,N_44510,N_44800);
or U45433 (N_45433,N_44548,N_44876);
and U45434 (N_45434,N_44950,N_44525);
nand U45435 (N_45435,N_44717,N_44731);
and U45436 (N_45436,N_44838,N_44504);
nor U45437 (N_45437,N_44773,N_44575);
and U45438 (N_45438,N_44971,N_44999);
or U45439 (N_45439,N_44688,N_44663);
and U45440 (N_45440,N_44991,N_44903);
xnor U45441 (N_45441,N_44613,N_44891);
and U45442 (N_45442,N_44903,N_44554);
and U45443 (N_45443,N_44524,N_44537);
or U45444 (N_45444,N_44939,N_44635);
xor U45445 (N_45445,N_44975,N_44527);
nor U45446 (N_45446,N_44817,N_44796);
nor U45447 (N_45447,N_44674,N_44995);
nor U45448 (N_45448,N_44992,N_44972);
xor U45449 (N_45449,N_44816,N_44738);
nand U45450 (N_45450,N_44689,N_44982);
or U45451 (N_45451,N_44797,N_44564);
xnor U45452 (N_45452,N_44837,N_44638);
and U45453 (N_45453,N_44687,N_44917);
and U45454 (N_45454,N_44557,N_44864);
and U45455 (N_45455,N_44898,N_44567);
nor U45456 (N_45456,N_44524,N_44549);
nand U45457 (N_45457,N_44910,N_44795);
xnor U45458 (N_45458,N_44895,N_44721);
nand U45459 (N_45459,N_44648,N_44831);
xor U45460 (N_45460,N_44965,N_44810);
nand U45461 (N_45461,N_44662,N_44998);
xor U45462 (N_45462,N_44590,N_44736);
nand U45463 (N_45463,N_44525,N_44864);
and U45464 (N_45464,N_44699,N_44929);
and U45465 (N_45465,N_44777,N_44630);
nand U45466 (N_45466,N_44740,N_44848);
xor U45467 (N_45467,N_44786,N_44699);
or U45468 (N_45468,N_44627,N_44785);
xor U45469 (N_45469,N_44532,N_44508);
xor U45470 (N_45470,N_44779,N_44547);
nand U45471 (N_45471,N_44963,N_44853);
xor U45472 (N_45472,N_44754,N_44620);
nand U45473 (N_45473,N_44519,N_44717);
or U45474 (N_45474,N_44795,N_44689);
xnor U45475 (N_45475,N_44863,N_44574);
nand U45476 (N_45476,N_44514,N_44638);
nand U45477 (N_45477,N_44650,N_44808);
or U45478 (N_45478,N_44934,N_44935);
xor U45479 (N_45479,N_44883,N_44907);
xor U45480 (N_45480,N_44812,N_44684);
nor U45481 (N_45481,N_44988,N_44852);
xnor U45482 (N_45482,N_44937,N_44530);
or U45483 (N_45483,N_44527,N_44704);
and U45484 (N_45484,N_44611,N_44877);
xnor U45485 (N_45485,N_44512,N_44702);
and U45486 (N_45486,N_44614,N_44994);
and U45487 (N_45487,N_44652,N_44696);
or U45488 (N_45488,N_44626,N_44727);
xor U45489 (N_45489,N_44597,N_44605);
or U45490 (N_45490,N_44765,N_44749);
nand U45491 (N_45491,N_44580,N_44723);
xnor U45492 (N_45492,N_44899,N_44645);
nand U45493 (N_45493,N_44791,N_44793);
or U45494 (N_45494,N_44983,N_44806);
and U45495 (N_45495,N_44610,N_44970);
and U45496 (N_45496,N_44723,N_44997);
or U45497 (N_45497,N_44666,N_44631);
xor U45498 (N_45498,N_44633,N_44849);
or U45499 (N_45499,N_44796,N_44679);
nand U45500 (N_45500,N_45090,N_45023);
nor U45501 (N_45501,N_45488,N_45497);
xor U45502 (N_45502,N_45399,N_45462);
or U45503 (N_45503,N_45321,N_45258);
nor U45504 (N_45504,N_45312,N_45133);
or U45505 (N_45505,N_45106,N_45481);
xnor U45506 (N_45506,N_45146,N_45173);
nor U45507 (N_45507,N_45262,N_45078);
or U45508 (N_45508,N_45231,N_45493);
and U45509 (N_45509,N_45408,N_45020);
and U45510 (N_45510,N_45216,N_45077);
and U45511 (N_45511,N_45252,N_45496);
and U45512 (N_45512,N_45355,N_45192);
xor U45513 (N_45513,N_45314,N_45453);
or U45514 (N_45514,N_45119,N_45297);
xor U45515 (N_45515,N_45084,N_45061);
and U45516 (N_45516,N_45148,N_45356);
nand U45517 (N_45517,N_45076,N_45011);
xor U45518 (N_45518,N_45140,N_45016);
or U45519 (N_45519,N_45423,N_45037);
and U45520 (N_45520,N_45160,N_45263);
nor U45521 (N_45521,N_45495,N_45281);
and U45522 (N_45522,N_45058,N_45034);
and U45523 (N_45523,N_45038,N_45449);
or U45524 (N_45524,N_45447,N_45112);
nor U45525 (N_45525,N_45006,N_45253);
and U45526 (N_45526,N_45157,N_45279);
nand U45527 (N_45527,N_45303,N_45190);
or U45528 (N_45528,N_45256,N_45284);
nand U45529 (N_45529,N_45341,N_45494);
nor U45530 (N_45530,N_45468,N_45144);
and U45531 (N_45531,N_45407,N_45487);
nand U45532 (N_45532,N_45396,N_45089);
or U45533 (N_45533,N_45461,N_45477);
nor U45534 (N_45534,N_45232,N_45154);
nand U45535 (N_45535,N_45002,N_45062);
xor U45536 (N_45536,N_45003,N_45234);
and U45537 (N_45537,N_45376,N_45042);
nand U45538 (N_45538,N_45437,N_45053);
and U45539 (N_45539,N_45172,N_45325);
xnor U45540 (N_45540,N_45385,N_45414);
xnor U45541 (N_45541,N_45442,N_45390);
nand U45542 (N_45542,N_45358,N_45127);
or U45543 (N_45543,N_45250,N_45309);
nor U45544 (N_45544,N_45413,N_45130);
or U45545 (N_45545,N_45125,N_45268);
xor U45546 (N_45546,N_45116,N_45412);
or U45547 (N_45547,N_45165,N_45168);
nor U45548 (N_45548,N_45159,N_45240);
or U45549 (N_45549,N_45107,N_45417);
or U45550 (N_45550,N_45402,N_45350);
nor U45551 (N_45551,N_45397,N_45083);
and U45552 (N_45552,N_45179,N_45409);
xor U45553 (N_45553,N_45132,N_45451);
or U45554 (N_45554,N_45180,N_45340);
or U45555 (N_45555,N_45415,N_45093);
and U45556 (N_45556,N_45104,N_45181);
or U45557 (N_45557,N_45043,N_45217);
and U45558 (N_45558,N_45259,N_45270);
nand U45559 (N_45559,N_45237,N_45117);
xor U45560 (N_45560,N_45290,N_45474);
or U45561 (N_45561,N_45103,N_45406);
nor U45562 (N_45562,N_45118,N_45212);
or U45563 (N_45563,N_45433,N_45087);
xnor U45564 (N_45564,N_45227,N_45244);
and U45565 (N_45565,N_45029,N_45334);
or U45566 (N_45566,N_45137,N_45289);
and U45567 (N_45567,N_45342,N_45299);
nand U45568 (N_45568,N_45004,N_45100);
xnor U45569 (N_45569,N_45143,N_45211);
or U45570 (N_45570,N_45219,N_45033);
and U45571 (N_45571,N_45072,N_45419);
and U45572 (N_45572,N_45193,N_45378);
or U45573 (N_45573,N_45114,N_45277);
nor U45574 (N_45574,N_45222,N_45007);
or U45575 (N_45575,N_45113,N_45470);
xor U45576 (N_45576,N_45275,N_45400);
xor U45577 (N_45577,N_45138,N_45257);
nor U45578 (N_45578,N_45201,N_45265);
and U45579 (N_45579,N_45241,N_45464);
or U45580 (N_45580,N_45318,N_45288);
and U45581 (N_45581,N_45455,N_45282);
xnor U45582 (N_45582,N_45060,N_45096);
xnor U45583 (N_45583,N_45392,N_45105);
nor U45584 (N_45584,N_45164,N_45291);
nor U45585 (N_45585,N_45071,N_45028);
or U45586 (N_45586,N_45178,N_45074);
nand U45587 (N_45587,N_45373,N_45343);
and U45588 (N_45588,N_45047,N_45088);
and U45589 (N_45589,N_45266,N_45264);
nand U45590 (N_45590,N_45332,N_45436);
or U45591 (N_45591,N_45422,N_45218);
nand U45592 (N_45592,N_45441,N_45388);
or U45593 (N_45593,N_45195,N_45050);
and U45594 (N_45594,N_45484,N_45425);
or U45595 (N_45595,N_45131,N_45018);
or U45596 (N_45596,N_45324,N_45359);
nand U45597 (N_45597,N_45121,N_45432);
or U45598 (N_45598,N_45025,N_45347);
and U45599 (N_45599,N_45041,N_45301);
or U45600 (N_45600,N_45313,N_45049);
nand U45601 (N_45601,N_45331,N_45039);
xor U45602 (N_45602,N_45055,N_45467);
nand U45603 (N_45603,N_45035,N_45075);
nand U45604 (N_45604,N_45368,N_45175);
and U45605 (N_45605,N_45357,N_45059);
and U45606 (N_45606,N_45184,N_45170);
nand U45607 (N_45607,N_45238,N_45465);
nand U45608 (N_45608,N_45457,N_45438);
or U45609 (N_45609,N_45210,N_45228);
nand U45610 (N_45610,N_45386,N_45308);
nor U45611 (N_45611,N_45403,N_45196);
nor U45612 (N_45612,N_45152,N_45239);
nor U45613 (N_45613,N_45208,N_45286);
nand U45614 (N_45614,N_45458,N_45445);
xor U45615 (N_45615,N_45024,N_45124);
or U45616 (N_45616,N_45176,N_45489);
and U45617 (N_45617,N_45189,N_45482);
or U45618 (N_45618,N_45478,N_45485);
xnor U45619 (N_45619,N_45097,N_45287);
or U45620 (N_45620,N_45327,N_45247);
xor U45621 (N_45621,N_45005,N_45254);
xor U45622 (N_45622,N_45323,N_45235);
xor U45623 (N_45623,N_45070,N_45197);
and U45624 (N_45624,N_45092,N_45293);
and U45625 (N_45625,N_45371,N_45285);
nor U45626 (N_45626,N_45479,N_45063);
nor U45627 (N_45627,N_45067,N_45151);
and U45628 (N_45628,N_45338,N_45242);
nand U45629 (N_45629,N_45404,N_45166);
nand U45630 (N_45630,N_45452,N_45294);
xnor U45631 (N_45631,N_45430,N_45026);
and U45632 (N_45632,N_45145,N_45186);
xor U45633 (N_45633,N_45246,N_45010);
nand U45634 (N_45634,N_45261,N_45080);
or U45635 (N_45635,N_45022,N_45079);
nor U45636 (N_45636,N_45048,N_45019);
xor U45637 (N_45637,N_45429,N_45233);
or U45638 (N_45638,N_45229,N_45008);
nor U45639 (N_45639,N_45272,N_45120);
nor U45640 (N_45640,N_45476,N_45395);
nand U45641 (N_45641,N_45204,N_45365);
and U45642 (N_45642,N_45202,N_45177);
and U45643 (N_45643,N_45206,N_45220);
nand U45644 (N_45644,N_45304,N_45435);
and U45645 (N_45645,N_45366,N_45123);
nand U45646 (N_45646,N_45446,N_45030);
or U45647 (N_45647,N_45046,N_45351);
xor U45648 (N_45648,N_45473,N_45139);
nor U45649 (N_45649,N_45295,N_45459);
or U45650 (N_45650,N_45337,N_45215);
and U45651 (N_45651,N_45469,N_45236);
xor U45652 (N_45652,N_45421,N_45099);
or U45653 (N_45653,N_45387,N_45491);
or U45654 (N_45654,N_45111,N_45182);
and U45655 (N_45655,N_45064,N_45086);
nor U45656 (N_45656,N_45167,N_45128);
nor U45657 (N_45657,N_45460,N_45187);
and U45658 (N_45658,N_45122,N_45012);
and U45659 (N_45659,N_45448,N_45360);
or U45660 (N_45660,N_45044,N_45095);
and U45661 (N_45661,N_45082,N_45101);
or U45662 (N_45662,N_45009,N_45283);
xnor U45663 (N_45663,N_45226,N_45162);
and U45664 (N_45664,N_45014,N_45426);
nand U45665 (N_45665,N_45115,N_45319);
xnor U45666 (N_45666,N_45230,N_45045);
or U45667 (N_45667,N_45134,N_45052);
nand U45668 (N_45668,N_45361,N_45149);
nor U45669 (N_45669,N_45156,N_45316);
nand U45670 (N_45670,N_45188,N_45031);
nand U45671 (N_45671,N_45013,N_45389);
nand U45672 (N_45672,N_45066,N_45370);
nand U45673 (N_45673,N_45249,N_45036);
and U45674 (N_45674,N_45381,N_45486);
nand U45675 (N_45675,N_45051,N_45276);
xor U45676 (N_45676,N_45367,N_45310);
nor U45677 (N_45677,N_45349,N_45335);
or U45678 (N_45678,N_45300,N_45069);
and U45679 (N_45679,N_45245,N_45068);
or U45680 (N_45680,N_45320,N_45490);
nor U45681 (N_45681,N_45135,N_45328);
nand U45682 (N_45682,N_45280,N_45379);
nor U45683 (N_45683,N_45384,N_45492);
xnor U45684 (N_45684,N_45364,N_45207);
or U45685 (N_45685,N_45383,N_45169);
or U45686 (N_45686,N_45317,N_45255);
xnor U45687 (N_45687,N_45375,N_45017);
and U45688 (N_45688,N_45410,N_45198);
nor U45689 (N_45689,N_45094,N_45183);
or U45690 (N_45690,N_45418,N_45102);
xnor U45691 (N_45691,N_45499,N_45380);
nand U45692 (N_45692,N_45269,N_45394);
xnor U45693 (N_45693,N_45085,N_45472);
nand U45694 (N_45694,N_45471,N_45155);
and U45695 (N_45695,N_45273,N_45440);
nand U45696 (N_45696,N_45091,N_45456);
or U45697 (N_45697,N_45306,N_45298);
nand U45698 (N_45698,N_45225,N_45296);
nand U45699 (N_45699,N_45163,N_45431);
nor U45700 (N_45700,N_45330,N_45311);
nor U45701 (N_45701,N_45110,N_45401);
and U45702 (N_45702,N_45065,N_45480);
nand U45703 (N_45703,N_45326,N_45021);
nor U45704 (N_45704,N_45032,N_45405);
nand U45705 (N_45705,N_45322,N_45411);
and U45706 (N_45706,N_45374,N_45466);
xor U45707 (N_45707,N_45372,N_45353);
nand U45708 (N_45708,N_45000,N_45129);
and U45709 (N_45709,N_45463,N_45428);
or U45710 (N_45710,N_45454,N_45475);
xnor U45711 (N_45711,N_45302,N_45305);
xor U45712 (N_45712,N_45398,N_45248);
and U45713 (N_45713,N_45307,N_45420);
nand U45714 (N_45714,N_45015,N_45362);
nand U45715 (N_45715,N_45057,N_45098);
and U45716 (N_45716,N_45027,N_45439);
or U45717 (N_45717,N_45224,N_45336);
nand U45718 (N_45718,N_45339,N_45251);
xor U45719 (N_45719,N_45205,N_45369);
nand U45720 (N_45720,N_45158,N_45214);
nand U45721 (N_45721,N_45382,N_45292);
nand U45722 (N_45722,N_45171,N_45213);
or U45723 (N_45723,N_45352,N_45450);
nand U45724 (N_45724,N_45271,N_45416);
nand U45725 (N_45725,N_45274,N_45278);
xor U45726 (N_45726,N_45223,N_45315);
nor U45727 (N_45727,N_45221,N_45108);
nor U45728 (N_45728,N_45260,N_45427);
xnor U45729 (N_45729,N_45109,N_45191);
nor U45730 (N_45730,N_45040,N_45346);
xor U45731 (N_45731,N_45393,N_45142);
nor U45732 (N_45732,N_45056,N_45136);
nor U45733 (N_45733,N_45354,N_45054);
or U45734 (N_45734,N_45267,N_45174);
nor U45735 (N_45735,N_45001,N_45344);
nand U45736 (N_45736,N_45345,N_45081);
nor U45737 (N_45737,N_45377,N_45329);
and U45738 (N_45738,N_45194,N_45150);
nor U45739 (N_45739,N_45200,N_45443);
nor U45740 (N_45740,N_45424,N_45141);
xor U45741 (N_45741,N_45209,N_45161);
nor U45742 (N_45742,N_45147,N_45391);
xnor U45743 (N_45743,N_45199,N_45073);
nand U45744 (N_45744,N_45153,N_45348);
nor U45745 (N_45745,N_45444,N_45126);
and U45746 (N_45746,N_45203,N_45185);
nor U45747 (N_45747,N_45243,N_45483);
xor U45748 (N_45748,N_45333,N_45434);
or U45749 (N_45749,N_45498,N_45363);
nand U45750 (N_45750,N_45034,N_45049);
and U45751 (N_45751,N_45110,N_45028);
and U45752 (N_45752,N_45450,N_45349);
or U45753 (N_45753,N_45310,N_45133);
or U45754 (N_45754,N_45481,N_45116);
or U45755 (N_45755,N_45171,N_45476);
nor U45756 (N_45756,N_45000,N_45496);
nor U45757 (N_45757,N_45285,N_45066);
or U45758 (N_45758,N_45077,N_45213);
or U45759 (N_45759,N_45339,N_45430);
or U45760 (N_45760,N_45355,N_45390);
nand U45761 (N_45761,N_45416,N_45478);
xnor U45762 (N_45762,N_45484,N_45337);
and U45763 (N_45763,N_45304,N_45400);
or U45764 (N_45764,N_45264,N_45329);
or U45765 (N_45765,N_45340,N_45082);
xor U45766 (N_45766,N_45151,N_45298);
nor U45767 (N_45767,N_45046,N_45197);
nor U45768 (N_45768,N_45021,N_45137);
or U45769 (N_45769,N_45017,N_45377);
and U45770 (N_45770,N_45270,N_45069);
nand U45771 (N_45771,N_45270,N_45114);
or U45772 (N_45772,N_45278,N_45018);
and U45773 (N_45773,N_45216,N_45005);
nor U45774 (N_45774,N_45420,N_45313);
xnor U45775 (N_45775,N_45402,N_45049);
or U45776 (N_45776,N_45378,N_45367);
xnor U45777 (N_45777,N_45088,N_45127);
or U45778 (N_45778,N_45268,N_45160);
and U45779 (N_45779,N_45343,N_45188);
xnor U45780 (N_45780,N_45289,N_45093);
nor U45781 (N_45781,N_45478,N_45490);
xnor U45782 (N_45782,N_45065,N_45123);
nor U45783 (N_45783,N_45022,N_45318);
xnor U45784 (N_45784,N_45431,N_45142);
or U45785 (N_45785,N_45130,N_45271);
and U45786 (N_45786,N_45470,N_45042);
nor U45787 (N_45787,N_45405,N_45106);
nand U45788 (N_45788,N_45430,N_45203);
xnor U45789 (N_45789,N_45020,N_45443);
or U45790 (N_45790,N_45301,N_45181);
and U45791 (N_45791,N_45272,N_45190);
or U45792 (N_45792,N_45368,N_45425);
nor U45793 (N_45793,N_45305,N_45190);
xnor U45794 (N_45794,N_45295,N_45224);
nand U45795 (N_45795,N_45177,N_45244);
or U45796 (N_45796,N_45244,N_45010);
and U45797 (N_45797,N_45300,N_45418);
xnor U45798 (N_45798,N_45222,N_45336);
and U45799 (N_45799,N_45166,N_45409);
nor U45800 (N_45800,N_45032,N_45329);
nor U45801 (N_45801,N_45310,N_45221);
xor U45802 (N_45802,N_45482,N_45284);
and U45803 (N_45803,N_45033,N_45158);
or U45804 (N_45804,N_45117,N_45321);
nand U45805 (N_45805,N_45210,N_45291);
or U45806 (N_45806,N_45475,N_45389);
xnor U45807 (N_45807,N_45180,N_45451);
nor U45808 (N_45808,N_45286,N_45257);
nand U45809 (N_45809,N_45192,N_45268);
nand U45810 (N_45810,N_45024,N_45424);
xnor U45811 (N_45811,N_45294,N_45044);
nor U45812 (N_45812,N_45251,N_45269);
and U45813 (N_45813,N_45206,N_45432);
or U45814 (N_45814,N_45335,N_45092);
or U45815 (N_45815,N_45498,N_45163);
or U45816 (N_45816,N_45431,N_45006);
nor U45817 (N_45817,N_45096,N_45315);
or U45818 (N_45818,N_45487,N_45178);
xor U45819 (N_45819,N_45232,N_45031);
xor U45820 (N_45820,N_45338,N_45199);
and U45821 (N_45821,N_45221,N_45280);
nor U45822 (N_45822,N_45111,N_45146);
nand U45823 (N_45823,N_45358,N_45269);
nand U45824 (N_45824,N_45341,N_45400);
or U45825 (N_45825,N_45174,N_45461);
or U45826 (N_45826,N_45016,N_45032);
and U45827 (N_45827,N_45497,N_45253);
xnor U45828 (N_45828,N_45366,N_45195);
and U45829 (N_45829,N_45183,N_45202);
nand U45830 (N_45830,N_45432,N_45216);
xor U45831 (N_45831,N_45055,N_45027);
and U45832 (N_45832,N_45086,N_45299);
xor U45833 (N_45833,N_45065,N_45431);
nor U45834 (N_45834,N_45089,N_45279);
nand U45835 (N_45835,N_45041,N_45413);
xnor U45836 (N_45836,N_45199,N_45275);
and U45837 (N_45837,N_45079,N_45271);
nand U45838 (N_45838,N_45176,N_45491);
nand U45839 (N_45839,N_45481,N_45010);
nand U45840 (N_45840,N_45407,N_45143);
or U45841 (N_45841,N_45091,N_45490);
and U45842 (N_45842,N_45487,N_45282);
nand U45843 (N_45843,N_45273,N_45215);
xnor U45844 (N_45844,N_45070,N_45476);
nor U45845 (N_45845,N_45424,N_45480);
or U45846 (N_45846,N_45440,N_45283);
nor U45847 (N_45847,N_45005,N_45165);
xnor U45848 (N_45848,N_45332,N_45428);
nand U45849 (N_45849,N_45247,N_45470);
xnor U45850 (N_45850,N_45446,N_45294);
xor U45851 (N_45851,N_45131,N_45353);
nor U45852 (N_45852,N_45483,N_45010);
nand U45853 (N_45853,N_45437,N_45004);
nand U45854 (N_45854,N_45356,N_45383);
nor U45855 (N_45855,N_45469,N_45305);
and U45856 (N_45856,N_45402,N_45303);
and U45857 (N_45857,N_45154,N_45362);
nor U45858 (N_45858,N_45301,N_45233);
nand U45859 (N_45859,N_45028,N_45375);
and U45860 (N_45860,N_45329,N_45304);
or U45861 (N_45861,N_45081,N_45058);
nor U45862 (N_45862,N_45368,N_45039);
nor U45863 (N_45863,N_45004,N_45401);
nand U45864 (N_45864,N_45293,N_45097);
nor U45865 (N_45865,N_45198,N_45477);
nor U45866 (N_45866,N_45353,N_45308);
xnor U45867 (N_45867,N_45258,N_45032);
xor U45868 (N_45868,N_45046,N_45163);
and U45869 (N_45869,N_45127,N_45148);
nand U45870 (N_45870,N_45300,N_45133);
nand U45871 (N_45871,N_45320,N_45114);
and U45872 (N_45872,N_45279,N_45020);
xnor U45873 (N_45873,N_45186,N_45456);
xor U45874 (N_45874,N_45371,N_45234);
nand U45875 (N_45875,N_45200,N_45479);
nor U45876 (N_45876,N_45290,N_45095);
or U45877 (N_45877,N_45223,N_45460);
and U45878 (N_45878,N_45108,N_45487);
nor U45879 (N_45879,N_45267,N_45161);
or U45880 (N_45880,N_45429,N_45292);
nand U45881 (N_45881,N_45029,N_45158);
and U45882 (N_45882,N_45103,N_45374);
or U45883 (N_45883,N_45291,N_45400);
and U45884 (N_45884,N_45208,N_45349);
xnor U45885 (N_45885,N_45257,N_45365);
xor U45886 (N_45886,N_45332,N_45339);
or U45887 (N_45887,N_45413,N_45126);
nor U45888 (N_45888,N_45027,N_45117);
nor U45889 (N_45889,N_45414,N_45398);
nand U45890 (N_45890,N_45077,N_45404);
and U45891 (N_45891,N_45131,N_45469);
nand U45892 (N_45892,N_45032,N_45446);
or U45893 (N_45893,N_45254,N_45365);
and U45894 (N_45894,N_45279,N_45419);
or U45895 (N_45895,N_45310,N_45123);
or U45896 (N_45896,N_45027,N_45495);
and U45897 (N_45897,N_45424,N_45048);
nor U45898 (N_45898,N_45131,N_45371);
nand U45899 (N_45899,N_45103,N_45475);
nand U45900 (N_45900,N_45283,N_45033);
nor U45901 (N_45901,N_45045,N_45085);
or U45902 (N_45902,N_45216,N_45409);
xnor U45903 (N_45903,N_45430,N_45327);
nor U45904 (N_45904,N_45264,N_45414);
xor U45905 (N_45905,N_45112,N_45264);
nand U45906 (N_45906,N_45380,N_45375);
nand U45907 (N_45907,N_45127,N_45159);
nand U45908 (N_45908,N_45420,N_45061);
and U45909 (N_45909,N_45438,N_45244);
nand U45910 (N_45910,N_45247,N_45274);
nor U45911 (N_45911,N_45479,N_45415);
nand U45912 (N_45912,N_45058,N_45407);
xor U45913 (N_45913,N_45066,N_45479);
or U45914 (N_45914,N_45389,N_45408);
nor U45915 (N_45915,N_45154,N_45072);
nor U45916 (N_45916,N_45303,N_45420);
or U45917 (N_45917,N_45418,N_45221);
nand U45918 (N_45918,N_45223,N_45313);
nor U45919 (N_45919,N_45461,N_45168);
nor U45920 (N_45920,N_45412,N_45465);
nand U45921 (N_45921,N_45396,N_45062);
nand U45922 (N_45922,N_45365,N_45044);
nand U45923 (N_45923,N_45480,N_45315);
nand U45924 (N_45924,N_45268,N_45149);
nand U45925 (N_45925,N_45224,N_45086);
nand U45926 (N_45926,N_45366,N_45182);
and U45927 (N_45927,N_45491,N_45036);
nand U45928 (N_45928,N_45270,N_45377);
and U45929 (N_45929,N_45216,N_45445);
nor U45930 (N_45930,N_45370,N_45279);
nor U45931 (N_45931,N_45372,N_45377);
xnor U45932 (N_45932,N_45487,N_45062);
and U45933 (N_45933,N_45101,N_45056);
or U45934 (N_45934,N_45135,N_45432);
nand U45935 (N_45935,N_45026,N_45340);
or U45936 (N_45936,N_45032,N_45084);
or U45937 (N_45937,N_45309,N_45335);
nand U45938 (N_45938,N_45310,N_45236);
or U45939 (N_45939,N_45225,N_45019);
or U45940 (N_45940,N_45281,N_45090);
xnor U45941 (N_45941,N_45486,N_45403);
nor U45942 (N_45942,N_45035,N_45198);
or U45943 (N_45943,N_45153,N_45017);
nor U45944 (N_45944,N_45389,N_45120);
or U45945 (N_45945,N_45129,N_45427);
nor U45946 (N_45946,N_45262,N_45318);
nor U45947 (N_45947,N_45415,N_45493);
xnor U45948 (N_45948,N_45064,N_45492);
nand U45949 (N_45949,N_45180,N_45277);
nand U45950 (N_45950,N_45446,N_45099);
or U45951 (N_45951,N_45393,N_45001);
or U45952 (N_45952,N_45246,N_45352);
nand U45953 (N_45953,N_45032,N_45070);
and U45954 (N_45954,N_45117,N_45182);
xor U45955 (N_45955,N_45421,N_45261);
nor U45956 (N_45956,N_45412,N_45023);
nor U45957 (N_45957,N_45362,N_45276);
and U45958 (N_45958,N_45073,N_45153);
nor U45959 (N_45959,N_45323,N_45122);
and U45960 (N_45960,N_45409,N_45055);
or U45961 (N_45961,N_45318,N_45088);
and U45962 (N_45962,N_45166,N_45180);
xor U45963 (N_45963,N_45242,N_45368);
or U45964 (N_45964,N_45263,N_45038);
nand U45965 (N_45965,N_45208,N_45007);
or U45966 (N_45966,N_45278,N_45131);
nand U45967 (N_45967,N_45455,N_45443);
nand U45968 (N_45968,N_45429,N_45052);
xor U45969 (N_45969,N_45291,N_45337);
and U45970 (N_45970,N_45064,N_45260);
or U45971 (N_45971,N_45192,N_45175);
nand U45972 (N_45972,N_45191,N_45476);
nor U45973 (N_45973,N_45341,N_45146);
nor U45974 (N_45974,N_45032,N_45074);
and U45975 (N_45975,N_45009,N_45318);
nand U45976 (N_45976,N_45283,N_45369);
nand U45977 (N_45977,N_45368,N_45413);
nand U45978 (N_45978,N_45296,N_45252);
nor U45979 (N_45979,N_45363,N_45305);
and U45980 (N_45980,N_45092,N_45288);
or U45981 (N_45981,N_45161,N_45389);
nand U45982 (N_45982,N_45335,N_45104);
nor U45983 (N_45983,N_45221,N_45492);
and U45984 (N_45984,N_45089,N_45259);
xnor U45985 (N_45985,N_45032,N_45119);
nor U45986 (N_45986,N_45196,N_45206);
and U45987 (N_45987,N_45175,N_45479);
xor U45988 (N_45988,N_45298,N_45003);
and U45989 (N_45989,N_45468,N_45110);
or U45990 (N_45990,N_45281,N_45076);
nand U45991 (N_45991,N_45261,N_45463);
nor U45992 (N_45992,N_45385,N_45149);
and U45993 (N_45993,N_45280,N_45499);
or U45994 (N_45994,N_45229,N_45059);
or U45995 (N_45995,N_45337,N_45486);
xnor U45996 (N_45996,N_45370,N_45262);
or U45997 (N_45997,N_45490,N_45048);
nand U45998 (N_45998,N_45469,N_45293);
xor U45999 (N_45999,N_45284,N_45058);
nor U46000 (N_46000,N_45738,N_45993);
nand U46001 (N_46001,N_45866,N_45750);
or U46002 (N_46002,N_45604,N_45907);
nor U46003 (N_46003,N_45904,N_45963);
nor U46004 (N_46004,N_45821,N_45930);
xnor U46005 (N_46005,N_45691,N_45775);
or U46006 (N_46006,N_45795,N_45803);
nor U46007 (N_46007,N_45862,N_45532);
or U46008 (N_46008,N_45847,N_45785);
or U46009 (N_46009,N_45662,N_45998);
nor U46010 (N_46010,N_45542,N_45936);
and U46011 (N_46011,N_45708,N_45741);
and U46012 (N_46012,N_45781,N_45910);
or U46013 (N_46013,N_45545,N_45576);
nor U46014 (N_46014,N_45796,N_45820);
or U46015 (N_46015,N_45724,N_45503);
xnor U46016 (N_46016,N_45509,N_45619);
or U46017 (N_46017,N_45739,N_45679);
xor U46018 (N_46018,N_45874,N_45506);
nor U46019 (N_46019,N_45835,N_45965);
nor U46020 (N_46020,N_45895,N_45642);
or U46021 (N_46021,N_45636,N_45653);
xor U46022 (N_46022,N_45972,N_45908);
or U46023 (N_46023,N_45746,N_45588);
xnor U46024 (N_46024,N_45892,N_45647);
nand U46025 (N_46025,N_45535,N_45769);
or U46026 (N_46026,N_45783,N_45685);
xor U46027 (N_46027,N_45712,N_45823);
or U46028 (N_46028,N_45810,N_45728);
and U46029 (N_46029,N_45664,N_45852);
xor U46030 (N_46030,N_45797,N_45901);
or U46031 (N_46031,N_45736,N_45782);
and U46032 (N_46032,N_45777,N_45707);
nor U46033 (N_46033,N_45540,N_45935);
and U46034 (N_46034,N_45857,N_45505);
and U46035 (N_46035,N_45853,N_45987);
nor U46036 (N_46036,N_45650,N_45523);
nor U46037 (N_46037,N_45673,N_45630);
xor U46038 (N_46038,N_45992,N_45859);
or U46039 (N_46039,N_45512,N_45861);
xor U46040 (N_46040,N_45511,N_45982);
and U46041 (N_46041,N_45787,N_45565);
and U46042 (N_46042,N_45966,N_45578);
or U46043 (N_46043,N_45942,N_45677);
xor U46044 (N_46044,N_45594,N_45549);
or U46045 (N_46045,N_45533,N_45557);
xor U46046 (N_46046,N_45695,N_45550);
nor U46047 (N_46047,N_45943,N_45669);
and U46048 (N_46048,N_45994,N_45985);
nor U46049 (N_46049,N_45706,N_45940);
nor U46050 (N_46050,N_45517,N_45825);
nor U46051 (N_46051,N_45784,N_45960);
nand U46052 (N_46052,N_45941,N_45589);
nand U46053 (N_46053,N_45932,N_45722);
xnor U46054 (N_46054,N_45951,N_45905);
xor U46055 (N_46055,N_45568,N_45926);
and U46056 (N_46056,N_45639,N_45661);
xor U46057 (N_46057,N_45928,N_45909);
nand U46058 (N_46058,N_45678,N_45916);
or U46059 (N_46059,N_45745,N_45969);
nor U46060 (N_46060,N_45897,N_45865);
nor U46061 (N_46061,N_45529,N_45676);
xor U46062 (N_46062,N_45592,N_45575);
nor U46063 (N_46063,N_45684,N_45502);
and U46064 (N_46064,N_45615,N_45889);
nor U46065 (N_46065,N_45875,N_45606);
or U46066 (N_46066,N_45863,N_45946);
nand U46067 (N_46067,N_45968,N_45513);
xnor U46068 (N_46068,N_45962,N_45717);
or U46069 (N_46069,N_45551,N_45776);
and U46070 (N_46070,N_45516,N_45806);
or U46071 (N_46071,N_45850,N_45885);
or U46072 (N_46072,N_45725,N_45629);
nand U46073 (N_46073,N_45976,N_45983);
nor U46074 (N_46074,N_45811,N_45559);
and U46075 (N_46075,N_45607,N_45819);
nand U46076 (N_46076,N_45918,N_45524);
xnor U46077 (N_46077,N_45666,N_45854);
or U46078 (N_46078,N_45543,N_45654);
or U46079 (N_46079,N_45881,N_45837);
and U46080 (N_46080,N_45772,N_45798);
and U46081 (N_46081,N_45700,N_45956);
nand U46082 (N_46082,N_45878,N_45729);
or U46083 (N_46083,N_45980,N_45743);
nor U46084 (N_46084,N_45974,N_45561);
nand U46085 (N_46085,N_45590,N_45698);
nand U46086 (N_46086,N_45912,N_45919);
nor U46087 (N_46087,N_45644,N_45933);
nand U46088 (N_46088,N_45587,N_45601);
nor U46089 (N_46089,N_45573,N_45947);
and U46090 (N_46090,N_45719,N_45760);
and U46091 (N_46091,N_45522,N_45788);
nand U46092 (N_46092,N_45582,N_45893);
and U46093 (N_46093,N_45789,N_45514);
and U46094 (N_46094,N_45714,N_45979);
nor U46095 (N_46095,N_45626,N_45780);
nand U46096 (N_46096,N_45603,N_45631);
nor U46097 (N_46097,N_45656,N_45556);
xnor U46098 (N_46098,N_45634,N_45842);
nand U46099 (N_46099,N_45884,N_45686);
nand U46100 (N_46100,N_45944,N_45655);
and U46101 (N_46101,N_45814,N_45975);
and U46102 (N_46102,N_45687,N_45816);
nand U46103 (N_46103,N_45703,N_45716);
or U46104 (N_46104,N_45681,N_45735);
xnor U46105 (N_46105,N_45931,N_45660);
and U46106 (N_46106,N_45574,N_45697);
nor U46107 (N_46107,N_45632,N_45737);
xor U46108 (N_46108,N_45710,N_45818);
nor U46109 (N_46109,N_45809,N_45709);
or U46110 (N_46110,N_45620,N_45824);
nor U46111 (N_46111,N_45637,N_45510);
and U46112 (N_46112,N_45548,N_45757);
xor U46113 (N_46113,N_45826,N_45732);
nor U46114 (N_46114,N_45845,N_45527);
or U46115 (N_46115,N_45900,N_45999);
nor U46116 (N_46116,N_45569,N_45558);
nor U46117 (N_46117,N_45635,N_45683);
and U46118 (N_46118,N_45733,N_45715);
nor U46119 (N_46119,N_45526,N_45793);
nor U46120 (N_46120,N_45720,N_45779);
xnor U46121 (N_46121,N_45856,N_45663);
or U46122 (N_46122,N_45989,N_45657);
nor U46123 (N_46123,N_45817,N_45829);
nor U46124 (N_46124,N_45536,N_45794);
and U46125 (N_46125,N_45538,N_45734);
nand U46126 (N_46126,N_45768,N_45896);
and U46127 (N_46127,N_45501,N_45858);
nor U46128 (N_46128,N_45830,N_45571);
or U46129 (N_46129,N_45581,N_45986);
xnor U46130 (N_46130,N_45713,N_45701);
or U46131 (N_46131,N_45831,N_45838);
nand U46132 (N_46132,N_45953,N_45903);
and U46133 (N_46133,N_45583,N_45723);
and U46134 (N_46134,N_45744,N_45843);
and U46135 (N_46135,N_45923,N_45751);
xor U46136 (N_46136,N_45566,N_45705);
and U46137 (N_46137,N_45537,N_45898);
nand U46138 (N_46138,N_45704,N_45572);
nand U46139 (N_46139,N_45761,N_45645);
or U46140 (N_46140,N_45579,N_45802);
nand U46141 (N_46141,N_45869,N_45890);
xnor U46142 (N_46142,N_45627,N_45786);
nand U46143 (N_46143,N_45871,N_45613);
or U46144 (N_46144,N_45860,N_45805);
or U46145 (N_46145,N_45959,N_45937);
xor U46146 (N_46146,N_45648,N_45879);
and U46147 (N_46147,N_45555,N_45675);
and U46148 (N_46148,N_45610,N_45602);
xnor U46149 (N_46149,N_45617,N_45870);
xnor U46150 (N_46150,N_45521,N_45597);
or U46151 (N_46151,N_45753,N_45585);
or U46152 (N_46152,N_45508,N_45833);
nor U46153 (N_46153,N_45696,N_45515);
xnor U46154 (N_46154,N_45528,N_45841);
or U46155 (N_46155,N_45808,N_45672);
and U46156 (N_46156,N_45518,N_45883);
and U46157 (N_46157,N_45880,N_45693);
nor U46158 (N_46158,N_45978,N_45546);
or U46159 (N_46159,N_45921,N_45608);
xnor U46160 (N_46160,N_45711,N_45766);
nand U46161 (N_46161,N_45873,N_45680);
nor U46162 (N_46162,N_45553,N_45544);
and U46163 (N_46163,N_45500,N_45665);
and U46164 (N_46164,N_45756,N_45752);
or U46165 (N_46165,N_45560,N_45564);
or U46166 (N_46166,N_45888,N_45957);
xor U46167 (N_46167,N_45844,N_45577);
and U46168 (N_46168,N_45682,N_45690);
xnor U46169 (N_46169,N_45834,N_45623);
and U46170 (N_46170,N_45727,N_45812);
xnor U46171 (N_46171,N_45770,N_45638);
and U46172 (N_46172,N_45902,N_45827);
nor U46173 (N_46173,N_45922,N_45791);
nor U46174 (N_46174,N_45547,N_45504);
xnor U46175 (N_46175,N_45598,N_45539);
nand U46176 (N_46176,N_45758,N_45882);
or U46177 (N_46177,N_45891,N_45764);
nand U46178 (N_46178,N_45939,N_45605);
xnor U46179 (N_46179,N_45997,N_45924);
and U46180 (N_46180,N_45584,N_45774);
nor U46181 (N_46181,N_45530,N_45990);
nand U46182 (N_46182,N_45804,N_45591);
or U46183 (N_46183,N_45967,N_45971);
xnor U46184 (N_46184,N_45649,N_45950);
xor U46185 (N_46185,N_45633,N_45984);
xnor U46186 (N_46186,N_45864,N_45920);
or U46187 (N_46187,N_45762,N_45815);
or U46188 (N_46188,N_45846,N_45973);
or U46189 (N_46189,N_45872,N_45507);
xor U46190 (N_46190,N_45541,N_45799);
or U46191 (N_46191,N_45894,N_45600);
xnor U46192 (N_46192,N_45927,N_45988);
and U46193 (N_46193,N_45742,N_45609);
or U46194 (N_46194,N_45567,N_45625);
xor U46195 (N_46195,N_45929,N_45913);
nand U46196 (N_46196,N_45915,N_45832);
and U46197 (N_46197,N_45778,N_45964);
or U46198 (N_46198,N_45658,N_45748);
and U46199 (N_46199,N_45595,N_45640);
xnor U46200 (N_46200,N_45887,N_45659);
xnor U46201 (N_46201,N_45612,N_45651);
xor U46202 (N_46202,N_45552,N_45749);
and U46203 (N_46203,N_45628,N_45828);
and U46204 (N_46204,N_45917,N_45840);
xor U46205 (N_46205,N_45955,N_45949);
or U46206 (N_46206,N_45689,N_45614);
nand U46207 (N_46207,N_45991,N_45580);
nor U46208 (N_46208,N_45755,N_45611);
and U46209 (N_46209,N_45970,N_45868);
nand U46210 (N_46210,N_45906,N_45934);
and U46211 (N_46211,N_45562,N_45643);
nand U46212 (N_46212,N_45876,N_45726);
or U46213 (N_46213,N_45867,N_45563);
or U46214 (N_46214,N_45622,N_45948);
or U46215 (N_46215,N_45822,N_45790);
nand U46216 (N_46216,N_45855,N_45740);
or U46217 (N_46217,N_45621,N_45702);
and U46218 (N_46218,N_45667,N_45886);
xnor U46219 (N_46219,N_45759,N_45995);
xnor U46220 (N_46220,N_45839,N_45747);
xor U46221 (N_46221,N_45773,N_45731);
xor U46222 (N_46222,N_45996,N_45848);
xor U46223 (N_46223,N_45914,N_45674);
or U46224 (N_46224,N_45618,N_45792);
nor U46225 (N_46225,N_45721,N_45670);
and U46226 (N_46226,N_45718,N_45925);
nor U46227 (N_46227,N_45671,N_45899);
nor U46228 (N_46228,N_45641,N_45765);
nor U46229 (N_46229,N_45570,N_45836);
nand U46230 (N_46230,N_45616,N_45730);
and U46231 (N_46231,N_45599,N_45813);
or U46232 (N_46232,N_45807,N_45694);
nor U46233 (N_46233,N_45877,N_45954);
nor U46234 (N_46234,N_45981,N_45624);
or U46235 (N_46235,N_45596,N_45534);
xnor U46236 (N_46236,N_45525,N_45531);
and U46237 (N_46237,N_45593,N_45668);
nand U46238 (N_46238,N_45646,N_45911);
nand U46239 (N_46239,N_45771,N_45938);
nand U46240 (N_46240,N_45692,N_45586);
and U46241 (N_46241,N_45763,N_45952);
nand U46242 (N_46242,N_45945,N_45958);
nand U46243 (N_46243,N_45800,N_45849);
nor U46244 (N_46244,N_45688,N_45554);
or U46245 (N_46245,N_45851,N_45754);
xor U46246 (N_46246,N_45520,N_45519);
and U46247 (N_46247,N_45801,N_45767);
nand U46248 (N_46248,N_45699,N_45961);
xor U46249 (N_46249,N_45652,N_45977);
xnor U46250 (N_46250,N_45580,N_45741);
or U46251 (N_46251,N_45624,N_45942);
and U46252 (N_46252,N_45519,N_45780);
nand U46253 (N_46253,N_45759,N_45697);
or U46254 (N_46254,N_45955,N_45775);
nor U46255 (N_46255,N_45853,N_45735);
and U46256 (N_46256,N_45966,N_45969);
nor U46257 (N_46257,N_45586,N_45688);
nand U46258 (N_46258,N_45546,N_45908);
or U46259 (N_46259,N_45815,N_45646);
nand U46260 (N_46260,N_45900,N_45690);
xnor U46261 (N_46261,N_45617,N_45965);
nand U46262 (N_46262,N_45605,N_45991);
or U46263 (N_46263,N_45876,N_45902);
and U46264 (N_46264,N_45897,N_45894);
nor U46265 (N_46265,N_45795,N_45953);
or U46266 (N_46266,N_45622,N_45831);
and U46267 (N_46267,N_45602,N_45530);
or U46268 (N_46268,N_45674,N_45939);
and U46269 (N_46269,N_45504,N_45688);
nor U46270 (N_46270,N_45959,N_45674);
or U46271 (N_46271,N_45730,N_45631);
xnor U46272 (N_46272,N_45898,N_45706);
xor U46273 (N_46273,N_45522,N_45676);
xor U46274 (N_46274,N_45764,N_45600);
xnor U46275 (N_46275,N_45609,N_45895);
xnor U46276 (N_46276,N_45710,N_45962);
nand U46277 (N_46277,N_45823,N_45506);
and U46278 (N_46278,N_45638,N_45986);
nor U46279 (N_46279,N_45840,N_45538);
nor U46280 (N_46280,N_45792,N_45560);
xor U46281 (N_46281,N_45646,N_45929);
xor U46282 (N_46282,N_45868,N_45888);
xor U46283 (N_46283,N_45905,N_45592);
nor U46284 (N_46284,N_45627,N_45592);
or U46285 (N_46285,N_45736,N_45546);
nor U46286 (N_46286,N_45961,N_45572);
nand U46287 (N_46287,N_45768,N_45647);
xnor U46288 (N_46288,N_45905,N_45695);
nand U46289 (N_46289,N_45676,N_45931);
xnor U46290 (N_46290,N_45817,N_45601);
nand U46291 (N_46291,N_45808,N_45620);
xor U46292 (N_46292,N_45854,N_45966);
or U46293 (N_46293,N_45873,N_45769);
and U46294 (N_46294,N_45713,N_45501);
nor U46295 (N_46295,N_45785,N_45741);
or U46296 (N_46296,N_45684,N_45633);
or U46297 (N_46297,N_45805,N_45637);
nand U46298 (N_46298,N_45937,N_45669);
xor U46299 (N_46299,N_45729,N_45525);
nand U46300 (N_46300,N_45801,N_45972);
or U46301 (N_46301,N_45872,N_45543);
nand U46302 (N_46302,N_45847,N_45672);
nand U46303 (N_46303,N_45895,N_45620);
xor U46304 (N_46304,N_45809,N_45589);
nor U46305 (N_46305,N_45564,N_45517);
or U46306 (N_46306,N_45716,N_45745);
nor U46307 (N_46307,N_45938,N_45939);
and U46308 (N_46308,N_45645,N_45693);
xor U46309 (N_46309,N_45788,N_45801);
and U46310 (N_46310,N_45587,N_45505);
nand U46311 (N_46311,N_45609,N_45590);
xor U46312 (N_46312,N_45816,N_45661);
xor U46313 (N_46313,N_45853,N_45889);
nor U46314 (N_46314,N_45823,N_45510);
nand U46315 (N_46315,N_45874,N_45661);
nor U46316 (N_46316,N_45553,N_45512);
and U46317 (N_46317,N_45794,N_45851);
nand U46318 (N_46318,N_45820,N_45624);
and U46319 (N_46319,N_45727,N_45774);
or U46320 (N_46320,N_45945,N_45727);
nor U46321 (N_46321,N_45665,N_45716);
nor U46322 (N_46322,N_45960,N_45584);
xnor U46323 (N_46323,N_45862,N_45640);
nor U46324 (N_46324,N_45941,N_45944);
nand U46325 (N_46325,N_45856,N_45586);
nor U46326 (N_46326,N_45683,N_45892);
nor U46327 (N_46327,N_45520,N_45544);
nand U46328 (N_46328,N_45709,N_45799);
and U46329 (N_46329,N_45871,N_45883);
and U46330 (N_46330,N_45518,N_45500);
and U46331 (N_46331,N_45924,N_45764);
and U46332 (N_46332,N_45847,N_45618);
nand U46333 (N_46333,N_45698,N_45597);
or U46334 (N_46334,N_45666,N_45571);
or U46335 (N_46335,N_45976,N_45531);
nor U46336 (N_46336,N_45944,N_45823);
and U46337 (N_46337,N_45807,N_45965);
and U46338 (N_46338,N_45711,N_45827);
xor U46339 (N_46339,N_45929,N_45581);
and U46340 (N_46340,N_45636,N_45887);
nand U46341 (N_46341,N_45920,N_45625);
nor U46342 (N_46342,N_45584,N_45553);
nand U46343 (N_46343,N_45691,N_45730);
xor U46344 (N_46344,N_45565,N_45919);
xor U46345 (N_46345,N_45541,N_45579);
or U46346 (N_46346,N_45584,N_45716);
and U46347 (N_46347,N_45765,N_45909);
or U46348 (N_46348,N_45626,N_45532);
nand U46349 (N_46349,N_45997,N_45672);
and U46350 (N_46350,N_45788,N_45830);
xnor U46351 (N_46351,N_45984,N_45996);
or U46352 (N_46352,N_45786,N_45704);
xnor U46353 (N_46353,N_45793,N_45880);
xnor U46354 (N_46354,N_45567,N_45973);
xnor U46355 (N_46355,N_45638,N_45903);
or U46356 (N_46356,N_45537,N_45822);
xnor U46357 (N_46357,N_45824,N_45674);
nand U46358 (N_46358,N_45944,N_45801);
or U46359 (N_46359,N_45610,N_45700);
and U46360 (N_46360,N_45618,N_45558);
or U46361 (N_46361,N_45656,N_45503);
or U46362 (N_46362,N_45792,N_45955);
xor U46363 (N_46363,N_45786,N_45651);
xor U46364 (N_46364,N_45512,N_45567);
or U46365 (N_46365,N_45929,N_45975);
and U46366 (N_46366,N_45956,N_45897);
xnor U46367 (N_46367,N_45759,N_45816);
or U46368 (N_46368,N_45742,N_45831);
or U46369 (N_46369,N_45702,N_45830);
nand U46370 (N_46370,N_45555,N_45803);
or U46371 (N_46371,N_45981,N_45519);
nor U46372 (N_46372,N_45873,N_45714);
xnor U46373 (N_46373,N_45973,N_45839);
nand U46374 (N_46374,N_45716,N_45706);
nand U46375 (N_46375,N_45525,N_45719);
or U46376 (N_46376,N_45773,N_45713);
and U46377 (N_46377,N_45730,N_45579);
nand U46378 (N_46378,N_45616,N_45778);
and U46379 (N_46379,N_45595,N_45782);
and U46380 (N_46380,N_45616,N_45555);
nor U46381 (N_46381,N_45644,N_45597);
nor U46382 (N_46382,N_45860,N_45933);
xnor U46383 (N_46383,N_45650,N_45589);
or U46384 (N_46384,N_45794,N_45559);
or U46385 (N_46385,N_45526,N_45726);
nor U46386 (N_46386,N_45925,N_45558);
xnor U46387 (N_46387,N_45604,N_45915);
or U46388 (N_46388,N_45573,N_45677);
nand U46389 (N_46389,N_45877,N_45914);
xnor U46390 (N_46390,N_45966,N_45963);
nand U46391 (N_46391,N_45846,N_45608);
nor U46392 (N_46392,N_45737,N_45561);
nor U46393 (N_46393,N_45606,N_45637);
nor U46394 (N_46394,N_45555,N_45827);
and U46395 (N_46395,N_45681,N_45887);
nor U46396 (N_46396,N_45695,N_45869);
and U46397 (N_46397,N_45856,N_45744);
nand U46398 (N_46398,N_45535,N_45901);
and U46399 (N_46399,N_45943,N_45581);
nand U46400 (N_46400,N_45941,N_45832);
nor U46401 (N_46401,N_45822,N_45871);
xor U46402 (N_46402,N_45621,N_45800);
or U46403 (N_46403,N_45994,N_45526);
xnor U46404 (N_46404,N_45982,N_45999);
nand U46405 (N_46405,N_45548,N_45745);
nand U46406 (N_46406,N_45945,N_45633);
xor U46407 (N_46407,N_45686,N_45570);
xor U46408 (N_46408,N_45993,N_45964);
nor U46409 (N_46409,N_45738,N_45641);
nand U46410 (N_46410,N_45543,N_45896);
nor U46411 (N_46411,N_45661,N_45955);
or U46412 (N_46412,N_45699,N_45665);
xnor U46413 (N_46413,N_45939,N_45889);
xor U46414 (N_46414,N_45841,N_45662);
nor U46415 (N_46415,N_45660,N_45613);
and U46416 (N_46416,N_45566,N_45509);
nor U46417 (N_46417,N_45854,N_45662);
nand U46418 (N_46418,N_45746,N_45607);
xnor U46419 (N_46419,N_45768,N_45751);
or U46420 (N_46420,N_45731,N_45934);
nand U46421 (N_46421,N_45702,N_45965);
nor U46422 (N_46422,N_45967,N_45536);
xnor U46423 (N_46423,N_45970,N_45743);
nor U46424 (N_46424,N_45512,N_45848);
xor U46425 (N_46425,N_45998,N_45711);
nand U46426 (N_46426,N_45820,N_45952);
or U46427 (N_46427,N_45662,N_45997);
nand U46428 (N_46428,N_45560,N_45809);
xor U46429 (N_46429,N_45824,N_45702);
and U46430 (N_46430,N_45916,N_45817);
nor U46431 (N_46431,N_45788,N_45865);
nand U46432 (N_46432,N_45509,N_45742);
or U46433 (N_46433,N_45523,N_45844);
xnor U46434 (N_46434,N_45507,N_45820);
or U46435 (N_46435,N_45662,N_45630);
or U46436 (N_46436,N_45768,N_45874);
xor U46437 (N_46437,N_45908,N_45968);
and U46438 (N_46438,N_45882,N_45726);
nor U46439 (N_46439,N_45527,N_45906);
xor U46440 (N_46440,N_45941,N_45959);
nor U46441 (N_46441,N_45638,N_45803);
nand U46442 (N_46442,N_45631,N_45672);
or U46443 (N_46443,N_45522,N_45770);
nor U46444 (N_46444,N_45513,N_45777);
nand U46445 (N_46445,N_45831,N_45695);
or U46446 (N_46446,N_45804,N_45619);
xnor U46447 (N_46447,N_45784,N_45896);
xnor U46448 (N_46448,N_45513,N_45835);
xor U46449 (N_46449,N_45915,N_45760);
and U46450 (N_46450,N_45957,N_45637);
and U46451 (N_46451,N_45820,N_45785);
nor U46452 (N_46452,N_45697,N_45709);
and U46453 (N_46453,N_45523,N_45945);
xnor U46454 (N_46454,N_45552,N_45763);
xnor U46455 (N_46455,N_45567,N_45558);
xnor U46456 (N_46456,N_45799,N_45722);
xor U46457 (N_46457,N_45952,N_45940);
xnor U46458 (N_46458,N_45577,N_45662);
nand U46459 (N_46459,N_45707,N_45789);
and U46460 (N_46460,N_45690,N_45517);
or U46461 (N_46461,N_45504,N_45999);
xnor U46462 (N_46462,N_45514,N_45969);
xnor U46463 (N_46463,N_45590,N_45872);
nand U46464 (N_46464,N_45787,N_45718);
nor U46465 (N_46465,N_45634,N_45644);
and U46466 (N_46466,N_45662,N_45507);
or U46467 (N_46467,N_45698,N_45621);
nand U46468 (N_46468,N_45855,N_45816);
nand U46469 (N_46469,N_45628,N_45857);
and U46470 (N_46470,N_45792,N_45728);
nand U46471 (N_46471,N_45689,N_45752);
or U46472 (N_46472,N_45799,N_45935);
xnor U46473 (N_46473,N_45891,N_45815);
nand U46474 (N_46474,N_45546,N_45927);
nand U46475 (N_46475,N_45724,N_45676);
nand U46476 (N_46476,N_45615,N_45684);
nand U46477 (N_46477,N_45774,N_45697);
and U46478 (N_46478,N_45897,N_45529);
or U46479 (N_46479,N_45990,N_45921);
nor U46480 (N_46480,N_45796,N_45853);
nor U46481 (N_46481,N_45816,N_45956);
nand U46482 (N_46482,N_45845,N_45721);
nor U46483 (N_46483,N_45680,N_45669);
xor U46484 (N_46484,N_45737,N_45825);
nor U46485 (N_46485,N_45624,N_45703);
xnor U46486 (N_46486,N_45798,N_45932);
nand U46487 (N_46487,N_45800,N_45644);
nand U46488 (N_46488,N_45530,N_45580);
nand U46489 (N_46489,N_45935,N_45992);
or U46490 (N_46490,N_45549,N_45896);
and U46491 (N_46491,N_45993,N_45827);
xor U46492 (N_46492,N_45545,N_45810);
and U46493 (N_46493,N_45830,N_45785);
and U46494 (N_46494,N_45791,N_45614);
nand U46495 (N_46495,N_45869,N_45953);
nor U46496 (N_46496,N_45952,N_45690);
xnor U46497 (N_46497,N_45574,N_45743);
and U46498 (N_46498,N_45509,N_45901);
or U46499 (N_46499,N_45839,N_45513);
nor U46500 (N_46500,N_46066,N_46359);
and U46501 (N_46501,N_46170,N_46014);
nor U46502 (N_46502,N_46379,N_46012);
xnor U46503 (N_46503,N_46243,N_46380);
nand U46504 (N_46504,N_46462,N_46072);
nor U46505 (N_46505,N_46005,N_46038);
xor U46506 (N_46506,N_46445,N_46307);
nor U46507 (N_46507,N_46259,N_46371);
nand U46508 (N_46508,N_46401,N_46326);
nand U46509 (N_46509,N_46203,N_46087);
xnor U46510 (N_46510,N_46328,N_46024);
and U46511 (N_46511,N_46331,N_46162);
nand U46512 (N_46512,N_46316,N_46270);
nor U46513 (N_46513,N_46245,N_46150);
or U46514 (N_46514,N_46062,N_46323);
nor U46515 (N_46515,N_46443,N_46232);
xor U46516 (N_46516,N_46350,N_46406);
nor U46517 (N_46517,N_46099,N_46455);
nand U46518 (N_46518,N_46258,N_46273);
and U46519 (N_46519,N_46219,N_46132);
and U46520 (N_46520,N_46497,N_46105);
nand U46521 (N_46521,N_46277,N_46059);
xor U46522 (N_46522,N_46297,N_46266);
xnor U46523 (N_46523,N_46222,N_46398);
and U46524 (N_46524,N_46374,N_46465);
nand U46525 (N_46525,N_46185,N_46019);
or U46526 (N_46526,N_46021,N_46128);
xor U46527 (N_46527,N_46125,N_46360);
nor U46528 (N_46528,N_46269,N_46116);
or U46529 (N_46529,N_46134,N_46491);
nand U46530 (N_46530,N_46364,N_46302);
nor U46531 (N_46531,N_46177,N_46475);
nor U46532 (N_46532,N_46400,N_46375);
nor U46533 (N_46533,N_46130,N_46015);
xnor U46534 (N_46534,N_46474,N_46133);
nand U46535 (N_46535,N_46054,N_46168);
and U46536 (N_46536,N_46184,N_46339);
or U46537 (N_46537,N_46340,N_46405);
and U46538 (N_46538,N_46317,N_46182);
and U46539 (N_46539,N_46319,N_46220);
or U46540 (N_46540,N_46187,N_46104);
nand U46541 (N_46541,N_46093,N_46322);
and U46542 (N_46542,N_46395,N_46229);
nand U46543 (N_46543,N_46094,N_46394);
or U46544 (N_46544,N_46068,N_46438);
nor U46545 (N_46545,N_46179,N_46180);
or U46546 (N_46546,N_46321,N_46031);
nand U46547 (N_46547,N_46240,N_46428);
nand U46548 (N_46548,N_46075,N_46310);
or U46549 (N_46549,N_46109,N_46223);
and U46550 (N_46550,N_46020,N_46139);
nor U46551 (N_46551,N_46152,N_46211);
nand U46552 (N_46552,N_46188,N_46431);
nor U46553 (N_46553,N_46047,N_46444);
nand U46554 (N_46554,N_46227,N_46027);
xor U46555 (N_46555,N_46107,N_46189);
nor U46556 (N_46556,N_46231,N_46214);
xnor U46557 (N_46557,N_46305,N_46457);
nand U46558 (N_46558,N_46251,N_46479);
nor U46559 (N_46559,N_46309,N_46076);
nor U46560 (N_46560,N_46241,N_46142);
and U46561 (N_46561,N_46115,N_46124);
nand U46562 (N_46562,N_46417,N_46077);
nor U46563 (N_46563,N_46486,N_46354);
nor U46564 (N_46564,N_46420,N_46329);
or U46565 (N_46565,N_46469,N_46291);
nor U46566 (N_46566,N_46349,N_46070);
nand U46567 (N_46567,N_46034,N_46347);
nand U46568 (N_46568,N_46299,N_46064);
nor U46569 (N_46569,N_46007,N_46055);
nor U46570 (N_46570,N_46278,N_46352);
xor U46571 (N_46571,N_46373,N_46143);
nor U46572 (N_46572,N_46197,N_46101);
and U46573 (N_46573,N_46255,N_46301);
xnor U46574 (N_46574,N_46221,N_46110);
nand U46575 (N_46575,N_46199,N_46216);
and U46576 (N_46576,N_46372,N_46092);
nand U46577 (N_46577,N_46201,N_46242);
xnor U46578 (N_46578,N_46370,N_46281);
nor U46579 (N_46579,N_46228,N_46052);
or U46580 (N_46580,N_46114,N_46451);
and U46581 (N_46581,N_46493,N_46033);
xnor U46582 (N_46582,N_46207,N_46282);
nand U46583 (N_46583,N_46256,N_46244);
xnor U46584 (N_46584,N_46454,N_46106);
nand U46585 (N_46585,N_46144,N_46345);
nand U46586 (N_46586,N_46238,N_46391);
nand U46587 (N_46587,N_46009,N_46045);
and U46588 (N_46588,N_46122,N_46463);
xor U46589 (N_46589,N_46046,N_46293);
nand U46590 (N_46590,N_46334,N_46164);
nand U46591 (N_46591,N_46058,N_46433);
xor U46592 (N_46592,N_46103,N_46169);
and U46593 (N_46593,N_46308,N_46022);
xnor U46594 (N_46594,N_46261,N_46096);
xor U46595 (N_46595,N_46381,N_46191);
or U46596 (N_46596,N_46217,N_46487);
and U46597 (N_46597,N_46167,N_46165);
and U46598 (N_46598,N_46267,N_46421);
or U46599 (N_46599,N_46489,N_46423);
or U46600 (N_46600,N_46225,N_46247);
nor U46601 (N_46601,N_46237,N_46037);
nand U46602 (N_46602,N_46468,N_46275);
nor U46603 (N_46603,N_46082,N_46336);
or U46604 (N_46604,N_46304,N_46215);
xnor U46605 (N_46605,N_46289,N_46212);
or U46606 (N_46606,N_46410,N_46393);
and U46607 (N_46607,N_46138,N_46284);
or U46608 (N_46608,N_46135,N_46378);
nor U46609 (N_46609,N_46018,N_46426);
xnor U46610 (N_46610,N_46265,N_46344);
xnor U46611 (N_46611,N_46436,N_46461);
or U46612 (N_46612,N_46030,N_46292);
or U46613 (N_46613,N_46496,N_46264);
xor U46614 (N_46614,N_46100,N_46362);
or U46615 (N_46615,N_46154,N_46396);
nand U46616 (N_46616,N_46157,N_46147);
nor U46617 (N_46617,N_46063,N_46298);
nand U46618 (N_46618,N_46171,N_46499);
or U46619 (N_46619,N_46091,N_46363);
xnor U46620 (N_46620,N_46482,N_46069);
or U46621 (N_46621,N_46205,N_46392);
or U46622 (N_46622,N_46413,N_46422);
and U46623 (N_46623,N_46198,N_46314);
xor U46624 (N_46624,N_46358,N_46383);
nand U46625 (N_46625,N_46286,N_46271);
and U46626 (N_46626,N_46011,N_46357);
nand U46627 (N_46627,N_46290,N_46161);
nor U46628 (N_46628,N_46209,N_46263);
or U46629 (N_46629,N_46181,N_46361);
nand U46630 (N_46630,N_46006,N_46173);
and U46631 (N_46631,N_46382,N_46126);
nand U46632 (N_46632,N_46306,N_46043);
or U46633 (N_46633,N_46039,N_46324);
nand U46634 (N_46634,N_46248,N_46262);
xnor U46635 (N_46635,N_46353,N_46194);
nand U46636 (N_46636,N_46050,N_46206);
xnor U46637 (N_46637,N_46355,N_46153);
nand U46638 (N_46638,N_46086,N_46095);
and U46639 (N_46639,N_46384,N_46246);
nor U46640 (N_46640,N_46449,N_46366);
and U46641 (N_46641,N_46313,N_46208);
or U46642 (N_46642,N_46236,N_46196);
nand U46643 (N_46643,N_46174,N_46409);
nor U46644 (N_46644,N_46473,N_46008);
nor U46645 (N_46645,N_46272,N_46166);
nor U46646 (N_46646,N_46137,N_46140);
nand U46647 (N_46647,N_46470,N_46253);
nor U46648 (N_46648,N_46003,N_46408);
and U46649 (N_46649,N_46476,N_46178);
xnor U46650 (N_46650,N_46343,N_46478);
nor U46651 (N_46651,N_46480,N_46419);
xnor U46652 (N_46652,N_46071,N_46294);
nand U46653 (N_46653,N_46459,N_46001);
nor U46654 (N_46654,N_46494,N_46123);
xor U46655 (N_46655,N_46234,N_46342);
nor U46656 (N_46656,N_46388,N_46440);
nand U46657 (N_46657,N_46017,N_46471);
and U46658 (N_46658,N_46485,N_46163);
xor U46659 (N_46659,N_46260,N_46159);
nor U46660 (N_46660,N_46283,N_46156);
or U46661 (N_46661,N_46320,N_46028);
or U46662 (N_46662,N_46442,N_46403);
or U46663 (N_46663,N_46333,N_46083);
xor U46664 (N_46664,N_46202,N_46367);
nor U46665 (N_46665,N_46010,N_46330);
nand U46666 (N_46666,N_46040,N_46112);
nand U46667 (N_46667,N_46484,N_46466);
or U46668 (N_46668,N_46233,N_46108);
nor U46669 (N_46669,N_46368,N_46252);
and U46670 (N_46670,N_46318,N_46315);
or U46671 (N_46671,N_46032,N_46439);
or U46672 (N_46672,N_46254,N_46160);
nand U46673 (N_46673,N_46200,N_46356);
xor U46674 (N_46674,N_46190,N_46056);
nand U46675 (N_46675,N_46312,N_46186);
xor U46676 (N_46676,N_46441,N_46285);
nor U46677 (N_46677,N_46016,N_46450);
and U46678 (N_46678,N_46386,N_46287);
nand U46679 (N_46679,N_46193,N_46080);
xor U46680 (N_46680,N_46427,N_46035);
nor U46681 (N_46681,N_46213,N_46183);
and U46682 (N_46682,N_46102,N_46295);
or U46683 (N_46683,N_46057,N_46498);
and U46684 (N_46684,N_46460,N_46404);
nor U46685 (N_46685,N_46131,N_46415);
and U46686 (N_46686,N_46276,N_46337);
or U46687 (N_46687,N_46488,N_46136);
xnor U46688 (N_46688,N_46335,N_46432);
nand U46689 (N_46689,N_46074,N_46430);
and U46690 (N_46690,N_46414,N_46411);
nor U46691 (N_46691,N_46483,N_46210);
xnor U46692 (N_46692,N_46060,N_46418);
or U46693 (N_46693,N_46452,N_46274);
and U46694 (N_46694,N_46141,N_46097);
or U46695 (N_46695,N_46042,N_46397);
or U46696 (N_46696,N_46048,N_46172);
and U46697 (N_46697,N_46280,N_46117);
or U46698 (N_46698,N_46158,N_46025);
xnor U46699 (N_46699,N_46303,N_46495);
or U46700 (N_46700,N_46036,N_46332);
and U46701 (N_46701,N_46296,N_46387);
nor U46702 (N_46702,N_46448,N_46226);
and U46703 (N_46703,N_46085,N_46311);
or U46704 (N_46704,N_46377,N_46079);
or U46705 (N_46705,N_46044,N_46088);
or U46706 (N_46706,N_46389,N_46218);
and U46707 (N_46707,N_46000,N_46149);
xor U46708 (N_46708,N_46446,N_46458);
xor U46709 (N_46709,N_46472,N_46002);
nor U46710 (N_46710,N_46053,N_46155);
xnor U46711 (N_46711,N_46148,N_46204);
nor U46712 (N_46712,N_46369,N_46004);
or U46713 (N_46713,N_46425,N_46453);
or U46714 (N_46714,N_46447,N_46481);
nand U46715 (N_46715,N_46051,N_46327);
nor U46716 (N_46716,N_46073,N_46090);
nor U46717 (N_46717,N_46084,N_46250);
xor U46718 (N_46718,N_46477,N_46127);
xor U46719 (N_46719,N_46257,N_46078);
xnor U46720 (N_46720,N_46029,N_46429);
and U46721 (N_46721,N_46113,N_46111);
nor U46722 (N_46722,N_46325,N_46041);
and U46723 (N_46723,N_46121,N_46402);
xnor U46724 (N_46724,N_46437,N_46145);
xor U46725 (N_46725,N_46239,N_46346);
xnor U46726 (N_46726,N_46376,N_46026);
nor U46727 (N_46727,N_46023,N_46365);
nor U46728 (N_46728,N_46399,N_46279);
and U46729 (N_46729,N_46467,N_46089);
xnor U46730 (N_46730,N_46434,N_46416);
nand U46731 (N_46731,N_46341,N_46435);
xnor U46732 (N_46732,N_46351,N_46492);
nand U46733 (N_46733,N_46338,N_46151);
or U46734 (N_46734,N_46065,N_46098);
nor U46735 (N_46735,N_46464,N_46490);
nor U46736 (N_46736,N_46390,N_46192);
nand U46737 (N_46737,N_46235,N_46081);
nor U46738 (N_46738,N_46456,N_46013);
xnor U46739 (N_46739,N_46049,N_46118);
xnor U46740 (N_46740,N_46129,N_46195);
nor U46741 (N_46741,N_46224,N_46230);
or U46742 (N_46742,N_46412,N_46249);
or U46743 (N_46743,N_46407,N_46119);
xnor U46744 (N_46744,N_46385,N_46268);
nand U46745 (N_46745,N_46061,N_46288);
or U46746 (N_46746,N_46175,N_46176);
xor U46747 (N_46747,N_46424,N_46348);
and U46748 (N_46748,N_46067,N_46300);
and U46749 (N_46749,N_46120,N_46146);
nor U46750 (N_46750,N_46209,N_46321);
xor U46751 (N_46751,N_46132,N_46448);
nor U46752 (N_46752,N_46203,N_46419);
nand U46753 (N_46753,N_46392,N_46449);
nand U46754 (N_46754,N_46431,N_46016);
nor U46755 (N_46755,N_46331,N_46182);
and U46756 (N_46756,N_46250,N_46254);
nor U46757 (N_46757,N_46446,N_46226);
nand U46758 (N_46758,N_46082,N_46144);
and U46759 (N_46759,N_46221,N_46132);
nand U46760 (N_46760,N_46378,N_46357);
nor U46761 (N_46761,N_46199,N_46307);
xnor U46762 (N_46762,N_46107,N_46246);
nor U46763 (N_46763,N_46419,N_46075);
nor U46764 (N_46764,N_46381,N_46285);
xnor U46765 (N_46765,N_46487,N_46374);
nor U46766 (N_46766,N_46090,N_46039);
nand U46767 (N_46767,N_46384,N_46387);
nand U46768 (N_46768,N_46267,N_46088);
xor U46769 (N_46769,N_46038,N_46390);
nand U46770 (N_46770,N_46054,N_46269);
and U46771 (N_46771,N_46452,N_46128);
nand U46772 (N_46772,N_46331,N_46263);
and U46773 (N_46773,N_46363,N_46451);
and U46774 (N_46774,N_46487,N_46020);
nand U46775 (N_46775,N_46398,N_46299);
and U46776 (N_46776,N_46009,N_46428);
nor U46777 (N_46777,N_46340,N_46274);
and U46778 (N_46778,N_46012,N_46074);
nand U46779 (N_46779,N_46218,N_46312);
xor U46780 (N_46780,N_46191,N_46371);
nor U46781 (N_46781,N_46412,N_46043);
or U46782 (N_46782,N_46414,N_46154);
xor U46783 (N_46783,N_46169,N_46439);
xnor U46784 (N_46784,N_46019,N_46428);
xor U46785 (N_46785,N_46137,N_46253);
nor U46786 (N_46786,N_46185,N_46239);
or U46787 (N_46787,N_46104,N_46033);
xnor U46788 (N_46788,N_46265,N_46223);
nand U46789 (N_46789,N_46481,N_46431);
nor U46790 (N_46790,N_46106,N_46025);
xor U46791 (N_46791,N_46059,N_46129);
or U46792 (N_46792,N_46174,N_46434);
xnor U46793 (N_46793,N_46157,N_46180);
and U46794 (N_46794,N_46364,N_46328);
or U46795 (N_46795,N_46296,N_46397);
nand U46796 (N_46796,N_46200,N_46339);
and U46797 (N_46797,N_46141,N_46066);
or U46798 (N_46798,N_46173,N_46489);
xnor U46799 (N_46799,N_46255,N_46030);
nand U46800 (N_46800,N_46265,N_46352);
nand U46801 (N_46801,N_46084,N_46286);
nor U46802 (N_46802,N_46200,N_46016);
nand U46803 (N_46803,N_46168,N_46311);
xnor U46804 (N_46804,N_46392,N_46478);
and U46805 (N_46805,N_46370,N_46293);
xor U46806 (N_46806,N_46238,N_46441);
nor U46807 (N_46807,N_46015,N_46455);
and U46808 (N_46808,N_46119,N_46250);
nor U46809 (N_46809,N_46200,N_46484);
nor U46810 (N_46810,N_46388,N_46180);
and U46811 (N_46811,N_46287,N_46039);
or U46812 (N_46812,N_46228,N_46328);
nand U46813 (N_46813,N_46469,N_46007);
nor U46814 (N_46814,N_46031,N_46407);
nor U46815 (N_46815,N_46437,N_46209);
and U46816 (N_46816,N_46431,N_46216);
xor U46817 (N_46817,N_46098,N_46310);
xor U46818 (N_46818,N_46333,N_46380);
or U46819 (N_46819,N_46125,N_46198);
nand U46820 (N_46820,N_46452,N_46406);
xor U46821 (N_46821,N_46441,N_46350);
nor U46822 (N_46822,N_46050,N_46489);
or U46823 (N_46823,N_46345,N_46302);
or U46824 (N_46824,N_46093,N_46014);
nor U46825 (N_46825,N_46458,N_46276);
nand U46826 (N_46826,N_46106,N_46024);
nand U46827 (N_46827,N_46375,N_46044);
xnor U46828 (N_46828,N_46251,N_46236);
xnor U46829 (N_46829,N_46181,N_46486);
nor U46830 (N_46830,N_46266,N_46180);
nor U46831 (N_46831,N_46358,N_46446);
nand U46832 (N_46832,N_46122,N_46412);
or U46833 (N_46833,N_46146,N_46364);
xnor U46834 (N_46834,N_46382,N_46044);
and U46835 (N_46835,N_46373,N_46052);
nor U46836 (N_46836,N_46341,N_46491);
and U46837 (N_46837,N_46372,N_46183);
nand U46838 (N_46838,N_46214,N_46331);
nor U46839 (N_46839,N_46363,N_46327);
or U46840 (N_46840,N_46334,N_46317);
xor U46841 (N_46841,N_46218,N_46317);
xnor U46842 (N_46842,N_46197,N_46442);
xnor U46843 (N_46843,N_46089,N_46337);
xnor U46844 (N_46844,N_46373,N_46310);
nand U46845 (N_46845,N_46292,N_46143);
xnor U46846 (N_46846,N_46456,N_46137);
nand U46847 (N_46847,N_46087,N_46214);
nand U46848 (N_46848,N_46003,N_46243);
or U46849 (N_46849,N_46453,N_46185);
and U46850 (N_46850,N_46238,N_46047);
or U46851 (N_46851,N_46030,N_46012);
and U46852 (N_46852,N_46005,N_46385);
nor U46853 (N_46853,N_46192,N_46130);
xor U46854 (N_46854,N_46033,N_46198);
and U46855 (N_46855,N_46367,N_46093);
nand U46856 (N_46856,N_46005,N_46395);
or U46857 (N_46857,N_46198,N_46245);
nor U46858 (N_46858,N_46342,N_46064);
nor U46859 (N_46859,N_46294,N_46352);
or U46860 (N_46860,N_46113,N_46264);
or U46861 (N_46861,N_46468,N_46481);
xor U46862 (N_46862,N_46415,N_46073);
and U46863 (N_46863,N_46488,N_46340);
nand U46864 (N_46864,N_46369,N_46230);
xnor U46865 (N_46865,N_46424,N_46421);
and U46866 (N_46866,N_46000,N_46126);
and U46867 (N_46867,N_46336,N_46098);
xor U46868 (N_46868,N_46079,N_46169);
xor U46869 (N_46869,N_46129,N_46302);
nor U46870 (N_46870,N_46163,N_46027);
xor U46871 (N_46871,N_46127,N_46321);
nand U46872 (N_46872,N_46377,N_46010);
and U46873 (N_46873,N_46350,N_46276);
xor U46874 (N_46874,N_46027,N_46206);
nand U46875 (N_46875,N_46472,N_46018);
xnor U46876 (N_46876,N_46286,N_46218);
nand U46877 (N_46877,N_46196,N_46209);
and U46878 (N_46878,N_46328,N_46448);
or U46879 (N_46879,N_46424,N_46142);
nor U46880 (N_46880,N_46292,N_46186);
nand U46881 (N_46881,N_46088,N_46489);
xor U46882 (N_46882,N_46312,N_46277);
and U46883 (N_46883,N_46332,N_46251);
nor U46884 (N_46884,N_46114,N_46013);
and U46885 (N_46885,N_46328,N_46120);
or U46886 (N_46886,N_46391,N_46107);
or U46887 (N_46887,N_46327,N_46003);
nand U46888 (N_46888,N_46198,N_46405);
or U46889 (N_46889,N_46081,N_46208);
xor U46890 (N_46890,N_46412,N_46044);
nand U46891 (N_46891,N_46135,N_46367);
or U46892 (N_46892,N_46359,N_46476);
and U46893 (N_46893,N_46273,N_46338);
xor U46894 (N_46894,N_46016,N_46190);
nand U46895 (N_46895,N_46390,N_46077);
or U46896 (N_46896,N_46244,N_46482);
nor U46897 (N_46897,N_46261,N_46459);
nand U46898 (N_46898,N_46404,N_46060);
nor U46899 (N_46899,N_46223,N_46396);
nand U46900 (N_46900,N_46061,N_46474);
and U46901 (N_46901,N_46222,N_46254);
nand U46902 (N_46902,N_46409,N_46009);
and U46903 (N_46903,N_46184,N_46342);
xnor U46904 (N_46904,N_46116,N_46257);
xor U46905 (N_46905,N_46447,N_46361);
nand U46906 (N_46906,N_46461,N_46069);
or U46907 (N_46907,N_46313,N_46388);
or U46908 (N_46908,N_46351,N_46016);
and U46909 (N_46909,N_46233,N_46322);
nand U46910 (N_46910,N_46311,N_46015);
and U46911 (N_46911,N_46303,N_46219);
or U46912 (N_46912,N_46265,N_46382);
or U46913 (N_46913,N_46435,N_46169);
or U46914 (N_46914,N_46179,N_46146);
xnor U46915 (N_46915,N_46317,N_46189);
and U46916 (N_46916,N_46159,N_46282);
nand U46917 (N_46917,N_46479,N_46191);
and U46918 (N_46918,N_46101,N_46170);
and U46919 (N_46919,N_46204,N_46055);
nand U46920 (N_46920,N_46209,N_46486);
nand U46921 (N_46921,N_46124,N_46154);
and U46922 (N_46922,N_46421,N_46347);
nor U46923 (N_46923,N_46434,N_46162);
nand U46924 (N_46924,N_46105,N_46000);
or U46925 (N_46925,N_46115,N_46269);
nor U46926 (N_46926,N_46159,N_46477);
nand U46927 (N_46927,N_46040,N_46383);
nand U46928 (N_46928,N_46318,N_46323);
or U46929 (N_46929,N_46101,N_46254);
and U46930 (N_46930,N_46227,N_46203);
and U46931 (N_46931,N_46320,N_46472);
nor U46932 (N_46932,N_46009,N_46308);
nand U46933 (N_46933,N_46210,N_46413);
nor U46934 (N_46934,N_46163,N_46494);
xor U46935 (N_46935,N_46459,N_46009);
or U46936 (N_46936,N_46312,N_46012);
xor U46937 (N_46937,N_46176,N_46277);
nand U46938 (N_46938,N_46407,N_46132);
xnor U46939 (N_46939,N_46417,N_46423);
xor U46940 (N_46940,N_46291,N_46446);
xnor U46941 (N_46941,N_46275,N_46238);
and U46942 (N_46942,N_46314,N_46276);
nand U46943 (N_46943,N_46402,N_46021);
and U46944 (N_46944,N_46102,N_46199);
xor U46945 (N_46945,N_46046,N_46199);
and U46946 (N_46946,N_46479,N_46077);
nand U46947 (N_46947,N_46220,N_46154);
xor U46948 (N_46948,N_46244,N_46309);
nor U46949 (N_46949,N_46015,N_46105);
or U46950 (N_46950,N_46340,N_46389);
nor U46951 (N_46951,N_46099,N_46310);
and U46952 (N_46952,N_46430,N_46291);
xnor U46953 (N_46953,N_46422,N_46374);
and U46954 (N_46954,N_46287,N_46053);
nor U46955 (N_46955,N_46404,N_46063);
xnor U46956 (N_46956,N_46369,N_46423);
nand U46957 (N_46957,N_46098,N_46035);
and U46958 (N_46958,N_46070,N_46364);
nand U46959 (N_46959,N_46107,N_46167);
and U46960 (N_46960,N_46249,N_46197);
nor U46961 (N_46961,N_46287,N_46276);
nor U46962 (N_46962,N_46195,N_46345);
or U46963 (N_46963,N_46124,N_46067);
or U46964 (N_46964,N_46417,N_46114);
xor U46965 (N_46965,N_46173,N_46432);
nor U46966 (N_46966,N_46365,N_46435);
and U46967 (N_46967,N_46327,N_46446);
nor U46968 (N_46968,N_46220,N_46473);
xnor U46969 (N_46969,N_46189,N_46208);
nand U46970 (N_46970,N_46109,N_46473);
nor U46971 (N_46971,N_46411,N_46320);
xor U46972 (N_46972,N_46474,N_46433);
and U46973 (N_46973,N_46155,N_46045);
or U46974 (N_46974,N_46059,N_46209);
and U46975 (N_46975,N_46431,N_46066);
xor U46976 (N_46976,N_46367,N_46186);
and U46977 (N_46977,N_46447,N_46263);
or U46978 (N_46978,N_46299,N_46244);
nand U46979 (N_46979,N_46464,N_46406);
and U46980 (N_46980,N_46354,N_46436);
nor U46981 (N_46981,N_46281,N_46294);
and U46982 (N_46982,N_46444,N_46390);
or U46983 (N_46983,N_46000,N_46351);
and U46984 (N_46984,N_46497,N_46087);
nand U46985 (N_46985,N_46182,N_46202);
xnor U46986 (N_46986,N_46203,N_46199);
and U46987 (N_46987,N_46139,N_46224);
and U46988 (N_46988,N_46485,N_46220);
nand U46989 (N_46989,N_46119,N_46155);
xor U46990 (N_46990,N_46309,N_46166);
nor U46991 (N_46991,N_46471,N_46463);
xnor U46992 (N_46992,N_46043,N_46343);
nor U46993 (N_46993,N_46470,N_46047);
xnor U46994 (N_46994,N_46386,N_46350);
and U46995 (N_46995,N_46495,N_46048);
nand U46996 (N_46996,N_46095,N_46470);
nand U46997 (N_46997,N_46317,N_46256);
xor U46998 (N_46998,N_46403,N_46259);
and U46999 (N_46999,N_46383,N_46072);
xor U47000 (N_47000,N_46655,N_46527);
xnor U47001 (N_47001,N_46604,N_46873);
or U47002 (N_47002,N_46832,N_46552);
xor U47003 (N_47003,N_46553,N_46710);
and U47004 (N_47004,N_46607,N_46917);
nor U47005 (N_47005,N_46722,N_46922);
nor U47006 (N_47006,N_46714,N_46538);
nand U47007 (N_47007,N_46747,N_46926);
or U47008 (N_47008,N_46988,N_46773);
xor U47009 (N_47009,N_46909,N_46811);
or U47010 (N_47010,N_46690,N_46588);
or U47011 (N_47011,N_46903,N_46709);
and U47012 (N_47012,N_46776,N_46644);
nand U47013 (N_47013,N_46693,N_46591);
nand U47014 (N_47014,N_46931,N_46763);
and U47015 (N_47015,N_46646,N_46558);
and U47016 (N_47016,N_46682,N_46566);
nor U47017 (N_47017,N_46636,N_46534);
nand U47018 (N_47018,N_46716,N_46501);
and U47019 (N_47019,N_46904,N_46984);
xor U47020 (N_47020,N_46932,N_46828);
nand U47021 (N_47021,N_46741,N_46844);
or U47022 (N_47022,N_46820,N_46704);
nor U47023 (N_47023,N_46898,N_46833);
nand U47024 (N_47024,N_46895,N_46748);
nand U47025 (N_47025,N_46500,N_46826);
xor U47026 (N_47026,N_46575,N_46940);
or U47027 (N_47027,N_46729,N_46994);
and U47028 (N_47028,N_46517,N_46881);
nand U47029 (N_47029,N_46705,N_46692);
nand U47030 (N_47030,N_46869,N_46681);
xor U47031 (N_47031,N_46595,N_46952);
nor U47032 (N_47032,N_46698,N_46831);
xor U47033 (N_47033,N_46562,N_46995);
nor U47034 (N_47034,N_46887,N_46980);
xnor U47035 (N_47035,N_46613,N_46586);
nor U47036 (N_47036,N_46505,N_46579);
xor U47037 (N_47037,N_46711,N_46884);
nor U47038 (N_47038,N_46663,N_46933);
and U47039 (N_47039,N_46805,N_46576);
nor U47040 (N_47040,N_46949,N_46719);
xnor U47041 (N_47041,N_46790,N_46648);
or U47042 (N_47042,N_46982,N_46539);
nand U47043 (N_47043,N_46674,N_46945);
and U47044 (N_47044,N_46676,N_46985);
nor U47045 (N_47045,N_46807,N_46894);
or U47046 (N_47046,N_46574,N_46630);
xnor U47047 (N_47047,N_46866,N_46863);
and U47048 (N_47048,N_46715,N_46752);
nand U47049 (N_47049,N_46612,N_46855);
and U47050 (N_47050,N_46789,N_46649);
nand U47051 (N_47051,N_46919,N_46787);
xor U47052 (N_47052,N_46685,N_46783);
xnor U47053 (N_47053,N_46925,N_46876);
xnor U47054 (N_47054,N_46930,N_46688);
and U47055 (N_47055,N_46993,N_46978);
nand U47056 (N_47056,N_46969,N_46587);
xnor U47057 (N_47057,N_46590,N_46572);
xnor U47058 (N_47058,N_46986,N_46975);
or U47059 (N_47059,N_46700,N_46583);
xnor U47060 (N_47060,N_46998,N_46751);
nand U47061 (N_47061,N_46843,N_46542);
xor U47062 (N_47062,N_46921,N_46816);
xor U47063 (N_47063,N_46684,N_46502);
or U47064 (N_47064,N_46775,N_46707);
and U47065 (N_47065,N_46537,N_46554);
nand U47066 (N_47066,N_46860,N_46778);
and U47067 (N_47067,N_46717,N_46523);
nand U47068 (N_47068,N_46964,N_46788);
or U47069 (N_47069,N_46525,N_46724);
xnor U47070 (N_47070,N_46518,N_46971);
xnor U47071 (N_47071,N_46600,N_46912);
and U47072 (N_47072,N_46515,N_46829);
nor U47073 (N_47073,N_46699,N_46734);
and U47074 (N_47074,N_46520,N_46943);
nand U47075 (N_47075,N_46670,N_46508);
xnor U47076 (N_47076,N_46606,N_46611);
xor U47077 (N_47077,N_46581,N_46896);
nor U47078 (N_47078,N_46666,N_46742);
and U47079 (N_47079,N_46506,N_46678);
or U47080 (N_47080,N_46673,N_46963);
nand U47081 (N_47081,N_46610,N_46871);
xor U47082 (N_47082,N_46792,N_46797);
nor U47083 (N_47083,N_46750,N_46849);
and U47084 (N_47084,N_46765,N_46910);
nor U47085 (N_47085,N_46735,N_46937);
nand U47086 (N_47086,N_46578,N_46555);
nand U47087 (N_47087,N_46745,N_46882);
nand U47088 (N_47088,N_46946,N_46640);
nor U47089 (N_47089,N_46777,N_46879);
nor U47090 (N_47090,N_46927,N_46740);
nand U47091 (N_47091,N_46598,N_46997);
nand U47092 (N_47092,N_46989,N_46565);
or U47093 (N_47093,N_46771,N_46924);
and U47094 (N_47094,N_46758,N_46799);
nand U47095 (N_47095,N_46850,N_46618);
and U47096 (N_47096,N_46535,N_46979);
xnor U47097 (N_47097,N_46633,N_46880);
nand U47098 (N_47098,N_46512,N_46614);
and U47099 (N_47099,N_46522,N_46920);
nor U47100 (N_47100,N_46677,N_46712);
nor U47101 (N_47101,N_46804,N_46838);
or U47102 (N_47102,N_46760,N_46645);
or U47103 (N_47103,N_46701,N_46802);
and U47104 (N_47104,N_46647,N_46798);
nand U47105 (N_47105,N_46872,N_46749);
or U47106 (N_47106,N_46540,N_46793);
nand U47107 (N_47107,N_46511,N_46594);
nand U47108 (N_47108,N_46658,N_46835);
and U47109 (N_47109,N_46996,N_46801);
nand U47110 (N_47110,N_46603,N_46687);
nand U47111 (N_47111,N_46827,N_46652);
or U47112 (N_47112,N_46597,N_46947);
nand U47113 (N_47113,N_46956,N_46948);
and U47114 (N_47114,N_46780,N_46503);
nor U47115 (N_47115,N_46533,N_46786);
and U47116 (N_47116,N_46839,N_46509);
and U47117 (N_47117,N_46563,N_46635);
nor U47118 (N_47118,N_46974,N_46695);
nor U47119 (N_47119,N_46864,N_46756);
nor U47120 (N_47120,N_46738,N_46661);
and U47121 (N_47121,N_46638,N_46836);
and U47122 (N_47122,N_46718,N_46764);
xnor U47123 (N_47123,N_46962,N_46950);
or U47124 (N_47124,N_46939,N_46733);
or U47125 (N_47125,N_46991,N_46754);
or U47126 (N_47126,N_46886,N_46601);
xor U47127 (N_47127,N_46620,N_46817);
nor U47128 (N_47128,N_46551,N_46965);
or U47129 (N_47129,N_46852,N_46592);
and U47130 (N_47130,N_46548,N_46672);
nor U47131 (N_47131,N_46885,N_46809);
xnor U47132 (N_47132,N_46893,N_46696);
nand U47133 (N_47133,N_46840,N_46536);
or U47134 (N_47134,N_46821,N_46642);
and U47135 (N_47135,N_46890,N_46936);
or U47136 (N_47136,N_46743,N_46957);
and U47137 (N_47137,N_46570,N_46641);
nor U47138 (N_47138,N_46941,N_46627);
nand U47139 (N_47139,N_46524,N_46862);
and U47140 (N_47140,N_46605,N_46589);
xnor U47141 (N_47141,N_46766,N_46813);
or U47142 (N_47142,N_46637,N_46761);
xnor U47143 (N_47143,N_46883,N_46823);
and U47144 (N_47144,N_46732,N_46713);
xnor U47145 (N_47145,N_46739,N_46772);
xor U47146 (N_47146,N_46526,N_46585);
nand U47147 (N_47147,N_46731,N_46992);
or U47148 (N_47148,N_46608,N_46720);
nor U47149 (N_47149,N_46609,N_46617);
or U47150 (N_47150,N_46762,N_46858);
or U47151 (N_47151,N_46721,N_46582);
nand U47152 (N_47152,N_46999,N_46504);
nand U47153 (N_47153,N_46623,N_46569);
or U47154 (N_47154,N_46942,N_46725);
nor U47155 (N_47155,N_46665,N_46657);
xnor U47156 (N_47156,N_46727,N_46878);
xnor U47157 (N_47157,N_46822,N_46529);
and U47158 (N_47158,N_46769,N_46651);
or U47159 (N_47159,N_46908,N_46867);
and U47160 (N_47160,N_46532,N_46768);
xnor U47161 (N_47161,N_46755,N_46889);
or U47162 (N_47162,N_46955,N_46865);
nor U47163 (N_47163,N_46736,N_46825);
or U47164 (N_47164,N_46779,N_46848);
and U47165 (N_47165,N_46958,N_46934);
nand U47166 (N_47166,N_46892,N_46653);
xnor U47167 (N_47167,N_46976,N_46691);
xnor U47168 (N_47168,N_46702,N_46824);
nor U47169 (N_47169,N_46906,N_46888);
and U47170 (N_47170,N_46803,N_46819);
nand U47171 (N_47171,N_46519,N_46560);
and U47172 (N_47172,N_46530,N_46853);
and U47173 (N_47173,N_46703,N_46983);
or U47174 (N_47174,N_46679,N_46818);
nor U47175 (N_47175,N_46774,N_46513);
and U47176 (N_47176,N_46669,N_46531);
nor U47177 (N_47177,N_46697,N_46784);
xor U47178 (N_47178,N_46664,N_46546);
and U47179 (N_47179,N_46854,N_46730);
nor U47180 (N_47180,N_46668,N_46660);
nand U47181 (N_47181,N_46859,N_46877);
nand U47182 (N_47182,N_46624,N_46913);
and U47183 (N_47183,N_46808,N_46510);
or U47184 (N_47184,N_46874,N_46683);
nand U47185 (N_47185,N_46905,N_46621);
and U47186 (N_47186,N_46899,N_46935);
and U47187 (N_47187,N_46796,N_46686);
nor U47188 (N_47188,N_46851,N_46845);
and U47189 (N_47189,N_46954,N_46753);
or U47190 (N_47190,N_46631,N_46770);
xnor U47191 (N_47191,N_46516,N_46841);
and U47192 (N_47192,N_46857,N_46966);
xnor U47193 (N_47193,N_46973,N_46911);
nor U47194 (N_47194,N_46907,N_46923);
nand U47195 (N_47195,N_46781,N_46891);
nor U47196 (N_47196,N_46616,N_46619);
or U47197 (N_47197,N_46547,N_46806);
nor U47198 (N_47198,N_46671,N_46938);
nand U47199 (N_47199,N_46708,N_46737);
nor U47200 (N_47200,N_46643,N_46902);
xor U47201 (N_47201,N_46556,N_46970);
xnor U47202 (N_47202,N_46521,N_46659);
xor U47203 (N_47203,N_46628,N_46901);
and U47204 (N_47204,N_46568,N_46959);
or U47205 (N_47205,N_46689,N_46814);
and U47206 (N_47206,N_46990,N_46667);
nor U47207 (N_47207,N_46928,N_46830);
nand U47208 (N_47208,N_46596,N_46650);
or U47209 (N_47209,N_46767,N_46654);
nand U47210 (N_47210,N_46856,N_46514);
nand U47211 (N_47211,N_46929,N_46744);
xor U47212 (N_47212,N_46875,N_46625);
xor U47213 (N_47213,N_46918,N_46593);
and U47214 (N_47214,N_46639,N_46549);
and U47215 (N_47215,N_46837,N_46916);
nand U47216 (N_47216,N_46599,N_46580);
xor U47217 (N_47217,N_46800,N_46567);
nand U47218 (N_47218,N_46951,N_46757);
or U47219 (N_47219,N_46626,N_46812);
and U47220 (N_47220,N_46561,N_46987);
xnor U47221 (N_47221,N_46541,N_46810);
nand U47222 (N_47222,N_46915,N_46632);
nor U47223 (N_47223,N_46694,N_46944);
nor U47224 (N_47224,N_46573,N_46615);
and U47225 (N_47225,N_46634,N_46543);
xnor U47226 (N_47226,N_46782,N_46981);
nor U47227 (N_47227,N_46953,N_46960);
nand U47228 (N_47228,N_46544,N_46584);
and U47229 (N_47229,N_46728,N_46868);
nand U47230 (N_47230,N_46967,N_46550);
and U47231 (N_47231,N_46785,N_46870);
and U47232 (N_47232,N_46706,N_46629);
or U47233 (N_47233,N_46795,N_46680);
nand U47234 (N_47234,N_46847,N_46746);
nor U47235 (N_47235,N_46972,N_46723);
xor U47236 (N_47236,N_46791,N_46897);
xnor U47237 (N_47237,N_46622,N_46571);
or U47238 (N_47238,N_46759,N_46577);
or U47239 (N_47239,N_46846,N_46961);
and U47240 (N_47240,N_46557,N_46602);
and U47241 (N_47241,N_46675,N_46507);
and U47242 (N_47242,N_46834,N_46815);
xnor U47243 (N_47243,N_46545,N_46559);
and U47244 (N_47244,N_46794,N_46861);
nand U47245 (N_47245,N_46914,N_46656);
or U47246 (N_47246,N_46726,N_46842);
and U47247 (N_47247,N_46968,N_46977);
nor U47248 (N_47248,N_46564,N_46528);
or U47249 (N_47249,N_46662,N_46900);
and U47250 (N_47250,N_46907,N_46620);
or U47251 (N_47251,N_46943,N_46774);
xor U47252 (N_47252,N_46923,N_46819);
and U47253 (N_47253,N_46605,N_46606);
or U47254 (N_47254,N_46653,N_46529);
nor U47255 (N_47255,N_46757,N_46675);
nand U47256 (N_47256,N_46813,N_46861);
or U47257 (N_47257,N_46971,N_46873);
nand U47258 (N_47258,N_46993,N_46534);
or U47259 (N_47259,N_46648,N_46609);
or U47260 (N_47260,N_46564,N_46906);
xor U47261 (N_47261,N_46695,N_46658);
nand U47262 (N_47262,N_46869,N_46901);
and U47263 (N_47263,N_46518,N_46750);
and U47264 (N_47264,N_46504,N_46600);
and U47265 (N_47265,N_46822,N_46921);
nor U47266 (N_47266,N_46501,N_46901);
and U47267 (N_47267,N_46839,N_46785);
or U47268 (N_47268,N_46758,N_46855);
and U47269 (N_47269,N_46744,N_46772);
nand U47270 (N_47270,N_46787,N_46873);
xor U47271 (N_47271,N_46720,N_46501);
nand U47272 (N_47272,N_46702,N_46563);
and U47273 (N_47273,N_46820,N_46594);
nor U47274 (N_47274,N_46989,N_46983);
xor U47275 (N_47275,N_46700,N_46784);
nor U47276 (N_47276,N_46907,N_46555);
nor U47277 (N_47277,N_46952,N_46503);
and U47278 (N_47278,N_46640,N_46567);
xnor U47279 (N_47279,N_46989,N_46708);
or U47280 (N_47280,N_46585,N_46755);
nor U47281 (N_47281,N_46713,N_46679);
nor U47282 (N_47282,N_46966,N_46892);
nand U47283 (N_47283,N_46834,N_46536);
xnor U47284 (N_47284,N_46569,N_46955);
or U47285 (N_47285,N_46908,N_46822);
and U47286 (N_47286,N_46955,N_46585);
nor U47287 (N_47287,N_46901,N_46896);
nor U47288 (N_47288,N_46745,N_46822);
or U47289 (N_47289,N_46565,N_46587);
nor U47290 (N_47290,N_46853,N_46519);
nor U47291 (N_47291,N_46914,N_46803);
nand U47292 (N_47292,N_46581,N_46739);
nor U47293 (N_47293,N_46851,N_46673);
xor U47294 (N_47294,N_46849,N_46579);
xnor U47295 (N_47295,N_46614,N_46924);
xor U47296 (N_47296,N_46513,N_46627);
or U47297 (N_47297,N_46717,N_46781);
xnor U47298 (N_47298,N_46569,N_46943);
or U47299 (N_47299,N_46600,N_46784);
and U47300 (N_47300,N_46902,N_46801);
and U47301 (N_47301,N_46890,N_46548);
nand U47302 (N_47302,N_46611,N_46729);
nor U47303 (N_47303,N_46504,N_46709);
or U47304 (N_47304,N_46725,N_46829);
or U47305 (N_47305,N_46709,N_46888);
or U47306 (N_47306,N_46555,N_46707);
xor U47307 (N_47307,N_46583,N_46627);
or U47308 (N_47308,N_46826,N_46694);
nor U47309 (N_47309,N_46519,N_46931);
or U47310 (N_47310,N_46986,N_46878);
and U47311 (N_47311,N_46671,N_46603);
or U47312 (N_47312,N_46900,N_46965);
and U47313 (N_47313,N_46975,N_46600);
nand U47314 (N_47314,N_46546,N_46589);
xnor U47315 (N_47315,N_46621,N_46551);
nor U47316 (N_47316,N_46784,N_46548);
xor U47317 (N_47317,N_46648,N_46589);
nand U47318 (N_47318,N_46883,N_46975);
or U47319 (N_47319,N_46662,N_46780);
xnor U47320 (N_47320,N_46677,N_46817);
and U47321 (N_47321,N_46958,N_46576);
xor U47322 (N_47322,N_46808,N_46600);
nand U47323 (N_47323,N_46883,N_46756);
nand U47324 (N_47324,N_46631,N_46873);
or U47325 (N_47325,N_46791,N_46542);
nor U47326 (N_47326,N_46649,N_46612);
nor U47327 (N_47327,N_46509,N_46737);
nor U47328 (N_47328,N_46605,N_46905);
xor U47329 (N_47329,N_46615,N_46707);
xor U47330 (N_47330,N_46654,N_46649);
nor U47331 (N_47331,N_46503,N_46837);
xnor U47332 (N_47332,N_46790,N_46904);
nand U47333 (N_47333,N_46559,N_46595);
and U47334 (N_47334,N_46689,N_46596);
nor U47335 (N_47335,N_46958,N_46638);
nor U47336 (N_47336,N_46930,N_46823);
nand U47337 (N_47337,N_46579,N_46768);
nor U47338 (N_47338,N_46638,N_46553);
nor U47339 (N_47339,N_46822,N_46675);
or U47340 (N_47340,N_46896,N_46591);
nor U47341 (N_47341,N_46730,N_46835);
and U47342 (N_47342,N_46740,N_46938);
nand U47343 (N_47343,N_46757,N_46623);
nor U47344 (N_47344,N_46590,N_46693);
nand U47345 (N_47345,N_46992,N_46979);
xnor U47346 (N_47346,N_46780,N_46793);
or U47347 (N_47347,N_46659,N_46629);
xnor U47348 (N_47348,N_46844,N_46631);
xor U47349 (N_47349,N_46803,N_46705);
nand U47350 (N_47350,N_46657,N_46581);
nor U47351 (N_47351,N_46707,N_46534);
xnor U47352 (N_47352,N_46624,N_46816);
and U47353 (N_47353,N_46895,N_46887);
nor U47354 (N_47354,N_46984,N_46977);
and U47355 (N_47355,N_46979,N_46784);
xnor U47356 (N_47356,N_46635,N_46862);
xor U47357 (N_47357,N_46742,N_46502);
or U47358 (N_47358,N_46659,N_46731);
nand U47359 (N_47359,N_46912,N_46900);
nand U47360 (N_47360,N_46594,N_46848);
or U47361 (N_47361,N_46780,N_46774);
nand U47362 (N_47362,N_46598,N_46531);
and U47363 (N_47363,N_46546,N_46929);
xnor U47364 (N_47364,N_46729,N_46620);
nor U47365 (N_47365,N_46999,N_46629);
nor U47366 (N_47366,N_46965,N_46749);
xor U47367 (N_47367,N_46996,N_46672);
or U47368 (N_47368,N_46756,N_46830);
or U47369 (N_47369,N_46962,N_46716);
nor U47370 (N_47370,N_46708,N_46576);
and U47371 (N_47371,N_46522,N_46759);
nand U47372 (N_47372,N_46604,N_46516);
nand U47373 (N_47373,N_46526,N_46582);
nand U47374 (N_47374,N_46714,N_46606);
or U47375 (N_47375,N_46764,N_46512);
or U47376 (N_47376,N_46667,N_46702);
or U47377 (N_47377,N_46787,N_46992);
nor U47378 (N_47378,N_46514,N_46645);
nor U47379 (N_47379,N_46933,N_46523);
nor U47380 (N_47380,N_46875,N_46879);
or U47381 (N_47381,N_46833,N_46687);
xor U47382 (N_47382,N_46764,N_46678);
nand U47383 (N_47383,N_46819,N_46935);
and U47384 (N_47384,N_46541,N_46607);
and U47385 (N_47385,N_46932,N_46553);
xor U47386 (N_47386,N_46612,N_46852);
or U47387 (N_47387,N_46822,N_46757);
nand U47388 (N_47388,N_46607,N_46888);
and U47389 (N_47389,N_46539,N_46709);
nand U47390 (N_47390,N_46822,N_46591);
nand U47391 (N_47391,N_46785,N_46631);
xnor U47392 (N_47392,N_46766,N_46524);
nor U47393 (N_47393,N_46593,N_46842);
xnor U47394 (N_47394,N_46658,N_46801);
nand U47395 (N_47395,N_46962,N_46867);
nand U47396 (N_47396,N_46536,N_46705);
xnor U47397 (N_47397,N_46558,N_46962);
nor U47398 (N_47398,N_46757,N_46805);
xnor U47399 (N_47399,N_46595,N_46695);
and U47400 (N_47400,N_46987,N_46618);
xnor U47401 (N_47401,N_46649,N_46524);
xnor U47402 (N_47402,N_46930,N_46754);
and U47403 (N_47403,N_46593,N_46689);
and U47404 (N_47404,N_46849,N_46537);
or U47405 (N_47405,N_46929,N_46548);
or U47406 (N_47406,N_46951,N_46621);
xnor U47407 (N_47407,N_46744,N_46813);
or U47408 (N_47408,N_46943,N_46804);
or U47409 (N_47409,N_46924,N_46581);
and U47410 (N_47410,N_46969,N_46596);
or U47411 (N_47411,N_46811,N_46728);
xnor U47412 (N_47412,N_46791,N_46506);
nor U47413 (N_47413,N_46723,N_46902);
xor U47414 (N_47414,N_46687,N_46908);
nor U47415 (N_47415,N_46881,N_46803);
nor U47416 (N_47416,N_46760,N_46742);
nor U47417 (N_47417,N_46809,N_46584);
xor U47418 (N_47418,N_46738,N_46663);
or U47419 (N_47419,N_46870,N_46854);
and U47420 (N_47420,N_46976,N_46626);
nand U47421 (N_47421,N_46609,N_46606);
nand U47422 (N_47422,N_46580,N_46629);
xnor U47423 (N_47423,N_46921,N_46843);
xor U47424 (N_47424,N_46798,N_46612);
xnor U47425 (N_47425,N_46871,N_46663);
and U47426 (N_47426,N_46721,N_46812);
and U47427 (N_47427,N_46527,N_46594);
or U47428 (N_47428,N_46993,N_46804);
and U47429 (N_47429,N_46518,N_46527);
or U47430 (N_47430,N_46680,N_46630);
or U47431 (N_47431,N_46553,N_46967);
nand U47432 (N_47432,N_46840,N_46675);
and U47433 (N_47433,N_46521,N_46542);
and U47434 (N_47434,N_46975,N_46806);
and U47435 (N_47435,N_46870,N_46889);
and U47436 (N_47436,N_46564,N_46900);
or U47437 (N_47437,N_46631,N_46687);
nor U47438 (N_47438,N_46857,N_46973);
xnor U47439 (N_47439,N_46862,N_46565);
nand U47440 (N_47440,N_46899,N_46726);
or U47441 (N_47441,N_46793,N_46897);
or U47442 (N_47442,N_46509,N_46592);
nor U47443 (N_47443,N_46851,N_46912);
and U47444 (N_47444,N_46573,N_46744);
or U47445 (N_47445,N_46720,N_46507);
nor U47446 (N_47446,N_46523,N_46886);
and U47447 (N_47447,N_46608,N_46777);
nor U47448 (N_47448,N_46583,N_46567);
nand U47449 (N_47449,N_46950,N_46739);
xor U47450 (N_47450,N_46623,N_46975);
and U47451 (N_47451,N_46593,N_46501);
nand U47452 (N_47452,N_46504,N_46907);
xnor U47453 (N_47453,N_46641,N_46569);
xor U47454 (N_47454,N_46673,N_46764);
or U47455 (N_47455,N_46800,N_46526);
nand U47456 (N_47456,N_46792,N_46559);
xnor U47457 (N_47457,N_46568,N_46596);
and U47458 (N_47458,N_46811,N_46759);
and U47459 (N_47459,N_46782,N_46693);
or U47460 (N_47460,N_46769,N_46952);
nor U47461 (N_47461,N_46551,N_46601);
xor U47462 (N_47462,N_46517,N_46683);
and U47463 (N_47463,N_46842,N_46924);
nand U47464 (N_47464,N_46852,N_46814);
or U47465 (N_47465,N_46841,N_46793);
xor U47466 (N_47466,N_46593,N_46711);
and U47467 (N_47467,N_46737,N_46504);
or U47468 (N_47468,N_46970,N_46830);
or U47469 (N_47469,N_46629,N_46600);
or U47470 (N_47470,N_46611,N_46643);
xor U47471 (N_47471,N_46735,N_46763);
xnor U47472 (N_47472,N_46945,N_46973);
nor U47473 (N_47473,N_46819,N_46978);
nand U47474 (N_47474,N_46734,N_46576);
nand U47475 (N_47475,N_46641,N_46961);
nand U47476 (N_47476,N_46947,N_46669);
nand U47477 (N_47477,N_46689,N_46647);
or U47478 (N_47478,N_46858,N_46709);
xnor U47479 (N_47479,N_46913,N_46570);
and U47480 (N_47480,N_46718,N_46975);
or U47481 (N_47481,N_46954,N_46604);
or U47482 (N_47482,N_46721,N_46758);
and U47483 (N_47483,N_46573,N_46790);
nor U47484 (N_47484,N_46704,N_46835);
nor U47485 (N_47485,N_46902,N_46638);
and U47486 (N_47486,N_46500,N_46750);
or U47487 (N_47487,N_46569,N_46780);
and U47488 (N_47488,N_46909,N_46748);
and U47489 (N_47489,N_46681,N_46964);
nor U47490 (N_47490,N_46934,N_46756);
xnor U47491 (N_47491,N_46618,N_46939);
nand U47492 (N_47492,N_46708,N_46695);
nor U47493 (N_47493,N_46543,N_46599);
or U47494 (N_47494,N_46600,N_46943);
nand U47495 (N_47495,N_46552,N_46913);
nand U47496 (N_47496,N_46708,N_46828);
nand U47497 (N_47497,N_46764,N_46750);
xor U47498 (N_47498,N_46664,N_46881);
nand U47499 (N_47499,N_46705,N_46961);
nand U47500 (N_47500,N_47484,N_47110);
or U47501 (N_47501,N_47023,N_47364);
and U47502 (N_47502,N_47374,N_47320);
nor U47503 (N_47503,N_47013,N_47306);
and U47504 (N_47504,N_47047,N_47359);
xnor U47505 (N_47505,N_47065,N_47379);
and U47506 (N_47506,N_47000,N_47020);
nand U47507 (N_47507,N_47042,N_47446);
nor U47508 (N_47508,N_47471,N_47436);
xor U47509 (N_47509,N_47039,N_47086);
nor U47510 (N_47510,N_47355,N_47369);
nand U47511 (N_47511,N_47327,N_47267);
and U47512 (N_47512,N_47053,N_47283);
nor U47513 (N_47513,N_47356,N_47411);
xor U47514 (N_47514,N_47277,N_47015);
nor U47515 (N_47515,N_47068,N_47498);
nand U47516 (N_47516,N_47298,N_47290);
xnor U47517 (N_47517,N_47438,N_47129);
xor U47518 (N_47518,N_47170,N_47222);
or U47519 (N_47519,N_47105,N_47066);
or U47520 (N_47520,N_47303,N_47198);
or U47521 (N_47521,N_47242,N_47445);
or U47522 (N_47522,N_47333,N_47378);
xnor U47523 (N_47523,N_47331,N_47187);
xnor U47524 (N_47524,N_47005,N_47370);
nand U47525 (N_47525,N_47224,N_47135);
or U47526 (N_47526,N_47447,N_47177);
nand U47527 (N_47527,N_47432,N_47060);
or U47528 (N_47528,N_47365,N_47274);
nand U47529 (N_47529,N_47402,N_47231);
xor U47530 (N_47530,N_47159,N_47300);
or U47531 (N_47531,N_47328,N_47263);
nand U47532 (N_47532,N_47044,N_47315);
nand U47533 (N_47533,N_47128,N_47470);
or U47534 (N_47534,N_47146,N_47190);
and U47535 (N_47535,N_47030,N_47323);
nor U47536 (N_47536,N_47390,N_47246);
or U47537 (N_47537,N_47382,N_47499);
xnor U47538 (N_47538,N_47305,N_47257);
nand U47539 (N_47539,N_47206,N_47161);
or U47540 (N_47540,N_47069,N_47118);
or U47541 (N_47541,N_47318,N_47237);
and U47542 (N_47542,N_47473,N_47130);
xnor U47543 (N_47543,N_47137,N_47405);
xnor U47544 (N_47544,N_47122,N_47464);
or U47545 (N_47545,N_47310,N_47002);
xor U47546 (N_47546,N_47099,N_47183);
nor U47547 (N_47547,N_47408,N_47101);
nor U47548 (N_47548,N_47063,N_47144);
or U47549 (N_47549,N_47397,N_47282);
nand U47550 (N_47550,N_47398,N_47311);
nor U47551 (N_47551,N_47149,N_47142);
nand U47552 (N_47552,N_47261,N_47450);
nor U47553 (N_47553,N_47084,N_47494);
nor U47554 (N_47554,N_47021,N_47387);
or U47555 (N_47555,N_47176,N_47091);
xor U47556 (N_47556,N_47103,N_47396);
and U47557 (N_47557,N_47280,N_47197);
or U47558 (N_47558,N_47191,N_47316);
xnor U47559 (N_47559,N_47071,N_47115);
or U47560 (N_47560,N_47260,N_47401);
nor U47561 (N_47561,N_47284,N_47182);
or U47562 (N_47562,N_47304,N_47482);
xor U47563 (N_47563,N_47472,N_47189);
or U47564 (N_47564,N_47286,N_47443);
and U47565 (N_47565,N_47407,N_47492);
nand U47566 (N_47566,N_47462,N_47287);
xor U47567 (N_47567,N_47228,N_47335);
or U47568 (N_47568,N_47100,N_47479);
and U47569 (N_47569,N_47095,N_47463);
and U47570 (N_47570,N_47330,N_47057);
nand U47571 (N_47571,N_47375,N_47388);
and U47572 (N_47572,N_47064,N_47302);
or U47573 (N_47573,N_47317,N_47234);
nand U47574 (N_47574,N_47451,N_47349);
xnor U47575 (N_47575,N_47239,N_47480);
nor U47576 (N_47576,N_47210,N_47029);
nand U47577 (N_47577,N_47121,N_47193);
nor U47578 (N_47578,N_47127,N_47037);
nor U47579 (N_47579,N_47452,N_47418);
and U47580 (N_47580,N_47423,N_47240);
and U47581 (N_47581,N_47226,N_47112);
xor U47582 (N_47582,N_47212,N_47141);
xor U47583 (N_47583,N_47377,N_47285);
and U47584 (N_47584,N_47439,N_47001);
or U47585 (N_47585,N_47295,N_47031);
nand U47586 (N_47586,N_47056,N_47324);
xor U47587 (N_47587,N_47448,N_47363);
xor U47588 (N_47588,N_47386,N_47460);
nor U47589 (N_47589,N_47162,N_47008);
xnor U47590 (N_47590,N_47314,N_47273);
nand U47591 (N_47591,N_47367,N_47139);
nor U47592 (N_47592,N_47107,N_47174);
xnor U47593 (N_47593,N_47026,N_47016);
xor U47594 (N_47594,N_47476,N_47169);
nor U47595 (N_47595,N_47133,N_47048);
xor U47596 (N_47596,N_47441,N_47481);
nand U47597 (N_47597,N_47173,N_47497);
or U47598 (N_47598,N_47389,N_47385);
or U47599 (N_47599,N_47250,N_47487);
or U47600 (N_47600,N_47461,N_47204);
and U47601 (N_47601,N_47061,N_47341);
or U47602 (N_47602,N_47252,N_47111);
and U47603 (N_47603,N_47490,N_47041);
nand U47604 (N_47604,N_47244,N_47458);
nor U47605 (N_47605,N_47166,N_47419);
or U47606 (N_47606,N_47213,N_47203);
nor U47607 (N_47607,N_47072,N_47268);
nor U47608 (N_47608,N_47296,N_47200);
xnor U47609 (N_47609,N_47120,N_47229);
or U47610 (N_47610,N_47098,N_47165);
nand U47611 (N_47611,N_47322,N_47357);
nor U47612 (N_47612,N_47087,N_47477);
xnor U47613 (N_47613,N_47054,N_47195);
and U47614 (N_47614,N_47449,N_47019);
and U47615 (N_47615,N_47465,N_47361);
nor U47616 (N_47616,N_47366,N_47171);
and U47617 (N_47617,N_47184,N_47453);
nand U47618 (N_47618,N_47154,N_47172);
xnor U47619 (N_47619,N_47395,N_47299);
xor U47620 (N_47620,N_47205,N_47058);
or U47621 (N_47621,N_47312,N_47368);
and U47622 (N_47622,N_47088,N_47342);
xnor U47623 (N_47623,N_47478,N_47483);
xor U47624 (N_47624,N_47475,N_47233);
and U47625 (N_47625,N_47114,N_47372);
nand U47626 (N_47626,N_47337,N_47215);
or U47627 (N_47627,N_47466,N_47288);
nand U47628 (N_47628,N_47308,N_47394);
xor U47629 (N_47629,N_47352,N_47126);
xnor U47630 (N_47630,N_47278,N_47093);
nand U47631 (N_47631,N_47256,N_47409);
nand U47632 (N_47632,N_47254,N_47362);
and U47633 (N_47633,N_47426,N_47208);
nor U47634 (N_47634,N_47345,N_47264);
and U47635 (N_47635,N_47491,N_47410);
xnor U47636 (N_47636,N_47415,N_47040);
nand U47637 (N_47637,N_47104,N_47247);
or U47638 (N_47638,N_47150,N_47433);
or U47639 (N_47639,N_47012,N_47313);
xor U47640 (N_47640,N_47148,N_47456);
or U47641 (N_47641,N_47329,N_47153);
xor U47642 (N_47642,N_47138,N_47262);
and U47643 (N_47643,N_47034,N_47004);
nor U47644 (N_47644,N_47297,N_47230);
nand U47645 (N_47645,N_47259,N_47348);
nor U47646 (N_47646,N_47444,N_47156);
or U47647 (N_47647,N_47334,N_47421);
or U47648 (N_47648,N_47014,N_47080);
nand U47649 (N_47649,N_47430,N_47003);
and U47650 (N_47650,N_47092,N_47336);
nor U47651 (N_47651,N_47151,N_47217);
or U47652 (N_47652,N_47249,N_47353);
xor U47653 (N_47653,N_47232,N_47108);
nand U47654 (N_47654,N_47202,N_47457);
and U47655 (N_47655,N_47258,N_47496);
nand U47656 (N_47656,N_47045,N_47028);
and U47657 (N_47657,N_47420,N_47218);
nor U47658 (N_47658,N_47227,N_47076);
and U47659 (N_47659,N_47134,N_47188);
or U47660 (N_47660,N_47049,N_47220);
or U47661 (N_47661,N_47413,N_47253);
xor U47662 (N_47662,N_47073,N_47245);
xor U47663 (N_47663,N_47123,N_47493);
nor U47664 (N_47664,N_47180,N_47293);
nand U47665 (N_47665,N_47155,N_47055);
xnor U47666 (N_47666,N_47131,N_47050);
nand U47667 (N_47667,N_47416,N_47081);
xnor U47668 (N_47668,N_47209,N_47332);
and U47669 (N_47669,N_47145,N_47163);
xnor U47670 (N_47670,N_47164,N_47292);
nand U47671 (N_47671,N_47235,N_47358);
or U47672 (N_47672,N_47158,N_47167);
or U47673 (N_47673,N_47143,N_47192);
nor U47674 (N_47674,N_47392,N_47216);
xor U47675 (N_47675,N_47168,N_47289);
xor U47676 (N_47676,N_47434,N_47340);
or U47677 (N_47677,N_47124,N_47351);
nand U47678 (N_47678,N_47010,N_47428);
xor U47679 (N_47679,N_47025,N_47321);
nor U47680 (N_47680,N_47024,N_47319);
and U47681 (N_47681,N_47412,N_47102);
nand U47682 (N_47682,N_47343,N_47291);
or U47683 (N_47683,N_47380,N_47116);
nor U47684 (N_47684,N_47083,N_47455);
nor U47685 (N_47685,N_47309,N_47185);
nand U47686 (N_47686,N_47179,N_47052);
or U47687 (N_47687,N_47011,N_47417);
xnor U47688 (N_47688,N_47294,N_47403);
xor U47689 (N_47689,N_47051,N_47178);
nor U47690 (N_47690,N_47241,N_47085);
or U47691 (N_47691,N_47059,N_47404);
nor U47692 (N_47692,N_47070,N_47425);
nand U47693 (N_47693,N_47136,N_47381);
nor U47694 (N_47694,N_47160,N_47399);
nand U47695 (N_47695,N_47400,N_47035);
xor U47696 (N_47696,N_47307,N_47468);
nor U47697 (N_47697,N_47238,N_47442);
xor U47698 (N_47698,N_47422,N_47032);
and U47699 (N_47699,N_47344,N_47199);
nand U47700 (N_47700,N_47006,N_47270);
nor U47701 (N_47701,N_47090,N_47459);
nor U47702 (N_47702,N_47113,N_47219);
nand U47703 (N_47703,N_47094,N_47437);
xor U47704 (N_47704,N_47435,N_47017);
nand U47705 (N_47705,N_47406,N_47339);
nor U47706 (N_47706,N_47251,N_47075);
and U47707 (N_47707,N_47194,N_47036);
xor U47708 (N_47708,N_47009,N_47269);
or U47709 (N_47709,N_47175,N_47474);
nand U47710 (N_47710,N_47207,N_47214);
or U47711 (N_47711,N_47489,N_47371);
or U47712 (N_47712,N_47007,N_47427);
nand U47713 (N_47713,N_47376,N_47326);
or U47714 (N_47714,N_47486,N_47275);
or U47715 (N_47715,N_47152,N_47354);
nand U47716 (N_47716,N_47384,N_47033);
xnor U47717 (N_47717,N_47393,N_47022);
xor U47718 (N_47718,N_47391,N_47196);
and U47719 (N_47719,N_47067,N_47360);
or U47720 (N_47720,N_47281,N_47440);
or U47721 (N_47721,N_47431,N_47078);
and U47722 (N_47722,N_47106,N_47488);
and U47723 (N_47723,N_47221,N_47429);
nor U47724 (N_47724,N_47186,N_47109);
or U47725 (N_47725,N_47097,N_47414);
xor U47726 (N_47726,N_47495,N_47276);
or U47727 (N_47727,N_47469,N_47181);
nor U47728 (N_47728,N_47485,N_47350);
nor U47729 (N_47729,N_47347,N_47082);
nand U47730 (N_47730,N_47096,N_47266);
xor U47731 (N_47731,N_47117,N_47027);
or U47732 (N_47732,N_47248,N_47467);
nor U47733 (N_47733,N_47236,N_47265);
xor U47734 (N_47734,N_47089,N_47147);
nand U47735 (N_47735,N_47157,N_47225);
nor U47736 (N_47736,N_47038,N_47062);
nor U47737 (N_47737,N_47132,N_47243);
nand U47738 (N_47738,N_47454,N_47223);
nand U47739 (N_47739,N_47211,N_47046);
and U47740 (N_47740,N_47424,N_47018);
and U47741 (N_47741,N_47077,N_47255);
nand U47742 (N_47742,N_47279,N_47140);
nand U47743 (N_47743,N_47338,N_47079);
and U47744 (N_47744,N_47272,N_47383);
or U47745 (N_47745,N_47125,N_47043);
nor U47746 (N_47746,N_47201,N_47271);
and U47747 (N_47747,N_47074,N_47301);
nand U47748 (N_47748,N_47119,N_47373);
nor U47749 (N_47749,N_47325,N_47346);
or U47750 (N_47750,N_47211,N_47150);
or U47751 (N_47751,N_47142,N_47279);
xor U47752 (N_47752,N_47205,N_47143);
or U47753 (N_47753,N_47400,N_47044);
nand U47754 (N_47754,N_47189,N_47201);
xor U47755 (N_47755,N_47496,N_47379);
nand U47756 (N_47756,N_47068,N_47496);
nand U47757 (N_47757,N_47412,N_47291);
nand U47758 (N_47758,N_47309,N_47362);
nor U47759 (N_47759,N_47207,N_47176);
and U47760 (N_47760,N_47377,N_47038);
and U47761 (N_47761,N_47270,N_47180);
nand U47762 (N_47762,N_47339,N_47150);
and U47763 (N_47763,N_47066,N_47373);
xnor U47764 (N_47764,N_47468,N_47052);
or U47765 (N_47765,N_47118,N_47106);
nand U47766 (N_47766,N_47258,N_47383);
xnor U47767 (N_47767,N_47131,N_47422);
and U47768 (N_47768,N_47228,N_47206);
nor U47769 (N_47769,N_47237,N_47294);
or U47770 (N_47770,N_47041,N_47301);
or U47771 (N_47771,N_47129,N_47289);
or U47772 (N_47772,N_47018,N_47208);
and U47773 (N_47773,N_47161,N_47061);
or U47774 (N_47774,N_47016,N_47099);
nand U47775 (N_47775,N_47461,N_47467);
nand U47776 (N_47776,N_47092,N_47210);
or U47777 (N_47777,N_47306,N_47005);
xor U47778 (N_47778,N_47091,N_47476);
or U47779 (N_47779,N_47326,N_47422);
nand U47780 (N_47780,N_47011,N_47339);
and U47781 (N_47781,N_47470,N_47208);
and U47782 (N_47782,N_47030,N_47458);
and U47783 (N_47783,N_47218,N_47349);
xnor U47784 (N_47784,N_47498,N_47460);
xnor U47785 (N_47785,N_47049,N_47127);
or U47786 (N_47786,N_47217,N_47365);
and U47787 (N_47787,N_47446,N_47300);
nand U47788 (N_47788,N_47480,N_47178);
nor U47789 (N_47789,N_47050,N_47109);
xnor U47790 (N_47790,N_47015,N_47460);
or U47791 (N_47791,N_47193,N_47341);
xor U47792 (N_47792,N_47455,N_47322);
or U47793 (N_47793,N_47303,N_47407);
xor U47794 (N_47794,N_47030,N_47439);
xnor U47795 (N_47795,N_47005,N_47462);
and U47796 (N_47796,N_47494,N_47469);
nor U47797 (N_47797,N_47135,N_47479);
or U47798 (N_47798,N_47385,N_47051);
xnor U47799 (N_47799,N_47371,N_47051);
or U47800 (N_47800,N_47415,N_47190);
or U47801 (N_47801,N_47119,N_47380);
or U47802 (N_47802,N_47441,N_47127);
or U47803 (N_47803,N_47080,N_47197);
nor U47804 (N_47804,N_47415,N_47031);
nand U47805 (N_47805,N_47235,N_47041);
nor U47806 (N_47806,N_47483,N_47146);
or U47807 (N_47807,N_47190,N_47187);
or U47808 (N_47808,N_47201,N_47397);
and U47809 (N_47809,N_47436,N_47171);
nor U47810 (N_47810,N_47289,N_47093);
nand U47811 (N_47811,N_47440,N_47487);
or U47812 (N_47812,N_47255,N_47327);
or U47813 (N_47813,N_47478,N_47095);
nor U47814 (N_47814,N_47456,N_47407);
nand U47815 (N_47815,N_47332,N_47045);
xnor U47816 (N_47816,N_47145,N_47177);
or U47817 (N_47817,N_47387,N_47129);
or U47818 (N_47818,N_47293,N_47468);
or U47819 (N_47819,N_47168,N_47472);
nor U47820 (N_47820,N_47295,N_47377);
nor U47821 (N_47821,N_47271,N_47112);
xor U47822 (N_47822,N_47099,N_47111);
nor U47823 (N_47823,N_47251,N_47214);
nand U47824 (N_47824,N_47237,N_47039);
xor U47825 (N_47825,N_47054,N_47219);
xnor U47826 (N_47826,N_47187,N_47122);
or U47827 (N_47827,N_47397,N_47342);
xor U47828 (N_47828,N_47124,N_47209);
nor U47829 (N_47829,N_47261,N_47224);
xnor U47830 (N_47830,N_47320,N_47264);
and U47831 (N_47831,N_47256,N_47488);
nor U47832 (N_47832,N_47077,N_47094);
nand U47833 (N_47833,N_47360,N_47238);
nor U47834 (N_47834,N_47490,N_47015);
xnor U47835 (N_47835,N_47358,N_47471);
xor U47836 (N_47836,N_47247,N_47386);
nand U47837 (N_47837,N_47093,N_47294);
nand U47838 (N_47838,N_47002,N_47472);
or U47839 (N_47839,N_47362,N_47218);
or U47840 (N_47840,N_47251,N_47023);
nor U47841 (N_47841,N_47387,N_47281);
nor U47842 (N_47842,N_47178,N_47290);
nor U47843 (N_47843,N_47421,N_47085);
nor U47844 (N_47844,N_47422,N_47407);
nand U47845 (N_47845,N_47428,N_47004);
and U47846 (N_47846,N_47301,N_47314);
xnor U47847 (N_47847,N_47377,N_47177);
nand U47848 (N_47848,N_47362,N_47044);
nor U47849 (N_47849,N_47440,N_47184);
nor U47850 (N_47850,N_47018,N_47458);
or U47851 (N_47851,N_47439,N_47422);
and U47852 (N_47852,N_47303,N_47135);
nor U47853 (N_47853,N_47299,N_47268);
nand U47854 (N_47854,N_47237,N_47047);
and U47855 (N_47855,N_47115,N_47056);
nand U47856 (N_47856,N_47093,N_47264);
or U47857 (N_47857,N_47057,N_47220);
or U47858 (N_47858,N_47169,N_47314);
and U47859 (N_47859,N_47174,N_47246);
xnor U47860 (N_47860,N_47445,N_47129);
nand U47861 (N_47861,N_47206,N_47401);
and U47862 (N_47862,N_47112,N_47157);
xor U47863 (N_47863,N_47387,N_47006);
nor U47864 (N_47864,N_47423,N_47188);
and U47865 (N_47865,N_47326,N_47196);
nand U47866 (N_47866,N_47033,N_47427);
nand U47867 (N_47867,N_47193,N_47498);
or U47868 (N_47868,N_47395,N_47453);
and U47869 (N_47869,N_47364,N_47308);
or U47870 (N_47870,N_47400,N_47401);
or U47871 (N_47871,N_47236,N_47154);
nand U47872 (N_47872,N_47355,N_47098);
or U47873 (N_47873,N_47259,N_47012);
nor U47874 (N_47874,N_47079,N_47113);
xnor U47875 (N_47875,N_47112,N_47159);
xnor U47876 (N_47876,N_47298,N_47215);
nor U47877 (N_47877,N_47094,N_47059);
nand U47878 (N_47878,N_47169,N_47430);
or U47879 (N_47879,N_47446,N_47088);
nor U47880 (N_47880,N_47096,N_47367);
nor U47881 (N_47881,N_47335,N_47176);
or U47882 (N_47882,N_47352,N_47260);
nand U47883 (N_47883,N_47254,N_47279);
nor U47884 (N_47884,N_47352,N_47033);
nor U47885 (N_47885,N_47045,N_47316);
nor U47886 (N_47886,N_47120,N_47169);
and U47887 (N_47887,N_47408,N_47130);
nor U47888 (N_47888,N_47432,N_47084);
or U47889 (N_47889,N_47314,N_47098);
nand U47890 (N_47890,N_47430,N_47213);
or U47891 (N_47891,N_47408,N_47241);
nand U47892 (N_47892,N_47047,N_47131);
or U47893 (N_47893,N_47064,N_47443);
and U47894 (N_47894,N_47329,N_47471);
xor U47895 (N_47895,N_47401,N_47417);
and U47896 (N_47896,N_47290,N_47055);
xnor U47897 (N_47897,N_47260,N_47402);
and U47898 (N_47898,N_47427,N_47111);
or U47899 (N_47899,N_47176,N_47334);
nor U47900 (N_47900,N_47395,N_47414);
or U47901 (N_47901,N_47372,N_47485);
xnor U47902 (N_47902,N_47394,N_47241);
and U47903 (N_47903,N_47211,N_47132);
nand U47904 (N_47904,N_47373,N_47372);
xnor U47905 (N_47905,N_47325,N_47240);
nor U47906 (N_47906,N_47292,N_47122);
or U47907 (N_47907,N_47254,N_47061);
xor U47908 (N_47908,N_47400,N_47469);
nand U47909 (N_47909,N_47241,N_47076);
or U47910 (N_47910,N_47402,N_47286);
nor U47911 (N_47911,N_47457,N_47237);
and U47912 (N_47912,N_47148,N_47378);
xnor U47913 (N_47913,N_47058,N_47358);
and U47914 (N_47914,N_47300,N_47424);
and U47915 (N_47915,N_47451,N_47467);
and U47916 (N_47916,N_47441,N_47197);
nand U47917 (N_47917,N_47061,N_47373);
nor U47918 (N_47918,N_47230,N_47006);
nor U47919 (N_47919,N_47490,N_47130);
or U47920 (N_47920,N_47233,N_47044);
nor U47921 (N_47921,N_47018,N_47107);
and U47922 (N_47922,N_47454,N_47051);
nand U47923 (N_47923,N_47367,N_47497);
nand U47924 (N_47924,N_47428,N_47048);
nand U47925 (N_47925,N_47244,N_47375);
xor U47926 (N_47926,N_47369,N_47378);
and U47927 (N_47927,N_47473,N_47255);
xor U47928 (N_47928,N_47193,N_47218);
and U47929 (N_47929,N_47107,N_47094);
or U47930 (N_47930,N_47334,N_47062);
xor U47931 (N_47931,N_47426,N_47330);
xor U47932 (N_47932,N_47093,N_47013);
nor U47933 (N_47933,N_47217,N_47234);
nand U47934 (N_47934,N_47119,N_47424);
xor U47935 (N_47935,N_47043,N_47209);
nor U47936 (N_47936,N_47313,N_47288);
or U47937 (N_47937,N_47157,N_47366);
nand U47938 (N_47938,N_47025,N_47320);
xor U47939 (N_47939,N_47309,N_47023);
nand U47940 (N_47940,N_47269,N_47174);
nor U47941 (N_47941,N_47203,N_47258);
and U47942 (N_47942,N_47240,N_47064);
nor U47943 (N_47943,N_47319,N_47454);
nand U47944 (N_47944,N_47232,N_47294);
xnor U47945 (N_47945,N_47108,N_47444);
and U47946 (N_47946,N_47017,N_47380);
nand U47947 (N_47947,N_47216,N_47278);
xor U47948 (N_47948,N_47115,N_47496);
nor U47949 (N_47949,N_47298,N_47237);
and U47950 (N_47950,N_47332,N_47237);
xnor U47951 (N_47951,N_47463,N_47258);
or U47952 (N_47952,N_47470,N_47199);
xor U47953 (N_47953,N_47195,N_47003);
nor U47954 (N_47954,N_47335,N_47183);
nand U47955 (N_47955,N_47283,N_47131);
and U47956 (N_47956,N_47058,N_47407);
nor U47957 (N_47957,N_47231,N_47136);
nand U47958 (N_47958,N_47078,N_47250);
nand U47959 (N_47959,N_47032,N_47298);
xor U47960 (N_47960,N_47390,N_47048);
nand U47961 (N_47961,N_47011,N_47196);
or U47962 (N_47962,N_47027,N_47203);
and U47963 (N_47963,N_47068,N_47258);
or U47964 (N_47964,N_47080,N_47381);
nand U47965 (N_47965,N_47421,N_47058);
nand U47966 (N_47966,N_47185,N_47099);
and U47967 (N_47967,N_47112,N_47248);
and U47968 (N_47968,N_47239,N_47424);
nor U47969 (N_47969,N_47265,N_47181);
or U47970 (N_47970,N_47058,N_47203);
nor U47971 (N_47971,N_47081,N_47493);
and U47972 (N_47972,N_47081,N_47097);
or U47973 (N_47973,N_47302,N_47261);
or U47974 (N_47974,N_47411,N_47195);
and U47975 (N_47975,N_47001,N_47121);
and U47976 (N_47976,N_47052,N_47074);
xor U47977 (N_47977,N_47371,N_47477);
nor U47978 (N_47978,N_47096,N_47090);
nor U47979 (N_47979,N_47430,N_47487);
nand U47980 (N_47980,N_47245,N_47136);
or U47981 (N_47981,N_47139,N_47015);
or U47982 (N_47982,N_47259,N_47013);
nor U47983 (N_47983,N_47147,N_47251);
or U47984 (N_47984,N_47329,N_47288);
xor U47985 (N_47985,N_47157,N_47229);
and U47986 (N_47986,N_47405,N_47448);
nand U47987 (N_47987,N_47122,N_47334);
or U47988 (N_47988,N_47190,N_47116);
nand U47989 (N_47989,N_47283,N_47352);
or U47990 (N_47990,N_47434,N_47218);
nor U47991 (N_47991,N_47258,N_47337);
xnor U47992 (N_47992,N_47157,N_47256);
and U47993 (N_47993,N_47358,N_47167);
and U47994 (N_47994,N_47122,N_47188);
or U47995 (N_47995,N_47312,N_47225);
nand U47996 (N_47996,N_47029,N_47012);
or U47997 (N_47997,N_47097,N_47497);
or U47998 (N_47998,N_47418,N_47092);
or U47999 (N_47999,N_47256,N_47459);
and U48000 (N_48000,N_47802,N_47993);
and U48001 (N_48001,N_47641,N_47596);
nand U48002 (N_48002,N_47709,N_47728);
or U48003 (N_48003,N_47638,N_47605);
or U48004 (N_48004,N_47590,N_47897);
nor U48005 (N_48005,N_47547,N_47512);
xor U48006 (N_48006,N_47853,N_47881);
xnor U48007 (N_48007,N_47631,N_47732);
and U48008 (N_48008,N_47941,N_47684);
and U48009 (N_48009,N_47515,N_47565);
nor U48010 (N_48010,N_47519,N_47649);
or U48011 (N_48011,N_47910,N_47822);
and U48012 (N_48012,N_47757,N_47575);
and U48013 (N_48013,N_47989,N_47574);
and U48014 (N_48014,N_47609,N_47997);
xnor U48015 (N_48015,N_47685,N_47983);
xor U48016 (N_48016,N_47758,N_47751);
and U48017 (N_48017,N_47607,N_47604);
nand U48018 (N_48018,N_47667,N_47722);
nor U48019 (N_48019,N_47961,N_47659);
nand U48020 (N_48020,N_47894,N_47554);
xor U48021 (N_48021,N_47738,N_47524);
xnor U48022 (N_48022,N_47545,N_47896);
nor U48023 (N_48023,N_47697,N_47787);
xnor U48024 (N_48024,N_47959,N_47804);
xnor U48025 (N_48025,N_47527,N_47563);
nor U48026 (N_48026,N_47944,N_47522);
xor U48027 (N_48027,N_47692,N_47736);
nand U48028 (N_48028,N_47695,N_47798);
nor U48029 (N_48029,N_47980,N_47916);
or U48030 (N_48030,N_47591,N_47613);
nand U48031 (N_48031,N_47791,N_47955);
xnor U48032 (N_48032,N_47960,N_47805);
nand U48033 (N_48033,N_47840,N_47534);
xnor U48034 (N_48034,N_47964,N_47931);
xor U48035 (N_48035,N_47560,N_47755);
nand U48036 (N_48036,N_47674,N_47851);
xor U48037 (N_48037,N_47807,N_47525);
xor U48038 (N_48038,N_47516,N_47647);
and U48039 (N_48039,N_47686,N_47643);
nand U48040 (N_48040,N_47784,N_47918);
nor U48041 (N_48041,N_47905,N_47612);
nor U48042 (N_48042,N_47810,N_47837);
nor U48043 (N_48043,N_47922,N_47733);
nor U48044 (N_48044,N_47812,N_47937);
and U48045 (N_48045,N_47713,N_47539);
or U48046 (N_48046,N_47572,N_47657);
or U48047 (N_48047,N_47870,N_47999);
nand U48048 (N_48048,N_47611,N_47526);
or U48049 (N_48049,N_47530,N_47963);
nand U48050 (N_48050,N_47538,N_47835);
nand U48051 (N_48051,N_47585,N_47621);
xor U48052 (N_48052,N_47882,N_47834);
nor U48053 (N_48053,N_47592,N_47786);
and U48054 (N_48054,N_47749,N_47599);
nor U48055 (N_48055,N_47844,N_47873);
nand U48056 (N_48056,N_47676,N_47823);
nand U48057 (N_48057,N_47848,N_47769);
xnor U48058 (N_48058,N_47696,N_47943);
nand U48059 (N_48059,N_47533,N_47670);
xor U48060 (N_48060,N_47759,N_47829);
xnor U48061 (N_48061,N_47994,N_47741);
and U48062 (N_48062,N_47637,N_47932);
xnor U48063 (N_48063,N_47566,N_47588);
and U48064 (N_48064,N_47866,N_47675);
nand U48065 (N_48065,N_47818,N_47940);
and U48066 (N_48066,N_47614,N_47995);
and U48067 (N_48067,N_47507,N_47793);
nand U48068 (N_48068,N_47734,N_47962);
nor U48069 (N_48069,N_47903,N_47912);
or U48070 (N_48070,N_47648,N_47627);
xor U48071 (N_48071,N_47765,N_47562);
and U48072 (N_48072,N_47602,N_47981);
and U48073 (N_48073,N_47813,N_47699);
or U48074 (N_48074,N_47909,N_47714);
nor U48075 (N_48075,N_47788,N_47982);
nand U48076 (N_48076,N_47680,N_47620);
xor U48077 (N_48077,N_47785,N_47571);
nand U48078 (N_48078,N_47839,N_47671);
or U48079 (N_48079,N_47619,N_47958);
or U48080 (N_48080,N_47718,N_47708);
xnor U48081 (N_48081,N_47750,N_47966);
and U48082 (N_48082,N_47930,N_47712);
and U48083 (N_48083,N_47781,N_47908);
nor U48084 (N_48084,N_47814,N_47716);
nand U48085 (N_48085,N_47629,N_47664);
or U48086 (N_48086,N_47715,N_47639);
xor U48087 (N_48087,N_47886,N_47723);
and U48088 (N_48088,N_47795,N_47730);
and U48089 (N_48089,N_47957,N_47672);
nor U48090 (N_48090,N_47929,N_47770);
and U48091 (N_48091,N_47772,N_47863);
or U48092 (N_48092,N_47953,N_47622);
xnor U48093 (N_48093,N_47949,N_47846);
and U48094 (N_48094,N_47794,N_47871);
xor U48095 (N_48095,N_47917,N_47744);
nor U48096 (N_48096,N_47827,N_47831);
nand U48097 (N_48097,N_47862,N_47731);
xnor U48098 (N_48098,N_47603,N_47767);
or U48099 (N_48099,N_47901,N_47816);
and U48100 (N_48100,N_47669,N_47776);
and U48101 (N_48101,N_47880,N_47589);
nor U48102 (N_48102,N_47860,N_47690);
or U48103 (N_48103,N_47577,N_47617);
or U48104 (N_48104,N_47595,N_47973);
nor U48105 (N_48105,N_47655,N_47872);
nand U48106 (N_48106,N_47573,N_47766);
or U48107 (N_48107,N_47830,N_47606);
nor U48108 (N_48108,N_47698,N_47868);
xor U48109 (N_48109,N_47624,N_47864);
or U48110 (N_48110,N_47729,N_47551);
nor U48111 (N_48111,N_47884,N_47660);
and U48112 (N_48112,N_47998,N_47911);
xnor U48113 (N_48113,N_47557,N_47892);
and U48114 (N_48114,N_47878,N_47546);
nor U48115 (N_48115,N_47775,N_47646);
nor U48116 (N_48116,N_47842,N_47531);
xnor U48117 (N_48117,N_47645,N_47509);
and U48118 (N_48118,N_47771,N_47514);
nor U48119 (N_48119,N_47779,N_47703);
nand U48120 (N_48120,N_47825,N_47867);
xor U48121 (N_48121,N_47799,N_47707);
nand U48122 (N_48122,N_47623,N_47762);
or U48123 (N_48123,N_47986,N_47540);
or U48124 (N_48124,N_47920,N_47935);
nand U48125 (N_48125,N_47673,N_47833);
or U48126 (N_48126,N_47978,N_47518);
or U48127 (N_48127,N_47682,N_47735);
nand U48128 (N_48128,N_47567,N_47847);
nand U48129 (N_48129,N_47542,N_47858);
and U48130 (N_48130,N_47907,N_47536);
xor U48131 (N_48131,N_47663,N_47938);
or U48132 (N_48132,N_47511,N_47528);
nor U48133 (N_48133,N_47678,N_47817);
nand U48134 (N_48134,N_47824,N_47549);
nand U48135 (N_48135,N_47583,N_47826);
nand U48136 (N_48136,N_47876,N_47936);
nand U48137 (N_48137,N_47773,N_47927);
and U48138 (N_48138,N_47666,N_47656);
xnor U48139 (N_48139,N_47745,N_47569);
nor U48140 (N_48140,N_47946,N_47815);
nand U48141 (N_48141,N_47724,N_47581);
xor U48142 (N_48142,N_47568,N_47926);
xnor U48143 (N_48143,N_47504,N_47702);
xor U48144 (N_48144,N_47752,N_47598);
and U48145 (N_48145,N_47662,N_47644);
xor U48146 (N_48146,N_47869,N_47942);
nor U48147 (N_48147,N_47889,N_47501);
xnor U48148 (N_48148,N_47874,N_47933);
or U48149 (N_48149,N_47857,N_47742);
nand U48150 (N_48150,N_47548,N_47832);
nand U48151 (N_48151,N_47683,N_47888);
nand U48152 (N_48152,N_47701,N_47968);
or U48153 (N_48153,N_47821,N_47819);
nand U48154 (N_48154,N_47653,N_47502);
nor U48155 (N_48155,N_47820,N_47977);
xnor U48156 (N_48156,N_47754,N_47739);
nor U48157 (N_48157,N_47996,N_47768);
or U48158 (N_48158,N_47985,N_47520);
or U48159 (N_48159,N_47774,N_47600);
nand U48160 (N_48160,N_47780,N_47950);
or U48161 (N_48161,N_47618,N_47928);
or U48162 (N_48162,N_47838,N_47796);
and U48163 (N_48163,N_47992,N_47727);
and U48164 (N_48164,N_47934,N_47523);
xor U48165 (N_48165,N_47753,N_47921);
and U48166 (N_48166,N_47783,N_47665);
nor U48167 (N_48167,N_47505,N_47809);
xor U48168 (N_48168,N_47642,N_47763);
and U48169 (N_48169,N_47705,N_47891);
or U48170 (N_48170,N_47521,N_47679);
nor U48171 (N_48171,N_47850,N_47969);
nor U48172 (N_48172,N_47841,N_47803);
nand U48173 (N_48173,N_47597,N_47694);
nand U48174 (N_48174,N_47510,N_47865);
nand U48175 (N_48175,N_47601,N_47808);
and U48176 (N_48176,N_47984,N_47756);
and U48177 (N_48177,N_47651,N_47704);
nor U48178 (N_48178,N_47828,N_47726);
or U48179 (N_48179,N_47777,N_47800);
nor U48180 (N_48180,N_47974,N_47914);
nor U48181 (N_48181,N_47859,N_47576);
and U48182 (N_48182,N_47628,N_47843);
or U48183 (N_48183,N_47652,N_47550);
nor U48184 (N_48184,N_47845,N_47654);
nor U48185 (N_48185,N_47792,N_47508);
nand U48186 (N_48186,N_47893,N_47529);
and U48187 (N_48187,N_47668,N_47748);
nand U48188 (N_48188,N_47677,N_47939);
or U48189 (N_48189,N_47902,N_47717);
nor U48190 (N_48190,N_47877,N_47711);
xnor U48191 (N_48191,N_47500,N_47970);
nand U48192 (N_48192,N_47991,N_47887);
nor U48193 (N_48193,N_47951,N_47720);
or U48194 (N_48194,N_47615,N_47811);
or U48195 (N_48195,N_47885,N_47954);
nor U48196 (N_48196,N_47979,N_47658);
nand U48197 (N_48197,N_47552,N_47761);
nand U48198 (N_48198,N_47544,N_47913);
and U48199 (N_48199,N_47971,N_47789);
nand U48200 (N_48200,N_47710,N_47691);
and U48201 (N_48201,N_47608,N_47640);
nor U48202 (N_48202,N_47535,N_47513);
nor U48203 (N_48203,N_47760,N_47661);
xor U48204 (N_48204,N_47740,N_47559);
or U48205 (N_48205,N_47879,N_47923);
and U48206 (N_48206,N_47625,N_47584);
or U48207 (N_48207,N_47797,N_47537);
nor U48208 (N_48208,N_47790,N_47975);
nand U48209 (N_48209,N_47650,N_47616);
or U48210 (N_48210,N_47782,N_47737);
and U48211 (N_48211,N_47987,N_47919);
and U48212 (N_48212,N_47956,N_47555);
xor U48213 (N_48213,N_47561,N_47579);
nor U48214 (N_48214,N_47915,N_47972);
or U48215 (N_48215,N_47681,N_47634);
or U48216 (N_48216,N_47564,N_47635);
or U48217 (N_48217,N_47965,N_47594);
xnor U48218 (N_48218,N_47746,N_47700);
nor U48219 (N_48219,N_47688,N_47900);
and U48220 (N_48220,N_47693,N_47778);
nor U48221 (N_48221,N_47556,N_47553);
and U48222 (N_48222,N_47854,N_47747);
and U48223 (N_48223,N_47948,N_47630);
nand U48224 (N_48224,N_47806,N_47626);
nand U48225 (N_48225,N_47587,N_47578);
or U48226 (N_48226,N_47875,N_47904);
or U48227 (N_48227,N_47633,N_47976);
and U48228 (N_48228,N_47924,N_47593);
xor U48229 (N_48229,N_47586,N_47861);
nand U48230 (N_48230,N_47558,N_47988);
and U48231 (N_48231,N_47952,N_47895);
and U48232 (N_48232,N_47849,N_47725);
and U48233 (N_48233,N_47855,N_47764);
or U48234 (N_48234,N_47610,N_47990);
and U48235 (N_48235,N_47721,N_47689);
nor U48236 (N_48236,N_47856,N_47947);
xor U48237 (N_48237,N_47580,N_47883);
xnor U48238 (N_48238,N_47899,N_47582);
and U48239 (N_48239,N_47890,N_47967);
and U48240 (N_48240,N_47632,N_47570);
xor U48241 (N_48241,N_47532,N_47906);
xor U48242 (N_48242,N_47687,N_47719);
xnor U48243 (N_48243,N_47945,N_47517);
nand U48244 (N_48244,N_47636,N_47925);
or U48245 (N_48245,N_47706,N_47743);
nand U48246 (N_48246,N_47852,N_47898);
and U48247 (N_48247,N_47541,N_47801);
nor U48248 (N_48248,N_47506,N_47836);
xnor U48249 (N_48249,N_47543,N_47503);
nand U48250 (N_48250,N_47999,N_47584);
nand U48251 (N_48251,N_47869,N_47765);
and U48252 (N_48252,N_47609,N_47617);
nor U48253 (N_48253,N_47743,N_47507);
nor U48254 (N_48254,N_47938,N_47534);
xor U48255 (N_48255,N_47739,N_47929);
xor U48256 (N_48256,N_47527,N_47638);
or U48257 (N_48257,N_47709,N_47536);
nand U48258 (N_48258,N_47903,N_47886);
and U48259 (N_48259,N_47505,N_47640);
nand U48260 (N_48260,N_47856,N_47649);
and U48261 (N_48261,N_47872,N_47848);
and U48262 (N_48262,N_47811,N_47826);
or U48263 (N_48263,N_47655,N_47860);
xnor U48264 (N_48264,N_47972,N_47641);
xnor U48265 (N_48265,N_47802,N_47938);
nor U48266 (N_48266,N_47691,N_47787);
nand U48267 (N_48267,N_47955,N_47757);
nand U48268 (N_48268,N_47677,N_47948);
and U48269 (N_48269,N_47664,N_47999);
xor U48270 (N_48270,N_47938,N_47703);
and U48271 (N_48271,N_47871,N_47918);
nand U48272 (N_48272,N_47619,N_47501);
nand U48273 (N_48273,N_47921,N_47598);
nand U48274 (N_48274,N_47780,N_47532);
nand U48275 (N_48275,N_47798,N_47812);
and U48276 (N_48276,N_47873,N_47925);
nand U48277 (N_48277,N_47955,N_47646);
nand U48278 (N_48278,N_47964,N_47858);
xor U48279 (N_48279,N_47567,N_47621);
and U48280 (N_48280,N_47982,N_47881);
nor U48281 (N_48281,N_47580,N_47595);
nor U48282 (N_48282,N_47569,N_47652);
or U48283 (N_48283,N_47999,N_47990);
nand U48284 (N_48284,N_47643,N_47779);
nor U48285 (N_48285,N_47906,N_47979);
and U48286 (N_48286,N_47546,N_47789);
xnor U48287 (N_48287,N_47835,N_47516);
or U48288 (N_48288,N_47595,N_47570);
nor U48289 (N_48289,N_47638,N_47712);
xnor U48290 (N_48290,N_47854,N_47676);
nand U48291 (N_48291,N_47501,N_47748);
nor U48292 (N_48292,N_47753,N_47927);
nand U48293 (N_48293,N_47732,N_47623);
nand U48294 (N_48294,N_47671,N_47933);
or U48295 (N_48295,N_47723,N_47699);
nor U48296 (N_48296,N_47753,N_47811);
nand U48297 (N_48297,N_47924,N_47532);
xor U48298 (N_48298,N_47511,N_47540);
xor U48299 (N_48299,N_47596,N_47551);
and U48300 (N_48300,N_47836,N_47512);
and U48301 (N_48301,N_47798,N_47873);
or U48302 (N_48302,N_47982,N_47520);
xnor U48303 (N_48303,N_47912,N_47556);
xnor U48304 (N_48304,N_47624,N_47794);
nor U48305 (N_48305,N_47995,N_47792);
xor U48306 (N_48306,N_47734,N_47866);
xnor U48307 (N_48307,N_47925,N_47994);
and U48308 (N_48308,N_47810,N_47874);
or U48309 (N_48309,N_47609,N_47709);
or U48310 (N_48310,N_47583,N_47606);
nor U48311 (N_48311,N_47872,N_47719);
nand U48312 (N_48312,N_47809,N_47837);
nand U48313 (N_48313,N_47842,N_47855);
nor U48314 (N_48314,N_47700,N_47621);
xnor U48315 (N_48315,N_47603,N_47775);
and U48316 (N_48316,N_47535,N_47761);
xor U48317 (N_48317,N_47980,N_47722);
and U48318 (N_48318,N_47889,N_47511);
nor U48319 (N_48319,N_47661,N_47730);
or U48320 (N_48320,N_47898,N_47690);
or U48321 (N_48321,N_47860,N_47623);
nor U48322 (N_48322,N_47599,N_47798);
and U48323 (N_48323,N_47527,N_47700);
and U48324 (N_48324,N_47771,N_47776);
or U48325 (N_48325,N_47630,N_47781);
nand U48326 (N_48326,N_47504,N_47952);
and U48327 (N_48327,N_47509,N_47579);
and U48328 (N_48328,N_47577,N_47574);
xor U48329 (N_48329,N_47645,N_47721);
nor U48330 (N_48330,N_47502,N_47887);
xor U48331 (N_48331,N_47605,N_47578);
xor U48332 (N_48332,N_47666,N_47816);
and U48333 (N_48333,N_47715,N_47703);
or U48334 (N_48334,N_47601,N_47759);
nor U48335 (N_48335,N_47887,N_47654);
nand U48336 (N_48336,N_47922,N_47562);
nor U48337 (N_48337,N_47956,N_47724);
nor U48338 (N_48338,N_47563,N_47990);
nand U48339 (N_48339,N_47907,N_47822);
and U48340 (N_48340,N_47905,N_47809);
or U48341 (N_48341,N_47770,N_47846);
nand U48342 (N_48342,N_47971,N_47908);
nand U48343 (N_48343,N_47876,N_47896);
and U48344 (N_48344,N_47800,N_47926);
and U48345 (N_48345,N_47630,N_47535);
and U48346 (N_48346,N_47550,N_47547);
nor U48347 (N_48347,N_47844,N_47841);
and U48348 (N_48348,N_47634,N_47637);
or U48349 (N_48349,N_47833,N_47741);
xor U48350 (N_48350,N_47598,N_47711);
or U48351 (N_48351,N_47851,N_47653);
xnor U48352 (N_48352,N_47869,N_47633);
nor U48353 (N_48353,N_47788,N_47500);
xor U48354 (N_48354,N_47826,N_47809);
nor U48355 (N_48355,N_47583,N_47752);
or U48356 (N_48356,N_47808,N_47635);
nor U48357 (N_48357,N_47947,N_47878);
nand U48358 (N_48358,N_47772,N_47747);
nor U48359 (N_48359,N_47946,N_47990);
nand U48360 (N_48360,N_47719,N_47751);
and U48361 (N_48361,N_47938,N_47818);
nor U48362 (N_48362,N_47963,N_47653);
nor U48363 (N_48363,N_47509,N_47675);
and U48364 (N_48364,N_47871,N_47789);
or U48365 (N_48365,N_47610,N_47570);
and U48366 (N_48366,N_47629,N_47574);
and U48367 (N_48367,N_47672,N_47517);
nand U48368 (N_48368,N_47874,N_47739);
xor U48369 (N_48369,N_47740,N_47849);
nor U48370 (N_48370,N_47853,N_47790);
nor U48371 (N_48371,N_47960,N_47653);
xor U48372 (N_48372,N_47815,N_47715);
nor U48373 (N_48373,N_47584,N_47830);
nor U48374 (N_48374,N_47962,N_47953);
and U48375 (N_48375,N_47500,N_47882);
and U48376 (N_48376,N_47808,N_47590);
nor U48377 (N_48377,N_47849,N_47676);
or U48378 (N_48378,N_47951,N_47992);
or U48379 (N_48379,N_47770,N_47677);
or U48380 (N_48380,N_47912,N_47721);
xnor U48381 (N_48381,N_47742,N_47932);
nor U48382 (N_48382,N_47946,N_47594);
nor U48383 (N_48383,N_47734,N_47832);
nor U48384 (N_48384,N_47817,N_47584);
nor U48385 (N_48385,N_47704,N_47628);
xor U48386 (N_48386,N_47520,N_47885);
or U48387 (N_48387,N_47954,N_47859);
and U48388 (N_48388,N_47557,N_47656);
or U48389 (N_48389,N_47541,N_47670);
nand U48390 (N_48390,N_47864,N_47622);
nor U48391 (N_48391,N_47699,N_47508);
xnor U48392 (N_48392,N_47563,N_47939);
nand U48393 (N_48393,N_47925,N_47789);
xnor U48394 (N_48394,N_47525,N_47881);
and U48395 (N_48395,N_47744,N_47769);
nand U48396 (N_48396,N_47827,N_47571);
or U48397 (N_48397,N_47829,N_47558);
nand U48398 (N_48398,N_47773,N_47764);
nor U48399 (N_48399,N_47617,N_47839);
or U48400 (N_48400,N_47789,N_47967);
xnor U48401 (N_48401,N_47929,N_47531);
nor U48402 (N_48402,N_47563,N_47739);
nor U48403 (N_48403,N_47754,N_47995);
nand U48404 (N_48404,N_47519,N_47524);
xnor U48405 (N_48405,N_47912,N_47511);
or U48406 (N_48406,N_47896,N_47778);
and U48407 (N_48407,N_47638,N_47897);
nand U48408 (N_48408,N_47832,N_47619);
or U48409 (N_48409,N_47829,N_47627);
xor U48410 (N_48410,N_47857,N_47740);
and U48411 (N_48411,N_47798,N_47819);
nor U48412 (N_48412,N_47583,N_47545);
and U48413 (N_48413,N_47785,N_47984);
or U48414 (N_48414,N_47872,N_47617);
xor U48415 (N_48415,N_47992,N_47830);
xor U48416 (N_48416,N_47729,N_47552);
nand U48417 (N_48417,N_47629,N_47914);
or U48418 (N_48418,N_47605,N_47774);
nor U48419 (N_48419,N_47907,N_47619);
xor U48420 (N_48420,N_47839,N_47848);
xor U48421 (N_48421,N_47602,N_47801);
nor U48422 (N_48422,N_47894,N_47783);
xor U48423 (N_48423,N_47862,N_47573);
nor U48424 (N_48424,N_47577,N_47880);
nand U48425 (N_48425,N_47923,N_47984);
xnor U48426 (N_48426,N_47570,N_47584);
and U48427 (N_48427,N_47545,N_47705);
nand U48428 (N_48428,N_47942,N_47886);
or U48429 (N_48429,N_47995,N_47500);
nand U48430 (N_48430,N_47628,N_47992);
xnor U48431 (N_48431,N_47600,N_47984);
xnor U48432 (N_48432,N_47569,N_47943);
nor U48433 (N_48433,N_47997,N_47670);
and U48434 (N_48434,N_47505,N_47760);
and U48435 (N_48435,N_47716,N_47758);
and U48436 (N_48436,N_47546,N_47891);
nand U48437 (N_48437,N_47830,N_47840);
nor U48438 (N_48438,N_47910,N_47730);
xor U48439 (N_48439,N_47870,N_47506);
xor U48440 (N_48440,N_47650,N_47778);
and U48441 (N_48441,N_47843,N_47905);
nand U48442 (N_48442,N_47880,N_47847);
nand U48443 (N_48443,N_47860,N_47638);
nor U48444 (N_48444,N_47820,N_47891);
and U48445 (N_48445,N_47985,N_47576);
and U48446 (N_48446,N_47720,N_47746);
and U48447 (N_48447,N_47616,N_47618);
or U48448 (N_48448,N_47820,N_47901);
nand U48449 (N_48449,N_47934,N_47860);
and U48450 (N_48450,N_47598,N_47535);
or U48451 (N_48451,N_47525,N_47990);
nand U48452 (N_48452,N_47679,N_47765);
nor U48453 (N_48453,N_47951,N_47747);
nor U48454 (N_48454,N_47896,N_47585);
xnor U48455 (N_48455,N_47549,N_47771);
xor U48456 (N_48456,N_47810,N_47540);
or U48457 (N_48457,N_47606,N_47870);
or U48458 (N_48458,N_47548,N_47699);
nor U48459 (N_48459,N_47995,N_47703);
xnor U48460 (N_48460,N_47672,N_47627);
nand U48461 (N_48461,N_47927,N_47953);
nand U48462 (N_48462,N_47605,N_47566);
nand U48463 (N_48463,N_47861,N_47622);
xor U48464 (N_48464,N_47605,N_47827);
nand U48465 (N_48465,N_47773,N_47626);
nor U48466 (N_48466,N_47643,N_47585);
nand U48467 (N_48467,N_47915,N_47623);
and U48468 (N_48468,N_47606,N_47524);
and U48469 (N_48469,N_47604,N_47678);
or U48470 (N_48470,N_47898,N_47735);
xnor U48471 (N_48471,N_47752,N_47985);
nor U48472 (N_48472,N_47689,N_47722);
and U48473 (N_48473,N_47931,N_47694);
nand U48474 (N_48474,N_47905,N_47792);
nor U48475 (N_48475,N_47786,N_47524);
nand U48476 (N_48476,N_47872,N_47828);
and U48477 (N_48477,N_47533,N_47857);
nand U48478 (N_48478,N_47915,N_47769);
nor U48479 (N_48479,N_47944,N_47529);
xor U48480 (N_48480,N_47604,N_47873);
and U48481 (N_48481,N_47603,N_47564);
nand U48482 (N_48482,N_47777,N_47721);
xor U48483 (N_48483,N_47507,N_47770);
nand U48484 (N_48484,N_47899,N_47587);
xnor U48485 (N_48485,N_47664,N_47583);
or U48486 (N_48486,N_47885,N_47634);
nand U48487 (N_48487,N_47557,N_47917);
or U48488 (N_48488,N_47759,N_47516);
nor U48489 (N_48489,N_47938,N_47900);
nor U48490 (N_48490,N_47958,N_47895);
and U48491 (N_48491,N_47790,N_47949);
or U48492 (N_48492,N_47900,N_47563);
nor U48493 (N_48493,N_47605,N_47632);
xor U48494 (N_48494,N_47504,N_47542);
nand U48495 (N_48495,N_47575,N_47587);
nand U48496 (N_48496,N_47899,N_47613);
nor U48497 (N_48497,N_47962,N_47620);
or U48498 (N_48498,N_47899,N_47704);
and U48499 (N_48499,N_47775,N_47605);
or U48500 (N_48500,N_48146,N_48426);
and U48501 (N_48501,N_48471,N_48100);
and U48502 (N_48502,N_48419,N_48250);
xnor U48503 (N_48503,N_48230,N_48240);
or U48504 (N_48504,N_48402,N_48171);
or U48505 (N_48505,N_48179,N_48078);
and U48506 (N_48506,N_48049,N_48016);
xor U48507 (N_48507,N_48125,N_48097);
nor U48508 (N_48508,N_48497,N_48375);
nand U48509 (N_48509,N_48055,N_48270);
xnor U48510 (N_48510,N_48321,N_48103);
or U48511 (N_48511,N_48200,N_48355);
and U48512 (N_48512,N_48371,N_48027);
nor U48513 (N_48513,N_48357,N_48294);
and U48514 (N_48514,N_48316,N_48435);
nor U48515 (N_48515,N_48076,N_48350);
nor U48516 (N_48516,N_48346,N_48204);
nand U48517 (N_48517,N_48446,N_48279);
and U48518 (N_48518,N_48257,N_48247);
or U48519 (N_48519,N_48287,N_48434);
or U48520 (N_48520,N_48369,N_48113);
or U48521 (N_48521,N_48202,N_48351);
or U48522 (N_48522,N_48413,N_48326);
xor U48523 (N_48523,N_48408,N_48142);
and U48524 (N_48524,N_48391,N_48406);
or U48525 (N_48525,N_48198,N_48140);
and U48526 (N_48526,N_48001,N_48324);
nor U48527 (N_48527,N_48168,N_48129);
or U48528 (N_48528,N_48379,N_48207);
nand U48529 (N_48529,N_48105,N_48255);
nor U48530 (N_48530,N_48412,N_48327);
or U48531 (N_48531,N_48094,N_48348);
nand U48532 (N_48532,N_48024,N_48056);
xor U48533 (N_48533,N_48431,N_48482);
nand U48534 (N_48534,N_48491,N_48073);
xnor U48535 (N_48535,N_48269,N_48284);
nor U48536 (N_48536,N_48470,N_48116);
nand U48537 (N_48537,N_48158,N_48473);
or U48538 (N_48538,N_48295,N_48216);
nand U48539 (N_48539,N_48490,N_48147);
nand U48540 (N_48540,N_48188,N_48015);
nor U48541 (N_48541,N_48065,N_48062);
xor U48542 (N_48542,N_48311,N_48137);
nand U48543 (N_48543,N_48252,N_48494);
nand U48544 (N_48544,N_48017,N_48170);
and U48545 (N_48545,N_48231,N_48301);
xnor U48546 (N_48546,N_48075,N_48046);
nand U48547 (N_48547,N_48135,N_48084);
and U48548 (N_48548,N_48468,N_48091);
and U48549 (N_48549,N_48128,N_48288);
or U48550 (N_48550,N_48217,N_48254);
nand U48551 (N_48551,N_48127,N_48420);
nor U48552 (N_48552,N_48069,N_48475);
nor U48553 (N_48553,N_48203,N_48449);
nor U48554 (N_48554,N_48463,N_48349);
xnor U48555 (N_48555,N_48251,N_48368);
or U48556 (N_48556,N_48367,N_48278);
and U48557 (N_48557,N_48372,N_48423);
nand U48558 (N_48558,N_48498,N_48425);
and U48559 (N_48559,N_48436,N_48011);
or U48560 (N_48560,N_48193,N_48130);
or U48561 (N_48561,N_48362,N_48399);
and U48562 (N_48562,N_48150,N_48417);
nor U48563 (N_48563,N_48138,N_48438);
nand U48564 (N_48564,N_48249,N_48134);
or U48565 (N_48565,N_48096,N_48012);
and U48566 (N_48566,N_48044,N_48467);
or U48567 (N_48567,N_48325,N_48430);
and U48568 (N_48568,N_48074,N_48095);
nand U48569 (N_48569,N_48178,N_48403);
xor U48570 (N_48570,N_48256,N_48386);
xnor U48571 (N_48571,N_48364,N_48000);
and U48572 (N_48572,N_48212,N_48036);
and U48573 (N_48573,N_48304,N_48317);
or U48574 (N_48574,N_48154,N_48296);
nor U48575 (N_48575,N_48106,N_48263);
nand U48576 (N_48576,N_48281,N_48102);
or U48577 (N_48577,N_48280,N_48305);
and U48578 (N_48578,N_48159,N_48405);
xnor U48579 (N_48579,N_48167,N_48440);
or U48580 (N_48580,N_48035,N_48308);
nand U48581 (N_48581,N_48225,N_48117);
nand U48582 (N_48582,N_48443,N_48373);
and U48583 (N_48583,N_48291,N_48356);
nand U48584 (N_48584,N_48300,N_48239);
and U48585 (N_48585,N_48002,N_48079);
or U48586 (N_48586,N_48339,N_48397);
nor U48587 (N_48587,N_48233,N_48264);
nand U48588 (N_48588,N_48234,N_48174);
and U48589 (N_48589,N_48298,N_48136);
xnor U48590 (N_48590,N_48019,N_48433);
nor U48591 (N_48591,N_48236,N_48183);
and U48592 (N_48592,N_48465,N_48165);
and U48593 (N_48593,N_48260,N_48126);
or U48594 (N_48594,N_48220,N_48334);
nand U48595 (N_48595,N_48070,N_48029);
xnor U48596 (N_48596,N_48222,N_48041);
nor U48597 (N_48597,N_48336,N_48003);
nor U48598 (N_48598,N_48306,N_48331);
xor U48599 (N_48599,N_48184,N_48313);
xor U48600 (N_48600,N_48427,N_48445);
nand U48601 (N_48601,N_48141,N_48133);
or U48602 (N_48602,N_48424,N_48271);
or U48603 (N_48603,N_48072,N_48007);
nor U48604 (N_48604,N_48447,N_48124);
xor U48605 (N_48605,N_48387,N_48381);
or U48606 (N_48606,N_48428,N_48177);
nor U48607 (N_48607,N_48099,N_48131);
or U48608 (N_48608,N_48223,N_48152);
nor U48609 (N_48609,N_48090,N_48086);
nand U48610 (N_48610,N_48118,N_48458);
nand U48611 (N_48611,N_48378,N_48013);
or U48612 (N_48612,N_48322,N_48329);
xnor U48613 (N_48613,N_48243,N_48415);
and U48614 (N_48614,N_48031,N_48213);
and U48615 (N_48615,N_48196,N_48156);
nor U48616 (N_48616,N_48409,N_48479);
nor U48617 (N_48617,N_48276,N_48347);
xor U48618 (N_48618,N_48407,N_48437);
and U48619 (N_48619,N_48401,N_48476);
or U48620 (N_48620,N_48283,N_48454);
or U48621 (N_48621,N_48400,N_48485);
xor U48622 (N_48622,N_48309,N_48382);
nor U48623 (N_48623,N_48081,N_48089);
or U48624 (N_48624,N_48370,N_48237);
nand U48625 (N_48625,N_48020,N_48104);
nand U48626 (N_48626,N_48120,N_48345);
or U48627 (N_48627,N_48241,N_48459);
xnor U48628 (N_48628,N_48219,N_48008);
nor U48629 (N_48629,N_48450,N_48082);
xor U48630 (N_48630,N_48163,N_48022);
nor U48631 (N_48631,N_48341,N_48010);
or U48632 (N_48632,N_48289,N_48201);
or U48633 (N_48633,N_48277,N_48299);
xnor U48634 (N_48634,N_48330,N_48051);
or U48635 (N_48635,N_48175,N_48115);
nor U48636 (N_48636,N_48315,N_48166);
nand U48637 (N_48637,N_48411,N_48376);
and U48638 (N_48638,N_48366,N_48388);
and U48639 (N_48639,N_48009,N_48209);
or U48640 (N_48640,N_48224,N_48169);
xnor U48641 (N_48641,N_48208,N_48374);
nand U48642 (N_48642,N_48272,N_48048);
xnor U48643 (N_48643,N_48242,N_48034);
and U48644 (N_48644,N_48144,N_48226);
nand U48645 (N_48645,N_48332,N_48145);
nor U48646 (N_48646,N_48197,N_48452);
nor U48647 (N_48647,N_48123,N_48410);
or U48648 (N_48648,N_48395,N_48273);
or U48649 (N_48649,N_48404,N_48181);
nand U48650 (N_48650,N_48499,N_48109);
nor U48651 (N_48651,N_48328,N_48194);
or U48652 (N_48652,N_48229,N_48361);
xor U48653 (N_48653,N_48068,N_48187);
nand U48654 (N_48654,N_48245,N_48061);
and U48655 (N_48655,N_48218,N_48162);
nand U48656 (N_48656,N_48246,N_48121);
nor U48657 (N_48657,N_48492,N_48098);
nand U48658 (N_48658,N_48186,N_48088);
xor U48659 (N_48659,N_48045,N_48483);
xor U48660 (N_48660,N_48344,N_48460);
and U48661 (N_48661,N_48363,N_48032);
nor U48662 (N_48662,N_48195,N_48359);
or U48663 (N_48663,N_48484,N_48493);
xor U48664 (N_48664,N_48337,N_48282);
xor U48665 (N_48665,N_48268,N_48354);
or U48666 (N_48666,N_48478,N_48267);
nor U48667 (N_48667,N_48005,N_48139);
xor U48668 (N_48668,N_48114,N_48489);
nor U48669 (N_48669,N_48083,N_48253);
nor U48670 (N_48670,N_48360,N_48323);
xor U48671 (N_48671,N_48290,N_48108);
and U48672 (N_48672,N_48365,N_48004);
nand U48673 (N_48673,N_48261,N_48414);
or U48674 (N_48674,N_48432,N_48014);
nor U48675 (N_48675,N_48155,N_48066);
xnor U48676 (N_48676,N_48047,N_48172);
nor U48677 (N_48677,N_48101,N_48389);
nand U48678 (N_48678,N_48488,N_48421);
nand U48679 (N_48679,N_48384,N_48059);
xor U48680 (N_48680,N_48173,N_48418);
xor U48681 (N_48681,N_48383,N_48262);
nor U48682 (N_48682,N_48297,N_48353);
xor U48683 (N_48683,N_48235,N_48064);
xnor U48684 (N_48684,N_48248,N_48164);
nand U48685 (N_48685,N_48481,N_48192);
xor U48686 (N_48686,N_48302,N_48040);
and U48687 (N_48687,N_48259,N_48340);
xnor U48688 (N_48688,N_48119,N_48211);
or U48689 (N_48689,N_48333,N_48335);
nor U48690 (N_48690,N_48292,N_48033);
xnor U48691 (N_48691,N_48157,N_48444);
nor U48692 (N_48692,N_48238,N_48028);
nand U48693 (N_48693,N_48205,N_48477);
xnor U48694 (N_48694,N_48352,N_48092);
and U48695 (N_48695,N_48110,N_48451);
nand U48696 (N_48696,N_48377,N_48474);
xor U48697 (N_48697,N_48054,N_48026);
nor U48698 (N_48698,N_48077,N_48380);
nor U48699 (N_48699,N_48176,N_48060);
nor U48700 (N_48700,N_48457,N_48472);
nand U48701 (N_48701,N_48258,N_48416);
nand U48702 (N_48702,N_48053,N_48232);
xor U48703 (N_48703,N_48037,N_48067);
xnor U48704 (N_48704,N_48303,N_48057);
and U48705 (N_48705,N_48392,N_48314);
nor U48706 (N_48706,N_48085,N_48058);
nor U48707 (N_48707,N_48393,N_48151);
or U48708 (N_48708,N_48228,N_48441);
and U48709 (N_48709,N_48191,N_48496);
nand U48710 (N_48710,N_48358,N_48385);
and U48711 (N_48711,N_48453,N_48038);
and U48712 (N_48712,N_48122,N_48093);
and U48713 (N_48713,N_48180,N_48422);
and U48714 (N_48714,N_48265,N_48043);
and U48715 (N_48715,N_48486,N_48442);
and U48716 (N_48716,N_48462,N_48464);
or U48717 (N_48717,N_48244,N_48023);
and U48718 (N_48718,N_48466,N_48087);
or U48719 (N_48719,N_48455,N_48153);
or U48720 (N_48720,N_48293,N_48307);
xor U48721 (N_48721,N_48439,N_48342);
or U48722 (N_48722,N_48050,N_48149);
or U48723 (N_48723,N_48275,N_48111);
xor U48724 (N_48724,N_48206,N_48107);
and U48725 (N_48725,N_48274,N_48456);
xor U48726 (N_48726,N_48338,N_48487);
xnor U48727 (N_48727,N_48063,N_48018);
and U48728 (N_48728,N_48266,N_48461);
nand U48729 (N_48729,N_48030,N_48210);
or U48730 (N_48730,N_48189,N_48396);
or U48731 (N_48731,N_48132,N_48182);
or U48732 (N_48732,N_48319,N_48161);
nor U48733 (N_48733,N_48312,N_48480);
nor U48734 (N_48734,N_48185,N_48310);
xnor U48735 (N_48735,N_48039,N_48143);
and U48736 (N_48736,N_48080,N_48285);
or U48737 (N_48737,N_48221,N_48495);
nor U48738 (N_48738,N_48227,N_48112);
or U48739 (N_48739,N_48429,N_48286);
and U48740 (N_48740,N_48199,N_48021);
and U48741 (N_48741,N_48394,N_48390);
and U48742 (N_48742,N_48148,N_48006);
nand U48743 (N_48743,N_48025,N_48398);
xnor U48744 (N_48744,N_48320,N_48448);
xnor U48745 (N_48745,N_48190,N_48042);
xnor U48746 (N_48746,N_48071,N_48343);
nand U48747 (N_48747,N_48214,N_48052);
xnor U48748 (N_48748,N_48318,N_48160);
nor U48749 (N_48749,N_48469,N_48215);
or U48750 (N_48750,N_48129,N_48297);
or U48751 (N_48751,N_48261,N_48452);
or U48752 (N_48752,N_48459,N_48157);
or U48753 (N_48753,N_48001,N_48038);
nand U48754 (N_48754,N_48363,N_48004);
nand U48755 (N_48755,N_48450,N_48161);
nor U48756 (N_48756,N_48168,N_48429);
xnor U48757 (N_48757,N_48091,N_48029);
nand U48758 (N_48758,N_48096,N_48145);
nand U48759 (N_48759,N_48204,N_48162);
nor U48760 (N_48760,N_48171,N_48428);
nand U48761 (N_48761,N_48395,N_48144);
or U48762 (N_48762,N_48455,N_48173);
xor U48763 (N_48763,N_48055,N_48021);
or U48764 (N_48764,N_48119,N_48402);
xnor U48765 (N_48765,N_48493,N_48277);
or U48766 (N_48766,N_48038,N_48194);
nand U48767 (N_48767,N_48173,N_48027);
nand U48768 (N_48768,N_48323,N_48278);
nor U48769 (N_48769,N_48207,N_48277);
nor U48770 (N_48770,N_48305,N_48379);
xor U48771 (N_48771,N_48071,N_48421);
nand U48772 (N_48772,N_48131,N_48080);
xnor U48773 (N_48773,N_48102,N_48343);
nand U48774 (N_48774,N_48309,N_48410);
and U48775 (N_48775,N_48334,N_48350);
xnor U48776 (N_48776,N_48337,N_48499);
nand U48777 (N_48777,N_48014,N_48019);
xnor U48778 (N_48778,N_48307,N_48439);
nor U48779 (N_48779,N_48207,N_48018);
and U48780 (N_48780,N_48135,N_48430);
and U48781 (N_48781,N_48073,N_48250);
and U48782 (N_48782,N_48380,N_48478);
and U48783 (N_48783,N_48144,N_48048);
and U48784 (N_48784,N_48385,N_48424);
and U48785 (N_48785,N_48431,N_48155);
or U48786 (N_48786,N_48272,N_48168);
and U48787 (N_48787,N_48130,N_48067);
or U48788 (N_48788,N_48114,N_48212);
nor U48789 (N_48789,N_48004,N_48257);
and U48790 (N_48790,N_48089,N_48142);
and U48791 (N_48791,N_48200,N_48190);
xnor U48792 (N_48792,N_48356,N_48459);
xnor U48793 (N_48793,N_48036,N_48268);
or U48794 (N_48794,N_48228,N_48240);
xnor U48795 (N_48795,N_48380,N_48356);
or U48796 (N_48796,N_48098,N_48373);
nor U48797 (N_48797,N_48484,N_48156);
xor U48798 (N_48798,N_48240,N_48252);
xor U48799 (N_48799,N_48439,N_48403);
and U48800 (N_48800,N_48317,N_48242);
xor U48801 (N_48801,N_48347,N_48034);
xor U48802 (N_48802,N_48204,N_48226);
nand U48803 (N_48803,N_48001,N_48213);
nand U48804 (N_48804,N_48032,N_48178);
or U48805 (N_48805,N_48099,N_48407);
and U48806 (N_48806,N_48126,N_48376);
nand U48807 (N_48807,N_48443,N_48413);
xor U48808 (N_48808,N_48308,N_48156);
nor U48809 (N_48809,N_48480,N_48197);
and U48810 (N_48810,N_48097,N_48320);
nand U48811 (N_48811,N_48043,N_48218);
and U48812 (N_48812,N_48290,N_48397);
nand U48813 (N_48813,N_48124,N_48082);
xor U48814 (N_48814,N_48063,N_48130);
and U48815 (N_48815,N_48383,N_48359);
xnor U48816 (N_48816,N_48332,N_48005);
xor U48817 (N_48817,N_48279,N_48061);
and U48818 (N_48818,N_48170,N_48254);
xnor U48819 (N_48819,N_48322,N_48155);
nand U48820 (N_48820,N_48261,N_48486);
and U48821 (N_48821,N_48371,N_48436);
and U48822 (N_48822,N_48009,N_48413);
nor U48823 (N_48823,N_48328,N_48048);
or U48824 (N_48824,N_48386,N_48300);
xnor U48825 (N_48825,N_48306,N_48352);
and U48826 (N_48826,N_48437,N_48077);
nor U48827 (N_48827,N_48229,N_48257);
and U48828 (N_48828,N_48050,N_48473);
xor U48829 (N_48829,N_48323,N_48469);
nor U48830 (N_48830,N_48060,N_48399);
or U48831 (N_48831,N_48472,N_48043);
or U48832 (N_48832,N_48080,N_48290);
xnor U48833 (N_48833,N_48200,N_48385);
nor U48834 (N_48834,N_48213,N_48279);
and U48835 (N_48835,N_48362,N_48037);
xnor U48836 (N_48836,N_48328,N_48391);
nand U48837 (N_48837,N_48152,N_48232);
and U48838 (N_48838,N_48124,N_48490);
nand U48839 (N_48839,N_48432,N_48468);
xnor U48840 (N_48840,N_48093,N_48466);
xor U48841 (N_48841,N_48208,N_48328);
and U48842 (N_48842,N_48267,N_48017);
nand U48843 (N_48843,N_48252,N_48224);
nor U48844 (N_48844,N_48461,N_48341);
xnor U48845 (N_48845,N_48495,N_48346);
xnor U48846 (N_48846,N_48329,N_48097);
or U48847 (N_48847,N_48359,N_48450);
xnor U48848 (N_48848,N_48052,N_48058);
xor U48849 (N_48849,N_48312,N_48464);
and U48850 (N_48850,N_48077,N_48429);
or U48851 (N_48851,N_48060,N_48266);
nand U48852 (N_48852,N_48103,N_48303);
nand U48853 (N_48853,N_48099,N_48389);
xnor U48854 (N_48854,N_48047,N_48152);
xnor U48855 (N_48855,N_48395,N_48349);
and U48856 (N_48856,N_48414,N_48367);
nand U48857 (N_48857,N_48388,N_48104);
nor U48858 (N_48858,N_48031,N_48167);
or U48859 (N_48859,N_48411,N_48374);
nand U48860 (N_48860,N_48174,N_48097);
and U48861 (N_48861,N_48380,N_48425);
or U48862 (N_48862,N_48081,N_48486);
nor U48863 (N_48863,N_48207,N_48426);
and U48864 (N_48864,N_48494,N_48015);
xor U48865 (N_48865,N_48220,N_48358);
nor U48866 (N_48866,N_48074,N_48356);
nor U48867 (N_48867,N_48430,N_48357);
nand U48868 (N_48868,N_48164,N_48367);
nor U48869 (N_48869,N_48284,N_48277);
nand U48870 (N_48870,N_48004,N_48021);
nor U48871 (N_48871,N_48468,N_48430);
and U48872 (N_48872,N_48310,N_48357);
nor U48873 (N_48873,N_48272,N_48080);
nor U48874 (N_48874,N_48193,N_48276);
nor U48875 (N_48875,N_48188,N_48294);
nand U48876 (N_48876,N_48038,N_48182);
and U48877 (N_48877,N_48399,N_48407);
or U48878 (N_48878,N_48375,N_48408);
xnor U48879 (N_48879,N_48361,N_48139);
or U48880 (N_48880,N_48346,N_48444);
xor U48881 (N_48881,N_48221,N_48228);
and U48882 (N_48882,N_48246,N_48410);
nor U48883 (N_48883,N_48056,N_48072);
and U48884 (N_48884,N_48329,N_48444);
or U48885 (N_48885,N_48472,N_48076);
nor U48886 (N_48886,N_48071,N_48095);
nand U48887 (N_48887,N_48427,N_48450);
nor U48888 (N_48888,N_48255,N_48250);
xnor U48889 (N_48889,N_48006,N_48333);
and U48890 (N_48890,N_48106,N_48289);
nand U48891 (N_48891,N_48389,N_48470);
and U48892 (N_48892,N_48271,N_48371);
xnor U48893 (N_48893,N_48307,N_48163);
or U48894 (N_48894,N_48393,N_48351);
and U48895 (N_48895,N_48008,N_48227);
xnor U48896 (N_48896,N_48357,N_48000);
xor U48897 (N_48897,N_48047,N_48440);
nand U48898 (N_48898,N_48360,N_48134);
or U48899 (N_48899,N_48463,N_48311);
xnor U48900 (N_48900,N_48234,N_48171);
nor U48901 (N_48901,N_48172,N_48116);
nand U48902 (N_48902,N_48152,N_48196);
nand U48903 (N_48903,N_48147,N_48474);
and U48904 (N_48904,N_48313,N_48390);
or U48905 (N_48905,N_48390,N_48298);
xor U48906 (N_48906,N_48071,N_48490);
and U48907 (N_48907,N_48175,N_48476);
nor U48908 (N_48908,N_48499,N_48311);
nand U48909 (N_48909,N_48210,N_48376);
and U48910 (N_48910,N_48398,N_48420);
xnor U48911 (N_48911,N_48378,N_48446);
and U48912 (N_48912,N_48245,N_48361);
xnor U48913 (N_48913,N_48347,N_48475);
nor U48914 (N_48914,N_48493,N_48374);
nand U48915 (N_48915,N_48152,N_48072);
nand U48916 (N_48916,N_48092,N_48149);
nand U48917 (N_48917,N_48058,N_48192);
nor U48918 (N_48918,N_48192,N_48030);
xnor U48919 (N_48919,N_48405,N_48125);
nand U48920 (N_48920,N_48011,N_48479);
xnor U48921 (N_48921,N_48158,N_48315);
xor U48922 (N_48922,N_48252,N_48298);
xnor U48923 (N_48923,N_48016,N_48474);
or U48924 (N_48924,N_48007,N_48029);
and U48925 (N_48925,N_48439,N_48325);
and U48926 (N_48926,N_48315,N_48397);
xnor U48927 (N_48927,N_48452,N_48115);
xnor U48928 (N_48928,N_48419,N_48298);
xor U48929 (N_48929,N_48200,N_48131);
or U48930 (N_48930,N_48183,N_48303);
or U48931 (N_48931,N_48310,N_48149);
and U48932 (N_48932,N_48063,N_48353);
or U48933 (N_48933,N_48342,N_48252);
or U48934 (N_48934,N_48488,N_48180);
nand U48935 (N_48935,N_48236,N_48318);
and U48936 (N_48936,N_48186,N_48018);
and U48937 (N_48937,N_48080,N_48225);
nand U48938 (N_48938,N_48143,N_48373);
nor U48939 (N_48939,N_48373,N_48333);
or U48940 (N_48940,N_48446,N_48120);
and U48941 (N_48941,N_48435,N_48485);
and U48942 (N_48942,N_48407,N_48451);
nand U48943 (N_48943,N_48190,N_48328);
or U48944 (N_48944,N_48078,N_48053);
nor U48945 (N_48945,N_48254,N_48462);
and U48946 (N_48946,N_48107,N_48054);
nor U48947 (N_48947,N_48040,N_48365);
nand U48948 (N_48948,N_48292,N_48116);
xnor U48949 (N_48949,N_48002,N_48094);
or U48950 (N_48950,N_48340,N_48234);
nor U48951 (N_48951,N_48372,N_48019);
or U48952 (N_48952,N_48473,N_48384);
nor U48953 (N_48953,N_48438,N_48312);
or U48954 (N_48954,N_48444,N_48393);
or U48955 (N_48955,N_48426,N_48338);
xor U48956 (N_48956,N_48122,N_48004);
or U48957 (N_48957,N_48482,N_48393);
and U48958 (N_48958,N_48490,N_48138);
nand U48959 (N_48959,N_48070,N_48462);
or U48960 (N_48960,N_48015,N_48369);
and U48961 (N_48961,N_48348,N_48083);
nor U48962 (N_48962,N_48220,N_48064);
and U48963 (N_48963,N_48378,N_48125);
xnor U48964 (N_48964,N_48364,N_48292);
or U48965 (N_48965,N_48023,N_48442);
nand U48966 (N_48966,N_48004,N_48458);
nor U48967 (N_48967,N_48224,N_48404);
xor U48968 (N_48968,N_48219,N_48237);
nor U48969 (N_48969,N_48198,N_48476);
nand U48970 (N_48970,N_48271,N_48339);
nand U48971 (N_48971,N_48068,N_48189);
or U48972 (N_48972,N_48095,N_48265);
nand U48973 (N_48973,N_48262,N_48441);
nand U48974 (N_48974,N_48390,N_48281);
nand U48975 (N_48975,N_48273,N_48283);
and U48976 (N_48976,N_48107,N_48113);
and U48977 (N_48977,N_48172,N_48404);
or U48978 (N_48978,N_48374,N_48042);
or U48979 (N_48979,N_48259,N_48203);
and U48980 (N_48980,N_48067,N_48428);
and U48981 (N_48981,N_48326,N_48269);
or U48982 (N_48982,N_48367,N_48347);
xor U48983 (N_48983,N_48113,N_48256);
nor U48984 (N_48984,N_48396,N_48192);
xor U48985 (N_48985,N_48212,N_48342);
xor U48986 (N_48986,N_48264,N_48343);
nor U48987 (N_48987,N_48155,N_48114);
or U48988 (N_48988,N_48365,N_48311);
nor U48989 (N_48989,N_48395,N_48436);
and U48990 (N_48990,N_48042,N_48446);
xnor U48991 (N_48991,N_48353,N_48140);
xnor U48992 (N_48992,N_48399,N_48386);
nor U48993 (N_48993,N_48257,N_48272);
nand U48994 (N_48994,N_48344,N_48353);
xnor U48995 (N_48995,N_48306,N_48491);
xor U48996 (N_48996,N_48098,N_48210);
nor U48997 (N_48997,N_48489,N_48469);
and U48998 (N_48998,N_48363,N_48228);
and U48999 (N_48999,N_48330,N_48409);
nor U49000 (N_49000,N_48713,N_48707);
nand U49001 (N_49001,N_48855,N_48644);
xor U49002 (N_49002,N_48723,N_48887);
nand U49003 (N_49003,N_48654,N_48826);
nor U49004 (N_49004,N_48685,N_48577);
nor U49005 (N_49005,N_48763,N_48529);
xnor U49006 (N_49006,N_48594,N_48878);
nor U49007 (N_49007,N_48542,N_48963);
nor U49008 (N_49008,N_48992,N_48614);
and U49009 (N_49009,N_48744,N_48828);
xnor U49010 (N_49010,N_48576,N_48846);
and U49011 (N_49011,N_48906,N_48950);
and U49012 (N_49012,N_48708,N_48725);
nand U49013 (N_49013,N_48908,N_48554);
nor U49014 (N_49014,N_48520,N_48555);
xor U49015 (N_49015,N_48595,N_48622);
xnor U49016 (N_49016,N_48543,N_48778);
and U49017 (N_49017,N_48736,N_48871);
and U49018 (N_49018,N_48754,N_48663);
or U49019 (N_49019,N_48626,N_48757);
xor U49020 (N_49020,N_48877,N_48617);
nand U49021 (N_49021,N_48774,N_48519);
nor U49022 (N_49022,N_48735,N_48539);
nor U49023 (N_49023,N_48661,N_48967);
nand U49024 (N_49024,N_48810,N_48732);
and U49025 (N_49025,N_48639,N_48602);
or U49026 (N_49026,N_48743,N_48546);
and U49027 (N_49027,N_48730,N_48733);
nand U49028 (N_49028,N_48691,N_48947);
and U49029 (N_49029,N_48958,N_48724);
and U49030 (N_49030,N_48684,N_48690);
and U49031 (N_49031,N_48505,N_48624);
xnor U49032 (N_49032,N_48786,N_48653);
and U49033 (N_49033,N_48728,N_48604);
and U49034 (N_49034,N_48720,N_48836);
nand U49035 (N_49035,N_48775,N_48934);
nor U49036 (N_49036,N_48656,N_48897);
and U49037 (N_49037,N_48813,N_48514);
nor U49038 (N_49038,N_48538,N_48954);
nand U49039 (N_49039,N_48790,N_48985);
nor U49040 (N_49040,N_48640,N_48573);
xor U49041 (N_49041,N_48613,N_48637);
and U49042 (N_49042,N_48843,N_48930);
nor U49043 (N_49043,N_48889,N_48808);
nor U49044 (N_49044,N_48811,N_48799);
or U49045 (N_49045,N_48633,N_48531);
nand U49046 (N_49046,N_48619,N_48578);
nor U49047 (N_49047,N_48581,N_48647);
nand U49048 (N_49048,N_48527,N_48524);
nor U49049 (N_49049,N_48983,N_48590);
and U49050 (N_49050,N_48507,N_48562);
or U49051 (N_49051,N_48956,N_48872);
xor U49052 (N_49052,N_48705,N_48762);
nand U49053 (N_49053,N_48965,N_48829);
nand U49054 (N_49054,N_48945,N_48882);
or U49055 (N_49055,N_48991,N_48921);
nand U49056 (N_49056,N_48847,N_48920);
xor U49057 (N_49057,N_48675,N_48974);
or U49058 (N_49058,N_48597,N_48525);
nor U49059 (N_49059,N_48949,N_48850);
or U49060 (N_49060,N_48816,N_48536);
or U49061 (N_49061,N_48780,N_48839);
xnor U49062 (N_49062,N_48782,N_48729);
nor U49063 (N_49063,N_48596,N_48873);
xor U49064 (N_49064,N_48997,N_48630);
or U49065 (N_49065,N_48643,N_48722);
nand U49066 (N_49066,N_48993,N_48781);
nand U49067 (N_49067,N_48611,N_48669);
and U49068 (N_49068,N_48972,N_48758);
nor U49069 (N_49069,N_48940,N_48900);
xnor U49070 (N_49070,N_48575,N_48612);
and U49071 (N_49071,N_48698,N_48513);
xor U49072 (N_49072,N_48574,N_48794);
nand U49073 (N_49073,N_48541,N_48697);
xnor U49074 (N_49074,N_48858,N_48870);
nand U49075 (N_49075,N_48552,N_48702);
nor U49076 (N_49076,N_48533,N_48506);
xor U49077 (N_49077,N_48941,N_48864);
and U49078 (N_49078,N_48534,N_48608);
nor U49079 (N_49079,N_48986,N_48923);
nor U49080 (N_49080,N_48831,N_48692);
nand U49081 (N_49081,N_48932,N_48746);
nand U49082 (N_49082,N_48951,N_48823);
nand U49083 (N_49083,N_48523,N_48927);
nor U49084 (N_49084,N_48931,N_48634);
and U49085 (N_49085,N_48701,N_48962);
or U49086 (N_49086,N_48571,N_48504);
nor U49087 (N_49087,N_48642,N_48880);
nor U49088 (N_49088,N_48779,N_48838);
and U49089 (N_49089,N_48710,N_48891);
and U49090 (N_49090,N_48537,N_48501);
xor U49091 (N_49091,N_48903,N_48907);
nand U49092 (N_49092,N_48863,N_48544);
xor U49093 (N_49093,N_48756,N_48764);
or U49094 (N_49094,N_48511,N_48977);
nor U49095 (N_49095,N_48586,N_48750);
and U49096 (N_49096,N_48984,N_48600);
or U49097 (N_49097,N_48717,N_48580);
or U49098 (N_49098,N_48579,N_48771);
xnor U49099 (N_49099,N_48645,N_48902);
xnor U49100 (N_49100,N_48973,N_48748);
nand U49101 (N_49101,N_48709,N_48638);
nand U49102 (N_49102,N_48801,N_48671);
xnor U49103 (N_49103,N_48535,N_48752);
xnor U49104 (N_49104,N_48564,N_48959);
nor U49105 (N_49105,N_48727,N_48686);
and U49106 (N_49106,N_48584,N_48960);
and U49107 (N_49107,N_48944,N_48568);
xnor U49108 (N_49108,N_48726,N_48910);
nor U49109 (N_49109,N_48755,N_48500);
nand U49110 (N_49110,N_48657,N_48696);
nand U49111 (N_49111,N_48901,N_48857);
and U49112 (N_49112,N_48936,N_48812);
nand U49113 (N_49113,N_48526,N_48515);
nand U49114 (N_49114,N_48912,N_48517);
xor U49115 (N_49115,N_48933,N_48817);
and U49116 (N_49116,N_48745,N_48769);
and U49117 (N_49117,N_48737,N_48770);
xnor U49118 (N_49118,N_48946,N_48704);
or U49119 (N_49119,N_48868,N_48678);
nand U49120 (N_49120,N_48673,N_48913);
xor U49121 (N_49121,N_48740,N_48783);
nor U49122 (N_49122,N_48802,N_48818);
nor U49123 (N_49123,N_48522,N_48830);
or U49124 (N_49124,N_48618,N_48567);
xor U49125 (N_49125,N_48674,N_48650);
or U49126 (N_49126,N_48942,N_48588);
nand U49127 (N_49127,N_48854,N_48917);
nand U49128 (N_49128,N_48631,N_48648);
and U49129 (N_49129,N_48890,N_48844);
nand U49130 (N_49130,N_48841,N_48955);
xnor U49131 (N_49131,N_48978,N_48593);
or U49132 (N_49132,N_48919,N_48659);
xnor U49133 (N_49133,N_48556,N_48591);
or U49134 (N_49134,N_48925,N_48609);
xnor U49135 (N_49135,N_48892,N_48687);
and U49136 (N_49136,N_48582,N_48821);
or U49137 (N_49137,N_48845,N_48560);
and U49138 (N_49138,N_48970,N_48881);
nand U49139 (N_49139,N_48558,N_48865);
and U49140 (N_49140,N_48867,N_48952);
nor U49141 (N_49141,N_48918,N_48767);
nand U49142 (N_49142,N_48738,N_48939);
xnor U49143 (N_49143,N_48922,N_48599);
nand U49144 (N_49144,N_48512,N_48566);
xnor U49145 (N_49145,N_48924,N_48785);
nor U49146 (N_49146,N_48563,N_48875);
nand U49147 (N_49147,N_48979,N_48834);
and U49148 (N_49148,N_48587,N_48787);
xnor U49149 (N_49149,N_48603,N_48721);
and U49150 (N_49150,N_48893,N_48625);
xor U49151 (N_49151,N_48565,N_48938);
or U49152 (N_49152,N_48937,N_48935);
and U49153 (N_49153,N_48928,N_48646);
nand U49154 (N_49154,N_48916,N_48885);
or U49155 (N_49155,N_48607,N_48987);
nand U49156 (N_49156,N_48876,N_48549);
nor U49157 (N_49157,N_48888,N_48852);
and U49158 (N_49158,N_48508,N_48683);
and U49159 (N_49159,N_48688,N_48840);
or U49160 (N_49160,N_48861,N_48716);
xor U49161 (N_49161,N_48772,N_48976);
nor U49162 (N_49162,N_48825,N_48996);
xor U49163 (N_49163,N_48819,N_48518);
nor U49164 (N_49164,N_48773,N_48814);
xnor U49165 (N_49165,N_48589,N_48851);
nor U49166 (N_49166,N_48966,N_48975);
nor U49167 (N_49167,N_48712,N_48879);
xor U49168 (N_49168,N_48895,N_48585);
nor U49169 (N_49169,N_48667,N_48820);
or U49170 (N_49170,N_48760,N_48822);
nand U49171 (N_49171,N_48793,N_48884);
or U49172 (N_49172,N_48551,N_48547);
xnor U49173 (N_49173,N_48766,N_48695);
or U49174 (N_49174,N_48809,N_48741);
and U49175 (N_49175,N_48957,N_48968);
or U49176 (N_49176,N_48789,N_48623);
and U49177 (N_49177,N_48776,N_48605);
nand U49178 (N_49178,N_48896,N_48971);
and U49179 (N_49179,N_48929,N_48768);
nor U49180 (N_49180,N_48503,N_48718);
xor U49181 (N_49181,N_48693,N_48849);
xor U49182 (N_49182,N_48570,N_48837);
or U49183 (N_49183,N_48824,N_48502);
or U49184 (N_49184,N_48635,N_48886);
or U49185 (N_49185,N_48805,N_48699);
nor U49186 (N_49186,N_48677,N_48679);
nor U49187 (N_49187,N_48550,N_48859);
xor U49188 (N_49188,N_48803,N_48703);
nand U49189 (N_49189,N_48636,N_48649);
nor U49190 (N_49190,N_48689,N_48658);
nand U49191 (N_49191,N_48791,N_48777);
xnor U49192 (N_49192,N_48681,N_48714);
or U49193 (N_49193,N_48860,N_48797);
nand U49194 (N_49194,N_48989,N_48516);
and U49195 (N_49195,N_48761,N_48994);
nor U49196 (N_49196,N_48827,N_48628);
xor U49197 (N_49197,N_48682,N_48530);
or U49198 (N_49198,N_48795,N_48545);
nand U49199 (N_49199,N_48742,N_48680);
xnor U49200 (N_49200,N_48660,N_48666);
and U49201 (N_49201,N_48751,N_48601);
or U49202 (N_49202,N_48842,N_48961);
xor U49203 (N_49203,N_48853,N_48981);
nor U49204 (N_49204,N_48615,N_48665);
nand U49205 (N_49205,N_48784,N_48672);
nand U49206 (N_49206,N_48806,N_48610);
or U49207 (N_49207,N_48909,N_48749);
nor U49208 (N_49208,N_48676,N_48598);
nand U49209 (N_49209,N_48969,N_48641);
nor U49210 (N_49210,N_48739,N_48670);
or U49211 (N_49211,N_48548,N_48583);
or U49212 (N_49212,N_48621,N_48627);
xnor U49213 (N_49213,N_48964,N_48606);
or U49214 (N_49214,N_48616,N_48796);
and U49215 (N_49215,N_48798,N_48668);
xor U49216 (N_49216,N_48528,N_48553);
and U49217 (N_49217,N_48804,N_48559);
nand U49218 (N_49218,N_48700,N_48835);
or U49219 (N_49219,N_48569,N_48800);
nor U49220 (N_49220,N_48655,N_48572);
nor U49221 (N_49221,N_48869,N_48731);
xnor U49222 (N_49222,N_48561,N_48894);
nand U49223 (N_49223,N_48747,N_48651);
xor U49224 (N_49224,N_48982,N_48532);
nand U49225 (N_49225,N_48943,N_48706);
nor U49226 (N_49226,N_48856,N_48899);
and U49227 (N_49227,N_48664,N_48914);
nor U49228 (N_49228,N_48832,N_48629);
xor U49229 (N_49229,N_48711,N_48521);
and U49230 (N_49230,N_48620,N_48948);
nor U49231 (N_49231,N_48999,N_48995);
nand U49232 (N_49232,N_48765,N_48848);
nor U49233 (N_49233,N_48874,N_48990);
or U49234 (N_49234,N_48915,N_48592);
nand U49235 (N_49235,N_48557,N_48862);
xnor U49236 (N_49236,N_48807,N_48926);
nor U49237 (N_49237,N_48734,N_48998);
nand U49238 (N_49238,N_48815,N_48883);
nand U49239 (N_49239,N_48980,N_48759);
and U49240 (N_49240,N_48866,N_48905);
nand U49241 (N_49241,N_48715,N_48652);
nand U49242 (N_49242,N_48898,N_48719);
nand U49243 (N_49243,N_48833,N_48509);
nor U49244 (N_49244,N_48911,N_48904);
nand U49245 (N_49245,N_48988,N_48540);
and U49246 (N_49246,N_48510,N_48662);
or U49247 (N_49247,N_48792,N_48694);
xor U49248 (N_49248,N_48953,N_48632);
xnor U49249 (N_49249,N_48788,N_48753);
and U49250 (N_49250,N_48941,N_48681);
nand U49251 (N_49251,N_48869,N_48607);
or U49252 (N_49252,N_48598,N_48698);
nand U49253 (N_49253,N_48937,N_48548);
nor U49254 (N_49254,N_48543,N_48970);
xor U49255 (N_49255,N_48728,N_48787);
xnor U49256 (N_49256,N_48546,N_48500);
nand U49257 (N_49257,N_48927,N_48673);
nor U49258 (N_49258,N_48701,N_48606);
and U49259 (N_49259,N_48604,N_48528);
nand U49260 (N_49260,N_48742,N_48660);
or U49261 (N_49261,N_48875,N_48787);
nor U49262 (N_49262,N_48843,N_48772);
or U49263 (N_49263,N_48679,N_48794);
nand U49264 (N_49264,N_48999,N_48583);
or U49265 (N_49265,N_48726,N_48582);
nand U49266 (N_49266,N_48921,N_48755);
xnor U49267 (N_49267,N_48945,N_48755);
nor U49268 (N_49268,N_48845,N_48767);
nand U49269 (N_49269,N_48724,N_48911);
nor U49270 (N_49270,N_48708,N_48805);
nor U49271 (N_49271,N_48892,N_48712);
or U49272 (N_49272,N_48549,N_48935);
xnor U49273 (N_49273,N_48691,N_48587);
and U49274 (N_49274,N_48536,N_48854);
nand U49275 (N_49275,N_48718,N_48664);
and U49276 (N_49276,N_48667,N_48912);
and U49277 (N_49277,N_48944,N_48906);
nor U49278 (N_49278,N_48736,N_48501);
xor U49279 (N_49279,N_48723,N_48576);
and U49280 (N_49280,N_48706,N_48721);
nor U49281 (N_49281,N_48671,N_48641);
nand U49282 (N_49282,N_48580,N_48755);
xnor U49283 (N_49283,N_48549,N_48917);
nand U49284 (N_49284,N_48875,N_48560);
and U49285 (N_49285,N_48759,N_48725);
nand U49286 (N_49286,N_48881,N_48804);
xor U49287 (N_49287,N_48928,N_48581);
or U49288 (N_49288,N_48826,N_48942);
and U49289 (N_49289,N_48797,N_48850);
and U49290 (N_49290,N_48724,N_48764);
nor U49291 (N_49291,N_48803,N_48814);
and U49292 (N_49292,N_48562,N_48794);
and U49293 (N_49293,N_48874,N_48964);
and U49294 (N_49294,N_48752,N_48698);
xnor U49295 (N_49295,N_48725,N_48818);
or U49296 (N_49296,N_48836,N_48601);
xnor U49297 (N_49297,N_48606,N_48556);
and U49298 (N_49298,N_48756,N_48941);
and U49299 (N_49299,N_48535,N_48662);
or U49300 (N_49300,N_48640,N_48950);
nand U49301 (N_49301,N_48984,N_48752);
or U49302 (N_49302,N_48866,N_48544);
nor U49303 (N_49303,N_48876,N_48994);
nor U49304 (N_49304,N_48709,N_48726);
nand U49305 (N_49305,N_48831,N_48766);
and U49306 (N_49306,N_48945,N_48598);
xnor U49307 (N_49307,N_48936,N_48593);
xor U49308 (N_49308,N_48678,N_48782);
xor U49309 (N_49309,N_48823,N_48761);
nand U49310 (N_49310,N_48670,N_48592);
or U49311 (N_49311,N_48807,N_48826);
nand U49312 (N_49312,N_48597,N_48512);
and U49313 (N_49313,N_48550,N_48566);
and U49314 (N_49314,N_48740,N_48742);
xor U49315 (N_49315,N_48863,N_48905);
nor U49316 (N_49316,N_48629,N_48815);
or U49317 (N_49317,N_48906,N_48788);
nand U49318 (N_49318,N_48830,N_48788);
nand U49319 (N_49319,N_48913,N_48637);
xor U49320 (N_49320,N_48763,N_48989);
or U49321 (N_49321,N_48877,N_48811);
xnor U49322 (N_49322,N_48613,N_48622);
nor U49323 (N_49323,N_48668,N_48710);
or U49324 (N_49324,N_48509,N_48605);
nor U49325 (N_49325,N_48830,N_48787);
and U49326 (N_49326,N_48690,N_48849);
or U49327 (N_49327,N_48896,N_48590);
and U49328 (N_49328,N_48519,N_48823);
and U49329 (N_49329,N_48896,N_48652);
nand U49330 (N_49330,N_48662,N_48955);
or U49331 (N_49331,N_48795,N_48993);
xnor U49332 (N_49332,N_48562,N_48941);
nand U49333 (N_49333,N_48890,N_48756);
xor U49334 (N_49334,N_48798,N_48889);
nor U49335 (N_49335,N_48812,N_48754);
nand U49336 (N_49336,N_48778,N_48985);
and U49337 (N_49337,N_48942,N_48720);
and U49338 (N_49338,N_48596,N_48517);
and U49339 (N_49339,N_48899,N_48568);
xor U49340 (N_49340,N_48919,N_48547);
and U49341 (N_49341,N_48833,N_48607);
nand U49342 (N_49342,N_48950,N_48690);
nand U49343 (N_49343,N_48909,N_48779);
or U49344 (N_49344,N_48841,N_48866);
xor U49345 (N_49345,N_48756,N_48913);
nor U49346 (N_49346,N_48560,N_48796);
and U49347 (N_49347,N_48780,N_48801);
or U49348 (N_49348,N_48718,N_48859);
xnor U49349 (N_49349,N_48509,N_48626);
and U49350 (N_49350,N_48889,N_48566);
and U49351 (N_49351,N_48506,N_48532);
nor U49352 (N_49352,N_48506,N_48818);
xnor U49353 (N_49353,N_48669,N_48896);
or U49354 (N_49354,N_48853,N_48518);
or U49355 (N_49355,N_48783,N_48598);
nand U49356 (N_49356,N_48719,N_48587);
nor U49357 (N_49357,N_48672,N_48743);
nor U49358 (N_49358,N_48607,N_48956);
xor U49359 (N_49359,N_48746,N_48941);
nor U49360 (N_49360,N_48864,N_48881);
nor U49361 (N_49361,N_48873,N_48641);
nor U49362 (N_49362,N_48704,N_48526);
and U49363 (N_49363,N_48519,N_48695);
or U49364 (N_49364,N_48872,N_48600);
and U49365 (N_49365,N_48605,N_48548);
and U49366 (N_49366,N_48872,N_48599);
nand U49367 (N_49367,N_48750,N_48597);
or U49368 (N_49368,N_48662,N_48749);
nor U49369 (N_49369,N_48556,N_48868);
or U49370 (N_49370,N_48623,N_48726);
and U49371 (N_49371,N_48608,N_48630);
xor U49372 (N_49372,N_48607,N_48523);
nand U49373 (N_49373,N_48938,N_48944);
xor U49374 (N_49374,N_48572,N_48948);
and U49375 (N_49375,N_48641,N_48636);
nand U49376 (N_49376,N_48904,N_48640);
and U49377 (N_49377,N_48936,N_48783);
nand U49378 (N_49378,N_48900,N_48526);
and U49379 (N_49379,N_48859,N_48816);
or U49380 (N_49380,N_48690,N_48947);
nor U49381 (N_49381,N_48516,N_48661);
nor U49382 (N_49382,N_48794,N_48942);
nor U49383 (N_49383,N_48555,N_48995);
and U49384 (N_49384,N_48871,N_48713);
nor U49385 (N_49385,N_48976,N_48752);
and U49386 (N_49386,N_48768,N_48775);
nand U49387 (N_49387,N_48529,N_48941);
nor U49388 (N_49388,N_48854,N_48639);
xnor U49389 (N_49389,N_48904,N_48521);
or U49390 (N_49390,N_48640,N_48988);
xor U49391 (N_49391,N_48896,N_48897);
and U49392 (N_49392,N_48980,N_48714);
or U49393 (N_49393,N_48590,N_48903);
nor U49394 (N_49394,N_48828,N_48908);
xor U49395 (N_49395,N_48859,N_48768);
nand U49396 (N_49396,N_48943,N_48514);
or U49397 (N_49397,N_48937,N_48952);
or U49398 (N_49398,N_48547,N_48582);
and U49399 (N_49399,N_48535,N_48700);
and U49400 (N_49400,N_48530,N_48930);
xnor U49401 (N_49401,N_48755,N_48797);
or U49402 (N_49402,N_48641,N_48537);
and U49403 (N_49403,N_48960,N_48520);
nand U49404 (N_49404,N_48630,N_48983);
and U49405 (N_49405,N_48940,N_48575);
or U49406 (N_49406,N_48567,N_48570);
or U49407 (N_49407,N_48526,N_48795);
or U49408 (N_49408,N_48765,N_48651);
or U49409 (N_49409,N_48794,N_48984);
nor U49410 (N_49410,N_48717,N_48568);
xor U49411 (N_49411,N_48640,N_48656);
or U49412 (N_49412,N_48639,N_48536);
or U49413 (N_49413,N_48870,N_48748);
xor U49414 (N_49414,N_48719,N_48759);
nand U49415 (N_49415,N_48790,N_48771);
xnor U49416 (N_49416,N_48782,N_48600);
nand U49417 (N_49417,N_48876,N_48633);
nor U49418 (N_49418,N_48585,N_48905);
and U49419 (N_49419,N_48863,N_48736);
nor U49420 (N_49420,N_48790,N_48703);
xor U49421 (N_49421,N_48990,N_48841);
and U49422 (N_49422,N_48666,N_48977);
xnor U49423 (N_49423,N_48993,N_48843);
xnor U49424 (N_49424,N_48694,N_48702);
nand U49425 (N_49425,N_48952,N_48812);
and U49426 (N_49426,N_48957,N_48986);
or U49427 (N_49427,N_48510,N_48886);
and U49428 (N_49428,N_48862,N_48980);
or U49429 (N_49429,N_48686,N_48852);
and U49430 (N_49430,N_48661,N_48836);
nor U49431 (N_49431,N_48616,N_48870);
or U49432 (N_49432,N_48745,N_48705);
or U49433 (N_49433,N_48519,N_48822);
nor U49434 (N_49434,N_48512,N_48778);
nand U49435 (N_49435,N_48616,N_48923);
xor U49436 (N_49436,N_48768,N_48757);
or U49437 (N_49437,N_48500,N_48942);
and U49438 (N_49438,N_48604,N_48713);
nor U49439 (N_49439,N_48620,N_48552);
nand U49440 (N_49440,N_48573,N_48788);
xor U49441 (N_49441,N_48500,N_48791);
or U49442 (N_49442,N_48800,N_48647);
nor U49443 (N_49443,N_48983,N_48707);
nand U49444 (N_49444,N_48958,N_48508);
and U49445 (N_49445,N_48560,N_48896);
nand U49446 (N_49446,N_48553,N_48686);
or U49447 (N_49447,N_48852,N_48764);
xor U49448 (N_49448,N_48549,N_48502);
and U49449 (N_49449,N_48795,N_48701);
nand U49450 (N_49450,N_48823,N_48974);
nor U49451 (N_49451,N_48635,N_48556);
xor U49452 (N_49452,N_48545,N_48555);
nand U49453 (N_49453,N_48916,N_48881);
or U49454 (N_49454,N_48726,N_48802);
nor U49455 (N_49455,N_48568,N_48606);
and U49456 (N_49456,N_48959,N_48784);
and U49457 (N_49457,N_48996,N_48754);
and U49458 (N_49458,N_48702,N_48510);
and U49459 (N_49459,N_48588,N_48768);
nand U49460 (N_49460,N_48685,N_48895);
nor U49461 (N_49461,N_48886,N_48800);
or U49462 (N_49462,N_48854,N_48690);
xnor U49463 (N_49463,N_48649,N_48593);
and U49464 (N_49464,N_48518,N_48622);
and U49465 (N_49465,N_48936,N_48866);
or U49466 (N_49466,N_48897,N_48932);
and U49467 (N_49467,N_48551,N_48624);
and U49468 (N_49468,N_48564,N_48602);
nand U49469 (N_49469,N_48655,N_48778);
or U49470 (N_49470,N_48727,N_48827);
and U49471 (N_49471,N_48755,N_48683);
and U49472 (N_49472,N_48842,N_48882);
or U49473 (N_49473,N_48845,N_48509);
xnor U49474 (N_49474,N_48918,N_48822);
nand U49475 (N_49475,N_48977,N_48659);
nor U49476 (N_49476,N_48963,N_48810);
nand U49477 (N_49477,N_48910,N_48766);
nand U49478 (N_49478,N_48605,N_48958);
or U49479 (N_49479,N_48929,N_48842);
nor U49480 (N_49480,N_48900,N_48854);
or U49481 (N_49481,N_48900,N_48517);
and U49482 (N_49482,N_48572,N_48654);
nor U49483 (N_49483,N_48607,N_48558);
nor U49484 (N_49484,N_48558,N_48949);
xnor U49485 (N_49485,N_48825,N_48619);
xor U49486 (N_49486,N_48655,N_48964);
and U49487 (N_49487,N_48993,N_48531);
or U49488 (N_49488,N_48755,N_48896);
or U49489 (N_49489,N_48699,N_48550);
nand U49490 (N_49490,N_48961,N_48591);
and U49491 (N_49491,N_48917,N_48831);
nand U49492 (N_49492,N_48876,N_48631);
and U49493 (N_49493,N_48759,N_48584);
nor U49494 (N_49494,N_48575,N_48705);
nand U49495 (N_49495,N_48962,N_48957);
or U49496 (N_49496,N_48645,N_48726);
nor U49497 (N_49497,N_48620,N_48950);
nor U49498 (N_49498,N_48670,N_48685);
or U49499 (N_49499,N_48926,N_48654);
or U49500 (N_49500,N_49067,N_49027);
xor U49501 (N_49501,N_49118,N_49452);
or U49502 (N_49502,N_49229,N_49456);
xor U49503 (N_49503,N_49003,N_49465);
or U49504 (N_49504,N_49442,N_49000);
nand U49505 (N_49505,N_49315,N_49162);
nor U49506 (N_49506,N_49417,N_49158);
and U49507 (N_49507,N_49490,N_49254);
and U49508 (N_49508,N_49450,N_49266);
nor U49509 (N_49509,N_49097,N_49296);
nand U49510 (N_49510,N_49121,N_49291);
and U49511 (N_49511,N_49420,N_49068);
xor U49512 (N_49512,N_49077,N_49086);
nand U49513 (N_49513,N_49186,N_49089);
nand U49514 (N_49514,N_49279,N_49478);
xor U49515 (N_49515,N_49366,N_49409);
nor U49516 (N_49516,N_49245,N_49183);
xnor U49517 (N_49517,N_49455,N_49047);
or U49518 (N_49518,N_49091,N_49081);
or U49519 (N_49519,N_49459,N_49070);
and U49520 (N_49520,N_49334,N_49428);
nand U49521 (N_49521,N_49078,N_49221);
xnor U49522 (N_49522,N_49485,N_49104);
and U49523 (N_49523,N_49230,N_49395);
xnor U49524 (N_49524,N_49069,N_49298);
and U49525 (N_49525,N_49423,N_49033);
and U49526 (N_49526,N_49458,N_49481);
nor U49527 (N_49527,N_49405,N_49177);
xnor U49528 (N_49528,N_49484,N_49325);
nor U49529 (N_49529,N_49468,N_49361);
nand U49530 (N_49530,N_49055,N_49140);
nor U49531 (N_49531,N_49268,N_49176);
nand U49532 (N_49532,N_49493,N_49318);
nand U49533 (N_49533,N_49333,N_49220);
nand U49534 (N_49534,N_49382,N_49276);
nor U49535 (N_49535,N_49256,N_49253);
or U49536 (N_49536,N_49262,N_49107);
nand U49537 (N_49537,N_49153,N_49208);
or U49538 (N_49538,N_49150,N_49083);
xor U49539 (N_49539,N_49397,N_49402);
xnor U49540 (N_49540,N_49418,N_49320);
xnor U49541 (N_49541,N_49377,N_49356);
nand U49542 (N_49542,N_49426,N_49292);
nor U49543 (N_49543,N_49005,N_49168);
and U49544 (N_49544,N_49084,N_49042);
xor U49545 (N_49545,N_49330,N_49212);
nor U49546 (N_49546,N_49322,N_49011);
xnor U49547 (N_49547,N_49421,N_49358);
nand U49548 (N_49548,N_49443,N_49057);
nor U49549 (N_49549,N_49154,N_49191);
nand U49550 (N_49550,N_49036,N_49437);
and U49551 (N_49551,N_49235,N_49422);
nor U49552 (N_49552,N_49317,N_49297);
and U49553 (N_49553,N_49149,N_49102);
nor U49554 (N_49554,N_49441,N_49095);
xor U49555 (N_49555,N_49270,N_49376);
xor U49556 (N_49556,N_49280,N_49314);
nand U49557 (N_49557,N_49157,N_49406);
nand U49558 (N_49558,N_49049,N_49407);
nor U49559 (N_49559,N_49217,N_49136);
nor U49560 (N_49560,N_49006,N_49340);
nor U49561 (N_49561,N_49338,N_49213);
nand U49562 (N_49562,N_49277,N_49462);
and U49563 (N_49563,N_49088,N_49483);
nor U49564 (N_49564,N_49263,N_49093);
xor U49565 (N_49565,N_49174,N_49375);
or U49566 (N_49566,N_49160,N_49087);
or U49567 (N_49567,N_49211,N_49059);
nand U49568 (N_49568,N_49147,N_49109);
or U49569 (N_49569,N_49165,N_49449);
nor U49570 (N_49570,N_49497,N_49223);
and U49571 (N_49571,N_49299,N_49438);
and U49572 (N_49572,N_49373,N_49415);
nor U49573 (N_49573,N_49370,N_49400);
and U49574 (N_49574,N_49075,N_49085);
xor U49575 (N_49575,N_49020,N_49013);
or U49576 (N_49576,N_49463,N_49066);
or U49577 (N_49577,N_49293,N_49196);
nand U49578 (N_49578,N_49192,N_49264);
or U49579 (N_49579,N_49362,N_49473);
and U49580 (N_49580,N_49024,N_49106);
nand U49581 (N_49581,N_49274,N_49134);
nor U49582 (N_49582,N_49239,N_49344);
nor U49583 (N_49583,N_49319,N_49430);
nand U49584 (N_49584,N_49404,N_49275);
or U49585 (N_49585,N_49349,N_49294);
xor U49586 (N_49586,N_49413,N_49265);
nor U49587 (N_49587,N_49019,N_49058);
xnor U49588 (N_49588,N_49489,N_49152);
and U49589 (N_49589,N_49328,N_49063);
xor U49590 (N_49590,N_49074,N_49123);
xor U49591 (N_49591,N_49201,N_49359);
xnor U49592 (N_49592,N_49092,N_49453);
xnor U49593 (N_49593,N_49060,N_49243);
nand U49594 (N_49594,N_49311,N_49030);
xnor U49595 (N_49595,N_49210,N_49342);
or U49596 (N_49596,N_49029,N_49414);
nand U49597 (N_49597,N_49015,N_49278);
nor U49598 (N_49598,N_49146,N_49203);
nor U49599 (N_49599,N_49495,N_49159);
and U49600 (N_49600,N_49371,N_49347);
and U49601 (N_49601,N_49491,N_49173);
nor U49602 (N_49602,N_49145,N_49480);
nor U49603 (N_49603,N_49002,N_49339);
and U49604 (N_49604,N_49304,N_49166);
xor U49605 (N_49605,N_49050,N_49008);
and U49606 (N_49606,N_49215,N_49143);
or U49607 (N_49607,N_49350,N_49197);
xnor U49608 (N_49608,N_49130,N_49273);
xnor U49609 (N_49609,N_49228,N_49242);
nand U49610 (N_49610,N_49431,N_49269);
nand U49611 (N_49611,N_49044,N_49206);
nor U49612 (N_49612,N_49290,N_49461);
nand U49613 (N_49613,N_49064,N_49188);
or U49614 (N_49614,N_49101,N_49281);
nor U49615 (N_49615,N_49255,N_49457);
nand U49616 (N_49616,N_49026,N_49062);
nor U49617 (N_49617,N_49259,N_49378);
and U49618 (N_49618,N_49038,N_49045);
nor U49619 (N_49619,N_49393,N_49306);
nand U49620 (N_49620,N_49122,N_49351);
xnor U49621 (N_49621,N_49394,N_49469);
or U49622 (N_49622,N_49194,N_49240);
and U49623 (N_49623,N_49103,N_49261);
and U49624 (N_49624,N_49331,N_49301);
nor U49625 (N_49625,N_49224,N_49336);
or U49626 (N_49626,N_49127,N_49303);
xnor U49627 (N_49627,N_49234,N_49267);
nand U49628 (N_49628,N_49392,N_49214);
and U49629 (N_49629,N_49028,N_49182);
nor U49630 (N_49630,N_49219,N_49079);
xor U49631 (N_49631,N_49094,N_49238);
xor U49632 (N_49632,N_49052,N_49425);
or U49633 (N_49633,N_49360,N_49236);
nor U49634 (N_49634,N_49329,N_49148);
xor U49635 (N_49635,N_49039,N_49445);
xor U49636 (N_49636,N_49424,N_49372);
nand U49637 (N_49637,N_49113,N_49477);
nand U49638 (N_49638,N_49040,N_49471);
or U49639 (N_49639,N_49337,N_49341);
xor U49640 (N_49640,N_49482,N_49218);
nor U49641 (N_49641,N_49385,N_49499);
and U49642 (N_49642,N_49369,N_49383);
and U49643 (N_49643,N_49009,N_49012);
or U49644 (N_49644,N_49169,N_49429);
or U49645 (N_49645,N_49401,N_49053);
and U49646 (N_49646,N_49111,N_49474);
and U49647 (N_49647,N_49467,N_49312);
xnor U49648 (N_49648,N_49161,N_49117);
nor U49649 (N_49649,N_49454,N_49380);
nor U49650 (N_49650,N_49014,N_49048);
nor U49651 (N_49651,N_49129,N_49295);
nand U49652 (N_49652,N_49357,N_49248);
xnor U49653 (N_49653,N_49282,N_49171);
and U49654 (N_49654,N_49017,N_49225);
nor U49655 (N_49655,N_49112,N_49387);
xnor U49656 (N_49656,N_49080,N_49151);
or U49657 (N_49657,N_49435,N_49163);
nor U49658 (N_49658,N_49105,N_49323);
nand U49659 (N_49659,N_49249,N_49226);
nand U49660 (N_49660,N_49410,N_49364);
or U49661 (N_49661,N_49302,N_49142);
nand U49662 (N_49662,N_49260,N_49365);
xor U49663 (N_49663,N_49222,N_49326);
or U49664 (N_49664,N_49004,N_49444);
nor U49665 (N_49665,N_49185,N_49283);
nor U49666 (N_49666,N_49167,N_49252);
nand U49667 (N_49667,N_49175,N_49309);
and U49668 (N_49668,N_49300,N_49310);
or U49669 (N_49669,N_49355,N_49195);
nor U49670 (N_49670,N_49436,N_49204);
xnor U49671 (N_49671,N_49416,N_49324);
xor U49672 (N_49672,N_49216,N_49287);
and U49673 (N_49673,N_49363,N_49272);
and U49674 (N_49674,N_49466,N_49010);
and U49675 (N_49675,N_49018,N_49200);
or U49676 (N_49676,N_49403,N_49479);
nor U49677 (N_49677,N_49021,N_49498);
and U49678 (N_49678,N_49396,N_49247);
and U49679 (N_49679,N_49427,N_49389);
xor U49680 (N_49680,N_49419,N_49307);
nor U49681 (N_49681,N_49205,N_49139);
or U49682 (N_49682,N_49155,N_49446);
nor U49683 (N_49683,N_49316,N_49284);
or U49684 (N_49684,N_49043,N_49348);
nand U49685 (N_49685,N_49335,N_49072);
or U49686 (N_49686,N_49390,N_49022);
nor U49687 (N_49687,N_49286,N_49170);
and U49688 (N_49688,N_49031,N_49202);
nor U49689 (N_49689,N_49232,N_49399);
and U49690 (N_49690,N_49308,N_49007);
nor U49691 (N_49691,N_49156,N_49061);
nor U49692 (N_49692,N_49354,N_49180);
xor U49693 (N_49693,N_49076,N_49189);
nor U49694 (N_49694,N_49071,N_49131);
and U49695 (N_49695,N_49037,N_49411);
and U49696 (N_49696,N_49137,N_49001);
and U49697 (N_49697,N_49190,N_49492);
or U49698 (N_49698,N_49016,N_49487);
and U49699 (N_49699,N_49073,N_49164);
and U49700 (N_49700,N_49486,N_49090);
xnor U49701 (N_49701,N_49332,N_49096);
or U49702 (N_49702,N_49246,N_49198);
nor U49703 (N_49703,N_49138,N_49110);
or U49704 (N_49704,N_49126,N_49367);
and U49705 (N_49705,N_49046,N_49115);
xnor U49706 (N_49706,N_49470,N_49231);
nand U49707 (N_49707,N_49132,N_49250);
and U49708 (N_49708,N_49381,N_49114);
or U49709 (N_49709,N_49434,N_49108);
or U49710 (N_49710,N_49035,N_49451);
and U49711 (N_49711,N_49464,N_49432);
and U49712 (N_49712,N_49305,N_49209);
or U49713 (N_49713,N_49041,N_49288);
nand U49714 (N_49714,N_49244,N_49345);
nand U49715 (N_49715,N_49368,N_49120);
or U49716 (N_49716,N_49135,N_49447);
nor U49717 (N_49717,N_49352,N_49379);
nor U49718 (N_49718,N_49374,N_49193);
xor U49719 (N_49719,N_49321,N_49082);
xor U49720 (N_49720,N_49472,N_49271);
xnor U49721 (N_49721,N_49125,N_49099);
nand U49722 (N_49722,N_49475,N_49181);
xor U49723 (N_49723,N_49448,N_49119);
or U49724 (N_49724,N_49388,N_49440);
xnor U49725 (N_49725,N_49051,N_49386);
and U49726 (N_49726,N_49285,N_49133);
or U49727 (N_49727,N_49172,N_49384);
xor U49728 (N_49728,N_49241,N_49144);
and U49729 (N_49729,N_49025,N_49289);
nor U49730 (N_49730,N_49098,N_49343);
or U49731 (N_49731,N_49227,N_49128);
nand U49732 (N_49732,N_49065,N_49353);
or U49733 (N_49733,N_49054,N_49257);
and U49734 (N_49734,N_49398,N_49187);
nor U49735 (N_49735,N_49141,N_49460);
nand U49736 (N_49736,N_49179,N_49346);
and U49737 (N_49737,N_49391,N_49207);
nand U49738 (N_49738,N_49496,N_49476);
nor U49739 (N_49739,N_49034,N_49032);
nor U49740 (N_49740,N_49199,N_49313);
xor U49741 (N_49741,N_49433,N_49116);
and U49742 (N_49742,N_49439,N_49251);
and U49743 (N_49743,N_49258,N_49124);
or U49744 (N_49744,N_49100,N_49327);
nand U49745 (N_49745,N_49056,N_49488);
nand U49746 (N_49746,N_49233,N_49494);
nand U49747 (N_49747,N_49178,N_49412);
xor U49748 (N_49748,N_49184,N_49237);
xnor U49749 (N_49749,N_49023,N_49408);
and U49750 (N_49750,N_49126,N_49263);
or U49751 (N_49751,N_49440,N_49123);
and U49752 (N_49752,N_49061,N_49233);
xnor U49753 (N_49753,N_49292,N_49187);
or U49754 (N_49754,N_49226,N_49254);
nor U49755 (N_49755,N_49370,N_49279);
xnor U49756 (N_49756,N_49259,N_49054);
and U49757 (N_49757,N_49318,N_49337);
nand U49758 (N_49758,N_49496,N_49480);
and U49759 (N_49759,N_49208,N_49032);
xnor U49760 (N_49760,N_49072,N_49200);
nor U49761 (N_49761,N_49495,N_49239);
nand U49762 (N_49762,N_49272,N_49111);
or U49763 (N_49763,N_49042,N_49232);
nand U49764 (N_49764,N_49408,N_49378);
nor U49765 (N_49765,N_49241,N_49313);
nor U49766 (N_49766,N_49434,N_49286);
and U49767 (N_49767,N_49234,N_49416);
nand U49768 (N_49768,N_49461,N_49202);
nand U49769 (N_49769,N_49160,N_49389);
nor U49770 (N_49770,N_49014,N_49206);
nor U49771 (N_49771,N_49116,N_49328);
xnor U49772 (N_49772,N_49409,N_49432);
and U49773 (N_49773,N_49456,N_49168);
xor U49774 (N_49774,N_49324,N_49151);
nor U49775 (N_49775,N_49426,N_49366);
nor U49776 (N_49776,N_49112,N_49046);
nor U49777 (N_49777,N_49418,N_49324);
nand U49778 (N_49778,N_49415,N_49081);
and U49779 (N_49779,N_49179,N_49078);
or U49780 (N_49780,N_49208,N_49320);
or U49781 (N_49781,N_49402,N_49351);
nand U49782 (N_49782,N_49234,N_49031);
xnor U49783 (N_49783,N_49473,N_49207);
xor U49784 (N_49784,N_49242,N_49348);
or U49785 (N_49785,N_49211,N_49307);
nand U49786 (N_49786,N_49269,N_49479);
and U49787 (N_49787,N_49330,N_49153);
nor U49788 (N_49788,N_49265,N_49267);
xor U49789 (N_49789,N_49475,N_49228);
and U49790 (N_49790,N_49060,N_49408);
and U49791 (N_49791,N_49465,N_49489);
xnor U49792 (N_49792,N_49435,N_49242);
and U49793 (N_49793,N_49222,N_49473);
nor U49794 (N_49794,N_49462,N_49192);
or U49795 (N_49795,N_49361,N_49078);
nand U49796 (N_49796,N_49137,N_49114);
nor U49797 (N_49797,N_49409,N_49385);
nor U49798 (N_49798,N_49129,N_49128);
or U49799 (N_49799,N_49311,N_49029);
and U49800 (N_49800,N_49227,N_49385);
nand U49801 (N_49801,N_49130,N_49419);
xor U49802 (N_49802,N_49369,N_49043);
nand U49803 (N_49803,N_49188,N_49478);
or U49804 (N_49804,N_49207,N_49458);
nor U49805 (N_49805,N_49104,N_49273);
nand U49806 (N_49806,N_49405,N_49421);
or U49807 (N_49807,N_49179,N_49257);
nand U49808 (N_49808,N_49423,N_49371);
nor U49809 (N_49809,N_49394,N_49118);
xnor U49810 (N_49810,N_49207,N_49248);
and U49811 (N_49811,N_49372,N_49316);
nand U49812 (N_49812,N_49340,N_49106);
or U49813 (N_49813,N_49131,N_49037);
nand U49814 (N_49814,N_49138,N_49003);
xor U49815 (N_49815,N_49265,N_49019);
xnor U49816 (N_49816,N_49052,N_49253);
nand U49817 (N_49817,N_49025,N_49332);
nand U49818 (N_49818,N_49358,N_49428);
or U49819 (N_49819,N_49222,N_49031);
and U49820 (N_49820,N_49256,N_49469);
nand U49821 (N_49821,N_49347,N_49017);
xnor U49822 (N_49822,N_49425,N_49047);
nor U49823 (N_49823,N_49182,N_49246);
xor U49824 (N_49824,N_49139,N_49090);
or U49825 (N_49825,N_49257,N_49260);
or U49826 (N_49826,N_49033,N_49007);
nand U49827 (N_49827,N_49227,N_49008);
nand U49828 (N_49828,N_49145,N_49285);
and U49829 (N_49829,N_49267,N_49000);
xnor U49830 (N_49830,N_49108,N_49340);
or U49831 (N_49831,N_49428,N_49213);
xor U49832 (N_49832,N_49429,N_49431);
nand U49833 (N_49833,N_49246,N_49380);
nor U49834 (N_49834,N_49207,N_49227);
nand U49835 (N_49835,N_49028,N_49018);
and U49836 (N_49836,N_49341,N_49419);
xor U49837 (N_49837,N_49446,N_49429);
nor U49838 (N_49838,N_49093,N_49143);
nor U49839 (N_49839,N_49335,N_49017);
nand U49840 (N_49840,N_49435,N_49484);
or U49841 (N_49841,N_49161,N_49266);
or U49842 (N_49842,N_49139,N_49429);
or U49843 (N_49843,N_49097,N_49162);
nor U49844 (N_49844,N_49166,N_49326);
xor U49845 (N_49845,N_49111,N_49378);
nand U49846 (N_49846,N_49003,N_49488);
nor U49847 (N_49847,N_49343,N_49485);
xnor U49848 (N_49848,N_49313,N_49299);
nor U49849 (N_49849,N_49181,N_49078);
and U49850 (N_49850,N_49042,N_49348);
xnor U49851 (N_49851,N_49230,N_49197);
and U49852 (N_49852,N_49245,N_49147);
and U49853 (N_49853,N_49485,N_49243);
and U49854 (N_49854,N_49209,N_49343);
or U49855 (N_49855,N_49113,N_49459);
xnor U49856 (N_49856,N_49264,N_49153);
xnor U49857 (N_49857,N_49360,N_49484);
nand U49858 (N_49858,N_49489,N_49191);
nor U49859 (N_49859,N_49405,N_49357);
nand U49860 (N_49860,N_49350,N_49016);
or U49861 (N_49861,N_49228,N_49075);
nand U49862 (N_49862,N_49389,N_49350);
nand U49863 (N_49863,N_49261,N_49358);
nand U49864 (N_49864,N_49467,N_49222);
nor U49865 (N_49865,N_49271,N_49350);
and U49866 (N_49866,N_49480,N_49016);
nor U49867 (N_49867,N_49072,N_49471);
nand U49868 (N_49868,N_49190,N_49290);
and U49869 (N_49869,N_49466,N_49452);
xor U49870 (N_49870,N_49231,N_49236);
xor U49871 (N_49871,N_49032,N_49073);
xor U49872 (N_49872,N_49272,N_49059);
and U49873 (N_49873,N_49429,N_49399);
nand U49874 (N_49874,N_49480,N_49435);
nor U49875 (N_49875,N_49001,N_49129);
nor U49876 (N_49876,N_49174,N_49263);
or U49877 (N_49877,N_49097,N_49489);
or U49878 (N_49878,N_49177,N_49219);
xor U49879 (N_49879,N_49053,N_49269);
nor U49880 (N_49880,N_49261,N_49440);
xnor U49881 (N_49881,N_49371,N_49427);
or U49882 (N_49882,N_49141,N_49122);
and U49883 (N_49883,N_49348,N_49361);
nor U49884 (N_49884,N_49358,N_49278);
nor U49885 (N_49885,N_49218,N_49125);
and U49886 (N_49886,N_49495,N_49245);
nand U49887 (N_49887,N_49312,N_49164);
xnor U49888 (N_49888,N_49180,N_49290);
xor U49889 (N_49889,N_49430,N_49190);
nor U49890 (N_49890,N_49179,N_49453);
and U49891 (N_49891,N_49361,N_49282);
xnor U49892 (N_49892,N_49338,N_49254);
nand U49893 (N_49893,N_49252,N_49021);
nor U49894 (N_49894,N_49025,N_49123);
and U49895 (N_49895,N_49012,N_49138);
nor U49896 (N_49896,N_49397,N_49250);
nor U49897 (N_49897,N_49057,N_49083);
nand U49898 (N_49898,N_49184,N_49361);
xor U49899 (N_49899,N_49106,N_49355);
xnor U49900 (N_49900,N_49241,N_49173);
and U49901 (N_49901,N_49228,N_49008);
nor U49902 (N_49902,N_49389,N_49001);
or U49903 (N_49903,N_49292,N_49430);
and U49904 (N_49904,N_49143,N_49239);
xor U49905 (N_49905,N_49086,N_49302);
or U49906 (N_49906,N_49498,N_49294);
or U49907 (N_49907,N_49355,N_49214);
nor U49908 (N_49908,N_49083,N_49425);
nor U49909 (N_49909,N_49453,N_49170);
xor U49910 (N_49910,N_49126,N_49143);
nand U49911 (N_49911,N_49309,N_49442);
and U49912 (N_49912,N_49196,N_49381);
nor U49913 (N_49913,N_49219,N_49113);
nand U49914 (N_49914,N_49257,N_49070);
and U49915 (N_49915,N_49279,N_49008);
xnor U49916 (N_49916,N_49235,N_49400);
xnor U49917 (N_49917,N_49048,N_49414);
or U49918 (N_49918,N_49419,N_49270);
or U49919 (N_49919,N_49031,N_49409);
or U49920 (N_49920,N_49212,N_49394);
or U49921 (N_49921,N_49457,N_49279);
xnor U49922 (N_49922,N_49231,N_49183);
xnor U49923 (N_49923,N_49206,N_49438);
nor U49924 (N_49924,N_49058,N_49339);
nand U49925 (N_49925,N_49104,N_49319);
nand U49926 (N_49926,N_49325,N_49349);
or U49927 (N_49927,N_49206,N_49004);
or U49928 (N_49928,N_49026,N_49005);
and U49929 (N_49929,N_49347,N_49225);
or U49930 (N_49930,N_49271,N_49078);
and U49931 (N_49931,N_49424,N_49351);
nor U49932 (N_49932,N_49405,N_49218);
nand U49933 (N_49933,N_49404,N_49066);
xor U49934 (N_49934,N_49189,N_49455);
nand U49935 (N_49935,N_49059,N_49214);
or U49936 (N_49936,N_49012,N_49136);
nand U49937 (N_49937,N_49261,N_49077);
and U49938 (N_49938,N_49070,N_49068);
or U49939 (N_49939,N_49263,N_49272);
and U49940 (N_49940,N_49092,N_49149);
xnor U49941 (N_49941,N_49448,N_49253);
and U49942 (N_49942,N_49471,N_49153);
and U49943 (N_49943,N_49376,N_49499);
nand U49944 (N_49944,N_49237,N_49338);
xor U49945 (N_49945,N_49481,N_49411);
nor U49946 (N_49946,N_49355,N_49140);
or U49947 (N_49947,N_49263,N_49176);
xnor U49948 (N_49948,N_49194,N_49199);
and U49949 (N_49949,N_49362,N_49041);
and U49950 (N_49950,N_49110,N_49486);
nand U49951 (N_49951,N_49350,N_49272);
nor U49952 (N_49952,N_49122,N_49242);
xnor U49953 (N_49953,N_49203,N_49326);
or U49954 (N_49954,N_49443,N_49001);
xor U49955 (N_49955,N_49132,N_49046);
xnor U49956 (N_49956,N_49349,N_49282);
and U49957 (N_49957,N_49285,N_49380);
or U49958 (N_49958,N_49480,N_49443);
nand U49959 (N_49959,N_49343,N_49225);
nand U49960 (N_49960,N_49481,N_49018);
and U49961 (N_49961,N_49073,N_49247);
nor U49962 (N_49962,N_49005,N_49182);
nand U49963 (N_49963,N_49055,N_49189);
nand U49964 (N_49964,N_49112,N_49173);
nand U49965 (N_49965,N_49305,N_49013);
or U49966 (N_49966,N_49258,N_49111);
xnor U49967 (N_49967,N_49403,N_49434);
or U49968 (N_49968,N_49370,N_49203);
or U49969 (N_49969,N_49236,N_49489);
nand U49970 (N_49970,N_49155,N_49186);
xnor U49971 (N_49971,N_49091,N_49359);
and U49972 (N_49972,N_49452,N_49391);
nand U49973 (N_49973,N_49182,N_49290);
nand U49974 (N_49974,N_49170,N_49236);
xnor U49975 (N_49975,N_49095,N_49333);
nand U49976 (N_49976,N_49407,N_49334);
xnor U49977 (N_49977,N_49307,N_49325);
or U49978 (N_49978,N_49185,N_49449);
and U49979 (N_49979,N_49101,N_49413);
nor U49980 (N_49980,N_49244,N_49214);
xor U49981 (N_49981,N_49453,N_49381);
nand U49982 (N_49982,N_49344,N_49374);
xnor U49983 (N_49983,N_49186,N_49084);
and U49984 (N_49984,N_49236,N_49130);
xnor U49985 (N_49985,N_49320,N_49165);
xnor U49986 (N_49986,N_49445,N_49103);
and U49987 (N_49987,N_49085,N_49111);
nand U49988 (N_49988,N_49157,N_49455);
xor U49989 (N_49989,N_49200,N_49025);
or U49990 (N_49990,N_49378,N_49416);
or U49991 (N_49991,N_49032,N_49419);
xnor U49992 (N_49992,N_49359,N_49489);
nand U49993 (N_49993,N_49245,N_49134);
nor U49994 (N_49994,N_49379,N_49205);
or U49995 (N_49995,N_49179,N_49014);
and U49996 (N_49996,N_49085,N_49158);
nor U49997 (N_49997,N_49349,N_49217);
nand U49998 (N_49998,N_49130,N_49193);
or U49999 (N_49999,N_49412,N_49225);
xor UO_0 (O_0,N_49958,N_49899);
xor UO_1 (O_1,N_49860,N_49625);
xnor UO_2 (O_2,N_49685,N_49840);
nand UO_3 (O_3,N_49930,N_49824);
or UO_4 (O_4,N_49921,N_49852);
or UO_5 (O_5,N_49572,N_49853);
nand UO_6 (O_6,N_49874,N_49695);
nand UO_7 (O_7,N_49769,N_49708);
or UO_8 (O_8,N_49931,N_49894);
or UO_9 (O_9,N_49993,N_49841);
nand UO_10 (O_10,N_49754,N_49650);
nor UO_11 (O_11,N_49526,N_49870);
nand UO_12 (O_12,N_49546,N_49888);
and UO_13 (O_13,N_49823,N_49801);
nor UO_14 (O_14,N_49503,N_49987);
nand UO_15 (O_15,N_49822,N_49770);
and UO_16 (O_16,N_49764,N_49953);
nor UO_17 (O_17,N_49863,N_49879);
nor UO_18 (O_18,N_49937,N_49532);
nor UO_19 (O_19,N_49776,N_49590);
xor UO_20 (O_20,N_49976,N_49678);
xor UO_21 (O_21,N_49654,N_49765);
and UO_22 (O_22,N_49825,N_49715);
xnor UO_23 (O_23,N_49703,N_49665);
nand UO_24 (O_24,N_49965,N_49522);
and UO_25 (O_25,N_49548,N_49595);
nor UO_26 (O_26,N_49712,N_49839);
or UO_27 (O_27,N_49615,N_49726);
and UO_28 (O_28,N_49621,N_49566);
nand UO_29 (O_29,N_49861,N_49677);
xnor UO_30 (O_30,N_49926,N_49794);
nor UO_31 (O_31,N_49913,N_49842);
nor UO_32 (O_32,N_49938,N_49549);
nand UO_33 (O_33,N_49602,N_49688);
xnor UO_34 (O_34,N_49727,N_49858);
nand UO_35 (O_35,N_49772,N_49810);
or UO_36 (O_36,N_49831,N_49989);
xor UO_37 (O_37,N_49828,N_49607);
xnor UO_38 (O_38,N_49576,N_49799);
nor UO_39 (O_39,N_49835,N_49785);
nand UO_40 (O_40,N_49543,N_49783);
nor UO_41 (O_41,N_49714,N_49960);
xor UO_42 (O_42,N_49529,N_49959);
and UO_43 (O_43,N_49671,N_49922);
nand UO_44 (O_44,N_49504,N_49721);
nor UO_45 (O_45,N_49649,N_49713);
and UO_46 (O_46,N_49652,N_49838);
nand UO_47 (O_47,N_49539,N_49758);
nand UO_48 (O_48,N_49686,N_49571);
and UO_49 (O_49,N_49626,N_49743);
and UO_50 (O_50,N_49533,N_49547);
nor UO_51 (O_51,N_49982,N_49568);
xor UO_52 (O_52,N_49779,N_49979);
xnor UO_53 (O_53,N_49747,N_49717);
and UO_54 (O_54,N_49847,N_49844);
nor UO_55 (O_55,N_49573,N_49709);
nand UO_56 (O_56,N_49676,N_49943);
nor UO_57 (O_57,N_49633,N_49911);
xnor UO_58 (O_58,N_49800,N_49986);
or UO_59 (O_59,N_49682,N_49978);
and UO_60 (O_60,N_49508,N_49559);
nor UO_61 (O_61,N_49704,N_49638);
nand UO_62 (O_62,N_49803,N_49701);
or UO_63 (O_63,N_49591,N_49971);
and UO_64 (O_64,N_49977,N_49789);
nand UO_65 (O_65,N_49804,N_49541);
nor UO_66 (O_66,N_49718,N_49927);
and UO_67 (O_67,N_49890,N_49683);
nand UO_68 (O_68,N_49616,N_49812);
xor UO_69 (O_69,N_49700,N_49855);
xor UO_70 (O_70,N_49939,N_49788);
and UO_71 (O_71,N_49759,N_49581);
or UO_72 (O_72,N_49784,N_49643);
nand UO_73 (O_73,N_49620,N_49837);
and UO_74 (O_74,N_49903,N_49735);
and UO_75 (O_75,N_49862,N_49906);
or UO_76 (O_76,N_49728,N_49535);
nor UO_77 (O_77,N_49944,N_49796);
xnor UO_78 (O_78,N_49955,N_49946);
and UO_79 (O_79,N_49511,N_49883);
and UO_80 (O_80,N_49694,N_49962);
nand UO_81 (O_81,N_49974,N_49645);
xnor UO_82 (O_82,N_49745,N_49928);
nand UO_83 (O_83,N_49947,N_49768);
or UO_84 (O_84,N_49790,N_49640);
nor UO_85 (O_85,N_49540,N_49952);
nand UO_86 (O_86,N_49603,N_49707);
or UO_87 (O_87,N_49691,N_49739);
and UO_88 (O_88,N_49793,N_49725);
nor UO_89 (O_89,N_49820,N_49570);
xor UO_90 (O_90,N_49669,N_49629);
or UO_91 (O_91,N_49580,N_49599);
xnor UO_92 (O_92,N_49527,N_49752);
nand UO_93 (O_93,N_49916,N_49613);
xnor UO_94 (O_94,N_49990,N_49923);
xnor UO_95 (O_95,N_49867,N_49587);
or UO_96 (O_96,N_49802,N_49856);
nand UO_97 (O_97,N_49775,N_49663);
or UO_98 (O_98,N_49639,N_49687);
and UO_99 (O_99,N_49562,N_49817);
nand UO_100 (O_100,N_49675,N_49872);
nor UO_101 (O_101,N_49729,N_49614);
and UO_102 (O_102,N_49693,N_49997);
and UO_103 (O_103,N_49732,N_49884);
nor UO_104 (O_104,N_49617,N_49632);
xor UO_105 (O_105,N_49918,N_49821);
nor UO_106 (O_106,N_49807,N_49791);
nand UO_107 (O_107,N_49980,N_49935);
and UO_108 (O_108,N_49763,N_49720);
xor UO_109 (O_109,N_49521,N_49734);
and UO_110 (O_110,N_49628,N_49753);
xor UO_111 (O_111,N_49505,N_49967);
or UO_112 (O_112,N_49648,N_49904);
nand UO_113 (O_113,N_49778,N_49597);
nand UO_114 (O_114,N_49780,N_49667);
and UO_115 (O_115,N_49895,N_49956);
xnor UO_116 (O_116,N_49742,N_49545);
xor UO_117 (O_117,N_49689,N_49538);
nand UO_118 (O_118,N_49898,N_49975);
or UO_119 (O_119,N_49588,N_49644);
nand UO_120 (O_120,N_49600,N_49887);
nor UO_121 (O_121,N_49605,N_49530);
and UO_122 (O_122,N_49968,N_49954);
and UO_123 (O_123,N_49555,N_49854);
and UO_124 (O_124,N_49710,N_49698);
xor UO_125 (O_125,N_49659,N_49813);
nor UO_126 (O_126,N_49762,N_49751);
xnor UO_127 (O_127,N_49963,N_49738);
and UO_128 (O_128,N_49557,N_49582);
and UO_129 (O_129,N_49900,N_49934);
xor UO_130 (O_130,N_49501,N_49544);
xnor UO_131 (O_131,N_49950,N_49907);
xnor UO_132 (O_132,N_49716,N_49896);
or UO_133 (O_133,N_49814,N_49586);
xnor UO_134 (O_134,N_49619,N_49750);
xnor UO_135 (O_135,N_49513,N_49848);
xor UO_136 (O_136,N_49843,N_49552);
xor UO_137 (O_137,N_49551,N_49542);
nor UO_138 (O_138,N_49520,N_49664);
nor UO_139 (O_139,N_49809,N_49696);
and UO_140 (O_140,N_49563,N_49740);
nor UO_141 (O_141,N_49951,N_49897);
and UO_142 (O_142,N_49681,N_49636);
xnor UO_143 (O_143,N_49601,N_49849);
xor UO_144 (O_144,N_49658,N_49558);
or UO_145 (O_145,N_49635,N_49737);
nor UO_146 (O_146,N_49606,N_49631);
or UO_147 (O_147,N_49512,N_49630);
nor UO_148 (O_148,N_49827,N_49949);
nand UO_149 (O_149,N_49502,N_49866);
nand UO_150 (O_150,N_49875,N_49692);
and UO_151 (O_151,N_49583,N_49819);
or UO_152 (O_152,N_49942,N_49711);
nand UO_153 (O_153,N_49992,N_49749);
and UO_154 (O_154,N_49973,N_49961);
xor UO_155 (O_155,N_49553,N_49579);
nor UO_156 (O_156,N_49519,N_49797);
nand UO_157 (O_157,N_49966,N_49920);
nand UO_158 (O_158,N_49661,N_49932);
xor UO_159 (O_159,N_49670,N_49656);
nor UO_160 (O_160,N_49845,N_49892);
xor UO_161 (O_161,N_49537,N_49748);
and UO_162 (O_162,N_49550,N_49724);
nand UO_163 (O_163,N_49510,N_49651);
xor UO_164 (O_164,N_49984,N_49612);
or UO_165 (O_165,N_49868,N_49878);
and UO_166 (O_166,N_49585,N_49876);
and UO_167 (O_167,N_49627,N_49924);
and UO_168 (O_168,N_49516,N_49915);
and UO_169 (O_169,N_49972,N_49910);
nor UO_170 (O_170,N_49531,N_49657);
nor UO_171 (O_171,N_49554,N_49941);
and UO_172 (O_172,N_49988,N_49592);
nand UO_173 (O_173,N_49981,N_49705);
xnor UO_174 (O_174,N_49830,N_49850);
and UO_175 (O_175,N_49746,N_49826);
or UO_176 (O_176,N_49761,N_49885);
nand UO_177 (O_177,N_49564,N_49859);
and UO_178 (O_178,N_49919,N_49518);
and UO_179 (O_179,N_49808,N_49970);
nor UO_180 (O_180,N_49755,N_49873);
and UO_181 (O_181,N_49893,N_49925);
or UO_182 (O_182,N_49706,N_49757);
nor UO_183 (O_183,N_49642,N_49575);
nand UO_184 (O_184,N_49598,N_49741);
nand UO_185 (O_185,N_49864,N_49829);
nand UO_186 (O_186,N_49699,N_49994);
or UO_187 (O_187,N_49936,N_49806);
nand UO_188 (O_188,N_49731,N_49787);
or UO_189 (O_189,N_49507,N_49851);
nand UO_190 (O_190,N_49760,N_49945);
nor UO_191 (O_191,N_49836,N_49567);
xor UO_192 (O_192,N_49891,N_49506);
nand UO_193 (O_193,N_49834,N_49795);
nand UO_194 (O_194,N_49996,N_49865);
nand UO_195 (O_195,N_49589,N_49983);
or UO_196 (O_196,N_49905,N_49815);
or UO_197 (O_197,N_49917,N_49957);
nand UO_198 (O_198,N_49697,N_49869);
xnor UO_199 (O_199,N_49912,N_49569);
and UO_200 (O_200,N_49624,N_49881);
or UO_201 (O_201,N_49781,N_49882);
nor UO_202 (O_202,N_49514,N_49515);
nand UO_203 (O_203,N_49623,N_49914);
nand UO_204 (O_204,N_49618,N_49766);
nor UO_205 (O_205,N_49933,N_49889);
nand UO_206 (O_206,N_49886,N_49901);
xnor UO_207 (O_207,N_49684,N_49798);
xor UO_208 (O_208,N_49647,N_49608);
xnor UO_209 (O_209,N_49909,N_49880);
or UO_210 (O_210,N_49560,N_49611);
xor UO_211 (O_211,N_49517,N_49871);
xor UO_212 (O_212,N_49622,N_49736);
or UO_213 (O_213,N_49782,N_49964);
xnor UO_214 (O_214,N_49672,N_49637);
or UO_215 (O_215,N_49846,N_49674);
and UO_216 (O_216,N_49995,N_49767);
xnor UO_217 (O_217,N_49730,N_49771);
and UO_218 (O_218,N_49940,N_49577);
and UO_219 (O_219,N_49733,N_49660);
xnor UO_220 (O_220,N_49833,N_49998);
or UO_221 (O_221,N_49723,N_49500);
and UO_222 (O_222,N_49610,N_49774);
nor UO_223 (O_223,N_49985,N_49509);
xor UO_224 (O_224,N_49662,N_49534);
and UO_225 (O_225,N_49594,N_49634);
nand UO_226 (O_226,N_49578,N_49584);
and UO_227 (O_227,N_49609,N_49786);
nor UO_228 (O_228,N_49641,N_49604);
or UO_229 (O_229,N_49561,N_49679);
and UO_230 (O_230,N_49857,N_49969);
xnor UO_231 (O_231,N_49818,N_49646);
nand UO_232 (O_232,N_49702,N_49574);
or UO_233 (O_233,N_49756,N_49948);
xnor UO_234 (O_234,N_49680,N_49690);
nand UO_235 (O_235,N_49777,N_49525);
and UO_236 (O_236,N_49668,N_49593);
and UO_237 (O_237,N_49929,N_49565);
xnor UO_238 (O_238,N_49523,N_49773);
and UO_239 (O_239,N_49596,N_49811);
or UO_240 (O_240,N_49832,N_49719);
nor UO_241 (O_241,N_49999,N_49902);
or UO_242 (O_242,N_49536,N_49666);
or UO_243 (O_243,N_49673,N_49524);
and UO_244 (O_244,N_49744,N_49528);
and UO_245 (O_245,N_49816,N_49792);
nand UO_246 (O_246,N_49805,N_49653);
nand UO_247 (O_247,N_49877,N_49722);
or UO_248 (O_248,N_49655,N_49556);
nor UO_249 (O_249,N_49991,N_49908);
nand UO_250 (O_250,N_49783,N_49866);
xnor UO_251 (O_251,N_49823,N_49923);
nor UO_252 (O_252,N_49713,N_49916);
and UO_253 (O_253,N_49602,N_49643);
or UO_254 (O_254,N_49765,N_49773);
xor UO_255 (O_255,N_49903,N_49599);
xnor UO_256 (O_256,N_49908,N_49735);
and UO_257 (O_257,N_49820,N_49569);
or UO_258 (O_258,N_49702,N_49818);
nand UO_259 (O_259,N_49745,N_49648);
nor UO_260 (O_260,N_49645,N_49649);
nand UO_261 (O_261,N_49681,N_49999);
or UO_262 (O_262,N_49883,N_49574);
and UO_263 (O_263,N_49504,N_49853);
and UO_264 (O_264,N_49808,N_49929);
nand UO_265 (O_265,N_49965,N_49774);
and UO_266 (O_266,N_49995,N_49723);
nand UO_267 (O_267,N_49932,N_49968);
or UO_268 (O_268,N_49679,N_49597);
nor UO_269 (O_269,N_49876,N_49847);
or UO_270 (O_270,N_49664,N_49668);
and UO_271 (O_271,N_49993,N_49676);
xnor UO_272 (O_272,N_49731,N_49583);
xnor UO_273 (O_273,N_49863,N_49571);
and UO_274 (O_274,N_49845,N_49673);
nand UO_275 (O_275,N_49920,N_49593);
nor UO_276 (O_276,N_49613,N_49655);
nand UO_277 (O_277,N_49937,N_49517);
nand UO_278 (O_278,N_49938,N_49966);
or UO_279 (O_279,N_49674,N_49983);
nand UO_280 (O_280,N_49859,N_49842);
nand UO_281 (O_281,N_49969,N_49562);
nand UO_282 (O_282,N_49897,N_49781);
or UO_283 (O_283,N_49519,N_49768);
xnor UO_284 (O_284,N_49903,N_49909);
xor UO_285 (O_285,N_49534,N_49879);
or UO_286 (O_286,N_49672,N_49533);
nand UO_287 (O_287,N_49503,N_49676);
or UO_288 (O_288,N_49741,N_49694);
nor UO_289 (O_289,N_49944,N_49943);
and UO_290 (O_290,N_49545,N_49989);
or UO_291 (O_291,N_49527,N_49920);
nor UO_292 (O_292,N_49804,N_49924);
or UO_293 (O_293,N_49998,N_49627);
or UO_294 (O_294,N_49697,N_49765);
xor UO_295 (O_295,N_49672,N_49570);
nand UO_296 (O_296,N_49614,N_49786);
and UO_297 (O_297,N_49700,N_49887);
and UO_298 (O_298,N_49736,N_49647);
nor UO_299 (O_299,N_49996,N_49905);
nor UO_300 (O_300,N_49685,N_49642);
or UO_301 (O_301,N_49551,N_49666);
nand UO_302 (O_302,N_49726,N_49829);
and UO_303 (O_303,N_49739,N_49975);
nor UO_304 (O_304,N_49641,N_49602);
xnor UO_305 (O_305,N_49583,N_49853);
xnor UO_306 (O_306,N_49845,N_49831);
xnor UO_307 (O_307,N_49799,N_49840);
xor UO_308 (O_308,N_49798,N_49903);
nor UO_309 (O_309,N_49707,N_49845);
xnor UO_310 (O_310,N_49531,N_49665);
and UO_311 (O_311,N_49949,N_49761);
and UO_312 (O_312,N_49890,N_49550);
xnor UO_313 (O_313,N_49614,N_49556);
xor UO_314 (O_314,N_49898,N_49758);
and UO_315 (O_315,N_49966,N_49693);
nand UO_316 (O_316,N_49692,N_49972);
or UO_317 (O_317,N_49841,N_49807);
nor UO_318 (O_318,N_49842,N_49633);
and UO_319 (O_319,N_49507,N_49676);
nand UO_320 (O_320,N_49764,N_49820);
nor UO_321 (O_321,N_49718,N_49573);
or UO_322 (O_322,N_49886,N_49971);
xor UO_323 (O_323,N_49614,N_49508);
or UO_324 (O_324,N_49579,N_49952);
and UO_325 (O_325,N_49671,N_49515);
xor UO_326 (O_326,N_49808,N_49767);
or UO_327 (O_327,N_49615,N_49597);
and UO_328 (O_328,N_49758,N_49954);
nand UO_329 (O_329,N_49754,N_49792);
and UO_330 (O_330,N_49620,N_49902);
and UO_331 (O_331,N_49809,N_49755);
and UO_332 (O_332,N_49753,N_49631);
nand UO_333 (O_333,N_49964,N_49607);
xnor UO_334 (O_334,N_49927,N_49609);
and UO_335 (O_335,N_49766,N_49843);
xor UO_336 (O_336,N_49859,N_49753);
and UO_337 (O_337,N_49742,N_49537);
nand UO_338 (O_338,N_49931,N_49594);
xor UO_339 (O_339,N_49647,N_49826);
xor UO_340 (O_340,N_49851,N_49779);
xor UO_341 (O_341,N_49752,N_49589);
and UO_342 (O_342,N_49893,N_49617);
xor UO_343 (O_343,N_49648,N_49948);
or UO_344 (O_344,N_49543,N_49691);
nor UO_345 (O_345,N_49557,N_49985);
xor UO_346 (O_346,N_49704,N_49937);
nand UO_347 (O_347,N_49683,N_49914);
nand UO_348 (O_348,N_49812,N_49865);
and UO_349 (O_349,N_49515,N_49846);
xor UO_350 (O_350,N_49756,N_49760);
and UO_351 (O_351,N_49756,N_49971);
xor UO_352 (O_352,N_49684,N_49924);
nor UO_353 (O_353,N_49800,N_49619);
nor UO_354 (O_354,N_49845,N_49959);
nor UO_355 (O_355,N_49596,N_49595);
nand UO_356 (O_356,N_49917,N_49620);
and UO_357 (O_357,N_49772,N_49942);
or UO_358 (O_358,N_49667,N_49966);
or UO_359 (O_359,N_49942,N_49751);
nand UO_360 (O_360,N_49856,N_49561);
and UO_361 (O_361,N_49565,N_49833);
or UO_362 (O_362,N_49766,N_49801);
xnor UO_363 (O_363,N_49876,N_49849);
or UO_364 (O_364,N_49624,N_49638);
nor UO_365 (O_365,N_49757,N_49623);
or UO_366 (O_366,N_49911,N_49739);
and UO_367 (O_367,N_49745,N_49679);
nor UO_368 (O_368,N_49672,N_49546);
nor UO_369 (O_369,N_49510,N_49841);
or UO_370 (O_370,N_49559,N_49584);
xor UO_371 (O_371,N_49509,N_49669);
and UO_372 (O_372,N_49621,N_49576);
and UO_373 (O_373,N_49621,N_49661);
nand UO_374 (O_374,N_49674,N_49813);
and UO_375 (O_375,N_49600,N_49994);
nand UO_376 (O_376,N_49930,N_49536);
nor UO_377 (O_377,N_49653,N_49560);
nor UO_378 (O_378,N_49789,N_49817);
nor UO_379 (O_379,N_49632,N_49757);
or UO_380 (O_380,N_49679,N_49885);
nand UO_381 (O_381,N_49840,N_49982);
nand UO_382 (O_382,N_49694,N_49893);
nor UO_383 (O_383,N_49679,N_49550);
nor UO_384 (O_384,N_49513,N_49728);
nand UO_385 (O_385,N_49523,N_49951);
xnor UO_386 (O_386,N_49523,N_49601);
nand UO_387 (O_387,N_49897,N_49997);
nor UO_388 (O_388,N_49971,N_49539);
or UO_389 (O_389,N_49701,N_49878);
or UO_390 (O_390,N_49930,N_49533);
nand UO_391 (O_391,N_49658,N_49975);
xor UO_392 (O_392,N_49856,N_49880);
nor UO_393 (O_393,N_49573,N_49860);
nand UO_394 (O_394,N_49840,N_49917);
nor UO_395 (O_395,N_49926,N_49688);
xnor UO_396 (O_396,N_49961,N_49965);
or UO_397 (O_397,N_49802,N_49936);
and UO_398 (O_398,N_49552,N_49736);
and UO_399 (O_399,N_49542,N_49831);
nand UO_400 (O_400,N_49850,N_49597);
xor UO_401 (O_401,N_49802,N_49946);
nor UO_402 (O_402,N_49677,N_49916);
and UO_403 (O_403,N_49906,N_49517);
and UO_404 (O_404,N_49540,N_49796);
and UO_405 (O_405,N_49819,N_49518);
nand UO_406 (O_406,N_49961,N_49554);
nand UO_407 (O_407,N_49844,N_49679);
and UO_408 (O_408,N_49640,N_49842);
nand UO_409 (O_409,N_49736,N_49967);
and UO_410 (O_410,N_49855,N_49828);
nor UO_411 (O_411,N_49962,N_49849);
nor UO_412 (O_412,N_49532,N_49827);
nor UO_413 (O_413,N_49758,N_49555);
nand UO_414 (O_414,N_49811,N_49635);
nand UO_415 (O_415,N_49735,N_49663);
xor UO_416 (O_416,N_49981,N_49758);
or UO_417 (O_417,N_49802,N_49731);
nor UO_418 (O_418,N_49759,N_49974);
or UO_419 (O_419,N_49685,N_49851);
nand UO_420 (O_420,N_49711,N_49648);
xnor UO_421 (O_421,N_49507,N_49862);
nand UO_422 (O_422,N_49641,N_49980);
nand UO_423 (O_423,N_49651,N_49547);
nand UO_424 (O_424,N_49995,N_49966);
xnor UO_425 (O_425,N_49977,N_49581);
xor UO_426 (O_426,N_49724,N_49585);
nor UO_427 (O_427,N_49909,N_49865);
or UO_428 (O_428,N_49949,N_49854);
nand UO_429 (O_429,N_49705,N_49818);
and UO_430 (O_430,N_49777,N_49552);
and UO_431 (O_431,N_49861,N_49650);
nand UO_432 (O_432,N_49672,N_49972);
and UO_433 (O_433,N_49785,N_49983);
xnor UO_434 (O_434,N_49513,N_49745);
xor UO_435 (O_435,N_49688,N_49700);
nor UO_436 (O_436,N_49928,N_49654);
or UO_437 (O_437,N_49703,N_49533);
xnor UO_438 (O_438,N_49532,N_49753);
and UO_439 (O_439,N_49584,N_49921);
nor UO_440 (O_440,N_49533,N_49845);
and UO_441 (O_441,N_49653,N_49934);
xnor UO_442 (O_442,N_49981,N_49847);
xnor UO_443 (O_443,N_49522,N_49822);
nor UO_444 (O_444,N_49523,N_49851);
or UO_445 (O_445,N_49694,N_49940);
and UO_446 (O_446,N_49707,N_49706);
and UO_447 (O_447,N_49638,N_49858);
xnor UO_448 (O_448,N_49918,N_49901);
and UO_449 (O_449,N_49773,N_49810);
and UO_450 (O_450,N_49604,N_49617);
nand UO_451 (O_451,N_49690,N_49529);
nor UO_452 (O_452,N_49624,N_49876);
xnor UO_453 (O_453,N_49968,N_49793);
nand UO_454 (O_454,N_49503,N_49875);
and UO_455 (O_455,N_49879,N_49661);
nor UO_456 (O_456,N_49541,N_49893);
nand UO_457 (O_457,N_49637,N_49871);
xor UO_458 (O_458,N_49919,N_49587);
and UO_459 (O_459,N_49756,N_49802);
nor UO_460 (O_460,N_49999,N_49868);
and UO_461 (O_461,N_49930,N_49781);
nor UO_462 (O_462,N_49890,N_49873);
and UO_463 (O_463,N_49988,N_49724);
nand UO_464 (O_464,N_49513,N_49674);
nand UO_465 (O_465,N_49795,N_49791);
nand UO_466 (O_466,N_49764,N_49745);
or UO_467 (O_467,N_49929,N_49665);
and UO_468 (O_468,N_49553,N_49795);
xor UO_469 (O_469,N_49702,N_49708);
nor UO_470 (O_470,N_49564,N_49818);
nor UO_471 (O_471,N_49779,N_49721);
or UO_472 (O_472,N_49993,N_49669);
nor UO_473 (O_473,N_49812,N_49562);
xor UO_474 (O_474,N_49883,N_49704);
nand UO_475 (O_475,N_49764,N_49574);
nor UO_476 (O_476,N_49584,N_49774);
nand UO_477 (O_477,N_49523,N_49689);
nor UO_478 (O_478,N_49566,N_49580);
nor UO_479 (O_479,N_49842,N_49507);
or UO_480 (O_480,N_49836,N_49893);
or UO_481 (O_481,N_49617,N_49620);
and UO_482 (O_482,N_49739,N_49827);
xnor UO_483 (O_483,N_49622,N_49958);
nand UO_484 (O_484,N_49835,N_49602);
and UO_485 (O_485,N_49722,N_49804);
nand UO_486 (O_486,N_49939,N_49655);
and UO_487 (O_487,N_49661,N_49542);
and UO_488 (O_488,N_49636,N_49847);
nor UO_489 (O_489,N_49653,N_49717);
nor UO_490 (O_490,N_49931,N_49628);
and UO_491 (O_491,N_49643,N_49612);
nand UO_492 (O_492,N_49970,N_49925);
and UO_493 (O_493,N_49651,N_49632);
or UO_494 (O_494,N_49911,N_49773);
xnor UO_495 (O_495,N_49852,N_49570);
nor UO_496 (O_496,N_49694,N_49927);
or UO_497 (O_497,N_49711,N_49632);
or UO_498 (O_498,N_49513,N_49819);
and UO_499 (O_499,N_49900,N_49571);
or UO_500 (O_500,N_49626,N_49917);
xor UO_501 (O_501,N_49672,N_49635);
nand UO_502 (O_502,N_49519,N_49592);
nand UO_503 (O_503,N_49512,N_49879);
nor UO_504 (O_504,N_49694,N_49910);
or UO_505 (O_505,N_49966,N_49890);
or UO_506 (O_506,N_49861,N_49708);
nand UO_507 (O_507,N_49656,N_49625);
xor UO_508 (O_508,N_49704,N_49538);
xor UO_509 (O_509,N_49770,N_49581);
nand UO_510 (O_510,N_49613,N_49836);
nand UO_511 (O_511,N_49544,N_49736);
and UO_512 (O_512,N_49777,N_49991);
nand UO_513 (O_513,N_49728,N_49905);
or UO_514 (O_514,N_49568,N_49661);
or UO_515 (O_515,N_49515,N_49609);
nor UO_516 (O_516,N_49516,N_49700);
nor UO_517 (O_517,N_49730,N_49686);
nor UO_518 (O_518,N_49890,N_49778);
nor UO_519 (O_519,N_49677,N_49838);
nand UO_520 (O_520,N_49575,N_49834);
or UO_521 (O_521,N_49674,N_49609);
nor UO_522 (O_522,N_49922,N_49807);
or UO_523 (O_523,N_49947,N_49807);
nor UO_524 (O_524,N_49863,N_49832);
nor UO_525 (O_525,N_49513,N_49708);
nor UO_526 (O_526,N_49793,N_49728);
and UO_527 (O_527,N_49577,N_49992);
nor UO_528 (O_528,N_49759,N_49574);
or UO_529 (O_529,N_49830,N_49562);
and UO_530 (O_530,N_49785,N_49980);
and UO_531 (O_531,N_49695,N_49508);
and UO_532 (O_532,N_49845,N_49550);
or UO_533 (O_533,N_49646,N_49859);
xnor UO_534 (O_534,N_49680,N_49709);
and UO_535 (O_535,N_49568,N_49518);
and UO_536 (O_536,N_49741,N_49910);
and UO_537 (O_537,N_49661,N_49554);
or UO_538 (O_538,N_49595,N_49720);
and UO_539 (O_539,N_49895,N_49518);
or UO_540 (O_540,N_49778,N_49807);
and UO_541 (O_541,N_49833,N_49959);
and UO_542 (O_542,N_49672,N_49879);
xor UO_543 (O_543,N_49934,N_49759);
and UO_544 (O_544,N_49949,N_49880);
nand UO_545 (O_545,N_49687,N_49523);
nand UO_546 (O_546,N_49753,N_49960);
nand UO_547 (O_547,N_49893,N_49832);
or UO_548 (O_548,N_49777,N_49883);
and UO_549 (O_549,N_49622,N_49850);
nor UO_550 (O_550,N_49955,N_49711);
nor UO_551 (O_551,N_49558,N_49868);
or UO_552 (O_552,N_49582,N_49923);
nand UO_553 (O_553,N_49954,N_49915);
nand UO_554 (O_554,N_49650,N_49823);
xor UO_555 (O_555,N_49547,N_49765);
and UO_556 (O_556,N_49925,N_49982);
or UO_557 (O_557,N_49990,N_49735);
and UO_558 (O_558,N_49902,N_49534);
and UO_559 (O_559,N_49939,N_49617);
nand UO_560 (O_560,N_49930,N_49649);
nand UO_561 (O_561,N_49581,N_49699);
nand UO_562 (O_562,N_49715,N_49532);
xnor UO_563 (O_563,N_49728,N_49662);
nand UO_564 (O_564,N_49631,N_49933);
or UO_565 (O_565,N_49575,N_49989);
nand UO_566 (O_566,N_49746,N_49562);
nor UO_567 (O_567,N_49844,N_49596);
nand UO_568 (O_568,N_49591,N_49592);
nand UO_569 (O_569,N_49741,N_49708);
nand UO_570 (O_570,N_49558,N_49854);
and UO_571 (O_571,N_49506,N_49627);
or UO_572 (O_572,N_49591,N_49579);
nor UO_573 (O_573,N_49645,N_49733);
nand UO_574 (O_574,N_49751,N_49793);
nand UO_575 (O_575,N_49947,N_49510);
xnor UO_576 (O_576,N_49741,N_49510);
nor UO_577 (O_577,N_49873,N_49769);
and UO_578 (O_578,N_49812,N_49541);
or UO_579 (O_579,N_49523,N_49504);
nor UO_580 (O_580,N_49721,N_49931);
or UO_581 (O_581,N_49634,N_49758);
or UO_582 (O_582,N_49737,N_49968);
xor UO_583 (O_583,N_49534,N_49835);
nor UO_584 (O_584,N_49992,N_49513);
xnor UO_585 (O_585,N_49715,N_49860);
xnor UO_586 (O_586,N_49910,N_49643);
nand UO_587 (O_587,N_49795,N_49743);
nor UO_588 (O_588,N_49510,N_49689);
and UO_589 (O_589,N_49960,N_49892);
xor UO_590 (O_590,N_49936,N_49777);
xnor UO_591 (O_591,N_49834,N_49804);
and UO_592 (O_592,N_49838,N_49558);
nor UO_593 (O_593,N_49855,N_49888);
or UO_594 (O_594,N_49914,N_49609);
xnor UO_595 (O_595,N_49813,N_49633);
nand UO_596 (O_596,N_49947,N_49712);
nand UO_597 (O_597,N_49621,N_49689);
nor UO_598 (O_598,N_49637,N_49766);
and UO_599 (O_599,N_49602,N_49507);
and UO_600 (O_600,N_49906,N_49547);
nand UO_601 (O_601,N_49716,N_49911);
nor UO_602 (O_602,N_49506,N_49823);
nor UO_603 (O_603,N_49937,N_49871);
and UO_604 (O_604,N_49808,N_49985);
xnor UO_605 (O_605,N_49582,N_49746);
nor UO_606 (O_606,N_49954,N_49550);
and UO_607 (O_607,N_49857,N_49722);
or UO_608 (O_608,N_49988,N_49660);
xor UO_609 (O_609,N_49941,N_49745);
nor UO_610 (O_610,N_49519,N_49668);
xor UO_611 (O_611,N_49666,N_49763);
xnor UO_612 (O_612,N_49582,N_49882);
nand UO_613 (O_613,N_49576,N_49778);
nor UO_614 (O_614,N_49861,N_49552);
xor UO_615 (O_615,N_49580,N_49881);
or UO_616 (O_616,N_49975,N_49999);
nand UO_617 (O_617,N_49593,N_49639);
and UO_618 (O_618,N_49743,N_49786);
nand UO_619 (O_619,N_49611,N_49925);
nand UO_620 (O_620,N_49789,N_49874);
nand UO_621 (O_621,N_49643,N_49902);
nor UO_622 (O_622,N_49627,N_49899);
xor UO_623 (O_623,N_49892,N_49861);
and UO_624 (O_624,N_49874,N_49842);
xnor UO_625 (O_625,N_49984,N_49850);
and UO_626 (O_626,N_49868,N_49588);
or UO_627 (O_627,N_49524,N_49655);
or UO_628 (O_628,N_49605,N_49960);
xor UO_629 (O_629,N_49819,N_49878);
and UO_630 (O_630,N_49896,N_49639);
xor UO_631 (O_631,N_49918,N_49596);
nor UO_632 (O_632,N_49930,N_49657);
and UO_633 (O_633,N_49818,N_49989);
xnor UO_634 (O_634,N_49924,N_49523);
or UO_635 (O_635,N_49762,N_49773);
nand UO_636 (O_636,N_49515,N_49600);
xnor UO_637 (O_637,N_49720,N_49746);
or UO_638 (O_638,N_49807,N_49630);
or UO_639 (O_639,N_49586,N_49950);
xor UO_640 (O_640,N_49718,N_49682);
and UO_641 (O_641,N_49568,N_49532);
or UO_642 (O_642,N_49563,N_49611);
or UO_643 (O_643,N_49835,N_49884);
nor UO_644 (O_644,N_49774,N_49884);
and UO_645 (O_645,N_49914,N_49582);
and UO_646 (O_646,N_49579,N_49828);
nand UO_647 (O_647,N_49713,N_49957);
nand UO_648 (O_648,N_49700,N_49571);
nor UO_649 (O_649,N_49542,N_49895);
nand UO_650 (O_650,N_49685,N_49975);
nand UO_651 (O_651,N_49626,N_49811);
nand UO_652 (O_652,N_49664,N_49812);
nor UO_653 (O_653,N_49860,N_49848);
nor UO_654 (O_654,N_49756,N_49803);
and UO_655 (O_655,N_49535,N_49595);
nand UO_656 (O_656,N_49645,N_49643);
and UO_657 (O_657,N_49864,N_49870);
and UO_658 (O_658,N_49560,N_49572);
and UO_659 (O_659,N_49504,N_49514);
nand UO_660 (O_660,N_49762,N_49634);
xor UO_661 (O_661,N_49986,N_49825);
and UO_662 (O_662,N_49834,N_49783);
and UO_663 (O_663,N_49561,N_49907);
nor UO_664 (O_664,N_49810,N_49664);
nand UO_665 (O_665,N_49658,N_49953);
or UO_666 (O_666,N_49691,N_49519);
nor UO_667 (O_667,N_49932,N_49765);
xor UO_668 (O_668,N_49768,N_49640);
xor UO_669 (O_669,N_49897,N_49504);
or UO_670 (O_670,N_49909,N_49567);
nand UO_671 (O_671,N_49740,N_49796);
and UO_672 (O_672,N_49568,N_49718);
xor UO_673 (O_673,N_49615,N_49510);
nor UO_674 (O_674,N_49748,N_49566);
and UO_675 (O_675,N_49917,N_49997);
or UO_676 (O_676,N_49734,N_49921);
and UO_677 (O_677,N_49504,N_49533);
or UO_678 (O_678,N_49821,N_49544);
nand UO_679 (O_679,N_49890,N_49548);
and UO_680 (O_680,N_49570,N_49754);
xnor UO_681 (O_681,N_49618,N_49800);
nand UO_682 (O_682,N_49850,N_49512);
or UO_683 (O_683,N_49986,N_49946);
and UO_684 (O_684,N_49744,N_49926);
nor UO_685 (O_685,N_49755,N_49885);
nor UO_686 (O_686,N_49546,N_49951);
and UO_687 (O_687,N_49711,N_49503);
nand UO_688 (O_688,N_49954,N_49649);
nand UO_689 (O_689,N_49503,N_49845);
or UO_690 (O_690,N_49711,N_49878);
xor UO_691 (O_691,N_49731,N_49665);
nor UO_692 (O_692,N_49958,N_49779);
or UO_693 (O_693,N_49583,N_49644);
nand UO_694 (O_694,N_49588,N_49708);
nor UO_695 (O_695,N_49615,N_49557);
or UO_696 (O_696,N_49725,N_49813);
and UO_697 (O_697,N_49595,N_49996);
nor UO_698 (O_698,N_49964,N_49787);
xor UO_699 (O_699,N_49955,N_49758);
nand UO_700 (O_700,N_49731,N_49540);
or UO_701 (O_701,N_49532,N_49820);
xor UO_702 (O_702,N_49534,N_49798);
xnor UO_703 (O_703,N_49728,N_49619);
nor UO_704 (O_704,N_49893,N_49750);
or UO_705 (O_705,N_49859,N_49605);
xor UO_706 (O_706,N_49981,N_49701);
nand UO_707 (O_707,N_49915,N_49853);
nand UO_708 (O_708,N_49595,N_49987);
or UO_709 (O_709,N_49944,N_49536);
nor UO_710 (O_710,N_49525,N_49710);
xor UO_711 (O_711,N_49602,N_49783);
and UO_712 (O_712,N_49857,N_49912);
nand UO_713 (O_713,N_49517,N_49818);
and UO_714 (O_714,N_49699,N_49658);
and UO_715 (O_715,N_49623,N_49771);
nor UO_716 (O_716,N_49747,N_49866);
xnor UO_717 (O_717,N_49893,N_49577);
and UO_718 (O_718,N_49865,N_49709);
xnor UO_719 (O_719,N_49976,N_49643);
nor UO_720 (O_720,N_49932,N_49531);
nand UO_721 (O_721,N_49522,N_49512);
or UO_722 (O_722,N_49667,N_49516);
xor UO_723 (O_723,N_49512,N_49943);
nor UO_724 (O_724,N_49635,N_49652);
nor UO_725 (O_725,N_49791,N_49669);
nor UO_726 (O_726,N_49686,N_49573);
nor UO_727 (O_727,N_49582,N_49663);
xor UO_728 (O_728,N_49535,N_49563);
xor UO_729 (O_729,N_49743,N_49722);
nor UO_730 (O_730,N_49515,N_49813);
and UO_731 (O_731,N_49807,N_49727);
nor UO_732 (O_732,N_49753,N_49542);
or UO_733 (O_733,N_49848,N_49727);
or UO_734 (O_734,N_49940,N_49943);
or UO_735 (O_735,N_49621,N_49978);
xor UO_736 (O_736,N_49952,N_49697);
or UO_737 (O_737,N_49602,N_49676);
nand UO_738 (O_738,N_49737,N_49711);
nor UO_739 (O_739,N_49913,N_49879);
or UO_740 (O_740,N_49673,N_49750);
and UO_741 (O_741,N_49601,N_49949);
nor UO_742 (O_742,N_49722,N_49619);
nand UO_743 (O_743,N_49799,N_49879);
nand UO_744 (O_744,N_49846,N_49754);
xnor UO_745 (O_745,N_49644,N_49647);
nand UO_746 (O_746,N_49668,N_49585);
xor UO_747 (O_747,N_49678,N_49857);
nor UO_748 (O_748,N_49959,N_49778);
and UO_749 (O_749,N_49675,N_49643);
or UO_750 (O_750,N_49676,N_49743);
nand UO_751 (O_751,N_49875,N_49992);
nand UO_752 (O_752,N_49915,N_49722);
or UO_753 (O_753,N_49688,N_49844);
nor UO_754 (O_754,N_49882,N_49616);
or UO_755 (O_755,N_49903,N_49801);
nor UO_756 (O_756,N_49699,N_49780);
xnor UO_757 (O_757,N_49521,N_49792);
and UO_758 (O_758,N_49557,N_49672);
nor UO_759 (O_759,N_49765,N_49567);
nor UO_760 (O_760,N_49544,N_49959);
nand UO_761 (O_761,N_49924,N_49676);
xor UO_762 (O_762,N_49511,N_49938);
nor UO_763 (O_763,N_49751,N_49920);
nand UO_764 (O_764,N_49990,N_49604);
nor UO_765 (O_765,N_49767,N_49586);
and UO_766 (O_766,N_49900,N_49876);
xor UO_767 (O_767,N_49943,N_49656);
nor UO_768 (O_768,N_49820,N_49556);
and UO_769 (O_769,N_49894,N_49510);
xor UO_770 (O_770,N_49673,N_49827);
xnor UO_771 (O_771,N_49863,N_49516);
and UO_772 (O_772,N_49875,N_49588);
and UO_773 (O_773,N_49840,N_49569);
nor UO_774 (O_774,N_49670,N_49595);
or UO_775 (O_775,N_49828,N_49830);
xor UO_776 (O_776,N_49898,N_49733);
xnor UO_777 (O_777,N_49709,N_49658);
or UO_778 (O_778,N_49797,N_49810);
and UO_779 (O_779,N_49897,N_49971);
or UO_780 (O_780,N_49890,N_49881);
nand UO_781 (O_781,N_49810,N_49709);
or UO_782 (O_782,N_49735,N_49967);
nor UO_783 (O_783,N_49616,N_49916);
xor UO_784 (O_784,N_49943,N_49523);
nor UO_785 (O_785,N_49612,N_49989);
nor UO_786 (O_786,N_49844,N_49655);
or UO_787 (O_787,N_49868,N_49711);
and UO_788 (O_788,N_49652,N_49705);
nor UO_789 (O_789,N_49614,N_49989);
nor UO_790 (O_790,N_49912,N_49644);
or UO_791 (O_791,N_49713,N_49641);
nand UO_792 (O_792,N_49537,N_49949);
nand UO_793 (O_793,N_49809,N_49597);
nand UO_794 (O_794,N_49652,N_49513);
nand UO_795 (O_795,N_49957,N_49865);
nand UO_796 (O_796,N_49990,N_49564);
xor UO_797 (O_797,N_49832,N_49779);
or UO_798 (O_798,N_49601,N_49999);
xnor UO_799 (O_799,N_49978,N_49508);
nor UO_800 (O_800,N_49617,N_49866);
and UO_801 (O_801,N_49977,N_49591);
and UO_802 (O_802,N_49644,N_49782);
and UO_803 (O_803,N_49969,N_49828);
xnor UO_804 (O_804,N_49806,N_49748);
xnor UO_805 (O_805,N_49772,N_49512);
or UO_806 (O_806,N_49908,N_49784);
and UO_807 (O_807,N_49933,N_49764);
nor UO_808 (O_808,N_49922,N_49573);
and UO_809 (O_809,N_49780,N_49982);
xnor UO_810 (O_810,N_49542,N_49730);
xor UO_811 (O_811,N_49557,N_49995);
nor UO_812 (O_812,N_49944,N_49823);
or UO_813 (O_813,N_49632,N_49703);
and UO_814 (O_814,N_49927,N_49884);
and UO_815 (O_815,N_49650,N_49574);
nor UO_816 (O_816,N_49698,N_49662);
and UO_817 (O_817,N_49677,N_49977);
xor UO_818 (O_818,N_49718,N_49883);
nor UO_819 (O_819,N_49583,N_49710);
nand UO_820 (O_820,N_49987,N_49682);
nand UO_821 (O_821,N_49616,N_49840);
xnor UO_822 (O_822,N_49837,N_49802);
nand UO_823 (O_823,N_49500,N_49852);
or UO_824 (O_824,N_49897,N_49657);
or UO_825 (O_825,N_49726,N_49607);
or UO_826 (O_826,N_49975,N_49518);
or UO_827 (O_827,N_49545,N_49623);
or UO_828 (O_828,N_49662,N_49590);
xnor UO_829 (O_829,N_49511,N_49812);
or UO_830 (O_830,N_49738,N_49978);
nor UO_831 (O_831,N_49942,N_49692);
nand UO_832 (O_832,N_49651,N_49715);
nand UO_833 (O_833,N_49531,N_49871);
or UO_834 (O_834,N_49697,N_49599);
nor UO_835 (O_835,N_49874,N_49903);
and UO_836 (O_836,N_49736,N_49567);
or UO_837 (O_837,N_49981,N_49855);
nor UO_838 (O_838,N_49808,N_49882);
nand UO_839 (O_839,N_49564,N_49741);
nand UO_840 (O_840,N_49663,N_49520);
and UO_841 (O_841,N_49559,N_49836);
and UO_842 (O_842,N_49945,N_49766);
nor UO_843 (O_843,N_49518,N_49801);
nor UO_844 (O_844,N_49685,N_49568);
nand UO_845 (O_845,N_49846,N_49821);
and UO_846 (O_846,N_49823,N_49850);
and UO_847 (O_847,N_49971,N_49806);
or UO_848 (O_848,N_49693,N_49983);
and UO_849 (O_849,N_49646,N_49629);
xor UO_850 (O_850,N_49734,N_49594);
and UO_851 (O_851,N_49961,N_49640);
nor UO_852 (O_852,N_49525,N_49657);
xor UO_853 (O_853,N_49696,N_49837);
and UO_854 (O_854,N_49537,N_49570);
xor UO_855 (O_855,N_49780,N_49871);
nor UO_856 (O_856,N_49751,N_49559);
nor UO_857 (O_857,N_49662,N_49847);
and UO_858 (O_858,N_49642,N_49724);
nand UO_859 (O_859,N_49617,N_49562);
and UO_860 (O_860,N_49619,N_49793);
and UO_861 (O_861,N_49944,N_49744);
and UO_862 (O_862,N_49805,N_49933);
nor UO_863 (O_863,N_49531,N_49847);
and UO_864 (O_864,N_49824,N_49643);
xnor UO_865 (O_865,N_49602,N_49604);
and UO_866 (O_866,N_49954,N_49589);
or UO_867 (O_867,N_49652,N_49611);
nor UO_868 (O_868,N_49556,N_49572);
and UO_869 (O_869,N_49890,N_49811);
nor UO_870 (O_870,N_49724,N_49743);
or UO_871 (O_871,N_49977,N_49948);
nor UO_872 (O_872,N_49743,N_49759);
or UO_873 (O_873,N_49626,N_49847);
nor UO_874 (O_874,N_49794,N_49715);
and UO_875 (O_875,N_49559,N_49536);
nand UO_876 (O_876,N_49995,N_49528);
nand UO_877 (O_877,N_49620,N_49525);
nand UO_878 (O_878,N_49604,N_49794);
nand UO_879 (O_879,N_49615,N_49715);
xor UO_880 (O_880,N_49795,N_49666);
nand UO_881 (O_881,N_49980,N_49777);
nor UO_882 (O_882,N_49574,N_49799);
and UO_883 (O_883,N_49653,N_49862);
and UO_884 (O_884,N_49754,N_49747);
nand UO_885 (O_885,N_49604,N_49647);
nand UO_886 (O_886,N_49579,N_49980);
xnor UO_887 (O_887,N_49828,N_49643);
nand UO_888 (O_888,N_49637,N_49908);
and UO_889 (O_889,N_49861,N_49891);
and UO_890 (O_890,N_49709,N_49803);
nor UO_891 (O_891,N_49829,N_49515);
or UO_892 (O_892,N_49701,N_49836);
or UO_893 (O_893,N_49870,N_49846);
and UO_894 (O_894,N_49720,N_49508);
nand UO_895 (O_895,N_49785,N_49665);
and UO_896 (O_896,N_49729,N_49764);
or UO_897 (O_897,N_49839,N_49743);
nand UO_898 (O_898,N_49555,N_49880);
nor UO_899 (O_899,N_49735,N_49654);
nor UO_900 (O_900,N_49832,N_49724);
and UO_901 (O_901,N_49917,N_49722);
xnor UO_902 (O_902,N_49522,N_49894);
xnor UO_903 (O_903,N_49507,N_49715);
and UO_904 (O_904,N_49571,N_49911);
xnor UO_905 (O_905,N_49606,N_49699);
and UO_906 (O_906,N_49565,N_49620);
nand UO_907 (O_907,N_49815,N_49796);
nand UO_908 (O_908,N_49589,N_49893);
and UO_909 (O_909,N_49779,N_49978);
or UO_910 (O_910,N_49771,N_49884);
and UO_911 (O_911,N_49831,N_49895);
nand UO_912 (O_912,N_49587,N_49860);
nor UO_913 (O_913,N_49524,N_49863);
and UO_914 (O_914,N_49635,N_49513);
xnor UO_915 (O_915,N_49528,N_49968);
xor UO_916 (O_916,N_49557,N_49963);
and UO_917 (O_917,N_49827,N_49629);
nor UO_918 (O_918,N_49979,N_49505);
xnor UO_919 (O_919,N_49537,N_49907);
nor UO_920 (O_920,N_49746,N_49529);
and UO_921 (O_921,N_49904,N_49699);
or UO_922 (O_922,N_49780,N_49561);
xor UO_923 (O_923,N_49789,N_49794);
nor UO_924 (O_924,N_49939,N_49638);
nor UO_925 (O_925,N_49819,N_49811);
xnor UO_926 (O_926,N_49916,N_49561);
nor UO_927 (O_927,N_49674,N_49589);
or UO_928 (O_928,N_49609,N_49834);
and UO_929 (O_929,N_49944,N_49820);
and UO_930 (O_930,N_49693,N_49902);
or UO_931 (O_931,N_49916,N_49953);
nand UO_932 (O_932,N_49814,N_49805);
nand UO_933 (O_933,N_49769,N_49713);
xnor UO_934 (O_934,N_49912,N_49903);
nand UO_935 (O_935,N_49929,N_49697);
nand UO_936 (O_936,N_49589,N_49717);
nand UO_937 (O_937,N_49859,N_49660);
xnor UO_938 (O_938,N_49816,N_49963);
nand UO_939 (O_939,N_49530,N_49633);
or UO_940 (O_940,N_49856,N_49532);
nor UO_941 (O_941,N_49995,N_49886);
nor UO_942 (O_942,N_49749,N_49748);
xnor UO_943 (O_943,N_49779,N_49941);
nor UO_944 (O_944,N_49811,N_49856);
nor UO_945 (O_945,N_49701,N_49620);
xor UO_946 (O_946,N_49951,N_49805);
xnor UO_947 (O_947,N_49892,N_49680);
xnor UO_948 (O_948,N_49824,N_49729);
or UO_949 (O_949,N_49624,N_49805);
xor UO_950 (O_950,N_49806,N_49538);
and UO_951 (O_951,N_49652,N_49993);
nor UO_952 (O_952,N_49755,N_49563);
nand UO_953 (O_953,N_49693,N_49863);
nor UO_954 (O_954,N_49711,N_49880);
xor UO_955 (O_955,N_49573,N_49753);
xor UO_956 (O_956,N_49903,N_49773);
and UO_957 (O_957,N_49875,N_49784);
or UO_958 (O_958,N_49537,N_49955);
nand UO_959 (O_959,N_49815,N_49574);
nor UO_960 (O_960,N_49750,N_49558);
nor UO_961 (O_961,N_49548,N_49654);
nand UO_962 (O_962,N_49573,N_49648);
nand UO_963 (O_963,N_49819,N_49751);
xnor UO_964 (O_964,N_49696,N_49687);
nor UO_965 (O_965,N_49890,N_49812);
nand UO_966 (O_966,N_49511,N_49538);
nand UO_967 (O_967,N_49663,N_49636);
or UO_968 (O_968,N_49603,N_49630);
nor UO_969 (O_969,N_49702,N_49810);
xor UO_970 (O_970,N_49642,N_49845);
xor UO_971 (O_971,N_49786,N_49596);
nor UO_972 (O_972,N_49622,N_49877);
or UO_973 (O_973,N_49917,N_49852);
and UO_974 (O_974,N_49956,N_49911);
nor UO_975 (O_975,N_49855,N_49701);
xor UO_976 (O_976,N_49909,N_49514);
nand UO_977 (O_977,N_49762,N_49983);
nor UO_978 (O_978,N_49510,N_49869);
or UO_979 (O_979,N_49754,N_49779);
and UO_980 (O_980,N_49602,N_49757);
nor UO_981 (O_981,N_49623,N_49507);
xnor UO_982 (O_982,N_49711,N_49541);
xor UO_983 (O_983,N_49619,N_49596);
and UO_984 (O_984,N_49814,N_49682);
and UO_985 (O_985,N_49976,N_49542);
nor UO_986 (O_986,N_49838,N_49841);
nand UO_987 (O_987,N_49686,N_49882);
and UO_988 (O_988,N_49580,N_49533);
nor UO_989 (O_989,N_49662,N_49809);
nor UO_990 (O_990,N_49592,N_49580);
xor UO_991 (O_991,N_49660,N_49735);
and UO_992 (O_992,N_49857,N_49705);
nand UO_993 (O_993,N_49919,N_49664);
xnor UO_994 (O_994,N_49952,N_49824);
xnor UO_995 (O_995,N_49772,N_49705);
nor UO_996 (O_996,N_49938,N_49643);
nor UO_997 (O_997,N_49881,N_49663);
xnor UO_998 (O_998,N_49905,N_49910);
nor UO_999 (O_999,N_49833,N_49760);
nand UO_1000 (O_1000,N_49652,N_49691);
nand UO_1001 (O_1001,N_49682,N_49924);
or UO_1002 (O_1002,N_49803,N_49724);
or UO_1003 (O_1003,N_49880,N_49879);
and UO_1004 (O_1004,N_49699,N_49663);
nand UO_1005 (O_1005,N_49987,N_49991);
and UO_1006 (O_1006,N_49786,N_49848);
or UO_1007 (O_1007,N_49631,N_49673);
nor UO_1008 (O_1008,N_49885,N_49731);
or UO_1009 (O_1009,N_49749,N_49953);
or UO_1010 (O_1010,N_49596,N_49547);
nor UO_1011 (O_1011,N_49783,N_49969);
nor UO_1012 (O_1012,N_49635,N_49666);
nand UO_1013 (O_1013,N_49698,N_49909);
nand UO_1014 (O_1014,N_49635,N_49889);
or UO_1015 (O_1015,N_49970,N_49774);
or UO_1016 (O_1016,N_49865,N_49595);
nor UO_1017 (O_1017,N_49878,N_49578);
xor UO_1018 (O_1018,N_49625,N_49821);
nor UO_1019 (O_1019,N_49865,N_49678);
or UO_1020 (O_1020,N_49610,N_49673);
nand UO_1021 (O_1021,N_49545,N_49725);
xor UO_1022 (O_1022,N_49591,N_49996);
xnor UO_1023 (O_1023,N_49821,N_49624);
and UO_1024 (O_1024,N_49682,N_49667);
nor UO_1025 (O_1025,N_49953,N_49506);
nand UO_1026 (O_1026,N_49555,N_49829);
and UO_1027 (O_1027,N_49888,N_49902);
and UO_1028 (O_1028,N_49808,N_49887);
xnor UO_1029 (O_1029,N_49961,N_49895);
or UO_1030 (O_1030,N_49785,N_49615);
nand UO_1031 (O_1031,N_49619,N_49752);
and UO_1032 (O_1032,N_49966,N_49805);
nor UO_1033 (O_1033,N_49909,N_49517);
nand UO_1034 (O_1034,N_49746,N_49780);
nand UO_1035 (O_1035,N_49950,N_49911);
or UO_1036 (O_1036,N_49892,N_49580);
nor UO_1037 (O_1037,N_49534,N_49725);
nor UO_1038 (O_1038,N_49698,N_49801);
or UO_1039 (O_1039,N_49702,N_49670);
nor UO_1040 (O_1040,N_49863,N_49887);
nor UO_1041 (O_1041,N_49729,N_49866);
and UO_1042 (O_1042,N_49720,N_49822);
xor UO_1043 (O_1043,N_49571,N_49829);
or UO_1044 (O_1044,N_49718,N_49533);
or UO_1045 (O_1045,N_49544,N_49541);
xor UO_1046 (O_1046,N_49510,N_49806);
nand UO_1047 (O_1047,N_49744,N_49897);
nor UO_1048 (O_1048,N_49630,N_49685);
and UO_1049 (O_1049,N_49754,N_49613);
xor UO_1050 (O_1050,N_49772,N_49948);
xor UO_1051 (O_1051,N_49933,N_49860);
and UO_1052 (O_1052,N_49794,N_49940);
nor UO_1053 (O_1053,N_49718,N_49837);
xor UO_1054 (O_1054,N_49730,N_49757);
and UO_1055 (O_1055,N_49561,N_49827);
or UO_1056 (O_1056,N_49655,N_49954);
and UO_1057 (O_1057,N_49631,N_49640);
nor UO_1058 (O_1058,N_49681,N_49628);
xnor UO_1059 (O_1059,N_49840,N_49529);
xnor UO_1060 (O_1060,N_49761,N_49522);
or UO_1061 (O_1061,N_49706,N_49527);
nor UO_1062 (O_1062,N_49800,N_49976);
nor UO_1063 (O_1063,N_49627,N_49939);
and UO_1064 (O_1064,N_49622,N_49671);
nand UO_1065 (O_1065,N_49535,N_49742);
nand UO_1066 (O_1066,N_49626,N_49560);
nand UO_1067 (O_1067,N_49749,N_49844);
and UO_1068 (O_1068,N_49564,N_49855);
xor UO_1069 (O_1069,N_49939,N_49589);
or UO_1070 (O_1070,N_49838,N_49944);
xor UO_1071 (O_1071,N_49543,N_49903);
nor UO_1072 (O_1072,N_49933,N_49918);
nor UO_1073 (O_1073,N_49539,N_49736);
xnor UO_1074 (O_1074,N_49918,N_49983);
nor UO_1075 (O_1075,N_49893,N_49596);
nor UO_1076 (O_1076,N_49528,N_49506);
nor UO_1077 (O_1077,N_49959,N_49694);
nor UO_1078 (O_1078,N_49511,N_49598);
nor UO_1079 (O_1079,N_49515,N_49912);
xor UO_1080 (O_1080,N_49938,N_49798);
and UO_1081 (O_1081,N_49779,N_49536);
xor UO_1082 (O_1082,N_49801,N_49500);
or UO_1083 (O_1083,N_49639,N_49899);
xor UO_1084 (O_1084,N_49915,N_49860);
nor UO_1085 (O_1085,N_49893,N_49625);
or UO_1086 (O_1086,N_49687,N_49661);
xnor UO_1087 (O_1087,N_49681,N_49879);
nor UO_1088 (O_1088,N_49902,N_49753);
nand UO_1089 (O_1089,N_49996,N_49536);
or UO_1090 (O_1090,N_49986,N_49848);
and UO_1091 (O_1091,N_49640,N_49615);
xor UO_1092 (O_1092,N_49939,N_49595);
nand UO_1093 (O_1093,N_49931,N_49609);
nor UO_1094 (O_1094,N_49507,N_49506);
xor UO_1095 (O_1095,N_49672,N_49673);
or UO_1096 (O_1096,N_49828,N_49918);
and UO_1097 (O_1097,N_49751,N_49569);
nand UO_1098 (O_1098,N_49719,N_49731);
and UO_1099 (O_1099,N_49688,N_49680);
and UO_1100 (O_1100,N_49919,N_49745);
or UO_1101 (O_1101,N_49707,N_49666);
nor UO_1102 (O_1102,N_49839,N_49581);
nand UO_1103 (O_1103,N_49862,N_49530);
xor UO_1104 (O_1104,N_49738,N_49846);
xnor UO_1105 (O_1105,N_49534,N_49531);
xor UO_1106 (O_1106,N_49868,N_49781);
xnor UO_1107 (O_1107,N_49828,N_49944);
nand UO_1108 (O_1108,N_49660,N_49691);
xor UO_1109 (O_1109,N_49982,N_49601);
nand UO_1110 (O_1110,N_49596,N_49890);
and UO_1111 (O_1111,N_49653,N_49741);
nand UO_1112 (O_1112,N_49747,N_49568);
xor UO_1113 (O_1113,N_49930,N_49659);
and UO_1114 (O_1114,N_49738,N_49787);
nand UO_1115 (O_1115,N_49776,N_49899);
xor UO_1116 (O_1116,N_49805,N_49934);
nand UO_1117 (O_1117,N_49727,N_49619);
nand UO_1118 (O_1118,N_49728,N_49792);
xor UO_1119 (O_1119,N_49915,N_49667);
and UO_1120 (O_1120,N_49847,N_49695);
nand UO_1121 (O_1121,N_49528,N_49749);
nor UO_1122 (O_1122,N_49761,N_49774);
nor UO_1123 (O_1123,N_49949,N_49517);
or UO_1124 (O_1124,N_49698,N_49621);
nor UO_1125 (O_1125,N_49782,N_49853);
xor UO_1126 (O_1126,N_49907,N_49913);
and UO_1127 (O_1127,N_49589,N_49777);
nand UO_1128 (O_1128,N_49532,N_49607);
xnor UO_1129 (O_1129,N_49569,N_49502);
nand UO_1130 (O_1130,N_49834,N_49646);
nor UO_1131 (O_1131,N_49606,N_49830);
nand UO_1132 (O_1132,N_49951,N_49646);
nand UO_1133 (O_1133,N_49743,N_49739);
and UO_1134 (O_1134,N_49721,N_49854);
nor UO_1135 (O_1135,N_49520,N_49928);
or UO_1136 (O_1136,N_49988,N_49644);
and UO_1137 (O_1137,N_49801,N_49842);
xor UO_1138 (O_1138,N_49693,N_49808);
nand UO_1139 (O_1139,N_49973,N_49782);
or UO_1140 (O_1140,N_49703,N_49623);
and UO_1141 (O_1141,N_49522,N_49867);
nand UO_1142 (O_1142,N_49666,N_49529);
or UO_1143 (O_1143,N_49818,N_49645);
or UO_1144 (O_1144,N_49966,N_49736);
xnor UO_1145 (O_1145,N_49649,N_49958);
nand UO_1146 (O_1146,N_49771,N_49726);
or UO_1147 (O_1147,N_49662,N_49848);
or UO_1148 (O_1148,N_49726,N_49556);
or UO_1149 (O_1149,N_49851,N_49794);
nand UO_1150 (O_1150,N_49661,N_49529);
xor UO_1151 (O_1151,N_49842,N_49745);
or UO_1152 (O_1152,N_49907,N_49912);
and UO_1153 (O_1153,N_49662,N_49692);
or UO_1154 (O_1154,N_49579,N_49546);
or UO_1155 (O_1155,N_49980,N_49915);
and UO_1156 (O_1156,N_49854,N_49931);
and UO_1157 (O_1157,N_49791,N_49709);
and UO_1158 (O_1158,N_49667,N_49687);
nand UO_1159 (O_1159,N_49736,N_49523);
xnor UO_1160 (O_1160,N_49657,N_49664);
and UO_1161 (O_1161,N_49869,N_49588);
and UO_1162 (O_1162,N_49640,N_49638);
and UO_1163 (O_1163,N_49525,N_49646);
xnor UO_1164 (O_1164,N_49521,N_49721);
nor UO_1165 (O_1165,N_49831,N_49589);
and UO_1166 (O_1166,N_49635,N_49668);
nand UO_1167 (O_1167,N_49548,N_49776);
nor UO_1168 (O_1168,N_49591,N_49718);
nand UO_1169 (O_1169,N_49751,N_49537);
and UO_1170 (O_1170,N_49645,N_49918);
nor UO_1171 (O_1171,N_49890,N_49809);
nor UO_1172 (O_1172,N_49787,N_49568);
or UO_1173 (O_1173,N_49829,N_49603);
and UO_1174 (O_1174,N_49823,N_49501);
nand UO_1175 (O_1175,N_49789,N_49785);
nor UO_1176 (O_1176,N_49582,N_49692);
or UO_1177 (O_1177,N_49628,N_49886);
xnor UO_1178 (O_1178,N_49546,N_49962);
xor UO_1179 (O_1179,N_49761,N_49992);
nor UO_1180 (O_1180,N_49948,N_49857);
or UO_1181 (O_1181,N_49658,N_49898);
nand UO_1182 (O_1182,N_49575,N_49836);
and UO_1183 (O_1183,N_49762,N_49769);
nand UO_1184 (O_1184,N_49647,N_49810);
nor UO_1185 (O_1185,N_49784,N_49599);
or UO_1186 (O_1186,N_49977,N_49522);
xnor UO_1187 (O_1187,N_49905,N_49671);
xnor UO_1188 (O_1188,N_49810,N_49853);
xor UO_1189 (O_1189,N_49931,N_49512);
or UO_1190 (O_1190,N_49689,N_49770);
and UO_1191 (O_1191,N_49893,N_49736);
nor UO_1192 (O_1192,N_49929,N_49759);
nor UO_1193 (O_1193,N_49810,N_49926);
or UO_1194 (O_1194,N_49562,N_49795);
and UO_1195 (O_1195,N_49856,N_49721);
and UO_1196 (O_1196,N_49960,N_49871);
or UO_1197 (O_1197,N_49582,N_49597);
xor UO_1198 (O_1198,N_49913,N_49679);
and UO_1199 (O_1199,N_49796,N_49500);
or UO_1200 (O_1200,N_49593,N_49560);
or UO_1201 (O_1201,N_49505,N_49574);
xor UO_1202 (O_1202,N_49500,N_49605);
or UO_1203 (O_1203,N_49764,N_49711);
nand UO_1204 (O_1204,N_49661,N_49543);
or UO_1205 (O_1205,N_49892,N_49853);
nand UO_1206 (O_1206,N_49977,N_49900);
or UO_1207 (O_1207,N_49975,N_49719);
xor UO_1208 (O_1208,N_49616,N_49805);
xnor UO_1209 (O_1209,N_49961,N_49516);
nor UO_1210 (O_1210,N_49616,N_49863);
nand UO_1211 (O_1211,N_49914,N_49986);
xor UO_1212 (O_1212,N_49839,N_49562);
or UO_1213 (O_1213,N_49516,N_49579);
xnor UO_1214 (O_1214,N_49646,N_49586);
nor UO_1215 (O_1215,N_49551,N_49578);
nor UO_1216 (O_1216,N_49502,N_49633);
nand UO_1217 (O_1217,N_49531,N_49809);
and UO_1218 (O_1218,N_49952,N_49872);
or UO_1219 (O_1219,N_49593,N_49646);
nor UO_1220 (O_1220,N_49546,N_49829);
nand UO_1221 (O_1221,N_49908,N_49886);
and UO_1222 (O_1222,N_49630,N_49714);
or UO_1223 (O_1223,N_49617,N_49762);
nor UO_1224 (O_1224,N_49639,N_49826);
and UO_1225 (O_1225,N_49808,N_49540);
xnor UO_1226 (O_1226,N_49548,N_49917);
nor UO_1227 (O_1227,N_49929,N_49904);
nand UO_1228 (O_1228,N_49924,N_49979);
or UO_1229 (O_1229,N_49911,N_49746);
and UO_1230 (O_1230,N_49694,N_49608);
nor UO_1231 (O_1231,N_49897,N_49658);
or UO_1232 (O_1232,N_49925,N_49511);
xor UO_1233 (O_1233,N_49934,N_49667);
and UO_1234 (O_1234,N_49768,N_49825);
xnor UO_1235 (O_1235,N_49811,N_49652);
and UO_1236 (O_1236,N_49948,N_49924);
and UO_1237 (O_1237,N_49606,N_49914);
nand UO_1238 (O_1238,N_49624,N_49522);
xnor UO_1239 (O_1239,N_49715,N_49528);
or UO_1240 (O_1240,N_49974,N_49986);
nor UO_1241 (O_1241,N_49838,N_49738);
and UO_1242 (O_1242,N_49554,N_49565);
nand UO_1243 (O_1243,N_49997,N_49871);
and UO_1244 (O_1244,N_49681,N_49700);
xnor UO_1245 (O_1245,N_49771,N_49632);
or UO_1246 (O_1246,N_49615,N_49642);
or UO_1247 (O_1247,N_49656,N_49627);
nand UO_1248 (O_1248,N_49897,N_49517);
and UO_1249 (O_1249,N_49936,N_49969);
nand UO_1250 (O_1250,N_49660,N_49997);
or UO_1251 (O_1251,N_49888,N_49598);
nand UO_1252 (O_1252,N_49502,N_49983);
xor UO_1253 (O_1253,N_49522,N_49876);
nand UO_1254 (O_1254,N_49802,N_49629);
xnor UO_1255 (O_1255,N_49979,N_49879);
or UO_1256 (O_1256,N_49841,N_49961);
nor UO_1257 (O_1257,N_49672,N_49963);
nor UO_1258 (O_1258,N_49815,N_49853);
nand UO_1259 (O_1259,N_49959,N_49974);
nor UO_1260 (O_1260,N_49625,N_49929);
xnor UO_1261 (O_1261,N_49541,N_49676);
or UO_1262 (O_1262,N_49565,N_49959);
and UO_1263 (O_1263,N_49628,N_49719);
nor UO_1264 (O_1264,N_49756,N_49728);
or UO_1265 (O_1265,N_49875,N_49793);
or UO_1266 (O_1266,N_49793,N_49578);
nor UO_1267 (O_1267,N_49566,N_49691);
xnor UO_1268 (O_1268,N_49622,N_49714);
nor UO_1269 (O_1269,N_49556,N_49650);
xor UO_1270 (O_1270,N_49629,N_49563);
nor UO_1271 (O_1271,N_49688,N_49789);
and UO_1272 (O_1272,N_49753,N_49597);
xor UO_1273 (O_1273,N_49986,N_49832);
or UO_1274 (O_1274,N_49775,N_49624);
or UO_1275 (O_1275,N_49648,N_49639);
nor UO_1276 (O_1276,N_49946,N_49987);
nor UO_1277 (O_1277,N_49970,N_49691);
and UO_1278 (O_1278,N_49731,N_49706);
xor UO_1279 (O_1279,N_49983,N_49614);
and UO_1280 (O_1280,N_49709,N_49699);
nand UO_1281 (O_1281,N_49676,N_49826);
nand UO_1282 (O_1282,N_49741,N_49744);
or UO_1283 (O_1283,N_49876,N_49831);
or UO_1284 (O_1284,N_49802,N_49688);
or UO_1285 (O_1285,N_49869,N_49987);
nand UO_1286 (O_1286,N_49935,N_49623);
xor UO_1287 (O_1287,N_49961,N_49815);
nand UO_1288 (O_1288,N_49694,N_49708);
or UO_1289 (O_1289,N_49964,N_49657);
or UO_1290 (O_1290,N_49578,N_49718);
nor UO_1291 (O_1291,N_49903,N_49800);
or UO_1292 (O_1292,N_49740,N_49628);
nor UO_1293 (O_1293,N_49895,N_49729);
nand UO_1294 (O_1294,N_49555,N_49572);
nand UO_1295 (O_1295,N_49811,N_49788);
or UO_1296 (O_1296,N_49721,N_49599);
or UO_1297 (O_1297,N_49864,N_49688);
nand UO_1298 (O_1298,N_49733,N_49792);
nor UO_1299 (O_1299,N_49797,N_49644);
nor UO_1300 (O_1300,N_49531,N_49662);
xor UO_1301 (O_1301,N_49865,N_49769);
nor UO_1302 (O_1302,N_49734,N_49758);
nor UO_1303 (O_1303,N_49741,N_49813);
nor UO_1304 (O_1304,N_49656,N_49613);
nand UO_1305 (O_1305,N_49864,N_49826);
and UO_1306 (O_1306,N_49913,N_49661);
nand UO_1307 (O_1307,N_49849,N_49598);
nor UO_1308 (O_1308,N_49797,N_49989);
nor UO_1309 (O_1309,N_49525,N_49825);
nand UO_1310 (O_1310,N_49584,N_49661);
nor UO_1311 (O_1311,N_49988,N_49776);
xnor UO_1312 (O_1312,N_49522,N_49635);
nor UO_1313 (O_1313,N_49780,N_49875);
xor UO_1314 (O_1314,N_49790,N_49615);
nor UO_1315 (O_1315,N_49758,N_49909);
nor UO_1316 (O_1316,N_49852,N_49652);
and UO_1317 (O_1317,N_49534,N_49952);
xor UO_1318 (O_1318,N_49849,N_49930);
and UO_1319 (O_1319,N_49525,N_49997);
or UO_1320 (O_1320,N_49670,N_49916);
nand UO_1321 (O_1321,N_49524,N_49936);
nand UO_1322 (O_1322,N_49642,N_49783);
nand UO_1323 (O_1323,N_49859,N_49807);
and UO_1324 (O_1324,N_49792,N_49641);
nand UO_1325 (O_1325,N_49964,N_49867);
xor UO_1326 (O_1326,N_49922,N_49878);
and UO_1327 (O_1327,N_49734,N_49547);
or UO_1328 (O_1328,N_49805,N_49612);
nand UO_1329 (O_1329,N_49705,N_49710);
or UO_1330 (O_1330,N_49681,N_49817);
nand UO_1331 (O_1331,N_49933,N_49991);
nor UO_1332 (O_1332,N_49543,N_49592);
nand UO_1333 (O_1333,N_49509,N_49760);
or UO_1334 (O_1334,N_49558,N_49916);
nand UO_1335 (O_1335,N_49843,N_49917);
and UO_1336 (O_1336,N_49564,N_49955);
nand UO_1337 (O_1337,N_49691,N_49515);
nor UO_1338 (O_1338,N_49959,N_49967);
nand UO_1339 (O_1339,N_49618,N_49878);
xor UO_1340 (O_1340,N_49529,N_49744);
and UO_1341 (O_1341,N_49535,N_49905);
or UO_1342 (O_1342,N_49832,N_49649);
xor UO_1343 (O_1343,N_49931,N_49582);
xor UO_1344 (O_1344,N_49728,N_49949);
nor UO_1345 (O_1345,N_49969,N_49785);
and UO_1346 (O_1346,N_49651,N_49686);
and UO_1347 (O_1347,N_49812,N_49786);
xnor UO_1348 (O_1348,N_49655,N_49578);
xnor UO_1349 (O_1349,N_49939,N_49794);
nand UO_1350 (O_1350,N_49977,N_49869);
xor UO_1351 (O_1351,N_49799,N_49608);
xnor UO_1352 (O_1352,N_49879,N_49878);
nor UO_1353 (O_1353,N_49573,N_49844);
and UO_1354 (O_1354,N_49716,N_49631);
xor UO_1355 (O_1355,N_49640,N_49689);
and UO_1356 (O_1356,N_49759,N_49815);
or UO_1357 (O_1357,N_49888,N_49813);
nor UO_1358 (O_1358,N_49702,N_49848);
nand UO_1359 (O_1359,N_49876,N_49634);
xor UO_1360 (O_1360,N_49785,N_49594);
xnor UO_1361 (O_1361,N_49964,N_49784);
and UO_1362 (O_1362,N_49933,N_49559);
xnor UO_1363 (O_1363,N_49956,N_49973);
xor UO_1364 (O_1364,N_49872,N_49848);
nor UO_1365 (O_1365,N_49827,N_49814);
xor UO_1366 (O_1366,N_49713,N_49772);
xor UO_1367 (O_1367,N_49692,N_49845);
or UO_1368 (O_1368,N_49782,N_49678);
nand UO_1369 (O_1369,N_49941,N_49665);
nand UO_1370 (O_1370,N_49694,N_49558);
and UO_1371 (O_1371,N_49764,N_49993);
xnor UO_1372 (O_1372,N_49899,N_49643);
nor UO_1373 (O_1373,N_49637,N_49721);
nor UO_1374 (O_1374,N_49878,N_49605);
nor UO_1375 (O_1375,N_49727,N_49936);
xnor UO_1376 (O_1376,N_49958,N_49791);
xnor UO_1377 (O_1377,N_49933,N_49654);
or UO_1378 (O_1378,N_49891,N_49559);
nor UO_1379 (O_1379,N_49997,N_49888);
xor UO_1380 (O_1380,N_49994,N_49683);
and UO_1381 (O_1381,N_49912,N_49993);
nor UO_1382 (O_1382,N_49871,N_49554);
xnor UO_1383 (O_1383,N_49666,N_49661);
nand UO_1384 (O_1384,N_49847,N_49972);
xor UO_1385 (O_1385,N_49745,N_49952);
xor UO_1386 (O_1386,N_49536,N_49711);
or UO_1387 (O_1387,N_49505,N_49904);
and UO_1388 (O_1388,N_49878,N_49658);
and UO_1389 (O_1389,N_49525,N_49568);
xnor UO_1390 (O_1390,N_49749,N_49628);
nand UO_1391 (O_1391,N_49775,N_49931);
and UO_1392 (O_1392,N_49554,N_49872);
or UO_1393 (O_1393,N_49513,N_49979);
xnor UO_1394 (O_1394,N_49694,N_49987);
nand UO_1395 (O_1395,N_49921,N_49724);
and UO_1396 (O_1396,N_49764,N_49889);
nand UO_1397 (O_1397,N_49530,N_49587);
or UO_1398 (O_1398,N_49728,N_49848);
nand UO_1399 (O_1399,N_49960,N_49500);
nand UO_1400 (O_1400,N_49835,N_49802);
nand UO_1401 (O_1401,N_49984,N_49892);
xor UO_1402 (O_1402,N_49942,N_49583);
or UO_1403 (O_1403,N_49878,N_49996);
xnor UO_1404 (O_1404,N_49566,N_49810);
xor UO_1405 (O_1405,N_49797,N_49849);
or UO_1406 (O_1406,N_49817,N_49801);
nand UO_1407 (O_1407,N_49692,N_49664);
nand UO_1408 (O_1408,N_49626,N_49952);
xor UO_1409 (O_1409,N_49955,N_49730);
nand UO_1410 (O_1410,N_49667,N_49596);
xor UO_1411 (O_1411,N_49700,N_49896);
xnor UO_1412 (O_1412,N_49763,N_49758);
nor UO_1413 (O_1413,N_49760,N_49564);
nor UO_1414 (O_1414,N_49619,N_49889);
nand UO_1415 (O_1415,N_49939,N_49593);
or UO_1416 (O_1416,N_49883,N_49671);
nand UO_1417 (O_1417,N_49870,N_49961);
nand UO_1418 (O_1418,N_49609,N_49537);
xor UO_1419 (O_1419,N_49901,N_49588);
xnor UO_1420 (O_1420,N_49782,N_49658);
xor UO_1421 (O_1421,N_49504,N_49569);
xor UO_1422 (O_1422,N_49528,N_49989);
nor UO_1423 (O_1423,N_49958,N_49832);
xor UO_1424 (O_1424,N_49594,N_49662);
or UO_1425 (O_1425,N_49931,N_49665);
nor UO_1426 (O_1426,N_49520,N_49889);
xor UO_1427 (O_1427,N_49855,N_49749);
nand UO_1428 (O_1428,N_49915,N_49544);
xor UO_1429 (O_1429,N_49791,N_49700);
and UO_1430 (O_1430,N_49510,N_49577);
or UO_1431 (O_1431,N_49784,N_49801);
or UO_1432 (O_1432,N_49763,N_49783);
xor UO_1433 (O_1433,N_49619,N_49881);
or UO_1434 (O_1434,N_49763,N_49796);
or UO_1435 (O_1435,N_49850,N_49680);
or UO_1436 (O_1436,N_49618,N_49938);
nor UO_1437 (O_1437,N_49706,N_49959);
nor UO_1438 (O_1438,N_49633,N_49708);
xnor UO_1439 (O_1439,N_49862,N_49781);
and UO_1440 (O_1440,N_49948,N_49710);
nand UO_1441 (O_1441,N_49972,N_49591);
nor UO_1442 (O_1442,N_49794,N_49925);
xnor UO_1443 (O_1443,N_49827,N_49640);
xnor UO_1444 (O_1444,N_49509,N_49888);
nor UO_1445 (O_1445,N_49745,N_49609);
nor UO_1446 (O_1446,N_49699,N_49828);
xnor UO_1447 (O_1447,N_49556,N_49707);
nor UO_1448 (O_1448,N_49970,N_49515);
nand UO_1449 (O_1449,N_49709,N_49581);
xnor UO_1450 (O_1450,N_49713,N_49664);
and UO_1451 (O_1451,N_49597,N_49637);
and UO_1452 (O_1452,N_49551,N_49933);
nand UO_1453 (O_1453,N_49942,N_49662);
and UO_1454 (O_1454,N_49715,N_49911);
and UO_1455 (O_1455,N_49907,N_49858);
nor UO_1456 (O_1456,N_49617,N_49821);
and UO_1457 (O_1457,N_49523,N_49590);
nand UO_1458 (O_1458,N_49943,N_49511);
nor UO_1459 (O_1459,N_49821,N_49663);
and UO_1460 (O_1460,N_49930,N_49747);
xnor UO_1461 (O_1461,N_49820,N_49926);
nand UO_1462 (O_1462,N_49827,N_49698);
xor UO_1463 (O_1463,N_49716,N_49777);
and UO_1464 (O_1464,N_49729,N_49763);
xnor UO_1465 (O_1465,N_49608,N_49915);
nand UO_1466 (O_1466,N_49640,N_49659);
nor UO_1467 (O_1467,N_49999,N_49775);
and UO_1468 (O_1468,N_49547,N_49934);
nor UO_1469 (O_1469,N_49779,N_49549);
or UO_1470 (O_1470,N_49610,N_49853);
nand UO_1471 (O_1471,N_49617,N_49981);
nand UO_1472 (O_1472,N_49961,N_49708);
xor UO_1473 (O_1473,N_49581,N_49534);
and UO_1474 (O_1474,N_49779,N_49842);
and UO_1475 (O_1475,N_49509,N_49593);
nand UO_1476 (O_1476,N_49893,N_49622);
nand UO_1477 (O_1477,N_49722,N_49555);
nor UO_1478 (O_1478,N_49640,N_49646);
xnor UO_1479 (O_1479,N_49747,N_49561);
or UO_1480 (O_1480,N_49915,N_49990);
nor UO_1481 (O_1481,N_49789,N_49612);
nor UO_1482 (O_1482,N_49592,N_49559);
and UO_1483 (O_1483,N_49789,N_49924);
or UO_1484 (O_1484,N_49687,N_49821);
or UO_1485 (O_1485,N_49660,N_49673);
nor UO_1486 (O_1486,N_49844,N_49955);
nor UO_1487 (O_1487,N_49742,N_49732);
xnor UO_1488 (O_1488,N_49754,N_49523);
nor UO_1489 (O_1489,N_49634,N_49865);
and UO_1490 (O_1490,N_49989,N_49802);
or UO_1491 (O_1491,N_49617,N_49788);
nand UO_1492 (O_1492,N_49841,N_49917);
nand UO_1493 (O_1493,N_49921,N_49983);
or UO_1494 (O_1494,N_49775,N_49657);
nand UO_1495 (O_1495,N_49531,N_49719);
xnor UO_1496 (O_1496,N_49864,N_49843);
and UO_1497 (O_1497,N_49660,N_49887);
nand UO_1498 (O_1498,N_49621,N_49922);
xor UO_1499 (O_1499,N_49992,N_49872);
and UO_1500 (O_1500,N_49565,N_49884);
nor UO_1501 (O_1501,N_49830,N_49597);
nor UO_1502 (O_1502,N_49814,N_49896);
and UO_1503 (O_1503,N_49784,N_49863);
and UO_1504 (O_1504,N_49846,N_49614);
xor UO_1505 (O_1505,N_49979,N_49695);
nand UO_1506 (O_1506,N_49852,N_49735);
or UO_1507 (O_1507,N_49997,N_49969);
and UO_1508 (O_1508,N_49933,N_49762);
nor UO_1509 (O_1509,N_49962,N_49911);
nand UO_1510 (O_1510,N_49759,N_49968);
nand UO_1511 (O_1511,N_49900,N_49777);
nor UO_1512 (O_1512,N_49948,N_49934);
and UO_1513 (O_1513,N_49643,N_49705);
and UO_1514 (O_1514,N_49574,N_49976);
and UO_1515 (O_1515,N_49541,N_49910);
and UO_1516 (O_1516,N_49752,N_49784);
and UO_1517 (O_1517,N_49747,N_49736);
and UO_1518 (O_1518,N_49739,N_49550);
nor UO_1519 (O_1519,N_49629,N_49834);
xnor UO_1520 (O_1520,N_49883,N_49635);
nor UO_1521 (O_1521,N_49950,N_49712);
or UO_1522 (O_1522,N_49670,N_49872);
and UO_1523 (O_1523,N_49766,N_49802);
nand UO_1524 (O_1524,N_49731,N_49770);
or UO_1525 (O_1525,N_49974,N_49585);
and UO_1526 (O_1526,N_49856,N_49916);
and UO_1527 (O_1527,N_49861,N_49695);
xnor UO_1528 (O_1528,N_49522,N_49958);
nor UO_1529 (O_1529,N_49917,N_49566);
nand UO_1530 (O_1530,N_49506,N_49641);
or UO_1531 (O_1531,N_49648,N_49757);
or UO_1532 (O_1532,N_49502,N_49570);
nor UO_1533 (O_1533,N_49539,N_49938);
xor UO_1534 (O_1534,N_49503,N_49728);
xnor UO_1535 (O_1535,N_49768,N_49821);
nor UO_1536 (O_1536,N_49962,N_49540);
xnor UO_1537 (O_1537,N_49748,N_49755);
or UO_1538 (O_1538,N_49735,N_49915);
nor UO_1539 (O_1539,N_49778,N_49837);
and UO_1540 (O_1540,N_49638,N_49948);
nand UO_1541 (O_1541,N_49555,N_49689);
nand UO_1542 (O_1542,N_49975,N_49802);
and UO_1543 (O_1543,N_49730,N_49769);
and UO_1544 (O_1544,N_49908,N_49547);
nand UO_1545 (O_1545,N_49651,N_49857);
nor UO_1546 (O_1546,N_49973,N_49932);
and UO_1547 (O_1547,N_49512,N_49818);
nor UO_1548 (O_1548,N_49944,N_49532);
or UO_1549 (O_1549,N_49966,N_49950);
and UO_1550 (O_1550,N_49936,N_49695);
nand UO_1551 (O_1551,N_49570,N_49785);
nor UO_1552 (O_1552,N_49847,N_49733);
or UO_1553 (O_1553,N_49972,N_49510);
or UO_1554 (O_1554,N_49525,N_49688);
and UO_1555 (O_1555,N_49949,N_49708);
xor UO_1556 (O_1556,N_49671,N_49733);
nand UO_1557 (O_1557,N_49726,N_49853);
or UO_1558 (O_1558,N_49578,N_49957);
and UO_1559 (O_1559,N_49691,N_49506);
nand UO_1560 (O_1560,N_49984,N_49613);
nor UO_1561 (O_1561,N_49786,N_49612);
and UO_1562 (O_1562,N_49676,N_49645);
and UO_1563 (O_1563,N_49819,N_49786);
nand UO_1564 (O_1564,N_49576,N_49673);
nor UO_1565 (O_1565,N_49962,N_49895);
and UO_1566 (O_1566,N_49569,N_49640);
nand UO_1567 (O_1567,N_49554,N_49544);
or UO_1568 (O_1568,N_49863,N_49764);
nand UO_1569 (O_1569,N_49837,N_49834);
and UO_1570 (O_1570,N_49833,N_49912);
or UO_1571 (O_1571,N_49680,N_49912);
xor UO_1572 (O_1572,N_49551,N_49729);
nor UO_1573 (O_1573,N_49559,N_49520);
nand UO_1574 (O_1574,N_49758,N_49870);
and UO_1575 (O_1575,N_49737,N_49674);
or UO_1576 (O_1576,N_49628,N_49999);
xnor UO_1577 (O_1577,N_49899,N_49762);
nand UO_1578 (O_1578,N_49917,N_49609);
nor UO_1579 (O_1579,N_49874,N_49865);
or UO_1580 (O_1580,N_49546,N_49500);
nor UO_1581 (O_1581,N_49608,N_49966);
nor UO_1582 (O_1582,N_49545,N_49568);
xor UO_1583 (O_1583,N_49810,N_49600);
or UO_1584 (O_1584,N_49657,N_49506);
and UO_1585 (O_1585,N_49778,N_49875);
or UO_1586 (O_1586,N_49560,N_49836);
and UO_1587 (O_1587,N_49761,N_49511);
nor UO_1588 (O_1588,N_49987,N_49616);
nor UO_1589 (O_1589,N_49792,N_49866);
nand UO_1590 (O_1590,N_49719,N_49830);
nand UO_1591 (O_1591,N_49540,N_49617);
or UO_1592 (O_1592,N_49624,N_49504);
and UO_1593 (O_1593,N_49650,N_49653);
xnor UO_1594 (O_1594,N_49617,N_49856);
nand UO_1595 (O_1595,N_49685,N_49944);
nand UO_1596 (O_1596,N_49819,N_49979);
xor UO_1597 (O_1597,N_49510,N_49963);
nand UO_1598 (O_1598,N_49620,N_49561);
and UO_1599 (O_1599,N_49949,N_49619);
and UO_1600 (O_1600,N_49750,N_49974);
nand UO_1601 (O_1601,N_49993,N_49897);
xnor UO_1602 (O_1602,N_49634,N_49649);
nand UO_1603 (O_1603,N_49820,N_49685);
xor UO_1604 (O_1604,N_49999,N_49570);
or UO_1605 (O_1605,N_49973,N_49824);
and UO_1606 (O_1606,N_49837,N_49606);
and UO_1607 (O_1607,N_49795,N_49778);
xor UO_1608 (O_1608,N_49632,N_49996);
or UO_1609 (O_1609,N_49940,N_49884);
nor UO_1610 (O_1610,N_49566,N_49830);
nand UO_1611 (O_1611,N_49917,N_49960);
xnor UO_1612 (O_1612,N_49624,N_49612);
xnor UO_1613 (O_1613,N_49518,N_49537);
nor UO_1614 (O_1614,N_49715,N_49620);
nand UO_1615 (O_1615,N_49767,N_49809);
nor UO_1616 (O_1616,N_49691,N_49947);
xor UO_1617 (O_1617,N_49667,N_49577);
nand UO_1618 (O_1618,N_49822,N_49579);
or UO_1619 (O_1619,N_49529,N_49993);
xor UO_1620 (O_1620,N_49656,N_49968);
nor UO_1621 (O_1621,N_49644,N_49913);
or UO_1622 (O_1622,N_49678,N_49918);
xor UO_1623 (O_1623,N_49983,N_49863);
or UO_1624 (O_1624,N_49914,N_49735);
or UO_1625 (O_1625,N_49722,N_49865);
and UO_1626 (O_1626,N_49867,N_49844);
xor UO_1627 (O_1627,N_49697,N_49949);
and UO_1628 (O_1628,N_49525,N_49529);
and UO_1629 (O_1629,N_49802,N_49790);
and UO_1630 (O_1630,N_49911,N_49613);
nand UO_1631 (O_1631,N_49957,N_49833);
nor UO_1632 (O_1632,N_49914,N_49547);
or UO_1633 (O_1633,N_49628,N_49549);
or UO_1634 (O_1634,N_49759,N_49943);
nor UO_1635 (O_1635,N_49684,N_49500);
nand UO_1636 (O_1636,N_49679,N_49592);
or UO_1637 (O_1637,N_49667,N_49617);
or UO_1638 (O_1638,N_49524,N_49624);
xor UO_1639 (O_1639,N_49719,N_49881);
and UO_1640 (O_1640,N_49748,N_49772);
nor UO_1641 (O_1641,N_49773,N_49643);
and UO_1642 (O_1642,N_49904,N_49822);
xnor UO_1643 (O_1643,N_49834,N_49622);
nand UO_1644 (O_1644,N_49634,N_49975);
nor UO_1645 (O_1645,N_49732,N_49567);
and UO_1646 (O_1646,N_49589,N_49811);
xor UO_1647 (O_1647,N_49715,N_49511);
nand UO_1648 (O_1648,N_49608,N_49678);
nand UO_1649 (O_1649,N_49714,N_49637);
nand UO_1650 (O_1650,N_49689,N_49806);
or UO_1651 (O_1651,N_49952,N_49665);
or UO_1652 (O_1652,N_49858,N_49579);
or UO_1653 (O_1653,N_49893,N_49742);
and UO_1654 (O_1654,N_49581,N_49901);
nor UO_1655 (O_1655,N_49652,N_49786);
xnor UO_1656 (O_1656,N_49576,N_49714);
or UO_1657 (O_1657,N_49626,N_49935);
or UO_1658 (O_1658,N_49908,N_49950);
xor UO_1659 (O_1659,N_49687,N_49703);
and UO_1660 (O_1660,N_49821,N_49527);
and UO_1661 (O_1661,N_49941,N_49713);
nand UO_1662 (O_1662,N_49574,N_49538);
nor UO_1663 (O_1663,N_49512,N_49792);
or UO_1664 (O_1664,N_49627,N_49702);
xor UO_1665 (O_1665,N_49560,N_49580);
nand UO_1666 (O_1666,N_49876,N_49553);
xnor UO_1667 (O_1667,N_49807,N_49891);
nor UO_1668 (O_1668,N_49585,N_49584);
or UO_1669 (O_1669,N_49592,N_49513);
or UO_1670 (O_1670,N_49580,N_49620);
and UO_1671 (O_1671,N_49800,N_49824);
xnor UO_1672 (O_1672,N_49651,N_49868);
xnor UO_1673 (O_1673,N_49735,N_49652);
xnor UO_1674 (O_1674,N_49809,N_49559);
and UO_1675 (O_1675,N_49890,N_49958);
or UO_1676 (O_1676,N_49764,N_49771);
nor UO_1677 (O_1677,N_49867,N_49521);
nor UO_1678 (O_1678,N_49814,N_49888);
nor UO_1679 (O_1679,N_49612,N_49577);
and UO_1680 (O_1680,N_49976,N_49844);
or UO_1681 (O_1681,N_49782,N_49767);
nor UO_1682 (O_1682,N_49819,N_49901);
or UO_1683 (O_1683,N_49931,N_49780);
xor UO_1684 (O_1684,N_49882,N_49866);
nor UO_1685 (O_1685,N_49758,N_49695);
or UO_1686 (O_1686,N_49536,N_49755);
nor UO_1687 (O_1687,N_49691,N_49990);
nand UO_1688 (O_1688,N_49915,N_49630);
xnor UO_1689 (O_1689,N_49578,N_49760);
nor UO_1690 (O_1690,N_49678,N_49752);
and UO_1691 (O_1691,N_49605,N_49677);
nor UO_1692 (O_1692,N_49506,N_49776);
and UO_1693 (O_1693,N_49561,N_49759);
and UO_1694 (O_1694,N_49571,N_49718);
or UO_1695 (O_1695,N_49853,N_49616);
xnor UO_1696 (O_1696,N_49852,N_49970);
xor UO_1697 (O_1697,N_49883,N_49701);
or UO_1698 (O_1698,N_49637,N_49903);
nand UO_1699 (O_1699,N_49835,N_49517);
nor UO_1700 (O_1700,N_49779,N_49776);
and UO_1701 (O_1701,N_49804,N_49836);
nand UO_1702 (O_1702,N_49945,N_49542);
xor UO_1703 (O_1703,N_49801,N_49662);
xor UO_1704 (O_1704,N_49587,N_49975);
nor UO_1705 (O_1705,N_49932,N_49819);
nand UO_1706 (O_1706,N_49655,N_49896);
or UO_1707 (O_1707,N_49681,N_49588);
and UO_1708 (O_1708,N_49987,N_49707);
nand UO_1709 (O_1709,N_49542,N_49990);
and UO_1710 (O_1710,N_49502,N_49887);
xnor UO_1711 (O_1711,N_49566,N_49661);
and UO_1712 (O_1712,N_49788,N_49954);
and UO_1713 (O_1713,N_49911,N_49783);
nor UO_1714 (O_1714,N_49825,N_49571);
or UO_1715 (O_1715,N_49756,N_49711);
and UO_1716 (O_1716,N_49628,N_49940);
or UO_1717 (O_1717,N_49851,N_49628);
and UO_1718 (O_1718,N_49640,N_49980);
and UO_1719 (O_1719,N_49574,N_49576);
nor UO_1720 (O_1720,N_49556,N_49992);
and UO_1721 (O_1721,N_49888,N_49524);
nor UO_1722 (O_1722,N_49670,N_49790);
nand UO_1723 (O_1723,N_49810,N_49856);
nand UO_1724 (O_1724,N_49720,N_49625);
xor UO_1725 (O_1725,N_49991,N_49922);
or UO_1726 (O_1726,N_49532,N_49742);
or UO_1727 (O_1727,N_49782,N_49554);
xnor UO_1728 (O_1728,N_49777,N_49913);
nand UO_1729 (O_1729,N_49806,N_49665);
nor UO_1730 (O_1730,N_49775,N_49571);
nor UO_1731 (O_1731,N_49618,N_49897);
xor UO_1732 (O_1732,N_49939,N_49848);
and UO_1733 (O_1733,N_49505,N_49870);
nand UO_1734 (O_1734,N_49679,N_49972);
or UO_1735 (O_1735,N_49915,N_49750);
nor UO_1736 (O_1736,N_49796,N_49973);
xor UO_1737 (O_1737,N_49641,N_49927);
nor UO_1738 (O_1738,N_49524,N_49677);
xor UO_1739 (O_1739,N_49909,N_49927);
or UO_1740 (O_1740,N_49504,N_49702);
nor UO_1741 (O_1741,N_49685,N_49965);
nor UO_1742 (O_1742,N_49752,N_49613);
nor UO_1743 (O_1743,N_49946,N_49515);
nor UO_1744 (O_1744,N_49513,N_49598);
or UO_1745 (O_1745,N_49565,N_49969);
xnor UO_1746 (O_1746,N_49945,N_49605);
xnor UO_1747 (O_1747,N_49661,N_49989);
and UO_1748 (O_1748,N_49683,N_49522);
and UO_1749 (O_1749,N_49603,N_49519);
nor UO_1750 (O_1750,N_49736,N_49728);
and UO_1751 (O_1751,N_49862,N_49831);
xnor UO_1752 (O_1752,N_49575,N_49747);
xnor UO_1753 (O_1753,N_49896,N_49550);
xnor UO_1754 (O_1754,N_49633,N_49631);
nor UO_1755 (O_1755,N_49784,N_49755);
or UO_1756 (O_1756,N_49585,N_49759);
or UO_1757 (O_1757,N_49768,N_49983);
nand UO_1758 (O_1758,N_49728,N_49762);
xor UO_1759 (O_1759,N_49618,N_49545);
xor UO_1760 (O_1760,N_49616,N_49586);
xnor UO_1761 (O_1761,N_49774,N_49996);
and UO_1762 (O_1762,N_49771,N_49815);
xor UO_1763 (O_1763,N_49573,N_49963);
or UO_1764 (O_1764,N_49516,N_49914);
and UO_1765 (O_1765,N_49694,N_49657);
xnor UO_1766 (O_1766,N_49535,N_49541);
nor UO_1767 (O_1767,N_49783,N_49789);
or UO_1768 (O_1768,N_49796,N_49742);
and UO_1769 (O_1769,N_49799,N_49624);
nand UO_1770 (O_1770,N_49833,N_49818);
nand UO_1771 (O_1771,N_49665,N_49848);
nor UO_1772 (O_1772,N_49592,N_49621);
nand UO_1773 (O_1773,N_49913,N_49926);
xor UO_1774 (O_1774,N_49635,N_49609);
nor UO_1775 (O_1775,N_49907,N_49617);
xnor UO_1776 (O_1776,N_49701,N_49929);
nand UO_1777 (O_1777,N_49819,N_49847);
and UO_1778 (O_1778,N_49745,N_49661);
xor UO_1779 (O_1779,N_49506,N_49575);
xor UO_1780 (O_1780,N_49707,N_49918);
and UO_1781 (O_1781,N_49560,N_49558);
nand UO_1782 (O_1782,N_49675,N_49687);
and UO_1783 (O_1783,N_49891,N_49852);
xnor UO_1784 (O_1784,N_49820,N_49918);
and UO_1785 (O_1785,N_49719,N_49714);
xor UO_1786 (O_1786,N_49788,N_49777);
xnor UO_1787 (O_1787,N_49560,N_49941);
nor UO_1788 (O_1788,N_49649,N_49836);
nand UO_1789 (O_1789,N_49731,N_49529);
xor UO_1790 (O_1790,N_49868,N_49672);
nor UO_1791 (O_1791,N_49609,N_49578);
or UO_1792 (O_1792,N_49713,N_49842);
or UO_1793 (O_1793,N_49694,N_49774);
xor UO_1794 (O_1794,N_49896,N_49707);
and UO_1795 (O_1795,N_49965,N_49550);
nor UO_1796 (O_1796,N_49645,N_49563);
and UO_1797 (O_1797,N_49991,N_49799);
and UO_1798 (O_1798,N_49699,N_49856);
nor UO_1799 (O_1799,N_49669,N_49522);
or UO_1800 (O_1800,N_49526,N_49962);
or UO_1801 (O_1801,N_49547,N_49500);
or UO_1802 (O_1802,N_49699,N_49583);
xnor UO_1803 (O_1803,N_49945,N_49505);
nor UO_1804 (O_1804,N_49537,N_49863);
or UO_1805 (O_1805,N_49879,N_49808);
nor UO_1806 (O_1806,N_49913,N_49878);
nor UO_1807 (O_1807,N_49573,N_49601);
nand UO_1808 (O_1808,N_49884,N_49595);
nor UO_1809 (O_1809,N_49553,N_49824);
xor UO_1810 (O_1810,N_49957,N_49530);
or UO_1811 (O_1811,N_49895,N_49849);
or UO_1812 (O_1812,N_49620,N_49628);
and UO_1813 (O_1813,N_49874,N_49654);
or UO_1814 (O_1814,N_49558,N_49773);
nand UO_1815 (O_1815,N_49987,N_49604);
xnor UO_1816 (O_1816,N_49748,N_49622);
nand UO_1817 (O_1817,N_49992,N_49664);
nand UO_1818 (O_1818,N_49930,N_49559);
or UO_1819 (O_1819,N_49969,N_49534);
nor UO_1820 (O_1820,N_49966,N_49660);
nor UO_1821 (O_1821,N_49889,N_49665);
nand UO_1822 (O_1822,N_49653,N_49854);
nand UO_1823 (O_1823,N_49530,N_49596);
nand UO_1824 (O_1824,N_49592,N_49771);
or UO_1825 (O_1825,N_49868,N_49705);
or UO_1826 (O_1826,N_49991,N_49508);
and UO_1827 (O_1827,N_49760,N_49873);
nand UO_1828 (O_1828,N_49533,N_49769);
nand UO_1829 (O_1829,N_49977,N_49973);
xor UO_1830 (O_1830,N_49517,N_49659);
or UO_1831 (O_1831,N_49842,N_49522);
xnor UO_1832 (O_1832,N_49863,N_49623);
or UO_1833 (O_1833,N_49748,N_49897);
nor UO_1834 (O_1834,N_49509,N_49636);
xor UO_1835 (O_1835,N_49539,N_49768);
or UO_1836 (O_1836,N_49866,N_49853);
or UO_1837 (O_1837,N_49810,N_49751);
nand UO_1838 (O_1838,N_49523,N_49598);
nor UO_1839 (O_1839,N_49650,N_49910);
and UO_1840 (O_1840,N_49635,N_49813);
or UO_1841 (O_1841,N_49947,N_49607);
nor UO_1842 (O_1842,N_49763,N_49935);
or UO_1843 (O_1843,N_49585,N_49628);
nor UO_1844 (O_1844,N_49719,N_49743);
xnor UO_1845 (O_1845,N_49716,N_49794);
nand UO_1846 (O_1846,N_49802,N_49635);
and UO_1847 (O_1847,N_49832,N_49657);
and UO_1848 (O_1848,N_49880,N_49617);
nor UO_1849 (O_1849,N_49540,N_49637);
nor UO_1850 (O_1850,N_49706,N_49921);
and UO_1851 (O_1851,N_49590,N_49898);
xnor UO_1852 (O_1852,N_49651,N_49505);
and UO_1853 (O_1853,N_49583,N_49871);
or UO_1854 (O_1854,N_49691,N_49707);
nand UO_1855 (O_1855,N_49943,N_49915);
nand UO_1856 (O_1856,N_49976,N_49569);
nor UO_1857 (O_1857,N_49656,N_49730);
nor UO_1858 (O_1858,N_49520,N_49501);
nor UO_1859 (O_1859,N_49895,N_49980);
or UO_1860 (O_1860,N_49527,N_49905);
or UO_1861 (O_1861,N_49609,N_49971);
nor UO_1862 (O_1862,N_49613,N_49868);
nand UO_1863 (O_1863,N_49838,N_49845);
or UO_1864 (O_1864,N_49569,N_49647);
or UO_1865 (O_1865,N_49941,N_49856);
nor UO_1866 (O_1866,N_49726,N_49756);
or UO_1867 (O_1867,N_49707,N_49627);
or UO_1868 (O_1868,N_49996,N_49888);
nand UO_1869 (O_1869,N_49511,N_49672);
nor UO_1870 (O_1870,N_49608,N_49548);
nor UO_1871 (O_1871,N_49664,N_49583);
or UO_1872 (O_1872,N_49929,N_49653);
and UO_1873 (O_1873,N_49572,N_49890);
or UO_1874 (O_1874,N_49892,N_49925);
xor UO_1875 (O_1875,N_49623,N_49542);
or UO_1876 (O_1876,N_49953,N_49728);
xor UO_1877 (O_1877,N_49546,N_49978);
or UO_1878 (O_1878,N_49790,N_49837);
and UO_1879 (O_1879,N_49949,N_49687);
nand UO_1880 (O_1880,N_49613,N_49944);
xnor UO_1881 (O_1881,N_49940,N_49960);
nor UO_1882 (O_1882,N_49856,N_49989);
xnor UO_1883 (O_1883,N_49742,N_49627);
or UO_1884 (O_1884,N_49905,N_49930);
nor UO_1885 (O_1885,N_49878,N_49902);
nor UO_1886 (O_1886,N_49885,N_49519);
xnor UO_1887 (O_1887,N_49820,N_49948);
or UO_1888 (O_1888,N_49561,N_49566);
nand UO_1889 (O_1889,N_49527,N_49511);
and UO_1890 (O_1890,N_49759,N_49754);
and UO_1891 (O_1891,N_49953,N_49672);
or UO_1892 (O_1892,N_49851,N_49573);
and UO_1893 (O_1893,N_49699,N_49986);
xnor UO_1894 (O_1894,N_49796,N_49779);
nand UO_1895 (O_1895,N_49800,N_49794);
and UO_1896 (O_1896,N_49848,N_49647);
nand UO_1897 (O_1897,N_49916,N_49899);
xnor UO_1898 (O_1898,N_49516,N_49569);
xor UO_1899 (O_1899,N_49817,N_49806);
xnor UO_1900 (O_1900,N_49587,N_49876);
and UO_1901 (O_1901,N_49979,N_49740);
xnor UO_1902 (O_1902,N_49976,N_49504);
or UO_1903 (O_1903,N_49620,N_49810);
and UO_1904 (O_1904,N_49937,N_49805);
or UO_1905 (O_1905,N_49885,N_49904);
xnor UO_1906 (O_1906,N_49753,N_49604);
xor UO_1907 (O_1907,N_49943,N_49609);
and UO_1908 (O_1908,N_49670,N_49532);
xor UO_1909 (O_1909,N_49825,N_49667);
and UO_1910 (O_1910,N_49958,N_49611);
xor UO_1911 (O_1911,N_49530,N_49986);
and UO_1912 (O_1912,N_49721,N_49678);
and UO_1913 (O_1913,N_49538,N_49546);
and UO_1914 (O_1914,N_49749,N_49808);
or UO_1915 (O_1915,N_49605,N_49665);
and UO_1916 (O_1916,N_49739,N_49900);
or UO_1917 (O_1917,N_49624,N_49989);
or UO_1918 (O_1918,N_49669,N_49695);
and UO_1919 (O_1919,N_49610,N_49660);
nor UO_1920 (O_1920,N_49572,N_49926);
nand UO_1921 (O_1921,N_49615,N_49526);
and UO_1922 (O_1922,N_49923,N_49993);
nor UO_1923 (O_1923,N_49984,N_49814);
and UO_1924 (O_1924,N_49776,N_49722);
or UO_1925 (O_1925,N_49736,N_49581);
nor UO_1926 (O_1926,N_49776,N_49593);
nand UO_1927 (O_1927,N_49576,N_49639);
xnor UO_1928 (O_1928,N_49788,N_49614);
xnor UO_1929 (O_1929,N_49686,N_49715);
nand UO_1930 (O_1930,N_49528,N_49702);
and UO_1931 (O_1931,N_49684,N_49833);
and UO_1932 (O_1932,N_49958,N_49995);
and UO_1933 (O_1933,N_49588,N_49952);
xor UO_1934 (O_1934,N_49857,N_49951);
nor UO_1935 (O_1935,N_49851,N_49781);
or UO_1936 (O_1936,N_49611,N_49555);
xnor UO_1937 (O_1937,N_49651,N_49971);
nor UO_1938 (O_1938,N_49558,N_49662);
nor UO_1939 (O_1939,N_49556,N_49691);
xnor UO_1940 (O_1940,N_49840,N_49874);
nor UO_1941 (O_1941,N_49848,N_49555);
xor UO_1942 (O_1942,N_49873,N_49998);
nor UO_1943 (O_1943,N_49945,N_49731);
or UO_1944 (O_1944,N_49799,N_49603);
or UO_1945 (O_1945,N_49693,N_49758);
nand UO_1946 (O_1946,N_49587,N_49914);
nor UO_1947 (O_1947,N_49523,N_49578);
nand UO_1948 (O_1948,N_49637,N_49828);
xnor UO_1949 (O_1949,N_49519,N_49541);
xnor UO_1950 (O_1950,N_49644,N_49607);
and UO_1951 (O_1951,N_49559,N_49823);
or UO_1952 (O_1952,N_49601,N_49785);
nand UO_1953 (O_1953,N_49670,N_49941);
xor UO_1954 (O_1954,N_49896,N_49582);
or UO_1955 (O_1955,N_49537,N_49519);
nor UO_1956 (O_1956,N_49845,N_49645);
and UO_1957 (O_1957,N_49864,N_49522);
nor UO_1958 (O_1958,N_49685,N_49952);
nand UO_1959 (O_1959,N_49976,N_49741);
and UO_1960 (O_1960,N_49891,N_49828);
or UO_1961 (O_1961,N_49522,N_49966);
xor UO_1962 (O_1962,N_49565,N_49943);
nor UO_1963 (O_1963,N_49731,N_49779);
nand UO_1964 (O_1964,N_49951,N_49958);
nor UO_1965 (O_1965,N_49852,N_49981);
and UO_1966 (O_1966,N_49722,N_49977);
nand UO_1967 (O_1967,N_49842,N_49675);
nor UO_1968 (O_1968,N_49508,N_49664);
xnor UO_1969 (O_1969,N_49728,N_49710);
or UO_1970 (O_1970,N_49887,N_49853);
xor UO_1971 (O_1971,N_49736,N_49955);
nor UO_1972 (O_1972,N_49683,N_49951);
and UO_1973 (O_1973,N_49634,N_49940);
nand UO_1974 (O_1974,N_49575,N_49868);
nor UO_1975 (O_1975,N_49915,N_49972);
nand UO_1976 (O_1976,N_49773,N_49747);
nand UO_1977 (O_1977,N_49914,N_49821);
nand UO_1978 (O_1978,N_49578,N_49847);
or UO_1979 (O_1979,N_49502,N_49584);
nand UO_1980 (O_1980,N_49701,N_49917);
nand UO_1981 (O_1981,N_49906,N_49656);
nor UO_1982 (O_1982,N_49939,N_49857);
xnor UO_1983 (O_1983,N_49546,N_49667);
nand UO_1984 (O_1984,N_49668,N_49547);
and UO_1985 (O_1985,N_49575,N_49832);
nand UO_1986 (O_1986,N_49640,N_49504);
and UO_1987 (O_1987,N_49638,N_49610);
and UO_1988 (O_1988,N_49868,N_49785);
xnor UO_1989 (O_1989,N_49703,N_49951);
xor UO_1990 (O_1990,N_49638,N_49970);
nor UO_1991 (O_1991,N_49930,N_49704);
nor UO_1992 (O_1992,N_49906,N_49981);
xnor UO_1993 (O_1993,N_49968,N_49781);
or UO_1994 (O_1994,N_49547,N_49957);
or UO_1995 (O_1995,N_49722,N_49981);
nand UO_1996 (O_1996,N_49591,N_49560);
or UO_1997 (O_1997,N_49558,N_49526);
nand UO_1998 (O_1998,N_49937,N_49514);
nand UO_1999 (O_1999,N_49795,N_49855);
nand UO_2000 (O_2000,N_49958,N_49618);
xnor UO_2001 (O_2001,N_49672,N_49924);
nand UO_2002 (O_2002,N_49966,N_49862);
xnor UO_2003 (O_2003,N_49952,N_49833);
or UO_2004 (O_2004,N_49704,N_49859);
and UO_2005 (O_2005,N_49708,N_49973);
or UO_2006 (O_2006,N_49566,N_49675);
xnor UO_2007 (O_2007,N_49810,N_49924);
or UO_2008 (O_2008,N_49981,N_49765);
nand UO_2009 (O_2009,N_49910,N_49825);
and UO_2010 (O_2010,N_49639,N_49773);
nor UO_2011 (O_2011,N_49825,N_49764);
or UO_2012 (O_2012,N_49949,N_49960);
xor UO_2013 (O_2013,N_49790,N_49546);
nand UO_2014 (O_2014,N_49507,N_49987);
or UO_2015 (O_2015,N_49746,N_49633);
xnor UO_2016 (O_2016,N_49525,N_49699);
xnor UO_2017 (O_2017,N_49656,N_49603);
nor UO_2018 (O_2018,N_49836,N_49508);
nand UO_2019 (O_2019,N_49880,N_49952);
nand UO_2020 (O_2020,N_49934,N_49619);
nor UO_2021 (O_2021,N_49920,N_49997);
and UO_2022 (O_2022,N_49769,N_49820);
or UO_2023 (O_2023,N_49895,N_49768);
or UO_2024 (O_2024,N_49528,N_49831);
nor UO_2025 (O_2025,N_49883,N_49528);
nand UO_2026 (O_2026,N_49868,N_49918);
nor UO_2027 (O_2027,N_49937,N_49791);
xor UO_2028 (O_2028,N_49847,N_49920);
xnor UO_2029 (O_2029,N_49845,N_49853);
or UO_2030 (O_2030,N_49677,N_49876);
nand UO_2031 (O_2031,N_49960,N_49873);
nor UO_2032 (O_2032,N_49978,N_49886);
nor UO_2033 (O_2033,N_49766,N_49673);
xnor UO_2034 (O_2034,N_49678,N_49892);
nand UO_2035 (O_2035,N_49861,N_49642);
and UO_2036 (O_2036,N_49604,N_49980);
and UO_2037 (O_2037,N_49910,N_49967);
nand UO_2038 (O_2038,N_49720,N_49670);
and UO_2039 (O_2039,N_49964,N_49729);
nor UO_2040 (O_2040,N_49646,N_49671);
and UO_2041 (O_2041,N_49699,N_49896);
or UO_2042 (O_2042,N_49619,N_49713);
or UO_2043 (O_2043,N_49528,N_49743);
or UO_2044 (O_2044,N_49796,N_49936);
nor UO_2045 (O_2045,N_49582,N_49913);
nor UO_2046 (O_2046,N_49682,N_49586);
xor UO_2047 (O_2047,N_49733,N_49928);
nor UO_2048 (O_2048,N_49580,N_49712);
nor UO_2049 (O_2049,N_49949,N_49834);
nand UO_2050 (O_2050,N_49834,N_49797);
or UO_2051 (O_2051,N_49729,N_49529);
and UO_2052 (O_2052,N_49543,N_49625);
and UO_2053 (O_2053,N_49695,N_49954);
nor UO_2054 (O_2054,N_49904,N_49662);
nor UO_2055 (O_2055,N_49594,N_49724);
nand UO_2056 (O_2056,N_49946,N_49929);
nor UO_2057 (O_2057,N_49816,N_49514);
nor UO_2058 (O_2058,N_49938,N_49693);
and UO_2059 (O_2059,N_49691,N_49902);
nor UO_2060 (O_2060,N_49622,N_49644);
and UO_2061 (O_2061,N_49505,N_49797);
or UO_2062 (O_2062,N_49751,N_49517);
nand UO_2063 (O_2063,N_49833,N_49723);
or UO_2064 (O_2064,N_49719,N_49786);
or UO_2065 (O_2065,N_49807,N_49827);
and UO_2066 (O_2066,N_49859,N_49956);
nand UO_2067 (O_2067,N_49592,N_49553);
and UO_2068 (O_2068,N_49864,N_49616);
xnor UO_2069 (O_2069,N_49924,N_49925);
nand UO_2070 (O_2070,N_49516,N_49932);
and UO_2071 (O_2071,N_49755,N_49579);
and UO_2072 (O_2072,N_49827,N_49937);
xor UO_2073 (O_2073,N_49867,N_49754);
xor UO_2074 (O_2074,N_49593,N_49838);
and UO_2075 (O_2075,N_49594,N_49733);
xnor UO_2076 (O_2076,N_49520,N_49592);
and UO_2077 (O_2077,N_49692,N_49935);
nand UO_2078 (O_2078,N_49510,N_49556);
nand UO_2079 (O_2079,N_49993,N_49732);
xnor UO_2080 (O_2080,N_49989,N_49705);
nor UO_2081 (O_2081,N_49772,N_49816);
or UO_2082 (O_2082,N_49707,N_49981);
and UO_2083 (O_2083,N_49592,N_49705);
nand UO_2084 (O_2084,N_49987,N_49637);
nor UO_2085 (O_2085,N_49624,N_49639);
or UO_2086 (O_2086,N_49843,N_49805);
or UO_2087 (O_2087,N_49575,N_49672);
xor UO_2088 (O_2088,N_49685,N_49700);
xnor UO_2089 (O_2089,N_49775,N_49610);
xor UO_2090 (O_2090,N_49554,N_49963);
or UO_2091 (O_2091,N_49606,N_49910);
nand UO_2092 (O_2092,N_49765,N_49651);
xnor UO_2093 (O_2093,N_49923,N_49626);
or UO_2094 (O_2094,N_49860,N_49979);
nor UO_2095 (O_2095,N_49996,N_49502);
xnor UO_2096 (O_2096,N_49888,N_49675);
and UO_2097 (O_2097,N_49686,N_49648);
nand UO_2098 (O_2098,N_49623,N_49857);
or UO_2099 (O_2099,N_49998,N_49943);
xnor UO_2100 (O_2100,N_49639,N_49700);
xnor UO_2101 (O_2101,N_49804,N_49781);
nor UO_2102 (O_2102,N_49878,N_49612);
xnor UO_2103 (O_2103,N_49932,N_49756);
and UO_2104 (O_2104,N_49691,N_49795);
nand UO_2105 (O_2105,N_49994,N_49607);
xnor UO_2106 (O_2106,N_49745,N_49858);
xnor UO_2107 (O_2107,N_49811,N_49951);
or UO_2108 (O_2108,N_49775,N_49527);
nand UO_2109 (O_2109,N_49605,N_49700);
and UO_2110 (O_2110,N_49756,N_49871);
nor UO_2111 (O_2111,N_49735,N_49570);
or UO_2112 (O_2112,N_49817,N_49788);
and UO_2113 (O_2113,N_49960,N_49895);
and UO_2114 (O_2114,N_49563,N_49982);
nand UO_2115 (O_2115,N_49776,N_49555);
nor UO_2116 (O_2116,N_49590,N_49978);
xnor UO_2117 (O_2117,N_49987,N_49858);
or UO_2118 (O_2118,N_49817,N_49758);
and UO_2119 (O_2119,N_49782,N_49726);
xor UO_2120 (O_2120,N_49820,N_49987);
xnor UO_2121 (O_2121,N_49572,N_49939);
or UO_2122 (O_2122,N_49681,N_49584);
xor UO_2123 (O_2123,N_49755,N_49720);
or UO_2124 (O_2124,N_49673,N_49948);
and UO_2125 (O_2125,N_49763,N_49977);
or UO_2126 (O_2126,N_49513,N_49643);
nand UO_2127 (O_2127,N_49595,N_49829);
and UO_2128 (O_2128,N_49974,N_49699);
or UO_2129 (O_2129,N_49714,N_49748);
nor UO_2130 (O_2130,N_49909,N_49952);
and UO_2131 (O_2131,N_49930,N_49712);
and UO_2132 (O_2132,N_49737,N_49812);
and UO_2133 (O_2133,N_49967,N_49775);
and UO_2134 (O_2134,N_49922,N_49940);
nand UO_2135 (O_2135,N_49836,N_49809);
xor UO_2136 (O_2136,N_49952,N_49521);
xor UO_2137 (O_2137,N_49933,N_49807);
or UO_2138 (O_2138,N_49619,N_49691);
nand UO_2139 (O_2139,N_49817,N_49690);
and UO_2140 (O_2140,N_49691,N_49748);
nand UO_2141 (O_2141,N_49529,N_49848);
and UO_2142 (O_2142,N_49901,N_49887);
or UO_2143 (O_2143,N_49729,N_49828);
nor UO_2144 (O_2144,N_49817,N_49722);
or UO_2145 (O_2145,N_49939,N_49663);
nand UO_2146 (O_2146,N_49624,N_49923);
xnor UO_2147 (O_2147,N_49887,N_49931);
nand UO_2148 (O_2148,N_49500,N_49663);
nor UO_2149 (O_2149,N_49864,N_49708);
nor UO_2150 (O_2150,N_49738,N_49718);
or UO_2151 (O_2151,N_49803,N_49795);
and UO_2152 (O_2152,N_49779,N_49903);
or UO_2153 (O_2153,N_49904,N_49818);
xnor UO_2154 (O_2154,N_49557,N_49580);
xnor UO_2155 (O_2155,N_49999,N_49783);
and UO_2156 (O_2156,N_49756,N_49744);
xnor UO_2157 (O_2157,N_49992,N_49808);
xnor UO_2158 (O_2158,N_49830,N_49512);
nand UO_2159 (O_2159,N_49549,N_49935);
or UO_2160 (O_2160,N_49719,N_49971);
nand UO_2161 (O_2161,N_49546,N_49535);
and UO_2162 (O_2162,N_49634,N_49517);
and UO_2163 (O_2163,N_49675,N_49665);
nand UO_2164 (O_2164,N_49501,N_49956);
xnor UO_2165 (O_2165,N_49573,N_49542);
xor UO_2166 (O_2166,N_49501,N_49663);
nand UO_2167 (O_2167,N_49938,N_49748);
or UO_2168 (O_2168,N_49806,N_49989);
or UO_2169 (O_2169,N_49919,N_49700);
xnor UO_2170 (O_2170,N_49923,N_49948);
nor UO_2171 (O_2171,N_49996,N_49576);
nand UO_2172 (O_2172,N_49663,N_49630);
nor UO_2173 (O_2173,N_49988,N_49697);
and UO_2174 (O_2174,N_49687,N_49751);
xor UO_2175 (O_2175,N_49969,N_49958);
nor UO_2176 (O_2176,N_49659,N_49811);
nor UO_2177 (O_2177,N_49511,N_49799);
xnor UO_2178 (O_2178,N_49737,N_49604);
xnor UO_2179 (O_2179,N_49937,N_49982);
and UO_2180 (O_2180,N_49668,N_49893);
xor UO_2181 (O_2181,N_49623,N_49535);
xnor UO_2182 (O_2182,N_49773,N_49978);
nand UO_2183 (O_2183,N_49924,N_49962);
nor UO_2184 (O_2184,N_49650,N_49601);
or UO_2185 (O_2185,N_49991,N_49593);
and UO_2186 (O_2186,N_49838,N_49751);
or UO_2187 (O_2187,N_49868,N_49730);
nor UO_2188 (O_2188,N_49676,N_49815);
xnor UO_2189 (O_2189,N_49710,N_49966);
nand UO_2190 (O_2190,N_49582,N_49912);
or UO_2191 (O_2191,N_49731,N_49668);
nor UO_2192 (O_2192,N_49716,N_49627);
nand UO_2193 (O_2193,N_49712,N_49563);
nand UO_2194 (O_2194,N_49768,N_49522);
nand UO_2195 (O_2195,N_49641,N_49686);
xnor UO_2196 (O_2196,N_49946,N_49805);
xnor UO_2197 (O_2197,N_49988,N_49921);
nand UO_2198 (O_2198,N_49751,N_49889);
or UO_2199 (O_2199,N_49580,N_49972);
or UO_2200 (O_2200,N_49662,N_49626);
and UO_2201 (O_2201,N_49564,N_49968);
nor UO_2202 (O_2202,N_49503,N_49645);
and UO_2203 (O_2203,N_49854,N_49728);
nor UO_2204 (O_2204,N_49533,N_49859);
nor UO_2205 (O_2205,N_49574,N_49777);
or UO_2206 (O_2206,N_49959,N_49933);
xor UO_2207 (O_2207,N_49883,N_49755);
nor UO_2208 (O_2208,N_49603,N_49823);
xnor UO_2209 (O_2209,N_49873,N_49511);
nand UO_2210 (O_2210,N_49688,N_49612);
nor UO_2211 (O_2211,N_49765,N_49544);
or UO_2212 (O_2212,N_49680,N_49813);
nand UO_2213 (O_2213,N_49697,N_49575);
nand UO_2214 (O_2214,N_49580,N_49683);
xor UO_2215 (O_2215,N_49890,N_49673);
nand UO_2216 (O_2216,N_49833,N_49923);
and UO_2217 (O_2217,N_49914,N_49709);
nor UO_2218 (O_2218,N_49956,N_49542);
and UO_2219 (O_2219,N_49734,N_49803);
xnor UO_2220 (O_2220,N_49572,N_49897);
xnor UO_2221 (O_2221,N_49869,N_49824);
nor UO_2222 (O_2222,N_49783,N_49784);
and UO_2223 (O_2223,N_49632,N_49993);
or UO_2224 (O_2224,N_49715,N_49602);
and UO_2225 (O_2225,N_49750,N_49651);
xnor UO_2226 (O_2226,N_49829,N_49677);
or UO_2227 (O_2227,N_49577,N_49555);
xnor UO_2228 (O_2228,N_49591,N_49769);
nand UO_2229 (O_2229,N_49885,N_49504);
nand UO_2230 (O_2230,N_49697,N_49928);
or UO_2231 (O_2231,N_49913,N_49984);
or UO_2232 (O_2232,N_49693,N_49551);
and UO_2233 (O_2233,N_49710,N_49578);
nor UO_2234 (O_2234,N_49927,N_49816);
nor UO_2235 (O_2235,N_49788,N_49904);
nor UO_2236 (O_2236,N_49679,N_49726);
xor UO_2237 (O_2237,N_49822,N_49729);
or UO_2238 (O_2238,N_49637,N_49768);
xor UO_2239 (O_2239,N_49522,N_49914);
or UO_2240 (O_2240,N_49766,N_49971);
xor UO_2241 (O_2241,N_49980,N_49633);
nor UO_2242 (O_2242,N_49924,N_49639);
or UO_2243 (O_2243,N_49897,N_49692);
or UO_2244 (O_2244,N_49519,N_49814);
or UO_2245 (O_2245,N_49780,N_49773);
or UO_2246 (O_2246,N_49527,N_49781);
nor UO_2247 (O_2247,N_49890,N_49803);
nand UO_2248 (O_2248,N_49555,N_49652);
and UO_2249 (O_2249,N_49779,N_49644);
and UO_2250 (O_2250,N_49749,N_49939);
or UO_2251 (O_2251,N_49695,N_49730);
or UO_2252 (O_2252,N_49857,N_49914);
and UO_2253 (O_2253,N_49559,N_49952);
and UO_2254 (O_2254,N_49571,N_49643);
nor UO_2255 (O_2255,N_49999,N_49784);
xnor UO_2256 (O_2256,N_49571,N_49881);
nand UO_2257 (O_2257,N_49832,N_49870);
xor UO_2258 (O_2258,N_49731,N_49972);
and UO_2259 (O_2259,N_49561,N_49503);
nand UO_2260 (O_2260,N_49567,N_49920);
xor UO_2261 (O_2261,N_49703,N_49967);
and UO_2262 (O_2262,N_49555,N_49912);
nand UO_2263 (O_2263,N_49675,N_49627);
xor UO_2264 (O_2264,N_49617,N_49890);
or UO_2265 (O_2265,N_49955,N_49577);
xnor UO_2266 (O_2266,N_49918,N_49960);
and UO_2267 (O_2267,N_49522,N_49754);
and UO_2268 (O_2268,N_49838,N_49816);
and UO_2269 (O_2269,N_49512,N_49937);
and UO_2270 (O_2270,N_49893,N_49602);
or UO_2271 (O_2271,N_49542,N_49991);
or UO_2272 (O_2272,N_49604,N_49684);
and UO_2273 (O_2273,N_49583,N_49650);
nand UO_2274 (O_2274,N_49748,N_49593);
and UO_2275 (O_2275,N_49885,N_49548);
xor UO_2276 (O_2276,N_49659,N_49602);
xnor UO_2277 (O_2277,N_49580,N_49853);
xor UO_2278 (O_2278,N_49524,N_49776);
xnor UO_2279 (O_2279,N_49837,N_49602);
xnor UO_2280 (O_2280,N_49656,N_49650);
xor UO_2281 (O_2281,N_49649,N_49619);
nand UO_2282 (O_2282,N_49795,N_49966);
xnor UO_2283 (O_2283,N_49850,N_49642);
or UO_2284 (O_2284,N_49872,N_49677);
xor UO_2285 (O_2285,N_49697,N_49512);
xor UO_2286 (O_2286,N_49534,N_49627);
nor UO_2287 (O_2287,N_49739,N_49572);
nor UO_2288 (O_2288,N_49914,N_49742);
nand UO_2289 (O_2289,N_49790,N_49553);
nor UO_2290 (O_2290,N_49853,N_49576);
nand UO_2291 (O_2291,N_49531,N_49989);
and UO_2292 (O_2292,N_49877,N_49878);
or UO_2293 (O_2293,N_49755,N_49677);
nor UO_2294 (O_2294,N_49959,N_49804);
nand UO_2295 (O_2295,N_49736,N_49748);
or UO_2296 (O_2296,N_49501,N_49737);
and UO_2297 (O_2297,N_49973,N_49574);
and UO_2298 (O_2298,N_49632,N_49566);
nand UO_2299 (O_2299,N_49814,N_49509);
nor UO_2300 (O_2300,N_49636,N_49576);
nor UO_2301 (O_2301,N_49675,N_49957);
nor UO_2302 (O_2302,N_49728,N_49612);
and UO_2303 (O_2303,N_49680,N_49681);
or UO_2304 (O_2304,N_49503,N_49509);
nand UO_2305 (O_2305,N_49772,N_49765);
xnor UO_2306 (O_2306,N_49572,N_49726);
nand UO_2307 (O_2307,N_49959,N_49801);
or UO_2308 (O_2308,N_49609,N_49994);
nor UO_2309 (O_2309,N_49944,N_49724);
and UO_2310 (O_2310,N_49640,N_49952);
nor UO_2311 (O_2311,N_49959,N_49787);
xnor UO_2312 (O_2312,N_49942,N_49963);
nand UO_2313 (O_2313,N_49591,N_49836);
or UO_2314 (O_2314,N_49618,N_49533);
nor UO_2315 (O_2315,N_49507,N_49830);
nor UO_2316 (O_2316,N_49649,N_49603);
nand UO_2317 (O_2317,N_49684,N_49687);
nand UO_2318 (O_2318,N_49779,N_49873);
and UO_2319 (O_2319,N_49509,N_49689);
or UO_2320 (O_2320,N_49914,N_49511);
nor UO_2321 (O_2321,N_49938,N_49523);
xnor UO_2322 (O_2322,N_49663,N_49527);
nor UO_2323 (O_2323,N_49870,N_49874);
or UO_2324 (O_2324,N_49799,N_49638);
or UO_2325 (O_2325,N_49823,N_49753);
nand UO_2326 (O_2326,N_49645,N_49505);
and UO_2327 (O_2327,N_49923,N_49943);
nand UO_2328 (O_2328,N_49963,N_49713);
and UO_2329 (O_2329,N_49886,N_49946);
nor UO_2330 (O_2330,N_49907,N_49870);
xor UO_2331 (O_2331,N_49872,N_49621);
xor UO_2332 (O_2332,N_49700,N_49805);
or UO_2333 (O_2333,N_49830,N_49755);
or UO_2334 (O_2334,N_49526,N_49974);
or UO_2335 (O_2335,N_49873,N_49545);
and UO_2336 (O_2336,N_49684,N_49896);
xor UO_2337 (O_2337,N_49638,N_49829);
and UO_2338 (O_2338,N_49886,N_49702);
or UO_2339 (O_2339,N_49870,N_49562);
xnor UO_2340 (O_2340,N_49865,N_49539);
or UO_2341 (O_2341,N_49772,N_49913);
xor UO_2342 (O_2342,N_49938,N_49736);
nor UO_2343 (O_2343,N_49878,N_49720);
nand UO_2344 (O_2344,N_49935,N_49671);
and UO_2345 (O_2345,N_49917,N_49817);
xnor UO_2346 (O_2346,N_49897,N_49519);
xnor UO_2347 (O_2347,N_49939,N_49731);
and UO_2348 (O_2348,N_49544,N_49740);
xor UO_2349 (O_2349,N_49676,N_49794);
nor UO_2350 (O_2350,N_49625,N_49863);
and UO_2351 (O_2351,N_49860,N_49683);
or UO_2352 (O_2352,N_49929,N_49756);
nor UO_2353 (O_2353,N_49983,N_49592);
nor UO_2354 (O_2354,N_49602,N_49911);
nand UO_2355 (O_2355,N_49760,N_49623);
nand UO_2356 (O_2356,N_49736,N_49568);
nand UO_2357 (O_2357,N_49703,N_49553);
and UO_2358 (O_2358,N_49810,N_49669);
xnor UO_2359 (O_2359,N_49820,N_49617);
nor UO_2360 (O_2360,N_49513,N_49560);
nand UO_2361 (O_2361,N_49735,N_49714);
and UO_2362 (O_2362,N_49638,N_49844);
nor UO_2363 (O_2363,N_49922,N_49877);
xor UO_2364 (O_2364,N_49531,N_49555);
or UO_2365 (O_2365,N_49745,N_49631);
xor UO_2366 (O_2366,N_49572,N_49649);
xor UO_2367 (O_2367,N_49804,N_49524);
nand UO_2368 (O_2368,N_49604,N_49895);
and UO_2369 (O_2369,N_49846,N_49828);
or UO_2370 (O_2370,N_49834,N_49887);
and UO_2371 (O_2371,N_49799,N_49964);
or UO_2372 (O_2372,N_49759,N_49829);
nand UO_2373 (O_2373,N_49765,N_49947);
xor UO_2374 (O_2374,N_49749,N_49625);
or UO_2375 (O_2375,N_49859,N_49744);
nand UO_2376 (O_2376,N_49973,N_49686);
or UO_2377 (O_2377,N_49570,N_49783);
xor UO_2378 (O_2378,N_49644,N_49558);
nand UO_2379 (O_2379,N_49542,N_49835);
xnor UO_2380 (O_2380,N_49746,N_49849);
or UO_2381 (O_2381,N_49793,N_49523);
and UO_2382 (O_2382,N_49865,N_49723);
and UO_2383 (O_2383,N_49625,N_49894);
xnor UO_2384 (O_2384,N_49722,N_49883);
nand UO_2385 (O_2385,N_49969,N_49756);
nand UO_2386 (O_2386,N_49763,N_49927);
or UO_2387 (O_2387,N_49635,N_49966);
or UO_2388 (O_2388,N_49787,N_49593);
nor UO_2389 (O_2389,N_49799,N_49749);
and UO_2390 (O_2390,N_49685,N_49817);
xnor UO_2391 (O_2391,N_49529,N_49641);
or UO_2392 (O_2392,N_49661,N_49679);
or UO_2393 (O_2393,N_49573,N_49978);
xor UO_2394 (O_2394,N_49785,N_49648);
or UO_2395 (O_2395,N_49536,N_49853);
xnor UO_2396 (O_2396,N_49841,N_49523);
and UO_2397 (O_2397,N_49685,N_49862);
or UO_2398 (O_2398,N_49513,N_49824);
nand UO_2399 (O_2399,N_49540,N_49846);
and UO_2400 (O_2400,N_49534,N_49668);
xnor UO_2401 (O_2401,N_49878,N_49752);
nand UO_2402 (O_2402,N_49713,N_49693);
and UO_2403 (O_2403,N_49641,N_49503);
nand UO_2404 (O_2404,N_49719,N_49964);
nand UO_2405 (O_2405,N_49943,N_49904);
or UO_2406 (O_2406,N_49682,N_49595);
nand UO_2407 (O_2407,N_49839,N_49836);
or UO_2408 (O_2408,N_49938,N_49568);
and UO_2409 (O_2409,N_49988,N_49520);
nor UO_2410 (O_2410,N_49883,N_49632);
nor UO_2411 (O_2411,N_49921,N_49900);
nand UO_2412 (O_2412,N_49714,N_49572);
nand UO_2413 (O_2413,N_49981,N_49684);
nor UO_2414 (O_2414,N_49837,N_49599);
xnor UO_2415 (O_2415,N_49777,N_49559);
xnor UO_2416 (O_2416,N_49610,N_49634);
xor UO_2417 (O_2417,N_49704,N_49934);
nand UO_2418 (O_2418,N_49511,N_49502);
and UO_2419 (O_2419,N_49507,N_49931);
or UO_2420 (O_2420,N_49794,N_49936);
and UO_2421 (O_2421,N_49747,N_49935);
nor UO_2422 (O_2422,N_49611,N_49533);
nand UO_2423 (O_2423,N_49905,N_49857);
or UO_2424 (O_2424,N_49592,N_49638);
and UO_2425 (O_2425,N_49543,N_49782);
xor UO_2426 (O_2426,N_49883,N_49842);
nand UO_2427 (O_2427,N_49589,N_49543);
and UO_2428 (O_2428,N_49919,N_49966);
xor UO_2429 (O_2429,N_49760,N_49712);
nand UO_2430 (O_2430,N_49942,N_49600);
or UO_2431 (O_2431,N_49917,N_49985);
nand UO_2432 (O_2432,N_49834,N_49824);
nand UO_2433 (O_2433,N_49723,N_49983);
or UO_2434 (O_2434,N_49534,N_49944);
xor UO_2435 (O_2435,N_49935,N_49714);
xor UO_2436 (O_2436,N_49695,N_49798);
nor UO_2437 (O_2437,N_49936,N_49716);
or UO_2438 (O_2438,N_49925,N_49571);
and UO_2439 (O_2439,N_49913,N_49681);
nor UO_2440 (O_2440,N_49520,N_49907);
xor UO_2441 (O_2441,N_49978,N_49671);
xnor UO_2442 (O_2442,N_49600,N_49532);
xor UO_2443 (O_2443,N_49944,N_49666);
xor UO_2444 (O_2444,N_49525,N_49718);
or UO_2445 (O_2445,N_49680,N_49956);
nor UO_2446 (O_2446,N_49988,N_49904);
nor UO_2447 (O_2447,N_49587,N_49996);
and UO_2448 (O_2448,N_49967,N_49714);
nor UO_2449 (O_2449,N_49934,N_49921);
nand UO_2450 (O_2450,N_49520,N_49610);
nor UO_2451 (O_2451,N_49978,N_49600);
and UO_2452 (O_2452,N_49979,N_49857);
and UO_2453 (O_2453,N_49908,N_49698);
xor UO_2454 (O_2454,N_49937,N_49902);
or UO_2455 (O_2455,N_49699,N_49862);
and UO_2456 (O_2456,N_49500,N_49849);
nand UO_2457 (O_2457,N_49859,N_49769);
xnor UO_2458 (O_2458,N_49609,N_49626);
and UO_2459 (O_2459,N_49979,N_49841);
or UO_2460 (O_2460,N_49729,N_49904);
and UO_2461 (O_2461,N_49987,N_49722);
or UO_2462 (O_2462,N_49788,N_49570);
nand UO_2463 (O_2463,N_49736,N_49633);
or UO_2464 (O_2464,N_49630,N_49515);
nor UO_2465 (O_2465,N_49543,N_49871);
or UO_2466 (O_2466,N_49555,N_49738);
nand UO_2467 (O_2467,N_49894,N_49637);
xor UO_2468 (O_2468,N_49716,N_49616);
or UO_2469 (O_2469,N_49816,N_49635);
nor UO_2470 (O_2470,N_49553,N_49814);
xor UO_2471 (O_2471,N_49603,N_49752);
or UO_2472 (O_2472,N_49680,N_49739);
xor UO_2473 (O_2473,N_49806,N_49884);
or UO_2474 (O_2474,N_49580,N_49830);
xor UO_2475 (O_2475,N_49966,N_49604);
nor UO_2476 (O_2476,N_49645,N_49872);
nor UO_2477 (O_2477,N_49729,N_49627);
nand UO_2478 (O_2478,N_49725,N_49690);
nand UO_2479 (O_2479,N_49889,N_49583);
nor UO_2480 (O_2480,N_49780,N_49961);
nor UO_2481 (O_2481,N_49528,N_49690);
nor UO_2482 (O_2482,N_49628,N_49706);
or UO_2483 (O_2483,N_49570,N_49530);
xor UO_2484 (O_2484,N_49558,N_49565);
or UO_2485 (O_2485,N_49918,N_49566);
or UO_2486 (O_2486,N_49808,N_49822);
xor UO_2487 (O_2487,N_49972,N_49853);
or UO_2488 (O_2488,N_49929,N_49893);
nand UO_2489 (O_2489,N_49504,N_49549);
nor UO_2490 (O_2490,N_49865,N_49633);
and UO_2491 (O_2491,N_49739,N_49512);
nor UO_2492 (O_2492,N_49923,N_49895);
and UO_2493 (O_2493,N_49785,N_49729);
xnor UO_2494 (O_2494,N_49547,N_49958);
xor UO_2495 (O_2495,N_49796,N_49507);
nand UO_2496 (O_2496,N_49729,N_49534);
or UO_2497 (O_2497,N_49759,N_49650);
nor UO_2498 (O_2498,N_49988,N_49909);
nor UO_2499 (O_2499,N_49646,N_49827);
and UO_2500 (O_2500,N_49896,N_49590);
nand UO_2501 (O_2501,N_49929,N_49683);
xor UO_2502 (O_2502,N_49692,N_49609);
nor UO_2503 (O_2503,N_49676,N_49732);
nor UO_2504 (O_2504,N_49963,N_49676);
xnor UO_2505 (O_2505,N_49817,N_49526);
or UO_2506 (O_2506,N_49979,N_49812);
xor UO_2507 (O_2507,N_49666,N_49955);
nor UO_2508 (O_2508,N_49801,N_49865);
and UO_2509 (O_2509,N_49599,N_49582);
and UO_2510 (O_2510,N_49587,N_49547);
nor UO_2511 (O_2511,N_49967,N_49508);
nor UO_2512 (O_2512,N_49993,N_49966);
and UO_2513 (O_2513,N_49658,N_49649);
nand UO_2514 (O_2514,N_49517,N_49691);
nand UO_2515 (O_2515,N_49851,N_49996);
and UO_2516 (O_2516,N_49553,N_49999);
nand UO_2517 (O_2517,N_49649,N_49817);
and UO_2518 (O_2518,N_49632,N_49730);
or UO_2519 (O_2519,N_49974,N_49990);
or UO_2520 (O_2520,N_49522,N_49564);
nand UO_2521 (O_2521,N_49653,N_49988);
and UO_2522 (O_2522,N_49560,N_49868);
or UO_2523 (O_2523,N_49526,N_49985);
xnor UO_2524 (O_2524,N_49577,N_49868);
nand UO_2525 (O_2525,N_49723,N_49612);
xnor UO_2526 (O_2526,N_49868,N_49869);
xor UO_2527 (O_2527,N_49748,N_49892);
nor UO_2528 (O_2528,N_49665,N_49825);
xor UO_2529 (O_2529,N_49831,N_49583);
and UO_2530 (O_2530,N_49917,N_49905);
nor UO_2531 (O_2531,N_49654,N_49972);
nor UO_2532 (O_2532,N_49580,N_49776);
and UO_2533 (O_2533,N_49987,N_49636);
or UO_2534 (O_2534,N_49970,N_49926);
nand UO_2535 (O_2535,N_49547,N_49925);
nor UO_2536 (O_2536,N_49527,N_49646);
xor UO_2537 (O_2537,N_49714,N_49631);
or UO_2538 (O_2538,N_49747,N_49842);
nand UO_2539 (O_2539,N_49865,N_49747);
or UO_2540 (O_2540,N_49980,N_49931);
nor UO_2541 (O_2541,N_49599,N_49940);
and UO_2542 (O_2542,N_49536,N_49513);
and UO_2543 (O_2543,N_49772,N_49867);
or UO_2544 (O_2544,N_49724,N_49954);
xor UO_2545 (O_2545,N_49618,N_49960);
xor UO_2546 (O_2546,N_49616,N_49643);
xnor UO_2547 (O_2547,N_49749,N_49683);
and UO_2548 (O_2548,N_49644,N_49531);
nand UO_2549 (O_2549,N_49894,N_49501);
nand UO_2550 (O_2550,N_49978,N_49727);
xnor UO_2551 (O_2551,N_49869,N_49526);
nand UO_2552 (O_2552,N_49523,N_49545);
or UO_2553 (O_2553,N_49913,N_49983);
nor UO_2554 (O_2554,N_49641,N_49856);
or UO_2555 (O_2555,N_49651,N_49937);
nor UO_2556 (O_2556,N_49972,N_49778);
or UO_2557 (O_2557,N_49894,N_49912);
xor UO_2558 (O_2558,N_49725,N_49817);
xnor UO_2559 (O_2559,N_49754,N_49877);
nor UO_2560 (O_2560,N_49957,N_49867);
nor UO_2561 (O_2561,N_49751,N_49964);
xor UO_2562 (O_2562,N_49744,N_49640);
nor UO_2563 (O_2563,N_49704,N_49992);
and UO_2564 (O_2564,N_49928,N_49799);
nand UO_2565 (O_2565,N_49952,N_49903);
or UO_2566 (O_2566,N_49985,N_49738);
nand UO_2567 (O_2567,N_49615,N_49829);
or UO_2568 (O_2568,N_49764,N_49748);
and UO_2569 (O_2569,N_49965,N_49616);
and UO_2570 (O_2570,N_49640,N_49847);
xnor UO_2571 (O_2571,N_49573,N_49742);
and UO_2572 (O_2572,N_49846,N_49983);
xnor UO_2573 (O_2573,N_49571,N_49968);
xnor UO_2574 (O_2574,N_49594,N_49583);
nand UO_2575 (O_2575,N_49937,N_49977);
nor UO_2576 (O_2576,N_49715,N_49633);
and UO_2577 (O_2577,N_49835,N_49837);
nor UO_2578 (O_2578,N_49852,N_49920);
xor UO_2579 (O_2579,N_49740,N_49774);
xor UO_2580 (O_2580,N_49946,N_49640);
nand UO_2581 (O_2581,N_49973,N_49558);
nand UO_2582 (O_2582,N_49773,N_49525);
and UO_2583 (O_2583,N_49583,N_49514);
and UO_2584 (O_2584,N_49915,N_49524);
or UO_2585 (O_2585,N_49557,N_49572);
or UO_2586 (O_2586,N_49926,N_49834);
xor UO_2587 (O_2587,N_49849,N_49814);
nand UO_2588 (O_2588,N_49951,N_49960);
nand UO_2589 (O_2589,N_49716,N_49643);
nand UO_2590 (O_2590,N_49677,N_49795);
nand UO_2591 (O_2591,N_49987,N_49543);
and UO_2592 (O_2592,N_49957,N_49592);
and UO_2593 (O_2593,N_49557,N_49702);
or UO_2594 (O_2594,N_49655,N_49733);
and UO_2595 (O_2595,N_49815,N_49855);
xnor UO_2596 (O_2596,N_49608,N_49685);
and UO_2597 (O_2597,N_49529,N_49994);
nand UO_2598 (O_2598,N_49559,N_49749);
nand UO_2599 (O_2599,N_49731,N_49753);
or UO_2600 (O_2600,N_49633,N_49659);
nor UO_2601 (O_2601,N_49836,N_49935);
nand UO_2602 (O_2602,N_49689,N_49866);
nand UO_2603 (O_2603,N_49836,N_49889);
or UO_2604 (O_2604,N_49612,N_49938);
nor UO_2605 (O_2605,N_49561,N_49575);
xor UO_2606 (O_2606,N_49774,N_49696);
nor UO_2607 (O_2607,N_49897,N_49826);
or UO_2608 (O_2608,N_49723,N_49534);
and UO_2609 (O_2609,N_49541,N_49556);
nand UO_2610 (O_2610,N_49659,N_49696);
and UO_2611 (O_2611,N_49566,N_49668);
xor UO_2612 (O_2612,N_49516,N_49577);
nor UO_2613 (O_2613,N_49983,N_49729);
nand UO_2614 (O_2614,N_49513,N_49557);
xnor UO_2615 (O_2615,N_49620,N_49879);
nor UO_2616 (O_2616,N_49899,N_49596);
nand UO_2617 (O_2617,N_49866,N_49928);
nand UO_2618 (O_2618,N_49576,N_49879);
xnor UO_2619 (O_2619,N_49783,N_49857);
and UO_2620 (O_2620,N_49984,N_49690);
nand UO_2621 (O_2621,N_49963,N_49911);
nand UO_2622 (O_2622,N_49766,N_49600);
xor UO_2623 (O_2623,N_49967,N_49551);
or UO_2624 (O_2624,N_49731,N_49785);
xnor UO_2625 (O_2625,N_49681,N_49834);
nor UO_2626 (O_2626,N_49632,N_49870);
or UO_2627 (O_2627,N_49790,N_49736);
nand UO_2628 (O_2628,N_49564,N_49544);
and UO_2629 (O_2629,N_49850,N_49727);
or UO_2630 (O_2630,N_49642,N_49953);
or UO_2631 (O_2631,N_49682,N_49857);
and UO_2632 (O_2632,N_49911,N_49686);
and UO_2633 (O_2633,N_49918,N_49690);
xnor UO_2634 (O_2634,N_49520,N_49602);
nand UO_2635 (O_2635,N_49985,N_49657);
and UO_2636 (O_2636,N_49612,N_49648);
or UO_2637 (O_2637,N_49686,N_49813);
and UO_2638 (O_2638,N_49912,N_49721);
nand UO_2639 (O_2639,N_49745,N_49754);
or UO_2640 (O_2640,N_49899,N_49572);
or UO_2641 (O_2641,N_49647,N_49762);
nand UO_2642 (O_2642,N_49632,N_49607);
nand UO_2643 (O_2643,N_49548,N_49661);
and UO_2644 (O_2644,N_49754,N_49661);
nand UO_2645 (O_2645,N_49814,N_49852);
and UO_2646 (O_2646,N_49521,N_49708);
and UO_2647 (O_2647,N_49623,N_49533);
and UO_2648 (O_2648,N_49641,N_49745);
or UO_2649 (O_2649,N_49684,N_49793);
xnor UO_2650 (O_2650,N_49634,N_49857);
and UO_2651 (O_2651,N_49659,N_49779);
and UO_2652 (O_2652,N_49806,N_49628);
and UO_2653 (O_2653,N_49877,N_49821);
nand UO_2654 (O_2654,N_49988,N_49826);
and UO_2655 (O_2655,N_49745,N_49519);
xnor UO_2656 (O_2656,N_49821,N_49747);
nor UO_2657 (O_2657,N_49803,N_49847);
and UO_2658 (O_2658,N_49510,N_49700);
nand UO_2659 (O_2659,N_49673,N_49976);
and UO_2660 (O_2660,N_49550,N_49691);
and UO_2661 (O_2661,N_49517,N_49994);
or UO_2662 (O_2662,N_49705,N_49845);
nor UO_2663 (O_2663,N_49663,N_49658);
nand UO_2664 (O_2664,N_49911,N_49875);
xnor UO_2665 (O_2665,N_49580,N_49657);
nand UO_2666 (O_2666,N_49798,N_49952);
nor UO_2667 (O_2667,N_49884,N_49629);
and UO_2668 (O_2668,N_49786,N_49970);
and UO_2669 (O_2669,N_49843,N_49563);
or UO_2670 (O_2670,N_49704,N_49511);
xor UO_2671 (O_2671,N_49857,N_49523);
nand UO_2672 (O_2672,N_49832,N_49624);
xor UO_2673 (O_2673,N_49912,N_49620);
and UO_2674 (O_2674,N_49648,N_49611);
or UO_2675 (O_2675,N_49641,N_49733);
xor UO_2676 (O_2676,N_49842,N_49539);
or UO_2677 (O_2677,N_49912,N_49879);
or UO_2678 (O_2678,N_49885,N_49523);
nor UO_2679 (O_2679,N_49775,N_49646);
nand UO_2680 (O_2680,N_49719,N_49826);
nand UO_2681 (O_2681,N_49835,N_49865);
xnor UO_2682 (O_2682,N_49820,N_49960);
and UO_2683 (O_2683,N_49571,N_49852);
xnor UO_2684 (O_2684,N_49979,N_49978);
and UO_2685 (O_2685,N_49726,N_49965);
nor UO_2686 (O_2686,N_49975,N_49664);
and UO_2687 (O_2687,N_49867,N_49733);
xor UO_2688 (O_2688,N_49879,N_49783);
or UO_2689 (O_2689,N_49742,N_49566);
nor UO_2690 (O_2690,N_49680,N_49768);
or UO_2691 (O_2691,N_49791,N_49733);
nor UO_2692 (O_2692,N_49591,N_49912);
or UO_2693 (O_2693,N_49580,N_49751);
or UO_2694 (O_2694,N_49735,N_49705);
xnor UO_2695 (O_2695,N_49704,N_49800);
nor UO_2696 (O_2696,N_49701,N_49600);
or UO_2697 (O_2697,N_49798,N_49779);
and UO_2698 (O_2698,N_49812,N_49711);
nand UO_2699 (O_2699,N_49868,N_49516);
nand UO_2700 (O_2700,N_49776,N_49805);
nand UO_2701 (O_2701,N_49754,N_49870);
nand UO_2702 (O_2702,N_49748,N_49930);
xnor UO_2703 (O_2703,N_49801,N_49867);
xnor UO_2704 (O_2704,N_49687,N_49759);
xnor UO_2705 (O_2705,N_49614,N_49988);
nand UO_2706 (O_2706,N_49522,N_49520);
and UO_2707 (O_2707,N_49745,N_49770);
and UO_2708 (O_2708,N_49967,N_49548);
nor UO_2709 (O_2709,N_49766,N_49720);
and UO_2710 (O_2710,N_49500,N_49850);
or UO_2711 (O_2711,N_49612,N_49636);
nand UO_2712 (O_2712,N_49513,N_49958);
xor UO_2713 (O_2713,N_49925,N_49544);
xnor UO_2714 (O_2714,N_49683,N_49893);
nor UO_2715 (O_2715,N_49709,N_49940);
or UO_2716 (O_2716,N_49687,N_49858);
nand UO_2717 (O_2717,N_49910,N_49667);
xor UO_2718 (O_2718,N_49719,N_49730);
or UO_2719 (O_2719,N_49637,N_49780);
or UO_2720 (O_2720,N_49560,N_49567);
nand UO_2721 (O_2721,N_49627,N_49556);
or UO_2722 (O_2722,N_49662,N_49889);
nor UO_2723 (O_2723,N_49689,N_49586);
or UO_2724 (O_2724,N_49713,N_49755);
or UO_2725 (O_2725,N_49592,N_49895);
xor UO_2726 (O_2726,N_49973,N_49634);
nor UO_2727 (O_2727,N_49792,N_49737);
nor UO_2728 (O_2728,N_49619,N_49996);
and UO_2729 (O_2729,N_49944,N_49530);
nor UO_2730 (O_2730,N_49602,N_49735);
nand UO_2731 (O_2731,N_49556,N_49964);
nor UO_2732 (O_2732,N_49509,N_49850);
nor UO_2733 (O_2733,N_49994,N_49588);
xor UO_2734 (O_2734,N_49541,N_49892);
or UO_2735 (O_2735,N_49759,N_49989);
or UO_2736 (O_2736,N_49958,N_49892);
and UO_2737 (O_2737,N_49911,N_49638);
nand UO_2738 (O_2738,N_49742,N_49512);
or UO_2739 (O_2739,N_49687,N_49723);
nor UO_2740 (O_2740,N_49782,N_49573);
nor UO_2741 (O_2741,N_49523,N_49586);
or UO_2742 (O_2742,N_49883,N_49526);
nor UO_2743 (O_2743,N_49655,N_49861);
xor UO_2744 (O_2744,N_49934,N_49773);
nand UO_2745 (O_2745,N_49683,N_49700);
and UO_2746 (O_2746,N_49928,N_49534);
nor UO_2747 (O_2747,N_49950,N_49972);
nor UO_2748 (O_2748,N_49581,N_49834);
xor UO_2749 (O_2749,N_49875,N_49903);
xor UO_2750 (O_2750,N_49541,N_49777);
xor UO_2751 (O_2751,N_49899,N_49504);
nor UO_2752 (O_2752,N_49734,N_49776);
nand UO_2753 (O_2753,N_49633,N_49873);
xor UO_2754 (O_2754,N_49740,N_49540);
nand UO_2755 (O_2755,N_49607,N_49705);
or UO_2756 (O_2756,N_49534,N_49913);
xor UO_2757 (O_2757,N_49857,N_49631);
xor UO_2758 (O_2758,N_49772,N_49749);
nor UO_2759 (O_2759,N_49520,N_49855);
nor UO_2760 (O_2760,N_49546,N_49973);
xnor UO_2761 (O_2761,N_49837,N_49582);
and UO_2762 (O_2762,N_49519,N_49822);
xnor UO_2763 (O_2763,N_49581,N_49545);
nor UO_2764 (O_2764,N_49572,N_49601);
nor UO_2765 (O_2765,N_49678,N_49590);
or UO_2766 (O_2766,N_49642,N_49824);
and UO_2767 (O_2767,N_49815,N_49584);
or UO_2768 (O_2768,N_49953,N_49995);
xnor UO_2769 (O_2769,N_49872,N_49775);
nor UO_2770 (O_2770,N_49926,N_49903);
nand UO_2771 (O_2771,N_49950,N_49557);
nand UO_2772 (O_2772,N_49777,N_49502);
nor UO_2773 (O_2773,N_49940,N_49605);
xor UO_2774 (O_2774,N_49531,N_49689);
xor UO_2775 (O_2775,N_49994,N_49521);
xnor UO_2776 (O_2776,N_49844,N_49690);
nand UO_2777 (O_2777,N_49690,N_49757);
nor UO_2778 (O_2778,N_49533,N_49861);
and UO_2779 (O_2779,N_49710,N_49748);
nor UO_2780 (O_2780,N_49858,N_49625);
nor UO_2781 (O_2781,N_49668,N_49853);
and UO_2782 (O_2782,N_49719,N_49863);
nand UO_2783 (O_2783,N_49676,N_49607);
nor UO_2784 (O_2784,N_49878,N_49924);
nand UO_2785 (O_2785,N_49749,N_49892);
nor UO_2786 (O_2786,N_49817,N_49944);
or UO_2787 (O_2787,N_49679,N_49656);
or UO_2788 (O_2788,N_49652,N_49971);
or UO_2789 (O_2789,N_49979,N_49985);
xor UO_2790 (O_2790,N_49675,N_49743);
and UO_2791 (O_2791,N_49896,N_49578);
and UO_2792 (O_2792,N_49759,N_49682);
or UO_2793 (O_2793,N_49810,N_49604);
nor UO_2794 (O_2794,N_49820,N_49590);
xnor UO_2795 (O_2795,N_49585,N_49828);
and UO_2796 (O_2796,N_49887,N_49774);
nor UO_2797 (O_2797,N_49886,N_49690);
nor UO_2798 (O_2798,N_49956,N_49688);
xor UO_2799 (O_2799,N_49864,N_49958);
and UO_2800 (O_2800,N_49771,N_49899);
or UO_2801 (O_2801,N_49620,N_49774);
nor UO_2802 (O_2802,N_49582,N_49629);
nand UO_2803 (O_2803,N_49636,N_49641);
and UO_2804 (O_2804,N_49529,N_49802);
or UO_2805 (O_2805,N_49610,N_49908);
nor UO_2806 (O_2806,N_49513,N_49761);
and UO_2807 (O_2807,N_49795,N_49751);
nand UO_2808 (O_2808,N_49775,N_49997);
nand UO_2809 (O_2809,N_49808,N_49712);
and UO_2810 (O_2810,N_49861,N_49503);
nand UO_2811 (O_2811,N_49791,N_49617);
xor UO_2812 (O_2812,N_49692,N_49791);
nor UO_2813 (O_2813,N_49681,N_49664);
nand UO_2814 (O_2814,N_49981,N_49881);
or UO_2815 (O_2815,N_49573,N_49847);
and UO_2816 (O_2816,N_49858,N_49983);
nor UO_2817 (O_2817,N_49533,N_49816);
nand UO_2818 (O_2818,N_49842,N_49543);
and UO_2819 (O_2819,N_49589,N_49528);
and UO_2820 (O_2820,N_49881,N_49976);
nor UO_2821 (O_2821,N_49521,N_49683);
or UO_2822 (O_2822,N_49780,N_49782);
and UO_2823 (O_2823,N_49608,N_49601);
or UO_2824 (O_2824,N_49587,N_49821);
nor UO_2825 (O_2825,N_49610,N_49655);
xnor UO_2826 (O_2826,N_49991,N_49931);
or UO_2827 (O_2827,N_49513,N_49927);
nor UO_2828 (O_2828,N_49621,N_49948);
nand UO_2829 (O_2829,N_49924,N_49670);
or UO_2830 (O_2830,N_49945,N_49886);
and UO_2831 (O_2831,N_49674,N_49574);
nand UO_2832 (O_2832,N_49552,N_49624);
nor UO_2833 (O_2833,N_49527,N_49737);
nor UO_2834 (O_2834,N_49540,N_49899);
or UO_2835 (O_2835,N_49643,N_49934);
nor UO_2836 (O_2836,N_49980,N_49802);
and UO_2837 (O_2837,N_49508,N_49612);
xnor UO_2838 (O_2838,N_49840,N_49502);
or UO_2839 (O_2839,N_49868,N_49629);
nand UO_2840 (O_2840,N_49684,N_49632);
or UO_2841 (O_2841,N_49765,N_49842);
xor UO_2842 (O_2842,N_49593,N_49834);
and UO_2843 (O_2843,N_49642,N_49706);
xnor UO_2844 (O_2844,N_49786,N_49955);
xor UO_2845 (O_2845,N_49571,N_49934);
nand UO_2846 (O_2846,N_49561,N_49828);
xor UO_2847 (O_2847,N_49767,N_49801);
or UO_2848 (O_2848,N_49959,N_49629);
nor UO_2849 (O_2849,N_49925,N_49710);
or UO_2850 (O_2850,N_49854,N_49978);
or UO_2851 (O_2851,N_49714,N_49780);
xor UO_2852 (O_2852,N_49734,N_49502);
and UO_2853 (O_2853,N_49810,N_49655);
nor UO_2854 (O_2854,N_49858,N_49869);
or UO_2855 (O_2855,N_49733,N_49824);
or UO_2856 (O_2856,N_49830,N_49979);
nor UO_2857 (O_2857,N_49766,N_49679);
nand UO_2858 (O_2858,N_49887,N_49638);
nand UO_2859 (O_2859,N_49543,N_49882);
xnor UO_2860 (O_2860,N_49695,N_49902);
xnor UO_2861 (O_2861,N_49642,N_49611);
and UO_2862 (O_2862,N_49935,N_49973);
nor UO_2863 (O_2863,N_49668,N_49970);
nor UO_2864 (O_2864,N_49869,N_49516);
or UO_2865 (O_2865,N_49517,N_49598);
xor UO_2866 (O_2866,N_49917,N_49580);
or UO_2867 (O_2867,N_49634,N_49693);
nor UO_2868 (O_2868,N_49579,N_49577);
or UO_2869 (O_2869,N_49907,N_49946);
nand UO_2870 (O_2870,N_49677,N_49693);
nand UO_2871 (O_2871,N_49979,N_49739);
or UO_2872 (O_2872,N_49531,N_49994);
and UO_2873 (O_2873,N_49900,N_49798);
xor UO_2874 (O_2874,N_49825,N_49543);
xnor UO_2875 (O_2875,N_49673,N_49605);
and UO_2876 (O_2876,N_49914,N_49964);
nand UO_2877 (O_2877,N_49816,N_49834);
nor UO_2878 (O_2878,N_49752,N_49796);
or UO_2879 (O_2879,N_49713,N_49525);
and UO_2880 (O_2880,N_49974,N_49756);
nor UO_2881 (O_2881,N_49513,N_49899);
xor UO_2882 (O_2882,N_49838,N_49884);
and UO_2883 (O_2883,N_49542,N_49819);
xor UO_2884 (O_2884,N_49706,N_49663);
nor UO_2885 (O_2885,N_49893,N_49641);
and UO_2886 (O_2886,N_49980,N_49819);
nand UO_2887 (O_2887,N_49780,N_49797);
xnor UO_2888 (O_2888,N_49509,N_49659);
nand UO_2889 (O_2889,N_49868,N_49953);
nor UO_2890 (O_2890,N_49528,N_49921);
xnor UO_2891 (O_2891,N_49888,N_49721);
nand UO_2892 (O_2892,N_49842,N_49987);
nor UO_2893 (O_2893,N_49512,N_49601);
or UO_2894 (O_2894,N_49711,N_49814);
nor UO_2895 (O_2895,N_49561,N_49625);
and UO_2896 (O_2896,N_49771,N_49525);
xnor UO_2897 (O_2897,N_49864,N_49565);
nand UO_2898 (O_2898,N_49521,N_49964);
xor UO_2899 (O_2899,N_49862,N_49791);
nand UO_2900 (O_2900,N_49980,N_49756);
and UO_2901 (O_2901,N_49617,N_49544);
nor UO_2902 (O_2902,N_49561,N_49843);
or UO_2903 (O_2903,N_49694,N_49805);
nor UO_2904 (O_2904,N_49538,N_49831);
nand UO_2905 (O_2905,N_49550,N_49547);
xor UO_2906 (O_2906,N_49909,N_49838);
and UO_2907 (O_2907,N_49806,N_49745);
nor UO_2908 (O_2908,N_49979,N_49828);
nand UO_2909 (O_2909,N_49939,N_49634);
and UO_2910 (O_2910,N_49970,N_49529);
or UO_2911 (O_2911,N_49846,N_49858);
and UO_2912 (O_2912,N_49848,N_49830);
nand UO_2913 (O_2913,N_49886,N_49740);
or UO_2914 (O_2914,N_49955,N_49880);
or UO_2915 (O_2915,N_49731,N_49630);
nor UO_2916 (O_2916,N_49604,N_49872);
nand UO_2917 (O_2917,N_49705,N_49764);
and UO_2918 (O_2918,N_49967,N_49673);
nand UO_2919 (O_2919,N_49646,N_49769);
or UO_2920 (O_2920,N_49884,N_49621);
xor UO_2921 (O_2921,N_49514,N_49880);
and UO_2922 (O_2922,N_49635,N_49759);
nand UO_2923 (O_2923,N_49613,N_49608);
xor UO_2924 (O_2924,N_49854,N_49916);
or UO_2925 (O_2925,N_49584,N_49593);
and UO_2926 (O_2926,N_49786,N_49543);
nor UO_2927 (O_2927,N_49870,N_49601);
xor UO_2928 (O_2928,N_49852,N_49765);
xor UO_2929 (O_2929,N_49634,N_49509);
or UO_2930 (O_2930,N_49926,N_49900);
xor UO_2931 (O_2931,N_49682,N_49639);
or UO_2932 (O_2932,N_49771,N_49863);
and UO_2933 (O_2933,N_49804,N_49810);
nand UO_2934 (O_2934,N_49512,N_49897);
nand UO_2935 (O_2935,N_49691,N_49552);
nand UO_2936 (O_2936,N_49892,N_49593);
nor UO_2937 (O_2937,N_49722,N_49892);
xnor UO_2938 (O_2938,N_49945,N_49559);
nand UO_2939 (O_2939,N_49913,N_49821);
nand UO_2940 (O_2940,N_49543,N_49640);
or UO_2941 (O_2941,N_49731,N_49760);
and UO_2942 (O_2942,N_49700,N_49858);
and UO_2943 (O_2943,N_49883,N_49968);
xnor UO_2944 (O_2944,N_49619,N_49970);
nand UO_2945 (O_2945,N_49535,N_49576);
and UO_2946 (O_2946,N_49694,N_49935);
or UO_2947 (O_2947,N_49767,N_49945);
nor UO_2948 (O_2948,N_49860,N_49867);
or UO_2949 (O_2949,N_49798,N_49786);
nand UO_2950 (O_2950,N_49508,N_49908);
and UO_2951 (O_2951,N_49905,N_49626);
nand UO_2952 (O_2952,N_49878,N_49725);
xnor UO_2953 (O_2953,N_49773,N_49836);
and UO_2954 (O_2954,N_49839,N_49759);
nor UO_2955 (O_2955,N_49915,N_49515);
nor UO_2956 (O_2956,N_49628,N_49581);
and UO_2957 (O_2957,N_49606,N_49884);
or UO_2958 (O_2958,N_49756,N_49833);
or UO_2959 (O_2959,N_49998,N_49966);
and UO_2960 (O_2960,N_49865,N_49779);
or UO_2961 (O_2961,N_49837,N_49913);
nand UO_2962 (O_2962,N_49782,N_49775);
and UO_2963 (O_2963,N_49689,N_49798);
and UO_2964 (O_2964,N_49655,N_49813);
or UO_2965 (O_2965,N_49508,N_49625);
nand UO_2966 (O_2966,N_49831,N_49847);
or UO_2967 (O_2967,N_49761,N_49865);
nand UO_2968 (O_2968,N_49715,N_49924);
xnor UO_2969 (O_2969,N_49642,N_49652);
nor UO_2970 (O_2970,N_49909,N_49835);
xnor UO_2971 (O_2971,N_49979,N_49932);
xnor UO_2972 (O_2972,N_49891,N_49799);
nand UO_2973 (O_2973,N_49992,N_49559);
or UO_2974 (O_2974,N_49746,N_49632);
xor UO_2975 (O_2975,N_49609,N_49633);
nand UO_2976 (O_2976,N_49583,N_49694);
or UO_2977 (O_2977,N_49631,N_49669);
xor UO_2978 (O_2978,N_49927,N_49996);
or UO_2979 (O_2979,N_49865,N_49622);
and UO_2980 (O_2980,N_49681,N_49896);
nor UO_2981 (O_2981,N_49638,N_49871);
and UO_2982 (O_2982,N_49771,N_49994);
xor UO_2983 (O_2983,N_49851,N_49753);
or UO_2984 (O_2984,N_49692,N_49650);
xnor UO_2985 (O_2985,N_49902,N_49647);
and UO_2986 (O_2986,N_49661,N_49708);
or UO_2987 (O_2987,N_49597,N_49931);
or UO_2988 (O_2988,N_49742,N_49923);
and UO_2989 (O_2989,N_49504,N_49855);
xor UO_2990 (O_2990,N_49951,N_49906);
nand UO_2991 (O_2991,N_49976,N_49882);
xor UO_2992 (O_2992,N_49683,N_49715);
nor UO_2993 (O_2993,N_49816,N_49846);
xnor UO_2994 (O_2994,N_49720,N_49735);
xor UO_2995 (O_2995,N_49908,N_49771);
nand UO_2996 (O_2996,N_49609,N_49908);
nor UO_2997 (O_2997,N_49731,N_49591);
nor UO_2998 (O_2998,N_49676,N_49616);
nor UO_2999 (O_2999,N_49533,N_49663);
nand UO_3000 (O_3000,N_49933,N_49951);
xnor UO_3001 (O_3001,N_49696,N_49897);
xor UO_3002 (O_3002,N_49530,N_49962);
and UO_3003 (O_3003,N_49603,N_49669);
xnor UO_3004 (O_3004,N_49804,N_49792);
nor UO_3005 (O_3005,N_49690,N_49979);
xor UO_3006 (O_3006,N_49627,N_49997);
or UO_3007 (O_3007,N_49568,N_49901);
or UO_3008 (O_3008,N_49661,N_49755);
xnor UO_3009 (O_3009,N_49717,N_49919);
and UO_3010 (O_3010,N_49790,N_49781);
xor UO_3011 (O_3011,N_49546,N_49578);
xnor UO_3012 (O_3012,N_49931,N_49801);
nand UO_3013 (O_3013,N_49555,N_49793);
or UO_3014 (O_3014,N_49929,N_49873);
or UO_3015 (O_3015,N_49939,N_49855);
nor UO_3016 (O_3016,N_49605,N_49891);
nor UO_3017 (O_3017,N_49523,N_49884);
nand UO_3018 (O_3018,N_49630,N_49615);
and UO_3019 (O_3019,N_49964,N_49884);
xnor UO_3020 (O_3020,N_49975,N_49937);
nand UO_3021 (O_3021,N_49756,N_49998);
or UO_3022 (O_3022,N_49920,N_49501);
nand UO_3023 (O_3023,N_49783,N_49792);
nand UO_3024 (O_3024,N_49775,N_49832);
and UO_3025 (O_3025,N_49728,N_49743);
or UO_3026 (O_3026,N_49631,N_49695);
or UO_3027 (O_3027,N_49754,N_49630);
nor UO_3028 (O_3028,N_49707,N_49973);
nor UO_3029 (O_3029,N_49967,N_49838);
nor UO_3030 (O_3030,N_49587,N_49572);
nand UO_3031 (O_3031,N_49653,N_49659);
nor UO_3032 (O_3032,N_49653,N_49985);
or UO_3033 (O_3033,N_49814,N_49617);
nor UO_3034 (O_3034,N_49894,N_49767);
and UO_3035 (O_3035,N_49636,N_49652);
nand UO_3036 (O_3036,N_49852,N_49728);
nor UO_3037 (O_3037,N_49803,N_49673);
xnor UO_3038 (O_3038,N_49945,N_49929);
xnor UO_3039 (O_3039,N_49929,N_49748);
and UO_3040 (O_3040,N_49787,N_49694);
nand UO_3041 (O_3041,N_49655,N_49586);
nand UO_3042 (O_3042,N_49987,N_49756);
xor UO_3043 (O_3043,N_49569,N_49936);
nor UO_3044 (O_3044,N_49624,N_49819);
and UO_3045 (O_3045,N_49830,N_49754);
and UO_3046 (O_3046,N_49843,N_49642);
nand UO_3047 (O_3047,N_49784,N_49720);
nand UO_3048 (O_3048,N_49907,N_49598);
or UO_3049 (O_3049,N_49506,N_49633);
or UO_3050 (O_3050,N_49601,N_49590);
and UO_3051 (O_3051,N_49510,N_49719);
nand UO_3052 (O_3052,N_49685,N_49652);
nor UO_3053 (O_3053,N_49540,N_49618);
xor UO_3054 (O_3054,N_49791,N_49951);
nand UO_3055 (O_3055,N_49718,N_49924);
xnor UO_3056 (O_3056,N_49766,N_49904);
or UO_3057 (O_3057,N_49618,N_49786);
nor UO_3058 (O_3058,N_49616,N_49537);
or UO_3059 (O_3059,N_49510,N_49877);
and UO_3060 (O_3060,N_49649,N_49952);
or UO_3061 (O_3061,N_49770,N_49845);
xor UO_3062 (O_3062,N_49767,N_49971);
and UO_3063 (O_3063,N_49766,N_49578);
xor UO_3064 (O_3064,N_49562,N_49907);
and UO_3065 (O_3065,N_49505,N_49648);
nor UO_3066 (O_3066,N_49962,N_49847);
nor UO_3067 (O_3067,N_49602,N_49622);
or UO_3068 (O_3068,N_49711,N_49963);
nor UO_3069 (O_3069,N_49822,N_49676);
nand UO_3070 (O_3070,N_49749,N_49889);
and UO_3071 (O_3071,N_49939,N_49955);
or UO_3072 (O_3072,N_49771,N_49524);
and UO_3073 (O_3073,N_49573,N_49828);
or UO_3074 (O_3074,N_49625,N_49611);
xor UO_3075 (O_3075,N_49692,N_49624);
or UO_3076 (O_3076,N_49915,N_49636);
xnor UO_3077 (O_3077,N_49998,N_49879);
or UO_3078 (O_3078,N_49674,N_49654);
nor UO_3079 (O_3079,N_49774,N_49727);
xor UO_3080 (O_3080,N_49668,N_49780);
nor UO_3081 (O_3081,N_49628,N_49923);
or UO_3082 (O_3082,N_49931,N_49872);
nand UO_3083 (O_3083,N_49523,N_49658);
nor UO_3084 (O_3084,N_49748,N_49669);
xnor UO_3085 (O_3085,N_49589,N_49837);
nand UO_3086 (O_3086,N_49603,N_49733);
nand UO_3087 (O_3087,N_49838,N_49885);
nor UO_3088 (O_3088,N_49629,N_49846);
xnor UO_3089 (O_3089,N_49906,N_49794);
xor UO_3090 (O_3090,N_49650,N_49761);
xor UO_3091 (O_3091,N_49799,N_49834);
xor UO_3092 (O_3092,N_49688,N_49930);
nor UO_3093 (O_3093,N_49999,N_49525);
or UO_3094 (O_3094,N_49973,N_49622);
or UO_3095 (O_3095,N_49666,N_49903);
or UO_3096 (O_3096,N_49652,N_49632);
nand UO_3097 (O_3097,N_49846,N_49690);
or UO_3098 (O_3098,N_49812,N_49652);
or UO_3099 (O_3099,N_49563,N_49516);
and UO_3100 (O_3100,N_49822,N_49575);
and UO_3101 (O_3101,N_49776,N_49608);
nor UO_3102 (O_3102,N_49637,N_49994);
and UO_3103 (O_3103,N_49939,N_49569);
and UO_3104 (O_3104,N_49708,N_49937);
nor UO_3105 (O_3105,N_49844,N_49887);
nor UO_3106 (O_3106,N_49942,N_49574);
nor UO_3107 (O_3107,N_49841,N_49764);
or UO_3108 (O_3108,N_49641,N_49650);
xor UO_3109 (O_3109,N_49730,N_49571);
or UO_3110 (O_3110,N_49715,N_49553);
nor UO_3111 (O_3111,N_49546,N_49772);
or UO_3112 (O_3112,N_49512,N_49815);
nor UO_3113 (O_3113,N_49886,N_49844);
xor UO_3114 (O_3114,N_49974,N_49792);
or UO_3115 (O_3115,N_49980,N_49605);
and UO_3116 (O_3116,N_49556,N_49612);
nor UO_3117 (O_3117,N_49966,N_49927);
xnor UO_3118 (O_3118,N_49932,N_49801);
nor UO_3119 (O_3119,N_49891,N_49606);
or UO_3120 (O_3120,N_49828,N_49693);
nand UO_3121 (O_3121,N_49895,N_49653);
nor UO_3122 (O_3122,N_49878,N_49653);
xnor UO_3123 (O_3123,N_49720,N_49814);
nor UO_3124 (O_3124,N_49502,N_49629);
xor UO_3125 (O_3125,N_49763,N_49877);
and UO_3126 (O_3126,N_49825,N_49777);
nor UO_3127 (O_3127,N_49540,N_49672);
or UO_3128 (O_3128,N_49947,N_49552);
nor UO_3129 (O_3129,N_49643,N_49964);
and UO_3130 (O_3130,N_49606,N_49994);
and UO_3131 (O_3131,N_49943,N_49801);
or UO_3132 (O_3132,N_49571,N_49516);
nand UO_3133 (O_3133,N_49610,N_49627);
or UO_3134 (O_3134,N_49613,N_49534);
or UO_3135 (O_3135,N_49787,N_49998);
or UO_3136 (O_3136,N_49556,N_49870);
or UO_3137 (O_3137,N_49699,N_49695);
nor UO_3138 (O_3138,N_49564,N_49742);
xnor UO_3139 (O_3139,N_49533,N_49949);
and UO_3140 (O_3140,N_49986,N_49520);
nand UO_3141 (O_3141,N_49527,N_49746);
nand UO_3142 (O_3142,N_49857,N_49640);
nor UO_3143 (O_3143,N_49897,N_49559);
nand UO_3144 (O_3144,N_49736,N_49833);
nand UO_3145 (O_3145,N_49549,N_49861);
or UO_3146 (O_3146,N_49744,N_49625);
nor UO_3147 (O_3147,N_49809,N_49740);
and UO_3148 (O_3148,N_49611,N_49527);
nand UO_3149 (O_3149,N_49818,N_49881);
nand UO_3150 (O_3150,N_49945,N_49977);
and UO_3151 (O_3151,N_49890,N_49989);
nand UO_3152 (O_3152,N_49654,N_49669);
and UO_3153 (O_3153,N_49658,N_49589);
nor UO_3154 (O_3154,N_49834,N_49831);
and UO_3155 (O_3155,N_49674,N_49979);
xor UO_3156 (O_3156,N_49544,N_49570);
or UO_3157 (O_3157,N_49886,N_49558);
nand UO_3158 (O_3158,N_49563,N_49666);
nand UO_3159 (O_3159,N_49594,N_49509);
nand UO_3160 (O_3160,N_49890,N_49834);
or UO_3161 (O_3161,N_49682,N_49725);
nand UO_3162 (O_3162,N_49912,N_49959);
and UO_3163 (O_3163,N_49968,N_49536);
or UO_3164 (O_3164,N_49951,N_49680);
xnor UO_3165 (O_3165,N_49712,N_49985);
and UO_3166 (O_3166,N_49901,N_49809);
or UO_3167 (O_3167,N_49679,N_49690);
and UO_3168 (O_3168,N_49726,N_49674);
xnor UO_3169 (O_3169,N_49699,N_49805);
and UO_3170 (O_3170,N_49702,N_49915);
xor UO_3171 (O_3171,N_49538,N_49596);
nand UO_3172 (O_3172,N_49665,N_49526);
xor UO_3173 (O_3173,N_49788,N_49514);
or UO_3174 (O_3174,N_49751,N_49683);
xor UO_3175 (O_3175,N_49897,N_49741);
xor UO_3176 (O_3176,N_49775,N_49531);
nand UO_3177 (O_3177,N_49662,N_49589);
xor UO_3178 (O_3178,N_49844,N_49594);
and UO_3179 (O_3179,N_49888,N_49939);
xor UO_3180 (O_3180,N_49668,N_49816);
xnor UO_3181 (O_3181,N_49780,N_49921);
or UO_3182 (O_3182,N_49785,N_49527);
nand UO_3183 (O_3183,N_49555,N_49580);
nor UO_3184 (O_3184,N_49737,N_49858);
nand UO_3185 (O_3185,N_49888,N_49649);
nand UO_3186 (O_3186,N_49851,N_49525);
and UO_3187 (O_3187,N_49865,N_49943);
nand UO_3188 (O_3188,N_49997,N_49722);
and UO_3189 (O_3189,N_49789,N_49780);
nand UO_3190 (O_3190,N_49920,N_49626);
nand UO_3191 (O_3191,N_49812,N_49662);
nor UO_3192 (O_3192,N_49698,N_49655);
nand UO_3193 (O_3193,N_49849,N_49631);
nand UO_3194 (O_3194,N_49618,N_49957);
or UO_3195 (O_3195,N_49890,N_49759);
nor UO_3196 (O_3196,N_49602,N_49638);
nor UO_3197 (O_3197,N_49633,N_49577);
nand UO_3198 (O_3198,N_49843,N_49790);
or UO_3199 (O_3199,N_49653,N_49729);
or UO_3200 (O_3200,N_49815,N_49967);
nand UO_3201 (O_3201,N_49822,N_49931);
or UO_3202 (O_3202,N_49999,N_49559);
nand UO_3203 (O_3203,N_49503,N_49966);
xor UO_3204 (O_3204,N_49635,N_49949);
nand UO_3205 (O_3205,N_49949,N_49513);
xor UO_3206 (O_3206,N_49653,N_49630);
nor UO_3207 (O_3207,N_49904,N_49975);
xnor UO_3208 (O_3208,N_49599,N_49705);
and UO_3209 (O_3209,N_49709,N_49809);
or UO_3210 (O_3210,N_49887,N_49697);
nor UO_3211 (O_3211,N_49957,N_49605);
nor UO_3212 (O_3212,N_49560,N_49682);
and UO_3213 (O_3213,N_49546,N_49719);
nor UO_3214 (O_3214,N_49593,N_49763);
xor UO_3215 (O_3215,N_49587,N_49870);
xor UO_3216 (O_3216,N_49765,N_49962);
nor UO_3217 (O_3217,N_49627,N_49816);
and UO_3218 (O_3218,N_49867,N_49571);
xnor UO_3219 (O_3219,N_49531,N_49617);
or UO_3220 (O_3220,N_49952,N_49766);
nor UO_3221 (O_3221,N_49783,N_49997);
and UO_3222 (O_3222,N_49928,N_49567);
nand UO_3223 (O_3223,N_49548,N_49980);
xnor UO_3224 (O_3224,N_49827,N_49674);
and UO_3225 (O_3225,N_49943,N_49503);
and UO_3226 (O_3226,N_49620,N_49962);
and UO_3227 (O_3227,N_49515,N_49569);
xnor UO_3228 (O_3228,N_49749,N_49930);
or UO_3229 (O_3229,N_49993,N_49925);
and UO_3230 (O_3230,N_49824,N_49606);
nand UO_3231 (O_3231,N_49500,N_49908);
nor UO_3232 (O_3232,N_49653,N_49821);
xnor UO_3233 (O_3233,N_49965,N_49681);
nand UO_3234 (O_3234,N_49792,N_49705);
nor UO_3235 (O_3235,N_49548,N_49756);
or UO_3236 (O_3236,N_49565,N_49676);
nand UO_3237 (O_3237,N_49812,N_49572);
nor UO_3238 (O_3238,N_49921,N_49539);
nand UO_3239 (O_3239,N_49504,N_49751);
xnor UO_3240 (O_3240,N_49530,N_49683);
nand UO_3241 (O_3241,N_49763,N_49876);
or UO_3242 (O_3242,N_49829,N_49852);
xor UO_3243 (O_3243,N_49875,N_49550);
and UO_3244 (O_3244,N_49585,N_49924);
and UO_3245 (O_3245,N_49716,N_49795);
nor UO_3246 (O_3246,N_49719,N_49980);
or UO_3247 (O_3247,N_49821,N_49926);
xor UO_3248 (O_3248,N_49933,N_49856);
and UO_3249 (O_3249,N_49598,N_49512);
or UO_3250 (O_3250,N_49992,N_49921);
or UO_3251 (O_3251,N_49707,N_49561);
and UO_3252 (O_3252,N_49895,N_49533);
nand UO_3253 (O_3253,N_49724,N_49955);
and UO_3254 (O_3254,N_49815,N_49556);
and UO_3255 (O_3255,N_49964,N_49814);
nand UO_3256 (O_3256,N_49564,N_49917);
and UO_3257 (O_3257,N_49661,N_49784);
nor UO_3258 (O_3258,N_49848,N_49932);
nand UO_3259 (O_3259,N_49527,N_49812);
or UO_3260 (O_3260,N_49744,N_49624);
nand UO_3261 (O_3261,N_49744,N_49850);
xnor UO_3262 (O_3262,N_49843,N_49534);
nor UO_3263 (O_3263,N_49971,N_49908);
or UO_3264 (O_3264,N_49699,N_49939);
nor UO_3265 (O_3265,N_49992,N_49549);
and UO_3266 (O_3266,N_49652,N_49798);
nand UO_3267 (O_3267,N_49898,N_49961);
and UO_3268 (O_3268,N_49626,N_49785);
nand UO_3269 (O_3269,N_49679,N_49577);
xnor UO_3270 (O_3270,N_49916,N_49717);
and UO_3271 (O_3271,N_49715,N_49979);
nor UO_3272 (O_3272,N_49869,N_49917);
or UO_3273 (O_3273,N_49543,N_49639);
nand UO_3274 (O_3274,N_49516,N_49716);
nand UO_3275 (O_3275,N_49672,N_49588);
and UO_3276 (O_3276,N_49971,N_49997);
nand UO_3277 (O_3277,N_49649,N_49739);
and UO_3278 (O_3278,N_49907,N_49625);
or UO_3279 (O_3279,N_49877,N_49702);
nor UO_3280 (O_3280,N_49998,N_49609);
and UO_3281 (O_3281,N_49763,N_49989);
or UO_3282 (O_3282,N_49534,N_49596);
or UO_3283 (O_3283,N_49850,N_49501);
xnor UO_3284 (O_3284,N_49937,N_49965);
nand UO_3285 (O_3285,N_49705,N_49903);
nand UO_3286 (O_3286,N_49628,N_49559);
nor UO_3287 (O_3287,N_49743,N_49941);
and UO_3288 (O_3288,N_49547,N_49960);
and UO_3289 (O_3289,N_49614,N_49714);
or UO_3290 (O_3290,N_49648,N_49723);
xnor UO_3291 (O_3291,N_49526,N_49512);
nor UO_3292 (O_3292,N_49673,N_49892);
xnor UO_3293 (O_3293,N_49894,N_49846);
nand UO_3294 (O_3294,N_49885,N_49946);
nand UO_3295 (O_3295,N_49604,N_49520);
or UO_3296 (O_3296,N_49865,N_49627);
or UO_3297 (O_3297,N_49863,N_49563);
nand UO_3298 (O_3298,N_49878,N_49994);
nor UO_3299 (O_3299,N_49758,N_49877);
xnor UO_3300 (O_3300,N_49891,N_49969);
xor UO_3301 (O_3301,N_49927,N_49968);
and UO_3302 (O_3302,N_49775,N_49974);
and UO_3303 (O_3303,N_49655,N_49700);
and UO_3304 (O_3304,N_49954,N_49905);
xnor UO_3305 (O_3305,N_49734,N_49695);
xnor UO_3306 (O_3306,N_49685,N_49509);
and UO_3307 (O_3307,N_49516,N_49778);
nor UO_3308 (O_3308,N_49513,N_49734);
nand UO_3309 (O_3309,N_49637,N_49800);
or UO_3310 (O_3310,N_49656,N_49945);
nor UO_3311 (O_3311,N_49542,N_49893);
nor UO_3312 (O_3312,N_49689,N_49746);
and UO_3313 (O_3313,N_49967,N_49598);
xor UO_3314 (O_3314,N_49892,N_49957);
or UO_3315 (O_3315,N_49721,N_49986);
or UO_3316 (O_3316,N_49610,N_49654);
nor UO_3317 (O_3317,N_49820,N_49961);
or UO_3318 (O_3318,N_49655,N_49527);
and UO_3319 (O_3319,N_49905,N_49853);
and UO_3320 (O_3320,N_49783,N_49504);
nor UO_3321 (O_3321,N_49806,N_49580);
and UO_3322 (O_3322,N_49650,N_49800);
and UO_3323 (O_3323,N_49913,N_49978);
nor UO_3324 (O_3324,N_49531,N_49770);
xnor UO_3325 (O_3325,N_49590,N_49727);
xnor UO_3326 (O_3326,N_49558,N_49798);
nand UO_3327 (O_3327,N_49745,N_49728);
or UO_3328 (O_3328,N_49623,N_49884);
nand UO_3329 (O_3329,N_49704,N_49591);
nor UO_3330 (O_3330,N_49805,N_49645);
and UO_3331 (O_3331,N_49584,N_49646);
nand UO_3332 (O_3332,N_49553,N_49870);
xnor UO_3333 (O_3333,N_49649,N_49962);
xor UO_3334 (O_3334,N_49841,N_49525);
nor UO_3335 (O_3335,N_49596,N_49803);
xnor UO_3336 (O_3336,N_49643,N_49819);
xnor UO_3337 (O_3337,N_49502,N_49710);
nand UO_3338 (O_3338,N_49552,N_49968);
nor UO_3339 (O_3339,N_49909,N_49649);
nand UO_3340 (O_3340,N_49666,N_49762);
and UO_3341 (O_3341,N_49699,N_49860);
nand UO_3342 (O_3342,N_49740,N_49673);
nand UO_3343 (O_3343,N_49503,N_49557);
nand UO_3344 (O_3344,N_49950,N_49781);
nor UO_3345 (O_3345,N_49653,N_49575);
and UO_3346 (O_3346,N_49963,N_49949);
nor UO_3347 (O_3347,N_49990,N_49926);
nand UO_3348 (O_3348,N_49734,N_49896);
and UO_3349 (O_3349,N_49992,N_49669);
xor UO_3350 (O_3350,N_49604,N_49950);
or UO_3351 (O_3351,N_49880,N_49983);
nor UO_3352 (O_3352,N_49548,N_49696);
xor UO_3353 (O_3353,N_49633,N_49761);
or UO_3354 (O_3354,N_49531,N_49637);
nor UO_3355 (O_3355,N_49653,N_49652);
nor UO_3356 (O_3356,N_49902,N_49559);
xnor UO_3357 (O_3357,N_49696,N_49846);
and UO_3358 (O_3358,N_49618,N_49987);
nand UO_3359 (O_3359,N_49759,N_49742);
xor UO_3360 (O_3360,N_49826,N_49710);
nor UO_3361 (O_3361,N_49961,N_49766);
nor UO_3362 (O_3362,N_49824,N_49928);
xnor UO_3363 (O_3363,N_49544,N_49784);
or UO_3364 (O_3364,N_49677,N_49819);
nand UO_3365 (O_3365,N_49723,N_49622);
nor UO_3366 (O_3366,N_49555,N_49952);
nor UO_3367 (O_3367,N_49878,N_49747);
nand UO_3368 (O_3368,N_49958,N_49685);
nor UO_3369 (O_3369,N_49781,N_49867);
or UO_3370 (O_3370,N_49919,N_49507);
or UO_3371 (O_3371,N_49505,N_49838);
and UO_3372 (O_3372,N_49581,N_49502);
xnor UO_3373 (O_3373,N_49568,N_49820);
or UO_3374 (O_3374,N_49720,N_49760);
nand UO_3375 (O_3375,N_49700,N_49725);
nand UO_3376 (O_3376,N_49932,N_49943);
nand UO_3377 (O_3377,N_49723,N_49986);
nand UO_3378 (O_3378,N_49575,N_49850);
or UO_3379 (O_3379,N_49645,N_49500);
nand UO_3380 (O_3380,N_49533,N_49746);
and UO_3381 (O_3381,N_49905,N_49859);
nand UO_3382 (O_3382,N_49561,N_49544);
and UO_3383 (O_3383,N_49955,N_49645);
xor UO_3384 (O_3384,N_49626,N_49688);
and UO_3385 (O_3385,N_49502,N_49600);
nor UO_3386 (O_3386,N_49799,N_49875);
and UO_3387 (O_3387,N_49827,N_49723);
nor UO_3388 (O_3388,N_49532,N_49690);
nor UO_3389 (O_3389,N_49845,N_49696);
nor UO_3390 (O_3390,N_49578,N_49794);
or UO_3391 (O_3391,N_49828,N_49594);
xnor UO_3392 (O_3392,N_49689,N_49645);
and UO_3393 (O_3393,N_49540,N_49526);
and UO_3394 (O_3394,N_49658,N_49921);
nor UO_3395 (O_3395,N_49816,N_49681);
or UO_3396 (O_3396,N_49852,N_49995);
or UO_3397 (O_3397,N_49815,N_49973);
or UO_3398 (O_3398,N_49769,N_49847);
and UO_3399 (O_3399,N_49631,N_49622);
or UO_3400 (O_3400,N_49854,N_49963);
nor UO_3401 (O_3401,N_49984,N_49888);
and UO_3402 (O_3402,N_49787,N_49917);
xnor UO_3403 (O_3403,N_49576,N_49552);
nor UO_3404 (O_3404,N_49819,N_49903);
nor UO_3405 (O_3405,N_49946,N_49879);
and UO_3406 (O_3406,N_49571,N_49617);
xnor UO_3407 (O_3407,N_49708,N_49860);
and UO_3408 (O_3408,N_49589,N_49933);
or UO_3409 (O_3409,N_49585,N_49612);
nand UO_3410 (O_3410,N_49929,N_49980);
nand UO_3411 (O_3411,N_49674,N_49843);
nand UO_3412 (O_3412,N_49506,N_49530);
nand UO_3413 (O_3413,N_49851,N_49903);
or UO_3414 (O_3414,N_49800,N_49533);
xor UO_3415 (O_3415,N_49970,N_49535);
nor UO_3416 (O_3416,N_49768,N_49972);
and UO_3417 (O_3417,N_49626,N_49587);
nor UO_3418 (O_3418,N_49870,N_49932);
and UO_3419 (O_3419,N_49880,N_49669);
nor UO_3420 (O_3420,N_49551,N_49560);
nor UO_3421 (O_3421,N_49649,N_49829);
nand UO_3422 (O_3422,N_49640,N_49560);
and UO_3423 (O_3423,N_49913,N_49979);
nor UO_3424 (O_3424,N_49878,N_49511);
and UO_3425 (O_3425,N_49903,N_49845);
or UO_3426 (O_3426,N_49976,N_49802);
and UO_3427 (O_3427,N_49745,N_49751);
nand UO_3428 (O_3428,N_49850,N_49624);
or UO_3429 (O_3429,N_49927,N_49690);
and UO_3430 (O_3430,N_49860,N_49920);
xnor UO_3431 (O_3431,N_49847,N_49805);
and UO_3432 (O_3432,N_49603,N_49705);
xor UO_3433 (O_3433,N_49657,N_49681);
nor UO_3434 (O_3434,N_49889,N_49875);
xnor UO_3435 (O_3435,N_49563,N_49828);
xnor UO_3436 (O_3436,N_49916,N_49515);
xor UO_3437 (O_3437,N_49644,N_49870);
nand UO_3438 (O_3438,N_49671,N_49942);
or UO_3439 (O_3439,N_49738,N_49510);
and UO_3440 (O_3440,N_49925,N_49650);
xnor UO_3441 (O_3441,N_49513,N_49780);
nand UO_3442 (O_3442,N_49937,N_49567);
xnor UO_3443 (O_3443,N_49853,N_49630);
and UO_3444 (O_3444,N_49565,N_49758);
and UO_3445 (O_3445,N_49997,N_49882);
nor UO_3446 (O_3446,N_49746,N_49588);
nand UO_3447 (O_3447,N_49914,N_49569);
nand UO_3448 (O_3448,N_49955,N_49663);
nor UO_3449 (O_3449,N_49862,N_49977);
xnor UO_3450 (O_3450,N_49632,N_49660);
nand UO_3451 (O_3451,N_49540,N_49626);
xor UO_3452 (O_3452,N_49556,N_49618);
nand UO_3453 (O_3453,N_49511,N_49806);
nor UO_3454 (O_3454,N_49971,N_49837);
nand UO_3455 (O_3455,N_49632,N_49519);
and UO_3456 (O_3456,N_49547,N_49588);
nor UO_3457 (O_3457,N_49602,N_49504);
and UO_3458 (O_3458,N_49882,N_49793);
or UO_3459 (O_3459,N_49657,N_49841);
nor UO_3460 (O_3460,N_49557,N_49523);
or UO_3461 (O_3461,N_49565,N_49505);
xnor UO_3462 (O_3462,N_49676,N_49726);
nand UO_3463 (O_3463,N_49985,N_49548);
xor UO_3464 (O_3464,N_49947,N_49996);
or UO_3465 (O_3465,N_49842,N_49738);
nor UO_3466 (O_3466,N_49995,N_49827);
xnor UO_3467 (O_3467,N_49683,N_49661);
xnor UO_3468 (O_3468,N_49623,N_49870);
xor UO_3469 (O_3469,N_49530,N_49508);
xor UO_3470 (O_3470,N_49670,N_49964);
nor UO_3471 (O_3471,N_49843,N_49667);
nor UO_3472 (O_3472,N_49875,N_49679);
nor UO_3473 (O_3473,N_49696,N_49744);
or UO_3474 (O_3474,N_49938,N_49532);
nand UO_3475 (O_3475,N_49943,N_49531);
nor UO_3476 (O_3476,N_49827,N_49812);
xnor UO_3477 (O_3477,N_49547,N_49564);
nand UO_3478 (O_3478,N_49783,N_49663);
nand UO_3479 (O_3479,N_49835,N_49575);
nand UO_3480 (O_3480,N_49671,N_49819);
and UO_3481 (O_3481,N_49672,N_49947);
nor UO_3482 (O_3482,N_49526,N_49829);
and UO_3483 (O_3483,N_49632,N_49797);
xnor UO_3484 (O_3484,N_49863,N_49899);
or UO_3485 (O_3485,N_49563,N_49743);
nor UO_3486 (O_3486,N_49946,N_49880);
xor UO_3487 (O_3487,N_49914,N_49886);
and UO_3488 (O_3488,N_49700,N_49551);
nor UO_3489 (O_3489,N_49986,N_49902);
xnor UO_3490 (O_3490,N_49701,N_49618);
or UO_3491 (O_3491,N_49561,N_49928);
and UO_3492 (O_3492,N_49966,N_49800);
nor UO_3493 (O_3493,N_49757,N_49824);
nor UO_3494 (O_3494,N_49531,N_49876);
xor UO_3495 (O_3495,N_49675,N_49635);
nor UO_3496 (O_3496,N_49686,N_49908);
or UO_3497 (O_3497,N_49569,N_49831);
or UO_3498 (O_3498,N_49633,N_49859);
and UO_3499 (O_3499,N_49562,N_49953);
nor UO_3500 (O_3500,N_49876,N_49770);
nand UO_3501 (O_3501,N_49662,N_49545);
nand UO_3502 (O_3502,N_49658,N_49666);
nand UO_3503 (O_3503,N_49791,N_49804);
xnor UO_3504 (O_3504,N_49971,N_49646);
nand UO_3505 (O_3505,N_49764,N_49569);
and UO_3506 (O_3506,N_49909,N_49968);
xnor UO_3507 (O_3507,N_49660,N_49672);
or UO_3508 (O_3508,N_49630,N_49925);
nand UO_3509 (O_3509,N_49975,N_49997);
nor UO_3510 (O_3510,N_49934,N_49778);
xor UO_3511 (O_3511,N_49568,N_49536);
and UO_3512 (O_3512,N_49557,N_49944);
and UO_3513 (O_3513,N_49708,N_49999);
or UO_3514 (O_3514,N_49858,N_49632);
nand UO_3515 (O_3515,N_49614,N_49613);
xor UO_3516 (O_3516,N_49631,N_49608);
xor UO_3517 (O_3517,N_49836,N_49580);
or UO_3518 (O_3518,N_49712,N_49780);
nor UO_3519 (O_3519,N_49863,N_49544);
xor UO_3520 (O_3520,N_49987,N_49638);
or UO_3521 (O_3521,N_49512,N_49948);
or UO_3522 (O_3522,N_49696,N_49720);
or UO_3523 (O_3523,N_49665,N_49613);
nor UO_3524 (O_3524,N_49615,N_49927);
xnor UO_3525 (O_3525,N_49626,N_49516);
nor UO_3526 (O_3526,N_49961,N_49755);
or UO_3527 (O_3527,N_49588,N_49622);
and UO_3528 (O_3528,N_49532,N_49508);
nor UO_3529 (O_3529,N_49843,N_49603);
and UO_3530 (O_3530,N_49597,N_49988);
or UO_3531 (O_3531,N_49571,N_49596);
and UO_3532 (O_3532,N_49718,N_49524);
nand UO_3533 (O_3533,N_49582,N_49825);
nor UO_3534 (O_3534,N_49737,N_49868);
or UO_3535 (O_3535,N_49626,N_49993);
and UO_3536 (O_3536,N_49506,N_49778);
xor UO_3537 (O_3537,N_49736,N_49603);
nor UO_3538 (O_3538,N_49968,N_49701);
and UO_3539 (O_3539,N_49715,N_49642);
nand UO_3540 (O_3540,N_49557,N_49882);
nand UO_3541 (O_3541,N_49691,N_49536);
nor UO_3542 (O_3542,N_49676,N_49844);
or UO_3543 (O_3543,N_49773,N_49753);
nand UO_3544 (O_3544,N_49953,N_49612);
and UO_3545 (O_3545,N_49821,N_49837);
and UO_3546 (O_3546,N_49974,N_49868);
xnor UO_3547 (O_3547,N_49581,N_49583);
nor UO_3548 (O_3548,N_49822,N_49763);
xnor UO_3549 (O_3549,N_49831,N_49601);
and UO_3550 (O_3550,N_49844,N_49879);
nand UO_3551 (O_3551,N_49885,N_49525);
nor UO_3552 (O_3552,N_49505,N_49850);
nand UO_3553 (O_3553,N_49832,N_49728);
xor UO_3554 (O_3554,N_49645,N_49610);
nor UO_3555 (O_3555,N_49928,N_49582);
nand UO_3556 (O_3556,N_49844,N_49815);
nor UO_3557 (O_3557,N_49662,N_49979);
or UO_3558 (O_3558,N_49663,N_49785);
and UO_3559 (O_3559,N_49688,N_49960);
and UO_3560 (O_3560,N_49942,N_49895);
or UO_3561 (O_3561,N_49737,N_49825);
and UO_3562 (O_3562,N_49521,N_49809);
or UO_3563 (O_3563,N_49762,N_49724);
or UO_3564 (O_3564,N_49813,N_49542);
nor UO_3565 (O_3565,N_49671,N_49585);
xor UO_3566 (O_3566,N_49996,N_49664);
xor UO_3567 (O_3567,N_49899,N_49682);
xnor UO_3568 (O_3568,N_49936,N_49835);
nand UO_3569 (O_3569,N_49996,N_49709);
and UO_3570 (O_3570,N_49839,N_49690);
and UO_3571 (O_3571,N_49848,N_49593);
and UO_3572 (O_3572,N_49666,N_49671);
nand UO_3573 (O_3573,N_49693,N_49741);
xor UO_3574 (O_3574,N_49506,N_49763);
nor UO_3575 (O_3575,N_49769,N_49772);
nor UO_3576 (O_3576,N_49792,N_49921);
or UO_3577 (O_3577,N_49708,N_49672);
or UO_3578 (O_3578,N_49866,N_49933);
nand UO_3579 (O_3579,N_49624,N_49547);
or UO_3580 (O_3580,N_49727,N_49693);
xor UO_3581 (O_3581,N_49735,N_49604);
and UO_3582 (O_3582,N_49740,N_49730);
xnor UO_3583 (O_3583,N_49847,N_49621);
or UO_3584 (O_3584,N_49680,N_49847);
nand UO_3585 (O_3585,N_49674,N_49781);
xnor UO_3586 (O_3586,N_49599,N_49733);
nand UO_3587 (O_3587,N_49638,N_49957);
xor UO_3588 (O_3588,N_49788,N_49723);
nand UO_3589 (O_3589,N_49576,N_49962);
or UO_3590 (O_3590,N_49802,N_49619);
and UO_3591 (O_3591,N_49710,N_49949);
and UO_3592 (O_3592,N_49654,N_49970);
nor UO_3593 (O_3593,N_49939,N_49835);
nand UO_3594 (O_3594,N_49808,N_49571);
xnor UO_3595 (O_3595,N_49624,N_49713);
nor UO_3596 (O_3596,N_49954,N_49940);
nand UO_3597 (O_3597,N_49502,N_49750);
and UO_3598 (O_3598,N_49725,N_49505);
xnor UO_3599 (O_3599,N_49830,N_49927);
and UO_3600 (O_3600,N_49916,N_49671);
and UO_3601 (O_3601,N_49940,N_49675);
and UO_3602 (O_3602,N_49702,N_49741);
nor UO_3603 (O_3603,N_49825,N_49915);
or UO_3604 (O_3604,N_49975,N_49879);
xnor UO_3605 (O_3605,N_49785,N_49776);
nand UO_3606 (O_3606,N_49610,N_49930);
nor UO_3607 (O_3607,N_49958,N_49976);
and UO_3608 (O_3608,N_49792,N_49828);
nor UO_3609 (O_3609,N_49677,N_49673);
nand UO_3610 (O_3610,N_49652,N_49524);
xor UO_3611 (O_3611,N_49694,N_49524);
or UO_3612 (O_3612,N_49813,N_49590);
or UO_3613 (O_3613,N_49993,N_49708);
and UO_3614 (O_3614,N_49976,N_49514);
and UO_3615 (O_3615,N_49553,N_49867);
xor UO_3616 (O_3616,N_49634,N_49888);
nor UO_3617 (O_3617,N_49610,N_49911);
and UO_3618 (O_3618,N_49888,N_49812);
nand UO_3619 (O_3619,N_49803,N_49571);
nor UO_3620 (O_3620,N_49588,N_49769);
nand UO_3621 (O_3621,N_49559,N_49662);
nor UO_3622 (O_3622,N_49691,N_49571);
xor UO_3623 (O_3623,N_49713,N_49960);
nand UO_3624 (O_3624,N_49983,N_49777);
nand UO_3625 (O_3625,N_49546,N_49824);
nor UO_3626 (O_3626,N_49713,N_49532);
nor UO_3627 (O_3627,N_49540,N_49691);
nand UO_3628 (O_3628,N_49569,N_49871);
nor UO_3629 (O_3629,N_49912,N_49875);
nand UO_3630 (O_3630,N_49582,N_49528);
and UO_3631 (O_3631,N_49862,N_49770);
nand UO_3632 (O_3632,N_49619,N_49670);
and UO_3633 (O_3633,N_49505,N_49903);
xor UO_3634 (O_3634,N_49828,N_49767);
nor UO_3635 (O_3635,N_49656,N_49781);
xor UO_3636 (O_3636,N_49692,N_49819);
nor UO_3637 (O_3637,N_49645,N_49726);
nand UO_3638 (O_3638,N_49795,N_49593);
xnor UO_3639 (O_3639,N_49834,N_49610);
nand UO_3640 (O_3640,N_49657,N_49760);
nor UO_3641 (O_3641,N_49763,N_49607);
nor UO_3642 (O_3642,N_49922,N_49797);
xnor UO_3643 (O_3643,N_49589,N_49691);
nor UO_3644 (O_3644,N_49646,N_49955);
xor UO_3645 (O_3645,N_49735,N_49700);
xnor UO_3646 (O_3646,N_49676,N_49819);
nand UO_3647 (O_3647,N_49590,N_49941);
nor UO_3648 (O_3648,N_49709,N_49607);
and UO_3649 (O_3649,N_49957,N_49946);
or UO_3650 (O_3650,N_49546,N_49845);
and UO_3651 (O_3651,N_49653,N_49587);
xor UO_3652 (O_3652,N_49531,N_49750);
xnor UO_3653 (O_3653,N_49867,N_49663);
nor UO_3654 (O_3654,N_49852,N_49508);
or UO_3655 (O_3655,N_49552,N_49627);
xnor UO_3656 (O_3656,N_49605,N_49617);
or UO_3657 (O_3657,N_49818,N_49974);
xnor UO_3658 (O_3658,N_49531,N_49925);
xor UO_3659 (O_3659,N_49775,N_49691);
and UO_3660 (O_3660,N_49628,N_49870);
nand UO_3661 (O_3661,N_49567,N_49865);
xnor UO_3662 (O_3662,N_49954,N_49845);
nand UO_3663 (O_3663,N_49533,N_49923);
and UO_3664 (O_3664,N_49525,N_49904);
and UO_3665 (O_3665,N_49706,N_49789);
and UO_3666 (O_3666,N_49675,N_49977);
xor UO_3667 (O_3667,N_49658,N_49923);
nand UO_3668 (O_3668,N_49533,N_49948);
xor UO_3669 (O_3669,N_49915,N_49946);
or UO_3670 (O_3670,N_49600,N_49915);
nand UO_3671 (O_3671,N_49893,N_49989);
nor UO_3672 (O_3672,N_49542,N_49938);
xor UO_3673 (O_3673,N_49710,N_49834);
or UO_3674 (O_3674,N_49766,N_49542);
nor UO_3675 (O_3675,N_49904,N_49980);
nand UO_3676 (O_3676,N_49695,N_49822);
xor UO_3677 (O_3677,N_49716,N_49990);
nand UO_3678 (O_3678,N_49693,N_49712);
xor UO_3679 (O_3679,N_49834,N_49812);
and UO_3680 (O_3680,N_49905,N_49869);
and UO_3681 (O_3681,N_49668,N_49509);
nand UO_3682 (O_3682,N_49672,N_49809);
nand UO_3683 (O_3683,N_49770,N_49606);
or UO_3684 (O_3684,N_49987,N_49568);
or UO_3685 (O_3685,N_49979,N_49580);
and UO_3686 (O_3686,N_49516,N_49635);
or UO_3687 (O_3687,N_49644,N_49996);
xor UO_3688 (O_3688,N_49563,N_49554);
nor UO_3689 (O_3689,N_49977,N_49701);
and UO_3690 (O_3690,N_49705,N_49790);
and UO_3691 (O_3691,N_49774,N_49775);
xor UO_3692 (O_3692,N_49511,N_49804);
xnor UO_3693 (O_3693,N_49502,N_49762);
or UO_3694 (O_3694,N_49792,N_49726);
or UO_3695 (O_3695,N_49527,N_49975);
or UO_3696 (O_3696,N_49628,N_49708);
nand UO_3697 (O_3697,N_49777,N_49976);
or UO_3698 (O_3698,N_49695,N_49852);
nor UO_3699 (O_3699,N_49722,N_49653);
and UO_3700 (O_3700,N_49644,N_49950);
xnor UO_3701 (O_3701,N_49600,N_49954);
nand UO_3702 (O_3702,N_49955,N_49983);
nand UO_3703 (O_3703,N_49618,N_49676);
or UO_3704 (O_3704,N_49996,N_49860);
and UO_3705 (O_3705,N_49757,N_49744);
nand UO_3706 (O_3706,N_49542,N_49872);
xnor UO_3707 (O_3707,N_49633,N_49637);
nand UO_3708 (O_3708,N_49942,N_49520);
xnor UO_3709 (O_3709,N_49598,N_49746);
xor UO_3710 (O_3710,N_49566,N_49564);
and UO_3711 (O_3711,N_49839,N_49627);
nand UO_3712 (O_3712,N_49880,N_49869);
and UO_3713 (O_3713,N_49589,N_49677);
nor UO_3714 (O_3714,N_49539,N_49927);
xor UO_3715 (O_3715,N_49961,N_49639);
nor UO_3716 (O_3716,N_49659,N_49690);
nor UO_3717 (O_3717,N_49741,N_49921);
xor UO_3718 (O_3718,N_49969,N_49575);
nand UO_3719 (O_3719,N_49753,N_49897);
and UO_3720 (O_3720,N_49753,N_49978);
nand UO_3721 (O_3721,N_49879,N_49958);
xor UO_3722 (O_3722,N_49825,N_49711);
nand UO_3723 (O_3723,N_49678,N_49939);
and UO_3724 (O_3724,N_49539,N_49545);
xor UO_3725 (O_3725,N_49802,N_49978);
nor UO_3726 (O_3726,N_49851,N_49875);
and UO_3727 (O_3727,N_49936,N_49542);
and UO_3728 (O_3728,N_49774,N_49861);
and UO_3729 (O_3729,N_49547,N_49755);
and UO_3730 (O_3730,N_49947,N_49675);
nor UO_3731 (O_3731,N_49782,N_49697);
or UO_3732 (O_3732,N_49689,N_49600);
nand UO_3733 (O_3733,N_49973,N_49524);
or UO_3734 (O_3734,N_49613,N_49511);
or UO_3735 (O_3735,N_49603,N_49801);
and UO_3736 (O_3736,N_49904,N_49759);
nor UO_3737 (O_3737,N_49974,N_49668);
nor UO_3738 (O_3738,N_49519,N_49973);
nor UO_3739 (O_3739,N_49870,N_49731);
and UO_3740 (O_3740,N_49500,N_49581);
or UO_3741 (O_3741,N_49593,N_49597);
xor UO_3742 (O_3742,N_49908,N_49745);
or UO_3743 (O_3743,N_49965,N_49956);
xnor UO_3744 (O_3744,N_49756,N_49585);
and UO_3745 (O_3745,N_49553,N_49953);
nand UO_3746 (O_3746,N_49597,N_49974);
nand UO_3747 (O_3747,N_49591,N_49858);
or UO_3748 (O_3748,N_49688,N_49929);
or UO_3749 (O_3749,N_49766,N_49678);
nand UO_3750 (O_3750,N_49822,N_49723);
or UO_3751 (O_3751,N_49678,N_49791);
nand UO_3752 (O_3752,N_49934,N_49542);
or UO_3753 (O_3753,N_49817,N_49850);
nor UO_3754 (O_3754,N_49514,N_49997);
nand UO_3755 (O_3755,N_49754,N_49618);
nor UO_3756 (O_3756,N_49695,N_49509);
or UO_3757 (O_3757,N_49931,N_49667);
nor UO_3758 (O_3758,N_49875,N_49518);
or UO_3759 (O_3759,N_49659,N_49727);
or UO_3760 (O_3760,N_49678,N_49728);
nand UO_3761 (O_3761,N_49861,N_49731);
xor UO_3762 (O_3762,N_49696,N_49536);
xor UO_3763 (O_3763,N_49730,N_49559);
nor UO_3764 (O_3764,N_49724,N_49946);
and UO_3765 (O_3765,N_49723,N_49518);
or UO_3766 (O_3766,N_49879,N_49579);
nor UO_3767 (O_3767,N_49866,N_49745);
and UO_3768 (O_3768,N_49813,N_49619);
and UO_3769 (O_3769,N_49689,N_49799);
and UO_3770 (O_3770,N_49668,N_49899);
xnor UO_3771 (O_3771,N_49502,N_49692);
or UO_3772 (O_3772,N_49736,N_49855);
xnor UO_3773 (O_3773,N_49743,N_49790);
xnor UO_3774 (O_3774,N_49658,N_49700);
nor UO_3775 (O_3775,N_49638,N_49907);
and UO_3776 (O_3776,N_49751,N_49685);
nand UO_3777 (O_3777,N_49648,N_49562);
and UO_3778 (O_3778,N_49505,N_49703);
nor UO_3779 (O_3779,N_49898,N_49974);
nand UO_3780 (O_3780,N_49693,N_49561);
or UO_3781 (O_3781,N_49953,N_49889);
nor UO_3782 (O_3782,N_49510,N_49634);
xnor UO_3783 (O_3783,N_49665,N_49904);
and UO_3784 (O_3784,N_49546,N_49911);
and UO_3785 (O_3785,N_49747,N_49523);
and UO_3786 (O_3786,N_49778,N_49517);
nand UO_3787 (O_3787,N_49532,N_49757);
nand UO_3788 (O_3788,N_49720,N_49583);
nand UO_3789 (O_3789,N_49946,N_49535);
nor UO_3790 (O_3790,N_49919,N_49724);
nor UO_3791 (O_3791,N_49694,N_49782);
nand UO_3792 (O_3792,N_49888,N_49936);
xnor UO_3793 (O_3793,N_49664,N_49671);
or UO_3794 (O_3794,N_49797,N_49805);
xnor UO_3795 (O_3795,N_49733,N_49870);
nand UO_3796 (O_3796,N_49616,N_49723);
xor UO_3797 (O_3797,N_49571,N_49780);
nor UO_3798 (O_3798,N_49790,N_49654);
nor UO_3799 (O_3799,N_49567,N_49604);
and UO_3800 (O_3800,N_49522,N_49649);
nor UO_3801 (O_3801,N_49959,N_49944);
or UO_3802 (O_3802,N_49627,N_49504);
nand UO_3803 (O_3803,N_49799,N_49581);
and UO_3804 (O_3804,N_49845,N_49656);
nor UO_3805 (O_3805,N_49905,N_49720);
and UO_3806 (O_3806,N_49880,N_49577);
or UO_3807 (O_3807,N_49633,N_49763);
nor UO_3808 (O_3808,N_49563,N_49737);
xnor UO_3809 (O_3809,N_49871,N_49878);
xnor UO_3810 (O_3810,N_49574,N_49572);
nand UO_3811 (O_3811,N_49890,N_49691);
and UO_3812 (O_3812,N_49590,N_49580);
nor UO_3813 (O_3813,N_49900,N_49963);
and UO_3814 (O_3814,N_49773,N_49796);
nor UO_3815 (O_3815,N_49951,N_49928);
and UO_3816 (O_3816,N_49663,N_49823);
or UO_3817 (O_3817,N_49618,N_49788);
nand UO_3818 (O_3818,N_49563,N_49979);
and UO_3819 (O_3819,N_49922,N_49882);
or UO_3820 (O_3820,N_49871,N_49679);
nor UO_3821 (O_3821,N_49504,N_49857);
xnor UO_3822 (O_3822,N_49665,N_49661);
and UO_3823 (O_3823,N_49879,N_49754);
nand UO_3824 (O_3824,N_49951,N_49684);
xor UO_3825 (O_3825,N_49507,N_49671);
and UO_3826 (O_3826,N_49745,N_49551);
nor UO_3827 (O_3827,N_49978,N_49796);
nand UO_3828 (O_3828,N_49745,N_49552);
and UO_3829 (O_3829,N_49863,N_49933);
and UO_3830 (O_3830,N_49955,N_49868);
and UO_3831 (O_3831,N_49915,N_49878);
nand UO_3832 (O_3832,N_49968,N_49875);
nor UO_3833 (O_3833,N_49527,N_49799);
nor UO_3834 (O_3834,N_49655,N_49851);
nor UO_3835 (O_3835,N_49512,N_49713);
and UO_3836 (O_3836,N_49597,N_49984);
xor UO_3837 (O_3837,N_49520,N_49825);
nand UO_3838 (O_3838,N_49977,N_49687);
or UO_3839 (O_3839,N_49940,N_49800);
and UO_3840 (O_3840,N_49517,N_49731);
xnor UO_3841 (O_3841,N_49939,N_49898);
nor UO_3842 (O_3842,N_49654,N_49989);
nor UO_3843 (O_3843,N_49813,N_49760);
nor UO_3844 (O_3844,N_49884,N_49991);
and UO_3845 (O_3845,N_49596,N_49735);
or UO_3846 (O_3846,N_49947,N_49825);
and UO_3847 (O_3847,N_49787,N_49754);
and UO_3848 (O_3848,N_49798,N_49634);
xor UO_3849 (O_3849,N_49740,N_49948);
nor UO_3850 (O_3850,N_49969,N_49824);
or UO_3851 (O_3851,N_49688,N_49767);
nor UO_3852 (O_3852,N_49807,N_49604);
nor UO_3853 (O_3853,N_49625,N_49542);
or UO_3854 (O_3854,N_49983,N_49749);
nand UO_3855 (O_3855,N_49666,N_49783);
nand UO_3856 (O_3856,N_49536,N_49578);
nand UO_3857 (O_3857,N_49758,N_49759);
or UO_3858 (O_3858,N_49712,N_49515);
or UO_3859 (O_3859,N_49706,N_49523);
and UO_3860 (O_3860,N_49937,N_49564);
xnor UO_3861 (O_3861,N_49940,N_49874);
nor UO_3862 (O_3862,N_49607,N_49553);
nand UO_3863 (O_3863,N_49707,N_49595);
or UO_3864 (O_3864,N_49719,N_49807);
xor UO_3865 (O_3865,N_49648,N_49722);
and UO_3866 (O_3866,N_49785,N_49848);
and UO_3867 (O_3867,N_49816,N_49857);
xor UO_3868 (O_3868,N_49902,N_49666);
or UO_3869 (O_3869,N_49725,N_49773);
nor UO_3870 (O_3870,N_49680,N_49794);
nand UO_3871 (O_3871,N_49770,N_49906);
nor UO_3872 (O_3872,N_49652,N_49621);
or UO_3873 (O_3873,N_49781,N_49636);
nand UO_3874 (O_3874,N_49935,N_49610);
and UO_3875 (O_3875,N_49917,N_49770);
or UO_3876 (O_3876,N_49651,N_49952);
or UO_3877 (O_3877,N_49707,N_49823);
and UO_3878 (O_3878,N_49761,N_49546);
nor UO_3879 (O_3879,N_49647,N_49691);
and UO_3880 (O_3880,N_49546,N_49656);
xor UO_3881 (O_3881,N_49682,N_49760);
xnor UO_3882 (O_3882,N_49553,N_49852);
xor UO_3883 (O_3883,N_49734,N_49779);
or UO_3884 (O_3884,N_49980,N_49680);
nor UO_3885 (O_3885,N_49646,N_49921);
and UO_3886 (O_3886,N_49509,N_49750);
xnor UO_3887 (O_3887,N_49595,N_49690);
nand UO_3888 (O_3888,N_49834,N_49956);
and UO_3889 (O_3889,N_49962,N_49661);
xnor UO_3890 (O_3890,N_49976,N_49566);
and UO_3891 (O_3891,N_49995,N_49565);
or UO_3892 (O_3892,N_49842,N_49882);
and UO_3893 (O_3893,N_49986,N_49552);
nand UO_3894 (O_3894,N_49921,N_49578);
nor UO_3895 (O_3895,N_49919,N_49828);
and UO_3896 (O_3896,N_49909,N_49786);
or UO_3897 (O_3897,N_49618,N_49636);
nand UO_3898 (O_3898,N_49674,N_49524);
xnor UO_3899 (O_3899,N_49999,N_49807);
or UO_3900 (O_3900,N_49892,N_49868);
nand UO_3901 (O_3901,N_49936,N_49580);
xnor UO_3902 (O_3902,N_49590,N_49886);
nand UO_3903 (O_3903,N_49942,N_49930);
nand UO_3904 (O_3904,N_49777,N_49838);
xor UO_3905 (O_3905,N_49732,N_49816);
nor UO_3906 (O_3906,N_49879,N_49833);
or UO_3907 (O_3907,N_49879,N_49631);
nand UO_3908 (O_3908,N_49880,N_49760);
and UO_3909 (O_3909,N_49920,N_49835);
or UO_3910 (O_3910,N_49594,N_49841);
xor UO_3911 (O_3911,N_49885,N_49558);
nor UO_3912 (O_3912,N_49887,N_49570);
nand UO_3913 (O_3913,N_49625,N_49688);
or UO_3914 (O_3914,N_49528,N_49785);
nand UO_3915 (O_3915,N_49527,N_49568);
nand UO_3916 (O_3916,N_49785,N_49669);
nor UO_3917 (O_3917,N_49531,N_49731);
nand UO_3918 (O_3918,N_49964,N_49806);
xor UO_3919 (O_3919,N_49825,N_49521);
nor UO_3920 (O_3920,N_49876,N_49722);
or UO_3921 (O_3921,N_49548,N_49874);
nand UO_3922 (O_3922,N_49789,N_49733);
and UO_3923 (O_3923,N_49928,N_49550);
nor UO_3924 (O_3924,N_49679,N_49761);
or UO_3925 (O_3925,N_49926,N_49888);
or UO_3926 (O_3926,N_49803,N_49668);
and UO_3927 (O_3927,N_49579,N_49876);
xor UO_3928 (O_3928,N_49951,N_49799);
nor UO_3929 (O_3929,N_49970,N_49781);
xor UO_3930 (O_3930,N_49792,N_49929);
xnor UO_3931 (O_3931,N_49717,N_49886);
xor UO_3932 (O_3932,N_49523,N_49915);
nand UO_3933 (O_3933,N_49807,N_49892);
nor UO_3934 (O_3934,N_49766,N_49762);
nand UO_3935 (O_3935,N_49757,N_49557);
and UO_3936 (O_3936,N_49987,N_49903);
and UO_3937 (O_3937,N_49671,N_49546);
nand UO_3938 (O_3938,N_49844,N_49760);
nand UO_3939 (O_3939,N_49528,N_49797);
xnor UO_3940 (O_3940,N_49605,N_49549);
and UO_3941 (O_3941,N_49856,N_49580);
nand UO_3942 (O_3942,N_49625,N_49589);
and UO_3943 (O_3943,N_49771,N_49902);
and UO_3944 (O_3944,N_49696,N_49726);
nand UO_3945 (O_3945,N_49575,N_49986);
xnor UO_3946 (O_3946,N_49566,N_49887);
or UO_3947 (O_3947,N_49710,N_49616);
nor UO_3948 (O_3948,N_49500,N_49627);
xnor UO_3949 (O_3949,N_49577,N_49592);
nor UO_3950 (O_3950,N_49933,N_49779);
xnor UO_3951 (O_3951,N_49985,N_49569);
xnor UO_3952 (O_3952,N_49747,N_49765);
and UO_3953 (O_3953,N_49640,N_49939);
or UO_3954 (O_3954,N_49656,N_49748);
xnor UO_3955 (O_3955,N_49773,N_49899);
nor UO_3956 (O_3956,N_49712,N_49908);
nand UO_3957 (O_3957,N_49834,N_49741);
or UO_3958 (O_3958,N_49900,N_49836);
nand UO_3959 (O_3959,N_49633,N_49943);
nand UO_3960 (O_3960,N_49945,N_49807);
nand UO_3961 (O_3961,N_49740,N_49826);
nand UO_3962 (O_3962,N_49872,N_49945);
and UO_3963 (O_3963,N_49908,N_49791);
xor UO_3964 (O_3964,N_49736,N_49777);
nand UO_3965 (O_3965,N_49537,N_49788);
and UO_3966 (O_3966,N_49911,N_49858);
xor UO_3967 (O_3967,N_49908,N_49884);
and UO_3968 (O_3968,N_49987,N_49799);
or UO_3969 (O_3969,N_49567,N_49935);
nand UO_3970 (O_3970,N_49584,N_49549);
xnor UO_3971 (O_3971,N_49859,N_49552);
or UO_3972 (O_3972,N_49522,N_49526);
or UO_3973 (O_3973,N_49887,N_49676);
nand UO_3974 (O_3974,N_49501,N_49796);
nand UO_3975 (O_3975,N_49648,N_49974);
nand UO_3976 (O_3976,N_49511,N_49732);
xnor UO_3977 (O_3977,N_49971,N_49890);
nand UO_3978 (O_3978,N_49882,N_49824);
xor UO_3979 (O_3979,N_49574,N_49605);
or UO_3980 (O_3980,N_49922,N_49704);
and UO_3981 (O_3981,N_49526,N_49555);
nand UO_3982 (O_3982,N_49792,N_49927);
nor UO_3983 (O_3983,N_49899,N_49810);
nand UO_3984 (O_3984,N_49990,N_49732);
xnor UO_3985 (O_3985,N_49965,N_49680);
and UO_3986 (O_3986,N_49993,N_49999);
and UO_3987 (O_3987,N_49657,N_49787);
xnor UO_3988 (O_3988,N_49928,N_49909);
xnor UO_3989 (O_3989,N_49983,N_49950);
nand UO_3990 (O_3990,N_49715,N_49661);
and UO_3991 (O_3991,N_49563,N_49774);
nand UO_3992 (O_3992,N_49892,N_49602);
nand UO_3993 (O_3993,N_49831,N_49957);
nand UO_3994 (O_3994,N_49721,N_49736);
nor UO_3995 (O_3995,N_49518,N_49551);
and UO_3996 (O_3996,N_49965,N_49504);
or UO_3997 (O_3997,N_49633,N_49925);
or UO_3998 (O_3998,N_49754,N_49627);
xor UO_3999 (O_3999,N_49734,N_49663);
nand UO_4000 (O_4000,N_49796,N_49546);
nor UO_4001 (O_4001,N_49508,N_49955);
and UO_4002 (O_4002,N_49994,N_49603);
nand UO_4003 (O_4003,N_49942,N_49994);
and UO_4004 (O_4004,N_49849,N_49983);
and UO_4005 (O_4005,N_49568,N_49657);
xor UO_4006 (O_4006,N_49596,N_49613);
xor UO_4007 (O_4007,N_49765,N_49647);
and UO_4008 (O_4008,N_49761,N_49937);
and UO_4009 (O_4009,N_49971,N_49760);
and UO_4010 (O_4010,N_49529,N_49506);
and UO_4011 (O_4011,N_49775,N_49577);
and UO_4012 (O_4012,N_49662,N_49504);
nand UO_4013 (O_4013,N_49746,N_49653);
nand UO_4014 (O_4014,N_49682,N_49549);
or UO_4015 (O_4015,N_49815,N_49635);
and UO_4016 (O_4016,N_49565,N_49728);
or UO_4017 (O_4017,N_49720,N_49672);
nand UO_4018 (O_4018,N_49769,N_49994);
xor UO_4019 (O_4019,N_49576,N_49793);
xnor UO_4020 (O_4020,N_49926,N_49651);
or UO_4021 (O_4021,N_49546,N_49767);
nor UO_4022 (O_4022,N_49610,N_49873);
and UO_4023 (O_4023,N_49886,N_49769);
xnor UO_4024 (O_4024,N_49850,N_49626);
nor UO_4025 (O_4025,N_49655,N_49949);
or UO_4026 (O_4026,N_49774,N_49866);
nand UO_4027 (O_4027,N_49510,N_49959);
nand UO_4028 (O_4028,N_49988,N_49962);
and UO_4029 (O_4029,N_49532,N_49973);
or UO_4030 (O_4030,N_49763,N_49591);
nor UO_4031 (O_4031,N_49633,N_49798);
and UO_4032 (O_4032,N_49774,N_49717);
nor UO_4033 (O_4033,N_49511,N_49713);
nand UO_4034 (O_4034,N_49918,N_49571);
nand UO_4035 (O_4035,N_49705,N_49711);
nand UO_4036 (O_4036,N_49815,N_49667);
or UO_4037 (O_4037,N_49631,N_49508);
nor UO_4038 (O_4038,N_49978,N_49677);
or UO_4039 (O_4039,N_49644,N_49682);
and UO_4040 (O_4040,N_49523,N_49877);
xor UO_4041 (O_4041,N_49599,N_49587);
xnor UO_4042 (O_4042,N_49922,N_49682);
nor UO_4043 (O_4043,N_49947,N_49501);
xnor UO_4044 (O_4044,N_49855,N_49816);
and UO_4045 (O_4045,N_49997,N_49604);
xnor UO_4046 (O_4046,N_49936,N_49606);
and UO_4047 (O_4047,N_49692,N_49962);
or UO_4048 (O_4048,N_49557,N_49617);
and UO_4049 (O_4049,N_49596,N_49643);
xnor UO_4050 (O_4050,N_49563,N_49530);
and UO_4051 (O_4051,N_49533,N_49632);
nor UO_4052 (O_4052,N_49979,N_49929);
nand UO_4053 (O_4053,N_49514,N_49930);
xnor UO_4054 (O_4054,N_49571,N_49568);
and UO_4055 (O_4055,N_49793,N_49851);
nor UO_4056 (O_4056,N_49614,N_49808);
nor UO_4057 (O_4057,N_49972,N_49668);
and UO_4058 (O_4058,N_49595,N_49643);
nand UO_4059 (O_4059,N_49695,N_49691);
nand UO_4060 (O_4060,N_49814,N_49589);
nor UO_4061 (O_4061,N_49559,N_49766);
xor UO_4062 (O_4062,N_49566,N_49741);
nor UO_4063 (O_4063,N_49681,N_49994);
or UO_4064 (O_4064,N_49895,N_49898);
xor UO_4065 (O_4065,N_49916,N_49964);
and UO_4066 (O_4066,N_49605,N_49561);
nand UO_4067 (O_4067,N_49642,N_49895);
nand UO_4068 (O_4068,N_49683,N_49815);
nand UO_4069 (O_4069,N_49850,N_49544);
nor UO_4070 (O_4070,N_49997,N_49563);
xor UO_4071 (O_4071,N_49813,N_49508);
xnor UO_4072 (O_4072,N_49528,N_49805);
or UO_4073 (O_4073,N_49937,N_49756);
or UO_4074 (O_4074,N_49680,N_49894);
nand UO_4075 (O_4075,N_49664,N_49600);
or UO_4076 (O_4076,N_49838,N_49794);
nand UO_4077 (O_4077,N_49957,N_49877);
nor UO_4078 (O_4078,N_49892,N_49784);
or UO_4079 (O_4079,N_49694,N_49624);
xnor UO_4080 (O_4080,N_49864,N_49533);
or UO_4081 (O_4081,N_49884,N_49714);
xor UO_4082 (O_4082,N_49637,N_49680);
xor UO_4083 (O_4083,N_49820,N_49656);
or UO_4084 (O_4084,N_49837,N_49757);
and UO_4085 (O_4085,N_49511,N_49567);
nor UO_4086 (O_4086,N_49628,N_49928);
nor UO_4087 (O_4087,N_49878,N_49896);
or UO_4088 (O_4088,N_49880,N_49635);
nand UO_4089 (O_4089,N_49715,N_49510);
and UO_4090 (O_4090,N_49889,N_49723);
xor UO_4091 (O_4091,N_49865,N_49863);
nor UO_4092 (O_4092,N_49971,N_49618);
nand UO_4093 (O_4093,N_49766,N_49815);
nand UO_4094 (O_4094,N_49655,N_49866);
and UO_4095 (O_4095,N_49811,N_49958);
nor UO_4096 (O_4096,N_49832,N_49957);
and UO_4097 (O_4097,N_49507,N_49960);
xor UO_4098 (O_4098,N_49788,N_49592);
and UO_4099 (O_4099,N_49923,N_49779);
or UO_4100 (O_4100,N_49855,N_49803);
nand UO_4101 (O_4101,N_49661,N_49836);
nor UO_4102 (O_4102,N_49550,N_49591);
or UO_4103 (O_4103,N_49809,N_49630);
or UO_4104 (O_4104,N_49984,N_49775);
or UO_4105 (O_4105,N_49783,N_49506);
and UO_4106 (O_4106,N_49862,N_49592);
nor UO_4107 (O_4107,N_49775,N_49861);
and UO_4108 (O_4108,N_49957,N_49669);
xor UO_4109 (O_4109,N_49705,N_49736);
nand UO_4110 (O_4110,N_49607,N_49846);
nand UO_4111 (O_4111,N_49963,N_49543);
xnor UO_4112 (O_4112,N_49843,N_49661);
or UO_4113 (O_4113,N_49717,N_49722);
nor UO_4114 (O_4114,N_49849,N_49685);
xor UO_4115 (O_4115,N_49927,N_49939);
and UO_4116 (O_4116,N_49563,N_49521);
or UO_4117 (O_4117,N_49550,N_49772);
or UO_4118 (O_4118,N_49555,N_49673);
and UO_4119 (O_4119,N_49677,N_49839);
or UO_4120 (O_4120,N_49921,N_49506);
nand UO_4121 (O_4121,N_49553,N_49537);
xor UO_4122 (O_4122,N_49955,N_49587);
or UO_4123 (O_4123,N_49860,N_49689);
or UO_4124 (O_4124,N_49572,N_49837);
and UO_4125 (O_4125,N_49654,N_49500);
xnor UO_4126 (O_4126,N_49646,N_49524);
nand UO_4127 (O_4127,N_49999,N_49942);
nor UO_4128 (O_4128,N_49660,N_49805);
xnor UO_4129 (O_4129,N_49567,N_49607);
or UO_4130 (O_4130,N_49574,N_49558);
and UO_4131 (O_4131,N_49711,N_49999);
nor UO_4132 (O_4132,N_49742,N_49930);
xnor UO_4133 (O_4133,N_49752,N_49822);
nor UO_4134 (O_4134,N_49513,N_49855);
nand UO_4135 (O_4135,N_49963,N_49802);
and UO_4136 (O_4136,N_49550,N_49909);
and UO_4137 (O_4137,N_49996,N_49933);
or UO_4138 (O_4138,N_49687,N_49701);
nor UO_4139 (O_4139,N_49965,N_49865);
nor UO_4140 (O_4140,N_49513,N_49509);
or UO_4141 (O_4141,N_49862,N_49548);
nand UO_4142 (O_4142,N_49786,N_49514);
and UO_4143 (O_4143,N_49868,N_49620);
nand UO_4144 (O_4144,N_49652,N_49665);
or UO_4145 (O_4145,N_49893,N_49977);
nor UO_4146 (O_4146,N_49706,N_49532);
and UO_4147 (O_4147,N_49578,N_49694);
and UO_4148 (O_4148,N_49556,N_49763);
xnor UO_4149 (O_4149,N_49609,N_49779);
and UO_4150 (O_4150,N_49554,N_49995);
nand UO_4151 (O_4151,N_49605,N_49683);
nand UO_4152 (O_4152,N_49696,N_49911);
or UO_4153 (O_4153,N_49798,N_49906);
nor UO_4154 (O_4154,N_49723,N_49689);
nor UO_4155 (O_4155,N_49628,N_49707);
nand UO_4156 (O_4156,N_49674,N_49734);
nand UO_4157 (O_4157,N_49919,N_49662);
xor UO_4158 (O_4158,N_49830,N_49572);
nand UO_4159 (O_4159,N_49752,N_49537);
and UO_4160 (O_4160,N_49754,N_49520);
and UO_4161 (O_4161,N_49929,N_49602);
nand UO_4162 (O_4162,N_49952,N_49529);
or UO_4163 (O_4163,N_49990,N_49516);
or UO_4164 (O_4164,N_49955,N_49887);
xor UO_4165 (O_4165,N_49822,N_49941);
xnor UO_4166 (O_4166,N_49937,N_49642);
xor UO_4167 (O_4167,N_49638,N_49794);
nor UO_4168 (O_4168,N_49568,N_49885);
or UO_4169 (O_4169,N_49898,N_49891);
and UO_4170 (O_4170,N_49519,N_49903);
xnor UO_4171 (O_4171,N_49533,N_49959);
xnor UO_4172 (O_4172,N_49539,N_49960);
nor UO_4173 (O_4173,N_49925,N_49748);
nand UO_4174 (O_4174,N_49872,N_49810);
nor UO_4175 (O_4175,N_49659,N_49506);
nor UO_4176 (O_4176,N_49545,N_49942);
nor UO_4177 (O_4177,N_49664,N_49602);
or UO_4178 (O_4178,N_49701,N_49631);
nand UO_4179 (O_4179,N_49741,N_49829);
nand UO_4180 (O_4180,N_49713,N_49732);
and UO_4181 (O_4181,N_49639,N_49734);
nor UO_4182 (O_4182,N_49933,N_49546);
nand UO_4183 (O_4183,N_49873,N_49931);
and UO_4184 (O_4184,N_49866,N_49824);
or UO_4185 (O_4185,N_49934,N_49787);
or UO_4186 (O_4186,N_49998,N_49584);
and UO_4187 (O_4187,N_49850,N_49570);
and UO_4188 (O_4188,N_49589,N_49952);
nor UO_4189 (O_4189,N_49877,N_49539);
xor UO_4190 (O_4190,N_49510,N_49631);
or UO_4191 (O_4191,N_49826,N_49945);
xnor UO_4192 (O_4192,N_49943,N_49762);
xor UO_4193 (O_4193,N_49760,N_49757);
nand UO_4194 (O_4194,N_49813,N_49909);
nand UO_4195 (O_4195,N_49594,N_49825);
nand UO_4196 (O_4196,N_49808,N_49743);
nand UO_4197 (O_4197,N_49951,N_49793);
xnor UO_4198 (O_4198,N_49750,N_49650);
nand UO_4199 (O_4199,N_49735,N_49971);
nor UO_4200 (O_4200,N_49667,N_49519);
or UO_4201 (O_4201,N_49514,N_49763);
nor UO_4202 (O_4202,N_49799,N_49645);
nor UO_4203 (O_4203,N_49740,N_49997);
or UO_4204 (O_4204,N_49853,N_49517);
or UO_4205 (O_4205,N_49941,N_49851);
and UO_4206 (O_4206,N_49812,N_49843);
and UO_4207 (O_4207,N_49927,N_49621);
or UO_4208 (O_4208,N_49833,N_49838);
or UO_4209 (O_4209,N_49559,N_49828);
nand UO_4210 (O_4210,N_49770,N_49809);
or UO_4211 (O_4211,N_49790,N_49993);
or UO_4212 (O_4212,N_49695,N_49898);
or UO_4213 (O_4213,N_49932,N_49651);
and UO_4214 (O_4214,N_49770,N_49782);
nand UO_4215 (O_4215,N_49682,N_49591);
xnor UO_4216 (O_4216,N_49781,N_49807);
or UO_4217 (O_4217,N_49917,N_49992);
nor UO_4218 (O_4218,N_49847,N_49536);
nand UO_4219 (O_4219,N_49678,N_49945);
nor UO_4220 (O_4220,N_49578,N_49775);
nand UO_4221 (O_4221,N_49830,N_49968);
and UO_4222 (O_4222,N_49503,N_49699);
nand UO_4223 (O_4223,N_49922,N_49658);
nand UO_4224 (O_4224,N_49913,N_49787);
and UO_4225 (O_4225,N_49859,N_49747);
or UO_4226 (O_4226,N_49742,N_49855);
and UO_4227 (O_4227,N_49556,N_49788);
nor UO_4228 (O_4228,N_49837,N_49842);
nor UO_4229 (O_4229,N_49750,N_49801);
nor UO_4230 (O_4230,N_49785,N_49653);
xnor UO_4231 (O_4231,N_49964,N_49950);
nand UO_4232 (O_4232,N_49838,N_49613);
or UO_4233 (O_4233,N_49658,N_49607);
or UO_4234 (O_4234,N_49799,N_49657);
and UO_4235 (O_4235,N_49935,N_49750);
nor UO_4236 (O_4236,N_49569,N_49760);
nand UO_4237 (O_4237,N_49653,N_49669);
nand UO_4238 (O_4238,N_49517,N_49795);
or UO_4239 (O_4239,N_49814,N_49744);
xor UO_4240 (O_4240,N_49751,N_49853);
xor UO_4241 (O_4241,N_49893,N_49959);
and UO_4242 (O_4242,N_49569,N_49731);
and UO_4243 (O_4243,N_49650,N_49595);
nand UO_4244 (O_4244,N_49785,N_49846);
nor UO_4245 (O_4245,N_49591,N_49913);
nand UO_4246 (O_4246,N_49712,N_49974);
xor UO_4247 (O_4247,N_49805,N_49690);
nor UO_4248 (O_4248,N_49955,N_49903);
nor UO_4249 (O_4249,N_49724,N_49953);
nand UO_4250 (O_4250,N_49780,N_49880);
and UO_4251 (O_4251,N_49845,N_49534);
or UO_4252 (O_4252,N_49828,N_49927);
xor UO_4253 (O_4253,N_49679,N_49506);
nand UO_4254 (O_4254,N_49671,N_49810);
nor UO_4255 (O_4255,N_49524,N_49783);
xor UO_4256 (O_4256,N_49841,N_49729);
xnor UO_4257 (O_4257,N_49953,N_49646);
nor UO_4258 (O_4258,N_49632,N_49843);
and UO_4259 (O_4259,N_49758,N_49969);
or UO_4260 (O_4260,N_49792,N_49881);
nor UO_4261 (O_4261,N_49805,N_49510);
xor UO_4262 (O_4262,N_49934,N_49928);
xnor UO_4263 (O_4263,N_49970,N_49669);
or UO_4264 (O_4264,N_49867,N_49900);
or UO_4265 (O_4265,N_49527,N_49907);
or UO_4266 (O_4266,N_49781,N_49669);
nor UO_4267 (O_4267,N_49646,N_49958);
or UO_4268 (O_4268,N_49721,N_49755);
and UO_4269 (O_4269,N_49945,N_49529);
nor UO_4270 (O_4270,N_49976,N_49578);
nor UO_4271 (O_4271,N_49611,N_49734);
nor UO_4272 (O_4272,N_49985,N_49746);
or UO_4273 (O_4273,N_49656,N_49902);
nor UO_4274 (O_4274,N_49626,N_49975);
and UO_4275 (O_4275,N_49597,N_49894);
and UO_4276 (O_4276,N_49532,N_49917);
or UO_4277 (O_4277,N_49683,N_49787);
nor UO_4278 (O_4278,N_49589,N_49645);
nand UO_4279 (O_4279,N_49887,N_49990);
and UO_4280 (O_4280,N_49602,N_49935);
and UO_4281 (O_4281,N_49506,N_49752);
and UO_4282 (O_4282,N_49831,N_49506);
nand UO_4283 (O_4283,N_49822,N_49908);
and UO_4284 (O_4284,N_49671,N_49768);
or UO_4285 (O_4285,N_49613,N_49782);
and UO_4286 (O_4286,N_49617,N_49727);
xor UO_4287 (O_4287,N_49535,N_49922);
or UO_4288 (O_4288,N_49638,N_49648);
or UO_4289 (O_4289,N_49506,N_49760);
nand UO_4290 (O_4290,N_49819,N_49526);
nand UO_4291 (O_4291,N_49996,N_49891);
nor UO_4292 (O_4292,N_49720,N_49880);
nand UO_4293 (O_4293,N_49643,N_49804);
nand UO_4294 (O_4294,N_49653,N_49745);
nand UO_4295 (O_4295,N_49662,N_49881);
nor UO_4296 (O_4296,N_49640,N_49884);
and UO_4297 (O_4297,N_49823,N_49729);
nor UO_4298 (O_4298,N_49797,N_49514);
and UO_4299 (O_4299,N_49859,N_49829);
xor UO_4300 (O_4300,N_49632,N_49700);
nor UO_4301 (O_4301,N_49598,N_49754);
xor UO_4302 (O_4302,N_49744,N_49708);
or UO_4303 (O_4303,N_49625,N_49853);
or UO_4304 (O_4304,N_49764,N_49962);
nand UO_4305 (O_4305,N_49810,N_49943);
nor UO_4306 (O_4306,N_49757,N_49508);
nor UO_4307 (O_4307,N_49820,N_49888);
xnor UO_4308 (O_4308,N_49931,N_49514);
nand UO_4309 (O_4309,N_49753,N_49999);
or UO_4310 (O_4310,N_49720,N_49704);
nand UO_4311 (O_4311,N_49706,N_49655);
nand UO_4312 (O_4312,N_49919,N_49818);
or UO_4313 (O_4313,N_49733,N_49805);
nor UO_4314 (O_4314,N_49720,N_49846);
nand UO_4315 (O_4315,N_49682,N_49732);
nor UO_4316 (O_4316,N_49851,N_49739);
and UO_4317 (O_4317,N_49973,N_49501);
or UO_4318 (O_4318,N_49528,N_49515);
nand UO_4319 (O_4319,N_49984,N_49893);
nand UO_4320 (O_4320,N_49975,N_49653);
and UO_4321 (O_4321,N_49844,N_49713);
and UO_4322 (O_4322,N_49848,N_49536);
nand UO_4323 (O_4323,N_49583,N_49872);
nor UO_4324 (O_4324,N_49592,N_49815);
or UO_4325 (O_4325,N_49618,N_49956);
and UO_4326 (O_4326,N_49588,N_49662);
nor UO_4327 (O_4327,N_49506,N_49722);
or UO_4328 (O_4328,N_49554,N_49705);
nand UO_4329 (O_4329,N_49858,N_49906);
nor UO_4330 (O_4330,N_49636,N_49504);
nand UO_4331 (O_4331,N_49978,N_49723);
and UO_4332 (O_4332,N_49988,N_49704);
nor UO_4333 (O_4333,N_49874,N_49542);
or UO_4334 (O_4334,N_49997,N_49749);
or UO_4335 (O_4335,N_49878,N_49963);
nand UO_4336 (O_4336,N_49933,N_49830);
or UO_4337 (O_4337,N_49867,N_49748);
and UO_4338 (O_4338,N_49998,N_49532);
nand UO_4339 (O_4339,N_49706,N_49588);
or UO_4340 (O_4340,N_49635,N_49683);
and UO_4341 (O_4341,N_49833,N_49786);
xor UO_4342 (O_4342,N_49852,N_49679);
nand UO_4343 (O_4343,N_49691,N_49877);
or UO_4344 (O_4344,N_49867,N_49717);
and UO_4345 (O_4345,N_49867,N_49573);
and UO_4346 (O_4346,N_49574,N_49847);
nand UO_4347 (O_4347,N_49641,N_49687);
xnor UO_4348 (O_4348,N_49622,N_49653);
xor UO_4349 (O_4349,N_49716,N_49646);
nor UO_4350 (O_4350,N_49691,N_49950);
or UO_4351 (O_4351,N_49922,N_49780);
and UO_4352 (O_4352,N_49572,N_49829);
nor UO_4353 (O_4353,N_49899,N_49609);
nand UO_4354 (O_4354,N_49835,N_49605);
or UO_4355 (O_4355,N_49543,N_49688);
or UO_4356 (O_4356,N_49952,N_49966);
nor UO_4357 (O_4357,N_49606,N_49510);
xor UO_4358 (O_4358,N_49617,N_49933);
or UO_4359 (O_4359,N_49896,N_49856);
nor UO_4360 (O_4360,N_49636,N_49696);
or UO_4361 (O_4361,N_49776,N_49605);
nand UO_4362 (O_4362,N_49843,N_49939);
and UO_4363 (O_4363,N_49963,N_49509);
and UO_4364 (O_4364,N_49809,N_49832);
nor UO_4365 (O_4365,N_49760,N_49642);
and UO_4366 (O_4366,N_49583,N_49833);
or UO_4367 (O_4367,N_49850,N_49931);
nor UO_4368 (O_4368,N_49978,N_49820);
nand UO_4369 (O_4369,N_49697,N_49885);
xor UO_4370 (O_4370,N_49951,N_49917);
xor UO_4371 (O_4371,N_49695,N_49513);
or UO_4372 (O_4372,N_49813,N_49617);
xnor UO_4373 (O_4373,N_49985,N_49663);
nand UO_4374 (O_4374,N_49953,N_49894);
nand UO_4375 (O_4375,N_49797,N_49861);
xor UO_4376 (O_4376,N_49500,N_49668);
xnor UO_4377 (O_4377,N_49716,N_49595);
or UO_4378 (O_4378,N_49727,N_49578);
and UO_4379 (O_4379,N_49952,N_49616);
and UO_4380 (O_4380,N_49901,N_49983);
nor UO_4381 (O_4381,N_49686,N_49858);
xnor UO_4382 (O_4382,N_49770,N_49850);
nor UO_4383 (O_4383,N_49767,N_49987);
nor UO_4384 (O_4384,N_49851,N_49708);
xor UO_4385 (O_4385,N_49779,N_49520);
xor UO_4386 (O_4386,N_49958,N_49560);
or UO_4387 (O_4387,N_49663,N_49511);
xnor UO_4388 (O_4388,N_49712,N_49941);
or UO_4389 (O_4389,N_49570,N_49507);
nor UO_4390 (O_4390,N_49612,N_49602);
xnor UO_4391 (O_4391,N_49548,N_49839);
and UO_4392 (O_4392,N_49976,N_49532);
or UO_4393 (O_4393,N_49520,N_49920);
nand UO_4394 (O_4394,N_49601,N_49991);
or UO_4395 (O_4395,N_49970,N_49914);
nor UO_4396 (O_4396,N_49681,N_49692);
nor UO_4397 (O_4397,N_49761,N_49563);
xnor UO_4398 (O_4398,N_49991,N_49945);
and UO_4399 (O_4399,N_49991,N_49658);
nor UO_4400 (O_4400,N_49812,N_49769);
nand UO_4401 (O_4401,N_49980,N_49712);
or UO_4402 (O_4402,N_49751,N_49607);
xor UO_4403 (O_4403,N_49531,N_49679);
nand UO_4404 (O_4404,N_49952,N_49957);
xnor UO_4405 (O_4405,N_49941,N_49720);
and UO_4406 (O_4406,N_49551,N_49959);
xor UO_4407 (O_4407,N_49520,N_49510);
xnor UO_4408 (O_4408,N_49973,N_49810);
xor UO_4409 (O_4409,N_49560,N_49989);
nand UO_4410 (O_4410,N_49690,N_49982);
nand UO_4411 (O_4411,N_49621,N_49501);
and UO_4412 (O_4412,N_49772,N_49589);
nor UO_4413 (O_4413,N_49606,N_49924);
and UO_4414 (O_4414,N_49840,N_49560);
and UO_4415 (O_4415,N_49514,N_49785);
xor UO_4416 (O_4416,N_49584,N_49784);
xnor UO_4417 (O_4417,N_49698,N_49520);
or UO_4418 (O_4418,N_49644,N_49919);
xor UO_4419 (O_4419,N_49780,N_49566);
nor UO_4420 (O_4420,N_49530,N_49899);
nand UO_4421 (O_4421,N_49542,N_49646);
nor UO_4422 (O_4422,N_49955,N_49734);
or UO_4423 (O_4423,N_49896,N_49660);
or UO_4424 (O_4424,N_49733,N_49524);
nor UO_4425 (O_4425,N_49743,N_49546);
xor UO_4426 (O_4426,N_49584,N_49557);
nor UO_4427 (O_4427,N_49565,N_49645);
and UO_4428 (O_4428,N_49717,N_49710);
xor UO_4429 (O_4429,N_49507,N_49513);
xnor UO_4430 (O_4430,N_49761,N_49946);
nor UO_4431 (O_4431,N_49821,N_49584);
xnor UO_4432 (O_4432,N_49784,N_49703);
xnor UO_4433 (O_4433,N_49647,N_49800);
nor UO_4434 (O_4434,N_49830,N_49536);
and UO_4435 (O_4435,N_49675,N_49536);
or UO_4436 (O_4436,N_49646,N_49500);
or UO_4437 (O_4437,N_49781,N_49769);
nand UO_4438 (O_4438,N_49593,N_49874);
nor UO_4439 (O_4439,N_49605,N_49741);
and UO_4440 (O_4440,N_49967,N_49685);
or UO_4441 (O_4441,N_49634,N_49952);
nand UO_4442 (O_4442,N_49639,N_49588);
and UO_4443 (O_4443,N_49678,N_49542);
xnor UO_4444 (O_4444,N_49561,N_49924);
or UO_4445 (O_4445,N_49925,N_49793);
or UO_4446 (O_4446,N_49713,N_49904);
nand UO_4447 (O_4447,N_49640,N_49991);
and UO_4448 (O_4448,N_49638,N_49900);
xnor UO_4449 (O_4449,N_49631,N_49985);
xnor UO_4450 (O_4450,N_49887,N_49606);
and UO_4451 (O_4451,N_49923,N_49631);
xor UO_4452 (O_4452,N_49920,N_49674);
and UO_4453 (O_4453,N_49623,N_49755);
and UO_4454 (O_4454,N_49534,N_49678);
and UO_4455 (O_4455,N_49540,N_49847);
or UO_4456 (O_4456,N_49522,N_49672);
or UO_4457 (O_4457,N_49855,N_49909);
nor UO_4458 (O_4458,N_49765,N_49895);
nor UO_4459 (O_4459,N_49695,N_49862);
nand UO_4460 (O_4460,N_49540,N_49822);
or UO_4461 (O_4461,N_49938,N_49926);
nand UO_4462 (O_4462,N_49909,N_49600);
xnor UO_4463 (O_4463,N_49790,N_49960);
nand UO_4464 (O_4464,N_49905,N_49638);
and UO_4465 (O_4465,N_49653,N_49613);
nand UO_4466 (O_4466,N_49755,N_49756);
and UO_4467 (O_4467,N_49578,N_49502);
nand UO_4468 (O_4468,N_49722,N_49990);
or UO_4469 (O_4469,N_49714,N_49661);
nor UO_4470 (O_4470,N_49876,N_49526);
xor UO_4471 (O_4471,N_49672,N_49936);
xor UO_4472 (O_4472,N_49588,N_49848);
or UO_4473 (O_4473,N_49555,N_49939);
nand UO_4474 (O_4474,N_49900,N_49711);
or UO_4475 (O_4475,N_49887,N_49615);
or UO_4476 (O_4476,N_49560,N_49529);
nor UO_4477 (O_4477,N_49881,N_49513);
nand UO_4478 (O_4478,N_49581,N_49903);
xnor UO_4479 (O_4479,N_49516,N_49987);
nor UO_4480 (O_4480,N_49815,N_49603);
or UO_4481 (O_4481,N_49996,N_49980);
nor UO_4482 (O_4482,N_49927,N_49709);
xnor UO_4483 (O_4483,N_49621,N_49577);
or UO_4484 (O_4484,N_49629,N_49907);
or UO_4485 (O_4485,N_49682,N_49664);
and UO_4486 (O_4486,N_49504,N_49931);
nand UO_4487 (O_4487,N_49569,N_49623);
xor UO_4488 (O_4488,N_49912,N_49772);
nand UO_4489 (O_4489,N_49913,N_49693);
or UO_4490 (O_4490,N_49903,N_49925);
nand UO_4491 (O_4491,N_49527,N_49818);
nor UO_4492 (O_4492,N_49759,N_49850);
and UO_4493 (O_4493,N_49801,N_49862);
nor UO_4494 (O_4494,N_49781,N_49750);
or UO_4495 (O_4495,N_49863,N_49691);
or UO_4496 (O_4496,N_49653,N_49829);
xnor UO_4497 (O_4497,N_49932,N_49917);
or UO_4498 (O_4498,N_49502,N_49877);
nand UO_4499 (O_4499,N_49901,N_49840);
and UO_4500 (O_4500,N_49892,N_49514);
and UO_4501 (O_4501,N_49858,N_49586);
or UO_4502 (O_4502,N_49936,N_49923);
nor UO_4503 (O_4503,N_49670,N_49797);
nor UO_4504 (O_4504,N_49954,N_49920);
or UO_4505 (O_4505,N_49961,N_49802);
nor UO_4506 (O_4506,N_49949,N_49519);
xor UO_4507 (O_4507,N_49978,N_49789);
or UO_4508 (O_4508,N_49685,N_49625);
xor UO_4509 (O_4509,N_49846,N_49682);
xnor UO_4510 (O_4510,N_49505,N_49624);
nor UO_4511 (O_4511,N_49809,N_49947);
nor UO_4512 (O_4512,N_49855,N_49625);
and UO_4513 (O_4513,N_49696,N_49527);
and UO_4514 (O_4514,N_49695,N_49686);
nor UO_4515 (O_4515,N_49983,N_49568);
or UO_4516 (O_4516,N_49853,N_49790);
or UO_4517 (O_4517,N_49793,N_49945);
nand UO_4518 (O_4518,N_49800,N_49644);
and UO_4519 (O_4519,N_49701,N_49877);
xnor UO_4520 (O_4520,N_49962,N_49705);
and UO_4521 (O_4521,N_49613,N_49889);
nor UO_4522 (O_4522,N_49964,N_49990);
nand UO_4523 (O_4523,N_49718,N_49753);
or UO_4524 (O_4524,N_49531,N_49973);
xor UO_4525 (O_4525,N_49918,N_49826);
and UO_4526 (O_4526,N_49552,N_49899);
nand UO_4527 (O_4527,N_49522,N_49676);
xnor UO_4528 (O_4528,N_49859,N_49942);
nor UO_4529 (O_4529,N_49668,N_49938);
nand UO_4530 (O_4530,N_49554,N_49571);
or UO_4531 (O_4531,N_49798,N_49925);
or UO_4532 (O_4532,N_49899,N_49717);
nor UO_4533 (O_4533,N_49554,N_49523);
xor UO_4534 (O_4534,N_49988,N_49580);
nor UO_4535 (O_4535,N_49530,N_49895);
and UO_4536 (O_4536,N_49654,N_49907);
xor UO_4537 (O_4537,N_49805,N_49995);
and UO_4538 (O_4538,N_49685,N_49949);
or UO_4539 (O_4539,N_49977,N_49616);
or UO_4540 (O_4540,N_49625,N_49817);
or UO_4541 (O_4541,N_49893,N_49687);
nor UO_4542 (O_4542,N_49933,N_49861);
and UO_4543 (O_4543,N_49960,N_49616);
or UO_4544 (O_4544,N_49951,N_49768);
nand UO_4545 (O_4545,N_49716,N_49507);
xor UO_4546 (O_4546,N_49550,N_49677);
xnor UO_4547 (O_4547,N_49629,N_49985);
xor UO_4548 (O_4548,N_49640,N_49951);
nor UO_4549 (O_4549,N_49979,N_49951);
xnor UO_4550 (O_4550,N_49854,N_49926);
xor UO_4551 (O_4551,N_49825,N_49663);
xor UO_4552 (O_4552,N_49798,N_49559);
or UO_4553 (O_4553,N_49634,N_49897);
nor UO_4554 (O_4554,N_49877,N_49814);
nand UO_4555 (O_4555,N_49618,N_49544);
nor UO_4556 (O_4556,N_49952,N_49681);
nand UO_4557 (O_4557,N_49563,N_49562);
nand UO_4558 (O_4558,N_49550,N_49578);
nor UO_4559 (O_4559,N_49664,N_49680);
xnor UO_4560 (O_4560,N_49553,N_49846);
nor UO_4561 (O_4561,N_49858,N_49758);
or UO_4562 (O_4562,N_49543,N_49620);
xnor UO_4563 (O_4563,N_49628,N_49863);
and UO_4564 (O_4564,N_49607,N_49903);
or UO_4565 (O_4565,N_49795,N_49959);
xnor UO_4566 (O_4566,N_49850,N_49933);
nor UO_4567 (O_4567,N_49866,N_49979);
and UO_4568 (O_4568,N_49786,N_49615);
or UO_4569 (O_4569,N_49668,N_49548);
or UO_4570 (O_4570,N_49587,N_49725);
xor UO_4571 (O_4571,N_49810,N_49999);
nand UO_4572 (O_4572,N_49641,N_49683);
or UO_4573 (O_4573,N_49804,N_49878);
nand UO_4574 (O_4574,N_49993,N_49544);
or UO_4575 (O_4575,N_49629,N_49705);
or UO_4576 (O_4576,N_49622,N_49788);
nor UO_4577 (O_4577,N_49736,N_49543);
nor UO_4578 (O_4578,N_49745,N_49936);
or UO_4579 (O_4579,N_49604,N_49722);
or UO_4580 (O_4580,N_49923,N_49675);
or UO_4581 (O_4581,N_49666,N_49599);
or UO_4582 (O_4582,N_49625,N_49521);
or UO_4583 (O_4583,N_49718,N_49671);
and UO_4584 (O_4584,N_49660,N_49696);
nand UO_4585 (O_4585,N_49862,N_49752);
and UO_4586 (O_4586,N_49577,N_49873);
nor UO_4587 (O_4587,N_49557,N_49642);
and UO_4588 (O_4588,N_49716,N_49864);
xnor UO_4589 (O_4589,N_49707,N_49875);
or UO_4590 (O_4590,N_49545,N_49610);
and UO_4591 (O_4591,N_49790,N_49905);
xnor UO_4592 (O_4592,N_49913,N_49962);
nand UO_4593 (O_4593,N_49915,N_49850);
and UO_4594 (O_4594,N_49698,N_49895);
nor UO_4595 (O_4595,N_49951,N_49869);
xor UO_4596 (O_4596,N_49549,N_49884);
or UO_4597 (O_4597,N_49720,N_49510);
and UO_4598 (O_4598,N_49898,N_49952);
nor UO_4599 (O_4599,N_49595,N_49696);
and UO_4600 (O_4600,N_49797,N_49547);
and UO_4601 (O_4601,N_49808,N_49617);
nand UO_4602 (O_4602,N_49600,N_49799);
nor UO_4603 (O_4603,N_49996,N_49697);
and UO_4604 (O_4604,N_49825,N_49511);
nor UO_4605 (O_4605,N_49659,N_49824);
nor UO_4606 (O_4606,N_49716,N_49579);
nor UO_4607 (O_4607,N_49951,N_49538);
or UO_4608 (O_4608,N_49880,N_49645);
and UO_4609 (O_4609,N_49884,N_49911);
and UO_4610 (O_4610,N_49690,N_49777);
nor UO_4611 (O_4611,N_49772,N_49525);
and UO_4612 (O_4612,N_49549,N_49851);
or UO_4613 (O_4613,N_49891,N_49813);
and UO_4614 (O_4614,N_49812,N_49836);
nand UO_4615 (O_4615,N_49896,N_49938);
nand UO_4616 (O_4616,N_49871,N_49907);
and UO_4617 (O_4617,N_49615,N_49564);
nor UO_4618 (O_4618,N_49785,N_49744);
or UO_4619 (O_4619,N_49546,N_49892);
nor UO_4620 (O_4620,N_49844,N_49516);
xnor UO_4621 (O_4621,N_49637,N_49741);
and UO_4622 (O_4622,N_49788,N_49559);
nand UO_4623 (O_4623,N_49682,N_49941);
or UO_4624 (O_4624,N_49831,N_49711);
nor UO_4625 (O_4625,N_49601,N_49857);
xnor UO_4626 (O_4626,N_49897,N_49556);
nand UO_4627 (O_4627,N_49549,N_49820);
nor UO_4628 (O_4628,N_49752,N_49758);
or UO_4629 (O_4629,N_49664,N_49870);
nor UO_4630 (O_4630,N_49950,N_49881);
xor UO_4631 (O_4631,N_49959,N_49802);
or UO_4632 (O_4632,N_49970,N_49951);
nand UO_4633 (O_4633,N_49766,N_49604);
nor UO_4634 (O_4634,N_49815,N_49555);
or UO_4635 (O_4635,N_49909,N_49978);
nor UO_4636 (O_4636,N_49722,N_49921);
and UO_4637 (O_4637,N_49869,N_49955);
xnor UO_4638 (O_4638,N_49859,N_49591);
nand UO_4639 (O_4639,N_49762,N_49642);
and UO_4640 (O_4640,N_49851,N_49860);
nand UO_4641 (O_4641,N_49958,N_49502);
xor UO_4642 (O_4642,N_49611,N_49503);
and UO_4643 (O_4643,N_49884,N_49864);
xnor UO_4644 (O_4644,N_49956,N_49990);
nor UO_4645 (O_4645,N_49532,N_49699);
or UO_4646 (O_4646,N_49895,N_49710);
xor UO_4647 (O_4647,N_49884,N_49988);
or UO_4648 (O_4648,N_49891,N_49881);
and UO_4649 (O_4649,N_49569,N_49873);
and UO_4650 (O_4650,N_49542,N_49739);
xnor UO_4651 (O_4651,N_49910,N_49686);
and UO_4652 (O_4652,N_49990,N_49724);
xor UO_4653 (O_4653,N_49783,N_49753);
xnor UO_4654 (O_4654,N_49764,N_49850);
and UO_4655 (O_4655,N_49660,N_49645);
nand UO_4656 (O_4656,N_49659,N_49627);
or UO_4657 (O_4657,N_49806,N_49900);
xor UO_4658 (O_4658,N_49859,N_49541);
nand UO_4659 (O_4659,N_49971,N_49595);
or UO_4660 (O_4660,N_49816,N_49750);
nand UO_4661 (O_4661,N_49882,N_49729);
nor UO_4662 (O_4662,N_49837,N_49666);
nor UO_4663 (O_4663,N_49659,N_49530);
xnor UO_4664 (O_4664,N_49673,N_49802);
and UO_4665 (O_4665,N_49505,N_49635);
or UO_4666 (O_4666,N_49566,N_49774);
or UO_4667 (O_4667,N_49904,N_49601);
or UO_4668 (O_4668,N_49511,N_49509);
nand UO_4669 (O_4669,N_49900,N_49694);
or UO_4670 (O_4670,N_49813,N_49504);
nand UO_4671 (O_4671,N_49744,N_49758);
and UO_4672 (O_4672,N_49732,N_49806);
xnor UO_4673 (O_4673,N_49802,N_49871);
and UO_4674 (O_4674,N_49657,N_49908);
nor UO_4675 (O_4675,N_49776,N_49851);
and UO_4676 (O_4676,N_49505,N_49886);
and UO_4677 (O_4677,N_49622,N_49984);
and UO_4678 (O_4678,N_49924,N_49681);
and UO_4679 (O_4679,N_49625,N_49692);
nor UO_4680 (O_4680,N_49688,N_49916);
and UO_4681 (O_4681,N_49929,N_49730);
nor UO_4682 (O_4682,N_49674,N_49796);
and UO_4683 (O_4683,N_49975,N_49793);
and UO_4684 (O_4684,N_49669,N_49601);
nand UO_4685 (O_4685,N_49884,N_49996);
nand UO_4686 (O_4686,N_49595,N_49691);
or UO_4687 (O_4687,N_49566,N_49700);
nand UO_4688 (O_4688,N_49818,N_49668);
nor UO_4689 (O_4689,N_49725,N_49859);
xor UO_4690 (O_4690,N_49795,N_49819);
and UO_4691 (O_4691,N_49847,N_49646);
nor UO_4692 (O_4692,N_49739,N_49760);
xor UO_4693 (O_4693,N_49983,N_49628);
xnor UO_4694 (O_4694,N_49947,N_49650);
nor UO_4695 (O_4695,N_49701,N_49843);
or UO_4696 (O_4696,N_49659,N_49667);
nor UO_4697 (O_4697,N_49802,N_49637);
nand UO_4698 (O_4698,N_49928,N_49669);
nor UO_4699 (O_4699,N_49725,N_49742);
nand UO_4700 (O_4700,N_49982,N_49718);
or UO_4701 (O_4701,N_49892,N_49805);
nand UO_4702 (O_4702,N_49506,N_49672);
or UO_4703 (O_4703,N_49755,N_49810);
nand UO_4704 (O_4704,N_49697,N_49604);
nand UO_4705 (O_4705,N_49512,N_49887);
or UO_4706 (O_4706,N_49804,N_49537);
and UO_4707 (O_4707,N_49528,N_49618);
nor UO_4708 (O_4708,N_49971,N_49644);
nand UO_4709 (O_4709,N_49967,N_49968);
nor UO_4710 (O_4710,N_49622,N_49611);
or UO_4711 (O_4711,N_49636,N_49567);
nand UO_4712 (O_4712,N_49700,N_49646);
xnor UO_4713 (O_4713,N_49835,N_49703);
xor UO_4714 (O_4714,N_49855,N_49974);
nor UO_4715 (O_4715,N_49991,N_49728);
and UO_4716 (O_4716,N_49582,N_49948);
or UO_4717 (O_4717,N_49935,N_49981);
nand UO_4718 (O_4718,N_49704,N_49904);
or UO_4719 (O_4719,N_49983,N_49747);
nor UO_4720 (O_4720,N_49975,N_49993);
and UO_4721 (O_4721,N_49753,N_49847);
xnor UO_4722 (O_4722,N_49609,N_49848);
and UO_4723 (O_4723,N_49943,N_49876);
or UO_4724 (O_4724,N_49791,N_49687);
nand UO_4725 (O_4725,N_49713,N_49500);
nand UO_4726 (O_4726,N_49608,N_49871);
nor UO_4727 (O_4727,N_49976,N_49584);
nor UO_4728 (O_4728,N_49834,N_49905);
and UO_4729 (O_4729,N_49898,N_49789);
nor UO_4730 (O_4730,N_49602,N_49894);
or UO_4731 (O_4731,N_49959,N_49617);
nand UO_4732 (O_4732,N_49734,N_49557);
nor UO_4733 (O_4733,N_49573,N_49921);
nand UO_4734 (O_4734,N_49843,N_49807);
or UO_4735 (O_4735,N_49863,N_49823);
and UO_4736 (O_4736,N_49737,N_49538);
xnor UO_4737 (O_4737,N_49738,N_49952);
xnor UO_4738 (O_4738,N_49648,N_49645);
and UO_4739 (O_4739,N_49861,N_49777);
nand UO_4740 (O_4740,N_49970,N_49886);
xnor UO_4741 (O_4741,N_49972,N_49727);
and UO_4742 (O_4742,N_49527,N_49630);
nor UO_4743 (O_4743,N_49670,N_49678);
and UO_4744 (O_4744,N_49803,N_49967);
xor UO_4745 (O_4745,N_49639,N_49552);
nor UO_4746 (O_4746,N_49795,N_49642);
or UO_4747 (O_4747,N_49898,N_49913);
nand UO_4748 (O_4748,N_49644,N_49533);
nor UO_4749 (O_4749,N_49721,N_49508);
or UO_4750 (O_4750,N_49561,N_49547);
or UO_4751 (O_4751,N_49528,N_49813);
xor UO_4752 (O_4752,N_49914,N_49947);
nor UO_4753 (O_4753,N_49951,N_49781);
and UO_4754 (O_4754,N_49830,N_49947);
and UO_4755 (O_4755,N_49906,N_49828);
nand UO_4756 (O_4756,N_49528,N_49929);
or UO_4757 (O_4757,N_49543,N_49828);
or UO_4758 (O_4758,N_49856,N_49570);
nor UO_4759 (O_4759,N_49972,N_49629);
and UO_4760 (O_4760,N_49926,N_49596);
nor UO_4761 (O_4761,N_49847,N_49767);
xnor UO_4762 (O_4762,N_49623,N_49949);
or UO_4763 (O_4763,N_49583,N_49673);
nor UO_4764 (O_4764,N_49595,N_49586);
nand UO_4765 (O_4765,N_49757,N_49954);
nand UO_4766 (O_4766,N_49915,N_49821);
xor UO_4767 (O_4767,N_49760,N_49719);
xor UO_4768 (O_4768,N_49698,N_49907);
nand UO_4769 (O_4769,N_49889,N_49614);
and UO_4770 (O_4770,N_49993,N_49947);
xnor UO_4771 (O_4771,N_49576,N_49822);
or UO_4772 (O_4772,N_49545,N_49665);
and UO_4773 (O_4773,N_49973,N_49537);
nor UO_4774 (O_4774,N_49982,N_49680);
and UO_4775 (O_4775,N_49622,N_49814);
or UO_4776 (O_4776,N_49522,N_49506);
xnor UO_4777 (O_4777,N_49591,N_49820);
xor UO_4778 (O_4778,N_49677,N_49737);
and UO_4779 (O_4779,N_49813,N_49584);
and UO_4780 (O_4780,N_49640,N_49577);
and UO_4781 (O_4781,N_49933,N_49506);
xnor UO_4782 (O_4782,N_49858,N_49734);
xor UO_4783 (O_4783,N_49786,N_49563);
or UO_4784 (O_4784,N_49547,N_49892);
or UO_4785 (O_4785,N_49692,N_49659);
or UO_4786 (O_4786,N_49573,N_49902);
nor UO_4787 (O_4787,N_49530,N_49905);
and UO_4788 (O_4788,N_49590,N_49829);
or UO_4789 (O_4789,N_49612,N_49509);
nor UO_4790 (O_4790,N_49543,N_49794);
xor UO_4791 (O_4791,N_49921,N_49695);
nand UO_4792 (O_4792,N_49914,N_49617);
nor UO_4793 (O_4793,N_49561,N_49832);
xor UO_4794 (O_4794,N_49737,N_49675);
nor UO_4795 (O_4795,N_49849,N_49902);
nand UO_4796 (O_4796,N_49709,N_49983);
nor UO_4797 (O_4797,N_49626,N_49799);
and UO_4798 (O_4798,N_49840,N_49553);
xor UO_4799 (O_4799,N_49503,N_49925);
nor UO_4800 (O_4800,N_49644,N_49905);
nand UO_4801 (O_4801,N_49805,N_49676);
xor UO_4802 (O_4802,N_49558,N_49971);
or UO_4803 (O_4803,N_49997,N_49892);
nor UO_4804 (O_4804,N_49583,N_49659);
xnor UO_4805 (O_4805,N_49732,N_49710);
nor UO_4806 (O_4806,N_49884,N_49672);
or UO_4807 (O_4807,N_49667,N_49984);
or UO_4808 (O_4808,N_49740,N_49784);
or UO_4809 (O_4809,N_49787,N_49997);
or UO_4810 (O_4810,N_49509,N_49680);
nor UO_4811 (O_4811,N_49778,N_49629);
nor UO_4812 (O_4812,N_49512,N_49881);
nor UO_4813 (O_4813,N_49889,N_49510);
and UO_4814 (O_4814,N_49663,N_49952);
and UO_4815 (O_4815,N_49979,N_49590);
nand UO_4816 (O_4816,N_49640,N_49969);
nor UO_4817 (O_4817,N_49596,N_49629);
or UO_4818 (O_4818,N_49690,N_49877);
xnor UO_4819 (O_4819,N_49550,N_49939);
xnor UO_4820 (O_4820,N_49863,N_49600);
nand UO_4821 (O_4821,N_49993,N_49891);
nand UO_4822 (O_4822,N_49933,N_49528);
xnor UO_4823 (O_4823,N_49789,N_49691);
and UO_4824 (O_4824,N_49711,N_49857);
nor UO_4825 (O_4825,N_49902,N_49623);
xor UO_4826 (O_4826,N_49847,N_49732);
or UO_4827 (O_4827,N_49836,N_49619);
or UO_4828 (O_4828,N_49637,N_49814);
nand UO_4829 (O_4829,N_49668,N_49557);
nand UO_4830 (O_4830,N_49890,N_49783);
xor UO_4831 (O_4831,N_49573,N_49825);
nand UO_4832 (O_4832,N_49506,N_49751);
nor UO_4833 (O_4833,N_49714,N_49867);
and UO_4834 (O_4834,N_49792,N_49906);
nor UO_4835 (O_4835,N_49812,N_49696);
and UO_4836 (O_4836,N_49761,N_49740);
nor UO_4837 (O_4837,N_49691,N_49724);
nor UO_4838 (O_4838,N_49767,N_49545);
or UO_4839 (O_4839,N_49856,N_49765);
nor UO_4840 (O_4840,N_49538,N_49728);
nand UO_4841 (O_4841,N_49549,N_49988);
or UO_4842 (O_4842,N_49682,N_49931);
nor UO_4843 (O_4843,N_49685,N_49579);
and UO_4844 (O_4844,N_49936,N_49646);
xnor UO_4845 (O_4845,N_49520,N_49901);
xor UO_4846 (O_4846,N_49713,N_49899);
or UO_4847 (O_4847,N_49533,N_49904);
xor UO_4848 (O_4848,N_49981,N_49801);
nor UO_4849 (O_4849,N_49750,N_49934);
nand UO_4850 (O_4850,N_49864,N_49793);
and UO_4851 (O_4851,N_49975,N_49998);
and UO_4852 (O_4852,N_49691,N_49569);
nand UO_4853 (O_4853,N_49551,N_49563);
nor UO_4854 (O_4854,N_49807,N_49662);
or UO_4855 (O_4855,N_49528,N_49517);
xnor UO_4856 (O_4856,N_49766,N_49667);
nor UO_4857 (O_4857,N_49650,N_49986);
and UO_4858 (O_4858,N_49534,N_49924);
nor UO_4859 (O_4859,N_49753,N_49502);
or UO_4860 (O_4860,N_49622,N_49965);
nand UO_4861 (O_4861,N_49939,N_49697);
or UO_4862 (O_4862,N_49777,N_49809);
nor UO_4863 (O_4863,N_49527,N_49582);
xnor UO_4864 (O_4864,N_49705,N_49839);
xnor UO_4865 (O_4865,N_49734,N_49703);
xor UO_4866 (O_4866,N_49761,N_49641);
or UO_4867 (O_4867,N_49629,N_49877);
and UO_4868 (O_4868,N_49929,N_49549);
or UO_4869 (O_4869,N_49883,N_49856);
nand UO_4870 (O_4870,N_49765,N_49700);
and UO_4871 (O_4871,N_49831,N_49953);
nand UO_4872 (O_4872,N_49746,N_49887);
nor UO_4873 (O_4873,N_49665,N_49700);
nand UO_4874 (O_4874,N_49636,N_49960);
nand UO_4875 (O_4875,N_49568,N_49739);
xnor UO_4876 (O_4876,N_49707,N_49642);
nand UO_4877 (O_4877,N_49944,N_49950);
xnor UO_4878 (O_4878,N_49635,N_49745);
and UO_4879 (O_4879,N_49855,N_49925);
nor UO_4880 (O_4880,N_49863,N_49534);
nor UO_4881 (O_4881,N_49535,N_49971);
or UO_4882 (O_4882,N_49748,N_49796);
nor UO_4883 (O_4883,N_49690,N_49749);
xnor UO_4884 (O_4884,N_49732,N_49621);
or UO_4885 (O_4885,N_49719,N_49639);
and UO_4886 (O_4886,N_49570,N_49615);
nand UO_4887 (O_4887,N_49662,N_49602);
and UO_4888 (O_4888,N_49731,N_49732);
nor UO_4889 (O_4889,N_49567,N_49906);
and UO_4890 (O_4890,N_49654,N_49545);
and UO_4891 (O_4891,N_49898,N_49558);
or UO_4892 (O_4892,N_49637,N_49935);
nor UO_4893 (O_4893,N_49831,N_49781);
nand UO_4894 (O_4894,N_49598,N_49979);
nand UO_4895 (O_4895,N_49824,N_49878);
and UO_4896 (O_4896,N_49700,N_49966);
nand UO_4897 (O_4897,N_49644,N_49754);
and UO_4898 (O_4898,N_49561,N_49897);
nand UO_4899 (O_4899,N_49594,N_49789);
or UO_4900 (O_4900,N_49642,N_49508);
nand UO_4901 (O_4901,N_49876,N_49593);
nand UO_4902 (O_4902,N_49777,N_49693);
nand UO_4903 (O_4903,N_49648,N_49574);
nor UO_4904 (O_4904,N_49630,N_49858);
and UO_4905 (O_4905,N_49766,N_49951);
nand UO_4906 (O_4906,N_49692,N_49957);
xor UO_4907 (O_4907,N_49691,N_49679);
and UO_4908 (O_4908,N_49601,N_49642);
and UO_4909 (O_4909,N_49594,N_49568);
and UO_4910 (O_4910,N_49951,N_49577);
nor UO_4911 (O_4911,N_49708,N_49732);
nand UO_4912 (O_4912,N_49588,N_49931);
or UO_4913 (O_4913,N_49827,N_49707);
or UO_4914 (O_4914,N_49725,N_49622);
nand UO_4915 (O_4915,N_49529,N_49827);
xnor UO_4916 (O_4916,N_49596,N_49796);
or UO_4917 (O_4917,N_49633,N_49654);
nand UO_4918 (O_4918,N_49886,N_49907);
xnor UO_4919 (O_4919,N_49856,N_49516);
or UO_4920 (O_4920,N_49700,N_49921);
or UO_4921 (O_4921,N_49869,N_49551);
xnor UO_4922 (O_4922,N_49501,N_49738);
nor UO_4923 (O_4923,N_49919,N_49624);
and UO_4924 (O_4924,N_49548,N_49546);
nand UO_4925 (O_4925,N_49769,N_49950);
or UO_4926 (O_4926,N_49709,N_49755);
or UO_4927 (O_4927,N_49834,N_49682);
xor UO_4928 (O_4928,N_49916,N_49700);
xor UO_4929 (O_4929,N_49992,N_49805);
and UO_4930 (O_4930,N_49617,N_49934);
and UO_4931 (O_4931,N_49902,N_49836);
nor UO_4932 (O_4932,N_49858,N_49764);
nor UO_4933 (O_4933,N_49951,N_49785);
or UO_4934 (O_4934,N_49856,N_49574);
and UO_4935 (O_4935,N_49986,N_49939);
nor UO_4936 (O_4936,N_49728,N_49952);
and UO_4937 (O_4937,N_49941,N_49854);
nand UO_4938 (O_4938,N_49761,N_49879);
nor UO_4939 (O_4939,N_49509,N_49952);
nor UO_4940 (O_4940,N_49770,N_49776);
or UO_4941 (O_4941,N_49669,N_49518);
nor UO_4942 (O_4942,N_49934,N_49955);
or UO_4943 (O_4943,N_49575,N_49517);
nand UO_4944 (O_4944,N_49905,N_49953);
nand UO_4945 (O_4945,N_49656,N_49942);
xor UO_4946 (O_4946,N_49880,N_49591);
nand UO_4947 (O_4947,N_49614,N_49677);
and UO_4948 (O_4948,N_49884,N_49791);
or UO_4949 (O_4949,N_49807,N_49506);
or UO_4950 (O_4950,N_49674,N_49794);
xor UO_4951 (O_4951,N_49632,N_49638);
and UO_4952 (O_4952,N_49586,N_49935);
nand UO_4953 (O_4953,N_49864,N_49756);
nor UO_4954 (O_4954,N_49740,N_49565);
nor UO_4955 (O_4955,N_49969,N_49840);
or UO_4956 (O_4956,N_49891,N_49781);
xor UO_4957 (O_4957,N_49894,N_49977);
nor UO_4958 (O_4958,N_49880,N_49862);
and UO_4959 (O_4959,N_49879,N_49649);
and UO_4960 (O_4960,N_49629,N_49897);
or UO_4961 (O_4961,N_49660,N_49693);
xnor UO_4962 (O_4962,N_49776,N_49725);
nor UO_4963 (O_4963,N_49539,N_49615);
or UO_4964 (O_4964,N_49735,N_49970);
and UO_4965 (O_4965,N_49710,N_49670);
nand UO_4966 (O_4966,N_49927,N_49920);
nor UO_4967 (O_4967,N_49648,N_49991);
or UO_4968 (O_4968,N_49572,N_49965);
xor UO_4969 (O_4969,N_49842,N_49943);
nand UO_4970 (O_4970,N_49569,N_49660);
xor UO_4971 (O_4971,N_49799,N_49980);
and UO_4972 (O_4972,N_49950,N_49541);
xnor UO_4973 (O_4973,N_49911,N_49779);
xor UO_4974 (O_4974,N_49791,N_49844);
nor UO_4975 (O_4975,N_49612,N_49894);
and UO_4976 (O_4976,N_49933,N_49765);
or UO_4977 (O_4977,N_49654,N_49601);
and UO_4978 (O_4978,N_49645,N_49612);
nor UO_4979 (O_4979,N_49515,N_49797);
nor UO_4980 (O_4980,N_49549,N_49625);
xor UO_4981 (O_4981,N_49870,N_49536);
xor UO_4982 (O_4982,N_49941,N_49607);
xor UO_4983 (O_4983,N_49754,N_49552);
or UO_4984 (O_4984,N_49655,N_49508);
nor UO_4985 (O_4985,N_49927,N_49822);
and UO_4986 (O_4986,N_49777,N_49978);
nor UO_4987 (O_4987,N_49738,N_49881);
nand UO_4988 (O_4988,N_49517,N_49747);
or UO_4989 (O_4989,N_49718,N_49765);
xnor UO_4990 (O_4990,N_49976,N_49744);
nand UO_4991 (O_4991,N_49583,N_49893);
or UO_4992 (O_4992,N_49610,N_49603);
and UO_4993 (O_4993,N_49946,N_49908);
or UO_4994 (O_4994,N_49825,N_49540);
nor UO_4995 (O_4995,N_49923,N_49526);
and UO_4996 (O_4996,N_49575,N_49965);
nand UO_4997 (O_4997,N_49900,N_49521);
nor UO_4998 (O_4998,N_49930,N_49701);
xnor UO_4999 (O_4999,N_49771,N_49627);
endmodule