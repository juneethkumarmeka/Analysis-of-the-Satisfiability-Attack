module basic_750_5000_1000_25_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_669,In_146);
nor U1 (N_1,In_735,In_41);
and U2 (N_2,In_581,In_496);
and U3 (N_3,In_598,In_387);
nand U4 (N_4,In_237,In_568);
nand U5 (N_5,In_455,In_9);
nand U6 (N_6,In_471,In_155);
and U7 (N_7,In_474,In_55);
nand U8 (N_8,In_677,In_484);
and U9 (N_9,In_222,In_532);
or U10 (N_10,In_621,In_319);
or U11 (N_11,In_630,In_352);
nor U12 (N_12,In_705,In_176);
or U13 (N_13,In_724,In_589);
nor U14 (N_14,In_715,In_304);
or U15 (N_15,In_683,In_593);
or U16 (N_16,In_173,In_157);
nor U17 (N_17,In_510,In_274);
or U18 (N_18,In_542,In_296);
nor U19 (N_19,In_311,In_341);
nor U20 (N_20,In_569,In_162);
nand U21 (N_21,In_125,In_14);
and U22 (N_22,In_689,In_137);
and U23 (N_23,In_343,In_385);
or U24 (N_24,In_430,In_670);
and U25 (N_25,In_269,In_134);
nand U26 (N_26,In_242,In_288);
nand U27 (N_27,In_442,In_577);
and U28 (N_28,In_410,In_25);
and U29 (N_29,In_239,In_720);
nand U30 (N_30,In_567,In_22);
nand U31 (N_31,In_616,In_167);
nand U32 (N_32,In_540,In_73);
or U33 (N_33,In_62,In_472);
and U34 (N_34,In_365,In_263);
nor U35 (N_35,In_641,In_245);
xnor U36 (N_36,In_128,In_210);
and U37 (N_37,In_556,In_537);
or U38 (N_38,In_721,In_583);
or U39 (N_39,In_250,In_283);
nand U40 (N_40,In_278,In_638);
or U41 (N_41,In_457,In_742);
or U42 (N_42,In_699,In_597);
nor U43 (N_43,In_129,In_694);
or U44 (N_44,In_637,In_511);
or U45 (N_45,In_646,In_733);
nor U46 (N_46,In_106,In_254);
nor U47 (N_47,In_315,In_46);
nor U48 (N_48,In_60,In_632);
nand U49 (N_49,In_656,In_30);
or U50 (N_50,In_132,In_276);
nor U51 (N_51,In_557,In_223);
and U52 (N_52,In_179,In_199);
and U53 (N_53,In_184,In_388);
or U54 (N_54,In_18,In_163);
xor U55 (N_55,In_518,In_224);
xnor U56 (N_56,In_688,In_204);
nand U57 (N_57,In_555,In_338);
nand U58 (N_58,In_533,In_57);
nor U59 (N_59,In_166,In_213);
nand U60 (N_60,In_560,In_684);
or U61 (N_61,In_333,In_428);
nand U62 (N_62,In_285,In_101);
nor U63 (N_63,In_329,In_396);
nand U64 (N_64,In_248,In_152);
nor U65 (N_65,In_290,In_494);
nor U66 (N_66,In_83,In_122);
nand U67 (N_67,In_215,In_5);
nor U68 (N_68,In_603,In_746);
nor U69 (N_69,In_371,In_447);
nor U70 (N_70,In_96,In_233);
nand U71 (N_71,In_139,In_2);
and U72 (N_72,In_231,In_727);
nand U73 (N_73,In_702,In_421);
nand U74 (N_74,In_287,In_153);
nand U75 (N_75,In_367,In_389);
nand U76 (N_76,In_413,In_726);
xnor U77 (N_77,In_397,In_402);
and U78 (N_78,In_160,In_99);
nand U79 (N_79,In_664,In_107);
or U80 (N_80,In_284,In_429);
or U81 (N_81,In_585,In_189);
or U82 (N_82,In_703,In_711);
or U83 (N_83,In_528,In_265);
nor U84 (N_84,In_325,In_196);
nand U85 (N_85,In_138,In_177);
nor U86 (N_86,In_16,In_690);
or U87 (N_87,In_282,In_501);
nor U88 (N_88,In_629,In_561);
or U89 (N_89,In_255,In_226);
nand U90 (N_90,In_574,In_227);
nand U91 (N_91,In_360,In_252);
nand U92 (N_92,In_20,In_431);
nor U93 (N_93,In_149,In_294);
and U94 (N_94,In_678,In_627);
or U95 (N_95,In_394,In_314);
or U96 (N_96,In_297,In_562);
xnor U97 (N_97,In_114,In_165);
nor U98 (N_98,In_258,In_181);
nand U99 (N_99,In_513,In_682);
and U100 (N_100,In_544,In_526);
and U101 (N_101,In_168,In_564);
or U102 (N_102,In_667,In_347);
and U103 (N_103,In_520,In_257);
and U104 (N_104,In_21,In_29);
and U105 (N_105,In_620,In_71);
and U106 (N_106,In_545,In_225);
nand U107 (N_107,In_470,In_645);
nand U108 (N_108,In_356,In_174);
nor U109 (N_109,In_707,In_626);
nor U110 (N_110,In_498,In_611);
nand U111 (N_111,In_147,In_58);
nor U112 (N_112,In_411,In_485);
and U113 (N_113,In_27,In_156);
and U114 (N_114,In_651,In_212);
nor U115 (N_115,In_441,In_92);
and U116 (N_116,In_148,In_64);
or U117 (N_117,In_698,In_710);
nand U118 (N_118,In_368,In_579);
or U119 (N_119,In_42,In_262);
and U120 (N_120,In_207,In_230);
or U121 (N_121,In_91,In_195);
nor U122 (N_122,In_514,In_384);
nand U123 (N_123,In_330,In_586);
nor U124 (N_124,In_640,In_466);
nor U125 (N_125,In_280,In_743);
nor U126 (N_126,In_539,In_456);
xor U127 (N_127,In_695,In_361);
or U128 (N_128,In_399,In_701);
and U129 (N_129,In_529,In_608);
nand U130 (N_130,In_37,In_191);
and U131 (N_131,In_382,In_551);
and U132 (N_132,In_673,In_435);
or U133 (N_133,In_301,In_159);
or U134 (N_134,In_639,In_89);
or U135 (N_135,In_580,In_261);
and U136 (N_136,In_183,In_595);
nand U137 (N_137,In_334,In_40);
or U138 (N_138,In_374,In_203);
nor U139 (N_139,In_732,In_578);
nand U140 (N_140,In_400,In_44);
or U141 (N_141,In_234,In_744);
or U142 (N_142,In_194,In_610);
and U143 (N_143,In_552,In_509);
nor U144 (N_144,In_105,In_693);
and U145 (N_145,In_481,In_398);
nor U146 (N_146,In_541,In_86);
nand U147 (N_147,In_324,In_522);
and U148 (N_148,In_607,In_469);
nor U149 (N_149,In_584,In_459);
or U150 (N_150,In_450,In_495);
and U151 (N_151,In_416,In_247);
and U152 (N_152,In_476,In_737);
and U153 (N_153,In_74,In_48);
xnor U154 (N_154,In_433,In_8);
and U155 (N_155,In_600,In_475);
or U156 (N_156,In_617,In_624);
nand U157 (N_157,In_351,In_604);
and U158 (N_158,In_504,In_605);
or U159 (N_159,In_205,In_536);
or U160 (N_160,In_477,In_686);
or U161 (N_161,In_363,In_45);
nand U162 (N_162,In_104,In_380);
nor U163 (N_163,In_427,In_650);
or U164 (N_164,In_90,In_658);
and U165 (N_165,In_103,In_590);
nor U166 (N_166,In_164,In_65);
and U167 (N_167,In_13,In_201);
or U168 (N_168,In_599,In_558);
and U169 (N_169,In_588,In_731);
xnor U170 (N_170,In_386,In_685);
nor U171 (N_171,In_644,In_436);
nor U172 (N_172,In_82,In_534);
and U173 (N_173,In_121,In_497);
and U174 (N_174,In_452,In_244);
nor U175 (N_175,In_349,In_381);
or U176 (N_176,In_256,In_525);
nand U177 (N_177,In_661,In_124);
or U178 (N_178,In_232,In_161);
and U179 (N_179,In_725,In_582);
nor U180 (N_180,In_369,In_706);
nand U181 (N_181,In_56,In_171);
nand U182 (N_182,In_749,In_316);
or U183 (N_183,In_505,In_337);
nor U184 (N_184,In_462,In_115);
and U185 (N_185,In_79,In_240);
or U186 (N_186,In_480,In_691);
nand U187 (N_187,In_364,In_328);
or U188 (N_188,In_446,In_359);
or U189 (N_189,In_358,In_424);
and U190 (N_190,In_454,In_591);
or U191 (N_191,In_310,In_523);
nor U192 (N_192,In_508,In_412);
nor U193 (N_193,In_408,In_663);
nor U194 (N_194,In_208,In_741);
nor U195 (N_195,In_649,In_186);
or U196 (N_196,In_521,In_216);
nand U197 (N_197,In_246,In_135);
or U198 (N_198,In_70,In_354);
or U199 (N_199,In_440,In_313);
xor U200 (N_200,N_29,In_559);
and U201 (N_201,In_323,In_643);
and U202 (N_202,In_573,In_415);
and U203 (N_203,N_41,N_48);
nand U204 (N_204,In_299,In_614);
nand U205 (N_205,In_339,In_331);
or U206 (N_206,N_150,In_81);
or U207 (N_207,In_403,In_723);
or U208 (N_208,In_549,N_53);
nand U209 (N_209,In_3,In_622);
nand U210 (N_210,In_185,In_85);
and U211 (N_211,In_492,N_144);
nand U212 (N_212,In_461,In_483);
and U213 (N_213,In_438,N_26);
nor U214 (N_214,In_679,In_652);
nand U215 (N_215,In_628,N_65);
or U216 (N_216,In_251,In_7);
and U217 (N_217,N_170,N_61);
or U218 (N_218,In_243,In_467);
nor U219 (N_219,N_145,In_547);
or U220 (N_220,N_91,N_9);
and U221 (N_221,N_125,In_123);
or U222 (N_222,N_155,N_126);
or U223 (N_223,In_432,N_151);
and U224 (N_224,In_113,N_63);
nor U225 (N_225,In_78,In_515);
nand U226 (N_226,In_175,In_437);
or U227 (N_227,N_105,N_103);
nor U228 (N_228,In_150,In_198);
or U229 (N_229,N_44,In_348);
or U230 (N_230,N_96,In_553);
nand U231 (N_231,In_220,In_214);
nor U232 (N_232,N_135,N_172);
or U233 (N_233,N_165,N_137);
nor U234 (N_234,In_500,N_2);
or U235 (N_235,In_434,N_195);
and U236 (N_236,In_546,In_332);
and U237 (N_237,In_708,N_197);
or U238 (N_238,In_728,In_606);
or U239 (N_239,In_68,In_502);
or U240 (N_240,N_79,In_506);
nor U241 (N_241,N_59,In_302);
nand U242 (N_242,N_85,N_56);
or U243 (N_243,In_266,N_181);
and U244 (N_244,In_671,N_188);
and U245 (N_245,In_322,N_106);
xnor U246 (N_246,In_321,N_175);
nand U247 (N_247,N_143,In_67);
nand U248 (N_248,In_35,N_184);
nand U249 (N_249,In_111,In_229);
and U250 (N_250,In_378,N_78);
or U251 (N_251,In_61,N_141);
nor U252 (N_252,In_426,In_709);
and U253 (N_253,In_393,N_185);
and U254 (N_254,In_53,In_405);
nand U255 (N_255,N_89,In_93);
nand U256 (N_256,N_111,N_30);
nor U257 (N_257,In_344,N_159);
nor U258 (N_258,N_120,N_20);
or U259 (N_259,N_77,In_38);
nor U260 (N_260,N_136,N_133);
or U261 (N_261,In_613,N_43);
and U262 (N_262,In_535,N_14);
and U263 (N_263,In_33,N_37);
nor U264 (N_264,In_102,In_141);
or U265 (N_265,In_31,N_199);
and U266 (N_266,In_370,In_383);
or U267 (N_267,In_260,In_26);
or U268 (N_268,N_113,In_193);
nor U269 (N_269,N_35,In_305);
or U270 (N_270,In_377,N_180);
and U271 (N_271,In_596,In_34);
nor U272 (N_272,In_681,N_109);
or U273 (N_273,In_267,In_503);
and U274 (N_274,In_264,N_154);
xor U275 (N_275,In_404,N_22);
or U276 (N_276,In_17,In_473);
or U277 (N_277,In_373,N_84);
nand U278 (N_278,In_722,In_704);
or U279 (N_279,In_298,N_134);
nor U280 (N_280,In_154,In_345);
nand U281 (N_281,In_118,In_443);
or U282 (N_282,In_392,N_47);
nor U283 (N_283,In_362,N_74);
and U284 (N_284,In_63,In_100);
nand U285 (N_285,In_674,N_87);
or U286 (N_286,In_327,In_675);
nand U287 (N_287,In_6,In_28);
and U288 (N_288,In_517,In_268);
nand U289 (N_289,N_176,In_635);
or U290 (N_290,N_112,In_43);
nand U291 (N_291,N_72,N_82);
nand U292 (N_292,In_131,In_592);
or U293 (N_293,N_116,N_194);
or U294 (N_294,In_145,N_39);
nand U295 (N_295,In_482,N_160);
nor U296 (N_296,In_340,N_54);
and U297 (N_297,In_587,In_407);
nor U298 (N_298,N_107,In_736);
and U299 (N_299,In_714,N_191);
nand U300 (N_300,In_217,In_444);
nand U301 (N_301,N_28,In_700);
and U302 (N_302,N_86,N_45);
xnor U303 (N_303,N_173,N_153);
nand U304 (N_304,In_178,In_94);
nor U305 (N_305,In_636,In_143);
nor U306 (N_306,In_543,N_34);
or U307 (N_307,In_187,In_401);
nand U308 (N_308,In_594,In_716);
and U309 (N_309,N_129,N_90);
nor U310 (N_310,N_23,In_306);
nor U311 (N_311,In_151,N_187);
nand U312 (N_312,In_487,N_66);
and U313 (N_313,In_293,N_193);
nand U314 (N_314,In_133,In_295);
nor U315 (N_315,In_36,In_524);
and U316 (N_316,N_15,In_647);
and U317 (N_317,In_672,In_712);
or U318 (N_318,N_92,N_156);
or U319 (N_319,In_576,In_376);
and U320 (N_320,N_3,N_52);
nand U321 (N_321,In_308,In_218);
nand U322 (N_322,In_309,N_161);
xor U323 (N_323,In_692,In_665);
nand U324 (N_324,In_357,N_139);
and U325 (N_325,In_271,In_75);
nor U326 (N_326,In_516,N_24);
nand U327 (N_327,In_238,In_420);
and U328 (N_328,In_318,In_655);
or U329 (N_329,In_300,In_219);
and U330 (N_330,N_36,In_575);
nand U331 (N_331,N_97,In_291);
nand U332 (N_332,In_448,In_565);
or U333 (N_333,N_83,N_110);
or U334 (N_334,N_179,N_162);
or U335 (N_335,In_303,In_668);
or U336 (N_336,In_372,In_519);
and U337 (N_337,In_192,N_6);
and U338 (N_338,N_131,N_75);
nand U339 (N_339,In_77,N_93);
and U340 (N_340,In_493,N_4);
or U341 (N_341,In_460,In_221);
nor U342 (N_342,In_414,N_12);
nand U343 (N_343,N_182,In_11);
nor U344 (N_344,N_158,In_117);
nor U345 (N_345,In_23,In_379);
nand U346 (N_346,In_142,In_72);
nand U347 (N_347,In_109,N_5);
and U348 (N_348,In_97,N_21);
nor U349 (N_349,In_634,In_696);
and U350 (N_350,In_479,N_152);
and U351 (N_351,N_147,In_188);
or U352 (N_352,N_186,In_307);
or U353 (N_353,In_618,In_734);
and U354 (N_354,N_114,N_101);
nor U355 (N_355,N_115,In_488);
nor U356 (N_356,N_17,In_601);
nand U357 (N_357,In_127,In_119);
and U358 (N_358,N_11,N_128);
and U359 (N_359,In_391,In_451);
nor U360 (N_360,In_24,In_654);
and U361 (N_361,In_418,In_463);
nor U362 (N_362,In_602,In_350);
and U363 (N_363,In_39,In_286);
and U364 (N_364,In_158,In_486);
nor U365 (N_365,In_312,In_648);
nor U366 (N_366,In_116,N_0);
nor U367 (N_367,In_530,In_619);
and U368 (N_368,In_490,In_98);
nand U369 (N_369,N_178,In_631);
nand U370 (N_370,In_687,N_168);
nand U371 (N_371,In_745,In_729);
nor U372 (N_372,In_680,N_98);
and U373 (N_373,In_211,In_609);
and U374 (N_374,N_16,In_642);
nor U375 (N_375,N_88,In_445);
or U376 (N_376,In_612,N_198);
nand U377 (N_377,N_94,In_52);
or U378 (N_378,In_275,N_130);
xnor U379 (N_379,N_190,N_76);
or U380 (N_380,N_149,N_68);
and U381 (N_381,N_146,N_1);
nand U382 (N_382,N_73,N_196);
xor U383 (N_383,In_228,In_144);
nand U384 (N_384,In_170,In_425);
or U385 (N_385,N_148,In_489);
and U386 (N_386,In_563,In_531);
and U387 (N_387,In_80,In_197);
nand U388 (N_388,In_84,N_122);
or U389 (N_389,In_130,In_281);
nand U390 (N_390,N_140,In_465);
nor U391 (N_391,In_657,N_99);
nor U392 (N_392,In_273,In_478);
nor U393 (N_393,In_550,In_253);
nor U394 (N_394,In_355,In_87);
xor U395 (N_395,In_659,In_317);
and U396 (N_396,In_88,N_18);
or U397 (N_397,In_320,N_127);
and U398 (N_398,N_7,In_59);
and U399 (N_399,In_747,In_458);
or U400 (N_400,N_95,N_390);
nand U401 (N_401,N_157,N_50);
xor U402 (N_402,N_358,In_277);
and U403 (N_403,N_142,N_300);
or U404 (N_404,N_366,N_204);
and U405 (N_405,In_548,N_216);
nand U406 (N_406,In_464,N_121);
nor U407 (N_407,N_307,N_362);
and U408 (N_408,N_119,N_236);
or U409 (N_409,N_33,N_203);
and U410 (N_410,In_623,N_229);
or U411 (N_411,In_615,N_340);
or U412 (N_412,N_388,N_250);
and U413 (N_413,N_341,N_269);
nand U414 (N_414,N_367,N_279);
or U415 (N_415,N_342,In_51);
and U416 (N_416,N_355,N_259);
and U417 (N_417,N_292,N_246);
and U418 (N_418,N_397,In_54);
nor U419 (N_419,N_365,N_169);
nand U420 (N_420,N_205,N_255);
or U421 (N_421,N_212,N_57);
nor U422 (N_422,N_396,N_379);
nor U423 (N_423,N_374,N_348);
nand U424 (N_424,In_417,In_66);
or U425 (N_425,In_10,N_380);
xor U426 (N_426,N_305,In_439);
nand U427 (N_427,N_253,N_167);
nor U428 (N_428,N_189,N_351);
nor U429 (N_429,N_226,N_104);
and U430 (N_430,N_240,N_274);
and U431 (N_431,In_172,In_346);
and U432 (N_432,N_306,N_349);
nand U433 (N_433,N_214,N_245);
or U434 (N_434,N_370,N_231);
or U435 (N_435,In_120,N_352);
and U436 (N_436,N_283,N_391);
nand U437 (N_437,N_252,N_293);
and U438 (N_438,In_270,N_49);
nand U439 (N_439,N_206,N_299);
and U440 (N_440,N_361,In_409);
or U441 (N_441,N_377,N_350);
nand U442 (N_442,In_140,N_32);
and U443 (N_443,N_369,N_67);
and U444 (N_444,N_249,In_719);
and U445 (N_445,N_164,N_27);
and U446 (N_446,In_713,In_395);
xnor U447 (N_447,N_46,N_398);
nor U448 (N_448,N_163,N_339);
and U449 (N_449,N_309,N_384);
nand U450 (N_450,N_210,In_390);
nand U451 (N_451,In_717,N_393);
and U452 (N_452,N_69,N_332);
and U453 (N_453,N_273,N_267);
nand U454 (N_454,N_108,In_571);
nand U455 (N_455,In_180,N_275);
nand U456 (N_456,In_47,N_171);
or U457 (N_457,N_266,In_512);
nor U458 (N_458,N_387,N_280);
nor U459 (N_459,N_364,In_108);
or U460 (N_460,N_321,In_730);
nand U461 (N_461,N_62,N_333);
and U462 (N_462,N_177,In_491);
xnor U463 (N_463,N_378,In_236);
nand U464 (N_464,N_227,N_359);
and U465 (N_465,N_234,N_346);
and U466 (N_466,N_219,N_385);
xnor U467 (N_467,In_272,N_308);
or U468 (N_468,N_301,N_200);
and U469 (N_469,N_356,N_276);
nand U470 (N_470,In_200,In_95);
nor U471 (N_471,N_264,N_237);
nand U472 (N_472,In_209,N_381);
or U473 (N_473,N_260,In_190);
and U474 (N_474,N_230,N_265);
nand U475 (N_475,N_208,N_372);
nor U476 (N_476,In_4,N_383);
nor U477 (N_477,N_242,In_666);
and U478 (N_478,N_217,N_256);
nand U479 (N_479,N_58,In_206);
nand U480 (N_480,In_50,N_296);
and U481 (N_481,In_653,N_289);
nor U482 (N_482,N_290,N_330);
or U483 (N_483,N_232,N_64);
or U484 (N_484,In_566,In_570);
nand U485 (N_485,N_284,N_331);
nor U486 (N_486,N_213,N_13);
nor U487 (N_487,N_25,In_366);
nor U488 (N_488,In_342,In_453);
or U489 (N_489,In_69,N_272);
and U490 (N_490,In_748,N_70);
nor U491 (N_491,N_288,In_292);
nand U492 (N_492,N_375,N_183);
nand U493 (N_493,N_353,N_211);
or U494 (N_494,N_257,N_286);
or U495 (N_495,N_258,N_123);
nor U496 (N_496,N_138,N_100);
and U497 (N_497,N_60,In_572);
nor U498 (N_498,N_360,N_357);
or U499 (N_499,In_32,N_271);
nor U500 (N_500,N_323,N_371);
nor U501 (N_501,N_251,N_295);
nor U502 (N_502,N_338,N_343);
nand U503 (N_503,N_285,N_220);
or U504 (N_504,N_319,In_633);
nor U505 (N_505,In_423,N_344);
and U506 (N_506,N_224,N_270);
nor U507 (N_507,N_268,N_354);
or U508 (N_508,N_399,N_336);
or U509 (N_509,N_313,N_337);
and U510 (N_510,N_55,In_676);
and U511 (N_511,In_49,In_110);
and U512 (N_512,In_259,In_739);
and U513 (N_513,N_102,N_202);
and U514 (N_514,In_15,N_124);
and U515 (N_515,N_317,N_373);
and U516 (N_516,N_38,N_225);
and U517 (N_517,N_223,N_81);
and U518 (N_518,N_40,N_118);
and U519 (N_519,N_117,N_310);
or U520 (N_520,N_324,N_315);
nor U521 (N_521,N_261,N_389);
nor U522 (N_522,N_302,N_218);
nor U523 (N_523,In_449,N_392);
nor U524 (N_524,N_262,In_76);
and U525 (N_525,In_112,In_182);
or U526 (N_526,N_241,N_376);
nand U527 (N_527,In_12,N_382);
nand U528 (N_528,In_241,In_335);
nand U529 (N_529,In_740,In_738);
or U530 (N_530,N_297,In_235);
and U531 (N_531,N_239,N_80);
or U532 (N_532,In_136,N_31);
or U533 (N_533,N_287,N_19);
nor U534 (N_534,In_660,In_422);
nor U535 (N_535,N_291,N_335);
or U536 (N_536,N_243,In_326);
and U537 (N_537,N_174,N_327);
or U538 (N_538,N_222,N_166);
nor U539 (N_539,N_395,N_254);
nand U540 (N_540,N_347,N_201);
nand U541 (N_541,N_345,In_507);
nand U542 (N_542,N_10,N_325);
nor U543 (N_543,In_19,In_625);
or U544 (N_544,In_406,N_278);
nand U545 (N_545,N_215,N_326);
and U546 (N_546,N_314,N_394);
or U547 (N_547,In_468,N_328);
and U548 (N_548,N_235,In_169);
and U549 (N_549,N_207,In_126);
nor U550 (N_550,N_363,N_71);
nor U551 (N_551,N_312,In_353);
nand U552 (N_552,N_238,In_289);
nand U553 (N_553,In_499,N_248);
nor U554 (N_554,N_311,In_0);
and U555 (N_555,In_202,In_249);
or U556 (N_556,In_554,N_42);
nor U557 (N_557,In_718,N_294);
or U558 (N_558,N_322,In_527);
nor U559 (N_559,N_303,N_316);
nand U560 (N_560,N_298,N_132);
nand U561 (N_561,N_8,N_277);
or U562 (N_562,N_192,N_320);
or U563 (N_563,N_318,N_329);
nor U564 (N_564,In_538,In_1);
nor U565 (N_565,N_368,N_282);
nand U566 (N_566,N_281,N_386);
nand U567 (N_567,N_209,In_279);
and U568 (N_568,N_263,In_419);
nor U569 (N_569,N_221,In_697);
nor U570 (N_570,N_334,In_375);
or U571 (N_571,In_336,N_233);
nand U572 (N_572,N_228,N_51);
and U573 (N_573,In_662,N_304);
and U574 (N_574,N_244,N_247);
nand U575 (N_575,N_359,In_676);
and U576 (N_576,N_118,N_192);
and U577 (N_577,N_237,N_305);
or U578 (N_578,N_399,N_214);
nor U579 (N_579,N_38,N_377);
nor U580 (N_580,N_358,N_235);
and U581 (N_581,N_286,In_666);
nor U582 (N_582,N_262,N_234);
nand U583 (N_583,N_370,In_548);
and U584 (N_584,In_110,N_349);
or U585 (N_585,In_464,N_189);
and U586 (N_586,In_47,N_100);
nand U587 (N_587,N_370,N_357);
xor U588 (N_588,N_374,In_449);
and U589 (N_589,N_380,N_228);
or U590 (N_590,In_235,N_254);
nor U591 (N_591,N_10,N_257);
and U592 (N_592,N_277,N_203);
or U593 (N_593,N_323,In_570);
and U594 (N_594,N_291,N_342);
and U595 (N_595,In_236,N_49);
nor U596 (N_596,N_367,In_353);
nand U597 (N_597,N_204,N_238);
and U598 (N_598,In_140,N_295);
or U599 (N_599,N_392,N_312);
and U600 (N_600,N_471,N_555);
and U601 (N_601,N_412,N_527);
nor U602 (N_602,N_481,N_566);
nand U603 (N_603,N_576,N_495);
nand U604 (N_604,N_493,N_515);
nor U605 (N_605,N_419,N_429);
and U606 (N_606,N_596,N_568);
nor U607 (N_607,N_451,N_465);
or U608 (N_608,N_500,N_552);
or U609 (N_609,N_525,N_414);
and U610 (N_610,N_469,N_501);
or U611 (N_611,N_562,N_446);
and U612 (N_612,N_406,N_430);
and U613 (N_613,N_557,N_483);
or U614 (N_614,N_559,N_537);
or U615 (N_615,N_427,N_470);
nand U616 (N_616,N_421,N_593);
and U617 (N_617,N_477,N_546);
and U618 (N_618,N_443,N_521);
and U619 (N_619,N_541,N_591);
and U620 (N_620,N_532,N_415);
and U621 (N_621,N_518,N_434);
nand U622 (N_622,N_458,N_487);
nor U623 (N_623,N_435,N_452);
nand U624 (N_624,N_597,N_550);
nand U625 (N_625,N_449,N_486);
nor U626 (N_626,N_503,N_575);
and U627 (N_627,N_491,N_570);
nor U628 (N_628,N_508,N_502);
nor U629 (N_629,N_519,N_578);
nor U630 (N_630,N_485,N_420);
and U631 (N_631,N_499,N_590);
or U632 (N_632,N_404,N_565);
nor U633 (N_633,N_450,N_544);
and U634 (N_634,N_492,N_585);
and U635 (N_635,N_558,N_594);
and U636 (N_636,N_447,N_440);
nor U637 (N_637,N_496,N_428);
xnor U638 (N_638,N_586,N_417);
and U639 (N_639,N_554,N_464);
and U640 (N_640,N_529,N_472);
and U641 (N_641,N_569,N_494);
nand U642 (N_642,N_456,N_516);
nor U643 (N_643,N_526,N_437);
nand U644 (N_644,N_520,N_507);
nand U645 (N_645,N_523,N_444);
and U646 (N_646,N_425,N_536);
nor U647 (N_647,N_462,N_422);
nand U648 (N_648,N_407,N_479);
nor U649 (N_649,N_438,N_461);
and U650 (N_650,N_574,N_432);
nor U651 (N_651,N_522,N_588);
and U652 (N_652,N_457,N_535);
nand U653 (N_653,N_478,N_548);
and U654 (N_654,N_580,N_466);
and U655 (N_655,N_563,N_488);
nor U656 (N_656,N_560,N_467);
nor U657 (N_657,N_573,N_468);
nor U658 (N_658,N_514,N_426);
nand U659 (N_659,N_572,N_405);
nand U660 (N_660,N_571,N_411);
or U661 (N_661,N_475,N_540);
nand U662 (N_662,N_581,N_402);
and U663 (N_663,N_513,N_403);
or U664 (N_664,N_531,N_592);
xnor U665 (N_665,N_595,N_598);
and U666 (N_666,N_431,N_455);
or U667 (N_667,N_413,N_439);
nor U668 (N_668,N_400,N_484);
or U669 (N_669,N_599,N_528);
or U670 (N_670,N_530,N_589);
or U671 (N_671,N_410,N_473);
nand U672 (N_672,N_476,N_459);
and U673 (N_673,N_482,N_480);
nor U674 (N_674,N_582,N_408);
or U675 (N_675,N_534,N_504);
nor U676 (N_676,N_509,N_533);
and U677 (N_677,N_401,N_542);
nand U678 (N_678,N_433,N_423);
or U679 (N_679,N_556,N_441);
and U680 (N_680,N_498,N_506);
or U681 (N_681,N_453,N_587);
nor U682 (N_682,N_510,N_567);
or U683 (N_683,N_418,N_497);
nand U684 (N_684,N_543,N_463);
or U685 (N_685,N_517,N_445);
nand U686 (N_686,N_584,N_545);
nor U687 (N_687,N_547,N_577);
nand U688 (N_688,N_489,N_512);
or U689 (N_689,N_553,N_416);
or U690 (N_690,N_539,N_409);
and U691 (N_691,N_549,N_442);
xor U692 (N_692,N_551,N_436);
nand U693 (N_693,N_454,N_524);
nor U694 (N_694,N_511,N_448);
nor U695 (N_695,N_490,N_505);
or U696 (N_696,N_564,N_583);
nor U697 (N_697,N_579,N_424);
and U698 (N_698,N_474,N_538);
nor U699 (N_699,N_561,N_460);
xor U700 (N_700,N_503,N_552);
nand U701 (N_701,N_522,N_405);
nor U702 (N_702,N_469,N_453);
nand U703 (N_703,N_534,N_549);
or U704 (N_704,N_405,N_504);
nor U705 (N_705,N_424,N_519);
and U706 (N_706,N_444,N_458);
or U707 (N_707,N_495,N_564);
nand U708 (N_708,N_455,N_591);
or U709 (N_709,N_406,N_533);
and U710 (N_710,N_448,N_590);
nor U711 (N_711,N_591,N_409);
or U712 (N_712,N_417,N_574);
nor U713 (N_713,N_411,N_524);
nor U714 (N_714,N_488,N_452);
nor U715 (N_715,N_550,N_485);
nand U716 (N_716,N_434,N_422);
xor U717 (N_717,N_496,N_415);
or U718 (N_718,N_582,N_492);
nor U719 (N_719,N_460,N_590);
or U720 (N_720,N_428,N_414);
nor U721 (N_721,N_534,N_509);
or U722 (N_722,N_425,N_558);
xor U723 (N_723,N_521,N_438);
xor U724 (N_724,N_579,N_470);
nand U725 (N_725,N_549,N_458);
or U726 (N_726,N_598,N_580);
or U727 (N_727,N_513,N_483);
nand U728 (N_728,N_423,N_570);
nor U729 (N_729,N_500,N_566);
and U730 (N_730,N_409,N_438);
or U731 (N_731,N_469,N_439);
nand U732 (N_732,N_569,N_562);
and U733 (N_733,N_454,N_495);
or U734 (N_734,N_447,N_498);
and U735 (N_735,N_428,N_480);
nor U736 (N_736,N_465,N_458);
or U737 (N_737,N_597,N_457);
nor U738 (N_738,N_593,N_489);
and U739 (N_739,N_443,N_470);
or U740 (N_740,N_505,N_467);
nor U741 (N_741,N_540,N_481);
and U742 (N_742,N_475,N_497);
nor U743 (N_743,N_577,N_511);
nand U744 (N_744,N_546,N_525);
and U745 (N_745,N_503,N_538);
nor U746 (N_746,N_508,N_461);
and U747 (N_747,N_441,N_511);
nor U748 (N_748,N_582,N_512);
nand U749 (N_749,N_506,N_532);
nand U750 (N_750,N_474,N_482);
nand U751 (N_751,N_541,N_546);
and U752 (N_752,N_552,N_525);
or U753 (N_753,N_421,N_503);
and U754 (N_754,N_478,N_493);
nand U755 (N_755,N_411,N_565);
and U756 (N_756,N_501,N_572);
nand U757 (N_757,N_406,N_445);
nor U758 (N_758,N_436,N_565);
nor U759 (N_759,N_571,N_475);
nand U760 (N_760,N_554,N_488);
nand U761 (N_761,N_558,N_596);
or U762 (N_762,N_475,N_424);
nor U763 (N_763,N_467,N_444);
nor U764 (N_764,N_490,N_502);
nor U765 (N_765,N_536,N_522);
or U766 (N_766,N_465,N_569);
and U767 (N_767,N_559,N_506);
nor U768 (N_768,N_568,N_416);
and U769 (N_769,N_513,N_465);
or U770 (N_770,N_578,N_410);
or U771 (N_771,N_457,N_464);
nor U772 (N_772,N_496,N_400);
nand U773 (N_773,N_457,N_548);
or U774 (N_774,N_497,N_478);
or U775 (N_775,N_437,N_597);
nand U776 (N_776,N_461,N_496);
and U777 (N_777,N_536,N_587);
and U778 (N_778,N_577,N_401);
nor U779 (N_779,N_467,N_550);
and U780 (N_780,N_442,N_591);
nor U781 (N_781,N_496,N_564);
nand U782 (N_782,N_465,N_583);
nor U783 (N_783,N_420,N_467);
nor U784 (N_784,N_486,N_469);
nand U785 (N_785,N_476,N_451);
or U786 (N_786,N_572,N_490);
nor U787 (N_787,N_468,N_412);
and U788 (N_788,N_519,N_575);
xnor U789 (N_789,N_597,N_580);
nor U790 (N_790,N_564,N_443);
or U791 (N_791,N_427,N_496);
or U792 (N_792,N_471,N_446);
or U793 (N_793,N_401,N_462);
xor U794 (N_794,N_414,N_477);
or U795 (N_795,N_574,N_523);
and U796 (N_796,N_462,N_500);
and U797 (N_797,N_535,N_471);
nand U798 (N_798,N_461,N_460);
or U799 (N_799,N_531,N_459);
or U800 (N_800,N_614,N_762);
or U801 (N_801,N_742,N_667);
nor U802 (N_802,N_746,N_787);
and U803 (N_803,N_726,N_773);
nor U804 (N_804,N_711,N_750);
or U805 (N_805,N_691,N_791);
nand U806 (N_806,N_648,N_702);
nor U807 (N_807,N_722,N_649);
nand U808 (N_808,N_724,N_659);
and U809 (N_809,N_754,N_658);
nand U810 (N_810,N_671,N_707);
or U811 (N_811,N_715,N_697);
nor U812 (N_812,N_605,N_765);
or U813 (N_813,N_731,N_768);
nand U814 (N_814,N_734,N_651);
or U815 (N_815,N_736,N_797);
nand U816 (N_816,N_607,N_712);
and U817 (N_817,N_680,N_673);
or U818 (N_818,N_704,N_662);
nand U819 (N_819,N_727,N_627);
and U820 (N_820,N_661,N_632);
or U821 (N_821,N_799,N_771);
or U822 (N_822,N_678,N_749);
nand U823 (N_823,N_751,N_774);
nor U824 (N_824,N_626,N_725);
and U825 (N_825,N_669,N_728);
and U826 (N_826,N_792,N_689);
nand U827 (N_827,N_709,N_675);
nand U828 (N_828,N_781,N_753);
or U829 (N_829,N_732,N_793);
and U830 (N_830,N_688,N_796);
and U831 (N_831,N_770,N_747);
or U832 (N_832,N_795,N_716);
or U833 (N_833,N_660,N_759);
nand U834 (N_834,N_636,N_763);
nand U835 (N_835,N_777,N_694);
or U836 (N_836,N_786,N_679);
and U837 (N_837,N_601,N_729);
nand U838 (N_838,N_790,N_618);
and U839 (N_839,N_630,N_617);
and U840 (N_840,N_681,N_776);
nand U841 (N_841,N_755,N_612);
and U842 (N_842,N_672,N_609);
or U843 (N_843,N_625,N_700);
nor U844 (N_844,N_647,N_708);
and U845 (N_845,N_615,N_705);
and U846 (N_846,N_757,N_611);
nor U847 (N_847,N_686,N_695);
nand U848 (N_848,N_703,N_758);
and U849 (N_849,N_794,N_645);
or U850 (N_850,N_655,N_687);
nand U851 (N_851,N_606,N_782);
nand U852 (N_852,N_644,N_616);
and U853 (N_853,N_699,N_785);
nand U854 (N_854,N_682,N_684);
or U855 (N_855,N_798,N_643);
or U856 (N_856,N_769,N_745);
nand U857 (N_857,N_657,N_635);
nand U858 (N_858,N_772,N_720);
or U859 (N_859,N_760,N_637);
nor U860 (N_860,N_652,N_641);
and U861 (N_861,N_628,N_650);
nor U862 (N_862,N_783,N_600);
nand U863 (N_863,N_775,N_743);
and U864 (N_864,N_719,N_698);
and U865 (N_865,N_621,N_610);
xor U866 (N_866,N_717,N_718);
nand U867 (N_867,N_654,N_608);
nor U868 (N_868,N_623,N_767);
or U869 (N_869,N_706,N_741);
or U870 (N_870,N_696,N_676);
nand U871 (N_871,N_735,N_714);
nor U872 (N_872,N_788,N_710);
nor U873 (N_873,N_646,N_737);
nand U874 (N_874,N_665,N_664);
nand U875 (N_875,N_764,N_730);
nand U876 (N_876,N_778,N_701);
and U877 (N_877,N_723,N_603);
and U878 (N_878,N_633,N_789);
and U879 (N_879,N_748,N_739);
nor U880 (N_880,N_638,N_602);
nand U881 (N_881,N_653,N_620);
nor U882 (N_882,N_631,N_690);
and U883 (N_883,N_752,N_634);
and U884 (N_884,N_639,N_668);
or U885 (N_885,N_656,N_613);
and U886 (N_886,N_622,N_604);
xor U887 (N_887,N_761,N_766);
nand U888 (N_888,N_721,N_663);
nand U889 (N_889,N_640,N_642);
and U890 (N_890,N_670,N_683);
or U891 (N_891,N_624,N_740);
nand U892 (N_892,N_629,N_713);
nor U893 (N_893,N_779,N_756);
nand U894 (N_894,N_784,N_738);
nand U895 (N_895,N_780,N_692);
nand U896 (N_896,N_693,N_744);
nand U897 (N_897,N_733,N_666);
and U898 (N_898,N_685,N_674);
and U899 (N_899,N_677,N_619);
nor U900 (N_900,N_749,N_748);
or U901 (N_901,N_635,N_794);
nor U902 (N_902,N_752,N_651);
nor U903 (N_903,N_732,N_658);
and U904 (N_904,N_666,N_649);
or U905 (N_905,N_776,N_602);
and U906 (N_906,N_601,N_673);
nor U907 (N_907,N_672,N_665);
nor U908 (N_908,N_732,N_684);
nand U909 (N_909,N_739,N_710);
or U910 (N_910,N_775,N_645);
and U911 (N_911,N_656,N_705);
nand U912 (N_912,N_669,N_684);
or U913 (N_913,N_772,N_612);
or U914 (N_914,N_782,N_655);
or U915 (N_915,N_686,N_670);
nor U916 (N_916,N_617,N_740);
xnor U917 (N_917,N_709,N_716);
nor U918 (N_918,N_660,N_699);
or U919 (N_919,N_756,N_621);
and U920 (N_920,N_775,N_720);
nor U921 (N_921,N_691,N_717);
and U922 (N_922,N_732,N_656);
and U923 (N_923,N_757,N_742);
nor U924 (N_924,N_666,N_702);
nor U925 (N_925,N_744,N_753);
or U926 (N_926,N_769,N_756);
nor U927 (N_927,N_777,N_704);
or U928 (N_928,N_672,N_662);
and U929 (N_929,N_701,N_611);
or U930 (N_930,N_650,N_671);
and U931 (N_931,N_776,N_788);
nand U932 (N_932,N_650,N_703);
or U933 (N_933,N_726,N_782);
and U934 (N_934,N_651,N_700);
or U935 (N_935,N_760,N_778);
nor U936 (N_936,N_776,N_773);
or U937 (N_937,N_663,N_738);
or U938 (N_938,N_736,N_752);
nand U939 (N_939,N_688,N_660);
nor U940 (N_940,N_616,N_721);
or U941 (N_941,N_678,N_799);
nand U942 (N_942,N_635,N_759);
and U943 (N_943,N_617,N_744);
and U944 (N_944,N_750,N_796);
or U945 (N_945,N_772,N_618);
nand U946 (N_946,N_721,N_796);
and U947 (N_947,N_792,N_747);
and U948 (N_948,N_629,N_644);
and U949 (N_949,N_601,N_668);
nand U950 (N_950,N_762,N_646);
nand U951 (N_951,N_693,N_751);
or U952 (N_952,N_794,N_605);
and U953 (N_953,N_706,N_720);
and U954 (N_954,N_637,N_657);
nand U955 (N_955,N_694,N_788);
nand U956 (N_956,N_724,N_656);
nor U957 (N_957,N_635,N_724);
nand U958 (N_958,N_709,N_696);
nand U959 (N_959,N_751,N_757);
and U960 (N_960,N_763,N_689);
nor U961 (N_961,N_609,N_761);
and U962 (N_962,N_773,N_631);
and U963 (N_963,N_672,N_669);
nand U964 (N_964,N_679,N_672);
nand U965 (N_965,N_603,N_799);
or U966 (N_966,N_675,N_616);
or U967 (N_967,N_707,N_753);
nand U968 (N_968,N_662,N_710);
or U969 (N_969,N_799,N_623);
or U970 (N_970,N_637,N_676);
and U971 (N_971,N_643,N_700);
nand U972 (N_972,N_768,N_744);
nor U973 (N_973,N_761,N_659);
and U974 (N_974,N_648,N_683);
and U975 (N_975,N_697,N_764);
or U976 (N_976,N_666,N_601);
nor U977 (N_977,N_728,N_761);
or U978 (N_978,N_743,N_731);
and U979 (N_979,N_674,N_602);
nand U980 (N_980,N_668,N_709);
nor U981 (N_981,N_664,N_693);
nand U982 (N_982,N_630,N_658);
nor U983 (N_983,N_672,N_729);
and U984 (N_984,N_774,N_698);
nor U985 (N_985,N_768,N_725);
or U986 (N_986,N_735,N_637);
or U987 (N_987,N_731,N_662);
nor U988 (N_988,N_756,N_784);
and U989 (N_989,N_769,N_785);
xor U990 (N_990,N_606,N_641);
nor U991 (N_991,N_779,N_680);
or U992 (N_992,N_732,N_790);
nor U993 (N_993,N_722,N_735);
nand U994 (N_994,N_703,N_715);
xor U995 (N_995,N_666,N_713);
or U996 (N_996,N_777,N_779);
nand U997 (N_997,N_712,N_782);
and U998 (N_998,N_755,N_669);
xnor U999 (N_999,N_659,N_792);
or U1000 (N_1000,N_916,N_893);
or U1001 (N_1001,N_865,N_828);
and U1002 (N_1002,N_856,N_859);
xor U1003 (N_1003,N_963,N_988);
nand U1004 (N_1004,N_940,N_817);
nand U1005 (N_1005,N_956,N_800);
and U1006 (N_1006,N_863,N_926);
or U1007 (N_1007,N_880,N_972);
and U1008 (N_1008,N_991,N_844);
and U1009 (N_1009,N_869,N_919);
and U1010 (N_1010,N_948,N_835);
and U1011 (N_1011,N_814,N_872);
nor U1012 (N_1012,N_962,N_876);
nand U1013 (N_1013,N_987,N_864);
or U1014 (N_1014,N_992,N_946);
nand U1015 (N_1015,N_917,N_974);
xor U1016 (N_1016,N_808,N_895);
or U1017 (N_1017,N_845,N_954);
nand U1018 (N_1018,N_887,N_997);
xor U1019 (N_1019,N_961,N_831);
nor U1020 (N_1020,N_878,N_951);
nand U1021 (N_1021,N_857,N_965);
and U1022 (N_1022,N_952,N_839);
nor U1023 (N_1023,N_821,N_907);
nand U1024 (N_1024,N_904,N_927);
nor U1025 (N_1025,N_882,N_801);
nor U1026 (N_1026,N_899,N_838);
xnor U1027 (N_1027,N_822,N_999);
nor U1028 (N_1028,N_861,N_906);
nor U1029 (N_1029,N_829,N_982);
nand U1030 (N_1030,N_921,N_943);
nor U1031 (N_1031,N_812,N_891);
or U1032 (N_1032,N_881,N_925);
nand U1033 (N_1033,N_932,N_815);
and U1034 (N_1034,N_967,N_873);
nor U1035 (N_1035,N_848,N_884);
and U1036 (N_1036,N_910,N_842);
and U1037 (N_1037,N_923,N_911);
nand U1038 (N_1038,N_913,N_939);
nor U1039 (N_1039,N_826,N_930);
nor U1040 (N_1040,N_854,N_840);
nand U1041 (N_1041,N_901,N_823);
nand U1042 (N_1042,N_998,N_806);
and U1043 (N_1043,N_849,N_900);
or U1044 (N_1044,N_970,N_903);
and U1045 (N_1045,N_983,N_964);
or U1046 (N_1046,N_888,N_867);
or U1047 (N_1047,N_986,N_990);
nor U1048 (N_1048,N_994,N_949);
nor U1049 (N_1049,N_920,N_804);
or U1050 (N_1050,N_915,N_933);
nor U1051 (N_1051,N_894,N_892);
and U1052 (N_1052,N_968,N_810);
nor U1053 (N_1053,N_996,N_837);
nor U1054 (N_1054,N_832,N_908);
nor U1055 (N_1055,N_862,N_860);
or U1056 (N_1056,N_905,N_825);
or U1057 (N_1057,N_942,N_813);
nand U1058 (N_1058,N_834,N_980);
or U1059 (N_1059,N_824,N_977);
or U1060 (N_1060,N_886,N_805);
and U1061 (N_1061,N_816,N_879);
nand U1062 (N_1062,N_885,N_827);
or U1063 (N_1063,N_938,N_936);
and U1064 (N_1064,N_978,N_833);
or U1065 (N_1065,N_960,N_924);
nor U1066 (N_1066,N_937,N_981);
or U1067 (N_1067,N_803,N_847);
and U1068 (N_1068,N_928,N_818);
and U1069 (N_1069,N_870,N_985);
nand U1070 (N_1070,N_896,N_971);
or U1071 (N_1071,N_989,N_958);
and U1072 (N_1072,N_807,N_897);
nand U1073 (N_1073,N_874,N_802);
nor U1074 (N_1074,N_950,N_866);
nand U1075 (N_1075,N_877,N_955);
and U1076 (N_1076,N_850,N_973);
nor U1077 (N_1077,N_852,N_858);
or U1078 (N_1078,N_935,N_898);
nor U1079 (N_1079,N_912,N_853);
or U1080 (N_1080,N_909,N_969);
and U1081 (N_1081,N_922,N_889);
nor U1082 (N_1082,N_941,N_966);
nand U1083 (N_1083,N_890,N_868);
and U1084 (N_1084,N_959,N_975);
or U1085 (N_1085,N_995,N_843);
or U1086 (N_1086,N_855,N_851);
nor U1087 (N_1087,N_947,N_841);
and U1088 (N_1088,N_931,N_984);
nor U1089 (N_1089,N_945,N_918);
nor U1090 (N_1090,N_929,N_846);
xor U1091 (N_1091,N_875,N_871);
and U1092 (N_1092,N_953,N_934);
and U1093 (N_1093,N_902,N_809);
nor U1094 (N_1094,N_914,N_957);
nand U1095 (N_1095,N_820,N_883);
and U1096 (N_1096,N_819,N_979);
nand U1097 (N_1097,N_976,N_836);
nand U1098 (N_1098,N_944,N_993);
or U1099 (N_1099,N_830,N_811);
nand U1100 (N_1100,N_892,N_966);
nand U1101 (N_1101,N_884,N_845);
nor U1102 (N_1102,N_943,N_808);
nor U1103 (N_1103,N_911,N_906);
or U1104 (N_1104,N_964,N_993);
and U1105 (N_1105,N_949,N_889);
nor U1106 (N_1106,N_839,N_945);
and U1107 (N_1107,N_895,N_924);
nand U1108 (N_1108,N_800,N_923);
nand U1109 (N_1109,N_975,N_964);
nand U1110 (N_1110,N_904,N_930);
nor U1111 (N_1111,N_886,N_986);
or U1112 (N_1112,N_830,N_902);
and U1113 (N_1113,N_989,N_994);
or U1114 (N_1114,N_959,N_956);
nor U1115 (N_1115,N_898,N_911);
or U1116 (N_1116,N_840,N_931);
and U1117 (N_1117,N_963,N_940);
nor U1118 (N_1118,N_993,N_988);
and U1119 (N_1119,N_904,N_882);
nor U1120 (N_1120,N_869,N_815);
and U1121 (N_1121,N_895,N_868);
nand U1122 (N_1122,N_848,N_849);
and U1123 (N_1123,N_918,N_888);
nor U1124 (N_1124,N_927,N_829);
nor U1125 (N_1125,N_906,N_833);
or U1126 (N_1126,N_976,N_945);
nand U1127 (N_1127,N_933,N_998);
nor U1128 (N_1128,N_885,N_952);
nand U1129 (N_1129,N_833,N_876);
nand U1130 (N_1130,N_830,N_849);
or U1131 (N_1131,N_955,N_962);
and U1132 (N_1132,N_910,N_999);
nor U1133 (N_1133,N_996,N_968);
nand U1134 (N_1134,N_903,N_990);
nand U1135 (N_1135,N_865,N_945);
and U1136 (N_1136,N_899,N_923);
and U1137 (N_1137,N_827,N_937);
nand U1138 (N_1138,N_822,N_993);
nand U1139 (N_1139,N_922,N_847);
or U1140 (N_1140,N_831,N_840);
nor U1141 (N_1141,N_895,N_939);
or U1142 (N_1142,N_999,N_896);
nand U1143 (N_1143,N_854,N_904);
and U1144 (N_1144,N_841,N_835);
or U1145 (N_1145,N_982,N_816);
and U1146 (N_1146,N_801,N_853);
or U1147 (N_1147,N_898,N_894);
nor U1148 (N_1148,N_858,N_828);
and U1149 (N_1149,N_876,N_985);
and U1150 (N_1150,N_945,N_989);
and U1151 (N_1151,N_856,N_968);
or U1152 (N_1152,N_864,N_917);
or U1153 (N_1153,N_960,N_991);
and U1154 (N_1154,N_812,N_999);
nand U1155 (N_1155,N_806,N_807);
or U1156 (N_1156,N_954,N_807);
nor U1157 (N_1157,N_927,N_915);
and U1158 (N_1158,N_958,N_898);
nand U1159 (N_1159,N_915,N_889);
nand U1160 (N_1160,N_843,N_909);
nor U1161 (N_1161,N_860,N_824);
nand U1162 (N_1162,N_881,N_803);
nand U1163 (N_1163,N_959,N_860);
or U1164 (N_1164,N_922,N_843);
or U1165 (N_1165,N_894,N_907);
nand U1166 (N_1166,N_886,N_947);
nand U1167 (N_1167,N_903,N_956);
nand U1168 (N_1168,N_836,N_937);
nand U1169 (N_1169,N_995,N_884);
nor U1170 (N_1170,N_886,N_983);
or U1171 (N_1171,N_866,N_924);
nand U1172 (N_1172,N_825,N_967);
nand U1173 (N_1173,N_986,N_805);
and U1174 (N_1174,N_864,N_923);
or U1175 (N_1175,N_858,N_831);
and U1176 (N_1176,N_900,N_962);
nor U1177 (N_1177,N_908,N_831);
and U1178 (N_1178,N_883,N_998);
or U1179 (N_1179,N_914,N_839);
nor U1180 (N_1180,N_889,N_956);
nor U1181 (N_1181,N_996,N_804);
or U1182 (N_1182,N_873,N_805);
and U1183 (N_1183,N_850,N_825);
or U1184 (N_1184,N_963,N_952);
nor U1185 (N_1185,N_961,N_929);
nand U1186 (N_1186,N_985,N_962);
xnor U1187 (N_1187,N_950,N_867);
or U1188 (N_1188,N_979,N_873);
nand U1189 (N_1189,N_996,N_913);
nor U1190 (N_1190,N_967,N_903);
nand U1191 (N_1191,N_868,N_939);
or U1192 (N_1192,N_995,N_900);
nor U1193 (N_1193,N_992,N_977);
and U1194 (N_1194,N_896,N_885);
nand U1195 (N_1195,N_938,N_844);
nand U1196 (N_1196,N_817,N_942);
nand U1197 (N_1197,N_867,N_916);
and U1198 (N_1198,N_917,N_889);
nand U1199 (N_1199,N_991,N_854);
and U1200 (N_1200,N_1036,N_1139);
or U1201 (N_1201,N_1146,N_1025);
and U1202 (N_1202,N_1045,N_1097);
nor U1203 (N_1203,N_1113,N_1166);
or U1204 (N_1204,N_1015,N_1073);
nor U1205 (N_1205,N_1169,N_1178);
and U1206 (N_1206,N_1168,N_1083);
or U1207 (N_1207,N_1125,N_1082);
nand U1208 (N_1208,N_1181,N_1034);
or U1209 (N_1209,N_1140,N_1011);
or U1210 (N_1210,N_1000,N_1076);
or U1211 (N_1211,N_1163,N_1198);
or U1212 (N_1212,N_1191,N_1131);
nand U1213 (N_1213,N_1144,N_1035);
and U1214 (N_1214,N_1127,N_1180);
nand U1215 (N_1215,N_1040,N_1137);
nand U1216 (N_1216,N_1043,N_1179);
nand U1217 (N_1217,N_1155,N_1121);
or U1218 (N_1218,N_1154,N_1012);
or U1219 (N_1219,N_1192,N_1152);
and U1220 (N_1220,N_1105,N_1069);
or U1221 (N_1221,N_1138,N_1136);
xor U1222 (N_1222,N_1128,N_1157);
and U1223 (N_1223,N_1088,N_1183);
or U1224 (N_1224,N_1053,N_1106);
or U1225 (N_1225,N_1118,N_1081);
nand U1226 (N_1226,N_1129,N_1078);
nand U1227 (N_1227,N_1020,N_1061);
and U1228 (N_1228,N_1063,N_1075);
or U1229 (N_1229,N_1182,N_1159);
nor U1230 (N_1230,N_1112,N_1199);
nand U1231 (N_1231,N_1017,N_1005);
and U1232 (N_1232,N_1188,N_1089);
and U1233 (N_1233,N_1109,N_1077);
or U1234 (N_1234,N_1156,N_1060);
nand U1235 (N_1235,N_1018,N_1067);
xnor U1236 (N_1236,N_1165,N_1068);
or U1237 (N_1237,N_1193,N_1009);
or U1238 (N_1238,N_1126,N_1044);
nand U1239 (N_1239,N_1119,N_1132);
xor U1240 (N_1240,N_1029,N_1087);
nor U1241 (N_1241,N_1133,N_1101);
nand U1242 (N_1242,N_1189,N_1064);
and U1243 (N_1243,N_1158,N_1123);
or U1244 (N_1244,N_1026,N_1177);
nand U1245 (N_1245,N_1066,N_1028);
or U1246 (N_1246,N_1037,N_1104);
nand U1247 (N_1247,N_1173,N_1098);
and U1248 (N_1248,N_1038,N_1055);
or U1249 (N_1249,N_1116,N_1008);
or U1250 (N_1250,N_1184,N_1016);
and U1251 (N_1251,N_1002,N_1031);
nor U1252 (N_1252,N_1046,N_1145);
or U1253 (N_1253,N_1122,N_1095);
nand U1254 (N_1254,N_1047,N_1007);
and U1255 (N_1255,N_1194,N_1057);
nor U1256 (N_1256,N_1141,N_1174);
or U1257 (N_1257,N_1090,N_1071);
or U1258 (N_1258,N_1092,N_1149);
and U1259 (N_1259,N_1187,N_1041);
and U1260 (N_1260,N_1062,N_1065);
nand U1261 (N_1261,N_1171,N_1019);
and U1262 (N_1262,N_1059,N_1124);
and U1263 (N_1263,N_1052,N_1110);
or U1264 (N_1264,N_1004,N_1084);
nor U1265 (N_1265,N_1014,N_1048);
nor U1266 (N_1266,N_1001,N_1054);
nor U1267 (N_1267,N_1024,N_1197);
nand U1268 (N_1268,N_1080,N_1027);
or U1269 (N_1269,N_1134,N_1111);
nor U1270 (N_1270,N_1190,N_1162);
and U1271 (N_1271,N_1058,N_1070);
or U1272 (N_1272,N_1039,N_1051);
and U1273 (N_1273,N_1170,N_1143);
nand U1274 (N_1274,N_1006,N_1079);
and U1275 (N_1275,N_1196,N_1120);
and U1276 (N_1276,N_1086,N_1023);
nor U1277 (N_1277,N_1167,N_1003);
nor U1278 (N_1278,N_1185,N_1091);
nand U1279 (N_1279,N_1010,N_1099);
and U1280 (N_1280,N_1103,N_1176);
nand U1281 (N_1281,N_1150,N_1195);
nor U1282 (N_1282,N_1050,N_1115);
and U1283 (N_1283,N_1142,N_1093);
xor U1284 (N_1284,N_1033,N_1074);
or U1285 (N_1285,N_1107,N_1186);
or U1286 (N_1286,N_1032,N_1022);
or U1287 (N_1287,N_1100,N_1094);
xor U1288 (N_1288,N_1096,N_1102);
nor U1289 (N_1289,N_1021,N_1161);
and U1290 (N_1290,N_1172,N_1130);
nand U1291 (N_1291,N_1153,N_1049);
nor U1292 (N_1292,N_1042,N_1114);
nand U1293 (N_1293,N_1117,N_1135);
xor U1294 (N_1294,N_1108,N_1013);
nor U1295 (N_1295,N_1147,N_1056);
nand U1296 (N_1296,N_1160,N_1175);
or U1297 (N_1297,N_1148,N_1085);
and U1298 (N_1298,N_1151,N_1164);
or U1299 (N_1299,N_1072,N_1030);
and U1300 (N_1300,N_1078,N_1031);
and U1301 (N_1301,N_1031,N_1022);
nand U1302 (N_1302,N_1015,N_1027);
nand U1303 (N_1303,N_1166,N_1029);
nand U1304 (N_1304,N_1023,N_1112);
nand U1305 (N_1305,N_1067,N_1153);
and U1306 (N_1306,N_1184,N_1139);
nor U1307 (N_1307,N_1195,N_1020);
or U1308 (N_1308,N_1030,N_1033);
nand U1309 (N_1309,N_1069,N_1128);
or U1310 (N_1310,N_1135,N_1120);
and U1311 (N_1311,N_1010,N_1066);
and U1312 (N_1312,N_1176,N_1129);
nor U1313 (N_1313,N_1024,N_1131);
nand U1314 (N_1314,N_1093,N_1105);
nor U1315 (N_1315,N_1013,N_1143);
and U1316 (N_1316,N_1102,N_1051);
or U1317 (N_1317,N_1009,N_1151);
and U1318 (N_1318,N_1071,N_1104);
nand U1319 (N_1319,N_1160,N_1051);
and U1320 (N_1320,N_1158,N_1050);
or U1321 (N_1321,N_1023,N_1142);
and U1322 (N_1322,N_1156,N_1062);
or U1323 (N_1323,N_1124,N_1046);
and U1324 (N_1324,N_1107,N_1076);
and U1325 (N_1325,N_1140,N_1176);
nand U1326 (N_1326,N_1155,N_1067);
nor U1327 (N_1327,N_1020,N_1184);
or U1328 (N_1328,N_1148,N_1109);
nand U1329 (N_1329,N_1155,N_1012);
or U1330 (N_1330,N_1056,N_1135);
nor U1331 (N_1331,N_1147,N_1086);
and U1332 (N_1332,N_1025,N_1188);
nand U1333 (N_1333,N_1167,N_1109);
nand U1334 (N_1334,N_1000,N_1004);
or U1335 (N_1335,N_1108,N_1156);
or U1336 (N_1336,N_1057,N_1082);
nor U1337 (N_1337,N_1013,N_1174);
or U1338 (N_1338,N_1175,N_1062);
nor U1339 (N_1339,N_1017,N_1091);
nor U1340 (N_1340,N_1036,N_1002);
nand U1341 (N_1341,N_1076,N_1125);
nand U1342 (N_1342,N_1197,N_1167);
nand U1343 (N_1343,N_1026,N_1046);
or U1344 (N_1344,N_1121,N_1148);
nand U1345 (N_1345,N_1065,N_1147);
and U1346 (N_1346,N_1038,N_1080);
and U1347 (N_1347,N_1088,N_1120);
and U1348 (N_1348,N_1122,N_1185);
or U1349 (N_1349,N_1159,N_1191);
and U1350 (N_1350,N_1189,N_1088);
and U1351 (N_1351,N_1148,N_1129);
nor U1352 (N_1352,N_1160,N_1082);
and U1353 (N_1353,N_1120,N_1128);
and U1354 (N_1354,N_1051,N_1145);
nor U1355 (N_1355,N_1047,N_1039);
nor U1356 (N_1356,N_1078,N_1052);
nor U1357 (N_1357,N_1190,N_1053);
nand U1358 (N_1358,N_1089,N_1020);
and U1359 (N_1359,N_1023,N_1017);
nor U1360 (N_1360,N_1068,N_1133);
or U1361 (N_1361,N_1097,N_1009);
and U1362 (N_1362,N_1012,N_1065);
or U1363 (N_1363,N_1157,N_1056);
or U1364 (N_1364,N_1097,N_1165);
and U1365 (N_1365,N_1175,N_1016);
nor U1366 (N_1366,N_1082,N_1187);
and U1367 (N_1367,N_1055,N_1107);
nor U1368 (N_1368,N_1004,N_1056);
nor U1369 (N_1369,N_1111,N_1075);
and U1370 (N_1370,N_1021,N_1047);
nor U1371 (N_1371,N_1078,N_1050);
nand U1372 (N_1372,N_1133,N_1056);
nor U1373 (N_1373,N_1167,N_1006);
and U1374 (N_1374,N_1007,N_1184);
or U1375 (N_1375,N_1050,N_1076);
and U1376 (N_1376,N_1127,N_1185);
nor U1377 (N_1377,N_1113,N_1120);
nor U1378 (N_1378,N_1069,N_1154);
nor U1379 (N_1379,N_1130,N_1095);
and U1380 (N_1380,N_1040,N_1170);
nand U1381 (N_1381,N_1193,N_1153);
nand U1382 (N_1382,N_1047,N_1124);
or U1383 (N_1383,N_1155,N_1187);
nand U1384 (N_1384,N_1112,N_1122);
or U1385 (N_1385,N_1046,N_1123);
nand U1386 (N_1386,N_1142,N_1040);
nor U1387 (N_1387,N_1188,N_1097);
or U1388 (N_1388,N_1193,N_1154);
nor U1389 (N_1389,N_1151,N_1183);
nor U1390 (N_1390,N_1178,N_1040);
nor U1391 (N_1391,N_1052,N_1109);
nand U1392 (N_1392,N_1036,N_1044);
nor U1393 (N_1393,N_1173,N_1012);
and U1394 (N_1394,N_1154,N_1196);
nand U1395 (N_1395,N_1118,N_1060);
or U1396 (N_1396,N_1121,N_1126);
xnor U1397 (N_1397,N_1158,N_1133);
nor U1398 (N_1398,N_1079,N_1186);
and U1399 (N_1399,N_1051,N_1038);
and U1400 (N_1400,N_1383,N_1327);
nor U1401 (N_1401,N_1365,N_1384);
nor U1402 (N_1402,N_1257,N_1289);
and U1403 (N_1403,N_1337,N_1261);
and U1404 (N_1404,N_1309,N_1204);
or U1405 (N_1405,N_1336,N_1276);
and U1406 (N_1406,N_1329,N_1360);
nor U1407 (N_1407,N_1251,N_1260);
nand U1408 (N_1408,N_1313,N_1215);
nor U1409 (N_1409,N_1208,N_1326);
or U1410 (N_1410,N_1382,N_1332);
xor U1411 (N_1411,N_1293,N_1268);
or U1412 (N_1412,N_1248,N_1224);
and U1413 (N_1413,N_1279,N_1380);
xnor U1414 (N_1414,N_1240,N_1294);
nand U1415 (N_1415,N_1223,N_1316);
and U1416 (N_1416,N_1236,N_1394);
nor U1417 (N_1417,N_1282,N_1302);
nor U1418 (N_1418,N_1271,N_1207);
nand U1419 (N_1419,N_1263,N_1232);
and U1420 (N_1420,N_1387,N_1391);
and U1421 (N_1421,N_1209,N_1255);
or U1422 (N_1422,N_1392,N_1395);
nor U1423 (N_1423,N_1375,N_1398);
or U1424 (N_1424,N_1212,N_1367);
nor U1425 (N_1425,N_1390,N_1333);
nor U1426 (N_1426,N_1311,N_1350);
and U1427 (N_1427,N_1330,N_1389);
and U1428 (N_1428,N_1272,N_1287);
or U1429 (N_1429,N_1300,N_1277);
nor U1430 (N_1430,N_1364,N_1220);
nand U1431 (N_1431,N_1270,N_1331);
nand U1432 (N_1432,N_1379,N_1250);
xor U1433 (N_1433,N_1227,N_1328);
and U1434 (N_1434,N_1352,N_1319);
nand U1435 (N_1435,N_1292,N_1299);
and U1436 (N_1436,N_1325,N_1310);
nand U1437 (N_1437,N_1372,N_1338);
and U1438 (N_1438,N_1211,N_1200);
and U1439 (N_1439,N_1393,N_1348);
nand U1440 (N_1440,N_1388,N_1249);
and U1441 (N_1441,N_1317,N_1222);
xor U1442 (N_1442,N_1245,N_1219);
and U1443 (N_1443,N_1347,N_1345);
nor U1444 (N_1444,N_1266,N_1386);
nand U1445 (N_1445,N_1253,N_1396);
nor U1446 (N_1446,N_1262,N_1363);
and U1447 (N_1447,N_1301,N_1286);
and U1448 (N_1448,N_1290,N_1339);
nand U1449 (N_1449,N_1320,N_1314);
nor U1450 (N_1450,N_1296,N_1228);
or U1451 (N_1451,N_1381,N_1259);
or U1452 (N_1452,N_1340,N_1354);
or U1453 (N_1453,N_1335,N_1291);
nor U1454 (N_1454,N_1288,N_1237);
or U1455 (N_1455,N_1210,N_1217);
nand U1456 (N_1456,N_1283,N_1298);
xor U1457 (N_1457,N_1233,N_1371);
nand U1458 (N_1458,N_1218,N_1346);
or U1459 (N_1459,N_1284,N_1213);
nand U1460 (N_1460,N_1201,N_1343);
nor U1461 (N_1461,N_1369,N_1357);
nand U1462 (N_1462,N_1376,N_1256);
nand U1463 (N_1463,N_1264,N_1362);
xor U1464 (N_1464,N_1221,N_1307);
or U1465 (N_1465,N_1214,N_1334);
nor U1466 (N_1466,N_1226,N_1374);
nand U1467 (N_1467,N_1274,N_1377);
and U1468 (N_1468,N_1359,N_1322);
and U1469 (N_1469,N_1355,N_1358);
nand U1470 (N_1470,N_1351,N_1370);
nand U1471 (N_1471,N_1303,N_1295);
or U1472 (N_1472,N_1399,N_1254);
or U1473 (N_1473,N_1203,N_1225);
nand U1474 (N_1474,N_1235,N_1281);
nand U1475 (N_1475,N_1285,N_1242);
nand U1476 (N_1476,N_1344,N_1378);
xor U1477 (N_1477,N_1206,N_1308);
nand U1478 (N_1478,N_1341,N_1368);
nor U1479 (N_1479,N_1239,N_1246);
or U1480 (N_1480,N_1252,N_1349);
nand U1481 (N_1481,N_1269,N_1273);
xnor U1482 (N_1482,N_1258,N_1321);
nor U1483 (N_1483,N_1366,N_1297);
nor U1484 (N_1484,N_1205,N_1305);
nor U1485 (N_1485,N_1361,N_1318);
nor U1486 (N_1486,N_1267,N_1306);
nand U1487 (N_1487,N_1241,N_1356);
and U1488 (N_1488,N_1234,N_1202);
nand U1489 (N_1489,N_1312,N_1216);
nand U1490 (N_1490,N_1304,N_1275);
or U1491 (N_1491,N_1244,N_1373);
nor U1492 (N_1492,N_1397,N_1265);
nand U1493 (N_1493,N_1230,N_1385);
and U1494 (N_1494,N_1231,N_1353);
nand U1495 (N_1495,N_1315,N_1278);
nand U1496 (N_1496,N_1243,N_1324);
nand U1497 (N_1497,N_1323,N_1238);
nor U1498 (N_1498,N_1229,N_1342);
nor U1499 (N_1499,N_1280,N_1247);
or U1500 (N_1500,N_1294,N_1346);
or U1501 (N_1501,N_1202,N_1255);
or U1502 (N_1502,N_1358,N_1235);
and U1503 (N_1503,N_1227,N_1302);
nor U1504 (N_1504,N_1320,N_1286);
nand U1505 (N_1505,N_1239,N_1379);
nor U1506 (N_1506,N_1226,N_1323);
and U1507 (N_1507,N_1205,N_1277);
nand U1508 (N_1508,N_1305,N_1250);
or U1509 (N_1509,N_1312,N_1393);
nand U1510 (N_1510,N_1367,N_1227);
nor U1511 (N_1511,N_1333,N_1222);
or U1512 (N_1512,N_1384,N_1344);
nand U1513 (N_1513,N_1335,N_1232);
nand U1514 (N_1514,N_1349,N_1242);
and U1515 (N_1515,N_1387,N_1214);
xnor U1516 (N_1516,N_1268,N_1265);
nand U1517 (N_1517,N_1249,N_1393);
nor U1518 (N_1518,N_1384,N_1358);
and U1519 (N_1519,N_1252,N_1258);
nand U1520 (N_1520,N_1208,N_1252);
or U1521 (N_1521,N_1258,N_1337);
or U1522 (N_1522,N_1314,N_1345);
and U1523 (N_1523,N_1211,N_1339);
nor U1524 (N_1524,N_1308,N_1245);
and U1525 (N_1525,N_1379,N_1216);
or U1526 (N_1526,N_1279,N_1246);
nand U1527 (N_1527,N_1304,N_1244);
nor U1528 (N_1528,N_1212,N_1280);
and U1529 (N_1529,N_1238,N_1303);
nand U1530 (N_1530,N_1243,N_1303);
and U1531 (N_1531,N_1270,N_1307);
nand U1532 (N_1532,N_1263,N_1398);
nor U1533 (N_1533,N_1255,N_1291);
nand U1534 (N_1534,N_1263,N_1271);
or U1535 (N_1535,N_1299,N_1286);
or U1536 (N_1536,N_1200,N_1386);
and U1537 (N_1537,N_1305,N_1370);
or U1538 (N_1538,N_1333,N_1218);
or U1539 (N_1539,N_1207,N_1326);
or U1540 (N_1540,N_1248,N_1334);
nor U1541 (N_1541,N_1247,N_1253);
or U1542 (N_1542,N_1382,N_1377);
and U1543 (N_1543,N_1272,N_1277);
nand U1544 (N_1544,N_1326,N_1293);
and U1545 (N_1545,N_1379,N_1316);
and U1546 (N_1546,N_1388,N_1284);
or U1547 (N_1547,N_1318,N_1388);
nor U1548 (N_1548,N_1398,N_1297);
and U1549 (N_1549,N_1348,N_1357);
and U1550 (N_1550,N_1232,N_1320);
or U1551 (N_1551,N_1239,N_1217);
and U1552 (N_1552,N_1384,N_1370);
and U1553 (N_1553,N_1293,N_1245);
or U1554 (N_1554,N_1209,N_1302);
or U1555 (N_1555,N_1225,N_1391);
xor U1556 (N_1556,N_1211,N_1220);
nor U1557 (N_1557,N_1353,N_1330);
or U1558 (N_1558,N_1287,N_1318);
nor U1559 (N_1559,N_1244,N_1381);
or U1560 (N_1560,N_1291,N_1251);
and U1561 (N_1561,N_1215,N_1252);
or U1562 (N_1562,N_1391,N_1236);
nand U1563 (N_1563,N_1364,N_1241);
nor U1564 (N_1564,N_1329,N_1247);
or U1565 (N_1565,N_1387,N_1323);
or U1566 (N_1566,N_1280,N_1210);
and U1567 (N_1567,N_1349,N_1378);
or U1568 (N_1568,N_1246,N_1270);
or U1569 (N_1569,N_1243,N_1267);
and U1570 (N_1570,N_1363,N_1274);
and U1571 (N_1571,N_1302,N_1314);
or U1572 (N_1572,N_1230,N_1341);
nand U1573 (N_1573,N_1348,N_1284);
and U1574 (N_1574,N_1336,N_1283);
and U1575 (N_1575,N_1258,N_1278);
or U1576 (N_1576,N_1205,N_1310);
and U1577 (N_1577,N_1230,N_1289);
nand U1578 (N_1578,N_1357,N_1206);
and U1579 (N_1579,N_1225,N_1284);
or U1580 (N_1580,N_1300,N_1394);
nor U1581 (N_1581,N_1304,N_1288);
nor U1582 (N_1582,N_1204,N_1317);
and U1583 (N_1583,N_1200,N_1245);
xnor U1584 (N_1584,N_1280,N_1267);
or U1585 (N_1585,N_1241,N_1239);
or U1586 (N_1586,N_1241,N_1295);
and U1587 (N_1587,N_1395,N_1326);
nand U1588 (N_1588,N_1244,N_1385);
and U1589 (N_1589,N_1340,N_1294);
nor U1590 (N_1590,N_1209,N_1324);
nand U1591 (N_1591,N_1293,N_1317);
nor U1592 (N_1592,N_1241,N_1318);
nand U1593 (N_1593,N_1269,N_1384);
nor U1594 (N_1594,N_1341,N_1303);
nand U1595 (N_1595,N_1269,N_1323);
nor U1596 (N_1596,N_1349,N_1206);
nand U1597 (N_1597,N_1362,N_1236);
or U1598 (N_1598,N_1227,N_1288);
nor U1599 (N_1599,N_1328,N_1295);
nand U1600 (N_1600,N_1491,N_1460);
nand U1601 (N_1601,N_1536,N_1587);
or U1602 (N_1602,N_1443,N_1465);
and U1603 (N_1603,N_1585,N_1597);
or U1604 (N_1604,N_1428,N_1412);
nand U1605 (N_1605,N_1568,N_1426);
nor U1606 (N_1606,N_1561,N_1575);
nand U1607 (N_1607,N_1478,N_1466);
or U1608 (N_1608,N_1554,N_1400);
nand U1609 (N_1609,N_1523,N_1446);
nor U1610 (N_1610,N_1545,N_1589);
nor U1611 (N_1611,N_1578,N_1504);
and U1612 (N_1612,N_1562,N_1419);
nor U1613 (N_1613,N_1517,N_1534);
and U1614 (N_1614,N_1579,N_1592);
and U1615 (N_1615,N_1512,N_1502);
or U1616 (N_1616,N_1548,N_1483);
xnor U1617 (N_1617,N_1450,N_1594);
and U1618 (N_1618,N_1401,N_1538);
and U1619 (N_1619,N_1557,N_1588);
xnor U1620 (N_1620,N_1529,N_1531);
nor U1621 (N_1621,N_1570,N_1429);
nor U1622 (N_1622,N_1447,N_1591);
nand U1623 (N_1623,N_1434,N_1449);
nor U1624 (N_1624,N_1406,N_1481);
nand U1625 (N_1625,N_1455,N_1461);
nand U1626 (N_1626,N_1537,N_1451);
or U1627 (N_1627,N_1532,N_1422);
nor U1628 (N_1628,N_1500,N_1555);
or U1629 (N_1629,N_1576,N_1431);
and U1630 (N_1630,N_1590,N_1509);
nand U1631 (N_1631,N_1402,N_1559);
nand U1632 (N_1632,N_1415,N_1490);
nor U1633 (N_1633,N_1563,N_1553);
nand U1634 (N_1634,N_1436,N_1598);
nor U1635 (N_1635,N_1586,N_1526);
nor U1636 (N_1636,N_1525,N_1540);
nor U1637 (N_1637,N_1417,N_1573);
or U1638 (N_1638,N_1433,N_1485);
or U1639 (N_1639,N_1445,N_1489);
or U1640 (N_1640,N_1518,N_1495);
and U1641 (N_1641,N_1499,N_1432);
nand U1642 (N_1642,N_1547,N_1410);
nor U1643 (N_1643,N_1498,N_1409);
nand U1644 (N_1644,N_1535,N_1533);
and U1645 (N_1645,N_1407,N_1497);
or U1646 (N_1646,N_1503,N_1564);
nor U1647 (N_1647,N_1459,N_1507);
or U1648 (N_1648,N_1473,N_1510);
xor U1649 (N_1649,N_1527,N_1549);
nand U1650 (N_1650,N_1569,N_1539);
or U1651 (N_1651,N_1550,N_1479);
or U1652 (N_1652,N_1482,N_1543);
or U1653 (N_1653,N_1467,N_1414);
nand U1654 (N_1654,N_1453,N_1593);
and U1655 (N_1655,N_1565,N_1444);
and U1656 (N_1656,N_1475,N_1505);
nand U1657 (N_1657,N_1437,N_1441);
or U1658 (N_1658,N_1520,N_1528);
or U1659 (N_1659,N_1556,N_1552);
nor U1660 (N_1660,N_1484,N_1580);
or U1661 (N_1661,N_1411,N_1581);
nand U1662 (N_1662,N_1572,N_1471);
xor U1663 (N_1663,N_1425,N_1566);
nand U1664 (N_1664,N_1416,N_1519);
or U1665 (N_1665,N_1452,N_1468);
nand U1666 (N_1666,N_1420,N_1427);
nand U1667 (N_1667,N_1522,N_1470);
xnor U1668 (N_1668,N_1442,N_1571);
and U1669 (N_1669,N_1474,N_1438);
and U1670 (N_1670,N_1493,N_1492);
or U1671 (N_1671,N_1423,N_1486);
nor U1672 (N_1672,N_1480,N_1477);
nor U1673 (N_1673,N_1599,N_1424);
nand U1674 (N_1674,N_1487,N_1558);
or U1675 (N_1675,N_1404,N_1530);
or U1676 (N_1676,N_1546,N_1508);
nor U1677 (N_1677,N_1582,N_1567);
and U1678 (N_1678,N_1513,N_1413);
and U1679 (N_1679,N_1542,N_1551);
and U1680 (N_1680,N_1440,N_1521);
nor U1681 (N_1681,N_1506,N_1577);
nand U1682 (N_1682,N_1515,N_1435);
nand U1683 (N_1683,N_1418,N_1524);
xnor U1684 (N_1684,N_1430,N_1541);
xnor U1685 (N_1685,N_1476,N_1488);
nor U1686 (N_1686,N_1544,N_1472);
nand U1687 (N_1687,N_1494,N_1463);
nand U1688 (N_1688,N_1448,N_1583);
and U1689 (N_1689,N_1511,N_1462);
nor U1690 (N_1690,N_1514,N_1560);
nor U1691 (N_1691,N_1439,N_1457);
nor U1692 (N_1692,N_1596,N_1496);
and U1693 (N_1693,N_1501,N_1464);
or U1694 (N_1694,N_1454,N_1456);
nor U1695 (N_1695,N_1595,N_1421);
nor U1696 (N_1696,N_1405,N_1574);
nor U1697 (N_1697,N_1458,N_1408);
and U1698 (N_1698,N_1469,N_1584);
or U1699 (N_1699,N_1403,N_1516);
nor U1700 (N_1700,N_1557,N_1488);
nand U1701 (N_1701,N_1484,N_1589);
xnor U1702 (N_1702,N_1549,N_1472);
nand U1703 (N_1703,N_1482,N_1485);
xnor U1704 (N_1704,N_1544,N_1461);
nand U1705 (N_1705,N_1436,N_1538);
nor U1706 (N_1706,N_1468,N_1557);
nand U1707 (N_1707,N_1525,N_1567);
and U1708 (N_1708,N_1427,N_1443);
and U1709 (N_1709,N_1439,N_1407);
xor U1710 (N_1710,N_1437,N_1491);
or U1711 (N_1711,N_1473,N_1403);
or U1712 (N_1712,N_1516,N_1598);
nand U1713 (N_1713,N_1470,N_1558);
and U1714 (N_1714,N_1591,N_1484);
nor U1715 (N_1715,N_1451,N_1579);
nor U1716 (N_1716,N_1461,N_1585);
nand U1717 (N_1717,N_1485,N_1498);
nand U1718 (N_1718,N_1448,N_1536);
and U1719 (N_1719,N_1498,N_1479);
or U1720 (N_1720,N_1556,N_1438);
and U1721 (N_1721,N_1466,N_1507);
and U1722 (N_1722,N_1564,N_1467);
nor U1723 (N_1723,N_1503,N_1477);
and U1724 (N_1724,N_1504,N_1425);
or U1725 (N_1725,N_1525,N_1523);
and U1726 (N_1726,N_1547,N_1444);
and U1727 (N_1727,N_1419,N_1565);
nor U1728 (N_1728,N_1417,N_1558);
nand U1729 (N_1729,N_1543,N_1545);
or U1730 (N_1730,N_1437,N_1593);
nor U1731 (N_1731,N_1470,N_1523);
nor U1732 (N_1732,N_1441,N_1549);
nor U1733 (N_1733,N_1408,N_1569);
or U1734 (N_1734,N_1551,N_1590);
nor U1735 (N_1735,N_1580,N_1494);
and U1736 (N_1736,N_1496,N_1493);
xor U1737 (N_1737,N_1562,N_1512);
nand U1738 (N_1738,N_1599,N_1434);
nand U1739 (N_1739,N_1526,N_1523);
nand U1740 (N_1740,N_1521,N_1412);
or U1741 (N_1741,N_1581,N_1503);
nor U1742 (N_1742,N_1565,N_1526);
nand U1743 (N_1743,N_1491,N_1480);
nor U1744 (N_1744,N_1430,N_1578);
nand U1745 (N_1745,N_1565,N_1557);
or U1746 (N_1746,N_1512,N_1407);
nor U1747 (N_1747,N_1514,N_1546);
nand U1748 (N_1748,N_1483,N_1428);
nand U1749 (N_1749,N_1401,N_1461);
nand U1750 (N_1750,N_1476,N_1507);
nand U1751 (N_1751,N_1524,N_1538);
nor U1752 (N_1752,N_1439,N_1429);
nor U1753 (N_1753,N_1500,N_1504);
and U1754 (N_1754,N_1532,N_1581);
nor U1755 (N_1755,N_1436,N_1420);
or U1756 (N_1756,N_1525,N_1532);
and U1757 (N_1757,N_1528,N_1440);
nor U1758 (N_1758,N_1592,N_1444);
and U1759 (N_1759,N_1466,N_1592);
or U1760 (N_1760,N_1494,N_1552);
or U1761 (N_1761,N_1509,N_1483);
and U1762 (N_1762,N_1438,N_1504);
or U1763 (N_1763,N_1551,N_1530);
and U1764 (N_1764,N_1464,N_1566);
nand U1765 (N_1765,N_1402,N_1544);
nand U1766 (N_1766,N_1535,N_1530);
and U1767 (N_1767,N_1426,N_1556);
nand U1768 (N_1768,N_1570,N_1423);
nand U1769 (N_1769,N_1579,N_1429);
and U1770 (N_1770,N_1412,N_1573);
or U1771 (N_1771,N_1551,N_1428);
nand U1772 (N_1772,N_1423,N_1415);
and U1773 (N_1773,N_1404,N_1422);
nand U1774 (N_1774,N_1468,N_1510);
and U1775 (N_1775,N_1543,N_1473);
nor U1776 (N_1776,N_1492,N_1517);
nand U1777 (N_1777,N_1515,N_1426);
nand U1778 (N_1778,N_1424,N_1561);
nand U1779 (N_1779,N_1496,N_1400);
and U1780 (N_1780,N_1475,N_1459);
or U1781 (N_1781,N_1579,N_1493);
nand U1782 (N_1782,N_1412,N_1506);
nor U1783 (N_1783,N_1528,N_1536);
and U1784 (N_1784,N_1465,N_1499);
nor U1785 (N_1785,N_1534,N_1450);
and U1786 (N_1786,N_1422,N_1587);
nand U1787 (N_1787,N_1401,N_1596);
xnor U1788 (N_1788,N_1599,N_1588);
nand U1789 (N_1789,N_1465,N_1431);
nand U1790 (N_1790,N_1451,N_1441);
or U1791 (N_1791,N_1581,N_1401);
or U1792 (N_1792,N_1433,N_1476);
nor U1793 (N_1793,N_1503,N_1550);
or U1794 (N_1794,N_1426,N_1552);
nand U1795 (N_1795,N_1587,N_1446);
nor U1796 (N_1796,N_1447,N_1561);
and U1797 (N_1797,N_1570,N_1507);
or U1798 (N_1798,N_1456,N_1593);
and U1799 (N_1799,N_1414,N_1543);
or U1800 (N_1800,N_1663,N_1703);
or U1801 (N_1801,N_1651,N_1622);
and U1802 (N_1802,N_1682,N_1673);
and U1803 (N_1803,N_1629,N_1716);
nor U1804 (N_1804,N_1798,N_1738);
or U1805 (N_1805,N_1636,N_1777);
or U1806 (N_1806,N_1652,N_1617);
or U1807 (N_1807,N_1700,N_1718);
and U1808 (N_1808,N_1721,N_1740);
nor U1809 (N_1809,N_1720,N_1706);
or U1810 (N_1810,N_1657,N_1632);
nor U1811 (N_1811,N_1790,N_1649);
nor U1812 (N_1812,N_1601,N_1633);
nand U1813 (N_1813,N_1638,N_1748);
or U1814 (N_1814,N_1793,N_1780);
nor U1815 (N_1815,N_1630,N_1726);
or U1816 (N_1816,N_1665,N_1676);
and U1817 (N_1817,N_1711,N_1705);
nor U1818 (N_1818,N_1723,N_1759);
or U1819 (N_1819,N_1786,N_1778);
nor U1820 (N_1820,N_1626,N_1749);
or U1821 (N_1821,N_1776,N_1719);
or U1822 (N_1822,N_1739,N_1717);
or U1823 (N_1823,N_1753,N_1693);
and U1824 (N_1824,N_1675,N_1770);
nor U1825 (N_1825,N_1733,N_1764);
and U1826 (N_1826,N_1757,N_1635);
or U1827 (N_1827,N_1795,N_1752);
nand U1828 (N_1828,N_1624,N_1732);
or U1829 (N_1829,N_1754,N_1600);
nor U1830 (N_1830,N_1713,N_1653);
nand U1831 (N_1831,N_1767,N_1607);
nor U1832 (N_1832,N_1688,N_1796);
nor U1833 (N_1833,N_1680,N_1619);
or U1834 (N_1834,N_1707,N_1667);
or U1835 (N_1835,N_1729,N_1620);
and U1836 (N_1836,N_1645,N_1775);
nand U1837 (N_1837,N_1612,N_1603);
nand U1838 (N_1838,N_1695,N_1664);
nand U1839 (N_1839,N_1779,N_1631);
nand U1840 (N_1840,N_1763,N_1677);
nand U1841 (N_1841,N_1737,N_1760);
nand U1842 (N_1842,N_1662,N_1605);
nor U1843 (N_1843,N_1730,N_1614);
nor U1844 (N_1844,N_1709,N_1687);
or U1845 (N_1845,N_1609,N_1715);
nand U1846 (N_1846,N_1608,N_1735);
nand U1847 (N_1847,N_1728,N_1613);
nand U1848 (N_1848,N_1616,N_1679);
and U1849 (N_1849,N_1771,N_1746);
nand U1850 (N_1850,N_1642,N_1644);
nor U1851 (N_1851,N_1625,N_1692);
xnor U1852 (N_1852,N_1772,N_1654);
or U1853 (N_1853,N_1646,N_1712);
nand U1854 (N_1854,N_1743,N_1751);
nand U1855 (N_1855,N_1736,N_1727);
or U1856 (N_1856,N_1648,N_1656);
or U1857 (N_1857,N_1742,N_1769);
nand U1858 (N_1858,N_1714,N_1750);
and U1859 (N_1859,N_1792,N_1690);
or U1860 (N_1860,N_1797,N_1666);
and U1861 (N_1861,N_1781,N_1758);
xnor U1862 (N_1862,N_1799,N_1783);
nor U1863 (N_1863,N_1710,N_1615);
xor U1864 (N_1864,N_1683,N_1761);
nand U1865 (N_1865,N_1747,N_1672);
and U1866 (N_1866,N_1789,N_1756);
nor U1867 (N_1867,N_1697,N_1725);
and U1868 (N_1868,N_1650,N_1643);
or U1869 (N_1869,N_1686,N_1610);
and U1870 (N_1870,N_1765,N_1744);
and U1871 (N_1871,N_1647,N_1791);
and U1872 (N_1872,N_1634,N_1702);
and U1873 (N_1873,N_1691,N_1671);
nand U1874 (N_1874,N_1661,N_1621);
or U1875 (N_1875,N_1658,N_1704);
nand U1876 (N_1876,N_1611,N_1731);
or U1877 (N_1877,N_1659,N_1787);
and U1878 (N_1878,N_1755,N_1724);
and U1879 (N_1879,N_1768,N_1681);
or U1880 (N_1880,N_1766,N_1762);
or U1881 (N_1881,N_1606,N_1641);
nand U1882 (N_1882,N_1685,N_1698);
nor U1883 (N_1883,N_1669,N_1640);
xnor U1884 (N_1884,N_1655,N_1628);
and U1885 (N_1885,N_1689,N_1623);
or U1886 (N_1886,N_1782,N_1794);
nand U1887 (N_1887,N_1684,N_1699);
nand U1888 (N_1888,N_1602,N_1722);
nor U1889 (N_1889,N_1734,N_1660);
nand U1890 (N_1890,N_1639,N_1788);
nor U1891 (N_1891,N_1784,N_1694);
and U1892 (N_1892,N_1678,N_1618);
nor U1893 (N_1893,N_1674,N_1668);
nand U1894 (N_1894,N_1627,N_1745);
nand U1895 (N_1895,N_1773,N_1708);
or U1896 (N_1896,N_1696,N_1785);
nor U1897 (N_1897,N_1604,N_1774);
and U1898 (N_1898,N_1741,N_1701);
nand U1899 (N_1899,N_1670,N_1637);
and U1900 (N_1900,N_1732,N_1706);
and U1901 (N_1901,N_1686,N_1620);
nand U1902 (N_1902,N_1600,N_1636);
or U1903 (N_1903,N_1662,N_1668);
or U1904 (N_1904,N_1781,N_1632);
or U1905 (N_1905,N_1795,N_1769);
nor U1906 (N_1906,N_1776,N_1746);
nor U1907 (N_1907,N_1667,N_1661);
and U1908 (N_1908,N_1695,N_1755);
or U1909 (N_1909,N_1662,N_1628);
and U1910 (N_1910,N_1638,N_1679);
and U1911 (N_1911,N_1672,N_1768);
nor U1912 (N_1912,N_1668,N_1655);
nor U1913 (N_1913,N_1772,N_1639);
and U1914 (N_1914,N_1786,N_1678);
and U1915 (N_1915,N_1700,N_1691);
nor U1916 (N_1916,N_1776,N_1615);
or U1917 (N_1917,N_1687,N_1618);
nor U1918 (N_1918,N_1675,N_1793);
and U1919 (N_1919,N_1773,N_1771);
nand U1920 (N_1920,N_1675,N_1637);
and U1921 (N_1921,N_1639,N_1728);
or U1922 (N_1922,N_1741,N_1618);
and U1923 (N_1923,N_1659,N_1715);
and U1924 (N_1924,N_1715,N_1696);
or U1925 (N_1925,N_1608,N_1603);
and U1926 (N_1926,N_1643,N_1670);
or U1927 (N_1927,N_1648,N_1790);
nor U1928 (N_1928,N_1788,N_1756);
or U1929 (N_1929,N_1692,N_1723);
xnor U1930 (N_1930,N_1717,N_1769);
nor U1931 (N_1931,N_1661,N_1630);
nand U1932 (N_1932,N_1607,N_1779);
nor U1933 (N_1933,N_1623,N_1625);
and U1934 (N_1934,N_1752,N_1742);
nor U1935 (N_1935,N_1691,N_1709);
nand U1936 (N_1936,N_1758,N_1625);
or U1937 (N_1937,N_1614,N_1792);
nor U1938 (N_1938,N_1663,N_1608);
nand U1939 (N_1939,N_1662,N_1646);
and U1940 (N_1940,N_1661,N_1703);
and U1941 (N_1941,N_1679,N_1646);
and U1942 (N_1942,N_1694,N_1755);
nor U1943 (N_1943,N_1648,N_1760);
and U1944 (N_1944,N_1735,N_1653);
nor U1945 (N_1945,N_1727,N_1678);
nor U1946 (N_1946,N_1721,N_1655);
or U1947 (N_1947,N_1746,N_1715);
xor U1948 (N_1948,N_1690,N_1681);
nand U1949 (N_1949,N_1626,N_1625);
or U1950 (N_1950,N_1700,N_1768);
nor U1951 (N_1951,N_1618,N_1694);
or U1952 (N_1952,N_1685,N_1600);
and U1953 (N_1953,N_1778,N_1606);
nor U1954 (N_1954,N_1796,N_1712);
and U1955 (N_1955,N_1611,N_1692);
nor U1956 (N_1956,N_1710,N_1700);
nand U1957 (N_1957,N_1756,N_1664);
or U1958 (N_1958,N_1604,N_1717);
nand U1959 (N_1959,N_1678,N_1698);
or U1960 (N_1960,N_1619,N_1750);
or U1961 (N_1961,N_1735,N_1696);
and U1962 (N_1962,N_1792,N_1738);
or U1963 (N_1963,N_1639,N_1670);
or U1964 (N_1964,N_1790,N_1679);
or U1965 (N_1965,N_1698,N_1621);
and U1966 (N_1966,N_1729,N_1771);
nand U1967 (N_1967,N_1777,N_1637);
nand U1968 (N_1968,N_1685,N_1634);
nor U1969 (N_1969,N_1781,N_1612);
xor U1970 (N_1970,N_1723,N_1704);
nor U1971 (N_1971,N_1643,N_1755);
and U1972 (N_1972,N_1730,N_1755);
nand U1973 (N_1973,N_1752,N_1623);
nand U1974 (N_1974,N_1629,N_1741);
and U1975 (N_1975,N_1623,N_1673);
or U1976 (N_1976,N_1791,N_1658);
or U1977 (N_1977,N_1695,N_1734);
or U1978 (N_1978,N_1722,N_1701);
nor U1979 (N_1979,N_1687,N_1762);
and U1980 (N_1980,N_1665,N_1641);
and U1981 (N_1981,N_1663,N_1792);
nand U1982 (N_1982,N_1787,N_1673);
nor U1983 (N_1983,N_1675,N_1657);
nor U1984 (N_1984,N_1666,N_1710);
nand U1985 (N_1985,N_1686,N_1661);
and U1986 (N_1986,N_1769,N_1775);
xor U1987 (N_1987,N_1600,N_1703);
and U1988 (N_1988,N_1736,N_1752);
nand U1989 (N_1989,N_1629,N_1718);
nand U1990 (N_1990,N_1690,N_1660);
nor U1991 (N_1991,N_1701,N_1735);
xnor U1992 (N_1992,N_1626,N_1712);
nor U1993 (N_1993,N_1692,N_1786);
and U1994 (N_1994,N_1765,N_1691);
and U1995 (N_1995,N_1775,N_1649);
and U1996 (N_1996,N_1643,N_1714);
or U1997 (N_1997,N_1690,N_1655);
or U1998 (N_1998,N_1669,N_1723);
xor U1999 (N_1999,N_1781,N_1715);
and U2000 (N_2000,N_1949,N_1924);
nand U2001 (N_2001,N_1913,N_1872);
or U2002 (N_2002,N_1864,N_1806);
or U2003 (N_2003,N_1940,N_1954);
nor U2004 (N_2004,N_1888,N_1901);
or U2005 (N_2005,N_1845,N_1813);
nand U2006 (N_2006,N_1848,N_1932);
or U2007 (N_2007,N_1836,N_1952);
nand U2008 (N_2008,N_1817,N_1909);
or U2009 (N_2009,N_1801,N_1958);
nor U2010 (N_2010,N_1802,N_1902);
nor U2011 (N_2011,N_1889,N_1972);
or U2012 (N_2012,N_1847,N_1970);
or U2013 (N_2013,N_1857,N_1910);
nand U2014 (N_2014,N_1965,N_1811);
or U2015 (N_2015,N_1804,N_1803);
and U2016 (N_2016,N_1807,N_1846);
and U2017 (N_2017,N_1808,N_1834);
nor U2018 (N_2018,N_1851,N_1859);
nor U2019 (N_2019,N_1985,N_1829);
nor U2020 (N_2020,N_1870,N_1850);
nand U2021 (N_2021,N_1860,N_1818);
nand U2022 (N_2022,N_1887,N_1998);
nand U2023 (N_2023,N_1964,N_1988);
or U2024 (N_2024,N_1911,N_1968);
nor U2025 (N_2025,N_1946,N_1884);
and U2026 (N_2026,N_1874,N_1925);
and U2027 (N_2027,N_1892,N_1896);
and U2028 (N_2028,N_1861,N_1900);
and U2029 (N_2029,N_1994,N_1904);
nor U2030 (N_2030,N_1977,N_1867);
nand U2031 (N_2031,N_1979,N_1879);
nor U2032 (N_2032,N_1993,N_1875);
nand U2033 (N_2033,N_1984,N_1894);
nand U2034 (N_2034,N_1844,N_1947);
or U2035 (N_2035,N_1939,N_1955);
nor U2036 (N_2036,N_1843,N_1908);
and U2037 (N_2037,N_1918,N_1961);
and U2038 (N_2038,N_1854,N_1996);
nor U2039 (N_2039,N_1926,N_1963);
and U2040 (N_2040,N_1839,N_1987);
nand U2041 (N_2041,N_1820,N_1999);
or U2042 (N_2042,N_1960,N_1944);
nand U2043 (N_2043,N_1828,N_1880);
nand U2044 (N_2044,N_1907,N_1842);
and U2045 (N_2045,N_1816,N_1812);
xnor U2046 (N_2046,N_1862,N_1876);
nand U2047 (N_2047,N_1890,N_1830);
and U2048 (N_2048,N_1922,N_1832);
and U2049 (N_2049,N_1883,N_1882);
or U2050 (N_2050,N_1903,N_1840);
nand U2051 (N_2051,N_1981,N_1953);
nand U2052 (N_2052,N_1814,N_1871);
and U2053 (N_2053,N_1923,N_1899);
and U2054 (N_2054,N_1935,N_1916);
nor U2055 (N_2055,N_1863,N_1868);
or U2056 (N_2056,N_1831,N_1917);
and U2057 (N_2057,N_1928,N_1805);
or U2058 (N_2058,N_1800,N_1856);
nor U2059 (N_2059,N_1967,N_1822);
or U2060 (N_2060,N_1942,N_1927);
or U2061 (N_2061,N_1980,N_1838);
nand U2062 (N_2062,N_1933,N_1891);
nor U2063 (N_2063,N_1826,N_1930);
and U2064 (N_2064,N_1991,N_1983);
nor U2065 (N_2065,N_1959,N_1938);
nor U2066 (N_2066,N_1943,N_1974);
nand U2067 (N_2067,N_1934,N_1971);
nor U2068 (N_2068,N_1941,N_1835);
or U2069 (N_2069,N_1827,N_1936);
and U2070 (N_2070,N_1920,N_1852);
and U2071 (N_2071,N_1858,N_1873);
and U2072 (N_2072,N_1929,N_1921);
and U2073 (N_2073,N_1962,N_1897);
and U2074 (N_2074,N_1914,N_1948);
nor U2075 (N_2075,N_1966,N_1824);
nand U2076 (N_2076,N_1995,N_1809);
nor U2077 (N_2077,N_1869,N_1997);
and U2078 (N_2078,N_1877,N_1912);
nor U2079 (N_2079,N_1893,N_1975);
and U2080 (N_2080,N_1849,N_1821);
and U2081 (N_2081,N_1986,N_1878);
nand U2082 (N_2082,N_1819,N_1950);
or U2083 (N_2083,N_1906,N_1837);
and U2084 (N_2084,N_1989,N_1973);
nor U2085 (N_2085,N_1992,N_1956);
or U2086 (N_2086,N_1898,N_1931);
or U2087 (N_2087,N_1810,N_1915);
and U2088 (N_2088,N_1865,N_1969);
nor U2089 (N_2089,N_1945,N_1825);
nor U2090 (N_2090,N_1881,N_1853);
and U2091 (N_2091,N_1841,N_1823);
nor U2092 (N_2092,N_1951,N_1833);
nand U2093 (N_2093,N_1990,N_1982);
nor U2094 (N_2094,N_1886,N_1919);
and U2095 (N_2095,N_1937,N_1895);
or U2096 (N_2096,N_1978,N_1866);
or U2097 (N_2097,N_1957,N_1855);
or U2098 (N_2098,N_1885,N_1976);
and U2099 (N_2099,N_1815,N_1905);
nor U2100 (N_2100,N_1820,N_1876);
nor U2101 (N_2101,N_1879,N_1912);
nor U2102 (N_2102,N_1836,N_1825);
nor U2103 (N_2103,N_1844,N_1942);
xnor U2104 (N_2104,N_1862,N_1929);
and U2105 (N_2105,N_1888,N_1988);
or U2106 (N_2106,N_1994,N_1909);
nor U2107 (N_2107,N_1802,N_1969);
and U2108 (N_2108,N_1946,N_1945);
and U2109 (N_2109,N_1878,N_1875);
nor U2110 (N_2110,N_1990,N_1847);
and U2111 (N_2111,N_1842,N_1921);
and U2112 (N_2112,N_1820,N_1823);
nor U2113 (N_2113,N_1875,N_1819);
nor U2114 (N_2114,N_1936,N_1985);
nand U2115 (N_2115,N_1896,N_1997);
nand U2116 (N_2116,N_1958,N_1900);
nor U2117 (N_2117,N_1909,N_1805);
and U2118 (N_2118,N_1826,N_1912);
xor U2119 (N_2119,N_1911,N_1863);
or U2120 (N_2120,N_1877,N_1861);
nor U2121 (N_2121,N_1859,N_1852);
xnor U2122 (N_2122,N_1885,N_1922);
nor U2123 (N_2123,N_1940,N_1960);
or U2124 (N_2124,N_1865,N_1857);
and U2125 (N_2125,N_1928,N_1800);
or U2126 (N_2126,N_1941,N_1982);
and U2127 (N_2127,N_1985,N_1819);
or U2128 (N_2128,N_1966,N_1847);
nand U2129 (N_2129,N_1801,N_1913);
and U2130 (N_2130,N_1899,N_1838);
or U2131 (N_2131,N_1837,N_1840);
nand U2132 (N_2132,N_1897,N_1824);
nor U2133 (N_2133,N_1960,N_1947);
nand U2134 (N_2134,N_1823,N_1933);
xnor U2135 (N_2135,N_1895,N_1804);
and U2136 (N_2136,N_1878,N_1848);
nor U2137 (N_2137,N_1807,N_1903);
nand U2138 (N_2138,N_1934,N_1813);
nand U2139 (N_2139,N_1887,N_1828);
and U2140 (N_2140,N_1942,N_1866);
nor U2141 (N_2141,N_1854,N_1936);
and U2142 (N_2142,N_1900,N_1989);
nand U2143 (N_2143,N_1982,N_1948);
nand U2144 (N_2144,N_1803,N_1968);
or U2145 (N_2145,N_1988,N_1973);
nor U2146 (N_2146,N_1947,N_1885);
or U2147 (N_2147,N_1958,N_1956);
and U2148 (N_2148,N_1851,N_1825);
or U2149 (N_2149,N_1899,N_1895);
or U2150 (N_2150,N_1882,N_1948);
nand U2151 (N_2151,N_1870,N_1978);
and U2152 (N_2152,N_1993,N_1961);
or U2153 (N_2153,N_1919,N_1995);
or U2154 (N_2154,N_1893,N_1995);
nand U2155 (N_2155,N_1894,N_1928);
or U2156 (N_2156,N_1982,N_1865);
nand U2157 (N_2157,N_1935,N_1951);
and U2158 (N_2158,N_1928,N_1963);
nor U2159 (N_2159,N_1817,N_1940);
or U2160 (N_2160,N_1839,N_1895);
nand U2161 (N_2161,N_1972,N_1853);
nand U2162 (N_2162,N_1990,N_1914);
nor U2163 (N_2163,N_1858,N_1835);
or U2164 (N_2164,N_1985,N_1951);
nor U2165 (N_2165,N_1842,N_1826);
or U2166 (N_2166,N_1862,N_1987);
and U2167 (N_2167,N_1933,N_1954);
nand U2168 (N_2168,N_1817,N_1887);
and U2169 (N_2169,N_1991,N_1970);
nand U2170 (N_2170,N_1953,N_1989);
and U2171 (N_2171,N_1958,N_1888);
nor U2172 (N_2172,N_1862,N_1893);
nand U2173 (N_2173,N_1934,N_1930);
nor U2174 (N_2174,N_1863,N_1924);
nand U2175 (N_2175,N_1926,N_1902);
nor U2176 (N_2176,N_1805,N_1826);
nand U2177 (N_2177,N_1848,N_1883);
nor U2178 (N_2178,N_1892,N_1822);
nand U2179 (N_2179,N_1807,N_1933);
nand U2180 (N_2180,N_1835,N_1947);
nand U2181 (N_2181,N_1876,N_1924);
nand U2182 (N_2182,N_1980,N_1817);
and U2183 (N_2183,N_1913,N_1935);
nand U2184 (N_2184,N_1971,N_1833);
nand U2185 (N_2185,N_1813,N_1927);
or U2186 (N_2186,N_1863,N_1920);
and U2187 (N_2187,N_1976,N_1946);
or U2188 (N_2188,N_1987,N_1935);
nand U2189 (N_2189,N_1857,N_1851);
nand U2190 (N_2190,N_1957,N_1821);
or U2191 (N_2191,N_1979,N_1871);
nand U2192 (N_2192,N_1870,N_1845);
nor U2193 (N_2193,N_1830,N_1925);
nand U2194 (N_2194,N_1893,N_1998);
and U2195 (N_2195,N_1907,N_1835);
or U2196 (N_2196,N_1819,N_1804);
xor U2197 (N_2197,N_1870,N_1982);
nor U2198 (N_2198,N_1992,N_1879);
nand U2199 (N_2199,N_1894,N_1946);
and U2200 (N_2200,N_2012,N_2194);
nor U2201 (N_2201,N_2029,N_2026);
nor U2202 (N_2202,N_2059,N_2170);
or U2203 (N_2203,N_2030,N_2176);
nand U2204 (N_2204,N_2169,N_2095);
nor U2205 (N_2205,N_2108,N_2145);
nor U2206 (N_2206,N_2002,N_2163);
and U2207 (N_2207,N_2111,N_2172);
nor U2208 (N_2208,N_2186,N_2189);
or U2209 (N_2209,N_2136,N_2043);
nand U2210 (N_2210,N_2123,N_2144);
or U2211 (N_2211,N_2178,N_2017);
xor U2212 (N_2212,N_2061,N_2128);
and U2213 (N_2213,N_2103,N_2031);
and U2214 (N_2214,N_2087,N_2159);
nor U2215 (N_2215,N_2143,N_2101);
and U2216 (N_2216,N_2166,N_2062);
or U2217 (N_2217,N_2140,N_2092);
nand U2218 (N_2218,N_2068,N_2179);
or U2219 (N_2219,N_2130,N_2047);
nand U2220 (N_2220,N_2120,N_2134);
and U2221 (N_2221,N_2078,N_2125);
nand U2222 (N_2222,N_2102,N_2053);
nand U2223 (N_2223,N_2018,N_2073);
and U2224 (N_2224,N_2162,N_2011);
or U2225 (N_2225,N_2024,N_2141);
or U2226 (N_2226,N_2138,N_2192);
nor U2227 (N_2227,N_2185,N_2109);
or U2228 (N_2228,N_2076,N_2075);
nor U2229 (N_2229,N_2124,N_2121);
nand U2230 (N_2230,N_2044,N_2175);
nor U2231 (N_2231,N_2028,N_2195);
nor U2232 (N_2232,N_2049,N_2187);
and U2233 (N_2233,N_2142,N_2063);
or U2234 (N_2234,N_2173,N_2065);
or U2235 (N_2235,N_2016,N_2045);
nor U2236 (N_2236,N_2070,N_2132);
nor U2237 (N_2237,N_2036,N_2131);
or U2238 (N_2238,N_2093,N_2054);
or U2239 (N_2239,N_2160,N_2048);
or U2240 (N_2240,N_2154,N_2098);
nand U2241 (N_2241,N_2196,N_2020);
nor U2242 (N_2242,N_2193,N_2199);
or U2243 (N_2243,N_2088,N_2085);
nand U2244 (N_2244,N_2114,N_2009);
nor U2245 (N_2245,N_2096,N_2082);
and U2246 (N_2246,N_2107,N_2083);
nor U2247 (N_2247,N_2023,N_2067);
and U2248 (N_2248,N_2071,N_2041);
or U2249 (N_2249,N_2034,N_2158);
nor U2250 (N_2250,N_2127,N_2090);
and U2251 (N_2251,N_2151,N_2003);
nor U2252 (N_2252,N_2021,N_2182);
and U2253 (N_2253,N_2072,N_2104);
and U2254 (N_2254,N_2097,N_2119);
nor U2255 (N_2255,N_2094,N_2190);
and U2256 (N_2256,N_2027,N_2035);
nor U2257 (N_2257,N_2010,N_2006);
and U2258 (N_2258,N_2046,N_2080);
nor U2259 (N_2259,N_2174,N_2013);
and U2260 (N_2260,N_2007,N_2115);
or U2261 (N_2261,N_2153,N_2064);
nand U2262 (N_2262,N_2042,N_2055);
or U2263 (N_2263,N_2008,N_2106);
nand U2264 (N_2264,N_2014,N_2148);
and U2265 (N_2265,N_2150,N_2032);
nor U2266 (N_2266,N_2079,N_2058);
xor U2267 (N_2267,N_2100,N_2060);
nor U2268 (N_2268,N_2081,N_2000);
and U2269 (N_2269,N_2117,N_2184);
or U2270 (N_2270,N_2105,N_2171);
and U2271 (N_2271,N_2180,N_2037);
xor U2272 (N_2272,N_2057,N_2167);
and U2273 (N_2273,N_2161,N_2001);
xnor U2274 (N_2274,N_2038,N_2015);
nor U2275 (N_2275,N_2146,N_2091);
nor U2276 (N_2276,N_2112,N_2116);
nand U2277 (N_2277,N_2156,N_2139);
or U2278 (N_2278,N_2147,N_2149);
nor U2279 (N_2279,N_2089,N_2033);
xnor U2280 (N_2280,N_2084,N_2052);
or U2281 (N_2281,N_2168,N_2039);
or U2282 (N_2282,N_2198,N_2164);
and U2283 (N_2283,N_2056,N_2152);
or U2284 (N_2284,N_2005,N_2188);
nor U2285 (N_2285,N_2004,N_2050);
or U2286 (N_2286,N_2137,N_2157);
or U2287 (N_2287,N_2177,N_2129);
nand U2288 (N_2288,N_2019,N_2066);
nor U2289 (N_2289,N_2133,N_2181);
nand U2290 (N_2290,N_2022,N_2099);
and U2291 (N_2291,N_2118,N_2122);
and U2292 (N_2292,N_2051,N_2040);
nor U2293 (N_2293,N_2155,N_2086);
and U2294 (N_2294,N_2165,N_2025);
nand U2295 (N_2295,N_2077,N_2183);
nor U2296 (N_2296,N_2135,N_2069);
nor U2297 (N_2297,N_2126,N_2191);
or U2298 (N_2298,N_2074,N_2197);
and U2299 (N_2299,N_2113,N_2110);
nor U2300 (N_2300,N_2042,N_2117);
or U2301 (N_2301,N_2071,N_2007);
nor U2302 (N_2302,N_2183,N_2193);
xnor U2303 (N_2303,N_2169,N_2110);
or U2304 (N_2304,N_2045,N_2059);
or U2305 (N_2305,N_2091,N_2019);
and U2306 (N_2306,N_2012,N_2088);
and U2307 (N_2307,N_2106,N_2125);
or U2308 (N_2308,N_2182,N_2091);
and U2309 (N_2309,N_2007,N_2059);
nor U2310 (N_2310,N_2168,N_2097);
or U2311 (N_2311,N_2074,N_2193);
and U2312 (N_2312,N_2123,N_2004);
and U2313 (N_2313,N_2140,N_2143);
and U2314 (N_2314,N_2004,N_2194);
nand U2315 (N_2315,N_2081,N_2124);
and U2316 (N_2316,N_2104,N_2194);
nor U2317 (N_2317,N_2076,N_2061);
or U2318 (N_2318,N_2016,N_2005);
nor U2319 (N_2319,N_2007,N_2095);
or U2320 (N_2320,N_2088,N_2187);
xnor U2321 (N_2321,N_2059,N_2024);
nor U2322 (N_2322,N_2081,N_2026);
nand U2323 (N_2323,N_2168,N_2100);
nor U2324 (N_2324,N_2194,N_2082);
nor U2325 (N_2325,N_2183,N_2088);
and U2326 (N_2326,N_2086,N_2140);
and U2327 (N_2327,N_2031,N_2093);
nor U2328 (N_2328,N_2012,N_2164);
nor U2329 (N_2329,N_2153,N_2118);
nor U2330 (N_2330,N_2108,N_2133);
and U2331 (N_2331,N_2192,N_2143);
or U2332 (N_2332,N_2197,N_2100);
nor U2333 (N_2333,N_2191,N_2094);
or U2334 (N_2334,N_2123,N_2030);
nand U2335 (N_2335,N_2050,N_2195);
nor U2336 (N_2336,N_2180,N_2029);
nor U2337 (N_2337,N_2170,N_2195);
or U2338 (N_2338,N_2047,N_2141);
and U2339 (N_2339,N_2133,N_2175);
nand U2340 (N_2340,N_2005,N_2026);
nor U2341 (N_2341,N_2038,N_2058);
nor U2342 (N_2342,N_2191,N_2136);
nor U2343 (N_2343,N_2169,N_2023);
nand U2344 (N_2344,N_2137,N_2198);
or U2345 (N_2345,N_2002,N_2145);
nand U2346 (N_2346,N_2043,N_2104);
nor U2347 (N_2347,N_2136,N_2033);
and U2348 (N_2348,N_2064,N_2172);
and U2349 (N_2349,N_2040,N_2104);
nand U2350 (N_2350,N_2054,N_2165);
nor U2351 (N_2351,N_2146,N_2081);
nor U2352 (N_2352,N_2111,N_2133);
and U2353 (N_2353,N_2076,N_2040);
and U2354 (N_2354,N_2186,N_2085);
nand U2355 (N_2355,N_2100,N_2166);
nand U2356 (N_2356,N_2020,N_2021);
or U2357 (N_2357,N_2095,N_2012);
or U2358 (N_2358,N_2011,N_2061);
nand U2359 (N_2359,N_2156,N_2035);
nand U2360 (N_2360,N_2186,N_2134);
nand U2361 (N_2361,N_2179,N_2150);
nor U2362 (N_2362,N_2141,N_2181);
nor U2363 (N_2363,N_2075,N_2119);
nand U2364 (N_2364,N_2151,N_2078);
nand U2365 (N_2365,N_2140,N_2010);
and U2366 (N_2366,N_2126,N_2145);
nor U2367 (N_2367,N_2154,N_2177);
and U2368 (N_2368,N_2178,N_2052);
nor U2369 (N_2369,N_2030,N_2024);
and U2370 (N_2370,N_2078,N_2060);
nand U2371 (N_2371,N_2069,N_2117);
or U2372 (N_2372,N_2080,N_2029);
nand U2373 (N_2373,N_2178,N_2089);
nand U2374 (N_2374,N_2021,N_2084);
nor U2375 (N_2375,N_2127,N_2137);
or U2376 (N_2376,N_2194,N_2053);
nor U2377 (N_2377,N_2087,N_2103);
nor U2378 (N_2378,N_2039,N_2198);
and U2379 (N_2379,N_2164,N_2086);
or U2380 (N_2380,N_2117,N_2137);
or U2381 (N_2381,N_2182,N_2060);
and U2382 (N_2382,N_2189,N_2087);
or U2383 (N_2383,N_2104,N_2007);
or U2384 (N_2384,N_2172,N_2117);
and U2385 (N_2385,N_2079,N_2066);
xor U2386 (N_2386,N_2177,N_2070);
nor U2387 (N_2387,N_2174,N_2063);
nand U2388 (N_2388,N_2100,N_2000);
nor U2389 (N_2389,N_2167,N_2093);
nor U2390 (N_2390,N_2169,N_2164);
and U2391 (N_2391,N_2174,N_2113);
or U2392 (N_2392,N_2037,N_2071);
and U2393 (N_2393,N_2069,N_2004);
nand U2394 (N_2394,N_2142,N_2091);
and U2395 (N_2395,N_2180,N_2115);
and U2396 (N_2396,N_2090,N_2002);
nand U2397 (N_2397,N_2078,N_2118);
or U2398 (N_2398,N_2142,N_2155);
nor U2399 (N_2399,N_2065,N_2049);
nand U2400 (N_2400,N_2394,N_2370);
nand U2401 (N_2401,N_2218,N_2327);
nand U2402 (N_2402,N_2239,N_2315);
nand U2403 (N_2403,N_2229,N_2364);
nor U2404 (N_2404,N_2219,N_2206);
and U2405 (N_2405,N_2220,N_2326);
nor U2406 (N_2406,N_2396,N_2307);
or U2407 (N_2407,N_2210,N_2328);
and U2408 (N_2408,N_2202,N_2245);
and U2409 (N_2409,N_2284,N_2278);
nand U2410 (N_2410,N_2244,N_2368);
or U2411 (N_2411,N_2213,N_2249);
and U2412 (N_2412,N_2322,N_2217);
or U2413 (N_2413,N_2321,N_2253);
or U2414 (N_2414,N_2332,N_2340);
and U2415 (N_2415,N_2200,N_2357);
nand U2416 (N_2416,N_2299,N_2345);
nand U2417 (N_2417,N_2386,N_2352);
or U2418 (N_2418,N_2361,N_2211);
nor U2419 (N_2419,N_2235,N_2308);
nor U2420 (N_2420,N_2221,N_2367);
nand U2421 (N_2421,N_2362,N_2260);
nand U2422 (N_2422,N_2379,N_2282);
and U2423 (N_2423,N_2359,N_2264);
or U2424 (N_2424,N_2360,N_2223);
and U2425 (N_2425,N_2304,N_2266);
nand U2426 (N_2426,N_2277,N_2392);
and U2427 (N_2427,N_2205,N_2300);
nand U2428 (N_2428,N_2283,N_2250);
nand U2429 (N_2429,N_2395,N_2366);
and U2430 (N_2430,N_2258,N_2240);
nand U2431 (N_2431,N_2377,N_2285);
nand U2432 (N_2432,N_2255,N_2346);
nor U2433 (N_2433,N_2269,N_2354);
or U2434 (N_2434,N_2373,N_2267);
nor U2435 (N_2435,N_2236,N_2323);
and U2436 (N_2436,N_2274,N_2333);
and U2437 (N_2437,N_2331,N_2265);
or U2438 (N_2438,N_2318,N_2261);
or U2439 (N_2439,N_2275,N_2288);
and U2440 (N_2440,N_2224,N_2311);
xor U2441 (N_2441,N_2393,N_2349);
xnor U2442 (N_2442,N_2252,N_2385);
nand U2443 (N_2443,N_2247,N_2263);
nor U2444 (N_2444,N_2317,N_2324);
nand U2445 (N_2445,N_2243,N_2376);
or U2446 (N_2446,N_2378,N_2207);
xor U2447 (N_2447,N_2389,N_2380);
or U2448 (N_2448,N_2351,N_2397);
nand U2449 (N_2449,N_2209,N_2348);
or U2450 (N_2450,N_2291,N_2384);
nand U2451 (N_2451,N_2214,N_2399);
nand U2452 (N_2452,N_2334,N_2344);
and U2453 (N_2453,N_2390,N_2295);
nor U2454 (N_2454,N_2391,N_2309);
nor U2455 (N_2455,N_2251,N_2358);
xor U2456 (N_2456,N_2382,N_2271);
nor U2457 (N_2457,N_2330,N_2293);
and U2458 (N_2458,N_2272,N_2303);
nor U2459 (N_2459,N_2301,N_2302);
nand U2460 (N_2460,N_2254,N_2298);
nor U2461 (N_2461,N_2287,N_2337);
or U2462 (N_2462,N_2374,N_2336);
nand U2463 (N_2463,N_2237,N_2335);
nor U2464 (N_2464,N_2371,N_2297);
nor U2465 (N_2465,N_2227,N_2216);
and U2466 (N_2466,N_2215,N_2204);
nand U2467 (N_2467,N_2343,N_2341);
or U2468 (N_2468,N_2203,N_2398);
nand U2469 (N_2469,N_2347,N_2286);
nand U2470 (N_2470,N_2270,N_2276);
and U2471 (N_2471,N_2381,N_2290);
or U2472 (N_2472,N_2387,N_2289);
nand U2473 (N_2473,N_2262,N_2234);
nor U2474 (N_2474,N_2257,N_2350);
nand U2475 (N_2475,N_2292,N_2268);
or U2476 (N_2476,N_2230,N_2256);
and U2477 (N_2477,N_2242,N_2313);
and U2478 (N_2478,N_2355,N_2226);
nor U2479 (N_2479,N_2363,N_2356);
or U2480 (N_2480,N_2212,N_2233);
nor U2481 (N_2481,N_2273,N_2353);
nor U2482 (N_2482,N_2388,N_2201);
or U2483 (N_2483,N_2225,N_2316);
nand U2484 (N_2484,N_2342,N_2222);
nor U2485 (N_2485,N_2228,N_2314);
nor U2486 (N_2486,N_2365,N_2232);
and U2487 (N_2487,N_2383,N_2310);
or U2488 (N_2488,N_2329,N_2375);
nand U2489 (N_2489,N_2294,N_2241);
nor U2490 (N_2490,N_2312,N_2306);
nor U2491 (N_2491,N_2238,N_2319);
or U2492 (N_2492,N_2325,N_2231);
nor U2493 (N_2493,N_2296,N_2372);
nor U2494 (N_2494,N_2259,N_2339);
and U2495 (N_2495,N_2305,N_2280);
nor U2496 (N_2496,N_2338,N_2369);
and U2497 (N_2497,N_2281,N_2320);
nor U2498 (N_2498,N_2208,N_2248);
nand U2499 (N_2499,N_2246,N_2279);
nor U2500 (N_2500,N_2354,N_2380);
nor U2501 (N_2501,N_2387,N_2364);
nand U2502 (N_2502,N_2209,N_2234);
or U2503 (N_2503,N_2317,N_2259);
nor U2504 (N_2504,N_2331,N_2221);
nand U2505 (N_2505,N_2389,N_2368);
nand U2506 (N_2506,N_2233,N_2308);
nor U2507 (N_2507,N_2305,N_2246);
or U2508 (N_2508,N_2304,N_2289);
and U2509 (N_2509,N_2356,N_2343);
and U2510 (N_2510,N_2367,N_2232);
and U2511 (N_2511,N_2294,N_2298);
nand U2512 (N_2512,N_2383,N_2268);
or U2513 (N_2513,N_2367,N_2251);
nor U2514 (N_2514,N_2330,N_2366);
nor U2515 (N_2515,N_2367,N_2265);
and U2516 (N_2516,N_2216,N_2348);
nor U2517 (N_2517,N_2372,N_2340);
or U2518 (N_2518,N_2372,N_2259);
nand U2519 (N_2519,N_2345,N_2387);
and U2520 (N_2520,N_2302,N_2248);
or U2521 (N_2521,N_2239,N_2264);
nor U2522 (N_2522,N_2216,N_2317);
and U2523 (N_2523,N_2248,N_2220);
nand U2524 (N_2524,N_2365,N_2302);
and U2525 (N_2525,N_2315,N_2350);
nor U2526 (N_2526,N_2201,N_2281);
nor U2527 (N_2527,N_2228,N_2327);
or U2528 (N_2528,N_2392,N_2274);
and U2529 (N_2529,N_2348,N_2306);
or U2530 (N_2530,N_2250,N_2258);
or U2531 (N_2531,N_2245,N_2335);
nand U2532 (N_2532,N_2380,N_2293);
nor U2533 (N_2533,N_2319,N_2341);
and U2534 (N_2534,N_2303,N_2236);
and U2535 (N_2535,N_2218,N_2290);
nand U2536 (N_2536,N_2389,N_2352);
nor U2537 (N_2537,N_2379,N_2253);
and U2538 (N_2538,N_2232,N_2252);
and U2539 (N_2539,N_2300,N_2309);
or U2540 (N_2540,N_2390,N_2378);
nand U2541 (N_2541,N_2377,N_2279);
nand U2542 (N_2542,N_2361,N_2281);
and U2543 (N_2543,N_2322,N_2336);
nand U2544 (N_2544,N_2398,N_2233);
nor U2545 (N_2545,N_2236,N_2318);
nor U2546 (N_2546,N_2379,N_2202);
nor U2547 (N_2547,N_2246,N_2377);
and U2548 (N_2548,N_2294,N_2233);
nor U2549 (N_2549,N_2328,N_2388);
or U2550 (N_2550,N_2336,N_2213);
nand U2551 (N_2551,N_2220,N_2207);
nor U2552 (N_2552,N_2325,N_2395);
nand U2553 (N_2553,N_2294,N_2254);
or U2554 (N_2554,N_2202,N_2325);
or U2555 (N_2555,N_2200,N_2339);
nor U2556 (N_2556,N_2248,N_2393);
and U2557 (N_2557,N_2390,N_2339);
nor U2558 (N_2558,N_2303,N_2281);
nor U2559 (N_2559,N_2213,N_2221);
nor U2560 (N_2560,N_2398,N_2264);
or U2561 (N_2561,N_2294,N_2314);
or U2562 (N_2562,N_2279,N_2393);
nor U2563 (N_2563,N_2238,N_2315);
or U2564 (N_2564,N_2254,N_2343);
and U2565 (N_2565,N_2228,N_2284);
or U2566 (N_2566,N_2238,N_2382);
nor U2567 (N_2567,N_2228,N_2321);
xor U2568 (N_2568,N_2360,N_2358);
nand U2569 (N_2569,N_2274,N_2276);
nand U2570 (N_2570,N_2281,N_2259);
and U2571 (N_2571,N_2349,N_2313);
or U2572 (N_2572,N_2341,N_2307);
and U2573 (N_2573,N_2263,N_2387);
and U2574 (N_2574,N_2279,N_2385);
nand U2575 (N_2575,N_2253,N_2250);
nand U2576 (N_2576,N_2249,N_2362);
nor U2577 (N_2577,N_2340,N_2315);
or U2578 (N_2578,N_2332,N_2369);
nand U2579 (N_2579,N_2359,N_2297);
nor U2580 (N_2580,N_2279,N_2255);
and U2581 (N_2581,N_2207,N_2324);
or U2582 (N_2582,N_2244,N_2306);
and U2583 (N_2583,N_2259,N_2370);
or U2584 (N_2584,N_2343,N_2358);
nor U2585 (N_2585,N_2367,N_2394);
or U2586 (N_2586,N_2307,N_2308);
nand U2587 (N_2587,N_2236,N_2253);
or U2588 (N_2588,N_2329,N_2303);
nor U2589 (N_2589,N_2228,N_2271);
nor U2590 (N_2590,N_2298,N_2349);
and U2591 (N_2591,N_2232,N_2300);
nand U2592 (N_2592,N_2262,N_2211);
nor U2593 (N_2593,N_2325,N_2284);
or U2594 (N_2594,N_2304,N_2348);
nand U2595 (N_2595,N_2307,N_2251);
nand U2596 (N_2596,N_2267,N_2301);
nor U2597 (N_2597,N_2206,N_2358);
nand U2598 (N_2598,N_2215,N_2320);
nor U2599 (N_2599,N_2257,N_2391);
and U2600 (N_2600,N_2585,N_2445);
nor U2601 (N_2601,N_2437,N_2463);
and U2602 (N_2602,N_2479,N_2519);
or U2603 (N_2603,N_2521,N_2443);
nand U2604 (N_2604,N_2476,N_2529);
or U2605 (N_2605,N_2403,N_2552);
nor U2606 (N_2606,N_2475,N_2511);
nor U2607 (N_2607,N_2419,N_2592);
or U2608 (N_2608,N_2594,N_2471);
and U2609 (N_2609,N_2535,N_2520);
nor U2610 (N_2610,N_2565,N_2559);
nor U2611 (N_2611,N_2566,N_2489);
nand U2612 (N_2612,N_2451,N_2409);
or U2613 (N_2613,N_2591,N_2539);
or U2614 (N_2614,N_2444,N_2408);
or U2615 (N_2615,N_2527,N_2428);
nand U2616 (N_2616,N_2424,N_2434);
and U2617 (N_2617,N_2481,N_2537);
and U2618 (N_2618,N_2568,N_2447);
nor U2619 (N_2619,N_2599,N_2401);
nor U2620 (N_2620,N_2423,N_2415);
nand U2621 (N_2621,N_2438,N_2429);
or U2622 (N_2622,N_2458,N_2554);
xnor U2623 (N_2623,N_2459,N_2582);
nand U2624 (N_2624,N_2493,N_2503);
nor U2625 (N_2625,N_2461,N_2420);
nand U2626 (N_2626,N_2567,N_2465);
nand U2627 (N_2627,N_2536,N_2462);
xor U2628 (N_2628,N_2542,N_2439);
nor U2629 (N_2629,N_2596,N_2517);
nand U2630 (N_2630,N_2581,N_2460);
or U2631 (N_2631,N_2467,N_2449);
nand U2632 (N_2632,N_2558,N_2470);
nor U2633 (N_2633,N_2544,N_2422);
nor U2634 (N_2634,N_2486,N_2495);
nand U2635 (N_2635,N_2499,N_2487);
xnor U2636 (N_2636,N_2482,N_2598);
and U2637 (N_2637,N_2501,N_2534);
and U2638 (N_2638,N_2589,N_2518);
nand U2639 (N_2639,N_2411,N_2526);
nand U2640 (N_2640,N_2490,N_2509);
nand U2641 (N_2641,N_2498,N_2427);
nand U2642 (N_2642,N_2576,N_2546);
nor U2643 (N_2643,N_2450,N_2477);
and U2644 (N_2644,N_2553,N_2578);
nor U2645 (N_2645,N_2412,N_2530);
nor U2646 (N_2646,N_2421,N_2595);
and U2647 (N_2647,N_2506,N_2478);
nor U2648 (N_2648,N_2418,N_2496);
and U2649 (N_2649,N_2547,N_2522);
nand U2650 (N_2650,N_2525,N_2480);
and U2651 (N_2651,N_2452,N_2548);
or U2652 (N_2652,N_2538,N_2502);
xnor U2653 (N_2653,N_2484,N_2413);
or U2654 (N_2654,N_2483,N_2562);
or U2655 (N_2655,N_2402,N_2454);
or U2656 (N_2656,N_2466,N_2497);
nand U2657 (N_2657,N_2574,N_2563);
xnor U2658 (N_2658,N_2446,N_2405);
and U2659 (N_2659,N_2550,N_2456);
nand U2660 (N_2660,N_2431,N_2491);
nand U2661 (N_2661,N_2593,N_2572);
nor U2662 (N_2662,N_2485,N_2426);
nand U2663 (N_2663,N_2570,N_2441);
nor U2664 (N_2664,N_2551,N_2575);
nand U2665 (N_2665,N_2528,N_2400);
and U2666 (N_2666,N_2588,N_2440);
nand U2667 (N_2667,N_2543,N_2457);
nand U2668 (N_2668,N_2590,N_2507);
nor U2669 (N_2669,N_2455,N_2494);
or U2670 (N_2670,N_2407,N_2514);
nor U2671 (N_2671,N_2573,N_2580);
or U2672 (N_2672,N_2417,N_2579);
nor U2673 (N_2673,N_2523,N_2584);
nand U2674 (N_2674,N_2533,N_2513);
or U2675 (N_2675,N_2508,N_2469);
nand U2676 (N_2676,N_2472,N_2432);
or U2677 (N_2677,N_2510,N_2492);
nand U2678 (N_2678,N_2560,N_2549);
nor U2679 (N_2679,N_2433,N_2597);
or U2680 (N_2680,N_2435,N_2404);
nand U2681 (N_2681,N_2556,N_2557);
nor U2682 (N_2682,N_2430,N_2504);
nor U2683 (N_2683,N_2515,N_2505);
or U2684 (N_2684,N_2545,N_2436);
and U2685 (N_2685,N_2531,N_2524);
or U2686 (N_2686,N_2569,N_2416);
nand U2687 (N_2687,N_2410,N_2564);
nand U2688 (N_2688,N_2512,N_2540);
nand U2689 (N_2689,N_2571,N_2532);
nand U2690 (N_2690,N_2473,N_2561);
xor U2691 (N_2691,N_2516,N_2464);
or U2692 (N_2692,N_2453,N_2577);
or U2693 (N_2693,N_2414,N_2406);
and U2694 (N_2694,N_2442,N_2500);
nand U2695 (N_2695,N_2555,N_2587);
or U2696 (N_2696,N_2448,N_2468);
nor U2697 (N_2697,N_2425,N_2586);
nor U2698 (N_2698,N_2488,N_2541);
nand U2699 (N_2699,N_2583,N_2474);
nand U2700 (N_2700,N_2432,N_2521);
nor U2701 (N_2701,N_2552,N_2597);
and U2702 (N_2702,N_2503,N_2435);
nand U2703 (N_2703,N_2522,N_2500);
and U2704 (N_2704,N_2567,N_2515);
nand U2705 (N_2705,N_2498,N_2570);
nor U2706 (N_2706,N_2556,N_2424);
nand U2707 (N_2707,N_2423,N_2503);
nor U2708 (N_2708,N_2525,N_2466);
or U2709 (N_2709,N_2577,N_2572);
nand U2710 (N_2710,N_2435,N_2588);
nand U2711 (N_2711,N_2544,N_2593);
or U2712 (N_2712,N_2523,N_2502);
and U2713 (N_2713,N_2564,N_2447);
nand U2714 (N_2714,N_2522,N_2425);
or U2715 (N_2715,N_2506,N_2539);
nand U2716 (N_2716,N_2554,N_2475);
nor U2717 (N_2717,N_2543,N_2494);
or U2718 (N_2718,N_2508,N_2595);
nand U2719 (N_2719,N_2556,N_2448);
nor U2720 (N_2720,N_2523,N_2425);
nor U2721 (N_2721,N_2450,N_2586);
or U2722 (N_2722,N_2455,N_2433);
nand U2723 (N_2723,N_2486,N_2405);
and U2724 (N_2724,N_2503,N_2472);
xnor U2725 (N_2725,N_2438,N_2565);
or U2726 (N_2726,N_2489,N_2491);
or U2727 (N_2727,N_2509,N_2425);
nor U2728 (N_2728,N_2478,N_2514);
nor U2729 (N_2729,N_2494,N_2404);
nor U2730 (N_2730,N_2408,N_2424);
or U2731 (N_2731,N_2443,N_2566);
and U2732 (N_2732,N_2578,N_2551);
or U2733 (N_2733,N_2474,N_2415);
nand U2734 (N_2734,N_2522,N_2474);
nor U2735 (N_2735,N_2431,N_2437);
nand U2736 (N_2736,N_2525,N_2430);
and U2737 (N_2737,N_2459,N_2406);
and U2738 (N_2738,N_2530,N_2586);
nand U2739 (N_2739,N_2404,N_2416);
and U2740 (N_2740,N_2571,N_2474);
and U2741 (N_2741,N_2405,N_2537);
nand U2742 (N_2742,N_2470,N_2406);
nor U2743 (N_2743,N_2448,N_2450);
nor U2744 (N_2744,N_2561,N_2438);
nor U2745 (N_2745,N_2432,N_2547);
or U2746 (N_2746,N_2433,N_2591);
and U2747 (N_2747,N_2520,N_2549);
and U2748 (N_2748,N_2491,N_2521);
and U2749 (N_2749,N_2565,N_2431);
and U2750 (N_2750,N_2559,N_2479);
or U2751 (N_2751,N_2462,N_2535);
or U2752 (N_2752,N_2481,N_2588);
and U2753 (N_2753,N_2426,N_2440);
and U2754 (N_2754,N_2402,N_2467);
nand U2755 (N_2755,N_2474,N_2546);
nor U2756 (N_2756,N_2598,N_2406);
nand U2757 (N_2757,N_2408,N_2406);
nor U2758 (N_2758,N_2559,N_2598);
or U2759 (N_2759,N_2448,N_2411);
nor U2760 (N_2760,N_2540,N_2436);
nor U2761 (N_2761,N_2456,N_2494);
and U2762 (N_2762,N_2464,N_2511);
and U2763 (N_2763,N_2574,N_2439);
nand U2764 (N_2764,N_2513,N_2559);
and U2765 (N_2765,N_2478,N_2475);
nand U2766 (N_2766,N_2419,N_2595);
nor U2767 (N_2767,N_2572,N_2451);
nand U2768 (N_2768,N_2535,N_2410);
or U2769 (N_2769,N_2545,N_2520);
nand U2770 (N_2770,N_2512,N_2500);
or U2771 (N_2771,N_2402,N_2423);
nand U2772 (N_2772,N_2508,N_2473);
nor U2773 (N_2773,N_2592,N_2461);
nand U2774 (N_2774,N_2578,N_2478);
nand U2775 (N_2775,N_2540,N_2536);
nand U2776 (N_2776,N_2401,N_2439);
and U2777 (N_2777,N_2411,N_2443);
nor U2778 (N_2778,N_2592,N_2540);
and U2779 (N_2779,N_2502,N_2452);
and U2780 (N_2780,N_2476,N_2437);
xor U2781 (N_2781,N_2580,N_2406);
and U2782 (N_2782,N_2489,N_2450);
and U2783 (N_2783,N_2507,N_2485);
nor U2784 (N_2784,N_2545,N_2488);
nor U2785 (N_2785,N_2435,N_2419);
nor U2786 (N_2786,N_2428,N_2588);
and U2787 (N_2787,N_2566,N_2553);
nand U2788 (N_2788,N_2428,N_2526);
or U2789 (N_2789,N_2518,N_2555);
nand U2790 (N_2790,N_2410,N_2400);
nor U2791 (N_2791,N_2508,N_2597);
nor U2792 (N_2792,N_2539,N_2523);
nor U2793 (N_2793,N_2431,N_2599);
or U2794 (N_2794,N_2474,N_2558);
nand U2795 (N_2795,N_2497,N_2412);
or U2796 (N_2796,N_2514,N_2586);
and U2797 (N_2797,N_2598,N_2419);
nand U2798 (N_2798,N_2504,N_2449);
or U2799 (N_2799,N_2590,N_2569);
or U2800 (N_2800,N_2714,N_2603);
and U2801 (N_2801,N_2708,N_2717);
nor U2802 (N_2802,N_2604,N_2713);
or U2803 (N_2803,N_2752,N_2686);
or U2804 (N_2804,N_2790,N_2632);
and U2805 (N_2805,N_2631,N_2762);
and U2806 (N_2806,N_2666,N_2719);
nor U2807 (N_2807,N_2763,N_2778);
nand U2808 (N_2808,N_2723,N_2797);
nor U2809 (N_2809,N_2637,N_2698);
nand U2810 (N_2810,N_2675,N_2730);
or U2811 (N_2811,N_2724,N_2626);
nand U2812 (N_2812,N_2645,N_2676);
or U2813 (N_2813,N_2772,N_2774);
nand U2814 (N_2814,N_2712,N_2733);
xnor U2815 (N_2815,N_2649,N_2636);
nand U2816 (N_2816,N_2607,N_2753);
or U2817 (N_2817,N_2760,N_2629);
nand U2818 (N_2818,N_2639,N_2764);
nor U2819 (N_2819,N_2740,N_2776);
nand U2820 (N_2820,N_2608,N_2618);
nor U2821 (N_2821,N_2710,N_2702);
and U2822 (N_2822,N_2766,N_2646);
nor U2823 (N_2823,N_2784,N_2690);
or U2824 (N_2824,N_2788,N_2693);
nand U2825 (N_2825,N_2726,N_2602);
and U2826 (N_2826,N_2703,N_2643);
or U2827 (N_2827,N_2749,N_2659);
nand U2828 (N_2828,N_2695,N_2630);
nand U2829 (N_2829,N_2673,N_2707);
and U2830 (N_2830,N_2731,N_2728);
xor U2831 (N_2831,N_2794,N_2669);
nor U2832 (N_2832,N_2779,N_2616);
nand U2833 (N_2833,N_2701,N_2692);
nand U2834 (N_2834,N_2633,N_2667);
and U2835 (N_2835,N_2743,N_2605);
nor U2836 (N_2836,N_2715,N_2665);
nor U2837 (N_2837,N_2781,N_2606);
and U2838 (N_2838,N_2746,N_2700);
nor U2839 (N_2839,N_2647,N_2624);
or U2840 (N_2840,N_2769,N_2642);
and U2841 (N_2841,N_2796,N_2687);
nor U2842 (N_2842,N_2737,N_2601);
and U2843 (N_2843,N_2689,N_2711);
and U2844 (N_2844,N_2663,N_2734);
nand U2845 (N_2845,N_2732,N_2610);
nor U2846 (N_2846,N_2748,N_2651);
xor U2847 (N_2847,N_2777,N_2634);
or U2848 (N_2848,N_2680,N_2783);
or U2849 (N_2849,N_2775,N_2627);
and U2850 (N_2850,N_2621,N_2696);
or U2851 (N_2851,N_2614,N_2600);
nor U2852 (N_2852,N_2684,N_2706);
nor U2853 (N_2853,N_2765,N_2652);
nor U2854 (N_2854,N_2661,N_2793);
or U2855 (N_2855,N_2742,N_2694);
nand U2856 (N_2856,N_2741,N_2725);
or U2857 (N_2857,N_2699,N_2685);
and U2858 (N_2858,N_2780,N_2767);
or U2859 (N_2859,N_2674,N_2628);
and U2860 (N_2860,N_2678,N_2738);
or U2861 (N_2861,N_2739,N_2619);
nor U2862 (N_2862,N_2720,N_2620);
or U2863 (N_2863,N_2757,N_2611);
and U2864 (N_2864,N_2705,N_2670);
nand U2865 (N_2865,N_2750,N_2682);
nand U2866 (N_2866,N_2789,N_2795);
and U2867 (N_2867,N_2735,N_2615);
xor U2868 (N_2868,N_2770,N_2716);
nor U2869 (N_2869,N_2751,N_2657);
and U2870 (N_2870,N_2727,N_2679);
or U2871 (N_2871,N_2623,N_2736);
nor U2872 (N_2872,N_2722,N_2745);
or U2873 (N_2873,N_2653,N_2761);
and U2874 (N_2874,N_2759,N_2617);
or U2875 (N_2875,N_2635,N_2625);
or U2876 (N_2876,N_2613,N_2656);
or U2877 (N_2877,N_2688,N_2671);
nand U2878 (N_2878,N_2773,N_2787);
or U2879 (N_2879,N_2744,N_2785);
or U2880 (N_2880,N_2747,N_2758);
nor U2881 (N_2881,N_2799,N_2798);
or U2882 (N_2882,N_2786,N_2662);
and U2883 (N_2883,N_2622,N_2648);
nand U2884 (N_2884,N_2640,N_2683);
nor U2885 (N_2885,N_2718,N_2756);
nor U2886 (N_2886,N_2612,N_2677);
nand U2887 (N_2887,N_2768,N_2755);
or U2888 (N_2888,N_2609,N_2697);
or U2889 (N_2889,N_2672,N_2654);
nand U2890 (N_2890,N_2655,N_2644);
or U2891 (N_2891,N_2691,N_2709);
and U2892 (N_2892,N_2650,N_2771);
or U2893 (N_2893,N_2638,N_2658);
or U2894 (N_2894,N_2681,N_2782);
nand U2895 (N_2895,N_2660,N_2754);
nand U2896 (N_2896,N_2792,N_2704);
and U2897 (N_2897,N_2641,N_2729);
nand U2898 (N_2898,N_2791,N_2664);
nand U2899 (N_2899,N_2668,N_2721);
and U2900 (N_2900,N_2611,N_2607);
nand U2901 (N_2901,N_2788,N_2761);
nand U2902 (N_2902,N_2761,N_2601);
or U2903 (N_2903,N_2618,N_2791);
and U2904 (N_2904,N_2611,N_2713);
and U2905 (N_2905,N_2605,N_2645);
nor U2906 (N_2906,N_2616,N_2689);
nor U2907 (N_2907,N_2793,N_2769);
nor U2908 (N_2908,N_2673,N_2646);
xor U2909 (N_2909,N_2764,N_2602);
or U2910 (N_2910,N_2750,N_2647);
and U2911 (N_2911,N_2611,N_2696);
nand U2912 (N_2912,N_2652,N_2728);
and U2913 (N_2913,N_2714,N_2726);
and U2914 (N_2914,N_2767,N_2716);
nand U2915 (N_2915,N_2622,N_2726);
nand U2916 (N_2916,N_2620,N_2716);
nand U2917 (N_2917,N_2780,N_2677);
and U2918 (N_2918,N_2625,N_2705);
xnor U2919 (N_2919,N_2713,N_2795);
or U2920 (N_2920,N_2739,N_2638);
and U2921 (N_2921,N_2625,N_2606);
nand U2922 (N_2922,N_2768,N_2776);
nor U2923 (N_2923,N_2778,N_2739);
or U2924 (N_2924,N_2738,N_2785);
nor U2925 (N_2925,N_2715,N_2763);
xor U2926 (N_2926,N_2731,N_2748);
or U2927 (N_2927,N_2769,N_2648);
nand U2928 (N_2928,N_2706,N_2609);
or U2929 (N_2929,N_2775,N_2617);
and U2930 (N_2930,N_2794,N_2667);
nand U2931 (N_2931,N_2736,N_2773);
nor U2932 (N_2932,N_2660,N_2676);
and U2933 (N_2933,N_2759,N_2676);
and U2934 (N_2934,N_2607,N_2625);
nand U2935 (N_2935,N_2676,N_2737);
or U2936 (N_2936,N_2652,N_2676);
and U2937 (N_2937,N_2694,N_2788);
nand U2938 (N_2938,N_2600,N_2758);
nand U2939 (N_2939,N_2792,N_2621);
nor U2940 (N_2940,N_2719,N_2623);
nor U2941 (N_2941,N_2773,N_2614);
nor U2942 (N_2942,N_2705,N_2757);
nor U2943 (N_2943,N_2659,N_2652);
and U2944 (N_2944,N_2708,N_2697);
and U2945 (N_2945,N_2742,N_2789);
nand U2946 (N_2946,N_2623,N_2754);
nand U2947 (N_2947,N_2795,N_2708);
and U2948 (N_2948,N_2609,N_2756);
or U2949 (N_2949,N_2637,N_2798);
nand U2950 (N_2950,N_2655,N_2600);
or U2951 (N_2951,N_2792,N_2747);
nand U2952 (N_2952,N_2616,N_2704);
nand U2953 (N_2953,N_2720,N_2665);
or U2954 (N_2954,N_2644,N_2713);
and U2955 (N_2955,N_2773,N_2777);
nand U2956 (N_2956,N_2693,N_2681);
and U2957 (N_2957,N_2774,N_2715);
nor U2958 (N_2958,N_2639,N_2715);
and U2959 (N_2959,N_2638,N_2641);
and U2960 (N_2960,N_2725,N_2640);
and U2961 (N_2961,N_2774,N_2736);
nor U2962 (N_2962,N_2784,N_2605);
nor U2963 (N_2963,N_2726,N_2723);
xnor U2964 (N_2964,N_2778,N_2605);
and U2965 (N_2965,N_2605,N_2681);
nor U2966 (N_2966,N_2690,N_2646);
and U2967 (N_2967,N_2714,N_2787);
and U2968 (N_2968,N_2751,N_2766);
nand U2969 (N_2969,N_2776,N_2648);
and U2970 (N_2970,N_2714,N_2612);
nor U2971 (N_2971,N_2762,N_2771);
nand U2972 (N_2972,N_2669,N_2641);
nand U2973 (N_2973,N_2607,N_2641);
and U2974 (N_2974,N_2635,N_2716);
nand U2975 (N_2975,N_2764,N_2735);
nor U2976 (N_2976,N_2643,N_2791);
nor U2977 (N_2977,N_2665,N_2703);
or U2978 (N_2978,N_2680,N_2726);
nor U2979 (N_2979,N_2772,N_2671);
nor U2980 (N_2980,N_2670,N_2738);
and U2981 (N_2981,N_2780,N_2667);
nand U2982 (N_2982,N_2786,N_2655);
nand U2983 (N_2983,N_2633,N_2651);
or U2984 (N_2984,N_2623,N_2739);
nand U2985 (N_2985,N_2704,N_2713);
nor U2986 (N_2986,N_2664,N_2735);
and U2987 (N_2987,N_2677,N_2769);
nand U2988 (N_2988,N_2758,N_2620);
nor U2989 (N_2989,N_2782,N_2728);
and U2990 (N_2990,N_2725,N_2737);
or U2991 (N_2991,N_2686,N_2652);
or U2992 (N_2992,N_2603,N_2728);
nor U2993 (N_2993,N_2609,N_2653);
or U2994 (N_2994,N_2641,N_2640);
and U2995 (N_2995,N_2617,N_2624);
or U2996 (N_2996,N_2721,N_2716);
or U2997 (N_2997,N_2695,N_2688);
or U2998 (N_2998,N_2661,N_2625);
nor U2999 (N_2999,N_2687,N_2648);
or U3000 (N_3000,N_2894,N_2898);
nand U3001 (N_3001,N_2833,N_2990);
nor U3002 (N_3002,N_2836,N_2913);
nand U3003 (N_3003,N_2828,N_2960);
and U3004 (N_3004,N_2962,N_2947);
nor U3005 (N_3005,N_2994,N_2955);
nor U3006 (N_3006,N_2937,N_2995);
or U3007 (N_3007,N_2840,N_2901);
nor U3008 (N_3008,N_2907,N_2897);
or U3009 (N_3009,N_2862,N_2817);
nand U3010 (N_3010,N_2920,N_2954);
or U3011 (N_3011,N_2977,N_2802);
nor U3012 (N_3012,N_2880,N_2972);
nand U3013 (N_3013,N_2905,N_2838);
or U3014 (N_3014,N_2826,N_2900);
and U3015 (N_3015,N_2858,N_2927);
nor U3016 (N_3016,N_2822,N_2861);
and U3017 (N_3017,N_2896,N_2850);
nor U3018 (N_3018,N_2957,N_2976);
or U3019 (N_3019,N_2866,N_2946);
and U3020 (N_3020,N_2971,N_2892);
or U3021 (N_3021,N_2811,N_2899);
or U3022 (N_3022,N_2909,N_2945);
nand U3023 (N_3023,N_2842,N_2872);
and U3024 (N_3024,N_2806,N_2925);
nor U3025 (N_3025,N_2846,N_2854);
nor U3026 (N_3026,N_2983,N_2928);
and U3027 (N_3027,N_2904,N_2871);
or U3028 (N_3028,N_2956,N_2870);
or U3029 (N_3029,N_2810,N_2986);
or U3030 (N_3030,N_2888,N_2875);
and U3031 (N_3031,N_2819,N_2936);
and U3032 (N_3032,N_2951,N_2996);
or U3033 (N_3033,N_2804,N_2939);
nand U3034 (N_3034,N_2910,N_2825);
nand U3035 (N_3035,N_2933,N_2938);
nand U3036 (N_3036,N_2919,N_2827);
nand U3037 (N_3037,N_2885,N_2863);
nand U3038 (N_3038,N_2815,N_2921);
nor U3039 (N_3039,N_2940,N_2856);
and U3040 (N_3040,N_2975,N_2845);
or U3041 (N_3041,N_2903,N_2834);
and U3042 (N_3042,N_2934,N_2948);
or U3043 (N_3043,N_2999,N_2969);
and U3044 (N_3044,N_2891,N_2997);
or U3045 (N_3045,N_2924,N_2857);
and U3046 (N_3046,N_2931,N_2916);
nor U3047 (N_3047,N_2941,N_2908);
and U3048 (N_3048,N_2922,N_2849);
nand U3049 (N_3049,N_2998,N_2816);
xor U3050 (N_3050,N_2841,N_2988);
nand U3051 (N_3051,N_2855,N_2984);
or U3052 (N_3052,N_2801,N_2805);
nor U3053 (N_3053,N_2967,N_2982);
nand U3054 (N_3054,N_2964,N_2843);
and U3055 (N_3055,N_2942,N_2832);
nand U3056 (N_3056,N_2800,N_2930);
nor U3057 (N_3057,N_2820,N_2873);
nand U3058 (N_3058,N_2869,N_2813);
nand U3059 (N_3059,N_2963,N_2879);
and U3060 (N_3060,N_2886,N_2902);
nor U3061 (N_3061,N_2917,N_2966);
nor U3062 (N_3062,N_2884,N_2914);
nor U3063 (N_3063,N_2821,N_2965);
or U3064 (N_3064,N_2835,N_2944);
nor U3065 (N_3065,N_2803,N_2868);
or U3066 (N_3066,N_2847,N_2809);
xnor U3067 (N_3067,N_2980,N_2959);
nor U3068 (N_3068,N_2915,N_2859);
and U3069 (N_3069,N_2895,N_2852);
and U3070 (N_3070,N_2961,N_2993);
nor U3071 (N_3071,N_2887,N_2987);
nand U3072 (N_3072,N_2818,N_2851);
nand U3073 (N_3073,N_2839,N_2974);
nand U3074 (N_3074,N_2853,N_2973);
and U3075 (N_3075,N_2932,N_2935);
and U3076 (N_3076,N_2923,N_2985);
and U3077 (N_3077,N_2848,N_2953);
nand U3078 (N_3078,N_2978,N_2949);
nor U3079 (N_3079,N_2989,N_2874);
and U3080 (N_3080,N_2883,N_2968);
and U3081 (N_3081,N_2808,N_2865);
nor U3082 (N_3082,N_2918,N_2970);
and U3083 (N_3083,N_2981,N_2889);
and U3084 (N_3084,N_2823,N_2824);
nand U3085 (N_3085,N_2814,N_2882);
nor U3086 (N_3086,N_2831,N_2844);
or U3087 (N_3087,N_2830,N_2890);
xnor U3088 (N_3088,N_2979,N_2992);
or U3089 (N_3089,N_2952,N_2829);
and U3090 (N_3090,N_2881,N_2929);
nor U3091 (N_3091,N_2860,N_2906);
or U3092 (N_3092,N_2837,N_2911);
or U3093 (N_3093,N_2893,N_2812);
nor U3094 (N_3094,N_2878,N_2867);
or U3095 (N_3095,N_2950,N_2877);
and U3096 (N_3096,N_2807,N_2958);
nand U3097 (N_3097,N_2876,N_2991);
nand U3098 (N_3098,N_2864,N_2943);
nand U3099 (N_3099,N_2926,N_2912);
or U3100 (N_3100,N_2961,N_2807);
nand U3101 (N_3101,N_2947,N_2955);
nor U3102 (N_3102,N_2804,N_2886);
xor U3103 (N_3103,N_2989,N_2814);
and U3104 (N_3104,N_2972,N_2818);
and U3105 (N_3105,N_2815,N_2881);
nor U3106 (N_3106,N_2875,N_2851);
and U3107 (N_3107,N_2865,N_2999);
nand U3108 (N_3108,N_2801,N_2993);
nand U3109 (N_3109,N_2810,N_2860);
nand U3110 (N_3110,N_2923,N_2984);
nor U3111 (N_3111,N_2932,N_2854);
xnor U3112 (N_3112,N_2950,N_2927);
or U3113 (N_3113,N_2898,N_2802);
nor U3114 (N_3114,N_2943,N_2818);
or U3115 (N_3115,N_2802,N_2833);
nor U3116 (N_3116,N_2868,N_2871);
and U3117 (N_3117,N_2825,N_2911);
nand U3118 (N_3118,N_2848,N_2820);
nor U3119 (N_3119,N_2906,N_2850);
or U3120 (N_3120,N_2923,N_2991);
or U3121 (N_3121,N_2959,N_2946);
or U3122 (N_3122,N_2835,N_2898);
nand U3123 (N_3123,N_2937,N_2856);
nor U3124 (N_3124,N_2993,N_2995);
xor U3125 (N_3125,N_2825,N_2916);
or U3126 (N_3126,N_2982,N_2819);
nand U3127 (N_3127,N_2953,N_2863);
and U3128 (N_3128,N_2907,N_2814);
nand U3129 (N_3129,N_2892,N_2872);
and U3130 (N_3130,N_2826,N_2843);
and U3131 (N_3131,N_2811,N_2881);
or U3132 (N_3132,N_2874,N_2992);
nand U3133 (N_3133,N_2917,N_2897);
nor U3134 (N_3134,N_2847,N_2825);
nand U3135 (N_3135,N_2831,N_2980);
or U3136 (N_3136,N_2927,N_2855);
nor U3137 (N_3137,N_2965,N_2959);
and U3138 (N_3138,N_2949,N_2970);
or U3139 (N_3139,N_2872,N_2826);
and U3140 (N_3140,N_2909,N_2873);
or U3141 (N_3141,N_2909,N_2951);
and U3142 (N_3142,N_2976,N_2829);
nor U3143 (N_3143,N_2800,N_2927);
nor U3144 (N_3144,N_2832,N_2847);
and U3145 (N_3145,N_2981,N_2859);
nand U3146 (N_3146,N_2958,N_2823);
nor U3147 (N_3147,N_2830,N_2862);
nor U3148 (N_3148,N_2851,N_2955);
or U3149 (N_3149,N_2810,N_2900);
and U3150 (N_3150,N_2999,N_2916);
or U3151 (N_3151,N_2947,N_2949);
or U3152 (N_3152,N_2903,N_2942);
nor U3153 (N_3153,N_2864,N_2984);
or U3154 (N_3154,N_2890,N_2962);
xnor U3155 (N_3155,N_2950,N_2962);
nor U3156 (N_3156,N_2977,N_2986);
nor U3157 (N_3157,N_2803,N_2866);
nand U3158 (N_3158,N_2829,N_2964);
nand U3159 (N_3159,N_2985,N_2827);
nor U3160 (N_3160,N_2967,N_2899);
and U3161 (N_3161,N_2844,N_2819);
or U3162 (N_3162,N_2954,N_2918);
nor U3163 (N_3163,N_2932,N_2997);
nor U3164 (N_3164,N_2867,N_2865);
xnor U3165 (N_3165,N_2908,N_2838);
or U3166 (N_3166,N_2938,N_2951);
and U3167 (N_3167,N_2952,N_2892);
and U3168 (N_3168,N_2930,N_2968);
nand U3169 (N_3169,N_2817,N_2897);
nand U3170 (N_3170,N_2933,N_2814);
nand U3171 (N_3171,N_2971,N_2907);
nand U3172 (N_3172,N_2995,N_2874);
and U3173 (N_3173,N_2950,N_2888);
nand U3174 (N_3174,N_2932,N_2861);
and U3175 (N_3175,N_2906,N_2896);
nand U3176 (N_3176,N_2946,N_2855);
and U3177 (N_3177,N_2903,N_2840);
nor U3178 (N_3178,N_2819,N_2988);
nor U3179 (N_3179,N_2887,N_2807);
nor U3180 (N_3180,N_2808,N_2983);
nand U3181 (N_3181,N_2959,N_2816);
nand U3182 (N_3182,N_2829,N_2833);
and U3183 (N_3183,N_2802,N_2896);
or U3184 (N_3184,N_2873,N_2801);
nor U3185 (N_3185,N_2907,N_2807);
and U3186 (N_3186,N_2853,N_2920);
and U3187 (N_3187,N_2905,N_2855);
or U3188 (N_3188,N_2845,N_2979);
nand U3189 (N_3189,N_2955,N_2978);
nor U3190 (N_3190,N_2912,N_2939);
nor U3191 (N_3191,N_2842,N_2822);
nor U3192 (N_3192,N_2877,N_2911);
and U3193 (N_3193,N_2832,N_2921);
nand U3194 (N_3194,N_2944,N_2985);
or U3195 (N_3195,N_2958,N_2940);
or U3196 (N_3196,N_2909,N_2935);
and U3197 (N_3197,N_2966,N_2842);
and U3198 (N_3198,N_2837,N_2868);
nand U3199 (N_3199,N_2892,N_2982);
or U3200 (N_3200,N_3124,N_3079);
or U3201 (N_3201,N_3107,N_3104);
and U3202 (N_3202,N_3047,N_3036);
nor U3203 (N_3203,N_3160,N_3067);
nand U3204 (N_3204,N_3078,N_3123);
or U3205 (N_3205,N_3140,N_3028);
or U3206 (N_3206,N_3093,N_3087);
and U3207 (N_3207,N_3086,N_3142);
xor U3208 (N_3208,N_3074,N_3152);
nand U3209 (N_3209,N_3131,N_3003);
nor U3210 (N_3210,N_3014,N_3026);
nand U3211 (N_3211,N_3133,N_3141);
nand U3212 (N_3212,N_3055,N_3072);
and U3213 (N_3213,N_3147,N_3061);
nor U3214 (N_3214,N_3151,N_3189);
or U3215 (N_3215,N_3020,N_3195);
nor U3216 (N_3216,N_3037,N_3029);
or U3217 (N_3217,N_3091,N_3044);
nor U3218 (N_3218,N_3135,N_3185);
or U3219 (N_3219,N_3052,N_3157);
or U3220 (N_3220,N_3143,N_3111);
or U3221 (N_3221,N_3166,N_3114);
and U3222 (N_3222,N_3184,N_3175);
and U3223 (N_3223,N_3009,N_3153);
nor U3224 (N_3224,N_3012,N_3005);
or U3225 (N_3225,N_3064,N_3176);
nor U3226 (N_3226,N_3181,N_3180);
nor U3227 (N_3227,N_3187,N_3042);
nor U3228 (N_3228,N_3008,N_3069);
nor U3229 (N_3229,N_3100,N_3034);
nor U3230 (N_3230,N_3198,N_3172);
and U3231 (N_3231,N_3109,N_3057);
or U3232 (N_3232,N_3173,N_3122);
nor U3233 (N_3233,N_3018,N_3070);
or U3234 (N_3234,N_3178,N_3040);
and U3235 (N_3235,N_3156,N_3154);
and U3236 (N_3236,N_3085,N_3048);
and U3237 (N_3237,N_3027,N_3144);
nand U3238 (N_3238,N_3098,N_3192);
nand U3239 (N_3239,N_3179,N_3056);
or U3240 (N_3240,N_3065,N_3138);
or U3241 (N_3241,N_3121,N_3102);
nor U3242 (N_3242,N_3108,N_3071);
nand U3243 (N_3243,N_3060,N_3148);
nand U3244 (N_3244,N_3115,N_3103);
nand U3245 (N_3245,N_3099,N_3063);
and U3246 (N_3246,N_3191,N_3168);
nor U3247 (N_3247,N_3149,N_3022);
nand U3248 (N_3248,N_3075,N_3088);
and U3249 (N_3249,N_3039,N_3132);
nor U3250 (N_3250,N_3158,N_3171);
and U3251 (N_3251,N_3053,N_3139);
or U3252 (N_3252,N_3011,N_3083);
or U3253 (N_3253,N_3177,N_3117);
or U3254 (N_3254,N_3013,N_3035);
or U3255 (N_3255,N_3095,N_3089);
or U3256 (N_3256,N_3193,N_3110);
and U3257 (N_3257,N_3119,N_3188);
or U3258 (N_3258,N_3167,N_3164);
or U3259 (N_3259,N_3186,N_3058);
xor U3260 (N_3260,N_3015,N_3162);
or U3261 (N_3261,N_3050,N_3054);
nand U3262 (N_3262,N_3082,N_3137);
or U3263 (N_3263,N_3182,N_3174);
or U3264 (N_3264,N_3031,N_3017);
and U3265 (N_3265,N_3010,N_3016);
xor U3266 (N_3266,N_3000,N_3112);
and U3267 (N_3267,N_3073,N_3023);
nand U3268 (N_3268,N_3116,N_3077);
or U3269 (N_3269,N_3183,N_3128);
and U3270 (N_3270,N_3006,N_3045);
and U3271 (N_3271,N_3066,N_3097);
or U3272 (N_3272,N_3190,N_3041);
or U3273 (N_3273,N_3076,N_3094);
nand U3274 (N_3274,N_3113,N_3051);
nor U3275 (N_3275,N_3106,N_3049);
or U3276 (N_3276,N_3062,N_3165);
nand U3277 (N_3277,N_3161,N_3118);
nor U3278 (N_3278,N_3136,N_3068);
nor U3279 (N_3279,N_3120,N_3197);
and U3280 (N_3280,N_3092,N_3130);
or U3281 (N_3281,N_3199,N_3025);
and U3282 (N_3282,N_3169,N_3038);
or U3283 (N_3283,N_3196,N_3163);
nor U3284 (N_3284,N_3134,N_3080);
nand U3285 (N_3285,N_3155,N_3125);
and U3286 (N_3286,N_3105,N_3101);
nor U3287 (N_3287,N_3150,N_3081);
nor U3288 (N_3288,N_3033,N_3001);
nand U3289 (N_3289,N_3059,N_3145);
or U3290 (N_3290,N_3194,N_3030);
and U3291 (N_3291,N_3021,N_3096);
and U3292 (N_3292,N_3032,N_3007);
nand U3293 (N_3293,N_3129,N_3084);
and U3294 (N_3294,N_3127,N_3024);
xnor U3295 (N_3295,N_3043,N_3004);
nor U3296 (N_3296,N_3126,N_3170);
and U3297 (N_3297,N_3046,N_3146);
nor U3298 (N_3298,N_3159,N_3090);
and U3299 (N_3299,N_3002,N_3019);
nand U3300 (N_3300,N_3044,N_3185);
and U3301 (N_3301,N_3053,N_3183);
nor U3302 (N_3302,N_3156,N_3135);
or U3303 (N_3303,N_3116,N_3194);
xor U3304 (N_3304,N_3154,N_3041);
and U3305 (N_3305,N_3146,N_3105);
and U3306 (N_3306,N_3012,N_3089);
or U3307 (N_3307,N_3095,N_3173);
or U3308 (N_3308,N_3195,N_3146);
and U3309 (N_3309,N_3158,N_3058);
nand U3310 (N_3310,N_3153,N_3000);
and U3311 (N_3311,N_3089,N_3056);
or U3312 (N_3312,N_3179,N_3051);
nor U3313 (N_3313,N_3046,N_3019);
nand U3314 (N_3314,N_3187,N_3169);
nand U3315 (N_3315,N_3086,N_3056);
and U3316 (N_3316,N_3131,N_3199);
nor U3317 (N_3317,N_3027,N_3100);
or U3318 (N_3318,N_3107,N_3180);
nand U3319 (N_3319,N_3010,N_3047);
nand U3320 (N_3320,N_3140,N_3054);
nand U3321 (N_3321,N_3134,N_3123);
nor U3322 (N_3322,N_3198,N_3136);
or U3323 (N_3323,N_3045,N_3000);
and U3324 (N_3324,N_3159,N_3099);
nor U3325 (N_3325,N_3075,N_3141);
nand U3326 (N_3326,N_3064,N_3016);
nor U3327 (N_3327,N_3185,N_3028);
nand U3328 (N_3328,N_3149,N_3036);
nor U3329 (N_3329,N_3151,N_3056);
or U3330 (N_3330,N_3106,N_3063);
nand U3331 (N_3331,N_3191,N_3149);
and U3332 (N_3332,N_3197,N_3155);
or U3333 (N_3333,N_3018,N_3007);
xor U3334 (N_3334,N_3013,N_3075);
and U3335 (N_3335,N_3165,N_3087);
and U3336 (N_3336,N_3105,N_3063);
or U3337 (N_3337,N_3160,N_3028);
or U3338 (N_3338,N_3046,N_3017);
or U3339 (N_3339,N_3180,N_3084);
nand U3340 (N_3340,N_3114,N_3025);
nand U3341 (N_3341,N_3161,N_3002);
nand U3342 (N_3342,N_3161,N_3155);
nor U3343 (N_3343,N_3059,N_3077);
nor U3344 (N_3344,N_3132,N_3066);
nor U3345 (N_3345,N_3085,N_3011);
nand U3346 (N_3346,N_3199,N_3039);
and U3347 (N_3347,N_3010,N_3141);
and U3348 (N_3348,N_3115,N_3137);
nand U3349 (N_3349,N_3067,N_3036);
and U3350 (N_3350,N_3127,N_3161);
nand U3351 (N_3351,N_3175,N_3021);
nor U3352 (N_3352,N_3192,N_3028);
nor U3353 (N_3353,N_3121,N_3022);
and U3354 (N_3354,N_3028,N_3029);
or U3355 (N_3355,N_3151,N_3114);
nor U3356 (N_3356,N_3091,N_3157);
nand U3357 (N_3357,N_3154,N_3024);
or U3358 (N_3358,N_3157,N_3080);
or U3359 (N_3359,N_3027,N_3069);
and U3360 (N_3360,N_3030,N_3145);
or U3361 (N_3361,N_3018,N_3020);
nor U3362 (N_3362,N_3022,N_3197);
or U3363 (N_3363,N_3030,N_3095);
or U3364 (N_3364,N_3182,N_3185);
and U3365 (N_3365,N_3126,N_3138);
or U3366 (N_3366,N_3074,N_3092);
nor U3367 (N_3367,N_3133,N_3082);
and U3368 (N_3368,N_3139,N_3103);
or U3369 (N_3369,N_3146,N_3040);
nand U3370 (N_3370,N_3111,N_3157);
or U3371 (N_3371,N_3116,N_3196);
nand U3372 (N_3372,N_3097,N_3182);
xor U3373 (N_3373,N_3078,N_3173);
and U3374 (N_3374,N_3047,N_3025);
nand U3375 (N_3375,N_3155,N_3111);
nand U3376 (N_3376,N_3000,N_3116);
and U3377 (N_3377,N_3146,N_3082);
or U3378 (N_3378,N_3110,N_3042);
nor U3379 (N_3379,N_3044,N_3134);
or U3380 (N_3380,N_3004,N_3011);
and U3381 (N_3381,N_3112,N_3045);
nand U3382 (N_3382,N_3140,N_3084);
or U3383 (N_3383,N_3022,N_3179);
or U3384 (N_3384,N_3039,N_3064);
nand U3385 (N_3385,N_3193,N_3095);
nor U3386 (N_3386,N_3055,N_3110);
nand U3387 (N_3387,N_3012,N_3074);
nand U3388 (N_3388,N_3114,N_3061);
or U3389 (N_3389,N_3136,N_3059);
nor U3390 (N_3390,N_3133,N_3062);
or U3391 (N_3391,N_3110,N_3065);
or U3392 (N_3392,N_3084,N_3112);
nor U3393 (N_3393,N_3157,N_3044);
or U3394 (N_3394,N_3079,N_3156);
nor U3395 (N_3395,N_3092,N_3190);
nand U3396 (N_3396,N_3126,N_3166);
nand U3397 (N_3397,N_3187,N_3007);
nor U3398 (N_3398,N_3132,N_3031);
nand U3399 (N_3399,N_3004,N_3087);
nand U3400 (N_3400,N_3318,N_3281);
and U3401 (N_3401,N_3364,N_3291);
nand U3402 (N_3402,N_3377,N_3201);
nor U3403 (N_3403,N_3257,N_3379);
nor U3404 (N_3404,N_3299,N_3380);
or U3405 (N_3405,N_3320,N_3374);
nor U3406 (N_3406,N_3242,N_3256);
and U3407 (N_3407,N_3203,N_3208);
or U3408 (N_3408,N_3362,N_3258);
nand U3409 (N_3409,N_3344,N_3333);
and U3410 (N_3410,N_3357,N_3298);
nand U3411 (N_3411,N_3313,N_3340);
nand U3412 (N_3412,N_3207,N_3370);
and U3413 (N_3413,N_3330,N_3202);
nor U3414 (N_3414,N_3285,N_3260);
and U3415 (N_3415,N_3269,N_3367);
xor U3416 (N_3416,N_3317,N_3388);
nor U3417 (N_3417,N_3225,N_3234);
or U3418 (N_3418,N_3227,N_3326);
nor U3419 (N_3419,N_3251,N_3384);
nand U3420 (N_3420,N_3275,N_3286);
nand U3421 (N_3421,N_3381,N_3372);
nor U3422 (N_3422,N_3343,N_3399);
nor U3423 (N_3423,N_3394,N_3383);
nand U3424 (N_3424,N_3355,N_3277);
or U3425 (N_3425,N_3352,N_3274);
xor U3426 (N_3426,N_3235,N_3241);
or U3427 (N_3427,N_3327,N_3324);
or U3428 (N_3428,N_3297,N_3224);
or U3429 (N_3429,N_3211,N_3284);
nand U3430 (N_3430,N_3263,N_3249);
nor U3431 (N_3431,N_3204,N_3378);
xor U3432 (N_3432,N_3243,N_3282);
xnor U3433 (N_3433,N_3215,N_3393);
nand U3434 (N_3434,N_3386,N_3230);
or U3435 (N_3435,N_3279,N_3398);
nor U3436 (N_3436,N_3329,N_3363);
nor U3437 (N_3437,N_3228,N_3319);
nor U3438 (N_3438,N_3237,N_3309);
and U3439 (N_3439,N_3345,N_3236);
nor U3440 (N_3440,N_3311,N_3238);
nor U3441 (N_3441,N_3390,N_3337);
nand U3442 (N_3442,N_3210,N_3356);
and U3443 (N_3443,N_3253,N_3255);
nand U3444 (N_3444,N_3233,N_3310);
and U3445 (N_3445,N_3273,N_3325);
nor U3446 (N_3446,N_3359,N_3396);
or U3447 (N_3447,N_3248,N_3358);
or U3448 (N_3448,N_3395,N_3302);
and U3449 (N_3449,N_3246,N_3371);
nand U3450 (N_3450,N_3220,N_3219);
and U3451 (N_3451,N_3290,N_3397);
xnor U3452 (N_3452,N_3217,N_3366);
and U3453 (N_3453,N_3240,N_3289);
nand U3454 (N_3454,N_3332,N_3308);
nor U3455 (N_3455,N_3369,N_3321);
nand U3456 (N_3456,N_3250,N_3296);
nand U3457 (N_3457,N_3247,N_3391);
nand U3458 (N_3458,N_3385,N_3365);
nand U3459 (N_3459,N_3259,N_3373);
and U3460 (N_3460,N_3331,N_3382);
or U3461 (N_3461,N_3209,N_3389);
and U3462 (N_3462,N_3295,N_3262);
xnor U3463 (N_3463,N_3288,N_3231);
nand U3464 (N_3464,N_3341,N_3301);
and U3465 (N_3465,N_3342,N_3205);
nand U3466 (N_3466,N_3351,N_3218);
nand U3467 (N_3467,N_3214,N_3361);
or U3468 (N_3468,N_3354,N_3283);
xor U3469 (N_3469,N_3254,N_3323);
xnor U3470 (N_3470,N_3307,N_3222);
nand U3471 (N_3471,N_3353,N_3270);
xnor U3472 (N_3472,N_3206,N_3347);
nand U3473 (N_3473,N_3272,N_3265);
and U3474 (N_3474,N_3264,N_3306);
nand U3475 (N_3475,N_3314,N_3293);
and U3476 (N_3476,N_3221,N_3223);
and U3477 (N_3477,N_3348,N_3267);
nand U3478 (N_3478,N_3280,N_3226);
and U3479 (N_3479,N_3316,N_3294);
nor U3480 (N_3480,N_3334,N_3244);
or U3481 (N_3481,N_3229,N_3252);
nor U3482 (N_3482,N_3276,N_3245);
and U3483 (N_3483,N_3305,N_3335);
nor U3484 (N_3484,N_3387,N_3315);
xnor U3485 (N_3485,N_3278,N_3216);
nand U3486 (N_3486,N_3349,N_3287);
nor U3487 (N_3487,N_3261,N_3322);
or U3488 (N_3488,N_3266,N_3338);
or U3489 (N_3489,N_3312,N_3303);
or U3490 (N_3490,N_3300,N_3368);
nand U3491 (N_3491,N_3328,N_3239);
nand U3492 (N_3492,N_3350,N_3376);
or U3493 (N_3493,N_3336,N_3339);
nand U3494 (N_3494,N_3360,N_3213);
xnor U3495 (N_3495,N_3346,N_3212);
or U3496 (N_3496,N_3392,N_3200);
nor U3497 (N_3497,N_3375,N_3232);
nor U3498 (N_3498,N_3292,N_3271);
nor U3499 (N_3499,N_3304,N_3268);
and U3500 (N_3500,N_3206,N_3392);
and U3501 (N_3501,N_3346,N_3224);
or U3502 (N_3502,N_3398,N_3364);
nand U3503 (N_3503,N_3247,N_3227);
xor U3504 (N_3504,N_3318,N_3309);
nor U3505 (N_3505,N_3330,N_3226);
nand U3506 (N_3506,N_3281,N_3203);
or U3507 (N_3507,N_3385,N_3276);
nand U3508 (N_3508,N_3385,N_3357);
and U3509 (N_3509,N_3369,N_3209);
nand U3510 (N_3510,N_3317,N_3280);
nand U3511 (N_3511,N_3274,N_3320);
or U3512 (N_3512,N_3222,N_3349);
or U3513 (N_3513,N_3311,N_3261);
and U3514 (N_3514,N_3318,N_3310);
nor U3515 (N_3515,N_3241,N_3315);
or U3516 (N_3516,N_3239,N_3319);
nor U3517 (N_3517,N_3338,N_3357);
or U3518 (N_3518,N_3387,N_3235);
or U3519 (N_3519,N_3224,N_3212);
or U3520 (N_3520,N_3244,N_3266);
nor U3521 (N_3521,N_3353,N_3372);
nand U3522 (N_3522,N_3300,N_3222);
nor U3523 (N_3523,N_3257,N_3363);
and U3524 (N_3524,N_3224,N_3273);
or U3525 (N_3525,N_3398,N_3280);
or U3526 (N_3526,N_3363,N_3399);
and U3527 (N_3527,N_3268,N_3335);
nand U3528 (N_3528,N_3308,N_3267);
nor U3529 (N_3529,N_3371,N_3297);
nand U3530 (N_3530,N_3369,N_3297);
or U3531 (N_3531,N_3308,N_3242);
and U3532 (N_3532,N_3201,N_3219);
or U3533 (N_3533,N_3303,N_3386);
nand U3534 (N_3534,N_3397,N_3366);
and U3535 (N_3535,N_3338,N_3269);
xnor U3536 (N_3536,N_3227,N_3220);
or U3537 (N_3537,N_3261,N_3317);
or U3538 (N_3538,N_3227,N_3206);
nand U3539 (N_3539,N_3320,N_3295);
and U3540 (N_3540,N_3276,N_3236);
or U3541 (N_3541,N_3282,N_3210);
nor U3542 (N_3542,N_3397,N_3301);
nand U3543 (N_3543,N_3230,N_3283);
or U3544 (N_3544,N_3397,N_3308);
nor U3545 (N_3545,N_3217,N_3349);
nor U3546 (N_3546,N_3245,N_3339);
nor U3547 (N_3547,N_3353,N_3236);
nand U3548 (N_3548,N_3218,N_3211);
nand U3549 (N_3549,N_3355,N_3270);
xor U3550 (N_3550,N_3334,N_3353);
and U3551 (N_3551,N_3289,N_3351);
and U3552 (N_3552,N_3384,N_3349);
or U3553 (N_3553,N_3337,N_3226);
nand U3554 (N_3554,N_3311,N_3249);
and U3555 (N_3555,N_3347,N_3342);
nand U3556 (N_3556,N_3307,N_3335);
or U3557 (N_3557,N_3384,N_3399);
and U3558 (N_3558,N_3233,N_3396);
nor U3559 (N_3559,N_3217,N_3312);
or U3560 (N_3560,N_3311,N_3213);
and U3561 (N_3561,N_3268,N_3203);
and U3562 (N_3562,N_3266,N_3347);
nor U3563 (N_3563,N_3336,N_3231);
nand U3564 (N_3564,N_3279,N_3351);
and U3565 (N_3565,N_3293,N_3357);
and U3566 (N_3566,N_3354,N_3372);
and U3567 (N_3567,N_3329,N_3381);
nand U3568 (N_3568,N_3235,N_3201);
and U3569 (N_3569,N_3267,N_3288);
nand U3570 (N_3570,N_3332,N_3394);
nor U3571 (N_3571,N_3255,N_3215);
or U3572 (N_3572,N_3224,N_3255);
or U3573 (N_3573,N_3241,N_3288);
nand U3574 (N_3574,N_3388,N_3219);
and U3575 (N_3575,N_3225,N_3277);
and U3576 (N_3576,N_3323,N_3205);
nor U3577 (N_3577,N_3233,N_3361);
nor U3578 (N_3578,N_3298,N_3201);
nand U3579 (N_3579,N_3314,N_3269);
nor U3580 (N_3580,N_3283,N_3324);
and U3581 (N_3581,N_3373,N_3283);
and U3582 (N_3582,N_3226,N_3233);
nor U3583 (N_3583,N_3327,N_3397);
and U3584 (N_3584,N_3279,N_3221);
and U3585 (N_3585,N_3277,N_3256);
nand U3586 (N_3586,N_3253,N_3338);
and U3587 (N_3587,N_3280,N_3203);
nand U3588 (N_3588,N_3222,N_3218);
nor U3589 (N_3589,N_3236,N_3376);
or U3590 (N_3590,N_3230,N_3382);
and U3591 (N_3591,N_3315,N_3203);
or U3592 (N_3592,N_3324,N_3374);
nand U3593 (N_3593,N_3278,N_3339);
and U3594 (N_3594,N_3278,N_3275);
or U3595 (N_3595,N_3294,N_3248);
nor U3596 (N_3596,N_3394,N_3364);
nor U3597 (N_3597,N_3349,N_3220);
or U3598 (N_3598,N_3233,N_3368);
and U3599 (N_3599,N_3340,N_3213);
nor U3600 (N_3600,N_3472,N_3560);
and U3601 (N_3601,N_3400,N_3407);
nor U3602 (N_3602,N_3480,N_3524);
nand U3603 (N_3603,N_3519,N_3551);
and U3604 (N_3604,N_3505,N_3457);
and U3605 (N_3605,N_3565,N_3578);
xor U3606 (N_3606,N_3464,N_3534);
and U3607 (N_3607,N_3430,N_3567);
nor U3608 (N_3608,N_3574,N_3433);
nand U3609 (N_3609,N_3585,N_3535);
nor U3610 (N_3610,N_3526,N_3413);
or U3611 (N_3611,N_3434,N_3583);
nand U3612 (N_3612,N_3414,N_3538);
and U3613 (N_3613,N_3552,N_3537);
and U3614 (N_3614,N_3426,N_3429);
and U3615 (N_3615,N_3509,N_3460);
or U3616 (N_3616,N_3401,N_3483);
or U3617 (N_3617,N_3445,N_3515);
nor U3618 (N_3618,N_3539,N_3594);
or U3619 (N_3619,N_3432,N_3488);
nor U3620 (N_3620,N_3571,N_3555);
or U3621 (N_3621,N_3529,N_3573);
and U3622 (N_3622,N_3446,N_3438);
nand U3623 (N_3623,N_3563,N_3566);
nor U3624 (N_3624,N_3531,N_3522);
nand U3625 (N_3625,N_3402,N_3506);
and U3626 (N_3626,N_3451,N_3554);
nor U3627 (N_3627,N_3495,N_3503);
nor U3628 (N_3628,N_3516,N_3454);
or U3629 (N_3629,N_3489,N_3449);
nor U3630 (N_3630,N_3553,N_3530);
or U3631 (N_3631,N_3425,N_3497);
nor U3632 (N_3632,N_3422,N_3403);
or U3633 (N_3633,N_3587,N_3410);
nand U3634 (N_3634,N_3479,N_3543);
nor U3635 (N_3635,N_3596,N_3478);
nand U3636 (N_3636,N_3588,N_3461);
nor U3637 (N_3637,N_3443,N_3517);
nand U3638 (N_3638,N_3595,N_3444);
nor U3639 (N_3639,N_3580,N_3456);
or U3640 (N_3640,N_3527,N_3424);
nand U3641 (N_3641,N_3542,N_3562);
or U3642 (N_3642,N_3484,N_3466);
and U3643 (N_3643,N_3589,N_3450);
or U3644 (N_3644,N_3540,N_3440);
or U3645 (N_3645,N_3408,N_3406);
nand U3646 (N_3646,N_3492,N_3570);
or U3647 (N_3647,N_3467,N_3452);
nand U3648 (N_3648,N_3427,N_3590);
or U3649 (N_3649,N_3547,N_3459);
nor U3650 (N_3650,N_3556,N_3511);
nor U3651 (N_3651,N_3415,N_3513);
or U3652 (N_3652,N_3514,N_3532);
nand U3653 (N_3653,N_3421,N_3441);
nand U3654 (N_3654,N_3493,N_3546);
nand U3655 (N_3655,N_3559,N_3463);
and U3656 (N_3656,N_3428,N_3496);
and U3657 (N_3657,N_3525,N_3417);
nor U3658 (N_3658,N_3557,N_3409);
xor U3659 (N_3659,N_3453,N_3584);
nand U3660 (N_3660,N_3564,N_3545);
nor U3661 (N_3661,N_3476,N_3598);
nand U3662 (N_3662,N_3419,N_3512);
or U3663 (N_3663,N_3468,N_3499);
and U3664 (N_3664,N_3416,N_3448);
or U3665 (N_3665,N_3593,N_3501);
nand U3666 (N_3666,N_3465,N_3504);
nand U3667 (N_3667,N_3458,N_3581);
nor U3668 (N_3668,N_3523,N_3412);
nand U3669 (N_3669,N_3439,N_3498);
or U3670 (N_3670,N_3521,N_3548);
or U3671 (N_3671,N_3592,N_3561);
and U3672 (N_3672,N_3591,N_3533);
nor U3673 (N_3673,N_3550,N_3490);
xnor U3674 (N_3674,N_3528,N_3405);
xor U3675 (N_3675,N_3485,N_3576);
nand U3676 (N_3676,N_3442,N_3481);
and U3677 (N_3677,N_3599,N_3502);
or U3678 (N_3678,N_3486,N_3541);
and U3679 (N_3679,N_3597,N_3586);
or U3680 (N_3680,N_3520,N_3569);
and U3681 (N_3681,N_3418,N_3558);
or U3682 (N_3682,N_3423,N_3500);
and U3683 (N_3683,N_3482,N_3568);
and U3684 (N_3684,N_3582,N_3475);
and U3685 (N_3685,N_3470,N_3404);
nand U3686 (N_3686,N_3575,N_3447);
and U3687 (N_3687,N_3469,N_3473);
xor U3688 (N_3688,N_3487,N_3431);
or U3689 (N_3689,N_3420,N_3507);
or U3690 (N_3690,N_3491,N_3544);
and U3691 (N_3691,N_3508,N_3411);
and U3692 (N_3692,N_3471,N_3536);
and U3693 (N_3693,N_3572,N_3462);
or U3694 (N_3694,N_3549,N_3577);
nor U3695 (N_3695,N_3494,N_3474);
or U3696 (N_3696,N_3435,N_3579);
nand U3697 (N_3697,N_3436,N_3455);
or U3698 (N_3698,N_3477,N_3510);
nand U3699 (N_3699,N_3437,N_3518);
or U3700 (N_3700,N_3543,N_3461);
nor U3701 (N_3701,N_3542,N_3482);
nor U3702 (N_3702,N_3518,N_3466);
or U3703 (N_3703,N_3452,N_3574);
and U3704 (N_3704,N_3554,N_3402);
nor U3705 (N_3705,N_3534,N_3589);
nand U3706 (N_3706,N_3485,N_3502);
nor U3707 (N_3707,N_3517,N_3402);
or U3708 (N_3708,N_3552,N_3524);
nor U3709 (N_3709,N_3465,N_3590);
nand U3710 (N_3710,N_3526,N_3414);
nor U3711 (N_3711,N_3451,N_3454);
nand U3712 (N_3712,N_3534,N_3505);
or U3713 (N_3713,N_3510,N_3475);
or U3714 (N_3714,N_3599,N_3469);
xor U3715 (N_3715,N_3503,N_3463);
nand U3716 (N_3716,N_3427,N_3588);
nand U3717 (N_3717,N_3584,N_3433);
or U3718 (N_3718,N_3415,N_3475);
nor U3719 (N_3719,N_3592,N_3535);
nor U3720 (N_3720,N_3574,N_3568);
nand U3721 (N_3721,N_3565,N_3522);
or U3722 (N_3722,N_3492,N_3543);
or U3723 (N_3723,N_3555,N_3553);
nand U3724 (N_3724,N_3400,N_3430);
nor U3725 (N_3725,N_3422,N_3534);
and U3726 (N_3726,N_3552,N_3443);
nor U3727 (N_3727,N_3542,N_3442);
and U3728 (N_3728,N_3561,N_3453);
nor U3729 (N_3729,N_3534,N_3591);
nand U3730 (N_3730,N_3478,N_3482);
and U3731 (N_3731,N_3565,N_3476);
nor U3732 (N_3732,N_3440,N_3576);
or U3733 (N_3733,N_3485,N_3411);
nor U3734 (N_3734,N_3445,N_3418);
nand U3735 (N_3735,N_3569,N_3595);
or U3736 (N_3736,N_3538,N_3549);
nor U3737 (N_3737,N_3413,N_3511);
and U3738 (N_3738,N_3535,N_3413);
nand U3739 (N_3739,N_3571,N_3516);
and U3740 (N_3740,N_3447,N_3513);
nor U3741 (N_3741,N_3499,N_3410);
or U3742 (N_3742,N_3415,N_3486);
and U3743 (N_3743,N_3572,N_3443);
and U3744 (N_3744,N_3576,N_3401);
nand U3745 (N_3745,N_3495,N_3558);
and U3746 (N_3746,N_3546,N_3520);
and U3747 (N_3747,N_3561,N_3490);
and U3748 (N_3748,N_3570,N_3593);
nand U3749 (N_3749,N_3452,N_3597);
nor U3750 (N_3750,N_3527,N_3449);
nor U3751 (N_3751,N_3528,N_3546);
nor U3752 (N_3752,N_3570,N_3482);
nand U3753 (N_3753,N_3402,N_3457);
nand U3754 (N_3754,N_3416,N_3422);
nand U3755 (N_3755,N_3430,N_3499);
nor U3756 (N_3756,N_3453,N_3550);
nand U3757 (N_3757,N_3562,N_3429);
or U3758 (N_3758,N_3580,N_3552);
nor U3759 (N_3759,N_3433,N_3445);
and U3760 (N_3760,N_3443,N_3582);
nor U3761 (N_3761,N_3476,N_3502);
xnor U3762 (N_3762,N_3405,N_3499);
nor U3763 (N_3763,N_3532,N_3417);
nor U3764 (N_3764,N_3464,N_3440);
and U3765 (N_3765,N_3467,N_3405);
nor U3766 (N_3766,N_3415,N_3521);
and U3767 (N_3767,N_3464,N_3406);
nand U3768 (N_3768,N_3486,N_3523);
and U3769 (N_3769,N_3430,N_3493);
nor U3770 (N_3770,N_3418,N_3469);
nand U3771 (N_3771,N_3513,N_3542);
and U3772 (N_3772,N_3489,N_3569);
or U3773 (N_3773,N_3420,N_3485);
nand U3774 (N_3774,N_3512,N_3506);
and U3775 (N_3775,N_3428,N_3592);
xnor U3776 (N_3776,N_3480,N_3435);
or U3777 (N_3777,N_3534,N_3521);
and U3778 (N_3778,N_3514,N_3414);
nor U3779 (N_3779,N_3545,N_3400);
and U3780 (N_3780,N_3573,N_3497);
or U3781 (N_3781,N_3403,N_3417);
nor U3782 (N_3782,N_3467,N_3565);
nand U3783 (N_3783,N_3501,N_3507);
nor U3784 (N_3784,N_3476,N_3516);
or U3785 (N_3785,N_3426,N_3436);
nor U3786 (N_3786,N_3533,N_3493);
and U3787 (N_3787,N_3472,N_3496);
or U3788 (N_3788,N_3474,N_3469);
nor U3789 (N_3789,N_3596,N_3525);
or U3790 (N_3790,N_3532,N_3491);
nor U3791 (N_3791,N_3452,N_3466);
and U3792 (N_3792,N_3468,N_3508);
and U3793 (N_3793,N_3457,N_3409);
nor U3794 (N_3794,N_3526,N_3424);
and U3795 (N_3795,N_3591,N_3455);
and U3796 (N_3796,N_3492,N_3574);
and U3797 (N_3797,N_3592,N_3556);
nor U3798 (N_3798,N_3517,N_3492);
nor U3799 (N_3799,N_3492,N_3406);
nor U3800 (N_3800,N_3726,N_3755);
nand U3801 (N_3801,N_3754,N_3714);
or U3802 (N_3802,N_3627,N_3760);
nand U3803 (N_3803,N_3635,N_3766);
or U3804 (N_3804,N_3630,N_3641);
nor U3805 (N_3805,N_3618,N_3672);
or U3806 (N_3806,N_3620,N_3600);
and U3807 (N_3807,N_3614,N_3772);
and U3808 (N_3808,N_3684,N_3659);
nand U3809 (N_3809,N_3791,N_3685);
nand U3810 (N_3810,N_3767,N_3645);
or U3811 (N_3811,N_3724,N_3773);
nand U3812 (N_3812,N_3699,N_3650);
nor U3813 (N_3813,N_3710,N_3715);
and U3814 (N_3814,N_3761,N_3654);
nand U3815 (N_3815,N_3794,N_3636);
and U3816 (N_3816,N_3688,N_3697);
or U3817 (N_3817,N_3705,N_3756);
nor U3818 (N_3818,N_3664,N_3666);
or U3819 (N_3819,N_3739,N_3712);
and U3820 (N_3820,N_3663,N_3677);
and U3821 (N_3821,N_3602,N_3747);
nor U3822 (N_3822,N_3655,N_3771);
and U3823 (N_3823,N_3787,N_3703);
nor U3824 (N_3824,N_3694,N_3701);
or U3825 (N_3825,N_3607,N_3689);
nor U3826 (N_3826,N_3695,N_3736);
nor U3827 (N_3827,N_3617,N_3613);
nand U3828 (N_3828,N_3683,N_3652);
nor U3829 (N_3829,N_3751,N_3783);
nor U3830 (N_3830,N_3745,N_3661);
nand U3831 (N_3831,N_3622,N_3723);
or U3832 (N_3832,N_3644,N_3716);
nor U3833 (N_3833,N_3642,N_3665);
nor U3834 (N_3834,N_3782,N_3660);
nand U3835 (N_3835,N_3759,N_3728);
or U3836 (N_3836,N_3744,N_3657);
nor U3837 (N_3837,N_3615,N_3608);
or U3838 (N_3838,N_3698,N_3626);
and U3839 (N_3839,N_3696,N_3798);
nor U3840 (N_3840,N_3648,N_3770);
or U3841 (N_3841,N_3776,N_3680);
and U3842 (N_3842,N_3729,N_3621);
nor U3843 (N_3843,N_3633,N_3675);
xor U3844 (N_3844,N_3757,N_3708);
and U3845 (N_3845,N_3640,N_3796);
nand U3846 (N_3846,N_3670,N_3681);
xor U3847 (N_3847,N_3780,N_3673);
nand U3848 (N_3848,N_3691,N_3738);
or U3849 (N_3849,N_3769,N_3762);
or U3850 (N_3850,N_3741,N_3734);
nand U3851 (N_3851,N_3662,N_3788);
nor U3852 (N_3852,N_3758,N_3679);
and U3853 (N_3853,N_3721,N_3669);
nand U3854 (N_3854,N_3727,N_3704);
nand U3855 (N_3855,N_3667,N_3611);
or U3856 (N_3856,N_3651,N_3735);
nand U3857 (N_3857,N_3737,N_3601);
and U3858 (N_3858,N_3763,N_3775);
or U3859 (N_3859,N_3732,N_3687);
and U3860 (N_3860,N_3717,N_3746);
nor U3861 (N_3861,N_3619,N_3718);
nand U3862 (N_3862,N_3742,N_3616);
nand U3863 (N_3863,N_3658,N_3764);
and U3864 (N_3864,N_3623,N_3790);
and U3865 (N_3865,N_3631,N_3674);
or U3866 (N_3866,N_3682,N_3647);
or U3867 (N_3867,N_3693,N_3656);
nor U3868 (N_3868,N_3639,N_3785);
or U3869 (N_3869,N_3711,N_3653);
or U3870 (N_3870,N_3743,N_3690);
or U3871 (N_3871,N_3678,N_3638);
and U3872 (N_3872,N_3713,N_3792);
and U3873 (N_3873,N_3748,N_3720);
nor U3874 (N_3874,N_3649,N_3668);
nand U3875 (N_3875,N_3702,N_3730);
nand U3876 (N_3876,N_3786,N_3646);
nand U3877 (N_3877,N_3604,N_3753);
and U3878 (N_3878,N_3700,N_3676);
and U3879 (N_3879,N_3609,N_3795);
or U3880 (N_3880,N_3628,N_3797);
nor U3881 (N_3881,N_3612,N_3793);
nor U3882 (N_3882,N_3784,N_3686);
and U3883 (N_3883,N_3603,N_3765);
and U3884 (N_3884,N_3692,N_3752);
or U3885 (N_3885,N_3707,N_3789);
or U3886 (N_3886,N_3606,N_3733);
nand U3887 (N_3887,N_3774,N_3750);
nand U3888 (N_3888,N_3643,N_3719);
or U3889 (N_3889,N_3610,N_3706);
or U3890 (N_3890,N_3632,N_3778);
and U3891 (N_3891,N_3709,N_3671);
nor U3892 (N_3892,N_3725,N_3624);
nand U3893 (N_3893,N_3634,N_3779);
nand U3894 (N_3894,N_3740,N_3781);
or U3895 (N_3895,N_3637,N_3731);
and U3896 (N_3896,N_3799,N_3749);
or U3897 (N_3897,N_3768,N_3625);
and U3898 (N_3898,N_3605,N_3629);
and U3899 (N_3899,N_3777,N_3722);
nor U3900 (N_3900,N_3731,N_3609);
or U3901 (N_3901,N_3669,N_3679);
nor U3902 (N_3902,N_3721,N_3760);
and U3903 (N_3903,N_3798,N_3709);
nor U3904 (N_3904,N_3721,N_3774);
or U3905 (N_3905,N_3604,N_3672);
nand U3906 (N_3906,N_3621,N_3742);
nor U3907 (N_3907,N_3775,N_3609);
and U3908 (N_3908,N_3636,N_3666);
nor U3909 (N_3909,N_3604,N_3619);
or U3910 (N_3910,N_3650,N_3734);
and U3911 (N_3911,N_3644,N_3645);
nor U3912 (N_3912,N_3787,N_3760);
nand U3913 (N_3913,N_3630,N_3734);
nor U3914 (N_3914,N_3605,N_3624);
nor U3915 (N_3915,N_3707,N_3608);
xnor U3916 (N_3916,N_3676,N_3648);
and U3917 (N_3917,N_3755,N_3738);
nand U3918 (N_3918,N_3747,N_3621);
and U3919 (N_3919,N_3673,N_3665);
and U3920 (N_3920,N_3794,N_3659);
nand U3921 (N_3921,N_3753,N_3732);
nor U3922 (N_3922,N_3769,N_3697);
nor U3923 (N_3923,N_3758,N_3740);
nor U3924 (N_3924,N_3793,N_3696);
nor U3925 (N_3925,N_3719,N_3757);
nor U3926 (N_3926,N_3674,N_3602);
nor U3927 (N_3927,N_3643,N_3731);
xnor U3928 (N_3928,N_3718,N_3672);
or U3929 (N_3929,N_3706,N_3696);
nor U3930 (N_3930,N_3733,N_3699);
nor U3931 (N_3931,N_3798,N_3757);
nor U3932 (N_3932,N_3628,N_3783);
and U3933 (N_3933,N_3730,N_3621);
and U3934 (N_3934,N_3798,N_3610);
or U3935 (N_3935,N_3779,N_3784);
xor U3936 (N_3936,N_3662,N_3794);
nand U3937 (N_3937,N_3624,N_3739);
or U3938 (N_3938,N_3605,N_3721);
nand U3939 (N_3939,N_3620,N_3712);
and U3940 (N_3940,N_3615,N_3765);
nand U3941 (N_3941,N_3776,N_3769);
nor U3942 (N_3942,N_3622,N_3707);
nor U3943 (N_3943,N_3746,N_3754);
or U3944 (N_3944,N_3649,N_3718);
nand U3945 (N_3945,N_3763,N_3787);
and U3946 (N_3946,N_3742,N_3796);
or U3947 (N_3947,N_3682,N_3770);
nand U3948 (N_3948,N_3770,N_3756);
or U3949 (N_3949,N_3613,N_3603);
nor U3950 (N_3950,N_3696,N_3618);
or U3951 (N_3951,N_3783,N_3763);
or U3952 (N_3952,N_3674,N_3736);
and U3953 (N_3953,N_3756,N_3667);
or U3954 (N_3954,N_3618,N_3747);
nor U3955 (N_3955,N_3638,N_3747);
nand U3956 (N_3956,N_3778,N_3723);
or U3957 (N_3957,N_3675,N_3767);
nor U3958 (N_3958,N_3735,N_3619);
and U3959 (N_3959,N_3753,N_3751);
or U3960 (N_3960,N_3642,N_3732);
nor U3961 (N_3961,N_3640,N_3759);
xnor U3962 (N_3962,N_3778,N_3732);
or U3963 (N_3963,N_3743,N_3691);
xnor U3964 (N_3964,N_3661,N_3699);
and U3965 (N_3965,N_3679,N_3789);
or U3966 (N_3966,N_3710,N_3638);
or U3967 (N_3967,N_3723,N_3631);
and U3968 (N_3968,N_3772,N_3619);
or U3969 (N_3969,N_3779,N_3662);
and U3970 (N_3970,N_3738,N_3687);
nand U3971 (N_3971,N_3763,N_3699);
nor U3972 (N_3972,N_3617,N_3668);
nor U3973 (N_3973,N_3636,N_3661);
nand U3974 (N_3974,N_3632,N_3665);
or U3975 (N_3975,N_3663,N_3644);
and U3976 (N_3976,N_3640,N_3647);
nand U3977 (N_3977,N_3640,N_3779);
nand U3978 (N_3978,N_3706,N_3674);
nor U3979 (N_3979,N_3739,N_3628);
and U3980 (N_3980,N_3693,N_3611);
and U3981 (N_3981,N_3703,N_3796);
or U3982 (N_3982,N_3689,N_3718);
or U3983 (N_3983,N_3732,N_3747);
nand U3984 (N_3984,N_3603,N_3650);
nor U3985 (N_3985,N_3690,N_3723);
nor U3986 (N_3986,N_3716,N_3623);
and U3987 (N_3987,N_3775,N_3669);
or U3988 (N_3988,N_3746,N_3771);
and U3989 (N_3989,N_3747,N_3616);
or U3990 (N_3990,N_3615,N_3711);
nand U3991 (N_3991,N_3702,N_3744);
nor U3992 (N_3992,N_3658,N_3630);
xnor U3993 (N_3993,N_3777,N_3604);
nand U3994 (N_3994,N_3717,N_3680);
nand U3995 (N_3995,N_3607,N_3662);
and U3996 (N_3996,N_3655,N_3671);
nor U3997 (N_3997,N_3744,N_3728);
and U3998 (N_3998,N_3688,N_3612);
or U3999 (N_3999,N_3654,N_3717);
or U4000 (N_4000,N_3826,N_3800);
nand U4001 (N_4001,N_3926,N_3861);
or U4002 (N_4002,N_3879,N_3875);
xnor U4003 (N_4003,N_3894,N_3930);
and U4004 (N_4004,N_3971,N_3811);
and U4005 (N_4005,N_3899,N_3805);
nand U4006 (N_4006,N_3977,N_3972);
nand U4007 (N_4007,N_3865,N_3927);
nor U4008 (N_4008,N_3802,N_3891);
nor U4009 (N_4009,N_3887,N_3834);
or U4010 (N_4010,N_3939,N_3911);
xnor U4011 (N_4011,N_3829,N_3849);
nor U4012 (N_4012,N_3856,N_3823);
nand U4013 (N_4013,N_3886,N_3965);
or U4014 (N_4014,N_3953,N_3909);
nand U4015 (N_4015,N_3801,N_3825);
nand U4016 (N_4016,N_3866,N_3841);
nor U4017 (N_4017,N_3985,N_3868);
nand U4018 (N_4018,N_3978,N_3846);
nor U4019 (N_4019,N_3905,N_3980);
nor U4020 (N_4020,N_3947,N_3827);
and U4021 (N_4021,N_3843,N_3943);
xnor U4022 (N_4022,N_3888,N_3983);
and U4023 (N_4023,N_3924,N_3874);
nand U4024 (N_4024,N_3839,N_3913);
nand U4025 (N_4025,N_3916,N_3844);
and U4026 (N_4026,N_3822,N_3995);
and U4027 (N_4027,N_3976,N_3878);
or U4028 (N_4028,N_3950,N_3949);
and U4029 (N_4029,N_3803,N_3842);
and U4030 (N_4030,N_3944,N_3966);
nor U4031 (N_4031,N_3994,N_3959);
and U4032 (N_4032,N_3836,N_3982);
nor U4033 (N_4033,N_3937,N_3857);
xnor U4034 (N_4034,N_3986,N_3948);
nor U4035 (N_4035,N_3897,N_3883);
or U4036 (N_4036,N_3923,N_3901);
or U4037 (N_4037,N_3915,N_3808);
and U4038 (N_4038,N_3970,N_3830);
and U4039 (N_4039,N_3845,N_3997);
nand U4040 (N_4040,N_3946,N_3867);
nor U4041 (N_4041,N_3906,N_3954);
nor U4042 (N_4042,N_3962,N_3912);
or U4043 (N_4043,N_3813,N_3896);
nand U4044 (N_4044,N_3872,N_3871);
and U4045 (N_4045,N_3991,N_3963);
xnor U4046 (N_4046,N_3812,N_3952);
or U4047 (N_4047,N_3884,N_3989);
nand U4048 (N_4048,N_3885,N_3824);
nor U4049 (N_4049,N_3935,N_3993);
nand U4050 (N_4050,N_3847,N_3904);
nand U4051 (N_4051,N_3804,N_3893);
nor U4052 (N_4052,N_3838,N_3869);
nor U4053 (N_4053,N_3929,N_3955);
and U4054 (N_4054,N_3870,N_3903);
and U4055 (N_4055,N_3992,N_3945);
nor U4056 (N_4056,N_3908,N_3851);
or U4057 (N_4057,N_3999,N_3876);
nand U4058 (N_4058,N_3968,N_3974);
or U4059 (N_4059,N_3925,N_3892);
and U4060 (N_4060,N_3837,N_3815);
nand U4061 (N_4061,N_3817,N_3979);
and U4062 (N_4062,N_3806,N_3910);
or U4063 (N_4063,N_3919,N_3855);
and U4064 (N_4064,N_3932,N_3964);
nand U4065 (N_4065,N_3996,N_3864);
or U4066 (N_4066,N_3940,N_3957);
nor U4067 (N_4067,N_3900,N_3918);
xor U4068 (N_4068,N_3928,N_3831);
nor U4069 (N_4069,N_3975,N_3895);
and U4070 (N_4070,N_3934,N_3863);
nand U4071 (N_4071,N_3941,N_3858);
and U4072 (N_4072,N_3898,N_3942);
nor U4073 (N_4073,N_3960,N_3832);
or U4074 (N_4074,N_3920,N_3853);
nand U4075 (N_4075,N_3973,N_3987);
or U4076 (N_4076,N_3914,N_3961);
and U4077 (N_4077,N_3833,N_3807);
and U4078 (N_4078,N_3810,N_3933);
nand U4079 (N_4079,N_3998,N_3984);
or U4080 (N_4080,N_3819,N_3862);
nand U4081 (N_4081,N_3835,N_3967);
nor U4082 (N_4082,N_3848,N_3936);
nand U4083 (N_4083,N_3818,N_3859);
nand U4084 (N_4084,N_3956,N_3881);
nor U4085 (N_4085,N_3981,N_3990);
nor U4086 (N_4086,N_3921,N_3890);
nor U4087 (N_4087,N_3809,N_3922);
nand U4088 (N_4088,N_3820,N_3907);
nor U4089 (N_4089,N_3814,N_3882);
nor U4090 (N_4090,N_3902,N_3880);
or U4091 (N_4091,N_3938,N_3958);
nand U4092 (N_4092,N_3873,N_3850);
nand U4093 (N_4093,N_3816,N_3840);
nand U4094 (N_4094,N_3860,N_3854);
nor U4095 (N_4095,N_3931,N_3821);
nand U4096 (N_4096,N_3988,N_3889);
nor U4097 (N_4097,N_3917,N_3852);
and U4098 (N_4098,N_3877,N_3828);
nor U4099 (N_4099,N_3951,N_3969);
or U4100 (N_4100,N_3871,N_3833);
or U4101 (N_4101,N_3866,N_3937);
or U4102 (N_4102,N_3948,N_3949);
nor U4103 (N_4103,N_3831,N_3930);
and U4104 (N_4104,N_3878,N_3978);
nand U4105 (N_4105,N_3951,N_3950);
and U4106 (N_4106,N_3987,N_3892);
nand U4107 (N_4107,N_3966,N_3846);
nand U4108 (N_4108,N_3957,N_3885);
or U4109 (N_4109,N_3880,N_3940);
or U4110 (N_4110,N_3814,N_3991);
nor U4111 (N_4111,N_3845,N_3911);
nand U4112 (N_4112,N_3974,N_3843);
or U4113 (N_4113,N_3811,N_3972);
or U4114 (N_4114,N_3801,N_3972);
nor U4115 (N_4115,N_3927,N_3856);
nand U4116 (N_4116,N_3987,N_3847);
and U4117 (N_4117,N_3921,N_3903);
and U4118 (N_4118,N_3885,N_3919);
xnor U4119 (N_4119,N_3921,N_3993);
and U4120 (N_4120,N_3915,N_3975);
and U4121 (N_4121,N_3867,N_3938);
nor U4122 (N_4122,N_3934,N_3980);
nor U4123 (N_4123,N_3863,N_3937);
and U4124 (N_4124,N_3970,N_3945);
nor U4125 (N_4125,N_3824,N_3853);
and U4126 (N_4126,N_3829,N_3975);
or U4127 (N_4127,N_3992,N_3820);
and U4128 (N_4128,N_3837,N_3816);
nand U4129 (N_4129,N_3954,N_3935);
xnor U4130 (N_4130,N_3961,N_3870);
nor U4131 (N_4131,N_3862,N_3944);
nand U4132 (N_4132,N_3925,N_3806);
and U4133 (N_4133,N_3905,N_3928);
nand U4134 (N_4134,N_3977,N_3837);
or U4135 (N_4135,N_3989,N_3853);
nor U4136 (N_4136,N_3807,N_3835);
nor U4137 (N_4137,N_3951,N_3885);
or U4138 (N_4138,N_3815,N_3852);
nor U4139 (N_4139,N_3965,N_3988);
and U4140 (N_4140,N_3938,N_3922);
nor U4141 (N_4141,N_3929,N_3918);
and U4142 (N_4142,N_3930,N_3875);
nor U4143 (N_4143,N_3978,N_3984);
or U4144 (N_4144,N_3850,N_3870);
and U4145 (N_4145,N_3995,N_3997);
nor U4146 (N_4146,N_3863,N_3899);
and U4147 (N_4147,N_3996,N_3894);
nand U4148 (N_4148,N_3806,N_3805);
or U4149 (N_4149,N_3842,N_3982);
xnor U4150 (N_4150,N_3949,N_3971);
nor U4151 (N_4151,N_3869,N_3870);
and U4152 (N_4152,N_3916,N_3974);
or U4153 (N_4153,N_3874,N_3981);
and U4154 (N_4154,N_3965,N_3838);
and U4155 (N_4155,N_3971,N_3970);
or U4156 (N_4156,N_3993,N_3958);
and U4157 (N_4157,N_3854,N_3909);
and U4158 (N_4158,N_3877,N_3896);
and U4159 (N_4159,N_3938,N_3832);
or U4160 (N_4160,N_3801,N_3887);
nand U4161 (N_4161,N_3935,N_3927);
nor U4162 (N_4162,N_3883,N_3862);
or U4163 (N_4163,N_3929,N_3911);
xnor U4164 (N_4164,N_3932,N_3907);
or U4165 (N_4165,N_3816,N_3982);
nand U4166 (N_4166,N_3846,N_3893);
nor U4167 (N_4167,N_3967,N_3958);
nor U4168 (N_4168,N_3886,N_3945);
and U4169 (N_4169,N_3910,N_3912);
or U4170 (N_4170,N_3881,N_3937);
xnor U4171 (N_4171,N_3878,N_3995);
nand U4172 (N_4172,N_3821,N_3841);
nand U4173 (N_4173,N_3961,N_3834);
nand U4174 (N_4174,N_3973,N_3896);
xor U4175 (N_4175,N_3871,N_3838);
or U4176 (N_4176,N_3920,N_3942);
nor U4177 (N_4177,N_3815,N_3888);
or U4178 (N_4178,N_3970,N_3882);
or U4179 (N_4179,N_3856,N_3996);
nor U4180 (N_4180,N_3831,N_3841);
or U4181 (N_4181,N_3870,N_3892);
nor U4182 (N_4182,N_3956,N_3948);
or U4183 (N_4183,N_3829,N_3901);
nand U4184 (N_4184,N_3838,N_3981);
nand U4185 (N_4185,N_3993,N_3946);
or U4186 (N_4186,N_3862,N_3927);
and U4187 (N_4187,N_3989,N_3933);
and U4188 (N_4188,N_3853,N_3857);
or U4189 (N_4189,N_3882,N_3896);
nand U4190 (N_4190,N_3914,N_3871);
nor U4191 (N_4191,N_3956,N_3846);
or U4192 (N_4192,N_3981,N_3835);
nor U4193 (N_4193,N_3883,N_3980);
nor U4194 (N_4194,N_3845,N_3915);
nand U4195 (N_4195,N_3818,N_3929);
and U4196 (N_4196,N_3892,N_3939);
nor U4197 (N_4197,N_3941,N_3992);
nor U4198 (N_4198,N_3909,N_3959);
and U4199 (N_4199,N_3897,N_3968);
or U4200 (N_4200,N_4117,N_4066);
nand U4201 (N_4201,N_4065,N_4026);
or U4202 (N_4202,N_4009,N_4159);
nor U4203 (N_4203,N_4136,N_4070);
nor U4204 (N_4204,N_4000,N_4190);
and U4205 (N_4205,N_4006,N_4074);
or U4206 (N_4206,N_4012,N_4067);
nor U4207 (N_4207,N_4104,N_4027);
and U4208 (N_4208,N_4036,N_4050);
or U4209 (N_4209,N_4124,N_4030);
or U4210 (N_4210,N_4018,N_4024);
nor U4211 (N_4211,N_4048,N_4084);
nand U4212 (N_4212,N_4062,N_4192);
or U4213 (N_4213,N_4183,N_4075);
nor U4214 (N_4214,N_4063,N_4138);
or U4215 (N_4215,N_4102,N_4080);
nand U4216 (N_4216,N_4165,N_4002);
and U4217 (N_4217,N_4088,N_4029);
or U4218 (N_4218,N_4035,N_4185);
nor U4219 (N_4219,N_4119,N_4096);
nor U4220 (N_4220,N_4121,N_4073);
nand U4221 (N_4221,N_4013,N_4044);
nor U4222 (N_4222,N_4139,N_4197);
and U4223 (N_4223,N_4010,N_4167);
or U4224 (N_4224,N_4163,N_4191);
nand U4225 (N_4225,N_4146,N_4015);
nand U4226 (N_4226,N_4155,N_4169);
nand U4227 (N_4227,N_4064,N_4153);
or U4228 (N_4228,N_4130,N_4069);
or U4229 (N_4229,N_4184,N_4058);
nor U4230 (N_4230,N_4051,N_4175);
or U4231 (N_4231,N_4160,N_4128);
nand U4232 (N_4232,N_4008,N_4193);
nand U4233 (N_4233,N_4157,N_4123);
nor U4234 (N_4234,N_4152,N_4077);
or U4235 (N_4235,N_4118,N_4017);
nor U4236 (N_4236,N_4034,N_4108);
nor U4237 (N_4237,N_4100,N_4105);
or U4238 (N_4238,N_4007,N_4141);
or U4239 (N_4239,N_4156,N_4187);
xnor U4240 (N_4240,N_4154,N_4039);
nand U4241 (N_4241,N_4173,N_4148);
nor U4242 (N_4242,N_4151,N_4086);
nor U4243 (N_4243,N_4122,N_4093);
or U4244 (N_4244,N_4092,N_4042);
and U4245 (N_4245,N_4149,N_4004);
or U4246 (N_4246,N_4171,N_4049);
or U4247 (N_4247,N_4003,N_4112);
nor U4248 (N_4248,N_4032,N_4145);
or U4249 (N_4249,N_4106,N_4158);
nand U4250 (N_4250,N_4179,N_4177);
and U4251 (N_4251,N_4110,N_4166);
nor U4252 (N_4252,N_4113,N_4014);
and U4253 (N_4253,N_4025,N_4043);
nand U4254 (N_4254,N_4164,N_4054);
or U4255 (N_4255,N_4144,N_4188);
nor U4256 (N_4256,N_4055,N_4140);
nor U4257 (N_4257,N_4031,N_4134);
nand U4258 (N_4258,N_4083,N_4198);
nor U4259 (N_4259,N_4143,N_4133);
nand U4260 (N_4260,N_4182,N_4150);
nor U4261 (N_4261,N_4016,N_4061);
nor U4262 (N_4262,N_4071,N_4126);
nor U4263 (N_4263,N_4085,N_4115);
and U4264 (N_4264,N_4195,N_4095);
or U4265 (N_4265,N_4019,N_4181);
nor U4266 (N_4266,N_4120,N_4132);
and U4267 (N_4267,N_4020,N_4101);
nor U4268 (N_4268,N_4028,N_4094);
nand U4269 (N_4269,N_4011,N_4194);
and U4270 (N_4270,N_4052,N_4131);
and U4271 (N_4271,N_4125,N_4098);
or U4272 (N_4272,N_4076,N_4103);
or U4273 (N_4273,N_4053,N_4135);
or U4274 (N_4274,N_4023,N_4041);
xor U4275 (N_4275,N_4089,N_4176);
xnor U4276 (N_4276,N_4059,N_4081);
nor U4277 (N_4277,N_4005,N_4037);
and U4278 (N_4278,N_4142,N_4090);
or U4279 (N_4279,N_4199,N_4091);
and U4280 (N_4280,N_4174,N_4180);
and U4281 (N_4281,N_4022,N_4046);
or U4282 (N_4282,N_4072,N_4178);
or U4283 (N_4283,N_4056,N_4196);
nand U4284 (N_4284,N_4001,N_4060);
nor U4285 (N_4285,N_4172,N_4161);
nor U4286 (N_4286,N_4082,N_4078);
or U4287 (N_4287,N_4057,N_4033);
nand U4288 (N_4288,N_4047,N_4109);
nor U4289 (N_4289,N_4038,N_4111);
nand U4290 (N_4290,N_4189,N_4147);
xor U4291 (N_4291,N_4045,N_4170);
or U4292 (N_4292,N_4168,N_4068);
nor U4293 (N_4293,N_4079,N_4099);
or U4294 (N_4294,N_4127,N_4107);
nor U4295 (N_4295,N_4186,N_4087);
nor U4296 (N_4296,N_4114,N_4021);
and U4297 (N_4297,N_4129,N_4097);
or U4298 (N_4298,N_4162,N_4040);
or U4299 (N_4299,N_4137,N_4116);
and U4300 (N_4300,N_4056,N_4197);
and U4301 (N_4301,N_4153,N_4120);
nor U4302 (N_4302,N_4049,N_4108);
nor U4303 (N_4303,N_4171,N_4120);
or U4304 (N_4304,N_4098,N_4036);
and U4305 (N_4305,N_4022,N_4126);
nand U4306 (N_4306,N_4102,N_4029);
and U4307 (N_4307,N_4170,N_4101);
nor U4308 (N_4308,N_4131,N_4105);
nor U4309 (N_4309,N_4043,N_4119);
nor U4310 (N_4310,N_4059,N_4006);
nand U4311 (N_4311,N_4030,N_4111);
nand U4312 (N_4312,N_4059,N_4129);
or U4313 (N_4313,N_4013,N_4194);
nor U4314 (N_4314,N_4106,N_4189);
or U4315 (N_4315,N_4187,N_4157);
and U4316 (N_4316,N_4020,N_4021);
nand U4317 (N_4317,N_4162,N_4126);
and U4318 (N_4318,N_4173,N_4134);
or U4319 (N_4319,N_4116,N_4143);
nor U4320 (N_4320,N_4061,N_4010);
nor U4321 (N_4321,N_4071,N_4149);
and U4322 (N_4322,N_4105,N_4058);
and U4323 (N_4323,N_4057,N_4059);
nor U4324 (N_4324,N_4136,N_4187);
nand U4325 (N_4325,N_4090,N_4028);
nand U4326 (N_4326,N_4162,N_4191);
and U4327 (N_4327,N_4013,N_4186);
or U4328 (N_4328,N_4050,N_4117);
or U4329 (N_4329,N_4167,N_4067);
nor U4330 (N_4330,N_4089,N_4062);
or U4331 (N_4331,N_4002,N_4038);
nor U4332 (N_4332,N_4138,N_4072);
or U4333 (N_4333,N_4080,N_4130);
and U4334 (N_4334,N_4164,N_4015);
and U4335 (N_4335,N_4137,N_4019);
nand U4336 (N_4336,N_4182,N_4089);
nand U4337 (N_4337,N_4079,N_4035);
nand U4338 (N_4338,N_4016,N_4024);
and U4339 (N_4339,N_4169,N_4043);
nand U4340 (N_4340,N_4118,N_4158);
nor U4341 (N_4341,N_4157,N_4120);
and U4342 (N_4342,N_4100,N_4189);
and U4343 (N_4343,N_4052,N_4085);
or U4344 (N_4344,N_4079,N_4033);
or U4345 (N_4345,N_4155,N_4064);
xnor U4346 (N_4346,N_4120,N_4129);
or U4347 (N_4347,N_4011,N_4136);
nand U4348 (N_4348,N_4188,N_4149);
and U4349 (N_4349,N_4080,N_4002);
nor U4350 (N_4350,N_4144,N_4050);
or U4351 (N_4351,N_4107,N_4158);
nor U4352 (N_4352,N_4074,N_4127);
or U4353 (N_4353,N_4081,N_4010);
xnor U4354 (N_4354,N_4032,N_4101);
and U4355 (N_4355,N_4184,N_4094);
and U4356 (N_4356,N_4102,N_4085);
nand U4357 (N_4357,N_4051,N_4136);
nand U4358 (N_4358,N_4054,N_4063);
or U4359 (N_4359,N_4071,N_4103);
and U4360 (N_4360,N_4040,N_4191);
nand U4361 (N_4361,N_4157,N_4034);
nand U4362 (N_4362,N_4024,N_4128);
xnor U4363 (N_4363,N_4026,N_4050);
or U4364 (N_4364,N_4006,N_4121);
nand U4365 (N_4365,N_4179,N_4105);
or U4366 (N_4366,N_4116,N_4088);
nand U4367 (N_4367,N_4116,N_4002);
nor U4368 (N_4368,N_4026,N_4119);
or U4369 (N_4369,N_4090,N_4098);
or U4370 (N_4370,N_4026,N_4081);
and U4371 (N_4371,N_4156,N_4009);
nand U4372 (N_4372,N_4138,N_4043);
or U4373 (N_4373,N_4183,N_4014);
nor U4374 (N_4374,N_4048,N_4116);
nor U4375 (N_4375,N_4011,N_4181);
or U4376 (N_4376,N_4042,N_4189);
or U4377 (N_4377,N_4076,N_4011);
nor U4378 (N_4378,N_4063,N_4062);
and U4379 (N_4379,N_4004,N_4028);
and U4380 (N_4380,N_4196,N_4130);
nand U4381 (N_4381,N_4178,N_4017);
and U4382 (N_4382,N_4179,N_4121);
nor U4383 (N_4383,N_4039,N_4057);
or U4384 (N_4384,N_4054,N_4027);
nor U4385 (N_4385,N_4026,N_4108);
nor U4386 (N_4386,N_4051,N_4188);
and U4387 (N_4387,N_4177,N_4060);
and U4388 (N_4388,N_4044,N_4114);
and U4389 (N_4389,N_4033,N_4114);
and U4390 (N_4390,N_4131,N_4081);
nor U4391 (N_4391,N_4181,N_4040);
and U4392 (N_4392,N_4081,N_4138);
or U4393 (N_4393,N_4014,N_4081);
or U4394 (N_4394,N_4069,N_4067);
nor U4395 (N_4395,N_4039,N_4032);
and U4396 (N_4396,N_4181,N_4026);
and U4397 (N_4397,N_4125,N_4063);
nor U4398 (N_4398,N_4017,N_4195);
nand U4399 (N_4399,N_4167,N_4068);
nand U4400 (N_4400,N_4247,N_4203);
nand U4401 (N_4401,N_4322,N_4268);
or U4402 (N_4402,N_4398,N_4227);
nor U4403 (N_4403,N_4257,N_4218);
nor U4404 (N_4404,N_4321,N_4201);
nor U4405 (N_4405,N_4380,N_4371);
and U4406 (N_4406,N_4339,N_4252);
or U4407 (N_4407,N_4200,N_4245);
and U4408 (N_4408,N_4210,N_4279);
nor U4409 (N_4409,N_4397,N_4246);
and U4410 (N_4410,N_4277,N_4358);
or U4411 (N_4411,N_4365,N_4242);
nor U4412 (N_4412,N_4293,N_4265);
or U4413 (N_4413,N_4312,N_4359);
and U4414 (N_4414,N_4328,N_4318);
nand U4415 (N_4415,N_4348,N_4212);
nor U4416 (N_4416,N_4248,N_4335);
nor U4417 (N_4417,N_4372,N_4391);
and U4418 (N_4418,N_4327,N_4229);
nor U4419 (N_4419,N_4346,N_4396);
or U4420 (N_4420,N_4206,N_4352);
or U4421 (N_4421,N_4336,N_4308);
nor U4422 (N_4422,N_4375,N_4357);
and U4423 (N_4423,N_4211,N_4319);
nand U4424 (N_4424,N_4306,N_4337);
nor U4425 (N_4425,N_4216,N_4385);
xor U4426 (N_4426,N_4373,N_4250);
and U4427 (N_4427,N_4368,N_4350);
nand U4428 (N_4428,N_4297,N_4292);
nand U4429 (N_4429,N_4342,N_4302);
and U4430 (N_4430,N_4361,N_4378);
and U4431 (N_4431,N_4228,N_4287);
xnor U4432 (N_4432,N_4225,N_4264);
nand U4433 (N_4433,N_4231,N_4275);
nor U4434 (N_4434,N_4299,N_4366);
nor U4435 (N_4435,N_4387,N_4219);
and U4436 (N_4436,N_4209,N_4217);
or U4437 (N_4437,N_4353,N_4333);
and U4438 (N_4438,N_4345,N_4395);
nor U4439 (N_4439,N_4389,N_4370);
and U4440 (N_4440,N_4239,N_4280);
or U4441 (N_4441,N_4313,N_4222);
xnor U4442 (N_4442,N_4258,N_4213);
nand U4443 (N_4443,N_4354,N_4224);
and U4444 (N_4444,N_4295,N_4338);
or U4445 (N_4445,N_4305,N_4329);
and U4446 (N_4446,N_4236,N_4301);
nor U4447 (N_4447,N_4273,N_4238);
and U4448 (N_4448,N_4267,N_4331);
and U4449 (N_4449,N_4261,N_4324);
or U4450 (N_4450,N_4388,N_4220);
or U4451 (N_4451,N_4215,N_4332);
nand U4452 (N_4452,N_4296,N_4379);
and U4453 (N_4453,N_4356,N_4382);
nand U4454 (N_4454,N_4294,N_4347);
and U4455 (N_4455,N_4386,N_4362);
or U4456 (N_4456,N_4369,N_4309);
nor U4457 (N_4457,N_4237,N_4226);
nand U4458 (N_4458,N_4235,N_4316);
or U4459 (N_4459,N_4255,N_4343);
xnor U4460 (N_4460,N_4286,N_4340);
or U4461 (N_4461,N_4284,N_4221);
nand U4462 (N_4462,N_4288,N_4240);
nand U4463 (N_4463,N_4314,N_4317);
and U4464 (N_4464,N_4307,N_4344);
nor U4465 (N_4465,N_4367,N_4266);
and U4466 (N_4466,N_4315,N_4205);
nand U4467 (N_4467,N_4381,N_4249);
and U4468 (N_4468,N_4298,N_4230);
nor U4469 (N_4469,N_4377,N_4270);
nand U4470 (N_4470,N_4207,N_4325);
nor U4471 (N_4471,N_4276,N_4360);
nand U4472 (N_4472,N_4253,N_4393);
or U4473 (N_4473,N_4269,N_4392);
or U4474 (N_4474,N_4355,N_4263);
nor U4475 (N_4475,N_4233,N_4289);
or U4476 (N_4476,N_4241,N_4399);
nand U4477 (N_4477,N_4363,N_4208);
or U4478 (N_4478,N_4374,N_4260);
and U4479 (N_4479,N_4214,N_4254);
nand U4480 (N_4480,N_4244,N_4326);
nand U4481 (N_4481,N_4278,N_4285);
or U4482 (N_4482,N_4243,N_4300);
nand U4483 (N_4483,N_4262,N_4334);
nand U4484 (N_4484,N_4330,N_4323);
nor U4485 (N_4485,N_4202,N_4283);
or U4486 (N_4486,N_4290,N_4304);
or U4487 (N_4487,N_4303,N_4256);
and U4488 (N_4488,N_4259,N_4376);
or U4489 (N_4489,N_4383,N_4251);
nand U4490 (N_4490,N_4204,N_4349);
or U4491 (N_4491,N_4291,N_4384);
or U4492 (N_4492,N_4390,N_4232);
or U4493 (N_4493,N_4223,N_4320);
nor U4494 (N_4494,N_4310,N_4234);
nand U4495 (N_4495,N_4282,N_4394);
nor U4496 (N_4496,N_4281,N_4272);
and U4497 (N_4497,N_4364,N_4311);
and U4498 (N_4498,N_4351,N_4341);
and U4499 (N_4499,N_4271,N_4274);
nor U4500 (N_4500,N_4301,N_4295);
and U4501 (N_4501,N_4369,N_4359);
and U4502 (N_4502,N_4353,N_4340);
or U4503 (N_4503,N_4246,N_4382);
or U4504 (N_4504,N_4371,N_4292);
and U4505 (N_4505,N_4345,N_4251);
and U4506 (N_4506,N_4386,N_4393);
and U4507 (N_4507,N_4313,N_4286);
and U4508 (N_4508,N_4267,N_4296);
or U4509 (N_4509,N_4209,N_4397);
or U4510 (N_4510,N_4328,N_4233);
nand U4511 (N_4511,N_4207,N_4215);
nor U4512 (N_4512,N_4224,N_4377);
nor U4513 (N_4513,N_4239,N_4225);
or U4514 (N_4514,N_4249,N_4294);
nand U4515 (N_4515,N_4316,N_4389);
and U4516 (N_4516,N_4223,N_4236);
nand U4517 (N_4517,N_4387,N_4353);
and U4518 (N_4518,N_4220,N_4334);
nand U4519 (N_4519,N_4317,N_4329);
or U4520 (N_4520,N_4312,N_4236);
and U4521 (N_4521,N_4277,N_4236);
or U4522 (N_4522,N_4329,N_4206);
nor U4523 (N_4523,N_4377,N_4207);
and U4524 (N_4524,N_4201,N_4323);
and U4525 (N_4525,N_4382,N_4261);
and U4526 (N_4526,N_4231,N_4307);
and U4527 (N_4527,N_4225,N_4206);
or U4528 (N_4528,N_4385,N_4366);
and U4529 (N_4529,N_4279,N_4212);
or U4530 (N_4530,N_4366,N_4378);
and U4531 (N_4531,N_4354,N_4297);
nor U4532 (N_4532,N_4236,N_4364);
nand U4533 (N_4533,N_4297,N_4367);
or U4534 (N_4534,N_4300,N_4246);
or U4535 (N_4535,N_4383,N_4245);
and U4536 (N_4536,N_4379,N_4361);
nor U4537 (N_4537,N_4240,N_4375);
nor U4538 (N_4538,N_4399,N_4358);
nor U4539 (N_4539,N_4358,N_4348);
and U4540 (N_4540,N_4348,N_4380);
nand U4541 (N_4541,N_4231,N_4305);
nand U4542 (N_4542,N_4378,N_4342);
nand U4543 (N_4543,N_4332,N_4322);
nand U4544 (N_4544,N_4254,N_4340);
and U4545 (N_4545,N_4393,N_4379);
nor U4546 (N_4546,N_4235,N_4207);
nand U4547 (N_4547,N_4201,N_4200);
or U4548 (N_4548,N_4373,N_4255);
nand U4549 (N_4549,N_4377,N_4397);
nor U4550 (N_4550,N_4262,N_4329);
and U4551 (N_4551,N_4365,N_4265);
nand U4552 (N_4552,N_4360,N_4341);
nand U4553 (N_4553,N_4231,N_4298);
and U4554 (N_4554,N_4272,N_4373);
nand U4555 (N_4555,N_4389,N_4297);
nand U4556 (N_4556,N_4341,N_4365);
nor U4557 (N_4557,N_4380,N_4230);
nor U4558 (N_4558,N_4219,N_4291);
or U4559 (N_4559,N_4305,N_4248);
or U4560 (N_4560,N_4382,N_4365);
nor U4561 (N_4561,N_4364,N_4339);
nor U4562 (N_4562,N_4367,N_4370);
and U4563 (N_4563,N_4298,N_4286);
nand U4564 (N_4564,N_4241,N_4216);
nor U4565 (N_4565,N_4335,N_4243);
nand U4566 (N_4566,N_4251,N_4268);
or U4567 (N_4567,N_4271,N_4239);
nand U4568 (N_4568,N_4398,N_4290);
and U4569 (N_4569,N_4260,N_4240);
or U4570 (N_4570,N_4309,N_4307);
or U4571 (N_4571,N_4283,N_4316);
and U4572 (N_4572,N_4305,N_4390);
or U4573 (N_4573,N_4239,N_4283);
nand U4574 (N_4574,N_4283,N_4268);
nand U4575 (N_4575,N_4266,N_4328);
nand U4576 (N_4576,N_4263,N_4209);
and U4577 (N_4577,N_4390,N_4238);
nor U4578 (N_4578,N_4281,N_4357);
nor U4579 (N_4579,N_4281,N_4381);
nor U4580 (N_4580,N_4337,N_4307);
and U4581 (N_4581,N_4324,N_4207);
and U4582 (N_4582,N_4393,N_4399);
and U4583 (N_4583,N_4301,N_4203);
and U4584 (N_4584,N_4276,N_4328);
nor U4585 (N_4585,N_4217,N_4385);
nor U4586 (N_4586,N_4306,N_4338);
nor U4587 (N_4587,N_4278,N_4306);
and U4588 (N_4588,N_4375,N_4296);
nor U4589 (N_4589,N_4209,N_4218);
and U4590 (N_4590,N_4200,N_4289);
nand U4591 (N_4591,N_4294,N_4318);
nand U4592 (N_4592,N_4332,N_4290);
nand U4593 (N_4593,N_4363,N_4373);
nand U4594 (N_4594,N_4339,N_4395);
or U4595 (N_4595,N_4302,N_4223);
xor U4596 (N_4596,N_4284,N_4328);
and U4597 (N_4597,N_4365,N_4235);
and U4598 (N_4598,N_4225,N_4289);
nand U4599 (N_4599,N_4210,N_4358);
nor U4600 (N_4600,N_4461,N_4586);
nand U4601 (N_4601,N_4472,N_4520);
or U4602 (N_4602,N_4409,N_4523);
nor U4603 (N_4603,N_4556,N_4438);
and U4604 (N_4604,N_4419,N_4506);
xnor U4605 (N_4605,N_4403,N_4540);
or U4606 (N_4606,N_4522,N_4598);
or U4607 (N_4607,N_4476,N_4532);
nand U4608 (N_4608,N_4538,N_4584);
nand U4609 (N_4609,N_4485,N_4565);
nand U4610 (N_4610,N_4544,N_4497);
or U4611 (N_4611,N_4549,N_4402);
nand U4612 (N_4612,N_4588,N_4559);
nor U4613 (N_4613,N_4487,N_4560);
and U4614 (N_4614,N_4516,N_4460);
nand U4615 (N_4615,N_4596,N_4443);
or U4616 (N_4616,N_4488,N_4589);
and U4617 (N_4617,N_4468,N_4441);
nand U4618 (N_4618,N_4495,N_4546);
or U4619 (N_4619,N_4452,N_4470);
and U4620 (N_4620,N_4545,N_4406);
nand U4621 (N_4621,N_4510,N_4491);
or U4622 (N_4622,N_4531,N_4496);
nand U4623 (N_4623,N_4494,N_4473);
nor U4624 (N_4624,N_4423,N_4412);
nor U4625 (N_4625,N_4416,N_4562);
nand U4626 (N_4626,N_4407,N_4555);
xnor U4627 (N_4627,N_4587,N_4534);
and U4628 (N_4628,N_4552,N_4554);
or U4629 (N_4629,N_4575,N_4542);
or U4630 (N_4630,N_4521,N_4459);
nor U4631 (N_4631,N_4400,N_4440);
nor U4632 (N_4632,N_4515,N_4401);
nand U4633 (N_4633,N_4502,N_4415);
nand U4634 (N_4634,N_4594,N_4424);
nor U4635 (N_4635,N_4498,N_4585);
xor U4636 (N_4636,N_4570,N_4539);
or U4637 (N_4637,N_4529,N_4478);
and U4638 (N_4638,N_4490,N_4527);
nor U4639 (N_4639,N_4535,N_4507);
nand U4640 (N_4640,N_4553,N_4493);
nand U4641 (N_4641,N_4404,N_4500);
nor U4642 (N_4642,N_4433,N_4482);
nor U4643 (N_4643,N_4595,N_4449);
and U4644 (N_4644,N_4526,N_4480);
and U4645 (N_4645,N_4450,N_4445);
and U4646 (N_4646,N_4574,N_4474);
or U4647 (N_4647,N_4489,N_4479);
nand U4648 (N_4648,N_4466,N_4467);
nor U4649 (N_4649,N_4557,N_4426);
nor U4650 (N_4650,N_4592,N_4519);
nand U4651 (N_4651,N_4590,N_4477);
nor U4652 (N_4652,N_4536,N_4503);
nor U4653 (N_4653,N_4517,N_4513);
nor U4654 (N_4654,N_4437,N_4505);
nor U4655 (N_4655,N_4469,N_4561);
or U4656 (N_4656,N_4564,N_4569);
and U4657 (N_4657,N_4548,N_4444);
and U4658 (N_4658,N_4448,N_4576);
nor U4659 (N_4659,N_4465,N_4573);
nand U4660 (N_4660,N_4411,N_4432);
nand U4661 (N_4661,N_4541,N_4434);
or U4662 (N_4662,N_4579,N_4446);
or U4663 (N_4663,N_4512,N_4525);
nor U4664 (N_4664,N_4453,N_4550);
or U4665 (N_4665,N_4435,N_4421);
and U4666 (N_4666,N_4431,N_4509);
nor U4667 (N_4667,N_4456,N_4457);
and U4668 (N_4668,N_4442,N_4577);
or U4669 (N_4669,N_4551,N_4566);
or U4670 (N_4670,N_4518,N_4583);
and U4671 (N_4671,N_4528,N_4563);
and U4672 (N_4672,N_4462,N_4501);
nand U4673 (N_4673,N_4414,N_4454);
xor U4674 (N_4674,N_4581,N_4410);
nand U4675 (N_4675,N_4405,N_4593);
and U4676 (N_4676,N_4486,N_4455);
or U4677 (N_4677,N_4475,N_4451);
or U4678 (N_4678,N_4547,N_4591);
nand U4679 (N_4679,N_4582,N_4483);
and U4680 (N_4680,N_4567,N_4417);
nor U4681 (N_4681,N_4499,N_4458);
nor U4682 (N_4682,N_4508,N_4537);
nor U4683 (N_4683,N_4420,N_4447);
nor U4684 (N_4684,N_4578,N_4533);
or U4685 (N_4685,N_4543,N_4439);
and U4686 (N_4686,N_4481,N_4571);
and U4687 (N_4687,N_4599,N_4524);
or U4688 (N_4688,N_4408,N_4413);
nor U4689 (N_4689,N_4597,N_4436);
or U4690 (N_4690,N_4464,N_4558);
nor U4691 (N_4691,N_4430,N_4511);
and U4692 (N_4692,N_4572,N_4471);
nand U4693 (N_4693,N_4422,N_4425);
xor U4694 (N_4694,N_4492,N_4429);
and U4695 (N_4695,N_4463,N_4418);
or U4696 (N_4696,N_4504,N_4427);
or U4697 (N_4697,N_4568,N_4484);
nor U4698 (N_4698,N_4530,N_4514);
nor U4699 (N_4699,N_4428,N_4580);
and U4700 (N_4700,N_4477,N_4478);
nand U4701 (N_4701,N_4479,N_4575);
nand U4702 (N_4702,N_4430,N_4550);
nand U4703 (N_4703,N_4488,N_4419);
and U4704 (N_4704,N_4560,N_4481);
xnor U4705 (N_4705,N_4473,N_4488);
or U4706 (N_4706,N_4587,N_4439);
or U4707 (N_4707,N_4593,N_4572);
or U4708 (N_4708,N_4450,N_4537);
nand U4709 (N_4709,N_4495,N_4433);
nor U4710 (N_4710,N_4534,N_4574);
nor U4711 (N_4711,N_4567,N_4536);
nand U4712 (N_4712,N_4473,N_4426);
nor U4713 (N_4713,N_4586,N_4546);
nand U4714 (N_4714,N_4453,N_4475);
nand U4715 (N_4715,N_4566,N_4483);
nand U4716 (N_4716,N_4419,N_4549);
or U4717 (N_4717,N_4558,N_4418);
and U4718 (N_4718,N_4496,N_4499);
nor U4719 (N_4719,N_4464,N_4483);
or U4720 (N_4720,N_4407,N_4459);
nor U4721 (N_4721,N_4401,N_4431);
and U4722 (N_4722,N_4556,N_4471);
xnor U4723 (N_4723,N_4545,N_4563);
or U4724 (N_4724,N_4535,N_4429);
and U4725 (N_4725,N_4414,N_4513);
and U4726 (N_4726,N_4560,N_4496);
or U4727 (N_4727,N_4475,N_4513);
and U4728 (N_4728,N_4593,N_4589);
or U4729 (N_4729,N_4563,N_4543);
nand U4730 (N_4730,N_4564,N_4491);
nand U4731 (N_4731,N_4455,N_4592);
nand U4732 (N_4732,N_4406,N_4478);
or U4733 (N_4733,N_4475,N_4495);
or U4734 (N_4734,N_4586,N_4414);
nor U4735 (N_4735,N_4409,N_4461);
nand U4736 (N_4736,N_4539,N_4416);
nor U4737 (N_4737,N_4471,N_4480);
or U4738 (N_4738,N_4490,N_4466);
or U4739 (N_4739,N_4470,N_4598);
nor U4740 (N_4740,N_4528,N_4469);
xor U4741 (N_4741,N_4586,N_4447);
nand U4742 (N_4742,N_4590,N_4419);
nand U4743 (N_4743,N_4455,N_4552);
and U4744 (N_4744,N_4586,N_4511);
or U4745 (N_4745,N_4485,N_4448);
or U4746 (N_4746,N_4432,N_4583);
and U4747 (N_4747,N_4432,N_4448);
and U4748 (N_4748,N_4594,N_4445);
nor U4749 (N_4749,N_4502,N_4480);
nor U4750 (N_4750,N_4420,N_4522);
nor U4751 (N_4751,N_4514,N_4409);
nor U4752 (N_4752,N_4455,N_4537);
or U4753 (N_4753,N_4509,N_4583);
and U4754 (N_4754,N_4505,N_4466);
or U4755 (N_4755,N_4599,N_4452);
nor U4756 (N_4756,N_4477,N_4495);
or U4757 (N_4757,N_4560,N_4519);
and U4758 (N_4758,N_4567,N_4401);
and U4759 (N_4759,N_4547,N_4438);
and U4760 (N_4760,N_4549,N_4531);
nor U4761 (N_4761,N_4545,N_4540);
nand U4762 (N_4762,N_4514,N_4567);
nand U4763 (N_4763,N_4418,N_4552);
and U4764 (N_4764,N_4522,N_4432);
or U4765 (N_4765,N_4400,N_4437);
nand U4766 (N_4766,N_4480,N_4407);
xnor U4767 (N_4767,N_4536,N_4514);
and U4768 (N_4768,N_4433,N_4412);
and U4769 (N_4769,N_4457,N_4414);
or U4770 (N_4770,N_4543,N_4454);
or U4771 (N_4771,N_4418,N_4442);
nor U4772 (N_4772,N_4479,N_4566);
nand U4773 (N_4773,N_4586,N_4434);
nand U4774 (N_4774,N_4491,N_4556);
nor U4775 (N_4775,N_4415,N_4589);
and U4776 (N_4776,N_4432,N_4571);
nand U4777 (N_4777,N_4532,N_4530);
and U4778 (N_4778,N_4414,N_4588);
xor U4779 (N_4779,N_4483,N_4578);
nor U4780 (N_4780,N_4404,N_4593);
xnor U4781 (N_4781,N_4467,N_4431);
or U4782 (N_4782,N_4524,N_4401);
nor U4783 (N_4783,N_4425,N_4544);
and U4784 (N_4784,N_4583,N_4496);
nand U4785 (N_4785,N_4539,N_4495);
and U4786 (N_4786,N_4511,N_4565);
nor U4787 (N_4787,N_4524,N_4451);
nand U4788 (N_4788,N_4534,N_4466);
or U4789 (N_4789,N_4500,N_4546);
nand U4790 (N_4790,N_4542,N_4547);
and U4791 (N_4791,N_4577,N_4491);
or U4792 (N_4792,N_4457,N_4466);
nand U4793 (N_4793,N_4418,N_4502);
and U4794 (N_4794,N_4485,N_4542);
nand U4795 (N_4795,N_4597,N_4538);
and U4796 (N_4796,N_4457,N_4460);
or U4797 (N_4797,N_4540,N_4429);
and U4798 (N_4798,N_4462,N_4539);
and U4799 (N_4799,N_4449,N_4548);
or U4800 (N_4800,N_4663,N_4711);
or U4801 (N_4801,N_4690,N_4698);
nand U4802 (N_4802,N_4620,N_4714);
or U4803 (N_4803,N_4798,N_4708);
nand U4804 (N_4804,N_4695,N_4748);
xor U4805 (N_4805,N_4785,N_4650);
or U4806 (N_4806,N_4769,N_4678);
or U4807 (N_4807,N_4693,N_4704);
and U4808 (N_4808,N_4749,N_4608);
nor U4809 (N_4809,N_4644,N_4709);
or U4810 (N_4810,N_4787,N_4659);
and U4811 (N_4811,N_4782,N_4655);
or U4812 (N_4812,N_4600,N_4673);
nand U4813 (N_4813,N_4780,N_4639);
and U4814 (N_4814,N_4736,N_4765);
nor U4815 (N_4815,N_4768,N_4689);
nor U4816 (N_4816,N_4773,N_4627);
nand U4817 (N_4817,N_4624,N_4640);
nor U4818 (N_4818,N_4633,N_4746);
and U4819 (N_4819,N_4604,N_4799);
or U4820 (N_4820,N_4617,N_4751);
or U4821 (N_4821,N_4646,N_4747);
nand U4822 (N_4822,N_4727,N_4665);
nand U4823 (N_4823,N_4792,N_4738);
nand U4824 (N_4824,N_4712,N_4767);
or U4825 (N_4825,N_4623,N_4726);
nand U4826 (N_4826,N_4734,N_4651);
and U4827 (N_4827,N_4752,N_4713);
nand U4828 (N_4828,N_4631,N_4789);
nand U4829 (N_4829,N_4664,N_4603);
and U4830 (N_4830,N_4696,N_4694);
and U4831 (N_4831,N_4705,N_4618);
and U4832 (N_4832,N_4697,N_4610);
nand U4833 (N_4833,N_4786,N_4615);
and U4834 (N_4834,N_4629,N_4756);
nor U4835 (N_4835,N_4759,N_4692);
nand U4836 (N_4836,N_4779,N_4670);
nor U4837 (N_4837,N_4757,N_4637);
nor U4838 (N_4838,N_4647,N_4741);
or U4839 (N_4839,N_4658,N_4775);
nor U4840 (N_4840,N_4662,N_4732);
nand U4841 (N_4841,N_4602,N_4717);
or U4842 (N_4842,N_4621,N_4794);
and U4843 (N_4843,N_4706,N_4703);
nor U4844 (N_4844,N_4636,N_4721);
nand U4845 (N_4845,N_4771,N_4700);
or U4846 (N_4846,N_4630,N_4777);
xnor U4847 (N_4847,N_4683,N_4761);
xor U4848 (N_4848,N_4722,N_4740);
and U4849 (N_4849,N_4686,N_4795);
and U4850 (N_4850,N_4657,N_4628);
and U4851 (N_4851,N_4681,N_4783);
or U4852 (N_4852,N_4677,N_4676);
nand U4853 (N_4853,N_4772,N_4605);
nand U4854 (N_4854,N_4774,N_4744);
and U4855 (N_4855,N_4601,N_4660);
or U4856 (N_4856,N_4754,N_4652);
and U4857 (N_4857,N_4720,N_4671);
and U4858 (N_4858,N_4674,N_4788);
and U4859 (N_4859,N_4725,N_4699);
and U4860 (N_4860,N_4762,N_4730);
and U4861 (N_4861,N_4619,N_4611);
nor U4862 (N_4862,N_4760,N_4764);
and U4863 (N_4863,N_4728,N_4638);
or U4864 (N_4864,N_4733,N_4763);
nand U4865 (N_4865,N_4632,N_4616);
nand U4866 (N_4866,N_4770,N_4743);
nor U4867 (N_4867,N_4641,N_4653);
nor U4868 (N_4868,N_4609,N_4626);
or U4869 (N_4869,N_4614,N_4622);
nor U4870 (N_4870,N_4680,N_4669);
or U4871 (N_4871,N_4634,N_4648);
or U4872 (N_4872,N_4635,N_4758);
and U4873 (N_4873,N_4766,N_4723);
and U4874 (N_4874,N_4750,N_4691);
or U4875 (N_4875,N_4642,N_4781);
xor U4876 (N_4876,N_4682,N_4643);
nor U4877 (N_4877,N_4745,N_4668);
or U4878 (N_4878,N_4729,N_4719);
and U4879 (N_4879,N_4612,N_4687);
nor U4880 (N_4880,N_4742,N_4702);
and U4881 (N_4881,N_4753,N_4716);
nor U4882 (N_4882,N_4649,N_4661);
nand U4883 (N_4883,N_4688,N_4797);
nor U4884 (N_4884,N_4613,N_4656);
xnor U4885 (N_4885,N_4684,N_4735);
and U4886 (N_4886,N_4778,N_4672);
nor U4887 (N_4887,N_4784,N_4731);
and U4888 (N_4888,N_4776,N_4606);
and U4889 (N_4889,N_4790,N_4654);
nor U4890 (N_4890,N_4737,N_4707);
nand U4891 (N_4891,N_4793,N_4685);
or U4892 (N_4892,N_4675,N_4724);
xor U4893 (N_4893,N_4645,N_4739);
nand U4894 (N_4894,N_4718,N_4701);
nand U4895 (N_4895,N_4796,N_4679);
nand U4896 (N_4896,N_4625,N_4667);
nand U4897 (N_4897,N_4710,N_4715);
or U4898 (N_4898,N_4755,N_4666);
and U4899 (N_4899,N_4607,N_4791);
or U4900 (N_4900,N_4674,N_4737);
nor U4901 (N_4901,N_4741,N_4676);
nand U4902 (N_4902,N_4659,N_4669);
nor U4903 (N_4903,N_4704,N_4736);
nor U4904 (N_4904,N_4690,N_4758);
and U4905 (N_4905,N_4752,N_4672);
xor U4906 (N_4906,N_4730,N_4656);
nor U4907 (N_4907,N_4752,N_4739);
and U4908 (N_4908,N_4760,N_4714);
xor U4909 (N_4909,N_4660,N_4623);
nand U4910 (N_4910,N_4649,N_4732);
nor U4911 (N_4911,N_4797,N_4671);
or U4912 (N_4912,N_4663,N_4641);
nor U4913 (N_4913,N_4761,N_4753);
nand U4914 (N_4914,N_4624,N_4625);
nand U4915 (N_4915,N_4740,N_4616);
or U4916 (N_4916,N_4611,N_4632);
nand U4917 (N_4917,N_4784,N_4687);
nand U4918 (N_4918,N_4731,N_4764);
or U4919 (N_4919,N_4788,N_4712);
nor U4920 (N_4920,N_4763,N_4608);
nand U4921 (N_4921,N_4785,N_4711);
and U4922 (N_4922,N_4710,N_4789);
nand U4923 (N_4923,N_4681,N_4683);
or U4924 (N_4924,N_4678,N_4761);
nor U4925 (N_4925,N_4662,N_4772);
nand U4926 (N_4926,N_4616,N_4648);
and U4927 (N_4927,N_4707,N_4668);
or U4928 (N_4928,N_4794,N_4675);
nand U4929 (N_4929,N_4682,N_4767);
or U4930 (N_4930,N_4781,N_4761);
nor U4931 (N_4931,N_4734,N_4752);
and U4932 (N_4932,N_4685,N_4727);
or U4933 (N_4933,N_4617,N_4629);
nand U4934 (N_4934,N_4692,N_4767);
nor U4935 (N_4935,N_4775,N_4692);
or U4936 (N_4936,N_4665,N_4735);
nand U4937 (N_4937,N_4754,N_4764);
nor U4938 (N_4938,N_4735,N_4621);
nand U4939 (N_4939,N_4606,N_4778);
or U4940 (N_4940,N_4736,N_4766);
nand U4941 (N_4941,N_4727,N_4642);
nor U4942 (N_4942,N_4720,N_4618);
or U4943 (N_4943,N_4661,N_4741);
or U4944 (N_4944,N_4711,N_4639);
nor U4945 (N_4945,N_4692,N_4611);
and U4946 (N_4946,N_4618,N_4643);
or U4947 (N_4947,N_4673,N_4694);
or U4948 (N_4948,N_4631,N_4742);
or U4949 (N_4949,N_4711,N_4779);
nand U4950 (N_4950,N_4735,N_4699);
nor U4951 (N_4951,N_4606,N_4740);
nor U4952 (N_4952,N_4699,N_4723);
or U4953 (N_4953,N_4747,N_4701);
nor U4954 (N_4954,N_4620,N_4783);
nor U4955 (N_4955,N_4617,N_4660);
nor U4956 (N_4956,N_4621,N_4662);
or U4957 (N_4957,N_4637,N_4684);
nand U4958 (N_4958,N_4748,N_4616);
nand U4959 (N_4959,N_4716,N_4762);
nor U4960 (N_4960,N_4716,N_4754);
or U4961 (N_4961,N_4675,N_4766);
nor U4962 (N_4962,N_4611,N_4778);
or U4963 (N_4963,N_4790,N_4751);
or U4964 (N_4964,N_4735,N_4773);
nand U4965 (N_4965,N_4682,N_4601);
nor U4966 (N_4966,N_4659,N_4672);
or U4967 (N_4967,N_4692,N_4670);
nor U4968 (N_4968,N_4609,N_4715);
nor U4969 (N_4969,N_4791,N_4712);
xor U4970 (N_4970,N_4666,N_4743);
nor U4971 (N_4971,N_4777,N_4699);
nor U4972 (N_4972,N_4749,N_4779);
and U4973 (N_4973,N_4775,N_4604);
nand U4974 (N_4974,N_4639,N_4799);
nand U4975 (N_4975,N_4657,N_4750);
nor U4976 (N_4976,N_4731,N_4707);
or U4977 (N_4977,N_4694,N_4645);
and U4978 (N_4978,N_4744,N_4717);
nor U4979 (N_4979,N_4742,N_4781);
or U4980 (N_4980,N_4697,N_4718);
and U4981 (N_4981,N_4681,N_4710);
nand U4982 (N_4982,N_4721,N_4613);
or U4983 (N_4983,N_4655,N_4675);
and U4984 (N_4984,N_4761,N_4695);
and U4985 (N_4985,N_4775,N_4712);
nor U4986 (N_4986,N_4776,N_4741);
or U4987 (N_4987,N_4757,N_4617);
and U4988 (N_4988,N_4755,N_4793);
or U4989 (N_4989,N_4693,N_4697);
or U4990 (N_4990,N_4636,N_4644);
nor U4991 (N_4991,N_4612,N_4775);
or U4992 (N_4992,N_4728,N_4661);
or U4993 (N_4993,N_4688,N_4609);
and U4994 (N_4994,N_4799,N_4706);
xor U4995 (N_4995,N_4725,N_4613);
and U4996 (N_4996,N_4755,N_4694);
or U4997 (N_4997,N_4731,N_4791);
or U4998 (N_4998,N_4717,N_4637);
and U4999 (N_4999,N_4665,N_4776);
nor UO_0 (O_0,N_4935,N_4887);
or UO_1 (O_1,N_4874,N_4856);
nand UO_2 (O_2,N_4995,N_4901);
nor UO_3 (O_3,N_4885,N_4976);
or UO_4 (O_4,N_4979,N_4884);
nand UO_5 (O_5,N_4883,N_4934);
nor UO_6 (O_6,N_4802,N_4951);
or UO_7 (O_7,N_4871,N_4906);
and UO_8 (O_8,N_4973,N_4959);
nand UO_9 (O_9,N_4994,N_4840);
nor UO_10 (O_10,N_4913,N_4866);
and UO_11 (O_11,N_4957,N_4952);
nor UO_12 (O_12,N_4836,N_4868);
xor UO_13 (O_13,N_4929,N_4851);
and UO_14 (O_14,N_4982,N_4997);
and UO_15 (O_15,N_4949,N_4841);
nand UO_16 (O_16,N_4872,N_4941);
nor UO_17 (O_17,N_4916,N_4947);
nor UO_18 (O_18,N_4939,N_4870);
or UO_19 (O_19,N_4818,N_4888);
nand UO_20 (O_20,N_4817,N_4930);
or UO_21 (O_21,N_4940,N_4953);
nor UO_22 (O_22,N_4920,N_4985);
or UO_23 (O_23,N_4805,N_4911);
nand UO_24 (O_24,N_4816,N_4926);
and UO_25 (O_25,N_4865,N_4830);
or UO_26 (O_26,N_4955,N_4891);
and UO_27 (O_27,N_4964,N_4900);
nand UO_28 (O_28,N_4855,N_4825);
nand UO_29 (O_29,N_4815,N_4958);
and UO_30 (O_30,N_4838,N_4873);
nand UO_31 (O_31,N_4814,N_4878);
or UO_32 (O_32,N_4806,N_4993);
or UO_33 (O_33,N_4936,N_4899);
nor UO_34 (O_34,N_4902,N_4864);
or UO_35 (O_35,N_4923,N_4835);
and UO_36 (O_36,N_4813,N_4827);
nand UO_37 (O_37,N_4989,N_4889);
xnor UO_38 (O_38,N_4962,N_4990);
nor UO_39 (O_39,N_4845,N_4998);
and UO_40 (O_40,N_4894,N_4974);
nand UO_41 (O_41,N_4892,N_4843);
or UO_42 (O_42,N_4984,N_4965);
nor UO_43 (O_43,N_4981,N_4980);
and UO_44 (O_44,N_4969,N_4839);
and UO_45 (O_45,N_4854,N_4919);
and UO_46 (O_46,N_4846,N_4876);
nand UO_47 (O_47,N_4967,N_4971);
or UO_48 (O_48,N_4860,N_4928);
nand UO_49 (O_49,N_4983,N_4869);
nor UO_50 (O_50,N_4831,N_4946);
nor UO_51 (O_51,N_4880,N_4897);
or UO_52 (O_52,N_4988,N_4963);
nor UO_53 (O_53,N_4890,N_4886);
or UO_54 (O_54,N_4862,N_4850);
nand UO_55 (O_55,N_4898,N_4937);
or UO_56 (O_56,N_4849,N_4822);
nor UO_57 (O_57,N_4833,N_4931);
or UO_58 (O_58,N_4942,N_4970);
and UO_59 (O_59,N_4853,N_4991);
nor UO_60 (O_60,N_4933,N_4832);
or UO_61 (O_61,N_4918,N_4948);
and UO_62 (O_62,N_4820,N_4895);
nor UO_63 (O_63,N_4924,N_4999);
nand UO_64 (O_64,N_4972,N_4800);
nor UO_65 (O_65,N_4803,N_4828);
or UO_66 (O_66,N_4807,N_4977);
nor UO_67 (O_67,N_4804,N_4961);
and UO_68 (O_68,N_4896,N_4821);
or UO_69 (O_69,N_4819,N_4861);
xor UO_70 (O_70,N_4914,N_4968);
nor UO_71 (O_71,N_4811,N_4944);
nand UO_72 (O_72,N_4875,N_4992);
nor UO_73 (O_73,N_4986,N_4954);
nor UO_74 (O_74,N_4812,N_4847);
nor UO_75 (O_75,N_4921,N_4823);
xnor UO_76 (O_76,N_4837,N_4829);
nor UO_77 (O_77,N_4996,N_4858);
or UO_78 (O_78,N_4917,N_4857);
nor UO_79 (O_79,N_4826,N_4960);
nand UO_80 (O_80,N_4882,N_4925);
nor UO_81 (O_81,N_4879,N_4943);
or UO_82 (O_82,N_4950,N_4867);
and UO_83 (O_83,N_4834,N_4844);
xor UO_84 (O_84,N_4910,N_4987);
or UO_85 (O_85,N_4848,N_4907);
nor UO_86 (O_86,N_4932,N_4842);
nor UO_87 (O_87,N_4809,N_4905);
and UO_88 (O_88,N_4801,N_4938);
xnor UO_89 (O_89,N_4893,N_4956);
or UO_90 (O_90,N_4945,N_4810);
nand UO_91 (O_91,N_4824,N_4915);
or UO_92 (O_92,N_4881,N_4859);
and UO_93 (O_93,N_4908,N_4912);
or UO_94 (O_94,N_4877,N_4978);
nor UO_95 (O_95,N_4863,N_4904);
or UO_96 (O_96,N_4852,N_4922);
nor UO_97 (O_97,N_4927,N_4808);
nor UO_98 (O_98,N_4903,N_4975);
nand UO_99 (O_99,N_4909,N_4966);
or UO_100 (O_100,N_4933,N_4885);
nand UO_101 (O_101,N_4880,N_4879);
nor UO_102 (O_102,N_4851,N_4913);
nor UO_103 (O_103,N_4958,N_4931);
or UO_104 (O_104,N_4987,N_4819);
and UO_105 (O_105,N_4810,N_4904);
and UO_106 (O_106,N_4948,N_4897);
nor UO_107 (O_107,N_4855,N_4930);
or UO_108 (O_108,N_4883,N_4901);
nor UO_109 (O_109,N_4896,N_4811);
nand UO_110 (O_110,N_4994,N_4877);
nand UO_111 (O_111,N_4986,N_4809);
nor UO_112 (O_112,N_4816,N_4930);
or UO_113 (O_113,N_4825,N_4856);
nor UO_114 (O_114,N_4884,N_4863);
nor UO_115 (O_115,N_4855,N_4916);
nor UO_116 (O_116,N_4870,N_4851);
or UO_117 (O_117,N_4880,N_4815);
nand UO_118 (O_118,N_4890,N_4841);
or UO_119 (O_119,N_4914,N_4960);
nor UO_120 (O_120,N_4886,N_4917);
and UO_121 (O_121,N_4990,N_4844);
or UO_122 (O_122,N_4927,N_4886);
and UO_123 (O_123,N_4980,N_4928);
or UO_124 (O_124,N_4964,N_4851);
nor UO_125 (O_125,N_4827,N_4930);
and UO_126 (O_126,N_4978,N_4884);
and UO_127 (O_127,N_4843,N_4905);
nand UO_128 (O_128,N_4860,N_4911);
nor UO_129 (O_129,N_4871,N_4932);
nand UO_130 (O_130,N_4876,N_4962);
nand UO_131 (O_131,N_4828,N_4843);
nand UO_132 (O_132,N_4860,N_4820);
or UO_133 (O_133,N_4813,N_4812);
xor UO_134 (O_134,N_4870,N_4844);
or UO_135 (O_135,N_4939,N_4905);
nand UO_136 (O_136,N_4992,N_4856);
nor UO_137 (O_137,N_4809,N_4836);
or UO_138 (O_138,N_4971,N_4861);
and UO_139 (O_139,N_4816,N_4949);
nor UO_140 (O_140,N_4926,N_4884);
nor UO_141 (O_141,N_4846,N_4890);
nand UO_142 (O_142,N_4874,N_4947);
or UO_143 (O_143,N_4813,N_4839);
nor UO_144 (O_144,N_4881,N_4807);
and UO_145 (O_145,N_4960,N_4888);
or UO_146 (O_146,N_4816,N_4947);
nor UO_147 (O_147,N_4852,N_4807);
nor UO_148 (O_148,N_4979,N_4829);
xnor UO_149 (O_149,N_4996,N_4862);
or UO_150 (O_150,N_4821,N_4945);
and UO_151 (O_151,N_4901,N_4969);
nor UO_152 (O_152,N_4893,N_4805);
and UO_153 (O_153,N_4881,N_4968);
or UO_154 (O_154,N_4906,N_4934);
nand UO_155 (O_155,N_4973,N_4934);
and UO_156 (O_156,N_4837,N_4976);
nand UO_157 (O_157,N_4815,N_4884);
nor UO_158 (O_158,N_4955,N_4805);
nand UO_159 (O_159,N_4800,N_4979);
nand UO_160 (O_160,N_4981,N_4938);
or UO_161 (O_161,N_4894,N_4825);
nand UO_162 (O_162,N_4908,N_4855);
or UO_163 (O_163,N_4855,N_4803);
and UO_164 (O_164,N_4961,N_4814);
nor UO_165 (O_165,N_4959,N_4825);
and UO_166 (O_166,N_4903,N_4983);
nand UO_167 (O_167,N_4846,N_4828);
nor UO_168 (O_168,N_4964,N_4818);
nor UO_169 (O_169,N_4860,N_4916);
nor UO_170 (O_170,N_4861,N_4865);
nand UO_171 (O_171,N_4869,N_4968);
and UO_172 (O_172,N_4939,N_4824);
or UO_173 (O_173,N_4985,N_4854);
nor UO_174 (O_174,N_4971,N_4883);
nand UO_175 (O_175,N_4822,N_4978);
and UO_176 (O_176,N_4978,N_4864);
and UO_177 (O_177,N_4917,N_4959);
nor UO_178 (O_178,N_4924,N_4839);
nor UO_179 (O_179,N_4804,N_4805);
nor UO_180 (O_180,N_4975,N_4933);
nand UO_181 (O_181,N_4876,N_4815);
and UO_182 (O_182,N_4833,N_4860);
and UO_183 (O_183,N_4858,N_4809);
and UO_184 (O_184,N_4823,N_4982);
or UO_185 (O_185,N_4899,N_4907);
nand UO_186 (O_186,N_4904,N_4941);
and UO_187 (O_187,N_4923,N_4921);
and UO_188 (O_188,N_4865,N_4835);
nand UO_189 (O_189,N_4840,N_4893);
nand UO_190 (O_190,N_4935,N_4854);
nor UO_191 (O_191,N_4989,N_4839);
nand UO_192 (O_192,N_4963,N_4930);
or UO_193 (O_193,N_4990,N_4957);
nand UO_194 (O_194,N_4937,N_4810);
and UO_195 (O_195,N_4992,N_4801);
or UO_196 (O_196,N_4915,N_4917);
nor UO_197 (O_197,N_4859,N_4992);
nor UO_198 (O_198,N_4929,N_4958);
or UO_199 (O_199,N_4887,N_4918);
nor UO_200 (O_200,N_4869,N_4804);
nor UO_201 (O_201,N_4944,N_4802);
or UO_202 (O_202,N_4887,N_4956);
nor UO_203 (O_203,N_4826,N_4988);
nor UO_204 (O_204,N_4801,N_4865);
xor UO_205 (O_205,N_4848,N_4846);
and UO_206 (O_206,N_4991,N_4952);
or UO_207 (O_207,N_4936,N_4804);
nor UO_208 (O_208,N_4816,N_4975);
and UO_209 (O_209,N_4901,N_4914);
and UO_210 (O_210,N_4909,N_4988);
nand UO_211 (O_211,N_4823,N_4918);
nor UO_212 (O_212,N_4836,N_4897);
and UO_213 (O_213,N_4801,N_4849);
or UO_214 (O_214,N_4803,N_4864);
and UO_215 (O_215,N_4932,N_4989);
nand UO_216 (O_216,N_4808,N_4937);
nand UO_217 (O_217,N_4932,N_4914);
nor UO_218 (O_218,N_4971,N_4814);
and UO_219 (O_219,N_4983,N_4833);
nor UO_220 (O_220,N_4948,N_4874);
and UO_221 (O_221,N_4983,N_4988);
nand UO_222 (O_222,N_4981,N_4991);
nand UO_223 (O_223,N_4838,N_4991);
nand UO_224 (O_224,N_4946,N_4918);
xnor UO_225 (O_225,N_4960,N_4933);
xnor UO_226 (O_226,N_4836,N_4934);
nor UO_227 (O_227,N_4878,N_4801);
nand UO_228 (O_228,N_4984,N_4883);
nor UO_229 (O_229,N_4803,N_4898);
nand UO_230 (O_230,N_4847,N_4972);
nand UO_231 (O_231,N_4812,N_4927);
nor UO_232 (O_232,N_4935,N_4925);
nand UO_233 (O_233,N_4972,N_4840);
nand UO_234 (O_234,N_4884,N_4824);
or UO_235 (O_235,N_4900,N_4857);
nor UO_236 (O_236,N_4800,N_4973);
or UO_237 (O_237,N_4977,N_4805);
nor UO_238 (O_238,N_4822,N_4816);
nor UO_239 (O_239,N_4940,N_4807);
or UO_240 (O_240,N_4898,N_4965);
nor UO_241 (O_241,N_4821,N_4881);
nand UO_242 (O_242,N_4932,N_4939);
nand UO_243 (O_243,N_4951,N_4889);
or UO_244 (O_244,N_4831,N_4819);
nand UO_245 (O_245,N_4937,N_4802);
or UO_246 (O_246,N_4884,N_4845);
xnor UO_247 (O_247,N_4919,N_4885);
nor UO_248 (O_248,N_4800,N_4940);
or UO_249 (O_249,N_4907,N_4909);
and UO_250 (O_250,N_4910,N_4905);
xor UO_251 (O_251,N_4836,N_4856);
and UO_252 (O_252,N_4944,N_4896);
nor UO_253 (O_253,N_4882,N_4861);
nor UO_254 (O_254,N_4811,N_4818);
nand UO_255 (O_255,N_4946,N_4823);
nor UO_256 (O_256,N_4993,N_4809);
and UO_257 (O_257,N_4882,N_4992);
or UO_258 (O_258,N_4871,N_4992);
or UO_259 (O_259,N_4822,N_4992);
nor UO_260 (O_260,N_4966,N_4821);
or UO_261 (O_261,N_4973,N_4913);
or UO_262 (O_262,N_4935,N_4996);
and UO_263 (O_263,N_4885,N_4997);
nor UO_264 (O_264,N_4880,N_4990);
or UO_265 (O_265,N_4806,N_4907);
and UO_266 (O_266,N_4861,N_4972);
nor UO_267 (O_267,N_4865,N_4984);
and UO_268 (O_268,N_4914,N_4994);
nor UO_269 (O_269,N_4971,N_4920);
and UO_270 (O_270,N_4891,N_4980);
or UO_271 (O_271,N_4916,N_4971);
or UO_272 (O_272,N_4965,N_4949);
nand UO_273 (O_273,N_4997,N_4922);
or UO_274 (O_274,N_4879,N_4934);
nand UO_275 (O_275,N_4934,N_4821);
or UO_276 (O_276,N_4964,N_4866);
and UO_277 (O_277,N_4966,N_4917);
nor UO_278 (O_278,N_4872,N_4819);
and UO_279 (O_279,N_4957,N_4869);
nor UO_280 (O_280,N_4951,N_4874);
or UO_281 (O_281,N_4808,N_4976);
nor UO_282 (O_282,N_4801,N_4819);
or UO_283 (O_283,N_4901,N_4880);
nor UO_284 (O_284,N_4806,N_4975);
and UO_285 (O_285,N_4823,N_4808);
xnor UO_286 (O_286,N_4800,N_4898);
nor UO_287 (O_287,N_4810,N_4834);
nor UO_288 (O_288,N_4877,N_4842);
nor UO_289 (O_289,N_4920,N_4914);
nand UO_290 (O_290,N_4826,N_4985);
or UO_291 (O_291,N_4951,N_4885);
nor UO_292 (O_292,N_4928,N_4920);
nor UO_293 (O_293,N_4967,N_4916);
or UO_294 (O_294,N_4965,N_4993);
nor UO_295 (O_295,N_4939,N_4834);
and UO_296 (O_296,N_4991,N_4975);
nand UO_297 (O_297,N_4823,N_4901);
or UO_298 (O_298,N_4834,N_4938);
and UO_299 (O_299,N_4905,N_4814);
or UO_300 (O_300,N_4858,N_4907);
nor UO_301 (O_301,N_4817,N_4919);
and UO_302 (O_302,N_4870,N_4909);
or UO_303 (O_303,N_4903,N_4867);
or UO_304 (O_304,N_4813,N_4886);
nor UO_305 (O_305,N_4831,N_4915);
nor UO_306 (O_306,N_4926,N_4983);
or UO_307 (O_307,N_4809,N_4872);
nor UO_308 (O_308,N_4803,N_4904);
and UO_309 (O_309,N_4921,N_4898);
nand UO_310 (O_310,N_4971,N_4965);
nand UO_311 (O_311,N_4912,N_4987);
or UO_312 (O_312,N_4924,N_4849);
nand UO_313 (O_313,N_4848,N_4925);
and UO_314 (O_314,N_4842,N_4990);
and UO_315 (O_315,N_4869,N_4909);
nand UO_316 (O_316,N_4963,N_4851);
and UO_317 (O_317,N_4998,N_4843);
nor UO_318 (O_318,N_4886,N_4881);
nor UO_319 (O_319,N_4880,N_4963);
nor UO_320 (O_320,N_4942,N_4813);
nand UO_321 (O_321,N_4890,N_4882);
or UO_322 (O_322,N_4830,N_4996);
nor UO_323 (O_323,N_4914,N_4849);
or UO_324 (O_324,N_4801,N_4915);
nor UO_325 (O_325,N_4887,N_4998);
nand UO_326 (O_326,N_4827,N_4862);
nor UO_327 (O_327,N_4906,N_4894);
or UO_328 (O_328,N_4985,N_4827);
and UO_329 (O_329,N_4828,N_4891);
nand UO_330 (O_330,N_4996,N_4916);
and UO_331 (O_331,N_4983,N_4867);
and UO_332 (O_332,N_4895,N_4948);
and UO_333 (O_333,N_4922,N_4949);
nand UO_334 (O_334,N_4937,N_4967);
nand UO_335 (O_335,N_4956,N_4809);
or UO_336 (O_336,N_4948,N_4870);
nand UO_337 (O_337,N_4937,N_4946);
nand UO_338 (O_338,N_4923,N_4853);
nand UO_339 (O_339,N_4804,N_4918);
and UO_340 (O_340,N_4942,N_4997);
nand UO_341 (O_341,N_4967,N_4949);
nand UO_342 (O_342,N_4982,N_4927);
nor UO_343 (O_343,N_4805,N_4921);
nor UO_344 (O_344,N_4894,N_4970);
nand UO_345 (O_345,N_4867,N_4830);
nand UO_346 (O_346,N_4912,N_4874);
nand UO_347 (O_347,N_4838,N_4907);
or UO_348 (O_348,N_4812,N_4922);
or UO_349 (O_349,N_4995,N_4892);
nor UO_350 (O_350,N_4893,N_4973);
or UO_351 (O_351,N_4983,N_4842);
and UO_352 (O_352,N_4922,N_4991);
nand UO_353 (O_353,N_4809,N_4890);
and UO_354 (O_354,N_4843,N_4829);
and UO_355 (O_355,N_4914,N_4909);
nand UO_356 (O_356,N_4956,N_4957);
and UO_357 (O_357,N_4831,N_4920);
or UO_358 (O_358,N_4900,N_4942);
or UO_359 (O_359,N_4873,N_4828);
nor UO_360 (O_360,N_4933,N_4881);
or UO_361 (O_361,N_4928,N_4879);
nand UO_362 (O_362,N_4889,N_4896);
nor UO_363 (O_363,N_4800,N_4857);
nand UO_364 (O_364,N_4943,N_4989);
and UO_365 (O_365,N_4872,N_4898);
nor UO_366 (O_366,N_4995,N_4881);
or UO_367 (O_367,N_4805,N_4941);
nor UO_368 (O_368,N_4964,N_4823);
nand UO_369 (O_369,N_4880,N_4854);
nor UO_370 (O_370,N_4993,N_4880);
and UO_371 (O_371,N_4876,N_4937);
or UO_372 (O_372,N_4950,N_4980);
nand UO_373 (O_373,N_4827,N_4885);
nor UO_374 (O_374,N_4965,N_4873);
nor UO_375 (O_375,N_4831,N_4972);
or UO_376 (O_376,N_4895,N_4801);
or UO_377 (O_377,N_4937,N_4827);
nor UO_378 (O_378,N_4851,N_4810);
nand UO_379 (O_379,N_4923,N_4914);
nor UO_380 (O_380,N_4910,N_4936);
nand UO_381 (O_381,N_4859,N_4833);
or UO_382 (O_382,N_4981,N_4924);
nand UO_383 (O_383,N_4823,N_4972);
and UO_384 (O_384,N_4814,N_4835);
nand UO_385 (O_385,N_4929,N_4908);
and UO_386 (O_386,N_4821,N_4964);
xnor UO_387 (O_387,N_4940,N_4948);
nand UO_388 (O_388,N_4883,N_4935);
nor UO_389 (O_389,N_4873,N_4810);
or UO_390 (O_390,N_4859,N_4901);
nor UO_391 (O_391,N_4818,N_4996);
nand UO_392 (O_392,N_4902,N_4957);
nand UO_393 (O_393,N_4985,N_4845);
and UO_394 (O_394,N_4913,N_4828);
or UO_395 (O_395,N_4804,N_4809);
or UO_396 (O_396,N_4857,N_4951);
or UO_397 (O_397,N_4813,N_4964);
nand UO_398 (O_398,N_4811,N_4954);
nor UO_399 (O_399,N_4957,N_4951);
nor UO_400 (O_400,N_4998,N_4940);
and UO_401 (O_401,N_4846,N_4996);
or UO_402 (O_402,N_4972,N_4818);
or UO_403 (O_403,N_4928,N_4946);
nand UO_404 (O_404,N_4808,N_4935);
nor UO_405 (O_405,N_4962,N_4830);
and UO_406 (O_406,N_4814,N_4817);
nand UO_407 (O_407,N_4878,N_4985);
nand UO_408 (O_408,N_4888,N_4823);
nand UO_409 (O_409,N_4969,N_4984);
nor UO_410 (O_410,N_4839,N_4821);
nand UO_411 (O_411,N_4807,N_4851);
xor UO_412 (O_412,N_4974,N_4834);
nand UO_413 (O_413,N_4839,N_4998);
nor UO_414 (O_414,N_4951,N_4937);
nor UO_415 (O_415,N_4806,N_4984);
nor UO_416 (O_416,N_4826,N_4872);
and UO_417 (O_417,N_4952,N_4939);
xnor UO_418 (O_418,N_4885,N_4935);
and UO_419 (O_419,N_4878,N_4969);
nand UO_420 (O_420,N_4982,N_4976);
and UO_421 (O_421,N_4879,N_4846);
nand UO_422 (O_422,N_4893,N_4966);
and UO_423 (O_423,N_4946,N_4879);
and UO_424 (O_424,N_4875,N_4989);
nor UO_425 (O_425,N_4809,N_4843);
or UO_426 (O_426,N_4988,N_4890);
nor UO_427 (O_427,N_4848,N_4804);
and UO_428 (O_428,N_4850,N_4951);
nand UO_429 (O_429,N_4887,N_4875);
nand UO_430 (O_430,N_4899,N_4873);
nor UO_431 (O_431,N_4851,N_4857);
nand UO_432 (O_432,N_4848,N_4918);
or UO_433 (O_433,N_4978,N_4876);
or UO_434 (O_434,N_4809,N_4813);
and UO_435 (O_435,N_4988,N_4834);
or UO_436 (O_436,N_4996,N_4912);
or UO_437 (O_437,N_4998,N_4860);
nor UO_438 (O_438,N_4959,N_4979);
and UO_439 (O_439,N_4821,N_4978);
or UO_440 (O_440,N_4990,N_4826);
and UO_441 (O_441,N_4857,N_4945);
nor UO_442 (O_442,N_4849,N_4903);
nand UO_443 (O_443,N_4974,N_4903);
and UO_444 (O_444,N_4877,N_4937);
nand UO_445 (O_445,N_4965,N_4979);
nand UO_446 (O_446,N_4871,N_4862);
nor UO_447 (O_447,N_4890,N_4830);
nor UO_448 (O_448,N_4847,N_4881);
nand UO_449 (O_449,N_4999,N_4822);
and UO_450 (O_450,N_4912,N_4984);
nand UO_451 (O_451,N_4808,N_4882);
or UO_452 (O_452,N_4818,N_4807);
and UO_453 (O_453,N_4820,N_4819);
and UO_454 (O_454,N_4854,N_4910);
nand UO_455 (O_455,N_4882,N_4933);
or UO_456 (O_456,N_4814,N_4900);
nor UO_457 (O_457,N_4815,N_4852);
or UO_458 (O_458,N_4921,N_4988);
and UO_459 (O_459,N_4953,N_4916);
nand UO_460 (O_460,N_4907,N_4885);
nand UO_461 (O_461,N_4977,N_4893);
nand UO_462 (O_462,N_4980,N_4967);
or UO_463 (O_463,N_4805,N_4964);
and UO_464 (O_464,N_4835,N_4840);
nor UO_465 (O_465,N_4998,N_4999);
or UO_466 (O_466,N_4895,N_4860);
or UO_467 (O_467,N_4870,N_4887);
nor UO_468 (O_468,N_4967,N_4884);
and UO_469 (O_469,N_4817,N_4947);
nor UO_470 (O_470,N_4857,N_4825);
and UO_471 (O_471,N_4821,N_4959);
or UO_472 (O_472,N_4921,N_4849);
and UO_473 (O_473,N_4856,N_4833);
or UO_474 (O_474,N_4847,N_4837);
and UO_475 (O_475,N_4949,N_4902);
nand UO_476 (O_476,N_4930,N_4885);
nand UO_477 (O_477,N_4988,N_4813);
and UO_478 (O_478,N_4908,N_4891);
and UO_479 (O_479,N_4925,N_4821);
nand UO_480 (O_480,N_4957,N_4943);
nand UO_481 (O_481,N_4888,N_4872);
and UO_482 (O_482,N_4833,N_4918);
or UO_483 (O_483,N_4889,N_4999);
xor UO_484 (O_484,N_4806,N_4947);
or UO_485 (O_485,N_4852,N_4885);
nand UO_486 (O_486,N_4974,N_4939);
and UO_487 (O_487,N_4944,N_4994);
nor UO_488 (O_488,N_4973,N_4821);
nor UO_489 (O_489,N_4829,N_4956);
nand UO_490 (O_490,N_4902,N_4976);
or UO_491 (O_491,N_4959,N_4927);
or UO_492 (O_492,N_4977,N_4961);
xor UO_493 (O_493,N_4828,N_4884);
nor UO_494 (O_494,N_4993,N_4934);
or UO_495 (O_495,N_4893,N_4897);
and UO_496 (O_496,N_4979,N_4956);
or UO_497 (O_497,N_4882,N_4956);
or UO_498 (O_498,N_4852,N_4993);
or UO_499 (O_499,N_4836,N_4891);
nand UO_500 (O_500,N_4932,N_4997);
nor UO_501 (O_501,N_4805,N_4980);
nand UO_502 (O_502,N_4864,N_4825);
or UO_503 (O_503,N_4802,N_4929);
or UO_504 (O_504,N_4820,N_4909);
nand UO_505 (O_505,N_4965,N_4927);
or UO_506 (O_506,N_4855,N_4971);
nor UO_507 (O_507,N_4889,N_4934);
and UO_508 (O_508,N_4980,N_4865);
and UO_509 (O_509,N_4946,N_4921);
nor UO_510 (O_510,N_4875,N_4866);
xor UO_511 (O_511,N_4855,N_4979);
nor UO_512 (O_512,N_4834,N_4906);
nor UO_513 (O_513,N_4969,N_4807);
nor UO_514 (O_514,N_4877,N_4899);
nand UO_515 (O_515,N_4886,N_4811);
nor UO_516 (O_516,N_4865,N_4800);
nand UO_517 (O_517,N_4919,N_4884);
or UO_518 (O_518,N_4941,N_4952);
nand UO_519 (O_519,N_4992,N_4919);
or UO_520 (O_520,N_4803,N_4893);
and UO_521 (O_521,N_4847,N_4900);
nor UO_522 (O_522,N_4899,N_4930);
and UO_523 (O_523,N_4973,N_4811);
or UO_524 (O_524,N_4904,N_4839);
or UO_525 (O_525,N_4869,N_4926);
and UO_526 (O_526,N_4937,N_4833);
and UO_527 (O_527,N_4844,N_4913);
nand UO_528 (O_528,N_4901,N_4841);
nand UO_529 (O_529,N_4944,N_4909);
nor UO_530 (O_530,N_4884,N_4870);
or UO_531 (O_531,N_4840,N_4979);
nand UO_532 (O_532,N_4847,N_4923);
or UO_533 (O_533,N_4838,N_4888);
nand UO_534 (O_534,N_4890,N_4807);
or UO_535 (O_535,N_4930,N_4886);
nor UO_536 (O_536,N_4906,N_4890);
or UO_537 (O_537,N_4987,N_4831);
nand UO_538 (O_538,N_4916,N_4878);
and UO_539 (O_539,N_4938,N_4804);
xor UO_540 (O_540,N_4863,N_4850);
or UO_541 (O_541,N_4981,N_4863);
or UO_542 (O_542,N_4843,N_4835);
or UO_543 (O_543,N_4864,N_4820);
and UO_544 (O_544,N_4982,N_4945);
nor UO_545 (O_545,N_4933,N_4894);
and UO_546 (O_546,N_4949,N_4979);
nand UO_547 (O_547,N_4923,N_4985);
or UO_548 (O_548,N_4981,N_4815);
nor UO_549 (O_549,N_4828,N_4905);
and UO_550 (O_550,N_4919,N_4947);
and UO_551 (O_551,N_4895,N_4861);
or UO_552 (O_552,N_4838,N_4968);
nand UO_553 (O_553,N_4914,N_4922);
and UO_554 (O_554,N_4932,N_4841);
nor UO_555 (O_555,N_4996,N_4885);
nand UO_556 (O_556,N_4829,N_4863);
and UO_557 (O_557,N_4886,N_4956);
or UO_558 (O_558,N_4849,N_4857);
and UO_559 (O_559,N_4895,N_4933);
or UO_560 (O_560,N_4917,N_4972);
nand UO_561 (O_561,N_4802,N_4898);
or UO_562 (O_562,N_4980,N_4848);
or UO_563 (O_563,N_4855,N_4986);
and UO_564 (O_564,N_4995,N_4959);
and UO_565 (O_565,N_4899,N_4993);
or UO_566 (O_566,N_4946,N_4801);
nand UO_567 (O_567,N_4894,N_4833);
and UO_568 (O_568,N_4812,N_4911);
nor UO_569 (O_569,N_4923,N_4964);
nor UO_570 (O_570,N_4810,N_4985);
and UO_571 (O_571,N_4878,N_4960);
nand UO_572 (O_572,N_4989,N_4974);
nor UO_573 (O_573,N_4832,N_4816);
or UO_574 (O_574,N_4966,N_4885);
and UO_575 (O_575,N_4801,N_4813);
and UO_576 (O_576,N_4823,N_4800);
and UO_577 (O_577,N_4993,N_4996);
nand UO_578 (O_578,N_4803,N_4916);
or UO_579 (O_579,N_4943,N_4995);
nand UO_580 (O_580,N_4962,N_4808);
nor UO_581 (O_581,N_4818,N_4835);
nand UO_582 (O_582,N_4856,N_4955);
and UO_583 (O_583,N_4993,N_4957);
and UO_584 (O_584,N_4945,N_4937);
nand UO_585 (O_585,N_4969,N_4847);
or UO_586 (O_586,N_4855,N_4836);
nand UO_587 (O_587,N_4888,N_4911);
nand UO_588 (O_588,N_4844,N_4863);
and UO_589 (O_589,N_4926,N_4856);
nor UO_590 (O_590,N_4881,N_4832);
or UO_591 (O_591,N_4916,N_4933);
or UO_592 (O_592,N_4809,N_4894);
nand UO_593 (O_593,N_4915,N_4821);
and UO_594 (O_594,N_4847,N_4815);
or UO_595 (O_595,N_4902,N_4845);
nand UO_596 (O_596,N_4912,N_4993);
or UO_597 (O_597,N_4910,N_4883);
nor UO_598 (O_598,N_4928,N_4818);
xnor UO_599 (O_599,N_4811,N_4841);
nor UO_600 (O_600,N_4896,N_4920);
nand UO_601 (O_601,N_4966,N_4959);
nor UO_602 (O_602,N_4859,N_4873);
and UO_603 (O_603,N_4951,N_4955);
and UO_604 (O_604,N_4925,N_4895);
nor UO_605 (O_605,N_4984,N_4813);
nor UO_606 (O_606,N_4918,N_4982);
and UO_607 (O_607,N_4947,N_4878);
nor UO_608 (O_608,N_4815,N_4854);
and UO_609 (O_609,N_4882,N_4869);
and UO_610 (O_610,N_4855,N_4858);
nand UO_611 (O_611,N_4877,N_4913);
nand UO_612 (O_612,N_4829,N_4968);
nand UO_613 (O_613,N_4844,N_4936);
nand UO_614 (O_614,N_4843,N_4916);
nand UO_615 (O_615,N_4962,N_4977);
nor UO_616 (O_616,N_4990,N_4800);
xor UO_617 (O_617,N_4830,N_4946);
nand UO_618 (O_618,N_4938,N_4952);
and UO_619 (O_619,N_4975,N_4950);
nand UO_620 (O_620,N_4883,N_4825);
and UO_621 (O_621,N_4994,N_4920);
nand UO_622 (O_622,N_4884,N_4822);
nand UO_623 (O_623,N_4897,N_4901);
or UO_624 (O_624,N_4996,N_4812);
or UO_625 (O_625,N_4994,N_4977);
nand UO_626 (O_626,N_4955,N_4847);
and UO_627 (O_627,N_4808,N_4854);
nand UO_628 (O_628,N_4836,N_4853);
nor UO_629 (O_629,N_4955,N_4833);
nand UO_630 (O_630,N_4977,N_4844);
nor UO_631 (O_631,N_4906,N_4911);
and UO_632 (O_632,N_4912,N_4864);
nor UO_633 (O_633,N_4826,N_4980);
and UO_634 (O_634,N_4821,N_4921);
or UO_635 (O_635,N_4847,N_4870);
or UO_636 (O_636,N_4979,N_4862);
nor UO_637 (O_637,N_4873,N_4812);
nand UO_638 (O_638,N_4919,N_4886);
and UO_639 (O_639,N_4841,N_4825);
or UO_640 (O_640,N_4812,N_4833);
nor UO_641 (O_641,N_4830,N_4904);
nor UO_642 (O_642,N_4976,N_4812);
and UO_643 (O_643,N_4835,N_4880);
nor UO_644 (O_644,N_4944,N_4827);
or UO_645 (O_645,N_4856,N_4845);
nand UO_646 (O_646,N_4857,N_4871);
xor UO_647 (O_647,N_4956,N_4895);
and UO_648 (O_648,N_4973,N_4877);
or UO_649 (O_649,N_4910,N_4988);
or UO_650 (O_650,N_4846,N_4821);
or UO_651 (O_651,N_4850,N_4846);
nor UO_652 (O_652,N_4963,N_4807);
nand UO_653 (O_653,N_4859,N_4806);
and UO_654 (O_654,N_4936,N_4878);
nor UO_655 (O_655,N_4965,N_4811);
and UO_656 (O_656,N_4956,N_4936);
nor UO_657 (O_657,N_4946,N_4999);
nand UO_658 (O_658,N_4880,N_4834);
and UO_659 (O_659,N_4840,N_4951);
and UO_660 (O_660,N_4953,N_4849);
nand UO_661 (O_661,N_4923,N_4958);
and UO_662 (O_662,N_4977,N_4814);
and UO_663 (O_663,N_4867,N_4943);
nand UO_664 (O_664,N_4930,N_4871);
nor UO_665 (O_665,N_4989,N_4818);
and UO_666 (O_666,N_4854,N_4944);
nor UO_667 (O_667,N_4890,N_4933);
nor UO_668 (O_668,N_4878,N_4942);
and UO_669 (O_669,N_4956,N_4942);
and UO_670 (O_670,N_4814,N_4920);
or UO_671 (O_671,N_4855,N_4842);
nor UO_672 (O_672,N_4826,N_4822);
nor UO_673 (O_673,N_4915,N_4818);
or UO_674 (O_674,N_4879,N_4914);
and UO_675 (O_675,N_4946,N_4994);
xnor UO_676 (O_676,N_4905,N_4887);
nor UO_677 (O_677,N_4821,N_4814);
or UO_678 (O_678,N_4936,N_4998);
nand UO_679 (O_679,N_4900,N_4981);
nor UO_680 (O_680,N_4813,N_4811);
and UO_681 (O_681,N_4908,N_4902);
nand UO_682 (O_682,N_4825,N_4866);
and UO_683 (O_683,N_4879,N_4985);
and UO_684 (O_684,N_4938,N_4891);
nor UO_685 (O_685,N_4937,N_4911);
nor UO_686 (O_686,N_4843,N_4917);
and UO_687 (O_687,N_4982,N_4923);
and UO_688 (O_688,N_4855,N_4923);
nand UO_689 (O_689,N_4819,N_4896);
and UO_690 (O_690,N_4811,N_4804);
nor UO_691 (O_691,N_4919,N_4815);
or UO_692 (O_692,N_4835,N_4975);
nand UO_693 (O_693,N_4903,N_4896);
and UO_694 (O_694,N_4815,N_4895);
nand UO_695 (O_695,N_4971,N_4822);
and UO_696 (O_696,N_4969,N_4832);
nor UO_697 (O_697,N_4847,N_4862);
and UO_698 (O_698,N_4838,N_4989);
nand UO_699 (O_699,N_4964,N_4982);
or UO_700 (O_700,N_4925,N_4914);
nor UO_701 (O_701,N_4815,N_4937);
or UO_702 (O_702,N_4875,N_4862);
nor UO_703 (O_703,N_4956,N_4876);
and UO_704 (O_704,N_4941,N_4914);
nand UO_705 (O_705,N_4984,N_4990);
nand UO_706 (O_706,N_4994,N_4859);
nand UO_707 (O_707,N_4806,N_4895);
nor UO_708 (O_708,N_4859,N_4899);
or UO_709 (O_709,N_4932,N_4902);
and UO_710 (O_710,N_4889,N_4970);
and UO_711 (O_711,N_4870,N_4822);
nor UO_712 (O_712,N_4809,N_4880);
nor UO_713 (O_713,N_4981,N_4804);
nor UO_714 (O_714,N_4919,N_4942);
or UO_715 (O_715,N_4922,N_4920);
nor UO_716 (O_716,N_4828,N_4943);
nor UO_717 (O_717,N_4953,N_4902);
or UO_718 (O_718,N_4998,N_4942);
and UO_719 (O_719,N_4889,N_4832);
or UO_720 (O_720,N_4914,N_4865);
nand UO_721 (O_721,N_4875,N_4847);
nand UO_722 (O_722,N_4937,N_4932);
or UO_723 (O_723,N_4987,N_4872);
nor UO_724 (O_724,N_4834,N_4983);
or UO_725 (O_725,N_4908,N_4989);
and UO_726 (O_726,N_4850,N_4840);
or UO_727 (O_727,N_4804,N_4853);
or UO_728 (O_728,N_4945,N_4899);
or UO_729 (O_729,N_4852,N_4978);
nor UO_730 (O_730,N_4818,N_4952);
nor UO_731 (O_731,N_4900,N_4804);
nand UO_732 (O_732,N_4980,N_4948);
nand UO_733 (O_733,N_4833,N_4974);
nor UO_734 (O_734,N_4992,N_4817);
nor UO_735 (O_735,N_4840,N_4865);
xor UO_736 (O_736,N_4979,N_4988);
nand UO_737 (O_737,N_4879,N_4986);
nor UO_738 (O_738,N_4945,N_4979);
xnor UO_739 (O_739,N_4883,N_4821);
and UO_740 (O_740,N_4926,N_4928);
or UO_741 (O_741,N_4950,N_4801);
nand UO_742 (O_742,N_4956,N_4949);
and UO_743 (O_743,N_4862,N_4825);
nand UO_744 (O_744,N_4926,N_4838);
xnor UO_745 (O_745,N_4813,N_4980);
and UO_746 (O_746,N_4817,N_4936);
nand UO_747 (O_747,N_4885,N_4927);
nand UO_748 (O_748,N_4837,N_4843);
nand UO_749 (O_749,N_4996,N_4980);
or UO_750 (O_750,N_4969,N_4820);
and UO_751 (O_751,N_4924,N_4844);
xor UO_752 (O_752,N_4905,N_4999);
or UO_753 (O_753,N_4943,N_4924);
nand UO_754 (O_754,N_4976,N_4893);
or UO_755 (O_755,N_4918,N_4925);
nand UO_756 (O_756,N_4829,N_4965);
and UO_757 (O_757,N_4843,N_4939);
and UO_758 (O_758,N_4846,N_4921);
nand UO_759 (O_759,N_4887,N_4820);
nor UO_760 (O_760,N_4898,N_4877);
nor UO_761 (O_761,N_4867,N_4970);
nor UO_762 (O_762,N_4958,N_4991);
nand UO_763 (O_763,N_4926,N_4860);
or UO_764 (O_764,N_4859,N_4841);
or UO_765 (O_765,N_4824,N_4813);
nor UO_766 (O_766,N_4879,N_4932);
or UO_767 (O_767,N_4860,N_4859);
or UO_768 (O_768,N_4934,N_4922);
or UO_769 (O_769,N_4970,N_4914);
and UO_770 (O_770,N_4985,N_4988);
xnor UO_771 (O_771,N_4814,N_4957);
and UO_772 (O_772,N_4845,N_4942);
nor UO_773 (O_773,N_4899,N_4837);
or UO_774 (O_774,N_4806,N_4841);
xnor UO_775 (O_775,N_4897,N_4826);
and UO_776 (O_776,N_4917,N_4882);
or UO_777 (O_777,N_4888,N_4977);
and UO_778 (O_778,N_4877,N_4953);
nand UO_779 (O_779,N_4851,N_4927);
nor UO_780 (O_780,N_4836,N_4938);
nor UO_781 (O_781,N_4820,N_4891);
and UO_782 (O_782,N_4965,N_4953);
or UO_783 (O_783,N_4943,N_4823);
nand UO_784 (O_784,N_4839,N_4845);
or UO_785 (O_785,N_4833,N_4938);
nand UO_786 (O_786,N_4816,N_4912);
nand UO_787 (O_787,N_4977,N_4827);
nand UO_788 (O_788,N_4892,N_4935);
or UO_789 (O_789,N_4839,N_4986);
and UO_790 (O_790,N_4877,N_4892);
nor UO_791 (O_791,N_4960,N_4847);
and UO_792 (O_792,N_4916,N_4870);
nand UO_793 (O_793,N_4942,N_4825);
and UO_794 (O_794,N_4978,N_4918);
nor UO_795 (O_795,N_4985,N_4965);
or UO_796 (O_796,N_4938,N_4843);
and UO_797 (O_797,N_4931,N_4872);
or UO_798 (O_798,N_4859,N_4852);
or UO_799 (O_799,N_4861,N_4973);
nand UO_800 (O_800,N_4843,N_4958);
nand UO_801 (O_801,N_4958,N_4824);
and UO_802 (O_802,N_4975,N_4815);
and UO_803 (O_803,N_4960,N_4812);
or UO_804 (O_804,N_4828,N_4993);
nor UO_805 (O_805,N_4995,N_4950);
xnor UO_806 (O_806,N_4921,N_4963);
nor UO_807 (O_807,N_4950,N_4942);
nor UO_808 (O_808,N_4858,N_4986);
or UO_809 (O_809,N_4975,N_4953);
nand UO_810 (O_810,N_4905,N_4942);
nor UO_811 (O_811,N_4914,N_4951);
nor UO_812 (O_812,N_4843,N_4919);
nand UO_813 (O_813,N_4837,N_4959);
nand UO_814 (O_814,N_4848,N_4937);
nand UO_815 (O_815,N_4956,N_4888);
or UO_816 (O_816,N_4954,N_4850);
nor UO_817 (O_817,N_4990,N_4843);
or UO_818 (O_818,N_4898,N_4996);
and UO_819 (O_819,N_4829,N_4847);
nand UO_820 (O_820,N_4921,N_4909);
and UO_821 (O_821,N_4963,N_4801);
nor UO_822 (O_822,N_4943,N_4816);
nor UO_823 (O_823,N_4937,N_4871);
and UO_824 (O_824,N_4979,N_4964);
or UO_825 (O_825,N_4920,N_4904);
nand UO_826 (O_826,N_4934,N_4894);
nand UO_827 (O_827,N_4913,N_4839);
and UO_828 (O_828,N_4909,N_4831);
and UO_829 (O_829,N_4820,N_4810);
or UO_830 (O_830,N_4989,N_4957);
or UO_831 (O_831,N_4996,N_4880);
nor UO_832 (O_832,N_4949,N_4839);
nor UO_833 (O_833,N_4885,N_4893);
or UO_834 (O_834,N_4955,N_4937);
or UO_835 (O_835,N_4856,N_4804);
nand UO_836 (O_836,N_4812,N_4845);
nor UO_837 (O_837,N_4809,N_4851);
nor UO_838 (O_838,N_4947,N_4839);
xnor UO_839 (O_839,N_4954,N_4862);
xor UO_840 (O_840,N_4810,N_4845);
nor UO_841 (O_841,N_4806,N_4810);
nand UO_842 (O_842,N_4974,N_4873);
nor UO_843 (O_843,N_4936,N_4917);
nand UO_844 (O_844,N_4899,N_4909);
nand UO_845 (O_845,N_4871,N_4845);
nor UO_846 (O_846,N_4967,N_4981);
nor UO_847 (O_847,N_4983,N_4818);
or UO_848 (O_848,N_4948,N_4814);
nor UO_849 (O_849,N_4815,N_4820);
and UO_850 (O_850,N_4956,N_4985);
or UO_851 (O_851,N_4889,N_4810);
and UO_852 (O_852,N_4887,N_4921);
nand UO_853 (O_853,N_4878,N_4876);
or UO_854 (O_854,N_4953,N_4838);
nand UO_855 (O_855,N_4895,N_4982);
nor UO_856 (O_856,N_4997,N_4857);
nand UO_857 (O_857,N_4931,N_4819);
or UO_858 (O_858,N_4984,N_4927);
nor UO_859 (O_859,N_4949,N_4831);
nand UO_860 (O_860,N_4809,N_4996);
or UO_861 (O_861,N_4820,N_4880);
nor UO_862 (O_862,N_4939,N_4830);
or UO_863 (O_863,N_4971,N_4884);
and UO_864 (O_864,N_4854,N_4898);
or UO_865 (O_865,N_4844,N_4906);
and UO_866 (O_866,N_4853,N_4848);
xor UO_867 (O_867,N_4962,N_4950);
or UO_868 (O_868,N_4947,N_4831);
and UO_869 (O_869,N_4810,N_4979);
or UO_870 (O_870,N_4951,N_4875);
or UO_871 (O_871,N_4815,N_4842);
and UO_872 (O_872,N_4906,N_4835);
or UO_873 (O_873,N_4956,N_4822);
or UO_874 (O_874,N_4862,N_4963);
and UO_875 (O_875,N_4825,N_4829);
and UO_876 (O_876,N_4835,N_4823);
or UO_877 (O_877,N_4870,N_4877);
nor UO_878 (O_878,N_4996,N_4804);
and UO_879 (O_879,N_4909,N_4962);
nand UO_880 (O_880,N_4806,N_4816);
nor UO_881 (O_881,N_4868,N_4949);
nand UO_882 (O_882,N_4944,N_4996);
or UO_883 (O_883,N_4866,N_4958);
nand UO_884 (O_884,N_4909,N_4994);
nor UO_885 (O_885,N_4847,N_4944);
nor UO_886 (O_886,N_4976,N_4896);
nand UO_887 (O_887,N_4935,N_4939);
xnor UO_888 (O_888,N_4828,N_4860);
and UO_889 (O_889,N_4876,N_4942);
or UO_890 (O_890,N_4854,N_4800);
or UO_891 (O_891,N_4892,N_4968);
nand UO_892 (O_892,N_4905,N_4842);
and UO_893 (O_893,N_4878,N_4818);
and UO_894 (O_894,N_4816,N_4941);
xor UO_895 (O_895,N_4952,N_4962);
nand UO_896 (O_896,N_4932,N_4970);
and UO_897 (O_897,N_4995,N_4830);
nand UO_898 (O_898,N_4812,N_4965);
nand UO_899 (O_899,N_4955,N_4992);
nand UO_900 (O_900,N_4805,N_4817);
or UO_901 (O_901,N_4894,N_4922);
nand UO_902 (O_902,N_4804,N_4852);
and UO_903 (O_903,N_4825,N_4824);
and UO_904 (O_904,N_4856,N_4941);
and UO_905 (O_905,N_4932,N_4829);
and UO_906 (O_906,N_4877,N_4805);
or UO_907 (O_907,N_4977,N_4972);
or UO_908 (O_908,N_4929,N_4980);
nand UO_909 (O_909,N_4894,N_4971);
or UO_910 (O_910,N_4810,N_4868);
and UO_911 (O_911,N_4850,N_4833);
nor UO_912 (O_912,N_4971,N_4821);
or UO_913 (O_913,N_4978,N_4921);
nor UO_914 (O_914,N_4890,N_4972);
nand UO_915 (O_915,N_4986,N_4913);
or UO_916 (O_916,N_4879,N_4849);
and UO_917 (O_917,N_4969,N_4853);
nand UO_918 (O_918,N_4830,N_4934);
and UO_919 (O_919,N_4882,N_4888);
and UO_920 (O_920,N_4960,N_4975);
nor UO_921 (O_921,N_4884,N_4897);
nand UO_922 (O_922,N_4901,N_4819);
nand UO_923 (O_923,N_4883,N_4865);
or UO_924 (O_924,N_4803,N_4802);
and UO_925 (O_925,N_4982,N_4879);
or UO_926 (O_926,N_4946,N_4939);
and UO_927 (O_927,N_4955,N_4814);
nand UO_928 (O_928,N_4848,N_4861);
or UO_929 (O_929,N_4883,N_4996);
nor UO_930 (O_930,N_4997,N_4955);
and UO_931 (O_931,N_4810,N_4941);
or UO_932 (O_932,N_4815,N_4883);
and UO_933 (O_933,N_4889,N_4930);
nor UO_934 (O_934,N_4866,N_4803);
nand UO_935 (O_935,N_4866,N_4939);
nand UO_936 (O_936,N_4982,N_4861);
or UO_937 (O_937,N_4908,N_4932);
xnor UO_938 (O_938,N_4878,N_4988);
nor UO_939 (O_939,N_4963,N_4947);
nand UO_940 (O_940,N_4983,N_4839);
nand UO_941 (O_941,N_4974,N_4997);
or UO_942 (O_942,N_4834,N_4930);
or UO_943 (O_943,N_4928,N_4832);
and UO_944 (O_944,N_4938,N_4959);
nand UO_945 (O_945,N_4807,N_4974);
nand UO_946 (O_946,N_4963,N_4956);
and UO_947 (O_947,N_4829,N_4926);
nand UO_948 (O_948,N_4884,N_4977);
nand UO_949 (O_949,N_4890,N_4949);
and UO_950 (O_950,N_4964,N_4929);
nand UO_951 (O_951,N_4866,N_4926);
nor UO_952 (O_952,N_4843,N_4877);
xnor UO_953 (O_953,N_4916,N_4812);
or UO_954 (O_954,N_4803,N_4962);
nand UO_955 (O_955,N_4915,N_4975);
nor UO_956 (O_956,N_4835,N_4930);
and UO_957 (O_957,N_4928,N_4942);
nor UO_958 (O_958,N_4877,N_4823);
and UO_959 (O_959,N_4885,N_4942);
nand UO_960 (O_960,N_4877,N_4821);
or UO_961 (O_961,N_4851,N_4849);
xor UO_962 (O_962,N_4978,N_4952);
or UO_963 (O_963,N_4878,N_4802);
xor UO_964 (O_964,N_4888,N_4841);
nand UO_965 (O_965,N_4905,N_4839);
or UO_966 (O_966,N_4905,N_4850);
or UO_967 (O_967,N_4838,N_4925);
or UO_968 (O_968,N_4913,N_4835);
xor UO_969 (O_969,N_4847,N_4964);
or UO_970 (O_970,N_4998,N_4997);
and UO_971 (O_971,N_4867,N_4961);
or UO_972 (O_972,N_4819,N_4833);
nand UO_973 (O_973,N_4928,N_4938);
nand UO_974 (O_974,N_4981,N_4800);
or UO_975 (O_975,N_4905,N_4979);
nor UO_976 (O_976,N_4865,N_4867);
nor UO_977 (O_977,N_4803,N_4845);
and UO_978 (O_978,N_4822,N_4850);
xnor UO_979 (O_979,N_4846,N_4851);
and UO_980 (O_980,N_4893,N_4819);
or UO_981 (O_981,N_4891,N_4894);
nor UO_982 (O_982,N_4982,N_4837);
or UO_983 (O_983,N_4934,N_4970);
nand UO_984 (O_984,N_4992,N_4946);
or UO_985 (O_985,N_4869,N_4886);
nor UO_986 (O_986,N_4908,N_4834);
or UO_987 (O_987,N_4859,N_4997);
or UO_988 (O_988,N_4894,N_4908);
nand UO_989 (O_989,N_4872,N_4929);
nor UO_990 (O_990,N_4864,N_4826);
and UO_991 (O_991,N_4984,N_4861);
nor UO_992 (O_992,N_4934,N_4947);
xor UO_993 (O_993,N_4822,N_4886);
and UO_994 (O_994,N_4809,N_4936);
or UO_995 (O_995,N_4837,N_4925);
nor UO_996 (O_996,N_4951,N_4918);
and UO_997 (O_997,N_4879,N_4828);
xor UO_998 (O_998,N_4849,N_4843);
nor UO_999 (O_999,N_4910,N_4979);
endmodule