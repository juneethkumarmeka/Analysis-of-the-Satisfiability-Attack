module basic_500_3000_500_40_levels_2xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_497,In_453);
nand U1 (N_1,In_486,In_162);
and U2 (N_2,In_476,In_372);
nor U3 (N_3,In_60,In_49);
or U4 (N_4,In_353,In_306);
xnor U5 (N_5,In_396,In_113);
and U6 (N_6,In_186,In_106);
and U7 (N_7,In_101,In_235);
nand U8 (N_8,In_446,In_442);
and U9 (N_9,In_490,In_339);
and U10 (N_10,In_82,In_38);
nand U11 (N_11,In_153,In_171);
nand U12 (N_12,In_105,In_359);
and U13 (N_13,In_0,In_410);
nand U14 (N_14,In_425,In_213);
or U15 (N_15,In_232,In_482);
nor U16 (N_16,In_472,In_483);
and U17 (N_17,In_237,In_36);
or U18 (N_18,In_471,In_244);
nand U19 (N_19,In_325,In_296);
and U20 (N_20,In_427,In_436);
nand U21 (N_21,In_177,In_447);
nor U22 (N_22,In_178,In_109);
or U23 (N_23,In_180,In_141);
nand U24 (N_24,In_269,In_115);
and U25 (N_25,In_161,In_110);
or U26 (N_26,In_347,In_438);
or U27 (N_27,In_48,In_418);
nor U28 (N_28,In_13,In_133);
and U29 (N_29,In_279,In_383);
nor U30 (N_30,In_64,In_228);
nor U31 (N_31,In_189,In_499);
and U32 (N_32,In_7,In_349);
and U33 (N_33,In_390,In_187);
and U34 (N_34,In_181,In_332);
or U35 (N_35,In_417,In_97);
nor U36 (N_36,In_465,In_479);
nor U37 (N_37,In_29,In_164);
and U38 (N_38,In_314,In_238);
and U39 (N_39,In_485,In_305);
and U40 (N_40,In_108,In_198);
and U41 (N_41,In_34,In_356);
and U42 (N_42,In_74,In_28);
nor U43 (N_43,In_39,In_317);
nor U44 (N_44,In_112,In_370);
nand U45 (N_45,In_3,In_464);
and U46 (N_46,In_315,In_124);
or U47 (N_47,In_58,In_489);
or U48 (N_48,In_369,In_392);
nor U49 (N_49,In_367,In_211);
nand U50 (N_50,In_365,In_413);
or U51 (N_51,In_88,In_111);
nor U52 (N_52,In_118,In_298);
or U53 (N_53,In_248,In_393);
and U54 (N_54,In_154,In_143);
or U55 (N_55,In_201,In_23);
and U56 (N_56,In_253,In_495);
or U57 (N_57,In_375,In_335);
or U58 (N_58,In_462,In_361);
or U59 (N_59,In_229,In_42);
nor U60 (N_60,In_329,In_94);
nand U61 (N_61,In_354,In_313);
nor U62 (N_62,In_160,In_146);
or U63 (N_63,In_289,In_196);
nand U64 (N_64,In_165,In_368);
and U65 (N_65,In_144,In_81);
nand U66 (N_66,In_57,In_126);
nand U67 (N_67,In_35,In_362);
nand U68 (N_68,In_131,In_15);
nor U69 (N_69,In_312,In_10);
nor U70 (N_70,In_342,In_226);
or U71 (N_71,In_333,In_318);
nor U72 (N_72,In_54,In_128);
and U73 (N_73,In_408,In_216);
nand U74 (N_74,In_307,In_348);
or U75 (N_75,In_304,In_429);
nand U76 (N_76,In_183,N_73);
or U77 (N_77,N_6,In_256);
or U78 (N_78,In_152,In_43);
or U79 (N_79,In_51,N_29);
nand U80 (N_80,N_9,In_89);
or U81 (N_81,N_53,In_84);
or U82 (N_82,In_374,In_85);
and U83 (N_83,In_72,In_340);
or U84 (N_84,In_323,N_74);
or U85 (N_85,N_49,In_364);
nand U86 (N_86,In_451,In_456);
or U87 (N_87,In_355,In_127);
or U88 (N_88,N_52,N_34);
and U89 (N_89,In_422,In_409);
or U90 (N_90,In_103,In_137);
nand U91 (N_91,N_32,In_439);
nand U92 (N_92,In_415,In_86);
nand U93 (N_93,In_378,In_437);
and U94 (N_94,In_397,In_430);
and U95 (N_95,In_249,In_431);
nor U96 (N_96,In_31,N_19);
or U97 (N_97,In_199,In_275);
nand U98 (N_98,N_25,In_241);
nand U99 (N_99,In_121,In_469);
nand U100 (N_100,In_338,In_405);
nand U101 (N_101,In_406,In_92);
nand U102 (N_102,In_322,In_252);
and U103 (N_103,In_283,In_480);
nor U104 (N_104,In_218,In_116);
nand U105 (N_105,In_208,In_292);
nor U106 (N_106,In_192,In_159);
nor U107 (N_107,In_428,In_276);
and U108 (N_108,In_475,In_40);
and U109 (N_109,In_351,In_93);
and U110 (N_110,In_387,In_231);
and U111 (N_111,N_38,In_227);
or U112 (N_112,In_247,In_386);
and U113 (N_113,In_260,In_225);
nand U114 (N_114,In_287,In_280);
and U115 (N_115,In_360,In_388);
or U116 (N_116,In_179,In_267);
nand U117 (N_117,In_440,In_481);
nand U118 (N_118,In_382,In_55);
and U119 (N_119,In_458,In_264);
and U120 (N_120,In_444,In_168);
nand U121 (N_121,N_58,In_414);
nor U122 (N_122,N_43,In_445);
nor U123 (N_123,In_303,In_197);
or U124 (N_124,In_316,In_157);
or U125 (N_125,N_71,In_345);
xor U126 (N_126,In_309,N_17);
or U127 (N_127,In_290,In_66);
and U128 (N_128,In_61,In_371);
or U129 (N_129,In_337,In_148);
or U130 (N_130,In_8,In_202);
or U131 (N_131,In_20,In_295);
nand U132 (N_132,In_373,In_254);
nand U133 (N_133,In_488,In_9);
nand U134 (N_134,In_65,In_284);
or U135 (N_135,In_461,In_381);
nor U136 (N_136,In_308,In_104);
and U137 (N_137,In_470,In_206);
nor U138 (N_138,N_5,In_73);
nor U139 (N_139,In_286,In_384);
and U140 (N_140,In_190,In_411);
nand U141 (N_141,In_250,In_310);
nor U142 (N_142,In_274,In_26);
or U143 (N_143,In_423,In_467);
or U144 (N_144,N_51,In_67);
nor U145 (N_145,In_150,In_380);
or U146 (N_146,In_100,N_64);
and U147 (N_147,In_448,In_343);
and U148 (N_148,N_18,In_158);
and U149 (N_149,N_10,In_321);
nand U150 (N_150,In_270,In_6);
or U151 (N_151,In_258,In_156);
and U152 (N_152,In_243,In_149);
nor U153 (N_153,In_385,In_130);
and U154 (N_154,In_271,In_83);
and U155 (N_155,In_291,In_334);
and U156 (N_156,In_394,N_16);
and U157 (N_157,In_173,In_277);
and U158 (N_158,In_155,N_93);
and U159 (N_159,N_62,N_39);
or U160 (N_160,N_80,In_403);
nand U161 (N_161,N_128,In_22);
and U162 (N_162,In_234,N_33);
or U163 (N_163,In_217,In_125);
nor U164 (N_164,In_212,In_478);
nor U165 (N_165,In_341,In_346);
or U166 (N_166,N_41,N_124);
or U167 (N_167,N_114,In_90);
or U168 (N_168,In_477,N_23);
nor U169 (N_169,In_240,N_106);
nand U170 (N_170,In_194,In_400);
or U171 (N_171,N_133,In_455);
nor U172 (N_172,In_328,In_459);
or U173 (N_173,In_433,In_151);
or U174 (N_174,N_118,In_262);
or U175 (N_175,N_12,N_27);
or U176 (N_176,In_221,N_98);
or U177 (N_177,N_15,In_395);
and U178 (N_178,N_14,N_138);
or U179 (N_179,In_350,N_121);
or U180 (N_180,In_46,In_87);
nand U181 (N_181,N_116,In_191);
nand U182 (N_182,In_327,N_63);
or U183 (N_183,N_84,In_358);
and U184 (N_184,In_294,N_4);
nand U185 (N_185,In_223,In_288);
nor U186 (N_186,In_98,N_88);
and U187 (N_187,N_112,N_142);
nand U188 (N_188,In_163,In_452);
xor U189 (N_189,In_389,In_412);
nor U190 (N_190,N_109,N_86);
and U191 (N_191,In_132,In_344);
nor U192 (N_192,N_139,In_434);
nor U193 (N_193,In_474,In_214);
or U194 (N_194,In_210,N_57);
nand U195 (N_195,N_125,In_419);
nor U196 (N_196,In_484,N_37);
and U197 (N_197,In_301,In_142);
nor U198 (N_198,In_435,N_26);
nand U199 (N_199,N_99,In_281);
nand U200 (N_200,In_302,In_402);
nand U201 (N_201,In_416,N_108);
or U202 (N_202,In_379,N_40);
and U203 (N_203,In_145,In_407);
and U204 (N_204,N_46,N_76);
nand U205 (N_205,In_246,In_80);
or U206 (N_206,In_47,N_48);
nand U207 (N_207,In_377,N_75);
nor U208 (N_208,In_170,In_468);
nand U209 (N_209,In_300,N_42);
nand U210 (N_210,N_7,In_11);
xor U211 (N_211,In_167,N_144);
and U212 (N_212,In_68,In_18);
and U213 (N_213,N_31,N_100);
or U214 (N_214,N_145,In_136);
and U215 (N_215,In_207,N_36);
nand U216 (N_216,In_76,In_432);
or U217 (N_217,In_172,In_122);
nand U218 (N_218,N_122,In_259);
nor U219 (N_219,In_117,In_219);
nand U220 (N_220,N_91,N_120);
and U221 (N_221,N_96,In_487);
and U222 (N_222,N_66,In_129);
or U223 (N_223,N_97,In_140);
nand U224 (N_224,N_78,In_441);
and U225 (N_225,N_8,In_139);
and U226 (N_226,N_187,In_493);
or U227 (N_227,N_126,N_167);
and U228 (N_228,N_214,In_95);
nand U229 (N_229,In_53,N_65);
and U230 (N_230,In_293,In_265);
nand U231 (N_231,In_114,In_215);
nand U232 (N_232,N_82,In_30);
or U233 (N_233,N_159,In_426);
and U234 (N_234,In_200,N_208);
or U235 (N_235,N_94,N_103);
or U236 (N_236,In_102,In_457);
and U237 (N_237,N_115,N_11);
or U238 (N_238,N_28,N_186);
and U239 (N_239,In_391,In_182);
or U240 (N_240,In_174,N_175);
nand U241 (N_241,N_90,In_331);
nor U242 (N_242,N_207,In_496);
or U243 (N_243,N_183,N_156);
nand U244 (N_244,N_164,N_60);
nor U245 (N_245,In_460,In_63);
nand U246 (N_246,In_282,In_230);
or U247 (N_247,In_17,N_3);
or U248 (N_248,N_182,N_193);
or U249 (N_249,N_221,N_153);
or U250 (N_250,In_204,N_181);
nand U251 (N_251,N_147,In_420);
and U252 (N_252,N_178,In_24);
nand U253 (N_253,In_203,N_166);
and U254 (N_254,In_119,In_62);
nand U255 (N_255,In_120,In_123);
nand U256 (N_256,N_176,In_1);
or U257 (N_257,N_201,N_203);
nor U258 (N_258,In_255,N_141);
nand U259 (N_259,In_398,N_204);
nand U260 (N_260,In_491,In_454);
nor U261 (N_261,N_102,In_319);
or U262 (N_262,In_99,In_266);
nor U263 (N_263,N_171,In_5);
nand U264 (N_264,N_161,In_401);
nor U265 (N_265,In_27,In_188);
and U266 (N_266,In_147,In_185);
or U267 (N_267,N_224,N_157);
nand U268 (N_268,N_218,N_45);
nand U269 (N_269,N_104,N_217);
nand U270 (N_270,N_2,N_30);
and U271 (N_271,N_132,In_245);
nand U272 (N_272,N_81,N_20);
nor U273 (N_273,In_44,N_163);
nand U274 (N_274,In_494,N_151);
nand U275 (N_275,N_210,N_89);
and U276 (N_276,In_466,N_61);
nor U277 (N_277,In_297,N_196);
or U278 (N_278,N_216,In_193);
nor U279 (N_279,In_205,N_195);
or U280 (N_280,In_278,N_107);
nor U281 (N_281,N_173,N_56);
nand U282 (N_282,N_129,N_143);
and U283 (N_283,N_212,In_239);
nand U284 (N_284,N_220,N_185);
nor U285 (N_285,In_424,N_170);
or U286 (N_286,In_134,In_251);
nor U287 (N_287,N_179,N_209);
and U288 (N_288,N_149,N_0);
nor U289 (N_289,N_69,N_59);
nand U290 (N_290,N_95,In_498);
nor U291 (N_291,N_205,In_492);
nand U292 (N_292,N_101,N_168);
and U293 (N_293,N_154,In_272);
nor U294 (N_294,In_336,In_421);
or U295 (N_295,N_130,N_223);
and U296 (N_296,N_111,N_135);
or U297 (N_297,N_68,N_35);
nor U298 (N_298,N_219,In_19);
or U299 (N_299,In_224,In_184);
nand U300 (N_300,N_54,N_148);
and U301 (N_301,N_233,In_242);
and U302 (N_302,N_184,N_117);
nand U303 (N_303,N_273,N_241);
nor U304 (N_304,In_135,N_55);
nand U305 (N_305,In_195,In_78);
and U306 (N_306,N_249,In_16);
nor U307 (N_307,N_294,N_230);
nand U308 (N_308,N_279,N_191);
nor U309 (N_309,N_215,N_238);
and U310 (N_310,N_264,N_270);
or U311 (N_311,N_269,N_262);
and U312 (N_312,N_188,N_162);
and U313 (N_313,N_50,In_273);
or U314 (N_314,In_107,In_2);
or U315 (N_315,N_293,N_21);
nand U316 (N_316,N_197,N_140);
nand U317 (N_317,In_91,N_276);
xor U318 (N_318,In_450,N_291);
nand U319 (N_319,N_275,N_260);
nor U320 (N_320,In_25,N_192);
or U321 (N_321,N_268,N_131);
or U322 (N_322,N_251,In_176);
or U323 (N_323,N_13,N_255);
nor U324 (N_324,N_229,N_105);
nor U325 (N_325,N_288,N_283);
or U326 (N_326,In_32,N_256);
and U327 (N_327,In_166,N_190);
nor U328 (N_328,N_243,N_160);
or U329 (N_329,In_326,N_165);
and U330 (N_330,N_246,N_299);
nand U331 (N_331,In_69,In_463);
and U332 (N_332,N_24,N_257);
nand U333 (N_333,N_284,N_286);
and U334 (N_334,In_75,N_236);
and U335 (N_335,N_281,N_146);
nand U336 (N_336,N_213,N_202);
nand U337 (N_337,N_79,In_71);
or U338 (N_338,N_150,N_199);
nand U339 (N_339,N_247,N_239);
nand U340 (N_340,N_169,In_257);
and U341 (N_341,N_22,N_174);
and U342 (N_342,N_253,N_211);
and U343 (N_343,In_169,N_240);
nor U344 (N_344,N_1,In_352);
nand U345 (N_345,N_194,N_172);
and U346 (N_346,N_136,N_155);
or U347 (N_347,N_134,N_232);
nor U348 (N_348,N_296,N_177);
xor U349 (N_349,N_67,N_77);
nor U350 (N_350,N_85,N_261);
nor U351 (N_351,In_70,N_250);
nor U352 (N_352,N_231,N_92);
and U353 (N_353,In_52,N_244);
or U354 (N_354,N_292,In_404);
nor U355 (N_355,N_248,N_72);
nor U356 (N_356,N_267,In_59);
nor U357 (N_357,In_285,N_87);
and U358 (N_358,In_320,In_376);
nor U359 (N_359,In_138,In_79);
nand U360 (N_360,N_245,N_290);
nand U361 (N_361,In_299,In_324);
or U362 (N_362,In_268,N_227);
or U363 (N_363,N_274,N_222);
nor U364 (N_364,In_41,N_271);
or U365 (N_365,In_473,N_47);
nor U366 (N_366,In_77,N_44);
nor U367 (N_367,In_233,In_14);
xor U368 (N_368,N_83,In_33);
and U369 (N_369,N_228,N_234);
nand U370 (N_370,N_113,N_158);
and U371 (N_371,In_45,In_366);
nand U372 (N_372,N_280,N_254);
or U373 (N_373,N_137,In_449);
nor U374 (N_374,N_127,In_222);
nand U375 (N_375,N_242,N_309);
or U376 (N_376,N_360,N_333);
nor U377 (N_377,N_344,N_364);
and U378 (N_378,N_352,N_225);
and U379 (N_379,In_220,N_287);
or U380 (N_380,N_374,N_336);
nand U381 (N_381,In_50,N_354);
nor U382 (N_382,N_305,In_443);
or U383 (N_383,In_37,N_258);
and U384 (N_384,N_278,N_335);
nand U385 (N_385,N_343,N_313);
and U386 (N_386,N_304,N_373);
nor U387 (N_387,N_189,N_285);
nor U388 (N_388,N_372,N_319);
or U389 (N_389,N_314,N_351);
nor U390 (N_390,N_263,N_308);
nand U391 (N_391,N_323,N_358);
nand U392 (N_392,N_295,N_363);
and U393 (N_393,N_330,N_332);
and U394 (N_394,N_347,N_369);
or U395 (N_395,In_175,In_209);
and U396 (N_396,N_350,N_356);
nand U397 (N_397,N_198,N_318);
nor U398 (N_398,N_180,N_70);
xor U399 (N_399,N_265,N_353);
and U400 (N_400,N_357,N_306);
nor U401 (N_401,N_361,N_362);
nand U402 (N_402,N_317,N_320);
and U403 (N_403,N_110,In_96);
and U404 (N_404,N_152,N_342);
nor U405 (N_405,N_345,N_259);
nand U406 (N_406,N_301,N_327);
nor U407 (N_407,In_263,N_302);
xnor U408 (N_408,N_300,N_316);
nor U409 (N_409,N_348,N_298);
or U410 (N_410,In_363,N_365);
nand U411 (N_411,N_307,N_334);
or U412 (N_412,N_123,In_236);
nor U413 (N_413,N_367,N_310);
nand U414 (N_414,N_119,N_338);
or U415 (N_415,In_357,N_311);
xnor U416 (N_416,N_252,In_4);
nor U417 (N_417,N_355,N_371);
nor U418 (N_418,In_21,N_282);
nor U419 (N_419,N_340,N_266);
nor U420 (N_420,N_370,N_272);
nand U421 (N_421,N_226,N_200);
nor U422 (N_422,N_206,In_399);
nor U423 (N_423,N_328,In_311);
nand U424 (N_424,N_237,N_329);
nand U425 (N_425,N_359,N_235);
and U426 (N_426,N_315,N_349);
or U427 (N_427,N_325,In_56);
xor U428 (N_428,N_289,N_322);
and U429 (N_429,N_366,In_12);
nor U430 (N_430,N_341,N_368);
nand U431 (N_431,In_261,N_324);
and U432 (N_432,N_339,N_303);
or U433 (N_433,N_312,N_297);
nor U434 (N_434,In_330,N_277);
or U435 (N_435,N_337,N_346);
xnor U436 (N_436,N_326,N_321);
nand U437 (N_437,N_331,N_312);
xnor U438 (N_438,N_356,N_335);
nor U439 (N_439,N_358,N_110);
or U440 (N_440,N_308,N_206);
nand U441 (N_441,N_282,N_119);
or U442 (N_442,N_198,N_341);
and U443 (N_443,N_307,N_123);
nand U444 (N_444,In_4,N_345);
nand U445 (N_445,N_366,N_189);
and U446 (N_446,N_356,N_206);
nand U447 (N_447,N_345,In_263);
and U448 (N_448,In_263,N_372);
nand U449 (N_449,N_226,N_277);
or U450 (N_450,N_376,N_425);
and U451 (N_451,N_405,N_406);
nand U452 (N_452,N_396,N_410);
or U453 (N_453,N_384,N_398);
xnor U454 (N_454,N_408,N_421);
nand U455 (N_455,N_423,N_412);
or U456 (N_456,N_422,N_401);
or U457 (N_457,N_435,N_385);
and U458 (N_458,N_429,N_414);
nor U459 (N_459,N_403,N_440);
nand U460 (N_460,N_443,N_386);
and U461 (N_461,N_399,N_393);
or U462 (N_462,N_428,N_409);
nor U463 (N_463,N_378,N_442);
or U464 (N_464,N_415,N_430);
nor U465 (N_465,N_431,N_404);
nand U466 (N_466,N_394,N_413);
and U467 (N_467,N_436,N_432);
nand U468 (N_468,N_424,N_395);
nand U469 (N_469,N_427,N_397);
and U470 (N_470,N_446,N_420);
and U471 (N_471,N_448,N_419);
or U472 (N_472,N_407,N_426);
nor U473 (N_473,N_402,N_445);
nor U474 (N_474,N_434,N_447);
nor U475 (N_475,N_379,N_444);
and U476 (N_476,N_417,N_416);
and U477 (N_477,N_390,N_441);
nand U478 (N_478,N_449,N_377);
nor U479 (N_479,N_391,N_411);
or U480 (N_480,N_438,N_383);
or U481 (N_481,N_418,N_400);
nand U482 (N_482,N_375,N_387);
or U483 (N_483,N_433,N_392);
nand U484 (N_484,N_437,N_389);
and U485 (N_485,N_381,N_439);
nor U486 (N_486,N_382,N_380);
and U487 (N_487,N_388,N_434);
or U488 (N_488,N_384,N_422);
nand U489 (N_489,N_395,N_449);
and U490 (N_490,N_422,N_407);
nand U491 (N_491,N_382,N_408);
and U492 (N_492,N_382,N_444);
and U493 (N_493,N_449,N_414);
nand U494 (N_494,N_441,N_443);
nand U495 (N_495,N_435,N_445);
nand U496 (N_496,N_415,N_388);
or U497 (N_497,N_391,N_419);
and U498 (N_498,N_440,N_433);
nor U499 (N_499,N_448,N_410);
and U500 (N_500,N_410,N_424);
nor U501 (N_501,N_384,N_412);
nor U502 (N_502,N_378,N_400);
nand U503 (N_503,N_437,N_410);
nand U504 (N_504,N_416,N_408);
nand U505 (N_505,N_416,N_414);
or U506 (N_506,N_401,N_428);
and U507 (N_507,N_377,N_383);
nor U508 (N_508,N_390,N_409);
and U509 (N_509,N_430,N_392);
nor U510 (N_510,N_385,N_397);
nand U511 (N_511,N_404,N_399);
nand U512 (N_512,N_377,N_425);
nand U513 (N_513,N_449,N_425);
nand U514 (N_514,N_392,N_422);
xor U515 (N_515,N_392,N_424);
or U516 (N_516,N_388,N_380);
nand U517 (N_517,N_415,N_418);
or U518 (N_518,N_442,N_390);
nor U519 (N_519,N_432,N_445);
or U520 (N_520,N_391,N_406);
nand U521 (N_521,N_428,N_432);
nor U522 (N_522,N_403,N_377);
or U523 (N_523,N_402,N_420);
nor U524 (N_524,N_447,N_427);
nand U525 (N_525,N_502,N_463);
or U526 (N_526,N_496,N_451);
and U527 (N_527,N_452,N_503);
nor U528 (N_528,N_516,N_478);
nand U529 (N_529,N_518,N_506);
nor U530 (N_530,N_487,N_515);
nor U531 (N_531,N_499,N_484);
and U532 (N_532,N_480,N_471);
nor U533 (N_533,N_454,N_458);
nor U534 (N_534,N_461,N_489);
or U535 (N_535,N_524,N_488);
nand U536 (N_536,N_467,N_457);
nor U537 (N_537,N_491,N_472);
nor U538 (N_538,N_509,N_462);
nor U539 (N_539,N_495,N_504);
and U540 (N_540,N_469,N_473);
or U541 (N_541,N_474,N_453);
or U542 (N_542,N_492,N_497);
xnor U543 (N_543,N_520,N_459);
nor U544 (N_544,N_501,N_513);
xor U545 (N_545,N_460,N_523);
and U546 (N_546,N_481,N_508);
nand U547 (N_547,N_522,N_486);
and U548 (N_548,N_521,N_507);
and U549 (N_549,N_465,N_511);
nand U550 (N_550,N_470,N_483);
nor U551 (N_551,N_468,N_476);
nand U552 (N_552,N_450,N_510);
xor U553 (N_553,N_475,N_494);
or U554 (N_554,N_482,N_493);
or U555 (N_555,N_479,N_505);
or U556 (N_556,N_485,N_466);
nor U557 (N_557,N_514,N_519);
and U558 (N_558,N_490,N_464);
or U559 (N_559,N_455,N_512);
or U560 (N_560,N_517,N_498);
nand U561 (N_561,N_477,N_456);
nand U562 (N_562,N_500,N_476);
or U563 (N_563,N_460,N_507);
and U564 (N_564,N_452,N_517);
or U565 (N_565,N_513,N_482);
nor U566 (N_566,N_475,N_480);
and U567 (N_567,N_472,N_504);
xor U568 (N_568,N_520,N_513);
nand U569 (N_569,N_451,N_511);
or U570 (N_570,N_504,N_503);
and U571 (N_571,N_494,N_487);
nor U572 (N_572,N_476,N_479);
or U573 (N_573,N_459,N_456);
nor U574 (N_574,N_479,N_501);
or U575 (N_575,N_516,N_461);
xnor U576 (N_576,N_499,N_464);
nor U577 (N_577,N_517,N_500);
or U578 (N_578,N_476,N_484);
or U579 (N_579,N_493,N_499);
nand U580 (N_580,N_499,N_486);
nand U581 (N_581,N_456,N_508);
nor U582 (N_582,N_474,N_519);
nor U583 (N_583,N_465,N_472);
or U584 (N_584,N_493,N_474);
and U585 (N_585,N_469,N_493);
nor U586 (N_586,N_486,N_507);
nor U587 (N_587,N_480,N_498);
nor U588 (N_588,N_458,N_515);
nor U589 (N_589,N_497,N_489);
and U590 (N_590,N_471,N_465);
nor U591 (N_591,N_516,N_497);
nand U592 (N_592,N_506,N_471);
or U593 (N_593,N_482,N_496);
nor U594 (N_594,N_518,N_484);
nand U595 (N_595,N_479,N_512);
nor U596 (N_596,N_498,N_500);
nor U597 (N_597,N_470,N_456);
or U598 (N_598,N_497,N_463);
nor U599 (N_599,N_497,N_519);
nand U600 (N_600,N_530,N_585);
nor U601 (N_601,N_541,N_552);
nand U602 (N_602,N_588,N_532);
nor U603 (N_603,N_525,N_538);
and U604 (N_604,N_578,N_558);
or U605 (N_605,N_597,N_598);
nor U606 (N_606,N_539,N_528);
or U607 (N_607,N_576,N_531);
or U608 (N_608,N_584,N_544);
and U609 (N_609,N_575,N_569);
nor U610 (N_610,N_591,N_589);
nand U611 (N_611,N_563,N_537);
nor U612 (N_612,N_572,N_529);
and U613 (N_613,N_573,N_540);
nor U614 (N_614,N_545,N_560);
or U615 (N_615,N_579,N_566);
nor U616 (N_616,N_526,N_581);
or U617 (N_617,N_595,N_587);
nand U618 (N_618,N_580,N_556);
nor U619 (N_619,N_548,N_547);
nand U620 (N_620,N_568,N_593);
and U621 (N_621,N_550,N_543);
nor U622 (N_622,N_596,N_534);
and U623 (N_623,N_527,N_557);
nor U624 (N_624,N_554,N_535);
and U625 (N_625,N_577,N_567);
or U626 (N_626,N_546,N_559);
or U627 (N_627,N_594,N_549);
nor U628 (N_628,N_561,N_582);
nand U629 (N_629,N_590,N_565);
nor U630 (N_630,N_592,N_571);
or U631 (N_631,N_599,N_553);
and U632 (N_632,N_536,N_562);
nor U633 (N_633,N_574,N_564);
nand U634 (N_634,N_542,N_555);
nor U635 (N_635,N_551,N_533);
nand U636 (N_636,N_586,N_583);
or U637 (N_637,N_570,N_532);
and U638 (N_638,N_553,N_589);
and U639 (N_639,N_572,N_587);
and U640 (N_640,N_545,N_539);
and U641 (N_641,N_560,N_543);
and U642 (N_642,N_582,N_589);
and U643 (N_643,N_588,N_541);
nand U644 (N_644,N_554,N_594);
nor U645 (N_645,N_550,N_597);
nor U646 (N_646,N_572,N_585);
nand U647 (N_647,N_538,N_580);
and U648 (N_648,N_565,N_574);
and U649 (N_649,N_598,N_579);
or U650 (N_650,N_527,N_574);
and U651 (N_651,N_590,N_550);
or U652 (N_652,N_596,N_597);
or U653 (N_653,N_586,N_581);
or U654 (N_654,N_572,N_553);
or U655 (N_655,N_574,N_546);
nor U656 (N_656,N_565,N_534);
or U657 (N_657,N_530,N_592);
nor U658 (N_658,N_563,N_577);
nor U659 (N_659,N_526,N_541);
and U660 (N_660,N_566,N_560);
nand U661 (N_661,N_578,N_525);
and U662 (N_662,N_572,N_528);
and U663 (N_663,N_587,N_532);
or U664 (N_664,N_536,N_594);
or U665 (N_665,N_545,N_586);
and U666 (N_666,N_559,N_532);
and U667 (N_667,N_579,N_574);
nand U668 (N_668,N_598,N_544);
nand U669 (N_669,N_582,N_586);
or U670 (N_670,N_562,N_560);
nor U671 (N_671,N_548,N_549);
nor U672 (N_672,N_558,N_577);
and U673 (N_673,N_596,N_571);
nor U674 (N_674,N_596,N_567);
and U675 (N_675,N_643,N_668);
nor U676 (N_676,N_613,N_609);
nor U677 (N_677,N_642,N_617);
nand U678 (N_678,N_611,N_600);
or U679 (N_679,N_627,N_651);
and U680 (N_680,N_614,N_623);
nor U681 (N_681,N_659,N_621);
nand U682 (N_682,N_622,N_650);
and U683 (N_683,N_641,N_601);
nand U684 (N_684,N_639,N_633);
and U685 (N_685,N_672,N_628);
nand U686 (N_686,N_615,N_667);
nand U687 (N_687,N_666,N_671);
nand U688 (N_688,N_602,N_664);
or U689 (N_689,N_655,N_608);
nor U690 (N_690,N_632,N_616);
nand U691 (N_691,N_656,N_644);
nor U692 (N_692,N_661,N_604);
and U693 (N_693,N_610,N_624);
or U694 (N_694,N_670,N_640);
nand U695 (N_695,N_618,N_612);
nor U696 (N_696,N_648,N_605);
and U697 (N_697,N_673,N_665);
nand U698 (N_698,N_654,N_663);
or U699 (N_699,N_606,N_638);
nor U700 (N_700,N_674,N_607);
or U701 (N_701,N_662,N_669);
and U702 (N_702,N_645,N_635);
and U703 (N_703,N_660,N_634);
or U704 (N_704,N_649,N_603);
or U705 (N_705,N_658,N_626);
and U706 (N_706,N_629,N_620);
or U707 (N_707,N_625,N_646);
and U708 (N_708,N_619,N_652);
or U709 (N_709,N_647,N_653);
nor U710 (N_710,N_637,N_630);
or U711 (N_711,N_657,N_631);
nand U712 (N_712,N_636,N_617);
and U713 (N_713,N_634,N_659);
and U714 (N_714,N_643,N_618);
or U715 (N_715,N_614,N_661);
and U716 (N_716,N_622,N_654);
or U717 (N_717,N_605,N_636);
nand U718 (N_718,N_670,N_661);
or U719 (N_719,N_611,N_647);
and U720 (N_720,N_655,N_663);
and U721 (N_721,N_607,N_656);
nor U722 (N_722,N_668,N_670);
or U723 (N_723,N_653,N_627);
nand U724 (N_724,N_667,N_672);
and U725 (N_725,N_605,N_607);
nor U726 (N_726,N_617,N_601);
and U727 (N_727,N_632,N_620);
or U728 (N_728,N_603,N_656);
or U729 (N_729,N_622,N_602);
nand U730 (N_730,N_650,N_659);
nor U731 (N_731,N_660,N_652);
or U732 (N_732,N_602,N_650);
nand U733 (N_733,N_629,N_667);
nor U734 (N_734,N_625,N_647);
nand U735 (N_735,N_609,N_658);
xor U736 (N_736,N_607,N_640);
nand U737 (N_737,N_659,N_626);
nand U738 (N_738,N_608,N_650);
nand U739 (N_739,N_665,N_600);
xor U740 (N_740,N_635,N_646);
nor U741 (N_741,N_621,N_672);
and U742 (N_742,N_618,N_674);
or U743 (N_743,N_600,N_649);
and U744 (N_744,N_613,N_667);
or U745 (N_745,N_630,N_623);
nand U746 (N_746,N_645,N_628);
nor U747 (N_747,N_637,N_666);
and U748 (N_748,N_643,N_621);
and U749 (N_749,N_672,N_637);
nand U750 (N_750,N_705,N_694);
and U751 (N_751,N_723,N_678);
and U752 (N_752,N_719,N_685);
and U753 (N_753,N_686,N_729);
and U754 (N_754,N_680,N_725);
or U755 (N_755,N_720,N_735);
or U756 (N_756,N_692,N_681);
nor U757 (N_757,N_711,N_701);
or U758 (N_758,N_675,N_727);
nor U759 (N_759,N_682,N_733);
nor U760 (N_760,N_713,N_715);
nand U761 (N_761,N_708,N_745);
and U762 (N_762,N_740,N_737);
and U763 (N_763,N_742,N_722);
and U764 (N_764,N_743,N_747);
nand U765 (N_765,N_704,N_736);
nor U766 (N_766,N_697,N_699);
nor U767 (N_767,N_691,N_709);
nand U768 (N_768,N_702,N_676);
nand U769 (N_769,N_732,N_748);
and U770 (N_770,N_698,N_687);
and U771 (N_771,N_683,N_739);
nand U772 (N_772,N_677,N_693);
and U773 (N_773,N_749,N_706);
or U774 (N_774,N_741,N_731);
nor U775 (N_775,N_724,N_710);
nor U776 (N_776,N_700,N_746);
nor U777 (N_777,N_734,N_712);
and U778 (N_778,N_721,N_717);
and U779 (N_779,N_728,N_716);
and U780 (N_780,N_684,N_696);
and U781 (N_781,N_714,N_738);
and U782 (N_782,N_690,N_688);
or U783 (N_783,N_679,N_718);
or U784 (N_784,N_744,N_703);
or U785 (N_785,N_707,N_726);
or U786 (N_786,N_730,N_695);
or U787 (N_787,N_689,N_698);
nor U788 (N_788,N_683,N_685);
nand U789 (N_789,N_736,N_709);
nor U790 (N_790,N_708,N_715);
nand U791 (N_791,N_687,N_700);
nand U792 (N_792,N_688,N_714);
or U793 (N_793,N_734,N_694);
or U794 (N_794,N_736,N_711);
or U795 (N_795,N_687,N_688);
and U796 (N_796,N_686,N_705);
nand U797 (N_797,N_719,N_713);
nand U798 (N_798,N_710,N_747);
or U799 (N_799,N_693,N_675);
nor U800 (N_800,N_723,N_715);
nor U801 (N_801,N_722,N_684);
nor U802 (N_802,N_726,N_727);
or U803 (N_803,N_748,N_728);
nor U804 (N_804,N_701,N_733);
nand U805 (N_805,N_690,N_722);
and U806 (N_806,N_748,N_744);
and U807 (N_807,N_733,N_700);
and U808 (N_808,N_692,N_685);
nand U809 (N_809,N_732,N_676);
nand U810 (N_810,N_691,N_739);
or U811 (N_811,N_736,N_715);
nand U812 (N_812,N_726,N_685);
nor U813 (N_813,N_704,N_724);
or U814 (N_814,N_690,N_721);
nor U815 (N_815,N_680,N_689);
and U816 (N_816,N_694,N_707);
or U817 (N_817,N_705,N_692);
and U818 (N_818,N_702,N_678);
nand U819 (N_819,N_694,N_740);
and U820 (N_820,N_714,N_692);
and U821 (N_821,N_732,N_706);
and U822 (N_822,N_683,N_678);
and U823 (N_823,N_739,N_682);
nand U824 (N_824,N_728,N_722);
nor U825 (N_825,N_769,N_805);
and U826 (N_826,N_759,N_808);
or U827 (N_827,N_796,N_792);
or U828 (N_828,N_765,N_754);
and U829 (N_829,N_806,N_816);
nand U830 (N_830,N_811,N_800);
or U831 (N_831,N_820,N_763);
nor U832 (N_832,N_752,N_823);
and U833 (N_833,N_812,N_795);
nand U834 (N_834,N_815,N_780);
or U835 (N_835,N_767,N_790);
and U836 (N_836,N_777,N_804);
nor U837 (N_837,N_751,N_785);
nand U838 (N_838,N_778,N_755);
or U839 (N_839,N_818,N_794);
nor U840 (N_840,N_781,N_791);
and U841 (N_841,N_757,N_766);
and U842 (N_842,N_779,N_758);
xor U843 (N_843,N_775,N_753);
nor U844 (N_844,N_750,N_810);
and U845 (N_845,N_776,N_797);
nand U846 (N_846,N_773,N_807);
and U847 (N_847,N_798,N_771);
nor U848 (N_848,N_799,N_762);
and U849 (N_849,N_782,N_809);
or U850 (N_850,N_783,N_813);
nand U851 (N_851,N_760,N_819);
nand U852 (N_852,N_802,N_761);
and U853 (N_853,N_770,N_772);
nand U854 (N_854,N_824,N_793);
nand U855 (N_855,N_821,N_803);
nand U856 (N_856,N_789,N_801);
nor U857 (N_857,N_784,N_822);
nand U858 (N_858,N_768,N_764);
or U859 (N_859,N_814,N_756);
and U860 (N_860,N_787,N_817);
nand U861 (N_861,N_786,N_788);
nand U862 (N_862,N_774,N_784);
nand U863 (N_863,N_811,N_813);
nor U864 (N_864,N_782,N_789);
nor U865 (N_865,N_763,N_778);
and U866 (N_866,N_766,N_752);
nand U867 (N_867,N_808,N_796);
nand U868 (N_868,N_781,N_812);
nor U869 (N_869,N_799,N_816);
or U870 (N_870,N_813,N_796);
nor U871 (N_871,N_815,N_806);
or U872 (N_872,N_789,N_786);
and U873 (N_873,N_822,N_763);
and U874 (N_874,N_818,N_819);
nand U875 (N_875,N_816,N_775);
nand U876 (N_876,N_793,N_809);
xnor U877 (N_877,N_757,N_758);
and U878 (N_878,N_750,N_789);
nor U879 (N_879,N_780,N_820);
nor U880 (N_880,N_803,N_772);
or U881 (N_881,N_795,N_780);
or U882 (N_882,N_785,N_755);
and U883 (N_883,N_812,N_805);
xnor U884 (N_884,N_812,N_820);
nor U885 (N_885,N_766,N_795);
and U886 (N_886,N_808,N_790);
nand U887 (N_887,N_772,N_819);
and U888 (N_888,N_802,N_759);
and U889 (N_889,N_788,N_791);
nand U890 (N_890,N_814,N_764);
nor U891 (N_891,N_805,N_821);
nor U892 (N_892,N_800,N_767);
or U893 (N_893,N_779,N_768);
or U894 (N_894,N_774,N_812);
and U895 (N_895,N_760,N_803);
nand U896 (N_896,N_807,N_796);
nor U897 (N_897,N_770,N_776);
nor U898 (N_898,N_756,N_801);
nand U899 (N_899,N_767,N_787);
or U900 (N_900,N_879,N_882);
or U901 (N_901,N_831,N_870);
nand U902 (N_902,N_884,N_865);
and U903 (N_903,N_896,N_866);
or U904 (N_904,N_826,N_859);
or U905 (N_905,N_864,N_868);
nand U906 (N_906,N_841,N_880);
nor U907 (N_907,N_860,N_847);
and U908 (N_908,N_839,N_849);
or U909 (N_909,N_881,N_834);
nor U910 (N_910,N_852,N_837);
nor U911 (N_911,N_892,N_878);
and U912 (N_912,N_846,N_833);
nor U913 (N_913,N_827,N_891);
nor U914 (N_914,N_851,N_874);
or U915 (N_915,N_856,N_899);
or U916 (N_916,N_883,N_840);
and U917 (N_917,N_832,N_886);
nand U918 (N_918,N_875,N_889);
nand U919 (N_919,N_871,N_830);
or U920 (N_920,N_854,N_863);
xor U921 (N_921,N_848,N_897);
and U922 (N_922,N_887,N_843);
and U923 (N_923,N_850,N_844);
nand U924 (N_924,N_872,N_853);
nor U925 (N_925,N_855,N_862);
nor U926 (N_926,N_845,N_893);
and U927 (N_927,N_888,N_838);
nor U928 (N_928,N_858,N_885);
or U929 (N_929,N_873,N_829);
nor U930 (N_930,N_869,N_894);
nor U931 (N_931,N_895,N_828);
nand U932 (N_932,N_867,N_857);
nor U933 (N_933,N_836,N_835);
nand U934 (N_934,N_890,N_842);
or U935 (N_935,N_825,N_898);
nand U936 (N_936,N_876,N_877);
nand U937 (N_937,N_861,N_853);
and U938 (N_938,N_897,N_832);
nor U939 (N_939,N_883,N_898);
or U940 (N_940,N_892,N_840);
nand U941 (N_941,N_825,N_857);
nor U942 (N_942,N_896,N_892);
nor U943 (N_943,N_896,N_894);
nand U944 (N_944,N_827,N_867);
nor U945 (N_945,N_863,N_839);
and U946 (N_946,N_866,N_849);
and U947 (N_947,N_847,N_878);
nand U948 (N_948,N_865,N_839);
and U949 (N_949,N_850,N_870);
nor U950 (N_950,N_897,N_882);
nor U951 (N_951,N_874,N_844);
nand U952 (N_952,N_829,N_897);
and U953 (N_953,N_883,N_884);
nor U954 (N_954,N_854,N_875);
nand U955 (N_955,N_854,N_830);
nand U956 (N_956,N_899,N_834);
or U957 (N_957,N_898,N_892);
or U958 (N_958,N_896,N_862);
or U959 (N_959,N_873,N_882);
nand U960 (N_960,N_876,N_873);
nor U961 (N_961,N_854,N_838);
nor U962 (N_962,N_879,N_863);
nor U963 (N_963,N_839,N_836);
nor U964 (N_964,N_872,N_835);
or U965 (N_965,N_877,N_852);
and U966 (N_966,N_872,N_837);
nor U967 (N_967,N_862,N_889);
nor U968 (N_968,N_854,N_848);
nor U969 (N_969,N_897,N_887);
and U970 (N_970,N_852,N_880);
or U971 (N_971,N_843,N_873);
nor U972 (N_972,N_829,N_894);
nor U973 (N_973,N_868,N_887);
nor U974 (N_974,N_833,N_849);
and U975 (N_975,N_909,N_931);
nand U976 (N_976,N_905,N_948);
nand U977 (N_977,N_923,N_971);
nor U978 (N_978,N_911,N_921);
nand U979 (N_979,N_957,N_962);
and U980 (N_980,N_970,N_901);
nor U981 (N_981,N_965,N_914);
or U982 (N_982,N_944,N_950);
nand U983 (N_983,N_928,N_919);
nand U984 (N_984,N_937,N_973);
or U985 (N_985,N_955,N_906);
or U986 (N_986,N_924,N_912);
and U987 (N_987,N_930,N_967);
or U988 (N_988,N_945,N_902);
nand U989 (N_989,N_900,N_907);
nor U990 (N_990,N_903,N_941);
and U991 (N_991,N_954,N_947);
and U992 (N_992,N_963,N_964);
or U993 (N_993,N_939,N_913);
nand U994 (N_994,N_974,N_949);
nand U995 (N_995,N_940,N_936);
and U996 (N_996,N_908,N_942);
or U997 (N_997,N_916,N_934);
and U998 (N_998,N_969,N_952);
and U999 (N_999,N_904,N_961);
nor U1000 (N_1000,N_953,N_956);
nand U1001 (N_1001,N_966,N_932);
or U1002 (N_1002,N_951,N_918);
or U1003 (N_1003,N_972,N_946);
or U1004 (N_1004,N_958,N_960);
nor U1005 (N_1005,N_943,N_917);
nor U1006 (N_1006,N_915,N_920);
xnor U1007 (N_1007,N_959,N_922);
or U1008 (N_1008,N_968,N_933);
nor U1009 (N_1009,N_938,N_910);
nor U1010 (N_1010,N_926,N_929);
or U1011 (N_1011,N_925,N_927);
nand U1012 (N_1012,N_935,N_954);
and U1013 (N_1013,N_913,N_908);
and U1014 (N_1014,N_911,N_927);
nor U1015 (N_1015,N_959,N_905);
nand U1016 (N_1016,N_961,N_962);
nand U1017 (N_1017,N_915,N_913);
and U1018 (N_1018,N_949,N_951);
and U1019 (N_1019,N_923,N_933);
nand U1020 (N_1020,N_948,N_969);
or U1021 (N_1021,N_910,N_967);
nand U1022 (N_1022,N_957,N_904);
nand U1023 (N_1023,N_963,N_948);
and U1024 (N_1024,N_964,N_959);
and U1025 (N_1025,N_932,N_972);
and U1026 (N_1026,N_907,N_921);
nor U1027 (N_1027,N_934,N_906);
nor U1028 (N_1028,N_943,N_964);
xnor U1029 (N_1029,N_935,N_939);
or U1030 (N_1030,N_940,N_966);
and U1031 (N_1031,N_970,N_921);
and U1032 (N_1032,N_953,N_932);
nor U1033 (N_1033,N_946,N_953);
nor U1034 (N_1034,N_968,N_916);
or U1035 (N_1035,N_919,N_964);
nand U1036 (N_1036,N_902,N_915);
nand U1037 (N_1037,N_965,N_948);
nor U1038 (N_1038,N_913,N_969);
nand U1039 (N_1039,N_948,N_943);
and U1040 (N_1040,N_944,N_942);
or U1041 (N_1041,N_968,N_953);
nor U1042 (N_1042,N_941,N_923);
nor U1043 (N_1043,N_967,N_947);
xor U1044 (N_1044,N_959,N_951);
or U1045 (N_1045,N_912,N_908);
and U1046 (N_1046,N_971,N_900);
nor U1047 (N_1047,N_968,N_909);
or U1048 (N_1048,N_902,N_935);
nor U1049 (N_1049,N_970,N_939);
nor U1050 (N_1050,N_1004,N_985);
and U1051 (N_1051,N_1019,N_1022);
and U1052 (N_1052,N_1037,N_990);
nor U1053 (N_1053,N_1013,N_1017);
and U1054 (N_1054,N_1031,N_1001);
nor U1055 (N_1055,N_1016,N_1038);
or U1056 (N_1056,N_976,N_999);
and U1057 (N_1057,N_1033,N_986);
xor U1058 (N_1058,N_1048,N_1029);
and U1059 (N_1059,N_991,N_1010);
or U1060 (N_1060,N_1021,N_1023);
nand U1061 (N_1061,N_1005,N_1006);
or U1062 (N_1062,N_1018,N_984);
or U1063 (N_1063,N_994,N_1049);
nand U1064 (N_1064,N_996,N_1047);
and U1065 (N_1065,N_997,N_1011);
nor U1066 (N_1066,N_1040,N_988);
nor U1067 (N_1067,N_1000,N_982);
and U1068 (N_1068,N_1030,N_1034);
and U1069 (N_1069,N_1025,N_998);
nor U1070 (N_1070,N_992,N_1046);
and U1071 (N_1071,N_1003,N_1044);
xnor U1072 (N_1072,N_993,N_975);
or U1073 (N_1073,N_979,N_981);
nor U1074 (N_1074,N_1012,N_1035);
nand U1075 (N_1075,N_1007,N_1002);
nor U1076 (N_1076,N_1041,N_1026);
nand U1077 (N_1077,N_983,N_1036);
or U1078 (N_1078,N_989,N_987);
and U1079 (N_1079,N_1009,N_1014);
xor U1080 (N_1080,N_1032,N_1043);
nand U1081 (N_1081,N_1028,N_1024);
xor U1082 (N_1082,N_1015,N_978);
nand U1083 (N_1083,N_1008,N_1042);
nor U1084 (N_1084,N_1020,N_977);
or U1085 (N_1085,N_980,N_1039);
or U1086 (N_1086,N_1045,N_995);
nand U1087 (N_1087,N_1027,N_1049);
or U1088 (N_1088,N_1012,N_1040);
and U1089 (N_1089,N_1044,N_1005);
and U1090 (N_1090,N_1000,N_975);
nand U1091 (N_1091,N_1009,N_1017);
and U1092 (N_1092,N_1034,N_1022);
and U1093 (N_1093,N_1010,N_981);
and U1094 (N_1094,N_1023,N_1024);
and U1095 (N_1095,N_983,N_1029);
nand U1096 (N_1096,N_1044,N_1002);
or U1097 (N_1097,N_990,N_1035);
nand U1098 (N_1098,N_994,N_1024);
nor U1099 (N_1099,N_1008,N_1021);
and U1100 (N_1100,N_1011,N_1021);
nand U1101 (N_1101,N_1024,N_987);
nand U1102 (N_1102,N_1045,N_975);
nor U1103 (N_1103,N_1021,N_986);
or U1104 (N_1104,N_975,N_1022);
and U1105 (N_1105,N_990,N_978);
nand U1106 (N_1106,N_1016,N_1010);
nor U1107 (N_1107,N_1013,N_1042);
and U1108 (N_1108,N_994,N_981);
nand U1109 (N_1109,N_984,N_997);
nor U1110 (N_1110,N_994,N_997);
nand U1111 (N_1111,N_1039,N_1019);
or U1112 (N_1112,N_1047,N_1046);
nor U1113 (N_1113,N_976,N_988);
nor U1114 (N_1114,N_1014,N_991);
and U1115 (N_1115,N_1013,N_1012);
nor U1116 (N_1116,N_1034,N_998);
or U1117 (N_1117,N_1016,N_1008);
and U1118 (N_1118,N_992,N_991);
nand U1119 (N_1119,N_1014,N_983);
or U1120 (N_1120,N_1023,N_999);
and U1121 (N_1121,N_1027,N_987);
and U1122 (N_1122,N_1025,N_1004);
or U1123 (N_1123,N_1034,N_1017);
nor U1124 (N_1124,N_1002,N_1043);
and U1125 (N_1125,N_1057,N_1097);
nor U1126 (N_1126,N_1105,N_1069);
nand U1127 (N_1127,N_1088,N_1121);
nand U1128 (N_1128,N_1124,N_1109);
nand U1129 (N_1129,N_1102,N_1112);
nor U1130 (N_1130,N_1090,N_1098);
nor U1131 (N_1131,N_1083,N_1093);
or U1132 (N_1132,N_1055,N_1052);
nand U1133 (N_1133,N_1117,N_1080);
nand U1134 (N_1134,N_1067,N_1095);
and U1135 (N_1135,N_1077,N_1075);
and U1136 (N_1136,N_1051,N_1110);
or U1137 (N_1137,N_1082,N_1059);
or U1138 (N_1138,N_1123,N_1100);
and U1139 (N_1139,N_1070,N_1061);
nand U1140 (N_1140,N_1074,N_1094);
or U1141 (N_1141,N_1116,N_1084);
nand U1142 (N_1142,N_1068,N_1104);
nand U1143 (N_1143,N_1118,N_1099);
or U1144 (N_1144,N_1087,N_1064);
nand U1145 (N_1145,N_1107,N_1065);
xnor U1146 (N_1146,N_1058,N_1111);
nand U1147 (N_1147,N_1092,N_1056);
nand U1148 (N_1148,N_1053,N_1122);
and U1149 (N_1149,N_1078,N_1108);
nand U1150 (N_1150,N_1101,N_1119);
and U1151 (N_1151,N_1050,N_1113);
nand U1152 (N_1152,N_1089,N_1071);
or U1153 (N_1153,N_1085,N_1066);
and U1154 (N_1154,N_1076,N_1115);
and U1155 (N_1155,N_1062,N_1086);
nor U1156 (N_1156,N_1120,N_1091);
nor U1157 (N_1157,N_1072,N_1054);
nand U1158 (N_1158,N_1063,N_1096);
nor U1159 (N_1159,N_1081,N_1079);
nor U1160 (N_1160,N_1106,N_1073);
and U1161 (N_1161,N_1114,N_1103);
nand U1162 (N_1162,N_1060,N_1090);
or U1163 (N_1163,N_1091,N_1076);
or U1164 (N_1164,N_1056,N_1078);
nor U1165 (N_1165,N_1084,N_1117);
and U1166 (N_1166,N_1075,N_1095);
nand U1167 (N_1167,N_1076,N_1088);
nand U1168 (N_1168,N_1058,N_1117);
nor U1169 (N_1169,N_1091,N_1052);
nand U1170 (N_1170,N_1108,N_1085);
nor U1171 (N_1171,N_1051,N_1082);
and U1172 (N_1172,N_1068,N_1101);
nor U1173 (N_1173,N_1090,N_1080);
and U1174 (N_1174,N_1100,N_1119);
nand U1175 (N_1175,N_1052,N_1058);
nand U1176 (N_1176,N_1084,N_1087);
nor U1177 (N_1177,N_1105,N_1086);
and U1178 (N_1178,N_1103,N_1059);
nor U1179 (N_1179,N_1110,N_1109);
or U1180 (N_1180,N_1083,N_1094);
nand U1181 (N_1181,N_1123,N_1103);
and U1182 (N_1182,N_1117,N_1071);
xnor U1183 (N_1183,N_1080,N_1073);
or U1184 (N_1184,N_1061,N_1090);
nor U1185 (N_1185,N_1079,N_1082);
nor U1186 (N_1186,N_1106,N_1084);
nor U1187 (N_1187,N_1121,N_1075);
and U1188 (N_1188,N_1085,N_1052);
nand U1189 (N_1189,N_1118,N_1103);
or U1190 (N_1190,N_1100,N_1077);
nand U1191 (N_1191,N_1116,N_1100);
or U1192 (N_1192,N_1055,N_1090);
and U1193 (N_1193,N_1108,N_1088);
nand U1194 (N_1194,N_1072,N_1077);
or U1195 (N_1195,N_1121,N_1086);
and U1196 (N_1196,N_1115,N_1077);
nand U1197 (N_1197,N_1093,N_1075);
and U1198 (N_1198,N_1089,N_1110);
nor U1199 (N_1199,N_1105,N_1123);
nand U1200 (N_1200,N_1194,N_1145);
nand U1201 (N_1201,N_1129,N_1177);
nand U1202 (N_1202,N_1187,N_1166);
nand U1203 (N_1203,N_1157,N_1134);
and U1204 (N_1204,N_1173,N_1197);
nand U1205 (N_1205,N_1127,N_1144);
nand U1206 (N_1206,N_1125,N_1161);
and U1207 (N_1207,N_1169,N_1138);
nor U1208 (N_1208,N_1151,N_1181);
or U1209 (N_1209,N_1179,N_1141);
nor U1210 (N_1210,N_1130,N_1153);
nand U1211 (N_1211,N_1176,N_1188);
nand U1212 (N_1212,N_1140,N_1147);
nand U1213 (N_1213,N_1193,N_1159);
or U1214 (N_1214,N_1178,N_1171);
nor U1215 (N_1215,N_1128,N_1150);
and U1216 (N_1216,N_1184,N_1149);
nand U1217 (N_1217,N_1155,N_1190);
nand U1218 (N_1218,N_1170,N_1135);
nor U1219 (N_1219,N_1175,N_1180);
nand U1220 (N_1220,N_1167,N_1126);
nand U1221 (N_1221,N_1196,N_1146);
nand U1222 (N_1222,N_1164,N_1199);
nand U1223 (N_1223,N_1191,N_1148);
and U1224 (N_1224,N_1186,N_1156);
nand U1225 (N_1225,N_1154,N_1131);
nor U1226 (N_1226,N_1165,N_1189);
nor U1227 (N_1227,N_1137,N_1174);
nand U1228 (N_1228,N_1172,N_1158);
nand U1229 (N_1229,N_1142,N_1133);
and U1230 (N_1230,N_1198,N_1168);
nor U1231 (N_1231,N_1143,N_1162);
and U1232 (N_1232,N_1132,N_1185);
and U1233 (N_1233,N_1139,N_1195);
nand U1234 (N_1234,N_1160,N_1152);
or U1235 (N_1235,N_1192,N_1183);
nor U1236 (N_1236,N_1182,N_1136);
or U1237 (N_1237,N_1163,N_1130);
nor U1238 (N_1238,N_1130,N_1175);
nand U1239 (N_1239,N_1174,N_1129);
and U1240 (N_1240,N_1141,N_1176);
nor U1241 (N_1241,N_1187,N_1145);
and U1242 (N_1242,N_1159,N_1153);
nor U1243 (N_1243,N_1186,N_1171);
and U1244 (N_1244,N_1165,N_1178);
and U1245 (N_1245,N_1176,N_1168);
and U1246 (N_1246,N_1177,N_1142);
and U1247 (N_1247,N_1131,N_1173);
nor U1248 (N_1248,N_1146,N_1161);
nand U1249 (N_1249,N_1158,N_1183);
nor U1250 (N_1250,N_1141,N_1157);
and U1251 (N_1251,N_1182,N_1154);
nor U1252 (N_1252,N_1158,N_1184);
nor U1253 (N_1253,N_1125,N_1136);
nand U1254 (N_1254,N_1167,N_1130);
nor U1255 (N_1255,N_1180,N_1199);
and U1256 (N_1256,N_1137,N_1153);
and U1257 (N_1257,N_1198,N_1150);
nand U1258 (N_1258,N_1131,N_1126);
xnor U1259 (N_1259,N_1196,N_1193);
nand U1260 (N_1260,N_1140,N_1177);
or U1261 (N_1261,N_1143,N_1146);
or U1262 (N_1262,N_1198,N_1125);
or U1263 (N_1263,N_1161,N_1191);
and U1264 (N_1264,N_1135,N_1153);
nor U1265 (N_1265,N_1167,N_1198);
or U1266 (N_1266,N_1129,N_1194);
and U1267 (N_1267,N_1185,N_1135);
nor U1268 (N_1268,N_1193,N_1198);
nand U1269 (N_1269,N_1163,N_1188);
or U1270 (N_1270,N_1156,N_1184);
nor U1271 (N_1271,N_1141,N_1185);
and U1272 (N_1272,N_1171,N_1133);
or U1273 (N_1273,N_1156,N_1151);
nor U1274 (N_1274,N_1156,N_1193);
or U1275 (N_1275,N_1265,N_1240);
and U1276 (N_1276,N_1207,N_1266);
nor U1277 (N_1277,N_1225,N_1203);
and U1278 (N_1278,N_1252,N_1258);
or U1279 (N_1279,N_1220,N_1245);
nor U1280 (N_1280,N_1218,N_1257);
and U1281 (N_1281,N_1224,N_1270);
nand U1282 (N_1282,N_1271,N_1204);
and U1283 (N_1283,N_1201,N_1211);
and U1284 (N_1284,N_1241,N_1248);
nor U1285 (N_1285,N_1230,N_1221);
nand U1286 (N_1286,N_1244,N_1261);
and U1287 (N_1287,N_1223,N_1234);
and U1288 (N_1288,N_1259,N_1216);
nor U1289 (N_1289,N_1226,N_1274);
and U1290 (N_1290,N_1254,N_1233);
nor U1291 (N_1291,N_1227,N_1267);
nor U1292 (N_1292,N_1229,N_1235);
nor U1293 (N_1293,N_1242,N_1262);
nand U1294 (N_1294,N_1209,N_1236);
nor U1295 (N_1295,N_1200,N_1251);
nand U1296 (N_1296,N_1250,N_1214);
or U1297 (N_1297,N_1217,N_1222);
and U1298 (N_1298,N_1268,N_1255);
nand U1299 (N_1299,N_1219,N_1213);
nor U1300 (N_1300,N_1272,N_1246);
nand U1301 (N_1301,N_1273,N_1247);
or U1302 (N_1302,N_1249,N_1205);
or U1303 (N_1303,N_1264,N_1206);
or U1304 (N_1304,N_1210,N_1237);
xnor U1305 (N_1305,N_1243,N_1238);
nand U1306 (N_1306,N_1260,N_1202);
xor U1307 (N_1307,N_1256,N_1208);
or U1308 (N_1308,N_1212,N_1253);
xor U1309 (N_1309,N_1263,N_1269);
and U1310 (N_1310,N_1215,N_1232);
or U1311 (N_1311,N_1231,N_1228);
nor U1312 (N_1312,N_1239,N_1238);
nand U1313 (N_1313,N_1261,N_1250);
nor U1314 (N_1314,N_1271,N_1250);
or U1315 (N_1315,N_1243,N_1268);
nor U1316 (N_1316,N_1220,N_1239);
nor U1317 (N_1317,N_1215,N_1269);
nand U1318 (N_1318,N_1223,N_1201);
and U1319 (N_1319,N_1224,N_1219);
or U1320 (N_1320,N_1221,N_1218);
or U1321 (N_1321,N_1240,N_1237);
nand U1322 (N_1322,N_1206,N_1204);
nor U1323 (N_1323,N_1205,N_1268);
nor U1324 (N_1324,N_1225,N_1226);
or U1325 (N_1325,N_1211,N_1263);
nand U1326 (N_1326,N_1200,N_1263);
nand U1327 (N_1327,N_1266,N_1216);
and U1328 (N_1328,N_1259,N_1258);
nor U1329 (N_1329,N_1209,N_1261);
or U1330 (N_1330,N_1266,N_1235);
xnor U1331 (N_1331,N_1214,N_1268);
and U1332 (N_1332,N_1256,N_1272);
nor U1333 (N_1333,N_1216,N_1200);
and U1334 (N_1334,N_1213,N_1233);
nor U1335 (N_1335,N_1252,N_1210);
and U1336 (N_1336,N_1217,N_1237);
and U1337 (N_1337,N_1257,N_1224);
or U1338 (N_1338,N_1213,N_1203);
or U1339 (N_1339,N_1247,N_1244);
nor U1340 (N_1340,N_1262,N_1224);
nor U1341 (N_1341,N_1220,N_1246);
nand U1342 (N_1342,N_1223,N_1263);
nand U1343 (N_1343,N_1200,N_1271);
nand U1344 (N_1344,N_1201,N_1274);
or U1345 (N_1345,N_1229,N_1205);
nand U1346 (N_1346,N_1234,N_1235);
xor U1347 (N_1347,N_1260,N_1262);
nor U1348 (N_1348,N_1234,N_1243);
or U1349 (N_1349,N_1222,N_1211);
or U1350 (N_1350,N_1286,N_1303);
and U1351 (N_1351,N_1347,N_1333);
or U1352 (N_1352,N_1329,N_1298);
or U1353 (N_1353,N_1339,N_1322);
xnor U1354 (N_1354,N_1314,N_1335);
nor U1355 (N_1355,N_1287,N_1295);
and U1356 (N_1356,N_1338,N_1330);
nand U1357 (N_1357,N_1316,N_1324);
or U1358 (N_1358,N_1307,N_1315);
or U1359 (N_1359,N_1275,N_1340);
nor U1360 (N_1360,N_1280,N_1323);
nand U1361 (N_1361,N_1334,N_1304);
or U1362 (N_1362,N_1299,N_1313);
and U1363 (N_1363,N_1344,N_1310);
nor U1364 (N_1364,N_1301,N_1281);
nand U1365 (N_1365,N_1331,N_1279);
nor U1366 (N_1366,N_1285,N_1327);
or U1367 (N_1367,N_1348,N_1342);
or U1368 (N_1368,N_1276,N_1312);
nor U1369 (N_1369,N_1332,N_1319);
nor U1370 (N_1370,N_1308,N_1282);
xor U1371 (N_1371,N_1320,N_1292);
nand U1372 (N_1372,N_1311,N_1288);
and U1373 (N_1373,N_1326,N_1337);
and U1374 (N_1374,N_1277,N_1349);
nor U1375 (N_1375,N_1317,N_1343);
and U1376 (N_1376,N_1321,N_1289);
or U1377 (N_1377,N_1284,N_1302);
and U1378 (N_1378,N_1296,N_1290);
nor U1379 (N_1379,N_1346,N_1309);
and U1380 (N_1380,N_1294,N_1341);
and U1381 (N_1381,N_1336,N_1345);
or U1382 (N_1382,N_1306,N_1297);
or U1383 (N_1383,N_1283,N_1328);
nor U1384 (N_1384,N_1305,N_1318);
and U1385 (N_1385,N_1325,N_1278);
nand U1386 (N_1386,N_1293,N_1300);
nand U1387 (N_1387,N_1291,N_1306);
nand U1388 (N_1388,N_1342,N_1330);
and U1389 (N_1389,N_1295,N_1338);
nand U1390 (N_1390,N_1346,N_1326);
nor U1391 (N_1391,N_1341,N_1338);
nand U1392 (N_1392,N_1332,N_1349);
nor U1393 (N_1393,N_1290,N_1345);
or U1394 (N_1394,N_1338,N_1276);
nand U1395 (N_1395,N_1288,N_1284);
and U1396 (N_1396,N_1286,N_1279);
and U1397 (N_1397,N_1277,N_1324);
and U1398 (N_1398,N_1285,N_1320);
and U1399 (N_1399,N_1281,N_1295);
nand U1400 (N_1400,N_1324,N_1279);
nor U1401 (N_1401,N_1323,N_1336);
xor U1402 (N_1402,N_1308,N_1338);
nor U1403 (N_1403,N_1342,N_1294);
xor U1404 (N_1404,N_1332,N_1348);
nand U1405 (N_1405,N_1310,N_1277);
nand U1406 (N_1406,N_1284,N_1327);
and U1407 (N_1407,N_1348,N_1291);
nand U1408 (N_1408,N_1325,N_1303);
or U1409 (N_1409,N_1286,N_1315);
or U1410 (N_1410,N_1301,N_1329);
or U1411 (N_1411,N_1346,N_1340);
nand U1412 (N_1412,N_1300,N_1336);
nor U1413 (N_1413,N_1319,N_1287);
or U1414 (N_1414,N_1323,N_1326);
nand U1415 (N_1415,N_1283,N_1275);
xnor U1416 (N_1416,N_1332,N_1314);
nand U1417 (N_1417,N_1337,N_1277);
nor U1418 (N_1418,N_1286,N_1288);
nor U1419 (N_1419,N_1280,N_1320);
nand U1420 (N_1420,N_1323,N_1285);
nor U1421 (N_1421,N_1288,N_1339);
nor U1422 (N_1422,N_1312,N_1323);
or U1423 (N_1423,N_1309,N_1301);
or U1424 (N_1424,N_1335,N_1318);
or U1425 (N_1425,N_1391,N_1411);
and U1426 (N_1426,N_1413,N_1382);
nor U1427 (N_1427,N_1372,N_1409);
nand U1428 (N_1428,N_1424,N_1367);
and U1429 (N_1429,N_1408,N_1400);
or U1430 (N_1430,N_1361,N_1395);
and U1431 (N_1431,N_1404,N_1373);
or U1432 (N_1432,N_1388,N_1379);
nor U1433 (N_1433,N_1397,N_1368);
and U1434 (N_1434,N_1358,N_1351);
and U1435 (N_1435,N_1393,N_1378);
nor U1436 (N_1436,N_1376,N_1410);
or U1437 (N_1437,N_1418,N_1377);
and U1438 (N_1438,N_1360,N_1399);
and U1439 (N_1439,N_1370,N_1403);
or U1440 (N_1440,N_1420,N_1421);
nor U1441 (N_1441,N_1354,N_1392);
nor U1442 (N_1442,N_1383,N_1419);
or U1443 (N_1443,N_1359,N_1381);
nand U1444 (N_1444,N_1380,N_1385);
nand U1445 (N_1445,N_1366,N_1375);
or U1446 (N_1446,N_1374,N_1394);
nor U1447 (N_1447,N_1364,N_1422);
nor U1448 (N_1448,N_1356,N_1398);
nand U1449 (N_1449,N_1384,N_1396);
or U1450 (N_1450,N_1401,N_1406);
nor U1451 (N_1451,N_1402,N_1386);
nor U1452 (N_1452,N_1415,N_1362);
or U1453 (N_1453,N_1407,N_1412);
nor U1454 (N_1454,N_1371,N_1416);
nor U1455 (N_1455,N_1405,N_1369);
or U1456 (N_1456,N_1352,N_1390);
nand U1457 (N_1457,N_1389,N_1350);
nand U1458 (N_1458,N_1363,N_1423);
and U1459 (N_1459,N_1357,N_1365);
nor U1460 (N_1460,N_1417,N_1353);
nor U1461 (N_1461,N_1387,N_1414);
or U1462 (N_1462,N_1355,N_1361);
nand U1463 (N_1463,N_1420,N_1377);
xor U1464 (N_1464,N_1365,N_1366);
or U1465 (N_1465,N_1379,N_1408);
xor U1466 (N_1466,N_1374,N_1350);
or U1467 (N_1467,N_1420,N_1402);
nor U1468 (N_1468,N_1364,N_1407);
nand U1469 (N_1469,N_1419,N_1378);
nor U1470 (N_1470,N_1350,N_1362);
or U1471 (N_1471,N_1379,N_1381);
nor U1472 (N_1472,N_1407,N_1384);
xor U1473 (N_1473,N_1358,N_1404);
nand U1474 (N_1474,N_1397,N_1369);
and U1475 (N_1475,N_1368,N_1417);
nor U1476 (N_1476,N_1385,N_1352);
or U1477 (N_1477,N_1421,N_1424);
nor U1478 (N_1478,N_1413,N_1392);
nor U1479 (N_1479,N_1420,N_1351);
xnor U1480 (N_1480,N_1357,N_1401);
xor U1481 (N_1481,N_1394,N_1371);
nor U1482 (N_1482,N_1396,N_1361);
or U1483 (N_1483,N_1370,N_1365);
nor U1484 (N_1484,N_1370,N_1412);
nand U1485 (N_1485,N_1408,N_1354);
nand U1486 (N_1486,N_1406,N_1363);
or U1487 (N_1487,N_1359,N_1354);
nand U1488 (N_1488,N_1408,N_1421);
or U1489 (N_1489,N_1356,N_1400);
nand U1490 (N_1490,N_1362,N_1360);
and U1491 (N_1491,N_1392,N_1407);
nand U1492 (N_1492,N_1419,N_1362);
and U1493 (N_1493,N_1371,N_1351);
or U1494 (N_1494,N_1366,N_1395);
nor U1495 (N_1495,N_1352,N_1388);
or U1496 (N_1496,N_1363,N_1413);
and U1497 (N_1497,N_1352,N_1421);
nand U1498 (N_1498,N_1383,N_1400);
and U1499 (N_1499,N_1413,N_1385);
nor U1500 (N_1500,N_1498,N_1446);
and U1501 (N_1501,N_1463,N_1434);
nand U1502 (N_1502,N_1426,N_1428);
and U1503 (N_1503,N_1431,N_1451);
nand U1504 (N_1504,N_1474,N_1475);
nand U1505 (N_1505,N_1488,N_1464);
and U1506 (N_1506,N_1437,N_1476);
or U1507 (N_1507,N_1441,N_1489);
nand U1508 (N_1508,N_1465,N_1471);
nor U1509 (N_1509,N_1462,N_1449);
nor U1510 (N_1510,N_1496,N_1461);
or U1511 (N_1511,N_1448,N_1433);
and U1512 (N_1512,N_1478,N_1468);
nand U1513 (N_1513,N_1479,N_1499);
or U1514 (N_1514,N_1460,N_1486);
or U1515 (N_1515,N_1454,N_1443);
or U1516 (N_1516,N_1438,N_1495);
or U1517 (N_1517,N_1481,N_1491);
nand U1518 (N_1518,N_1490,N_1445);
or U1519 (N_1519,N_1477,N_1456);
and U1520 (N_1520,N_1497,N_1485);
and U1521 (N_1521,N_1484,N_1473);
and U1522 (N_1522,N_1425,N_1436);
xor U1523 (N_1523,N_1470,N_1487);
nand U1524 (N_1524,N_1453,N_1455);
xnor U1525 (N_1525,N_1427,N_1452);
nor U1526 (N_1526,N_1429,N_1472);
or U1527 (N_1527,N_1480,N_1430);
nor U1528 (N_1528,N_1450,N_1457);
or U1529 (N_1529,N_1482,N_1439);
and U1530 (N_1530,N_1458,N_1493);
nand U1531 (N_1531,N_1466,N_1459);
or U1532 (N_1532,N_1442,N_1447);
or U1533 (N_1533,N_1440,N_1494);
and U1534 (N_1534,N_1432,N_1467);
or U1535 (N_1535,N_1435,N_1444);
nor U1536 (N_1536,N_1483,N_1469);
and U1537 (N_1537,N_1492,N_1459);
and U1538 (N_1538,N_1494,N_1455);
or U1539 (N_1539,N_1435,N_1499);
and U1540 (N_1540,N_1430,N_1451);
and U1541 (N_1541,N_1480,N_1487);
and U1542 (N_1542,N_1464,N_1442);
nor U1543 (N_1543,N_1485,N_1491);
nand U1544 (N_1544,N_1492,N_1444);
nor U1545 (N_1545,N_1498,N_1474);
nand U1546 (N_1546,N_1472,N_1482);
nand U1547 (N_1547,N_1496,N_1490);
nand U1548 (N_1548,N_1467,N_1476);
or U1549 (N_1549,N_1499,N_1430);
or U1550 (N_1550,N_1461,N_1447);
or U1551 (N_1551,N_1473,N_1448);
nand U1552 (N_1552,N_1470,N_1452);
nand U1553 (N_1553,N_1454,N_1471);
and U1554 (N_1554,N_1433,N_1449);
and U1555 (N_1555,N_1482,N_1454);
and U1556 (N_1556,N_1450,N_1487);
nand U1557 (N_1557,N_1462,N_1459);
nand U1558 (N_1558,N_1432,N_1453);
nand U1559 (N_1559,N_1432,N_1478);
nor U1560 (N_1560,N_1441,N_1464);
and U1561 (N_1561,N_1490,N_1436);
or U1562 (N_1562,N_1427,N_1466);
nand U1563 (N_1563,N_1466,N_1436);
and U1564 (N_1564,N_1497,N_1495);
nand U1565 (N_1565,N_1457,N_1453);
nor U1566 (N_1566,N_1475,N_1446);
xnor U1567 (N_1567,N_1455,N_1477);
nand U1568 (N_1568,N_1497,N_1434);
xor U1569 (N_1569,N_1495,N_1460);
nor U1570 (N_1570,N_1426,N_1478);
nand U1571 (N_1571,N_1427,N_1486);
or U1572 (N_1572,N_1475,N_1496);
and U1573 (N_1573,N_1433,N_1443);
and U1574 (N_1574,N_1476,N_1484);
and U1575 (N_1575,N_1500,N_1548);
and U1576 (N_1576,N_1530,N_1569);
nand U1577 (N_1577,N_1502,N_1568);
or U1578 (N_1578,N_1540,N_1503);
nand U1579 (N_1579,N_1553,N_1551);
and U1580 (N_1580,N_1556,N_1574);
and U1581 (N_1581,N_1504,N_1516);
and U1582 (N_1582,N_1537,N_1546);
nand U1583 (N_1583,N_1533,N_1506);
nor U1584 (N_1584,N_1550,N_1526);
and U1585 (N_1585,N_1567,N_1521);
nor U1586 (N_1586,N_1542,N_1563);
nand U1587 (N_1587,N_1527,N_1534);
nand U1588 (N_1588,N_1572,N_1543);
nand U1589 (N_1589,N_1519,N_1528);
and U1590 (N_1590,N_1512,N_1559);
or U1591 (N_1591,N_1549,N_1532);
nand U1592 (N_1592,N_1545,N_1547);
or U1593 (N_1593,N_1513,N_1541);
and U1594 (N_1594,N_1573,N_1562);
nor U1595 (N_1595,N_1511,N_1555);
or U1596 (N_1596,N_1531,N_1505);
and U1597 (N_1597,N_1560,N_1518);
and U1598 (N_1598,N_1524,N_1509);
and U1599 (N_1599,N_1523,N_1501);
and U1600 (N_1600,N_1514,N_1565);
and U1601 (N_1601,N_1507,N_1508);
and U1602 (N_1602,N_1529,N_1535);
or U1603 (N_1603,N_1558,N_1552);
or U1604 (N_1604,N_1525,N_1510);
nand U1605 (N_1605,N_1539,N_1520);
nand U1606 (N_1606,N_1564,N_1571);
and U1607 (N_1607,N_1517,N_1554);
nor U1608 (N_1608,N_1538,N_1566);
and U1609 (N_1609,N_1570,N_1522);
nor U1610 (N_1610,N_1515,N_1557);
and U1611 (N_1611,N_1536,N_1561);
nand U1612 (N_1612,N_1544,N_1522);
nor U1613 (N_1613,N_1537,N_1547);
or U1614 (N_1614,N_1526,N_1542);
nor U1615 (N_1615,N_1530,N_1535);
and U1616 (N_1616,N_1520,N_1541);
nor U1617 (N_1617,N_1561,N_1528);
and U1618 (N_1618,N_1535,N_1537);
or U1619 (N_1619,N_1554,N_1551);
nand U1620 (N_1620,N_1515,N_1516);
and U1621 (N_1621,N_1544,N_1500);
and U1622 (N_1622,N_1548,N_1556);
nor U1623 (N_1623,N_1509,N_1534);
nor U1624 (N_1624,N_1525,N_1521);
nand U1625 (N_1625,N_1573,N_1552);
or U1626 (N_1626,N_1505,N_1538);
nor U1627 (N_1627,N_1506,N_1561);
nand U1628 (N_1628,N_1562,N_1504);
and U1629 (N_1629,N_1509,N_1508);
nand U1630 (N_1630,N_1540,N_1506);
and U1631 (N_1631,N_1555,N_1572);
and U1632 (N_1632,N_1549,N_1539);
or U1633 (N_1633,N_1509,N_1571);
or U1634 (N_1634,N_1517,N_1515);
nand U1635 (N_1635,N_1522,N_1557);
nand U1636 (N_1636,N_1503,N_1511);
nor U1637 (N_1637,N_1528,N_1521);
or U1638 (N_1638,N_1520,N_1555);
nor U1639 (N_1639,N_1523,N_1545);
nor U1640 (N_1640,N_1555,N_1562);
nand U1641 (N_1641,N_1563,N_1500);
nor U1642 (N_1642,N_1513,N_1570);
nor U1643 (N_1643,N_1544,N_1502);
nand U1644 (N_1644,N_1558,N_1534);
and U1645 (N_1645,N_1501,N_1565);
or U1646 (N_1646,N_1527,N_1530);
nand U1647 (N_1647,N_1553,N_1554);
and U1648 (N_1648,N_1535,N_1536);
nand U1649 (N_1649,N_1526,N_1544);
nor U1650 (N_1650,N_1635,N_1579);
nand U1651 (N_1651,N_1591,N_1584);
and U1652 (N_1652,N_1641,N_1588);
nor U1653 (N_1653,N_1599,N_1592);
nand U1654 (N_1654,N_1645,N_1623);
and U1655 (N_1655,N_1642,N_1622);
and U1656 (N_1656,N_1644,N_1606);
and U1657 (N_1657,N_1616,N_1624);
xor U1658 (N_1658,N_1575,N_1643);
nor U1659 (N_1659,N_1583,N_1576);
or U1660 (N_1660,N_1603,N_1614);
nor U1661 (N_1661,N_1581,N_1621);
nor U1662 (N_1662,N_1613,N_1646);
nand U1663 (N_1663,N_1600,N_1605);
or U1664 (N_1664,N_1595,N_1577);
nor U1665 (N_1665,N_1582,N_1596);
nand U1666 (N_1666,N_1619,N_1632);
nand U1667 (N_1667,N_1629,N_1604);
nor U1668 (N_1668,N_1634,N_1627);
and U1669 (N_1669,N_1589,N_1607);
nand U1670 (N_1670,N_1640,N_1580);
xnor U1671 (N_1671,N_1648,N_1585);
and U1672 (N_1672,N_1638,N_1630);
nand U1673 (N_1673,N_1578,N_1617);
nand U1674 (N_1674,N_1625,N_1628);
and U1675 (N_1675,N_1637,N_1597);
or U1676 (N_1676,N_1594,N_1608);
nand U1677 (N_1677,N_1626,N_1609);
nor U1678 (N_1678,N_1633,N_1620);
nor U1679 (N_1679,N_1602,N_1611);
nand U1680 (N_1680,N_1610,N_1612);
nand U1681 (N_1681,N_1587,N_1601);
nor U1682 (N_1682,N_1647,N_1649);
or U1683 (N_1683,N_1590,N_1631);
or U1684 (N_1684,N_1639,N_1618);
and U1685 (N_1685,N_1586,N_1636);
or U1686 (N_1686,N_1593,N_1598);
xnor U1687 (N_1687,N_1615,N_1627);
and U1688 (N_1688,N_1627,N_1579);
or U1689 (N_1689,N_1601,N_1606);
nor U1690 (N_1690,N_1586,N_1581);
nand U1691 (N_1691,N_1584,N_1598);
or U1692 (N_1692,N_1644,N_1638);
nand U1693 (N_1693,N_1585,N_1578);
and U1694 (N_1694,N_1628,N_1598);
or U1695 (N_1695,N_1611,N_1582);
nand U1696 (N_1696,N_1611,N_1632);
or U1697 (N_1697,N_1592,N_1629);
xor U1698 (N_1698,N_1607,N_1629);
nand U1699 (N_1699,N_1610,N_1597);
nand U1700 (N_1700,N_1586,N_1606);
nor U1701 (N_1701,N_1627,N_1608);
or U1702 (N_1702,N_1575,N_1618);
and U1703 (N_1703,N_1596,N_1647);
nand U1704 (N_1704,N_1631,N_1637);
and U1705 (N_1705,N_1592,N_1644);
or U1706 (N_1706,N_1645,N_1603);
nand U1707 (N_1707,N_1604,N_1645);
or U1708 (N_1708,N_1597,N_1593);
and U1709 (N_1709,N_1618,N_1592);
or U1710 (N_1710,N_1646,N_1617);
or U1711 (N_1711,N_1614,N_1619);
and U1712 (N_1712,N_1624,N_1633);
nor U1713 (N_1713,N_1599,N_1619);
and U1714 (N_1714,N_1581,N_1603);
nand U1715 (N_1715,N_1629,N_1601);
nand U1716 (N_1716,N_1630,N_1632);
and U1717 (N_1717,N_1631,N_1634);
nand U1718 (N_1718,N_1585,N_1576);
xnor U1719 (N_1719,N_1611,N_1641);
nand U1720 (N_1720,N_1588,N_1604);
nor U1721 (N_1721,N_1615,N_1595);
nand U1722 (N_1722,N_1603,N_1619);
xor U1723 (N_1723,N_1598,N_1636);
nor U1724 (N_1724,N_1591,N_1600);
nand U1725 (N_1725,N_1715,N_1700);
or U1726 (N_1726,N_1651,N_1705);
nor U1727 (N_1727,N_1713,N_1662);
or U1728 (N_1728,N_1692,N_1685);
nand U1729 (N_1729,N_1693,N_1683);
or U1730 (N_1730,N_1711,N_1664);
nor U1731 (N_1731,N_1709,N_1708);
nor U1732 (N_1732,N_1722,N_1659);
nand U1733 (N_1733,N_1707,N_1714);
nand U1734 (N_1734,N_1704,N_1691);
nor U1735 (N_1735,N_1703,N_1696);
and U1736 (N_1736,N_1670,N_1697);
or U1737 (N_1737,N_1690,N_1668);
nand U1738 (N_1738,N_1702,N_1684);
or U1739 (N_1739,N_1723,N_1706);
and U1740 (N_1740,N_1653,N_1712);
nor U1741 (N_1741,N_1676,N_1681);
nand U1742 (N_1742,N_1694,N_1717);
and U1743 (N_1743,N_1671,N_1695);
or U1744 (N_1744,N_1699,N_1701);
or U1745 (N_1745,N_1688,N_1661);
or U1746 (N_1746,N_1679,N_1655);
nand U1747 (N_1747,N_1665,N_1675);
nand U1748 (N_1748,N_1652,N_1720);
or U1749 (N_1749,N_1687,N_1657);
or U1750 (N_1750,N_1654,N_1650);
and U1751 (N_1751,N_1673,N_1666);
nor U1752 (N_1752,N_1667,N_1669);
nor U1753 (N_1753,N_1686,N_1719);
and U1754 (N_1754,N_1672,N_1674);
and U1755 (N_1755,N_1718,N_1724);
or U1756 (N_1756,N_1682,N_1656);
nor U1757 (N_1757,N_1721,N_1658);
or U1758 (N_1758,N_1710,N_1680);
nand U1759 (N_1759,N_1677,N_1660);
or U1760 (N_1760,N_1716,N_1698);
nand U1761 (N_1761,N_1678,N_1663);
and U1762 (N_1762,N_1689,N_1718);
nor U1763 (N_1763,N_1723,N_1679);
nor U1764 (N_1764,N_1674,N_1700);
or U1765 (N_1765,N_1688,N_1686);
nand U1766 (N_1766,N_1690,N_1688);
or U1767 (N_1767,N_1656,N_1650);
or U1768 (N_1768,N_1710,N_1723);
or U1769 (N_1769,N_1704,N_1720);
or U1770 (N_1770,N_1669,N_1671);
or U1771 (N_1771,N_1695,N_1718);
or U1772 (N_1772,N_1669,N_1689);
or U1773 (N_1773,N_1709,N_1718);
nor U1774 (N_1774,N_1679,N_1656);
nor U1775 (N_1775,N_1655,N_1714);
or U1776 (N_1776,N_1668,N_1672);
and U1777 (N_1777,N_1666,N_1707);
nor U1778 (N_1778,N_1707,N_1700);
nand U1779 (N_1779,N_1695,N_1716);
nand U1780 (N_1780,N_1711,N_1653);
nand U1781 (N_1781,N_1651,N_1673);
or U1782 (N_1782,N_1677,N_1718);
nand U1783 (N_1783,N_1687,N_1713);
nand U1784 (N_1784,N_1670,N_1708);
xnor U1785 (N_1785,N_1683,N_1669);
nor U1786 (N_1786,N_1717,N_1689);
nor U1787 (N_1787,N_1698,N_1683);
nand U1788 (N_1788,N_1707,N_1658);
or U1789 (N_1789,N_1670,N_1661);
nor U1790 (N_1790,N_1706,N_1700);
nand U1791 (N_1791,N_1720,N_1679);
or U1792 (N_1792,N_1690,N_1703);
and U1793 (N_1793,N_1686,N_1652);
nor U1794 (N_1794,N_1702,N_1703);
and U1795 (N_1795,N_1659,N_1666);
or U1796 (N_1796,N_1690,N_1700);
or U1797 (N_1797,N_1669,N_1659);
or U1798 (N_1798,N_1672,N_1671);
and U1799 (N_1799,N_1671,N_1650);
nor U1800 (N_1800,N_1746,N_1763);
and U1801 (N_1801,N_1786,N_1750);
or U1802 (N_1802,N_1728,N_1731);
nor U1803 (N_1803,N_1767,N_1742);
or U1804 (N_1804,N_1735,N_1759);
nor U1805 (N_1805,N_1754,N_1730);
and U1806 (N_1806,N_1792,N_1797);
nor U1807 (N_1807,N_1782,N_1776);
or U1808 (N_1808,N_1785,N_1762);
nand U1809 (N_1809,N_1749,N_1769);
nand U1810 (N_1810,N_1780,N_1787);
nor U1811 (N_1811,N_1733,N_1745);
or U1812 (N_1812,N_1765,N_1778);
nor U1813 (N_1813,N_1751,N_1737);
nor U1814 (N_1814,N_1795,N_1779);
or U1815 (N_1815,N_1784,N_1740);
and U1816 (N_1816,N_1729,N_1756);
nor U1817 (N_1817,N_1771,N_1732);
nand U1818 (N_1818,N_1741,N_1770);
or U1819 (N_1819,N_1748,N_1725);
or U1820 (N_1820,N_1747,N_1753);
nand U1821 (N_1821,N_1772,N_1790);
nor U1822 (N_1822,N_1789,N_1758);
and U1823 (N_1823,N_1744,N_1739);
nor U1824 (N_1824,N_1734,N_1764);
and U1825 (N_1825,N_1773,N_1761);
and U1826 (N_1826,N_1757,N_1791);
nor U1827 (N_1827,N_1755,N_1794);
and U1828 (N_1828,N_1727,N_1752);
and U1829 (N_1829,N_1774,N_1775);
nor U1830 (N_1830,N_1726,N_1760);
nand U1831 (N_1831,N_1777,N_1796);
nand U1832 (N_1832,N_1766,N_1743);
nor U1833 (N_1833,N_1799,N_1793);
nand U1834 (N_1834,N_1783,N_1738);
or U1835 (N_1835,N_1798,N_1768);
and U1836 (N_1836,N_1736,N_1788);
or U1837 (N_1837,N_1781,N_1760);
nor U1838 (N_1838,N_1786,N_1755);
nor U1839 (N_1839,N_1745,N_1732);
nor U1840 (N_1840,N_1754,N_1799);
nor U1841 (N_1841,N_1784,N_1776);
xor U1842 (N_1842,N_1777,N_1750);
nor U1843 (N_1843,N_1767,N_1792);
nand U1844 (N_1844,N_1792,N_1778);
or U1845 (N_1845,N_1749,N_1793);
nand U1846 (N_1846,N_1778,N_1726);
nand U1847 (N_1847,N_1749,N_1730);
or U1848 (N_1848,N_1763,N_1748);
nand U1849 (N_1849,N_1728,N_1737);
nor U1850 (N_1850,N_1787,N_1743);
nand U1851 (N_1851,N_1783,N_1754);
nor U1852 (N_1852,N_1725,N_1740);
nor U1853 (N_1853,N_1752,N_1736);
nand U1854 (N_1854,N_1777,N_1778);
and U1855 (N_1855,N_1754,N_1729);
nand U1856 (N_1856,N_1744,N_1780);
and U1857 (N_1857,N_1753,N_1778);
nor U1858 (N_1858,N_1769,N_1740);
and U1859 (N_1859,N_1772,N_1783);
or U1860 (N_1860,N_1765,N_1742);
and U1861 (N_1861,N_1757,N_1758);
nand U1862 (N_1862,N_1752,N_1759);
or U1863 (N_1863,N_1734,N_1751);
nand U1864 (N_1864,N_1794,N_1778);
and U1865 (N_1865,N_1753,N_1786);
or U1866 (N_1866,N_1728,N_1739);
nor U1867 (N_1867,N_1783,N_1753);
nor U1868 (N_1868,N_1726,N_1727);
or U1869 (N_1869,N_1749,N_1758);
and U1870 (N_1870,N_1747,N_1733);
and U1871 (N_1871,N_1773,N_1727);
and U1872 (N_1872,N_1778,N_1766);
or U1873 (N_1873,N_1766,N_1775);
nand U1874 (N_1874,N_1740,N_1770);
nor U1875 (N_1875,N_1872,N_1832);
nand U1876 (N_1876,N_1812,N_1800);
and U1877 (N_1877,N_1840,N_1846);
nor U1878 (N_1878,N_1820,N_1824);
nand U1879 (N_1879,N_1858,N_1809);
nor U1880 (N_1880,N_1810,N_1829);
or U1881 (N_1881,N_1826,N_1815);
nor U1882 (N_1882,N_1852,N_1819);
and U1883 (N_1883,N_1838,N_1833);
and U1884 (N_1884,N_1861,N_1834);
and U1885 (N_1885,N_1860,N_1818);
or U1886 (N_1886,N_1847,N_1853);
or U1887 (N_1887,N_1864,N_1817);
nor U1888 (N_1888,N_1862,N_1842);
nand U1889 (N_1889,N_1843,N_1868);
nor U1890 (N_1890,N_1851,N_1831);
and U1891 (N_1891,N_1841,N_1823);
and U1892 (N_1892,N_1807,N_1863);
or U1893 (N_1893,N_1854,N_1828);
nor U1894 (N_1894,N_1857,N_1850);
and U1895 (N_1895,N_1848,N_1844);
xnor U1896 (N_1896,N_1821,N_1802);
and U1897 (N_1897,N_1811,N_1871);
or U1898 (N_1898,N_1866,N_1859);
nand U1899 (N_1899,N_1839,N_1822);
nand U1900 (N_1900,N_1845,N_1870);
nor U1901 (N_1901,N_1856,N_1805);
nor U1902 (N_1902,N_1865,N_1835);
nand U1903 (N_1903,N_1801,N_1873);
nand U1904 (N_1904,N_1855,N_1827);
or U1905 (N_1905,N_1808,N_1849);
or U1906 (N_1906,N_1806,N_1803);
nand U1907 (N_1907,N_1804,N_1814);
nor U1908 (N_1908,N_1874,N_1830);
nor U1909 (N_1909,N_1825,N_1836);
or U1910 (N_1910,N_1816,N_1837);
or U1911 (N_1911,N_1869,N_1867);
nor U1912 (N_1912,N_1813,N_1831);
nand U1913 (N_1913,N_1817,N_1856);
or U1914 (N_1914,N_1830,N_1816);
nor U1915 (N_1915,N_1859,N_1855);
nand U1916 (N_1916,N_1830,N_1815);
or U1917 (N_1917,N_1844,N_1850);
and U1918 (N_1918,N_1867,N_1855);
and U1919 (N_1919,N_1812,N_1845);
or U1920 (N_1920,N_1866,N_1870);
and U1921 (N_1921,N_1804,N_1843);
and U1922 (N_1922,N_1852,N_1826);
and U1923 (N_1923,N_1861,N_1811);
nand U1924 (N_1924,N_1804,N_1865);
or U1925 (N_1925,N_1841,N_1843);
nand U1926 (N_1926,N_1856,N_1854);
nand U1927 (N_1927,N_1839,N_1845);
nand U1928 (N_1928,N_1848,N_1863);
or U1929 (N_1929,N_1812,N_1848);
or U1930 (N_1930,N_1853,N_1806);
nand U1931 (N_1931,N_1858,N_1807);
and U1932 (N_1932,N_1801,N_1805);
and U1933 (N_1933,N_1832,N_1841);
nor U1934 (N_1934,N_1836,N_1821);
nand U1935 (N_1935,N_1864,N_1833);
or U1936 (N_1936,N_1866,N_1856);
and U1937 (N_1937,N_1813,N_1821);
or U1938 (N_1938,N_1810,N_1845);
and U1939 (N_1939,N_1813,N_1818);
or U1940 (N_1940,N_1821,N_1811);
nor U1941 (N_1941,N_1832,N_1865);
nor U1942 (N_1942,N_1836,N_1847);
or U1943 (N_1943,N_1859,N_1873);
and U1944 (N_1944,N_1863,N_1829);
and U1945 (N_1945,N_1830,N_1841);
and U1946 (N_1946,N_1821,N_1816);
and U1947 (N_1947,N_1830,N_1868);
nor U1948 (N_1948,N_1809,N_1860);
or U1949 (N_1949,N_1866,N_1862);
or U1950 (N_1950,N_1891,N_1895);
xnor U1951 (N_1951,N_1920,N_1905);
xor U1952 (N_1952,N_1927,N_1907);
and U1953 (N_1953,N_1933,N_1910);
nand U1954 (N_1954,N_1942,N_1939);
nand U1955 (N_1955,N_1893,N_1894);
and U1956 (N_1956,N_1930,N_1946);
nand U1957 (N_1957,N_1881,N_1949);
or U1958 (N_1958,N_1898,N_1931);
or U1959 (N_1959,N_1885,N_1892);
xor U1960 (N_1960,N_1896,N_1897);
nor U1961 (N_1961,N_1938,N_1882);
and U1962 (N_1962,N_1913,N_1944);
and U1963 (N_1963,N_1909,N_1904);
nand U1964 (N_1964,N_1875,N_1878);
or U1965 (N_1965,N_1932,N_1923);
nor U1966 (N_1966,N_1888,N_1890);
or U1967 (N_1967,N_1906,N_1914);
nand U1968 (N_1968,N_1948,N_1917);
nand U1969 (N_1969,N_1916,N_1876);
or U1970 (N_1970,N_1884,N_1908);
nand U1971 (N_1971,N_1937,N_1945);
and U1972 (N_1972,N_1936,N_1940);
or U1973 (N_1973,N_1887,N_1929);
nand U1974 (N_1974,N_1919,N_1934);
nor U1975 (N_1975,N_1899,N_1925);
nand U1976 (N_1976,N_1912,N_1924);
or U1977 (N_1977,N_1903,N_1886);
nor U1978 (N_1978,N_1880,N_1928);
nor U1979 (N_1979,N_1900,N_1935);
nor U1980 (N_1980,N_1915,N_1947);
nor U1981 (N_1981,N_1911,N_1902);
and U1982 (N_1982,N_1889,N_1918);
and U1983 (N_1983,N_1877,N_1922);
nand U1984 (N_1984,N_1883,N_1926);
nor U1985 (N_1985,N_1921,N_1879);
nand U1986 (N_1986,N_1901,N_1943);
nor U1987 (N_1987,N_1941,N_1911);
or U1988 (N_1988,N_1880,N_1878);
nand U1989 (N_1989,N_1919,N_1902);
nand U1990 (N_1990,N_1884,N_1917);
and U1991 (N_1991,N_1945,N_1915);
and U1992 (N_1992,N_1885,N_1949);
and U1993 (N_1993,N_1900,N_1949);
nand U1994 (N_1994,N_1899,N_1927);
nand U1995 (N_1995,N_1933,N_1944);
nand U1996 (N_1996,N_1905,N_1908);
or U1997 (N_1997,N_1911,N_1883);
nor U1998 (N_1998,N_1911,N_1938);
or U1999 (N_1999,N_1928,N_1901);
xnor U2000 (N_2000,N_1939,N_1947);
nor U2001 (N_2001,N_1912,N_1892);
or U2002 (N_2002,N_1941,N_1940);
nand U2003 (N_2003,N_1927,N_1928);
nand U2004 (N_2004,N_1943,N_1924);
nand U2005 (N_2005,N_1916,N_1918);
and U2006 (N_2006,N_1949,N_1907);
nor U2007 (N_2007,N_1930,N_1938);
or U2008 (N_2008,N_1938,N_1942);
nand U2009 (N_2009,N_1892,N_1889);
nand U2010 (N_2010,N_1901,N_1932);
or U2011 (N_2011,N_1931,N_1889);
or U2012 (N_2012,N_1914,N_1947);
nor U2013 (N_2013,N_1938,N_1885);
or U2014 (N_2014,N_1929,N_1888);
and U2015 (N_2015,N_1896,N_1933);
or U2016 (N_2016,N_1886,N_1893);
nor U2017 (N_2017,N_1944,N_1937);
or U2018 (N_2018,N_1881,N_1941);
and U2019 (N_2019,N_1907,N_1877);
and U2020 (N_2020,N_1929,N_1900);
nand U2021 (N_2021,N_1889,N_1934);
nor U2022 (N_2022,N_1889,N_1899);
xnor U2023 (N_2023,N_1931,N_1878);
or U2024 (N_2024,N_1912,N_1881);
nand U2025 (N_2025,N_1997,N_1960);
and U2026 (N_2026,N_1981,N_2000);
and U2027 (N_2027,N_1950,N_1992);
nand U2028 (N_2028,N_1959,N_2012);
and U2029 (N_2029,N_1993,N_1968);
and U2030 (N_2030,N_1985,N_1972);
nor U2031 (N_2031,N_1988,N_1980);
or U2032 (N_2032,N_1984,N_2004);
nor U2033 (N_2033,N_1991,N_1983);
nor U2034 (N_2034,N_2020,N_2007);
nand U2035 (N_2035,N_1971,N_1996);
nand U2036 (N_2036,N_1973,N_2014);
and U2037 (N_2037,N_2002,N_2003);
nor U2038 (N_2038,N_1975,N_1974);
nor U2039 (N_2039,N_2015,N_1990);
xor U2040 (N_2040,N_1986,N_1955);
and U2041 (N_2041,N_1958,N_2018);
nand U2042 (N_2042,N_2011,N_2022);
nor U2043 (N_2043,N_2021,N_1977);
nand U2044 (N_2044,N_1994,N_2019);
and U2045 (N_2045,N_1952,N_1970);
nand U2046 (N_2046,N_2009,N_1976);
or U2047 (N_2047,N_1962,N_1989);
nand U2048 (N_2048,N_2005,N_1967);
and U2049 (N_2049,N_2016,N_2024);
nand U2050 (N_2050,N_1969,N_1965);
nand U2051 (N_2051,N_1966,N_2017);
and U2052 (N_2052,N_1954,N_1995);
or U2053 (N_2053,N_1978,N_1964);
nor U2054 (N_2054,N_2013,N_1956);
xnor U2055 (N_2055,N_1999,N_2023);
or U2056 (N_2056,N_1961,N_1979);
nor U2057 (N_2057,N_2008,N_1957);
or U2058 (N_2058,N_1987,N_2006);
nor U2059 (N_2059,N_1951,N_1963);
nand U2060 (N_2060,N_1982,N_1998);
and U2061 (N_2061,N_1953,N_2001);
nand U2062 (N_2062,N_2010,N_1957);
and U2063 (N_2063,N_1992,N_2001);
nor U2064 (N_2064,N_2011,N_2015);
or U2065 (N_2065,N_2003,N_2009);
nor U2066 (N_2066,N_1980,N_2018);
nor U2067 (N_2067,N_1994,N_1989);
nor U2068 (N_2068,N_1969,N_2023);
nand U2069 (N_2069,N_1961,N_2021);
nand U2070 (N_2070,N_1988,N_1974);
and U2071 (N_2071,N_1974,N_2020);
nand U2072 (N_2072,N_1975,N_1951);
nand U2073 (N_2073,N_2005,N_2004);
or U2074 (N_2074,N_1991,N_1998);
and U2075 (N_2075,N_2024,N_1993);
nor U2076 (N_2076,N_2016,N_2014);
nand U2077 (N_2077,N_2023,N_1967);
xor U2078 (N_2078,N_1968,N_1950);
nand U2079 (N_2079,N_1965,N_1954);
xor U2080 (N_2080,N_2018,N_1963);
and U2081 (N_2081,N_1987,N_2010);
nand U2082 (N_2082,N_2003,N_2022);
nand U2083 (N_2083,N_1964,N_1963);
and U2084 (N_2084,N_1989,N_2002);
and U2085 (N_2085,N_1994,N_1984);
nand U2086 (N_2086,N_2007,N_1984);
nand U2087 (N_2087,N_1995,N_2003);
nand U2088 (N_2088,N_1970,N_1967);
and U2089 (N_2089,N_1951,N_2012);
or U2090 (N_2090,N_1962,N_1963);
or U2091 (N_2091,N_2004,N_1971);
xnor U2092 (N_2092,N_2023,N_1972);
nand U2093 (N_2093,N_2005,N_1991);
and U2094 (N_2094,N_2015,N_2023);
or U2095 (N_2095,N_1983,N_1958);
or U2096 (N_2096,N_2024,N_1953);
or U2097 (N_2097,N_1972,N_2008);
or U2098 (N_2098,N_1993,N_1997);
or U2099 (N_2099,N_2014,N_1952);
nand U2100 (N_2100,N_2086,N_2069);
nand U2101 (N_2101,N_2052,N_2081);
xor U2102 (N_2102,N_2058,N_2068);
nand U2103 (N_2103,N_2082,N_2046);
or U2104 (N_2104,N_2077,N_2094);
and U2105 (N_2105,N_2080,N_2053);
and U2106 (N_2106,N_2089,N_2073);
or U2107 (N_2107,N_2097,N_2064);
nor U2108 (N_2108,N_2049,N_2091);
nor U2109 (N_2109,N_2026,N_2029);
nor U2110 (N_2110,N_2027,N_2095);
nand U2111 (N_2111,N_2036,N_2066);
or U2112 (N_2112,N_2040,N_2051);
nor U2113 (N_2113,N_2079,N_2044);
or U2114 (N_2114,N_2060,N_2035);
or U2115 (N_2115,N_2057,N_2047);
and U2116 (N_2116,N_2045,N_2038);
or U2117 (N_2117,N_2032,N_2092);
nor U2118 (N_2118,N_2050,N_2070);
nor U2119 (N_2119,N_2088,N_2071);
and U2120 (N_2120,N_2063,N_2076);
or U2121 (N_2121,N_2034,N_2030);
or U2122 (N_2122,N_2098,N_2061);
nor U2123 (N_2123,N_2025,N_2037);
and U2124 (N_2124,N_2093,N_2072);
and U2125 (N_2125,N_2084,N_2056);
nor U2126 (N_2126,N_2078,N_2083);
or U2127 (N_2127,N_2033,N_2067);
nand U2128 (N_2128,N_2048,N_2065);
nor U2129 (N_2129,N_2042,N_2087);
or U2130 (N_2130,N_2075,N_2041);
and U2131 (N_2131,N_2059,N_2074);
nand U2132 (N_2132,N_2031,N_2062);
or U2133 (N_2133,N_2043,N_2054);
xor U2134 (N_2134,N_2028,N_2085);
nand U2135 (N_2135,N_2096,N_2099);
and U2136 (N_2136,N_2039,N_2055);
nand U2137 (N_2137,N_2090,N_2072);
nand U2138 (N_2138,N_2029,N_2089);
nand U2139 (N_2139,N_2032,N_2064);
and U2140 (N_2140,N_2040,N_2059);
nor U2141 (N_2141,N_2065,N_2041);
nor U2142 (N_2142,N_2084,N_2067);
nor U2143 (N_2143,N_2077,N_2095);
or U2144 (N_2144,N_2054,N_2034);
nand U2145 (N_2145,N_2064,N_2035);
nor U2146 (N_2146,N_2068,N_2071);
or U2147 (N_2147,N_2051,N_2029);
nor U2148 (N_2148,N_2081,N_2067);
and U2149 (N_2149,N_2092,N_2054);
nor U2150 (N_2150,N_2042,N_2075);
or U2151 (N_2151,N_2031,N_2073);
nand U2152 (N_2152,N_2063,N_2084);
nor U2153 (N_2153,N_2082,N_2041);
or U2154 (N_2154,N_2079,N_2052);
nor U2155 (N_2155,N_2098,N_2068);
and U2156 (N_2156,N_2071,N_2029);
nand U2157 (N_2157,N_2044,N_2081);
and U2158 (N_2158,N_2032,N_2098);
or U2159 (N_2159,N_2085,N_2082);
and U2160 (N_2160,N_2051,N_2035);
nand U2161 (N_2161,N_2050,N_2039);
or U2162 (N_2162,N_2050,N_2035);
or U2163 (N_2163,N_2048,N_2050);
nand U2164 (N_2164,N_2057,N_2058);
or U2165 (N_2165,N_2099,N_2060);
nor U2166 (N_2166,N_2028,N_2083);
and U2167 (N_2167,N_2028,N_2081);
nor U2168 (N_2168,N_2075,N_2038);
nand U2169 (N_2169,N_2068,N_2077);
nor U2170 (N_2170,N_2072,N_2045);
nor U2171 (N_2171,N_2048,N_2074);
or U2172 (N_2172,N_2071,N_2030);
nor U2173 (N_2173,N_2079,N_2099);
xnor U2174 (N_2174,N_2052,N_2041);
nand U2175 (N_2175,N_2106,N_2128);
and U2176 (N_2176,N_2133,N_2164);
xnor U2177 (N_2177,N_2155,N_2158);
nor U2178 (N_2178,N_2139,N_2147);
nand U2179 (N_2179,N_2118,N_2142);
nand U2180 (N_2180,N_2145,N_2125);
and U2181 (N_2181,N_2104,N_2110);
and U2182 (N_2182,N_2144,N_2132);
nand U2183 (N_2183,N_2103,N_2109);
nand U2184 (N_2184,N_2134,N_2169);
nand U2185 (N_2185,N_2166,N_2167);
nand U2186 (N_2186,N_2141,N_2162);
and U2187 (N_2187,N_2138,N_2159);
nor U2188 (N_2188,N_2126,N_2105);
nand U2189 (N_2189,N_2160,N_2116);
and U2190 (N_2190,N_2115,N_2113);
and U2191 (N_2191,N_2165,N_2168);
or U2192 (N_2192,N_2170,N_2120);
nand U2193 (N_2193,N_2173,N_2102);
or U2194 (N_2194,N_2117,N_2148);
and U2195 (N_2195,N_2111,N_2136);
and U2196 (N_2196,N_2174,N_2131);
nor U2197 (N_2197,N_2108,N_2123);
or U2198 (N_2198,N_2156,N_2121);
or U2199 (N_2199,N_2154,N_2161);
nor U2200 (N_2200,N_2127,N_2112);
xor U2201 (N_2201,N_2119,N_2163);
nor U2202 (N_2202,N_2124,N_2157);
or U2203 (N_2203,N_2171,N_2149);
or U2204 (N_2204,N_2143,N_2101);
xor U2205 (N_2205,N_2107,N_2130);
and U2206 (N_2206,N_2129,N_2152);
nor U2207 (N_2207,N_2153,N_2122);
and U2208 (N_2208,N_2172,N_2114);
or U2209 (N_2209,N_2146,N_2150);
nand U2210 (N_2210,N_2137,N_2135);
nand U2211 (N_2211,N_2140,N_2151);
nand U2212 (N_2212,N_2100,N_2138);
or U2213 (N_2213,N_2127,N_2140);
nand U2214 (N_2214,N_2144,N_2135);
and U2215 (N_2215,N_2157,N_2174);
or U2216 (N_2216,N_2140,N_2149);
xor U2217 (N_2217,N_2150,N_2129);
and U2218 (N_2218,N_2144,N_2119);
nor U2219 (N_2219,N_2148,N_2102);
or U2220 (N_2220,N_2137,N_2102);
or U2221 (N_2221,N_2128,N_2119);
and U2222 (N_2222,N_2111,N_2158);
nand U2223 (N_2223,N_2114,N_2159);
nor U2224 (N_2224,N_2156,N_2138);
and U2225 (N_2225,N_2151,N_2172);
or U2226 (N_2226,N_2142,N_2148);
or U2227 (N_2227,N_2127,N_2132);
nor U2228 (N_2228,N_2127,N_2152);
nor U2229 (N_2229,N_2118,N_2140);
and U2230 (N_2230,N_2149,N_2147);
nor U2231 (N_2231,N_2127,N_2158);
nor U2232 (N_2232,N_2119,N_2166);
nor U2233 (N_2233,N_2113,N_2162);
nor U2234 (N_2234,N_2117,N_2155);
nor U2235 (N_2235,N_2118,N_2174);
nand U2236 (N_2236,N_2113,N_2114);
or U2237 (N_2237,N_2174,N_2112);
nand U2238 (N_2238,N_2162,N_2159);
nor U2239 (N_2239,N_2123,N_2154);
or U2240 (N_2240,N_2150,N_2157);
nor U2241 (N_2241,N_2106,N_2130);
nor U2242 (N_2242,N_2125,N_2163);
nor U2243 (N_2243,N_2106,N_2113);
or U2244 (N_2244,N_2127,N_2170);
and U2245 (N_2245,N_2103,N_2115);
and U2246 (N_2246,N_2169,N_2160);
nor U2247 (N_2247,N_2104,N_2145);
and U2248 (N_2248,N_2153,N_2149);
xor U2249 (N_2249,N_2121,N_2116);
nand U2250 (N_2250,N_2202,N_2233);
nand U2251 (N_2251,N_2226,N_2221);
or U2252 (N_2252,N_2175,N_2198);
nand U2253 (N_2253,N_2245,N_2178);
nor U2254 (N_2254,N_2200,N_2186);
and U2255 (N_2255,N_2177,N_2214);
nand U2256 (N_2256,N_2248,N_2201);
or U2257 (N_2257,N_2238,N_2210);
or U2258 (N_2258,N_2208,N_2219);
or U2259 (N_2259,N_2244,N_2211);
nor U2260 (N_2260,N_2249,N_2217);
nor U2261 (N_2261,N_2187,N_2232);
and U2262 (N_2262,N_2176,N_2213);
nor U2263 (N_2263,N_2229,N_2216);
nor U2264 (N_2264,N_2239,N_2240);
or U2265 (N_2265,N_2247,N_2193);
or U2266 (N_2266,N_2246,N_2218);
or U2267 (N_2267,N_2206,N_2224);
nor U2268 (N_2268,N_2196,N_2197);
and U2269 (N_2269,N_2209,N_2227);
nand U2270 (N_2270,N_2185,N_2234);
nand U2271 (N_2271,N_2228,N_2236);
or U2272 (N_2272,N_2192,N_2243);
nand U2273 (N_2273,N_2179,N_2241);
nor U2274 (N_2274,N_2182,N_2199);
nand U2275 (N_2275,N_2204,N_2223);
nor U2276 (N_2276,N_2195,N_2189);
xor U2277 (N_2277,N_2203,N_2181);
nor U2278 (N_2278,N_2205,N_2207);
nor U2279 (N_2279,N_2191,N_2190);
nand U2280 (N_2280,N_2184,N_2235);
or U2281 (N_2281,N_2230,N_2225);
nor U2282 (N_2282,N_2188,N_2215);
and U2283 (N_2283,N_2222,N_2183);
nand U2284 (N_2284,N_2180,N_2220);
or U2285 (N_2285,N_2194,N_2242);
nand U2286 (N_2286,N_2212,N_2231);
nor U2287 (N_2287,N_2237,N_2202);
nand U2288 (N_2288,N_2219,N_2235);
nor U2289 (N_2289,N_2229,N_2188);
or U2290 (N_2290,N_2225,N_2238);
nor U2291 (N_2291,N_2221,N_2213);
and U2292 (N_2292,N_2214,N_2243);
and U2293 (N_2293,N_2227,N_2218);
nand U2294 (N_2294,N_2184,N_2236);
and U2295 (N_2295,N_2222,N_2205);
and U2296 (N_2296,N_2226,N_2225);
nand U2297 (N_2297,N_2218,N_2223);
nor U2298 (N_2298,N_2191,N_2230);
and U2299 (N_2299,N_2246,N_2234);
or U2300 (N_2300,N_2234,N_2179);
or U2301 (N_2301,N_2202,N_2221);
nand U2302 (N_2302,N_2222,N_2234);
and U2303 (N_2303,N_2199,N_2241);
nor U2304 (N_2304,N_2183,N_2229);
nand U2305 (N_2305,N_2215,N_2183);
nor U2306 (N_2306,N_2182,N_2230);
and U2307 (N_2307,N_2213,N_2231);
nand U2308 (N_2308,N_2233,N_2243);
xnor U2309 (N_2309,N_2248,N_2225);
nor U2310 (N_2310,N_2177,N_2236);
nor U2311 (N_2311,N_2213,N_2190);
nor U2312 (N_2312,N_2225,N_2243);
or U2313 (N_2313,N_2215,N_2206);
or U2314 (N_2314,N_2239,N_2229);
or U2315 (N_2315,N_2188,N_2218);
or U2316 (N_2316,N_2201,N_2176);
nand U2317 (N_2317,N_2229,N_2221);
and U2318 (N_2318,N_2225,N_2183);
or U2319 (N_2319,N_2178,N_2222);
or U2320 (N_2320,N_2203,N_2233);
nor U2321 (N_2321,N_2228,N_2195);
nor U2322 (N_2322,N_2204,N_2217);
nor U2323 (N_2323,N_2227,N_2226);
or U2324 (N_2324,N_2212,N_2177);
nor U2325 (N_2325,N_2253,N_2314);
or U2326 (N_2326,N_2309,N_2278);
nand U2327 (N_2327,N_2298,N_2305);
or U2328 (N_2328,N_2271,N_2311);
or U2329 (N_2329,N_2291,N_2324);
nor U2330 (N_2330,N_2269,N_2267);
or U2331 (N_2331,N_2276,N_2260);
nor U2332 (N_2332,N_2286,N_2300);
nand U2333 (N_2333,N_2255,N_2258);
and U2334 (N_2334,N_2262,N_2323);
nand U2335 (N_2335,N_2275,N_2293);
or U2336 (N_2336,N_2273,N_2304);
nand U2337 (N_2337,N_2279,N_2320);
or U2338 (N_2338,N_2312,N_2302);
and U2339 (N_2339,N_2261,N_2259);
or U2340 (N_2340,N_2321,N_2288);
or U2341 (N_2341,N_2296,N_2250);
nor U2342 (N_2342,N_2294,N_2257);
or U2343 (N_2343,N_2297,N_2301);
or U2344 (N_2344,N_2254,N_2285);
nor U2345 (N_2345,N_2256,N_2251);
or U2346 (N_2346,N_2313,N_2307);
and U2347 (N_2347,N_2284,N_2299);
and U2348 (N_2348,N_2252,N_2306);
xor U2349 (N_2349,N_2289,N_2264);
nand U2350 (N_2350,N_2274,N_2317);
or U2351 (N_2351,N_2281,N_2292);
or U2352 (N_2352,N_2282,N_2283);
or U2353 (N_2353,N_2265,N_2316);
and U2354 (N_2354,N_2268,N_2308);
and U2355 (N_2355,N_2290,N_2322);
and U2356 (N_2356,N_2287,N_2272);
and U2357 (N_2357,N_2270,N_2263);
nor U2358 (N_2358,N_2280,N_2315);
or U2359 (N_2359,N_2310,N_2318);
nand U2360 (N_2360,N_2266,N_2295);
or U2361 (N_2361,N_2303,N_2319);
or U2362 (N_2362,N_2277,N_2302);
nor U2363 (N_2363,N_2324,N_2269);
and U2364 (N_2364,N_2318,N_2257);
and U2365 (N_2365,N_2308,N_2309);
nand U2366 (N_2366,N_2262,N_2293);
or U2367 (N_2367,N_2302,N_2282);
nand U2368 (N_2368,N_2291,N_2282);
nor U2369 (N_2369,N_2287,N_2288);
nor U2370 (N_2370,N_2266,N_2306);
and U2371 (N_2371,N_2313,N_2255);
nand U2372 (N_2372,N_2264,N_2302);
or U2373 (N_2373,N_2269,N_2283);
and U2374 (N_2374,N_2298,N_2290);
nor U2375 (N_2375,N_2291,N_2310);
nor U2376 (N_2376,N_2282,N_2285);
nor U2377 (N_2377,N_2273,N_2269);
or U2378 (N_2378,N_2281,N_2258);
or U2379 (N_2379,N_2287,N_2258);
or U2380 (N_2380,N_2290,N_2268);
nor U2381 (N_2381,N_2273,N_2266);
nor U2382 (N_2382,N_2303,N_2271);
nand U2383 (N_2383,N_2293,N_2297);
nor U2384 (N_2384,N_2282,N_2294);
nor U2385 (N_2385,N_2293,N_2283);
xnor U2386 (N_2386,N_2269,N_2256);
or U2387 (N_2387,N_2257,N_2261);
or U2388 (N_2388,N_2259,N_2307);
or U2389 (N_2389,N_2285,N_2320);
xor U2390 (N_2390,N_2305,N_2292);
or U2391 (N_2391,N_2251,N_2309);
or U2392 (N_2392,N_2251,N_2260);
nand U2393 (N_2393,N_2272,N_2250);
or U2394 (N_2394,N_2297,N_2272);
and U2395 (N_2395,N_2290,N_2279);
nand U2396 (N_2396,N_2298,N_2302);
and U2397 (N_2397,N_2253,N_2322);
nand U2398 (N_2398,N_2305,N_2271);
and U2399 (N_2399,N_2299,N_2287);
and U2400 (N_2400,N_2340,N_2387);
or U2401 (N_2401,N_2365,N_2385);
or U2402 (N_2402,N_2397,N_2335);
or U2403 (N_2403,N_2368,N_2329);
nor U2404 (N_2404,N_2352,N_2366);
or U2405 (N_2405,N_2356,N_2393);
nor U2406 (N_2406,N_2388,N_2334);
nor U2407 (N_2407,N_2326,N_2371);
and U2408 (N_2408,N_2394,N_2351);
nor U2409 (N_2409,N_2337,N_2342);
nor U2410 (N_2410,N_2369,N_2373);
and U2411 (N_2411,N_2354,N_2399);
nand U2412 (N_2412,N_2346,N_2330);
nand U2413 (N_2413,N_2355,N_2395);
nand U2414 (N_2414,N_2375,N_2348);
or U2415 (N_2415,N_2325,N_2353);
or U2416 (N_2416,N_2398,N_2377);
and U2417 (N_2417,N_2396,N_2391);
nor U2418 (N_2418,N_2359,N_2343);
nand U2419 (N_2419,N_2327,N_2347);
nand U2420 (N_2420,N_2363,N_2382);
and U2421 (N_2421,N_2390,N_2332);
or U2422 (N_2422,N_2380,N_2389);
or U2423 (N_2423,N_2386,N_2338);
and U2424 (N_2424,N_2372,N_2379);
nor U2425 (N_2425,N_2378,N_2336);
nor U2426 (N_2426,N_2357,N_2344);
nor U2427 (N_2427,N_2367,N_2349);
or U2428 (N_2428,N_2345,N_2361);
and U2429 (N_2429,N_2374,N_2384);
or U2430 (N_2430,N_2333,N_2350);
nor U2431 (N_2431,N_2392,N_2362);
nand U2432 (N_2432,N_2381,N_2360);
or U2433 (N_2433,N_2341,N_2339);
or U2434 (N_2434,N_2370,N_2364);
and U2435 (N_2435,N_2328,N_2358);
nand U2436 (N_2436,N_2331,N_2376);
nor U2437 (N_2437,N_2383,N_2361);
nand U2438 (N_2438,N_2355,N_2357);
nand U2439 (N_2439,N_2327,N_2336);
nor U2440 (N_2440,N_2388,N_2375);
or U2441 (N_2441,N_2368,N_2344);
nor U2442 (N_2442,N_2342,N_2357);
or U2443 (N_2443,N_2360,N_2327);
nand U2444 (N_2444,N_2366,N_2374);
or U2445 (N_2445,N_2329,N_2389);
xnor U2446 (N_2446,N_2386,N_2356);
nand U2447 (N_2447,N_2379,N_2385);
or U2448 (N_2448,N_2330,N_2359);
and U2449 (N_2449,N_2378,N_2380);
and U2450 (N_2450,N_2360,N_2343);
nand U2451 (N_2451,N_2375,N_2330);
xnor U2452 (N_2452,N_2325,N_2381);
and U2453 (N_2453,N_2385,N_2383);
or U2454 (N_2454,N_2395,N_2331);
nor U2455 (N_2455,N_2389,N_2352);
or U2456 (N_2456,N_2382,N_2331);
nor U2457 (N_2457,N_2367,N_2370);
or U2458 (N_2458,N_2349,N_2381);
or U2459 (N_2459,N_2331,N_2354);
or U2460 (N_2460,N_2371,N_2359);
or U2461 (N_2461,N_2351,N_2382);
or U2462 (N_2462,N_2349,N_2391);
and U2463 (N_2463,N_2352,N_2348);
nand U2464 (N_2464,N_2375,N_2340);
and U2465 (N_2465,N_2389,N_2351);
nand U2466 (N_2466,N_2349,N_2355);
nand U2467 (N_2467,N_2364,N_2332);
nor U2468 (N_2468,N_2386,N_2343);
and U2469 (N_2469,N_2326,N_2379);
and U2470 (N_2470,N_2393,N_2378);
or U2471 (N_2471,N_2395,N_2327);
and U2472 (N_2472,N_2327,N_2380);
or U2473 (N_2473,N_2333,N_2362);
and U2474 (N_2474,N_2387,N_2389);
nand U2475 (N_2475,N_2420,N_2422);
and U2476 (N_2476,N_2457,N_2416);
nand U2477 (N_2477,N_2469,N_2406);
or U2478 (N_2478,N_2456,N_2411);
and U2479 (N_2479,N_2435,N_2419);
or U2480 (N_2480,N_2401,N_2462);
nand U2481 (N_2481,N_2428,N_2461);
and U2482 (N_2482,N_2447,N_2421);
and U2483 (N_2483,N_2466,N_2424);
nor U2484 (N_2484,N_2454,N_2407);
nor U2485 (N_2485,N_2467,N_2434);
xnor U2486 (N_2486,N_2470,N_2444);
or U2487 (N_2487,N_2452,N_2468);
nor U2488 (N_2488,N_2464,N_2438);
nand U2489 (N_2489,N_2433,N_2413);
or U2490 (N_2490,N_2414,N_2437);
xor U2491 (N_2491,N_2460,N_2451);
nand U2492 (N_2492,N_2427,N_2429);
and U2493 (N_2493,N_2408,N_2440);
and U2494 (N_2494,N_2453,N_2425);
and U2495 (N_2495,N_2432,N_2410);
and U2496 (N_2496,N_2403,N_2436);
and U2497 (N_2497,N_2426,N_2463);
nand U2498 (N_2498,N_2404,N_2465);
or U2499 (N_2499,N_2455,N_2448);
and U2500 (N_2500,N_2459,N_2439);
nor U2501 (N_2501,N_2450,N_2402);
or U2502 (N_2502,N_2442,N_2417);
nor U2503 (N_2503,N_2423,N_2445);
or U2504 (N_2504,N_2471,N_2441);
nor U2505 (N_2505,N_2415,N_2443);
xnor U2506 (N_2506,N_2430,N_2412);
nor U2507 (N_2507,N_2431,N_2449);
nor U2508 (N_2508,N_2472,N_2458);
or U2509 (N_2509,N_2446,N_2418);
or U2510 (N_2510,N_2473,N_2400);
or U2511 (N_2511,N_2409,N_2474);
or U2512 (N_2512,N_2405,N_2427);
or U2513 (N_2513,N_2418,N_2448);
nand U2514 (N_2514,N_2412,N_2448);
and U2515 (N_2515,N_2470,N_2474);
nand U2516 (N_2516,N_2452,N_2451);
nand U2517 (N_2517,N_2419,N_2420);
nor U2518 (N_2518,N_2437,N_2425);
and U2519 (N_2519,N_2413,N_2432);
nor U2520 (N_2520,N_2430,N_2466);
nor U2521 (N_2521,N_2455,N_2457);
nor U2522 (N_2522,N_2473,N_2411);
nor U2523 (N_2523,N_2458,N_2428);
or U2524 (N_2524,N_2429,N_2433);
nand U2525 (N_2525,N_2428,N_2442);
and U2526 (N_2526,N_2407,N_2411);
nor U2527 (N_2527,N_2470,N_2429);
and U2528 (N_2528,N_2413,N_2431);
and U2529 (N_2529,N_2454,N_2432);
or U2530 (N_2530,N_2442,N_2420);
and U2531 (N_2531,N_2447,N_2461);
and U2532 (N_2532,N_2458,N_2423);
or U2533 (N_2533,N_2418,N_2467);
nand U2534 (N_2534,N_2460,N_2462);
nor U2535 (N_2535,N_2401,N_2402);
or U2536 (N_2536,N_2439,N_2464);
or U2537 (N_2537,N_2440,N_2442);
or U2538 (N_2538,N_2457,N_2431);
xor U2539 (N_2539,N_2410,N_2422);
or U2540 (N_2540,N_2471,N_2464);
nand U2541 (N_2541,N_2431,N_2432);
nor U2542 (N_2542,N_2452,N_2448);
or U2543 (N_2543,N_2452,N_2402);
nor U2544 (N_2544,N_2474,N_2442);
and U2545 (N_2545,N_2413,N_2468);
nand U2546 (N_2546,N_2414,N_2461);
and U2547 (N_2547,N_2456,N_2459);
nor U2548 (N_2548,N_2405,N_2441);
nand U2549 (N_2549,N_2443,N_2421);
nand U2550 (N_2550,N_2518,N_2513);
nor U2551 (N_2551,N_2542,N_2484);
and U2552 (N_2552,N_2549,N_2547);
or U2553 (N_2553,N_2529,N_2536);
nand U2554 (N_2554,N_2510,N_2487);
or U2555 (N_2555,N_2535,N_2506);
nor U2556 (N_2556,N_2543,N_2530);
nand U2557 (N_2557,N_2541,N_2523);
nand U2558 (N_2558,N_2546,N_2525);
nand U2559 (N_2559,N_2532,N_2476);
or U2560 (N_2560,N_2515,N_2478);
and U2561 (N_2561,N_2534,N_2501);
nand U2562 (N_2562,N_2526,N_2498);
or U2563 (N_2563,N_2544,N_2519);
nor U2564 (N_2564,N_2521,N_2516);
nor U2565 (N_2565,N_2517,N_2482);
nand U2566 (N_2566,N_2499,N_2486);
and U2567 (N_2567,N_2514,N_2496);
and U2568 (N_2568,N_2485,N_2548);
or U2569 (N_2569,N_2537,N_2492);
and U2570 (N_2570,N_2512,N_2495);
nand U2571 (N_2571,N_2511,N_2493);
and U2572 (N_2572,N_2539,N_2540);
nand U2573 (N_2573,N_2507,N_2483);
or U2574 (N_2574,N_2502,N_2527);
and U2575 (N_2575,N_2538,N_2488);
and U2576 (N_2576,N_2508,N_2531);
or U2577 (N_2577,N_2533,N_2494);
or U2578 (N_2578,N_2505,N_2522);
and U2579 (N_2579,N_2528,N_2497);
or U2580 (N_2580,N_2520,N_2500);
and U2581 (N_2581,N_2503,N_2524);
nor U2582 (N_2582,N_2491,N_2490);
nor U2583 (N_2583,N_2509,N_2479);
or U2584 (N_2584,N_2504,N_2545);
and U2585 (N_2585,N_2480,N_2477);
and U2586 (N_2586,N_2489,N_2475);
xor U2587 (N_2587,N_2481,N_2506);
or U2588 (N_2588,N_2546,N_2485);
and U2589 (N_2589,N_2539,N_2520);
or U2590 (N_2590,N_2504,N_2525);
nand U2591 (N_2591,N_2487,N_2538);
or U2592 (N_2592,N_2503,N_2493);
and U2593 (N_2593,N_2529,N_2531);
or U2594 (N_2594,N_2514,N_2520);
and U2595 (N_2595,N_2484,N_2515);
or U2596 (N_2596,N_2488,N_2491);
nor U2597 (N_2597,N_2541,N_2549);
nand U2598 (N_2598,N_2518,N_2525);
nor U2599 (N_2599,N_2518,N_2533);
and U2600 (N_2600,N_2483,N_2479);
or U2601 (N_2601,N_2541,N_2533);
nand U2602 (N_2602,N_2524,N_2488);
nand U2603 (N_2603,N_2497,N_2494);
or U2604 (N_2604,N_2513,N_2494);
xor U2605 (N_2605,N_2506,N_2487);
nand U2606 (N_2606,N_2513,N_2479);
nor U2607 (N_2607,N_2487,N_2523);
nor U2608 (N_2608,N_2519,N_2478);
or U2609 (N_2609,N_2526,N_2530);
nand U2610 (N_2610,N_2489,N_2548);
nand U2611 (N_2611,N_2526,N_2537);
nor U2612 (N_2612,N_2525,N_2494);
or U2613 (N_2613,N_2507,N_2532);
nand U2614 (N_2614,N_2527,N_2482);
nor U2615 (N_2615,N_2489,N_2549);
nor U2616 (N_2616,N_2524,N_2509);
nand U2617 (N_2617,N_2507,N_2544);
and U2618 (N_2618,N_2494,N_2534);
or U2619 (N_2619,N_2543,N_2534);
nand U2620 (N_2620,N_2498,N_2536);
or U2621 (N_2621,N_2535,N_2486);
nand U2622 (N_2622,N_2509,N_2496);
and U2623 (N_2623,N_2501,N_2483);
nand U2624 (N_2624,N_2478,N_2526);
and U2625 (N_2625,N_2596,N_2577);
nand U2626 (N_2626,N_2556,N_2567);
nand U2627 (N_2627,N_2586,N_2589);
or U2628 (N_2628,N_2561,N_2624);
or U2629 (N_2629,N_2610,N_2566);
xor U2630 (N_2630,N_2550,N_2563);
nand U2631 (N_2631,N_2609,N_2614);
nor U2632 (N_2632,N_2574,N_2606);
nand U2633 (N_2633,N_2553,N_2617);
or U2634 (N_2634,N_2592,N_2555);
and U2635 (N_2635,N_2581,N_2579);
or U2636 (N_2636,N_2607,N_2557);
and U2637 (N_2637,N_2583,N_2554);
or U2638 (N_2638,N_2562,N_2582);
nand U2639 (N_2639,N_2573,N_2570);
nor U2640 (N_2640,N_2585,N_2552);
and U2641 (N_2641,N_2602,N_2580);
and U2642 (N_2642,N_2564,N_2595);
or U2643 (N_2643,N_2611,N_2588);
and U2644 (N_2644,N_2623,N_2559);
nand U2645 (N_2645,N_2615,N_2622);
nor U2646 (N_2646,N_2608,N_2598);
and U2647 (N_2647,N_2601,N_2578);
nand U2648 (N_2648,N_2603,N_2571);
or U2649 (N_2649,N_2600,N_2558);
or U2650 (N_2650,N_2551,N_2576);
or U2651 (N_2651,N_2597,N_2594);
or U2652 (N_2652,N_2591,N_2618);
nor U2653 (N_2653,N_2612,N_2621);
nand U2654 (N_2654,N_2568,N_2605);
nor U2655 (N_2655,N_2569,N_2575);
and U2656 (N_2656,N_2590,N_2584);
nand U2657 (N_2657,N_2619,N_2572);
or U2658 (N_2658,N_2620,N_2613);
nand U2659 (N_2659,N_2565,N_2599);
and U2660 (N_2660,N_2593,N_2587);
nand U2661 (N_2661,N_2616,N_2604);
nand U2662 (N_2662,N_2560,N_2617);
nand U2663 (N_2663,N_2561,N_2592);
or U2664 (N_2664,N_2566,N_2614);
nand U2665 (N_2665,N_2616,N_2582);
nor U2666 (N_2666,N_2624,N_2614);
nor U2667 (N_2667,N_2554,N_2616);
and U2668 (N_2668,N_2561,N_2602);
nor U2669 (N_2669,N_2604,N_2565);
and U2670 (N_2670,N_2619,N_2601);
nand U2671 (N_2671,N_2553,N_2571);
nor U2672 (N_2672,N_2595,N_2571);
xor U2673 (N_2673,N_2581,N_2580);
nor U2674 (N_2674,N_2602,N_2599);
or U2675 (N_2675,N_2566,N_2605);
and U2676 (N_2676,N_2557,N_2590);
nor U2677 (N_2677,N_2583,N_2553);
nor U2678 (N_2678,N_2597,N_2564);
nor U2679 (N_2679,N_2622,N_2613);
and U2680 (N_2680,N_2613,N_2583);
and U2681 (N_2681,N_2571,N_2622);
nand U2682 (N_2682,N_2556,N_2624);
or U2683 (N_2683,N_2616,N_2611);
nor U2684 (N_2684,N_2596,N_2624);
nand U2685 (N_2685,N_2570,N_2582);
or U2686 (N_2686,N_2585,N_2554);
nor U2687 (N_2687,N_2590,N_2607);
or U2688 (N_2688,N_2574,N_2562);
nor U2689 (N_2689,N_2559,N_2554);
or U2690 (N_2690,N_2613,N_2555);
nor U2691 (N_2691,N_2606,N_2591);
and U2692 (N_2692,N_2621,N_2585);
and U2693 (N_2693,N_2582,N_2622);
and U2694 (N_2694,N_2610,N_2579);
and U2695 (N_2695,N_2605,N_2571);
nor U2696 (N_2696,N_2596,N_2560);
nor U2697 (N_2697,N_2617,N_2561);
nor U2698 (N_2698,N_2609,N_2607);
and U2699 (N_2699,N_2578,N_2598);
or U2700 (N_2700,N_2659,N_2683);
or U2701 (N_2701,N_2662,N_2640);
or U2702 (N_2702,N_2698,N_2672);
or U2703 (N_2703,N_2679,N_2685);
nor U2704 (N_2704,N_2634,N_2664);
nand U2705 (N_2705,N_2684,N_2637);
nand U2706 (N_2706,N_2674,N_2629);
or U2707 (N_2707,N_2675,N_2686);
nand U2708 (N_2708,N_2669,N_2681);
nor U2709 (N_2709,N_2668,N_2677);
and U2710 (N_2710,N_2625,N_2654);
and U2711 (N_2711,N_2648,N_2643);
or U2712 (N_2712,N_2645,N_2636);
xnor U2713 (N_2713,N_2688,N_2666);
or U2714 (N_2714,N_2670,N_2653);
nor U2715 (N_2715,N_2649,N_2631);
nand U2716 (N_2716,N_2665,N_2699);
and U2717 (N_2717,N_2661,N_2690);
and U2718 (N_2718,N_2692,N_2627);
nor U2719 (N_2719,N_2647,N_2682);
or U2720 (N_2720,N_2673,N_2656);
or U2721 (N_2721,N_2657,N_2660);
xor U2722 (N_2722,N_2635,N_2658);
or U2723 (N_2723,N_2693,N_2678);
or U2724 (N_2724,N_2644,N_2663);
or U2725 (N_2725,N_2691,N_2642);
nand U2726 (N_2726,N_2628,N_2626);
nor U2727 (N_2727,N_2687,N_2694);
xor U2728 (N_2728,N_2646,N_2676);
and U2729 (N_2729,N_2689,N_2650);
nor U2730 (N_2730,N_2633,N_2639);
or U2731 (N_2731,N_2652,N_2696);
nand U2732 (N_2732,N_2671,N_2651);
nor U2733 (N_2733,N_2638,N_2695);
xor U2734 (N_2734,N_2630,N_2680);
and U2735 (N_2735,N_2655,N_2641);
and U2736 (N_2736,N_2667,N_2632);
nor U2737 (N_2737,N_2697,N_2699);
or U2738 (N_2738,N_2671,N_2686);
nand U2739 (N_2739,N_2625,N_2674);
and U2740 (N_2740,N_2678,N_2672);
nor U2741 (N_2741,N_2646,N_2684);
and U2742 (N_2742,N_2654,N_2638);
and U2743 (N_2743,N_2626,N_2674);
and U2744 (N_2744,N_2635,N_2627);
nand U2745 (N_2745,N_2684,N_2675);
and U2746 (N_2746,N_2671,N_2668);
nor U2747 (N_2747,N_2631,N_2668);
and U2748 (N_2748,N_2635,N_2685);
and U2749 (N_2749,N_2678,N_2689);
nand U2750 (N_2750,N_2696,N_2695);
or U2751 (N_2751,N_2640,N_2672);
nor U2752 (N_2752,N_2697,N_2626);
and U2753 (N_2753,N_2638,N_2673);
and U2754 (N_2754,N_2696,N_2650);
nor U2755 (N_2755,N_2674,N_2697);
or U2756 (N_2756,N_2636,N_2689);
and U2757 (N_2757,N_2676,N_2667);
and U2758 (N_2758,N_2690,N_2649);
nand U2759 (N_2759,N_2625,N_2662);
and U2760 (N_2760,N_2689,N_2634);
or U2761 (N_2761,N_2678,N_2641);
or U2762 (N_2762,N_2630,N_2636);
nor U2763 (N_2763,N_2686,N_2660);
nor U2764 (N_2764,N_2653,N_2675);
nor U2765 (N_2765,N_2631,N_2688);
xnor U2766 (N_2766,N_2689,N_2668);
or U2767 (N_2767,N_2633,N_2636);
or U2768 (N_2768,N_2667,N_2628);
and U2769 (N_2769,N_2688,N_2683);
or U2770 (N_2770,N_2658,N_2626);
nor U2771 (N_2771,N_2696,N_2699);
or U2772 (N_2772,N_2641,N_2644);
nand U2773 (N_2773,N_2692,N_2681);
and U2774 (N_2774,N_2662,N_2644);
and U2775 (N_2775,N_2746,N_2716);
nor U2776 (N_2776,N_2739,N_2755);
nand U2777 (N_2777,N_2773,N_2742);
and U2778 (N_2778,N_2753,N_2710);
nor U2779 (N_2779,N_2747,N_2723);
nand U2780 (N_2780,N_2706,N_2766);
or U2781 (N_2781,N_2703,N_2724);
nor U2782 (N_2782,N_2727,N_2735);
xor U2783 (N_2783,N_2761,N_2700);
and U2784 (N_2784,N_2744,N_2763);
or U2785 (N_2785,N_2707,N_2725);
and U2786 (N_2786,N_2774,N_2717);
and U2787 (N_2787,N_2752,N_2756);
nand U2788 (N_2788,N_2769,N_2709);
or U2789 (N_2789,N_2748,N_2750);
nand U2790 (N_2790,N_2743,N_2764);
and U2791 (N_2791,N_2741,N_2715);
and U2792 (N_2792,N_2719,N_2713);
or U2793 (N_2793,N_2770,N_2734);
nand U2794 (N_2794,N_2765,N_2721);
and U2795 (N_2795,N_2729,N_2749);
nand U2796 (N_2796,N_2745,N_2751);
and U2797 (N_2797,N_2731,N_2771);
and U2798 (N_2798,N_2736,N_2740);
nor U2799 (N_2799,N_2726,N_2759);
nor U2800 (N_2800,N_2738,N_2762);
nor U2801 (N_2801,N_2730,N_2758);
or U2802 (N_2802,N_2702,N_2712);
xor U2803 (N_2803,N_2737,N_2701);
and U2804 (N_2804,N_2733,N_2772);
and U2805 (N_2805,N_2757,N_2718);
and U2806 (N_2806,N_2704,N_2705);
nand U2807 (N_2807,N_2722,N_2754);
or U2808 (N_2808,N_2714,N_2728);
nand U2809 (N_2809,N_2711,N_2732);
nor U2810 (N_2810,N_2708,N_2760);
and U2811 (N_2811,N_2720,N_2767);
nand U2812 (N_2812,N_2768,N_2736);
and U2813 (N_2813,N_2764,N_2701);
nor U2814 (N_2814,N_2726,N_2716);
and U2815 (N_2815,N_2709,N_2711);
nand U2816 (N_2816,N_2770,N_2767);
and U2817 (N_2817,N_2706,N_2713);
and U2818 (N_2818,N_2735,N_2770);
nand U2819 (N_2819,N_2734,N_2739);
nor U2820 (N_2820,N_2709,N_2718);
nor U2821 (N_2821,N_2757,N_2731);
and U2822 (N_2822,N_2746,N_2725);
or U2823 (N_2823,N_2738,N_2748);
nor U2824 (N_2824,N_2706,N_2717);
or U2825 (N_2825,N_2754,N_2735);
and U2826 (N_2826,N_2753,N_2730);
xor U2827 (N_2827,N_2705,N_2721);
and U2828 (N_2828,N_2770,N_2758);
nor U2829 (N_2829,N_2724,N_2745);
nor U2830 (N_2830,N_2720,N_2745);
and U2831 (N_2831,N_2745,N_2747);
xnor U2832 (N_2832,N_2705,N_2735);
or U2833 (N_2833,N_2770,N_2719);
and U2834 (N_2834,N_2749,N_2774);
or U2835 (N_2835,N_2762,N_2760);
nor U2836 (N_2836,N_2719,N_2763);
or U2837 (N_2837,N_2714,N_2756);
or U2838 (N_2838,N_2700,N_2757);
nand U2839 (N_2839,N_2770,N_2716);
nand U2840 (N_2840,N_2736,N_2767);
or U2841 (N_2841,N_2766,N_2730);
and U2842 (N_2842,N_2702,N_2720);
or U2843 (N_2843,N_2748,N_2774);
nand U2844 (N_2844,N_2738,N_2740);
and U2845 (N_2845,N_2700,N_2706);
nand U2846 (N_2846,N_2722,N_2744);
xor U2847 (N_2847,N_2774,N_2767);
and U2848 (N_2848,N_2737,N_2768);
nand U2849 (N_2849,N_2751,N_2748);
nand U2850 (N_2850,N_2823,N_2829);
or U2851 (N_2851,N_2789,N_2780);
nand U2852 (N_2852,N_2788,N_2821);
nand U2853 (N_2853,N_2822,N_2801);
nor U2854 (N_2854,N_2824,N_2844);
or U2855 (N_2855,N_2832,N_2838);
or U2856 (N_2856,N_2799,N_2777);
or U2857 (N_2857,N_2794,N_2791);
nor U2858 (N_2858,N_2835,N_2796);
and U2859 (N_2859,N_2813,N_2781);
or U2860 (N_2860,N_2782,N_2828);
and U2861 (N_2861,N_2798,N_2802);
or U2862 (N_2862,N_2783,N_2809);
nor U2863 (N_2863,N_2834,N_2836);
nand U2864 (N_2864,N_2784,N_2825);
or U2865 (N_2865,N_2778,N_2775);
nor U2866 (N_2866,N_2833,N_2814);
and U2867 (N_2867,N_2803,N_2807);
or U2868 (N_2868,N_2847,N_2805);
nor U2869 (N_2869,N_2815,N_2826);
and U2870 (N_2870,N_2830,N_2811);
nor U2871 (N_2871,N_2831,N_2842);
or U2872 (N_2872,N_2839,N_2795);
nor U2873 (N_2873,N_2792,N_2779);
and U2874 (N_2874,N_2800,N_2816);
and U2875 (N_2875,N_2797,N_2837);
or U2876 (N_2876,N_2776,N_2827);
xnor U2877 (N_2877,N_2790,N_2817);
nand U2878 (N_2878,N_2787,N_2810);
or U2879 (N_2879,N_2818,N_2849);
and U2880 (N_2880,N_2819,N_2808);
and U2881 (N_2881,N_2846,N_2841);
nand U2882 (N_2882,N_2848,N_2845);
or U2883 (N_2883,N_2804,N_2793);
and U2884 (N_2884,N_2820,N_2786);
nor U2885 (N_2885,N_2806,N_2785);
and U2886 (N_2886,N_2840,N_2843);
nor U2887 (N_2887,N_2812,N_2806);
nand U2888 (N_2888,N_2829,N_2794);
nand U2889 (N_2889,N_2817,N_2827);
nand U2890 (N_2890,N_2827,N_2835);
and U2891 (N_2891,N_2841,N_2786);
nor U2892 (N_2892,N_2787,N_2815);
nand U2893 (N_2893,N_2848,N_2777);
and U2894 (N_2894,N_2802,N_2810);
or U2895 (N_2895,N_2836,N_2808);
or U2896 (N_2896,N_2775,N_2821);
and U2897 (N_2897,N_2845,N_2815);
or U2898 (N_2898,N_2789,N_2776);
and U2899 (N_2899,N_2781,N_2831);
or U2900 (N_2900,N_2844,N_2838);
nand U2901 (N_2901,N_2837,N_2821);
nor U2902 (N_2902,N_2781,N_2788);
nor U2903 (N_2903,N_2832,N_2829);
or U2904 (N_2904,N_2845,N_2841);
nand U2905 (N_2905,N_2844,N_2839);
or U2906 (N_2906,N_2791,N_2801);
and U2907 (N_2907,N_2787,N_2827);
or U2908 (N_2908,N_2823,N_2837);
or U2909 (N_2909,N_2776,N_2799);
or U2910 (N_2910,N_2791,N_2800);
nor U2911 (N_2911,N_2782,N_2798);
or U2912 (N_2912,N_2794,N_2790);
nor U2913 (N_2913,N_2799,N_2848);
or U2914 (N_2914,N_2784,N_2830);
or U2915 (N_2915,N_2789,N_2828);
nor U2916 (N_2916,N_2786,N_2808);
nand U2917 (N_2917,N_2775,N_2779);
nor U2918 (N_2918,N_2797,N_2844);
and U2919 (N_2919,N_2837,N_2822);
nand U2920 (N_2920,N_2840,N_2832);
nor U2921 (N_2921,N_2783,N_2784);
and U2922 (N_2922,N_2831,N_2813);
nand U2923 (N_2923,N_2782,N_2826);
nand U2924 (N_2924,N_2847,N_2796);
nor U2925 (N_2925,N_2864,N_2883);
and U2926 (N_2926,N_2867,N_2871);
nand U2927 (N_2927,N_2861,N_2878);
nor U2928 (N_2928,N_2856,N_2896);
and U2929 (N_2929,N_2907,N_2885);
or U2930 (N_2930,N_2873,N_2912);
nand U2931 (N_2931,N_2905,N_2881);
nor U2932 (N_2932,N_2868,N_2852);
or U2933 (N_2933,N_2892,N_2854);
and U2934 (N_2934,N_2920,N_2863);
nand U2935 (N_2935,N_2866,N_2914);
nor U2936 (N_2936,N_2870,N_2859);
nand U2937 (N_2937,N_2886,N_2918);
and U2938 (N_2938,N_2893,N_2862);
nor U2939 (N_2939,N_2874,N_2922);
or U2940 (N_2940,N_2913,N_2904);
or U2941 (N_2941,N_2901,N_2853);
xnor U2942 (N_2942,N_2899,N_2855);
or U2943 (N_2943,N_2915,N_2875);
and U2944 (N_2944,N_2879,N_2890);
and U2945 (N_2945,N_2910,N_2860);
nor U2946 (N_2946,N_2850,N_2887);
or U2947 (N_2947,N_2916,N_2909);
and U2948 (N_2948,N_2898,N_2902);
nand U2949 (N_2949,N_2894,N_2908);
and U2950 (N_2950,N_2884,N_2891);
nand U2951 (N_2951,N_2924,N_2888);
nand U2952 (N_2952,N_2877,N_2889);
and U2953 (N_2953,N_2919,N_2921);
or U2954 (N_2954,N_2897,N_2900);
and U2955 (N_2955,N_2882,N_2923);
or U2956 (N_2956,N_2865,N_2872);
and U2957 (N_2957,N_2895,N_2869);
or U2958 (N_2958,N_2903,N_2851);
and U2959 (N_2959,N_2876,N_2858);
nor U2960 (N_2960,N_2917,N_2857);
and U2961 (N_2961,N_2911,N_2880);
nand U2962 (N_2962,N_2906,N_2894);
nand U2963 (N_2963,N_2876,N_2866);
nor U2964 (N_2964,N_2854,N_2869);
and U2965 (N_2965,N_2906,N_2889);
nor U2966 (N_2966,N_2880,N_2872);
and U2967 (N_2967,N_2856,N_2913);
nor U2968 (N_2968,N_2853,N_2855);
and U2969 (N_2969,N_2850,N_2898);
nand U2970 (N_2970,N_2902,N_2862);
nor U2971 (N_2971,N_2924,N_2923);
nand U2972 (N_2972,N_2863,N_2867);
and U2973 (N_2973,N_2910,N_2884);
and U2974 (N_2974,N_2861,N_2874);
nor U2975 (N_2975,N_2876,N_2881);
and U2976 (N_2976,N_2856,N_2859);
nand U2977 (N_2977,N_2909,N_2852);
nor U2978 (N_2978,N_2896,N_2862);
nor U2979 (N_2979,N_2921,N_2859);
nand U2980 (N_2980,N_2884,N_2887);
or U2981 (N_2981,N_2850,N_2899);
xor U2982 (N_2982,N_2920,N_2856);
and U2983 (N_2983,N_2897,N_2923);
nand U2984 (N_2984,N_2874,N_2889);
or U2985 (N_2985,N_2895,N_2880);
or U2986 (N_2986,N_2863,N_2887);
or U2987 (N_2987,N_2873,N_2896);
nor U2988 (N_2988,N_2918,N_2877);
or U2989 (N_2989,N_2863,N_2856);
nor U2990 (N_2990,N_2866,N_2872);
nor U2991 (N_2991,N_2916,N_2881);
nand U2992 (N_2992,N_2882,N_2922);
nand U2993 (N_2993,N_2852,N_2894);
or U2994 (N_2994,N_2867,N_2893);
nand U2995 (N_2995,N_2904,N_2895);
nand U2996 (N_2996,N_2863,N_2915);
and U2997 (N_2997,N_2910,N_2902);
and U2998 (N_2998,N_2899,N_2862);
or U2999 (N_2999,N_2886,N_2924);
and UO_0 (O_0,N_2953,N_2927);
or UO_1 (O_1,N_2951,N_2987);
nand UO_2 (O_2,N_2942,N_2941);
and UO_3 (O_3,N_2932,N_2970);
and UO_4 (O_4,N_2940,N_2943);
or UO_5 (O_5,N_2966,N_2939);
or UO_6 (O_6,N_2983,N_2946);
nand UO_7 (O_7,N_2992,N_2952);
nor UO_8 (O_8,N_2934,N_2949);
and UO_9 (O_9,N_2994,N_2989);
or UO_10 (O_10,N_2985,N_2997);
and UO_11 (O_11,N_2998,N_2945);
or UO_12 (O_12,N_2982,N_2977);
nand UO_13 (O_13,N_2926,N_2990);
and UO_14 (O_14,N_2981,N_2930);
or UO_15 (O_15,N_2986,N_2929);
nand UO_16 (O_16,N_2957,N_2962);
and UO_17 (O_17,N_2954,N_2980);
nor UO_18 (O_18,N_2956,N_2928);
or UO_19 (O_19,N_2961,N_2944);
and UO_20 (O_20,N_2971,N_2969);
nand UO_21 (O_21,N_2936,N_2938);
nand UO_22 (O_22,N_2972,N_2948);
and UO_23 (O_23,N_2955,N_2975);
or UO_24 (O_24,N_2964,N_2959);
or UO_25 (O_25,N_2937,N_2976);
nand UO_26 (O_26,N_2991,N_2950);
or UO_27 (O_27,N_2935,N_2965);
or UO_28 (O_28,N_2974,N_2967);
or UO_29 (O_29,N_2960,N_2988);
or UO_30 (O_30,N_2925,N_2993);
nor UO_31 (O_31,N_2973,N_2958);
nand UO_32 (O_32,N_2996,N_2963);
xor UO_33 (O_33,N_2968,N_2999);
and UO_34 (O_34,N_2931,N_2933);
and UO_35 (O_35,N_2995,N_2984);
and UO_36 (O_36,N_2979,N_2978);
nor UO_37 (O_37,N_2947,N_2944);
nand UO_38 (O_38,N_2931,N_2940);
xnor UO_39 (O_39,N_2997,N_2996);
nand UO_40 (O_40,N_2954,N_2979);
nor UO_41 (O_41,N_2969,N_2966);
or UO_42 (O_42,N_2935,N_2985);
nand UO_43 (O_43,N_2983,N_2999);
nand UO_44 (O_44,N_2987,N_2966);
nand UO_45 (O_45,N_2927,N_2965);
and UO_46 (O_46,N_2994,N_2944);
and UO_47 (O_47,N_2950,N_2956);
or UO_48 (O_48,N_2969,N_2965);
nor UO_49 (O_49,N_2947,N_2926);
nand UO_50 (O_50,N_2951,N_2932);
nor UO_51 (O_51,N_2949,N_2999);
or UO_52 (O_52,N_2961,N_2954);
or UO_53 (O_53,N_2930,N_2943);
and UO_54 (O_54,N_2953,N_2961);
nand UO_55 (O_55,N_2976,N_2962);
nand UO_56 (O_56,N_2927,N_2962);
or UO_57 (O_57,N_2925,N_2994);
nand UO_58 (O_58,N_2980,N_2987);
xor UO_59 (O_59,N_2950,N_2938);
nand UO_60 (O_60,N_2988,N_2972);
nand UO_61 (O_61,N_2998,N_2959);
nand UO_62 (O_62,N_2937,N_2997);
and UO_63 (O_63,N_2987,N_2934);
xor UO_64 (O_64,N_2975,N_2972);
nand UO_65 (O_65,N_2948,N_2954);
nor UO_66 (O_66,N_2980,N_2937);
and UO_67 (O_67,N_2932,N_2955);
or UO_68 (O_68,N_2996,N_2954);
and UO_69 (O_69,N_2945,N_2995);
or UO_70 (O_70,N_2959,N_2941);
nand UO_71 (O_71,N_2966,N_2934);
nand UO_72 (O_72,N_2934,N_2970);
nor UO_73 (O_73,N_2946,N_2940);
and UO_74 (O_74,N_2963,N_2964);
nor UO_75 (O_75,N_2925,N_2960);
nand UO_76 (O_76,N_2969,N_2934);
and UO_77 (O_77,N_2938,N_2967);
or UO_78 (O_78,N_2945,N_2978);
nor UO_79 (O_79,N_2965,N_2950);
nor UO_80 (O_80,N_2953,N_2990);
nand UO_81 (O_81,N_2986,N_2956);
nand UO_82 (O_82,N_2998,N_2952);
and UO_83 (O_83,N_2937,N_2954);
nor UO_84 (O_84,N_2945,N_2967);
or UO_85 (O_85,N_2975,N_2971);
or UO_86 (O_86,N_2958,N_2990);
or UO_87 (O_87,N_2979,N_2965);
nor UO_88 (O_88,N_2947,N_2986);
nand UO_89 (O_89,N_2954,N_2946);
nand UO_90 (O_90,N_2998,N_2958);
nand UO_91 (O_91,N_2950,N_2957);
and UO_92 (O_92,N_2972,N_2932);
nand UO_93 (O_93,N_2993,N_2994);
and UO_94 (O_94,N_2993,N_2970);
and UO_95 (O_95,N_2933,N_2930);
and UO_96 (O_96,N_2958,N_2928);
nand UO_97 (O_97,N_2987,N_2969);
nor UO_98 (O_98,N_2944,N_2968);
nor UO_99 (O_99,N_2968,N_2958);
nand UO_100 (O_100,N_2952,N_2991);
nand UO_101 (O_101,N_2951,N_2994);
or UO_102 (O_102,N_2932,N_2944);
and UO_103 (O_103,N_2956,N_2951);
nand UO_104 (O_104,N_2976,N_2975);
nor UO_105 (O_105,N_2970,N_2935);
nand UO_106 (O_106,N_2956,N_2964);
or UO_107 (O_107,N_2930,N_2936);
and UO_108 (O_108,N_2949,N_2950);
or UO_109 (O_109,N_2955,N_2949);
or UO_110 (O_110,N_2997,N_2955);
nand UO_111 (O_111,N_2971,N_2934);
and UO_112 (O_112,N_2974,N_2989);
and UO_113 (O_113,N_2969,N_2949);
and UO_114 (O_114,N_2992,N_2957);
xor UO_115 (O_115,N_2958,N_2992);
or UO_116 (O_116,N_2937,N_2999);
nor UO_117 (O_117,N_2932,N_2966);
or UO_118 (O_118,N_2929,N_2967);
and UO_119 (O_119,N_2973,N_2955);
and UO_120 (O_120,N_2933,N_2980);
nand UO_121 (O_121,N_2970,N_2974);
or UO_122 (O_122,N_2948,N_2991);
and UO_123 (O_123,N_2974,N_2983);
and UO_124 (O_124,N_2940,N_2962);
or UO_125 (O_125,N_2954,N_2999);
nand UO_126 (O_126,N_2926,N_2953);
and UO_127 (O_127,N_2944,N_2965);
nand UO_128 (O_128,N_2987,N_2978);
nand UO_129 (O_129,N_2942,N_2928);
xnor UO_130 (O_130,N_2950,N_2971);
nand UO_131 (O_131,N_2998,N_2935);
or UO_132 (O_132,N_2989,N_2931);
or UO_133 (O_133,N_2971,N_2998);
nor UO_134 (O_134,N_2980,N_2947);
or UO_135 (O_135,N_2994,N_2976);
nand UO_136 (O_136,N_2985,N_2971);
or UO_137 (O_137,N_2948,N_2975);
nor UO_138 (O_138,N_2997,N_2954);
or UO_139 (O_139,N_2959,N_2986);
nor UO_140 (O_140,N_2951,N_2976);
or UO_141 (O_141,N_2969,N_2940);
and UO_142 (O_142,N_2969,N_2962);
nand UO_143 (O_143,N_2946,N_2977);
or UO_144 (O_144,N_2970,N_2928);
or UO_145 (O_145,N_2966,N_2981);
nor UO_146 (O_146,N_2952,N_2947);
and UO_147 (O_147,N_2995,N_2969);
and UO_148 (O_148,N_2933,N_2969);
nor UO_149 (O_149,N_2987,N_2989);
or UO_150 (O_150,N_2980,N_2943);
or UO_151 (O_151,N_2982,N_2990);
or UO_152 (O_152,N_2954,N_2972);
or UO_153 (O_153,N_2966,N_2958);
and UO_154 (O_154,N_2950,N_2931);
nand UO_155 (O_155,N_2974,N_2949);
nand UO_156 (O_156,N_2939,N_2934);
and UO_157 (O_157,N_2949,N_2940);
nor UO_158 (O_158,N_2967,N_2944);
or UO_159 (O_159,N_2951,N_2945);
nor UO_160 (O_160,N_2963,N_2982);
xor UO_161 (O_161,N_2965,N_2989);
or UO_162 (O_162,N_2950,N_2983);
or UO_163 (O_163,N_2930,N_2996);
xnor UO_164 (O_164,N_2966,N_2936);
and UO_165 (O_165,N_2997,N_2976);
nand UO_166 (O_166,N_2977,N_2936);
xnor UO_167 (O_167,N_2969,N_2950);
nor UO_168 (O_168,N_2977,N_2960);
nor UO_169 (O_169,N_2987,N_2964);
and UO_170 (O_170,N_2938,N_2949);
nand UO_171 (O_171,N_2984,N_2982);
nor UO_172 (O_172,N_2979,N_2941);
and UO_173 (O_173,N_2967,N_2926);
nand UO_174 (O_174,N_2956,N_2955);
nor UO_175 (O_175,N_2951,N_2958);
and UO_176 (O_176,N_2937,N_2978);
and UO_177 (O_177,N_2928,N_2972);
nor UO_178 (O_178,N_2931,N_2973);
or UO_179 (O_179,N_2928,N_2945);
nor UO_180 (O_180,N_2946,N_2952);
or UO_181 (O_181,N_2973,N_2996);
or UO_182 (O_182,N_2993,N_2941);
nand UO_183 (O_183,N_2978,N_2988);
or UO_184 (O_184,N_2997,N_2928);
or UO_185 (O_185,N_2965,N_2936);
and UO_186 (O_186,N_2967,N_2930);
nor UO_187 (O_187,N_2961,N_2972);
xnor UO_188 (O_188,N_2979,N_2945);
and UO_189 (O_189,N_2976,N_2953);
nor UO_190 (O_190,N_2955,N_2959);
nor UO_191 (O_191,N_2955,N_2988);
nand UO_192 (O_192,N_2993,N_2986);
nand UO_193 (O_193,N_2997,N_2932);
nor UO_194 (O_194,N_2999,N_2961);
and UO_195 (O_195,N_2982,N_2972);
and UO_196 (O_196,N_2977,N_2998);
or UO_197 (O_197,N_2928,N_2936);
nand UO_198 (O_198,N_2988,N_2953);
nand UO_199 (O_199,N_2980,N_2955);
or UO_200 (O_200,N_2974,N_2966);
nor UO_201 (O_201,N_2980,N_2998);
nand UO_202 (O_202,N_2990,N_2963);
nand UO_203 (O_203,N_2952,N_2929);
and UO_204 (O_204,N_2957,N_2980);
nor UO_205 (O_205,N_2940,N_2986);
nor UO_206 (O_206,N_2996,N_2986);
nor UO_207 (O_207,N_2941,N_2970);
or UO_208 (O_208,N_2949,N_2927);
or UO_209 (O_209,N_2937,N_2931);
nand UO_210 (O_210,N_2985,N_2949);
nand UO_211 (O_211,N_2947,N_2948);
or UO_212 (O_212,N_2976,N_2980);
or UO_213 (O_213,N_2980,N_2978);
or UO_214 (O_214,N_2960,N_2974);
or UO_215 (O_215,N_2981,N_2949);
or UO_216 (O_216,N_2937,N_2958);
nor UO_217 (O_217,N_2999,N_2962);
and UO_218 (O_218,N_2998,N_2989);
nor UO_219 (O_219,N_2975,N_2987);
or UO_220 (O_220,N_2944,N_2952);
nor UO_221 (O_221,N_2927,N_2928);
nor UO_222 (O_222,N_2975,N_2925);
nor UO_223 (O_223,N_2937,N_2957);
nor UO_224 (O_224,N_2983,N_2937);
and UO_225 (O_225,N_2961,N_2951);
or UO_226 (O_226,N_2970,N_2946);
and UO_227 (O_227,N_2975,N_2952);
nor UO_228 (O_228,N_2982,N_2976);
and UO_229 (O_229,N_2943,N_2925);
nand UO_230 (O_230,N_2952,N_2978);
nor UO_231 (O_231,N_2938,N_2940);
or UO_232 (O_232,N_2949,N_2932);
and UO_233 (O_233,N_2966,N_2943);
or UO_234 (O_234,N_2933,N_2945);
nand UO_235 (O_235,N_2985,N_2982);
or UO_236 (O_236,N_2950,N_2952);
nand UO_237 (O_237,N_2987,N_2943);
nand UO_238 (O_238,N_2997,N_2974);
and UO_239 (O_239,N_2962,N_2968);
nor UO_240 (O_240,N_2941,N_2936);
nand UO_241 (O_241,N_2990,N_2968);
nor UO_242 (O_242,N_2989,N_2939);
or UO_243 (O_243,N_2973,N_2945);
or UO_244 (O_244,N_2974,N_2948);
nor UO_245 (O_245,N_2946,N_2926);
nand UO_246 (O_246,N_2960,N_2971);
nand UO_247 (O_247,N_2973,N_2932);
or UO_248 (O_248,N_2994,N_2961);
or UO_249 (O_249,N_2970,N_2977);
nor UO_250 (O_250,N_2964,N_2955);
nor UO_251 (O_251,N_2965,N_2931);
nor UO_252 (O_252,N_2950,N_2937);
nor UO_253 (O_253,N_2975,N_2974);
or UO_254 (O_254,N_2963,N_2936);
nor UO_255 (O_255,N_2996,N_2961);
nor UO_256 (O_256,N_2939,N_2960);
nor UO_257 (O_257,N_2997,N_2945);
nor UO_258 (O_258,N_2955,N_2934);
nor UO_259 (O_259,N_2975,N_2993);
and UO_260 (O_260,N_2995,N_2976);
xor UO_261 (O_261,N_2968,N_2947);
nor UO_262 (O_262,N_2991,N_2963);
or UO_263 (O_263,N_2958,N_2925);
and UO_264 (O_264,N_2983,N_2930);
xor UO_265 (O_265,N_2949,N_2928);
nor UO_266 (O_266,N_2954,N_2983);
and UO_267 (O_267,N_2981,N_2968);
and UO_268 (O_268,N_2980,N_2946);
nor UO_269 (O_269,N_2951,N_2946);
nor UO_270 (O_270,N_2974,N_2979);
nor UO_271 (O_271,N_2944,N_2943);
nand UO_272 (O_272,N_2948,N_2977);
nand UO_273 (O_273,N_2983,N_2995);
nand UO_274 (O_274,N_2992,N_2925);
nand UO_275 (O_275,N_2954,N_2939);
xor UO_276 (O_276,N_2942,N_2965);
and UO_277 (O_277,N_2929,N_2992);
and UO_278 (O_278,N_2956,N_2946);
xnor UO_279 (O_279,N_2983,N_2970);
and UO_280 (O_280,N_2948,N_2963);
or UO_281 (O_281,N_2948,N_2931);
nor UO_282 (O_282,N_2943,N_2975);
nand UO_283 (O_283,N_2958,N_2954);
and UO_284 (O_284,N_2955,N_2943);
nand UO_285 (O_285,N_2939,N_2935);
nand UO_286 (O_286,N_2961,N_2962);
and UO_287 (O_287,N_2931,N_2974);
nand UO_288 (O_288,N_2940,N_2944);
nor UO_289 (O_289,N_2996,N_2955);
or UO_290 (O_290,N_2941,N_2978);
nand UO_291 (O_291,N_2959,N_2999);
or UO_292 (O_292,N_2993,N_2976);
nor UO_293 (O_293,N_2940,N_2992);
nor UO_294 (O_294,N_2995,N_2979);
nor UO_295 (O_295,N_2931,N_2953);
or UO_296 (O_296,N_2998,N_2949);
nand UO_297 (O_297,N_2948,N_2950);
and UO_298 (O_298,N_2982,N_2987);
nand UO_299 (O_299,N_2946,N_2993);
nand UO_300 (O_300,N_2942,N_2951);
nand UO_301 (O_301,N_2975,N_2937);
nand UO_302 (O_302,N_2953,N_2974);
and UO_303 (O_303,N_2927,N_2995);
nor UO_304 (O_304,N_2987,N_2974);
nand UO_305 (O_305,N_2983,N_2988);
nor UO_306 (O_306,N_2949,N_2977);
or UO_307 (O_307,N_2993,N_2991);
or UO_308 (O_308,N_2979,N_2953);
and UO_309 (O_309,N_2993,N_2951);
nand UO_310 (O_310,N_2926,N_2935);
nand UO_311 (O_311,N_2964,N_2977);
nand UO_312 (O_312,N_2980,N_2985);
nand UO_313 (O_313,N_2932,N_2965);
nand UO_314 (O_314,N_2967,N_2979);
or UO_315 (O_315,N_2954,N_2992);
or UO_316 (O_316,N_2968,N_2948);
nor UO_317 (O_317,N_2940,N_2993);
or UO_318 (O_318,N_2934,N_2958);
nor UO_319 (O_319,N_2969,N_2931);
and UO_320 (O_320,N_2997,N_2943);
or UO_321 (O_321,N_2941,N_2957);
nand UO_322 (O_322,N_2953,N_2954);
nor UO_323 (O_323,N_2936,N_2950);
xor UO_324 (O_324,N_2925,N_2990);
and UO_325 (O_325,N_2947,N_2949);
and UO_326 (O_326,N_2925,N_2964);
nor UO_327 (O_327,N_2933,N_2977);
and UO_328 (O_328,N_2972,N_2998);
or UO_329 (O_329,N_2990,N_2994);
nor UO_330 (O_330,N_2977,N_2961);
nand UO_331 (O_331,N_2952,N_2979);
nor UO_332 (O_332,N_2930,N_2925);
and UO_333 (O_333,N_2936,N_2981);
and UO_334 (O_334,N_2950,N_2961);
nor UO_335 (O_335,N_2978,N_2984);
nor UO_336 (O_336,N_2980,N_2969);
nand UO_337 (O_337,N_2976,N_2978);
nor UO_338 (O_338,N_2938,N_2996);
nor UO_339 (O_339,N_2986,N_2970);
or UO_340 (O_340,N_2989,N_2996);
nand UO_341 (O_341,N_2949,N_2962);
nor UO_342 (O_342,N_2969,N_2926);
or UO_343 (O_343,N_2984,N_2959);
nand UO_344 (O_344,N_2936,N_2952);
xor UO_345 (O_345,N_2990,N_2995);
xor UO_346 (O_346,N_2960,N_2986);
or UO_347 (O_347,N_2937,N_2977);
and UO_348 (O_348,N_2948,N_2987);
nand UO_349 (O_349,N_2984,N_2963);
or UO_350 (O_350,N_2969,N_2925);
nor UO_351 (O_351,N_2947,N_2932);
nand UO_352 (O_352,N_2946,N_2933);
or UO_353 (O_353,N_2989,N_2957);
nor UO_354 (O_354,N_2957,N_2993);
nor UO_355 (O_355,N_2937,N_2995);
xor UO_356 (O_356,N_2952,N_2968);
or UO_357 (O_357,N_2965,N_2962);
nor UO_358 (O_358,N_2975,N_2929);
or UO_359 (O_359,N_2970,N_2937);
nand UO_360 (O_360,N_2930,N_2976);
nand UO_361 (O_361,N_2951,N_2964);
and UO_362 (O_362,N_2993,N_2966);
nand UO_363 (O_363,N_2931,N_2951);
nand UO_364 (O_364,N_2958,N_2965);
nor UO_365 (O_365,N_2930,N_2972);
xnor UO_366 (O_366,N_2938,N_2941);
nor UO_367 (O_367,N_2988,N_2990);
and UO_368 (O_368,N_2944,N_2999);
nor UO_369 (O_369,N_2925,N_2945);
nand UO_370 (O_370,N_2928,N_2971);
or UO_371 (O_371,N_2947,N_2970);
nand UO_372 (O_372,N_2965,N_2998);
nand UO_373 (O_373,N_2982,N_2940);
or UO_374 (O_374,N_2956,N_2943);
and UO_375 (O_375,N_2928,N_2967);
or UO_376 (O_376,N_2991,N_2962);
and UO_377 (O_377,N_2941,N_2939);
nor UO_378 (O_378,N_2957,N_2936);
nor UO_379 (O_379,N_2953,N_2950);
nor UO_380 (O_380,N_2966,N_2991);
and UO_381 (O_381,N_2995,N_2974);
nand UO_382 (O_382,N_2961,N_2931);
nand UO_383 (O_383,N_2942,N_2958);
or UO_384 (O_384,N_2939,N_2956);
nor UO_385 (O_385,N_2960,N_2976);
and UO_386 (O_386,N_2982,N_2927);
and UO_387 (O_387,N_2955,N_2995);
and UO_388 (O_388,N_2996,N_2933);
nor UO_389 (O_389,N_2931,N_2970);
nor UO_390 (O_390,N_2971,N_2956);
or UO_391 (O_391,N_2938,N_2943);
nand UO_392 (O_392,N_2939,N_2998);
and UO_393 (O_393,N_2942,N_2997);
or UO_394 (O_394,N_2988,N_2937);
nand UO_395 (O_395,N_2929,N_2971);
or UO_396 (O_396,N_2990,N_2978);
nand UO_397 (O_397,N_2993,N_2987);
and UO_398 (O_398,N_2992,N_2966);
or UO_399 (O_399,N_2958,N_2977);
nor UO_400 (O_400,N_2963,N_2970);
or UO_401 (O_401,N_2976,N_2981);
and UO_402 (O_402,N_2960,N_2953);
nand UO_403 (O_403,N_2992,N_2981);
or UO_404 (O_404,N_2960,N_2997);
or UO_405 (O_405,N_2948,N_2980);
nand UO_406 (O_406,N_2928,N_2976);
nor UO_407 (O_407,N_2926,N_2963);
nor UO_408 (O_408,N_2989,N_2983);
and UO_409 (O_409,N_2980,N_2973);
or UO_410 (O_410,N_2928,N_2941);
and UO_411 (O_411,N_2932,N_2930);
nor UO_412 (O_412,N_2948,N_2990);
nor UO_413 (O_413,N_2978,N_2959);
and UO_414 (O_414,N_2949,N_2954);
nor UO_415 (O_415,N_2927,N_2948);
and UO_416 (O_416,N_2949,N_2944);
nand UO_417 (O_417,N_2934,N_2940);
nor UO_418 (O_418,N_2961,N_2992);
xor UO_419 (O_419,N_2938,N_2992);
and UO_420 (O_420,N_2951,N_2959);
or UO_421 (O_421,N_2927,N_2963);
nor UO_422 (O_422,N_2952,N_2997);
nor UO_423 (O_423,N_2951,N_2963);
or UO_424 (O_424,N_2926,N_2966);
nor UO_425 (O_425,N_2990,N_2973);
nand UO_426 (O_426,N_2954,N_2947);
or UO_427 (O_427,N_2963,N_2954);
nor UO_428 (O_428,N_2933,N_2974);
nand UO_429 (O_429,N_2931,N_2964);
and UO_430 (O_430,N_2944,N_2936);
and UO_431 (O_431,N_2938,N_2978);
or UO_432 (O_432,N_2989,N_2975);
nand UO_433 (O_433,N_2927,N_2956);
nor UO_434 (O_434,N_2998,N_2938);
xnor UO_435 (O_435,N_2967,N_2951);
and UO_436 (O_436,N_2948,N_2959);
nor UO_437 (O_437,N_2984,N_2975);
nand UO_438 (O_438,N_2972,N_2966);
nand UO_439 (O_439,N_2994,N_2980);
nor UO_440 (O_440,N_2945,N_2965);
or UO_441 (O_441,N_2949,N_2965);
xor UO_442 (O_442,N_2931,N_2952);
nor UO_443 (O_443,N_2979,N_2970);
nor UO_444 (O_444,N_2968,N_2930);
nor UO_445 (O_445,N_2967,N_2956);
and UO_446 (O_446,N_2974,N_2938);
or UO_447 (O_447,N_2950,N_2993);
nand UO_448 (O_448,N_2930,N_2965);
and UO_449 (O_449,N_2972,N_2943);
and UO_450 (O_450,N_2989,N_2970);
nor UO_451 (O_451,N_2965,N_2966);
nor UO_452 (O_452,N_2933,N_2960);
nand UO_453 (O_453,N_2986,N_2932);
nand UO_454 (O_454,N_2933,N_2928);
nand UO_455 (O_455,N_2959,N_2981);
or UO_456 (O_456,N_2963,N_2949);
xor UO_457 (O_457,N_2967,N_2989);
nand UO_458 (O_458,N_2950,N_2999);
or UO_459 (O_459,N_2945,N_2975);
or UO_460 (O_460,N_2963,N_2976);
and UO_461 (O_461,N_2941,N_2934);
and UO_462 (O_462,N_2935,N_2993);
or UO_463 (O_463,N_2966,N_2933);
or UO_464 (O_464,N_2959,N_2953);
or UO_465 (O_465,N_2989,N_2936);
and UO_466 (O_466,N_2999,N_2990);
nand UO_467 (O_467,N_2943,N_2937);
and UO_468 (O_468,N_2992,N_2994);
or UO_469 (O_469,N_2971,N_2931);
or UO_470 (O_470,N_2965,N_2994);
or UO_471 (O_471,N_2959,N_2960);
nand UO_472 (O_472,N_2955,N_2967);
and UO_473 (O_473,N_2945,N_2993);
nor UO_474 (O_474,N_2990,N_2987);
nor UO_475 (O_475,N_2937,N_2973);
and UO_476 (O_476,N_2935,N_2937);
or UO_477 (O_477,N_2989,N_2985);
or UO_478 (O_478,N_2932,N_2998);
nand UO_479 (O_479,N_2988,N_2944);
or UO_480 (O_480,N_2963,N_2968);
nand UO_481 (O_481,N_2979,N_2930);
nand UO_482 (O_482,N_2937,N_2932);
nand UO_483 (O_483,N_2940,N_2989);
nor UO_484 (O_484,N_2984,N_2931);
and UO_485 (O_485,N_2975,N_2963);
and UO_486 (O_486,N_2952,N_2938);
nand UO_487 (O_487,N_2978,N_2956);
or UO_488 (O_488,N_2988,N_2964);
nand UO_489 (O_489,N_2965,N_2941);
nand UO_490 (O_490,N_2941,N_2990);
or UO_491 (O_491,N_2974,N_2990);
or UO_492 (O_492,N_2957,N_2930);
and UO_493 (O_493,N_2953,N_2944);
xor UO_494 (O_494,N_2989,N_2963);
and UO_495 (O_495,N_2975,N_2933);
nand UO_496 (O_496,N_2933,N_2971);
nor UO_497 (O_497,N_2929,N_2959);
or UO_498 (O_498,N_2930,N_2926);
and UO_499 (O_499,N_2949,N_2987);
endmodule