module basic_500_3000_500_5_levels_1xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_15,In_200);
nor U1 (N_1,In_112,In_263);
nand U2 (N_2,In_34,In_226);
and U3 (N_3,In_285,In_238);
or U4 (N_4,In_356,In_295);
or U5 (N_5,In_355,In_360);
nor U6 (N_6,In_66,In_114);
nand U7 (N_7,In_10,In_385);
or U8 (N_8,In_165,In_202);
nand U9 (N_9,In_391,In_225);
or U10 (N_10,In_250,In_161);
and U11 (N_11,In_81,In_57);
nor U12 (N_12,In_466,In_462);
and U13 (N_13,In_231,In_369);
nand U14 (N_14,In_128,In_299);
and U15 (N_15,In_451,In_72);
or U16 (N_16,In_396,In_311);
and U17 (N_17,In_46,In_68);
nand U18 (N_18,In_418,In_472);
and U19 (N_19,In_327,In_48);
nand U20 (N_20,In_398,In_133);
nor U21 (N_21,In_42,In_292);
nor U22 (N_22,In_450,In_305);
or U23 (N_23,In_468,In_452);
and U24 (N_24,In_24,In_111);
and U25 (N_25,In_340,In_213);
and U26 (N_26,In_415,In_393);
or U27 (N_27,In_100,In_384);
nand U28 (N_28,In_125,In_307);
or U29 (N_29,In_475,In_117);
or U30 (N_30,In_409,In_363);
or U31 (N_31,In_245,In_493);
nand U32 (N_32,In_23,In_35);
nor U33 (N_33,In_487,In_205);
nor U34 (N_34,In_341,In_139);
and U35 (N_35,In_51,In_364);
and U36 (N_36,In_412,In_84);
nor U37 (N_37,In_346,In_416);
nor U38 (N_38,In_436,In_435);
or U39 (N_39,In_306,In_214);
and U40 (N_40,In_287,In_293);
and U41 (N_41,In_316,In_454);
or U42 (N_42,In_38,In_58);
nor U43 (N_43,In_300,In_65);
or U44 (N_44,In_290,In_267);
and U45 (N_45,In_163,In_473);
and U46 (N_46,In_484,In_60);
nor U47 (N_47,In_107,In_188);
nor U48 (N_48,In_234,In_130);
nand U49 (N_49,In_467,In_414);
or U50 (N_50,In_89,In_104);
nor U51 (N_51,In_144,In_464);
nor U52 (N_52,In_294,In_52);
nand U53 (N_53,In_434,In_322);
nand U54 (N_54,In_64,In_93);
and U55 (N_55,In_183,In_1);
or U56 (N_56,In_198,In_395);
nand U57 (N_57,In_430,In_116);
or U58 (N_58,In_349,In_187);
or U59 (N_59,In_439,In_204);
nand U60 (N_60,In_63,In_129);
and U61 (N_61,In_374,In_312);
nor U62 (N_62,In_173,In_304);
and U63 (N_63,In_315,In_458);
nor U64 (N_64,In_397,In_403);
nand U65 (N_65,In_386,In_195);
nand U66 (N_66,In_302,In_149);
nand U67 (N_67,In_266,In_309);
nor U68 (N_68,In_207,In_498);
and U69 (N_69,In_423,In_441);
or U70 (N_70,In_120,In_495);
nor U71 (N_71,In_275,In_438);
nand U72 (N_72,In_460,In_227);
and U73 (N_73,In_158,In_99);
or U74 (N_74,In_352,In_235);
nand U75 (N_75,In_419,In_79);
nand U76 (N_76,In_87,In_328);
or U77 (N_77,In_37,In_444);
nor U78 (N_78,In_206,In_478);
nand U79 (N_79,In_319,In_85);
nor U80 (N_80,In_69,In_445);
or U81 (N_81,In_230,In_176);
nand U82 (N_82,In_368,In_31);
nor U83 (N_83,In_494,In_102);
and U84 (N_84,In_210,In_410);
and U85 (N_85,In_110,In_83);
or U86 (N_86,In_192,In_255);
or U87 (N_87,In_407,In_461);
or U88 (N_88,In_481,In_406);
nand U89 (N_89,In_80,In_166);
or U90 (N_90,In_490,In_348);
or U91 (N_91,In_359,In_417);
and U92 (N_92,In_94,In_208);
nand U93 (N_93,In_443,In_145);
nor U94 (N_94,In_6,In_201);
nand U95 (N_95,In_103,In_193);
nand U96 (N_96,In_408,In_222);
nor U97 (N_97,In_279,In_218);
or U98 (N_98,In_480,In_215);
or U99 (N_99,In_182,In_345);
nor U100 (N_100,In_330,In_421);
and U101 (N_101,In_162,In_278);
and U102 (N_102,In_124,In_17);
or U103 (N_103,In_350,In_113);
and U104 (N_104,In_194,In_358);
nand U105 (N_105,In_269,In_197);
nand U106 (N_106,In_123,In_317);
or U107 (N_107,In_366,In_164);
or U108 (N_108,In_96,In_394);
nand U109 (N_109,In_339,In_171);
nor U110 (N_110,In_244,In_212);
and U111 (N_111,In_281,In_390);
nand U112 (N_112,In_282,In_26);
or U113 (N_113,In_343,In_224);
nor U114 (N_114,In_260,In_297);
and U115 (N_115,In_97,In_486);
xnor U116 (N_116,In_74,In_335);
or U117 (N_117,In_86,In_70);
and U118 (N_118,In_424,In_8);
or U119 (N_119,In_411,In_399);
and U120 (N_120,In_331,In_247);
nor U121 (N_121,In_361,In_453);
nor U122 (N_122,In_143,In_254);
and U123 (N_123,In_199,In_457);
or U124 (N_124,In_387,In_404);
or U125 (N_125,In_320,In_392);
and U126 (N_126,In_9,In_49);
nor U127 (N_127,In_376,In_431);
nor U128 (N_128,In_88,In_174);
nand U129 (N_129,In_463,In_177);
and U130 (N_130,In_126,In_39);
nand U131 (N_131,In_437,In_142);
or U132 (N_132,In_185,In_119);
nor U133 (N_133,In_179,In_11);
and U134 (N_134,In_14,In_334);
and U135 (N_135,In_134,In_379);
nand U136 (N_136,In_427,In_95);
and U137 (N_137,In_276,In_135);
nor U138 (N_138,In_242,In_347);
nor U139 (N_139,In_170,In_249);
or U140 (N_140,In_389,In_21);
nand U141 (N_141,In_483,In_273);
and U142 (N_142,In_258,In_20);
or U143 (N_143,In_301,In_122);
or U144 (N_144,In_474,In_61);
nand U145 (N_145,In_446,In_271);
nor U146 (N_146,In_148,In_105);
nand U147 (N_147,In_353,In_18);
nor U148 (N_148,In_367,In_108);
nand U149 (N_149,In_73,In_283);
or U150 (N_150,In_413,In_77);
nand U151 (N_151,In_455,In_132);
or U152 (N_152,In_286,In_45);
or U153 (N_153,In_448,In_482);
or U154 (N_154,In_190,In_370);
nor U155 (N_155,In_318,In_137);
xnor U156 (N_156,In_262,In_28);
or U157 (N_157,In_337,In_447);
nor U158 (N_158,In_402,In_47);
or U159 (N_159,In_30,In_67);
and U160 (N_160,In_338,In_203);
or U161 (N_161,In_155,In_90);
nor U162 (N_162,In_159,In_2);
xor U163 (N_163,In_496,In_432);
and U164 (N_164,In_19,In_118);
nor U165 (N_165,In_378,In_284);
or U166 (N_166,In_13,In_181);
or U167 (N_167,In_219,In_371);
or U168 (N_168,In_25,In_54);
or U169 (N_169,In_237,In_32);
and U170 (N_170,In_36,In_405);
nor U171 (N_171,In_167,In_138);
and U172 (N_172,In_157,In_153);
nand U173 (N_173,In_440,In_109);
or U174 (N_174,In_277,In_325);
nor U175 (N_175,In_296,In_429);
nor U176 (N_176,In_78,In_16);
and U177 (N_177,In_252,In_489);
nand U178 (N_178,In_485,In_336);
and U179 (N_179,In_229,In_146);
or U180 (N_180,In_33,In_92);
and U181 (N_181,In_191,In_426);
or U182 (N_182,In_127,In_27);
and U183 (N_183,In_469,In_324);
nand U184 (N_184,In_383,In_216);
nand U185 (N_185,In_470,In_270);
nand U186 (N_186,In_178,In_329);
nor U187 (N_187,In_168,In_131);
or U188 (N_188,In_43,In_420);
nor U189 (N_189,In_156,In_151);
nor U190 (N_190,In_152,In_442);
and U191 (N_191,In_180,In_459);
or U192 (N_192,In_3,In_248);
or U193 (N_193,In_140,In_209);
nor U194 (N_194,In_221,In_184);
nand U195 (N_195,In_56,In_351);
nand U196 (N_196,In_326,In_342);
and U197 (N_197,In_401,In_241);
and U198 (N_198,In_240,In_233);
nor U199 (N_199,In_53,In_465);
or U200 (N_200,In_422,In_253);
nand U201 (N_201,In_154,In_115);
and U202 (N_202,In_232,In_449);
or U203 (N_203,In_136,In_388);
or U204 (N_204,In_280,In_313);
and U205 (N_205,In_344,In_476);
nor U206 (N_206,In_332,In_62);
nor U207 (N_207,In_7,In_499);
or U208 (N_208,In_268,In_425);
or U209 (N_209,In_76,In_22);
or U210 (N_210,In_372,In_175);
nand U211 (N_211,In_217,In_75);
or U212 (N_212,In_354,In_196);
and U213 (N_213,In_259,In_186);
or U214 (N_214,In_4,In_5);
nand U215 (N_215,In_55,In_381);
or U216 (N_216,In_172,In_101);
and U217 (N_217,In_373,In_160);
nor U218 (N_218,In_479,In_121);
and U219 (N_219,In_380,In_223);
or U220 (N_220,In_492,In_147);
nor U221 (N_221,In_0,In_243);
and U222 (N_222,In_211,In_272);
nand U223 (N_223,In_323,In_497);
or U224 (N_224,In_98,In_236);
or U225 (N_225,In_433,In_264);
or U226 (N_226,In_428,In_357);
nor U227 (N_227,In_169,In_375);
or U228 (N_228,In_71,In_298);
nand U229 (N_229,In_456,In_29);
xor U230 (N_230,In_261,In_220);
and U231 (N_231,In_257,In_310);
nand U232 (N_232,In_106,In_12);
nand U233 (N_233,In_228,In_303);
or U234 (N_234,In_40,In_488);
or U235 (N_235,In_189,In_321);
or U236 (N_236,In_91,In_471);
and U237 (N_237,In_251,In_265);
and U238 (N_238,In_377,In_50);
or U239 (N_239,In_288,In_289);
or U240 (N_240,In_362,In_308);
nand U241 (N_241,In_382,In_491);
nand U242 (N_242,In_291,In_141);
and U243 (N_243,In_82,In_150);
nor U244 (N_244,In_365,In_41);
or U245 (N_245,In_274,In_477);
xnor U246 (N_246,In_239,In_59);
and U247 (N_247,In_256,In_400);
nor U248 (N_248,In_246,In_333);
and U249 (N_249,In_314,In_44);
or U250 (N_250,In_150,In_5);
and U251 (N_251,In_206,In_117);
or U252 (N_252,In_407,In_292);
and U253 (N_253,In_140,In_49);
or U254 (N_254,In_431,In_155);
or U255 (N_255,In_182,In_485);
nand U256 (N_256,In_475,In_262);
and U257 (N_257,In_108,In_141);
and U258 (N_258,In_10,In_125);
and U259 (N_259,In_107,In_493);
nor U260 (N_260,In_222,In_213);
and U261 (N_261,In_352,In_279);
or U262 (N_262,In_265,In_91);
nand U263 (N_263,In_319,In_30);
or U264 (N_264,In_320,In_207);
and U265 (N_265,In_409,In_118);
or U266 (N_266,In_271,In_96);
and U267 (N_267,In_292,In_481);
nand U268 (N_268,In_440,In_197);
and U269 (N_269,In_271,In_292);
or U270 (N_270,In_488,In_290);
nor U271 (N_271,In_460,In_325);
nor U272 (N_272,In_405,In_331);
and U273 (N_273,In_487,In_401);
and U274 (N_274,In_118,In_288);
and U275 (N_275,In_0,In_137);
and U276 (N_276,In_92,In_221);
nand U277 (N_277,In_123,In_398);
nor U278 (N_278,In_287,In_192);
and U279 (N_279,In_221,In_224);
nor U280 (N_280,In_344,In_304);
or U281 (N_281,In_484,In_22);
or U282 (N_282,In_376,In_458);
and U283 (N_283,In_43,In_280);
nor U284 (N_284,In_19,In_254);
nand U285 (N_285,In_203,In_319);
or U286 (N_286,In_228,In_481);
and U287 (N_287,In_291,In_179);
nor U288 (N_288,In_174,In_12);
nand U289 (N_289,In_244,In_287);
nor U290 (N_290,In_89,In_455);
nand U291 (N_291,In_106,In_308);
or U292 (N_292,In_423,In_475);
or U293 (N_293,In_360,In_398);
and U294 (N_294,In_55,In_430);
nand U295 (N_295,In_309,In_137);
nand U296 (N_296,In_291,In_209);
or U297 (N_297,In_274,In_45);
and U298 (N_298,In_65,In_97);
nand U299 (N_299,In_355,In_426);
and U300 (N_300,In_141,In_183);
or U301 (N_301,In_210,In_167);
nand U302 (N_302,In_204,In_153);
nand U303 (N_303,In_428,In_335);
nand U304 (N_304,In_360,In_106);
nand U305 (N_305,In_66,In_398);
and U306 (N_306,In_419,In_118);
nand U307 (N_307,In_84,In_93);
and U308 (N_308,In_331,In_13);
nor U309 (N_309,In_332,In_48);
nor U310 (N_310,In_36,In_245);
nand U311 (N_311,In_124,In_29);
or U312 (N_312,In_452,In_250);
nor U313 (N_313,In_186,In_263);
xor U314 (N_314,In_325,In_218);
nand U315 (N_315,In_470,In_267);
nand U316 (N_316,In_431,In_249);
nor U317 (N_317,In_163,In_264);
nor U318 (N_318,In_103,In_462);
and U319 (N_319,In_496,In_404);
nor U320 (N_320,In_462,In_137);
nor U321 (N_321,In_163,In_56);
nor U322 (N_322,In_262,In_25);
nor U323 (N_323,In_347,In_236);
or U324 (N_324,In_291,In_165);
nor U325 (N_325,In_296,In_197);
nor U326 (N_326,In_162,In_95);
nand U327 (N_327,In_418,In_409);
or U328 (N_328,In_368,In_432);
nand U329 (N_329,In_320,In_211);
or U330 (N_330,In_309,In_185);
nor U331 (N_331,In_238,In_63);
nand U332 (N_332,In_375,In_205);
nor U333 (N_333,In_182,In_474);
nor U334 (N_334,In_350,In_414);
nand U335 (N_335,In_450,In_14);
or U336 (N_336,In_233,In_247);
nand U337 (N_337,In_309,In_258);
nor U338 (N_338,In_89,In_139);
nand U339 (N_339,In_419,In_198);
and U340 (N_340,In_13,In_26);
nor U341 (N_341,In_126,In_80);
nand U342 (N_342,In_241,In_453);
nor U343 (N_343,In_230,In_47);
nor U344 (N_344,In_375,In_151);
nor U345 (N_345,In_472,In_64);
and U346 (N_346,In_317,In_95);
or U347 (N_347,In_381,In_88);
or U348 (N_348,In_444,In_143);
nand U349 (N_349,In_194,In_91);
nor U350 (N_350,In_139,In_206);
xor U351 (N_351,In_252,In_155);
nand U352 (N_352,In_109,In_412);
nor U353 (N_353,In_1,In_388);
or U354 (N_354,In_496,In_422);
and U355 (N_355,In_44,In_371);
and U356 (N_356,In_229,In_98);
nor U357 (N_357,In_431,In_135);
or U358 (N_358,In_276,In_422);
and U359 (N_359,In_12,In_391);
nand U360 (N_360,In_372,In_269);
nor U361 (N_361,In_212,In_246);
and U362 (N_362,In_342,In_329);
xor U363 (N_363,In_236,In_146);
nor U364 (N_364,In_140,In_67);
nand U365 (N_365,In_269,In_335);
nor U366 (N_366,In_200,In_52);
nand U367 (N_367,In_225,In_459);
nor U368 (N_368,In_120,In_165);
nor U369 (N_369,In_353,In_339);
or U370 (N_370,In_361,In_272);
and U371 (N_371,In_283,In_206);
nor U372 (N_372,In_136,In_399);
or U373 (N_373,In_20,In_58);
and U374 (N_374,In_198,In_281);
and U375 (N_375,In_365,In_441);
and U376 (N_376,In_454,In_458);
nand U377 (N_377,In_307,In_20);
or U378 (N_378,In_276,In_480);
nor U379 (N_379,In_23,In_343);
and U380 (N_380,In_370,In_227);
nor U381 (N_381,In_211,In_84);
or U382 (N_382,In_250,In_307);
and U383 (N_383,In_151,In_436);
or U384 (N_384,In_203,In_72);
and U385 (N_385,In_98,In_76);
nand U386 (N_386,In_184,In_289);
nor U387 (N_387,In_199,In_53);
and U388 (N_388,In_144,In_307);
and U389 (N_389,In_390,In_317);
or U390 (N_390,In_138,In_34);
or U391 (N_391,In_476,In_70);
and U392 (N_392,In_250,In_123);
nor U393 (N_393,In_27,In_391);
and U394 (N_394,In_39,In_307);
nor U395 (N_395,In_361,In_130);
nor U396 (N_396,In_32,In_267);
and U397 (N_397,In_322,In_113);
or U398 (N_398,In_383,In_247);
nor U399 (N_399,In_370,In_475);
and U400 (N_400,In_306,In_395);
nand U401 (N_401,In_437,In_80);
nand U402 (N_402,In_284,In_83);
nand U403 (N_403,In_398,In_6);
or U404 (N_404,In_26,In_394);
or U405 (N_405,In_403,In_380);
and U406 (N_406,In_22,In_331);
or U407 (N_407,In_298,In_105);
nor U408 (N_408,In_40,In_280);
or U409 (N_409,In_365,In_307);
or U410 (N_410,In_350,In_490);
nand U411 (N_411,In_94,In_146);
and U412 (N_412,In_394,In_25);
nand U413 (N_413,In_43,In_90);
nor U414 (N_414,In_273,In_65);
nand U415 (N_415,In_93,In_327);
nor U416 (N_416,In_359,In_294);
nand U417 (N_417,In_267,In_162);
nand U418 (N_418,In_439,In_1);
nor U419 (N_419,In_131,In_262);
or U420 (N_420,In_112,In_457);
and U421 (N_421,In_222,In_14);
nand U422 (N_422,In_171,In_189);
nand U423 (N_423,In_105,In_385);
or U424 (N_424,In_275,In_160);
and U425 (N_425,In_468,In_157);
and U426 (N_426,In_22,In_135);
nor U427 (N_427,In_448,In_338);
nand U428 (N_428,In_388,In_118);
nor U429 (N_429,In_227,In_402);
and U430 (N_430,In_183,In_300);
nand U431 (N_431,In_157,In_378);
nand U432 (N_432,In_10,In_452);
and U433 (N_433,In_287,In_209);
nor U434 (N_434,In_191,In_283);
nor U435 (N_435,In_398,In_117);
nand U436 (N_436,In_454,In_91);
nand U437 (N_437,In_165,In_320);
nand U438 (N_438,In_10,In_378);
or U439 (N_439,In_142,In_255);
nor U440 (N_440,In_265,In_470);
or U441 (N_441,In_98,In_240);
and U442 (N_442,In_384,In_472);
or U443 (N_443,In_490,In_329);
and U444 (N_444,In_435,In_209);
or U445 (N_445,In_423,In_376);
nor U446 (N_446,In_372,In_339);
nor U447 (N_447,In_72,In_332);
nand U448 (N_448,In_251,In_249);
nor U449 (N_449,In_151,In_434);
nand U450 (N_450,In_170,In_151);
and U451 (N_451,In_102,In_410);
nand U452 (N_452,In_175,In_279);
nand U453 (N_453,In_271,In_51);
nand U454 (N_454,In_428,In_188);
nand U455 (N_455,In_152,In_5);
or U456 (N_456,In_252,In_286);
nor U457 (N_457,In_490,In_102);
nand U458 (N_458,In_153,In_149);
or U459 (N_459,In_358,In_340);
nor U460 (N_460,In_443,In_389);
nor U461 (N_461,In_155,In_186);
or U462 (N_462,In_342,In_279);
or U463 (N_463,In_191,In_396);
nand U464 (N_464,In_445,In_432);
nand U465 (N_465,In_185,In_187);
nor U466 (N_466,In_196,In_82);
and U467 (N_467,In_491,In_40);
or U468 (N_468,In_50,In_366);
nor U469 (N_469,In_439,In_253);
nor U470 (N_470,In_24,In_110);
and U471 (N_471,In_443,In_284);
and U472 (N_472,In_259,In_388);
nand U473 (N_473,In_419,In_181);
or U474 (N_474,In_435,In_476);
nor U475 (N_475,In_449,In_441);
nand U476 (N_476,In_38,In_112);
nand U477 (N_477,In_304,In_445);
or U478 (N_478,In_135,In_92);
and U479 (N_479,In_311,In_228);
and U480 (N_480,In_304,In_342);
and U481 (N_481,In_226,In_299);
nor U482 (N_482,In_166,In_243);
nor U483 (N_483,In_96,In_387);
nor U484 (N_484,In_234,In_379);
nand U485 (N_485,In_320,In_1);
nor U486 (N_486,In_248,In_131);
or U487 (N_487,In_376,In_259);
or U488 (N_488,In_11,In_453);
and U489 (N_489,In_21,In_393);
or U490 (N_490,In_45,In_287);
or U491 (N_491,In_442,In_479);
or U492 (N_492,In_426,In_238);
nand U493 (N_493,In_140,In_223);
xor U494 (N_494,In_334,In_319);
nand U495 (N_495,In_250,In_279);
nor U496 (N_496,In_168,In_163);
nand U497 (N_497,In_261,In_110);
nand U498 (N_498,In_144,In_176);
or U499 (N_499,In_165,In_236);
and U500 (N_500,In_197,In_224);
nand U501 (N_501,In_429,In_15);
and U502 (N_502,In_250,In_105);
nor U503 (N_503,In_34,In_274);
nor U504 (N_504,In_50,In_51);
nor U505 (N_505,In_440,In_81);
nor U506 (N_506,In_426,In_470);
nand U507 (N_507,In_47,In_432);
or U508 (N_508,In_83,In_5);
nor U509 (N_509,In_330,In_65);
nor U510 (N_510,In_494,In_230);
nor U511 (N_511,In_208,In_2);
or U512 (N_512,In_36,In_287);
nor U513 (N_513,In_356,In_229);
nor U514 (N_514,In_230,In_229);
nand U515 (N_515,In_193,In_206);
and U516 (N_516,In_68,In_284);
nand U517 (N_517,In_143,In_160);
or U518 (N_518,In_70,In_354);
and U519 (N_519,In_409,In_308);
or U520 (N_520,In_424,In_494);
and U521 (N_521,In_280,In_147);
nand U522 (N_522,In_13,In_119);
and U523 (N_523,In_139,In_391);
nor U524 (N_524,In_143,In_2);
nor U525 (N_525,In_53,In_163);
nand U526 (N_526,In_480,In_141);
nand U527 (N_527,In_492,In_291);
xor U528 (N_528,In_377,In_491);
nand U529 (N_529,In_53,In_368);
nand U530 (N_530,In_482,In_383);
xor U531 (N_531,In_178,In_27);
nor U532 (N_532,In_4,In_468);
nor U533 (N_533,In_455,In_289);
nand U534 (N_534,In_158,In_367);
or U535 (N_535,In_173,In_156);
nand U536 (N_536,In_38,In_341);
or U537 (N_537,In_154,In_455);
and U538 (N_538,In_287,In_65);
and U539 (N_539,In_220,In_301);
or U540 (N_540,In_103,In_89);
or U541 (N_541,In_279,In_169);
nand U542 (N_542,In_335,In_254);
nand U543 (N_543,In_193,In_365);
nor U544 (N_544,In_237,In_262);
or U545 (N_545,In_484,In_273);
nand U546 (N_546,In_476,In_498);
or U547 (N_547,In_246,In_335);
nor U548 (N_548,In_325,In_350);
nor U549 (N_549,In_288,In_498);
nand U550 (N_550,In_495,In_160);
and U551 (N_551,In_346,In_467);
or U552 (N_552,In_302,In_376);
nor U553 (N_553,In_272,In_146);
or U554 (N_554,In_47,In_484);
and U555 (N_555,In_444,In_237);
and U556 (N_556,In_116,In_335);
or U557 (N_557,In_352,In_379);
nor U558 (N_558,In_46,In_488);
nand U559 (N_559,In_455,In_106);
and U560 (N_560,In_125,In_485);
or U561 (N_561,In_235,In_484);
nand U562 (N_562,In_234,In_335);
and U563 (N_563,In_29,In_323);
and U564 (N_564,In_291,In_56);
or U565 (N_565,In_77,In_254);
nor U566 (N_566,In_292,In_423);
or U567 (N_567,In_453,In_192);
and U568 (N_568,In_268,In_315);
and U569 (N_569,In_368,In_379);
nor U570 (N_570,In_86,In_37);
nand U571 (N_571,In_36,In_289);
or U572 (N_572,In_461,In_151);
and U573 (N_573,In_223,In_374);
nor U574 (N_574,In_164,In_487);
or U575 (N_575,In_116,In_459);
and U576 (N_576,In_195,In_456);
and U577 (N_577,In_278,In_193);
nand U578 (N_578,In_110,In_423);
or U579 (N_579,In_57,In_35);
or U580 (N_580,In_44,In_160);
nand U581 (N_581,In_28,In_58);
or U582 (N_582,In_17,In_227);
nand U583 (N_583,In_462,In_372);
and U584 (N_584,In_368,In_388);
nand U585 (N_585,In_405,In_9);
nand U586 (N_586,In_65,In_446);
or U587 (N_587,In_3,In_200);
and U588 (N_588,In_128,In_429);
or U589 (N_589,In_315,In_296);
nand U590 (N_590,In_294,In_484);
nor U591 (N_591,In_242,In_141);
nor U592 (N_592,In_23,In_137);
nand U593 (N_593,In_251,In_203);
nand U594 (N_594,In_193,In_346);
and U595 (N_595,In_195,In_186);
or U596 (N_596,In_323,In_239);
nand U597 (N_597,In_323,In_364);
or U598 (N_598,In_427,In_245);
or U599 (N_599,In_93,In_30);
nand U600 (N_600,N_85,N_567);
or U601 (N_601,N_137,N_460);
nor U602 (N_602,N_475,N_100);
nor U603 (N_603,N_305,N_283);
or U604 (N_604,N_144,N_483);
nand U605 (N_605,N_196,N_2);
nor U606 (N_606,N_353,N_220);
and U607 (N_607,N_117,N_288);
or U608 (N_608,N_159,N_20);
or U609 (N_609,N_512,N_214);
nor U610 (N_610,N_356,N_556);
nor U611 (N_611,N_366,N_435);
or U612 (N_612,N_420,N_527);
or U613 (N_613,N_273,N_439);
or U614 (N_614,N_393,N_42);
nor U615 (N_615,N_205,N_275);
nor U616 (N_616,N_184,N_230);
or U617 (N_617,N_339,N_331);
and U618 (N_618,N_583,N_368);
or U619 (N_619,N_412,N_555);
and U620 (N_620,N_183,N_354);
or U621 (N_621,N_156,N_161);
nand U622 (N_622,N_461,N_493);
nor U623 (N_623,N_396,N_350);
and U624 (N_624,N_302,N_223);
or U625 (N_625,N_232,N_581);
or U626 (N_626,N_180,N_484);
or U627 (N_627,N_456,N_268);
or U628 (N_628,N_375,N_434);
and U629 (N_629,N_4,N_291);
or U630 (N_630,N_332,N_152);
nor U631 (N_631,N_29,N_228);
and U632 (N_632,N_229,N_351);
nand U633 (N_633,N_433,N_364);
nor U634 (N_634,N_300,N_469);
nor U635 (N_635,N_150,N_127);
and U636 (N_636,N_316,N_132);
nand U637 (N_637,N_576,N_188);
nand U638 (N_638,N_352,N_432);
nor U639 (N_639,N_525,N_538);
nor U640 (N_640,N_546,N_245);
and U641 (N_641,N_450,N_293);
or U642 (N_642,N_187,N_67);
or U643 (N_643,N_145,N_406);
nor U644 (N_644,N_135,N_90);
nand U645 (N_645,N_219,N_358);
and U646 (N_646,N_410,N_570);
and U647 (N_647,N_382,N_598);
or U648 (N_648,N_215,N_237);
nor U649 (N_649,N_56,N_421);
nand U650 (N_650,N_343,N_249);
or U651 (N_651,N_338,N_348);
nor U652 (N_652,N_323,N_270);
and U653 (N_653,N_235,N_169);
nand U654 (N_654,N_349,N_592);
xnor U655 (N_655,N_22,N_513);
and U656 (N_656,N_458,N_203);
and U657 (N_657,N_381,N_129);
or U658 (N_658,N_7,N_44);
or U659 (N_659,N_492,N_560);
and U660 (N_660,N_191,N_51);
nand U661 (N_661,N_452,N_542);
and U662 (N_662,N_280,N_134);
and U663 (N_663,N_502,N_176);
nor U664 (N_664,N_45,N_199);
xnor U665 (N_665,N_447,N_562);
or U666 (N_666,N_247,N_102);
nand U667 (N_667,N_437,N_5);
or U668 (N_668,N_455,N_372);
or U669 (N_669,N_553,N_27);
and U670 (N_670,N_278,N_321);
or U671 (N_671,N_106,N_197);
nand U672 (N_672,N_408,N_238);
nand U673 (N_673,N_524,N_192);
or U674 (N_674,N_46,N_81);
nor U675 (N_675,N_17,N_66);
nand U676 (N_676,N_558,N_563);
or U677 (N_677,N_468,N_494);
or U678 (N_678,N_54,N_431);
or U679 (N_679,N_384,N_285);
or U680 (N_680,N_32,N_466);
nor U681 (N_681,N_387,N_39);
nor U682 (N_682,N_267,N_322);
or U683 (N_683,N_207,N_248);
or U684 (N_684,N_202,N_271);
and U685 (N_685,N_216,N_506);
nand U686 (N_686,N_599,N_70);
or U687 (N_687,N_251,N_367);
nand U688 (N_688,N_509,N_206);
or U689 (N_689,N_451,N_526);
nor U690 (N_690,N_21,N_260);
nand U691 (N_691,N_160,N_355);
and U692 (N_692,N_111,N_87);
and U693 (N_693,N_307,N_464);
or U694 (N_694,N_470,N_306);
or U695 (N_695,N_195,N_518);
nor U696 (N_696,N_496,N_49);
or U697 (N_697,N_279,N_378);
nor U698 (N_698,N_409,N_386);
nor U699 (N_699,N_93,N_16);
and U700 (N_700,N_573,N_165);
or U701 (N_701,N_110,N_97);
nand U702 (N_702,N_153,N_281);
nand U703 (N_703,N_566,N_374);
or U704 (N_704,N_244,N_26);
nor U705 (N_705,N_328,N_429);
or U706 (N_706,N_163,N_83);
nor U707 (N_707,N_320,N_341);
nand U708 (N_708,N_231,N_172);
or U709 (N_709,N_457,N_575);
or U710 (N_710,N_208,N_155);
or U711 (N_711,N_415,N_398);
nand U712 (N_712,N_535,N_73);
and U713 (N_713,N_37,N_91);
or U714 (N_714,N_211,N_139);
and U715 (N_715,N_52,N_463);
or U716 (N_716,N_257,N_376);
and U717 (N_717,N_69,N_1);
nor U718 (N_718,N_50,N_586);
or U719 (N_719,N_312,N_580);
or U720 (N_720,N_178,N_373);
nand U721 (N_721,N_28,N_43);
nand U722 (N_722,N_298,N_233);
nand U723 (N_723,N_78,N_400);
or U724 (N_724,N_385,N_318);
or U725 (N_725,N_564,N_179);
xor U726 (N_726,N_481,N_532);
nand U727 (N_727,N_465,N_241);
or U728 (N_728,N_327,N_116);
xnor U729 (N_729,N_571,N_55);
or U730 (N_730,N_379,N_541);
nor U731 (N_731,N_143,N_201);
or U732 (N_732,N_480,N_389);
or U733 (N_733,N_317,N_171);
and U734 (N_734,N_516,N_269);
or U735 (N_735,N_0,N_15);
nor U736 (N_736,N_121,N_505);
and U737 (N_737,N_529,N_108);
or U738 (N_738,N_53,N_333);
and U739 (N_739,N_397,N_335);
and U740 (N_740,N_86,N_234);
nand U741 (N_741,N_467,N_547);
nor U742 (N_742,N_151,N_404);
and U743 (N_743,N_98,N_361);
and U744 (N_744,N_499,N_304);
xnor U745 (N_745,N_200,N_182);
and U746 (N_746,N_63,N_530);
and U747 (N_747,N_193,N_25);
nand U748 (N_748,N_75,N_113);
or U749 (N_749,N_194,N_68);
or U750 (N_750,N_107,N_388);
or U751 (N_751,N_162,N_588);
or U752 (N_752,N_62,N_6);
nor U753 (N_753,N_277,N_487);
nor U754 (N_754,N_533,N_36);
nor U755 (N_755,N_65,N_218);
or U756 (N_756,N_242,N_282);
and U757 (N_757,N_272,N_276);
nor U758 (N_758,N_82,N_519);
or U759 (N_759,N_255,N_289);
nor U760 (N_760,N_572,N_337);
nor U761 (N_761,N_292,N_430);
or U762 (N_762,N_261,N_540);
or U763 (N_763,N_503,N_325);
nand U764 (N_764,N_297,N_9);
nand U765 (N_765,N_263,N_287);
nor U766 (N_766,N_539,N_545);
and U767 (N_767,N_498,N_308);
nor U768 (N_768,N_326,N_221);
nor U769 (N_769,N_147,N_423);
nand U770 (N_770,N_99,N_584);
and U771 (N_771,N_565,N_301);
and U772 (N_772,N_256,N_124);
nand U773 (N_773,N_284,N_164);
or U774 (N_774,N_189,N_427);
xor U775 (N_775,N_340,N_311);
and U776 (N_776,N_118,N_490);
or U777 (N_777,N_390,N_112);
xor U778 (N_778,N_595,N_357);
or U779 (N_779,N_174,N_64);
and U780 (N_780,N_444,N_13);
or U781 (N_781,N_462,N_265);
xor U782 (N_782,N_438,N_315);
or U783 (N_783,N_536,N_476);
nor U784 (N_784,N_130,N_294);
nor U785 (N_785,N_578,N_128);
and U786 (N_786,N_72,N_425);
or U787 (N_787,N_426,N_158);
and U788 (N_788,N_119,N_391);
or U789 (N_789,N_246,N_71);
and U790 (N_790,N_227,N_491);
nand U791 (N_791,N_407,N_523);
nand U792 (N_792,N_449,N_167);
nand U793 (N_793,N_266,N_103);
or U794 (N_794,N_38,N_531);
nand U795 (N_795,N_345,N_168);
and U796 (N_796,N_537,N_336);
and U797 (N_797,N_454,N_383);
nor U798 (N_798,N_508,N_101);
or U799 (N_799,N_359,N_262);
nand U800 (N_800,N_258,N_41);
nand U801 (N_801,N_370,N_126);
nor U802 (N_802,N_472,N_369);
or U803 (N_803,N_554,N_477);
and U804 (N_804,N_236,N_528);
and U805 (N_805,N_142,N_401);
nand U806 (N_806,N_122,N_587);
nor U807 (N_807,N_94,N_568);
nor U808 (N_808,N_173,N_346);
nand U809 (N_809,N_14,N_377);
and U810 (N_810,N_243,N_138);
nor U811 (N_811,N_264,N_35);
and U812 (N_812,N_290,N_34);
xor U813 (N_813,N_104,N_314);
and U814 (N_814,N_89,N_166);
nand U815 (N_815,N_190,N_574);
or U816 (N_816,N_120,N_125);
and U817 (N_817,N_109,N_482);
and U818 (N_818,N_92,N_80);
nor U819 (N_819,N_593,N_394);
nand U820 (N_820,N_517,N_18);
or U821 (N_821,N_253,N_31);
nand U822 (N_822,N_217,N_11);
nand U823 (N_823,N_371,N_224);
and U824 (N_824,N_403,N_250);
nand U825 (N_825,N_495,N_582);
nand U826 (N_826,N_488,N_33);
or U827 (N_827,N_299,N_181);
nor U828 (N_828,N_48,N_344);
nor U829 (N_829,N_79,N_40);
nor U830 (N_830,N_76,N_520);
and U831 (N_831,N_309,N_313);
and U832 (N_832,N_459,N_510);
and U833 (N_833,N_131,N_441);
or U834 (N_834,N_157,N_239);
or U835 (N_835,N_310,N_84);
or U836 (N_836,N_140,N_442);
nor U837 (N_837,N_324,N_413);
nor U838 (N_838,N_12,N_175);
nand U839 (N_839,N_170,N_596);
and U840 (N_840,N_522,N_534);
or U841 (N_841,N_416,N_252);
nand U842 (N_842,N_136,N_569);
and U843 (N_843,N_319,N_57);
nand U844 (N_844,N_330,N_579);
nand U845 (N_845,N_577,N_550);
nor U846 (N_846,N_226,N_177);
nand U847 (N_847,N_402,N_392);
nor U848 (N_848,N_10,N_417);
or U849 (N_849,N_428,N_95);
or U850 (N_850,N_286,N_365);
nor U851 (N_851,N_149,N_557);
nor U852 (N_852,N_473,N_424);
or U853 (N_853,N_186,N_148);
or U854 (N_854,N_204,N_114);
nand U855 (N_855,N_448,N_133);
and U856 (N_856,N_405,N_585);
nand U857 (N_857,N_591,N_210);
nand U858 (N_858,N_123,N_504);
nand U859 (N_859,N_225,N_77);
nor U860 (N_860,N_363,N_443);
and U861 (N_861,N_544,N_446);
nand U862 (N_862,N_561,N_497);
or U863 (N_863,N_471,N_212);
and U864 (N_864,N_559,N_419);
nand U865 (N_865,N_30,N_411);
or U866 (N_866,N_19,N_590);
or U867 (N_867,N_380,N_342);
or U868 (N_868,N_115,N_259);
nor U869 (N_869,N_254,N_96);
or U870 (N_870,N_515,N_296);
or U871 (N_871,N_594,N_507);
and U872 (N_872,N_23,N_60);
or U873 (N_873,N_347,N_418);
or U874 (N_874,N_549,N_489);
or U875 (N_875,N_59,N_303);
nand U876 (N_876,N_240,N_3);
xnor U877 (N_877,N_154,N_543);
nor U878 (N_878,N_399,N_360);
or U879 (N_879,N_213,N_440);
nand U880 (N_880,N_222,N_479);
nand U881 (N_881,N_501,N_141);
and U882 (N_882,N_485,N_274);
nand U883 (N_883,N_198,N_478);
or U884 (N_884,N_185,N_24);
nand U885 (N_885,N_422,N_589);
nor U886 (N_886,N_414,N_61);
nand U887 (N_887,N_334,N_74);
nor U888 (N_888,N_521,N_362);
and U889 (N_889,N_548,N_552);
nand U890 (N_890,N_597,N_295);
nand U891 (N_891,N_453,N_445);
or U892 (N_892,N_8,N_146);
or U893 (N_893,N_88,N_500);
nand U894 (N_894,N_486,N_514);
nor U895 (N_895,N_105,N_436);
nand U896 (N_896,N_329,N_395);
or U897 (N_897,N_511,N_474);
and U898 (N_898,N_209,N_58);
nor U899 (N_899,N_47,N_551);
and U900 (N_900,N_86,N_28);
nand U901 (N_901,N_525,N_239);
nor U902 (N_902,N_374,N_494);
and U903 (N_903,N_541,N_255);
nand U904 (N_904,N_333,N_519);
nor U905 (N_905,N_592,N_56);
and U906 (N_906,N_479,N_8);
or U907 (N_907,N_568,N_514);
nand U908 (N_908,N_22,N_146);
or U909 (N_909,N_280,N_62);
or U910 (N_910,N_125,N_161);
nor U911 (N_911,N_418,N_401);
and U912 (N_912,N_278,N_40);
and U913 (N_913,N_178,N_341);
nor U914 (N_914,N_64,N_139);
nand U915 (N_915,N_478,N_515);
and U916 (N_916,N_426,N_45);
or U917 (N_917,N_284,N_547);
nand U918 (N_918,N_231,N_310);
or U919 (N_919,N_549,N_207);
nand U920 (N_920,N_7,N_133);
nor U921 (N_921,N_398,N_513);
or U922 (N_922,N_44,N_440);
nor U923 (N_923,N_138,N_261);
nor U924 (N_924,N_333,N_32);
nor U925 (N_925,N_90,N_552);
nand U926 (N_926,N_420,N_500);
nand U927 (N_927,N_89,N_10);
or U928 (N_928,N_439,N_551);
nor U929 (N_929,N_106,N_39);
or U930 (N_930,N_107,N_482);
and U931 (N_931,N_334,N_539);
nand U932 (N_932,N_265,N_42);
nor U933 (N_933,N_128,N_412);
and U934 (N_934,N_172,N_363);
or U935 (N_935,N_85,N_300);
nor U936 (N_936,N_209,N_507);
or U937 (N_937,N_341,N_51);
or U938 (N_938,N_186,N_483);
or U939 (N_939,N_307,N_462);
and U940 (N_940,N_22,N_160);
and U941 (N_941,N_486,N_425);
or U942 (N_942,N_466,N_391);
and U943 (N_943,N_198,N_560);
or U944 (N_944,N_66,N_370);
xor U945 (N_945,N_472,N_291);
nor U946 (N_946,N_106,N_573);
nand U947 (N_947,N_243,N_69);
or U948 (N_948,N_264,N_178);
nor U949 (N_949,N_236,N_479);
nand U950 (N_950,N_4,N_130);
and U951 (N_951,N_145,N_113);
nor U952 (N_952,N_527,N_534);
nor U953 (N_953,N_286,N_108);
or U954 (N_954,N_235,N_300);
nor U955 (N_955,N_256,N_401);
nand U956 (N_956,N_479,N_434);
nand U957 (N_957,N_503,N_568);
nor U958 (N_958,N_115,N_505);
nand U959 (N_959,N_344,N_343);
nand U960 (N_960,N_248,N_599);
nand U961 (N_961,N_67,N_373);
and U962 (N_962,N_247,N_351);
and U963 (N_963,N_15,N_477);
or U964 (N_964,N_147,N_471);
or U965 (N_965,N_462,N_584);
and U966 (N_966,N_15,N_237);
or U967 (N_967,N_29,N_554);
nand U968 (N_968,N_199,N_588);
or U969 (N_969,N_475,N_51);
nor U970 (N_970,N_17,N_304);
and U971 (N_971,N_209,N_123);
and U972 (N_972,N_534,N_453);
nor U973 (N_973,N_256,N_391);
or U974 (N_974,N_243,N_49);
nand U975 (N_975,N_92,N_277);
nand U976 (N_976,N_77,N_427);
nand U977 (N_977,N_405,N_460);
or U978 (N_978,N_3,N_266);
and U979 (N_979,N_339,N_60);
nand U980 (N_980,N_400,N_129);
nand U981 (N_981,N_125,N_404);
nand U982 (N_982,N_110,N_565);
or U983 (N_983,N_441,N_216);
or U984 (N_984,N_4,N_469);
nor U985 (N_985,N_333,N_75);
nand U986 (N_986,N_487,N_128);
or U987 (N_987,N_343,N_510);
or U988 (N_988,N_368,N_425);
or U989 (N_989,N_111,N_447);
nor U990 (N_990,N_518,N_558);
nor U991 (N_991,N_490,N_336);
and U992 (N_992,N_336,N_237);
nor U993 (N_993,N_59,N_187);
or U994 (N_994,N_551,N_240);
or U995 (N_995,N_107,N_339);
nand U996 (N_996,N_187,N_312);
or U997 (N_997,N_323,N_328);
nand U998 (N_998,N_560,N_189);
and U999 (N_999,N_144,N_428);
or U1000 (N_1000,N_337,N_470);
nor U1001 (N_1001,N_268,N_300);
nor U1002 (N_1002,N_542,N_355);
nand U1003 (N_1003,N_487,N_521);
nor U1004 (N_1004,N_549,N_284);
and U1005 (N_1005,N_255,N_374);
nor U1006 (N_1006,N_314,N_460);
nand U1007 (N_1007,N_177,N_153);
or U1008 (N_1008,N_504,N_448);
or U1009 (N_1009,N_243,N_181);
or U1010 (N_1010,N_562,N_161);
nor U1011 (N_1011,N_301,N_87);
and U1012 (N_1012,N_398,N_50);
or U1013 (N_1013,N_344,N_260);
and U1014 (N_1014,N_118,N_217);
or U1015 (N_1015,N_165,N_83);
nand U1016 (N_1016,N_240,N_334);
or U1017 (N_1017,N_292,N_301);
and U1018 (N_1018,N_4,N_18);
and U1019 (N_1019,N_331,N_427);
nor U1020 (N_1020,N_67,N_361);
nand U1021 (N_1021,N_75,N_220);
nand U1022 (N_1022,N_203,N_217);
nand U1023 (N_1023,N_580,N_419);
or U1024 (N_1024,N_163,N_424);
and U1025 (N_1025,N_439,N_32);
and U1026 (N_1026,N_60,N_299);
or U1027 (N_1027,N_369,N_19);
and U1028 (N_1028,N_396,N_384);
nand U1029 (N_1029,N_429,N_312);
nor U1030 (N_1030,N_593,N_300);
nor U1031 (N_1031,N_340,N_342);
or U1032 (N_1032,N_351,N_28);
or U1033 (N_1033,N_149,N_246);
or U1034 (N_1034,N_400,N_160);
nor U1035 (N_1035,N_540,N_79);
nor U1036 (N_1036,N_40,N_372);
or U1037 (N_1037,N_390,N_370);
or U1038 (N_1038,N_550,N_166);
and U1039 (N_1039,N_199,N_526);
nor U1040 (N_1040,N_415,N_583);
nand U1041 (N_1041,N_523,N_493);
and U1042 (N_1042,N_369,N_21);
and U1043 (N_1043,N_145,N_213);
and U1044 (N_1044,N_203,N_109);
nor U1045 (N_1045,N_69,N_330);
and U1046 (N_1046,N_186,N_400);
nand U1047 (N_1047,N_93,N_561);
and U1048 (N_1048,N_446,N_103);
nand U1049 (N_1049,N_480,N_237);
or U1050 (N_1050,N_71,N_128);
nor U1051 (N_1051,N_397,N_34);
or U1052 (N_1052,N_142,N_387);
and U1053 (N_1053,N_375,N_411);
and U1054 (N_1054,N_177,N_137);
and U1055 (N_1055,N_586,N_245);
nor U1056 (N_1056,N_540,N_479);
and U1057 (N_1057,N_500,N_12);
and U1058 (N_1058,N_222,N_247);
or U1059 (N_1059,N_12,N_577);
or U1060 (N_1060,N_237,N_515);
or U1061 (N_1061,N_451,N_389);
nor U1062 (N_1062,N_62,N_111);
nor U1063 (N_1063,N_541,N_188);
nand U1064 (N_1064,N_280,N_82);
and U1065 (N_1065,N_131,N_310);
or U1066 (N_1066,N_41,N_591);
and U1067 (N_1067,N_163,N_223);
nand U1068 (N_1068,N_332,N_17);
or U1069 (N_1069,N_575,N_19);
or U1070 (N_1070,N_198,N_505);
nand U1071 (N_1071,N_109,N_270);
nand U1072 (N_1072,N_76,N_487);
nor U1073 (N_1073,N_402,N_260);
or U1074 (N_1074,N_264,N_390);
nand U1075 (N_1075,N_247,N_395);
or U1076 (N_1076,N_332,N_250);
or U1077 (N_1077,N_142,N_279);
nand U1078 (N_1078,N_314,N_577);
and U1079 (N_1079,N_284,N_158);
and U1080 (N_1080,N_323,N_367);
xor U1081 (N_1081,N_3,N_46);
and U1082 (N_1082,N_19,N_453);
nand U1083 (N_1083,N_77,N_162);
or U1084 (N_1084,N_538,N_341);
nand U1085 (N_1085,N_563,N_246);
nor U1086 (N_1086,N_330,N_238);
nand U1087 (N_1087,N_501,N_335);
nand U1088 (N_1088,N_530,N_592);
nor U1089 (N_1089,N_554,N_320);
and U1090 (N_1090,N_261,N_244);
nand U1091 (N_1091,N_532,N_588);
and U1092 (N_1092,N_303,N_112);
and U1093 (N_1093,N_266,N_367);
nor U1094 (N_1094,N_282,N_346);
xnor U1095 (N_1095,N_0,N_536);
and U1096 (N_1096,N_359,N_582);
nand U1097 (N_1097,N_66,N_537);
and U1098 (N_1098,N_63,N_136);
nor U1099 (N_1099,N_581,N_407);
nand U1100 (N_1100,N_84,N_494);
nor U1101 (N_1101,N_391,N_75);
and U1102 (N_1102,N_40,N_386);
or U1103 (N_1103,N_58,N_426);
nand U1104 (N_1104,N_302,N_353);
nand U1105 (N_1105,N_133,N_214);
nor U1106 (N_1106,N_566,N_403);
and U1107 (N_1107,N_181,N_263);
nor U1108 (N_1108,N_508,N_161);
nand U1109 (N_1109,N_536,N_528);
and U1110 (N_1110,N_265,N_398);
or U1111 (N_1111,N_221,N_293);
nand U1112 (N_1112,N_218,N_95);
xnor U1113 (N_1113,N_50,N_509);
nor U1114 (N_1114,N_546,N_32);
nor U1115 (N_1115,N_363,N_497);
and U1116 (N_1116,N_278,N_381);
nor U1117 (N_1117,N_331,N_222);
nand U1118 (N_1118,N_354,N_529);
nand U1119 (N_1119,N_329,N_437);
nor U1120 (N_1120,N_43,N_353);
and U1121 (N_1121,N_276,N_158);
or U1122 (N_1122,N_316,N_253);
nand U1123 (N_1123,N_361,N_431);
or U1124 (N_1124,N_176,N_493);
nand U1125 (N_1125,N_79,N_310);
nor U1126 (N_1126,N_420,N_8);
and U1127 (N_1127,N_161,N_313);
xor U1128 (N_1128,N_11,N_361);
and U1129 (N_1129,N_371,N_482);
and U1130 (N_1130,N_111,N_527);
nand U1131 (N_1131,N_396,N_98);
or U1132 (N_1132,N_453,N_314);
nor U1133 (N_1133,N_551,N_123);
or U1134 (N_1134,N_535,N_275);
nand U1135 (N_1135,N_476,N_419);
nand U1136 (N_1136,N_3,N_7);
and U1137 (N_1137,N_527,N_280);
nand U1138 (N_1138,N_170,N_250);
nor U1139 (N_1139,N_272,N_416);
and U1140 (N_1140,N_138,N_439);
xor U1141 (N_1141,N_344,N_112);
and U1142 (N_1142,N_133,N_172);
nand U1143 (N_1143,N_40,N_136);
or U1144 (N_1144,N_369,N_228);
or U1145 (N_1145,N_368,N_52);
or U1146 (N_1146,N_427,N_595);
xor U1147 (N_1147,N_94,N_187);
nor U1148 (N_1148,N_327,N_170);
and U1149 (N_1149,N_242,N_487);
nand U1150 (N_1150,N_231,N_428);
nand U1151 (N_1151,N_327,N_424);
nand U1152 (N_1152,N_469,N_380);
nand U1153 (N_1153,N_114,N_435);
nand U1154 (N_1154,N_224,N_568);
nand U1155 (N_1155,N_506,N_127);
nor U1156 (N_1156,N_233,N_339);
nand U1157 (N_1157,N_4,N_508);
nor U1158 (N_1158,N_363,N_426);
nor U1159 (N_1159,N_506,N_33);
nor U1160 (N_1160,N_237,N_315);
nor U1161 (N_1161,N_373,N_63);
nor U1162 (N_1162,N_491,N_108);
and U1163 (N_1163,N_385,N_538);
or U1164 (N_1164,N_334,N_388);
nor U1165 (N_1165,N_478,N_60);
and U1166 (N_1166,N_374,N_546);
and U1167 (N_1167,N_1,N_429);
nor U1168 (N_1168,N_53,N_401);
nand U1169 (N_1169,N_227,N_301);
nor U1170 (N_1170,N_406,N_53);
nor U1171 (N_1171,N_443,N_156);
nand U1172 (N_1172,N_298,N_387);
nand U1173 (N_1173,N_120,N_0);
or U1174 (N_1174,N_305,N_506);
nor U1175 (N_1175,N_529,N_278);
or U1176 (N_1176,N_144,N_427);
or U1177 (N_1177,N_443,N_254);
nor U1178 (N_1178,N_243,N_35);
or U1179 (N_1179,N_571,N_280);
nor U1180 (N_1180,N_166,N_590);
and U1181 (N_1181,N_265,N_228);
and U1182 (N_1182,N_191,N_84);
nand U1183 (N_1183,N_125,N_128);
nand U1184 (N_1184,N_379,N_234);
nor U1185 (N_1185,N_189,N_216);
and U1186 (N_1186,N_328,N_108);
nor U1187 (N_1187,N_69,N_208);
and U1188 (N_1188,N_339,N_454);
and U1189 (N_1189,N_286,N_23);
nor U1190 (N_1190,N_236,N_7);
nor U1191 (N_1191,N_325,N_431);
nand U1192 (N_1192,N_93,N_228);
and U1193 (N_1193,N_252,N_574);
nand U1194 (N_1194,N_61,N_513);
nand U1195 (N_1195,N_59,N_8);
or U1196 (N_1196,N_344,N_171);
or U1197 (N_1197,N_28,N_122);
or U1198 (N_1198,N_246,N_307);
and U1199 (N_1199,N_584,N_284);
or U1200 (N_1200,N_847,N_615);
nor U1201 (N_1201,N_1145,N_950);
and U1202 (N_1202,N_833,N_1012);
or U1203 (N_1203,N_620,N_744);
or U1204 (N_1204,N_1175,N_802);
and U1205 (N_1205,N_875,N_1182);
nor U1206 (N_1206,N_1162,N_1071);
and U1207 (N_1207,N_693,N_1160);
and U1208 (N_1208,N_708,N_716);
nand U1209 (N_1209,N_777,N_640);
nand U1210 (N_1210,N_688,N_961);
nand U1211 (N_1211,N_857,N_686);
nor U1212 (N_1212,N_1110,N_932);
or U1213 (N_1213,N_779,N_1049);
and U1214 (N_1214,N_1191,N_763);
and U1215 (N_1215,N_1031,N_1136);
nor U1216 (N_1216,N_846,N_1089);
and U1217 (N_1217,N_772,N_879);
nand U1218 (N_1218,N_1181,N_634);
and U1219 (N_1219,N_965,N_800);
and U1220 (N_1220,N_667,N_743);
nand U1221 (N_1221,N_1074,N_751);
and U1222 (N_1222,N_1015,N_909);
nor U1223 (N_1223,N_1114,N_1156);
nand U1224 (N_1224,N_788,N_1135);
or U1225 (N_1225,N_889,N_608);
nand U1226 (N_1226,N_741,N_982);
and U1227 (N_1227,N_1163,N_997);
nor U1228 (N_1228,N_639,N_1142);
and U1229 (N_1229,N_930,N_1034);
and U1230 (N_1230,N_881,N_709);
or U1231 (N_1231,N_918,N_643);
or U1232 (N_1232,N_759,N_995);
and U1233 (N_1233,N_1146,N_1102);
and U1234 (N_1234,N_765,N_869);
nor U1235 (N_1235,N_1047,N_1189);
or U1236 (N_1236,N_949,N_1024);
or U1237 (N_1237,N_897,N_1129);
or U1238 (N_1238,N_1178,N_905);
nor U1239 (N_1239,N_929,N_1121);
nand U1240 (N_1240,N_975,N_764);
nand U1241 (N_1241,N_633,N_618);
or U1242 (N_1242,N_637,N_753);
nor U1243 (N_1243,N_660,N_1143);
or U1244 (N_1244,N_818,N_960);
or U1245 (N_1245,N_1072,N_796);
nand U1246 (N_1246,N_670,N_648);
or U1247 (N_1247,N_1151,N_1009);
xnor U1248 (N_1248,N_1184,N_669);
nor U1249 (N_1249,N_1067,N_609);
or U1250 (N_1250,N_725,N_941);
nor U1251 (N_1251,N_1075,N_801);
or U1252 (N_1252,N_668,N_737);
and U1253 (N_1253,N_919,N_962);
nand U1254 (N_1254,N_821,N_1010);
or U1255 (N_1255,N_998,N_1101);
and U1256 (N_1256,N_845,N_673);
and U1257 (N_1257,N_735,N_601);
or U1258 (N_1258,N_1176,N_1123);
or U1259 (N_1259,N_815,N_679);
xor U1260 (N_1260,N_956,N_1007);
or U1261 (N_1261,N_1043,N_1056);
nor U1262 (N_1262,N_701,N_1016);
nand U1263 (N_1263,N_825,N_641);
or U1264 (N_1264,N_694,N_1134);
nor U1265 (N_1265,N_1157,N_646);
nor U1266 (N_1266,N_936,N_1005);
or U1267 (N_1267,N_1126,N_642);
and U1268 (N_1268,N_899,N_1173);
and U1269 (N_1269,N_692,N_682);
or U1270 (N_1270,N_614,N_1088);
or U1271 (N_1271,N_1138,N_698);
nor U1272 (N_1272,N_964,N_856);
nand U1273 (N_1273,N_795,N_671);
nor U1274 (N_1274,N_872,N_662);
nand U1275 (N_1275,N_1158,N_1168);
or U1276 (N_1276,N_977,N_848);
xnor U1277 (N_1277,N_697,N_798);
or U1278 (N_1278,N_675,N_696);
nor U1279 (N_1279,N_749,N_830);
xor U1280 (N_1280,N_858,N_923);
nor U1281 (N_1281,N_602,N_810);
or U1282 (N_1282,N_1028,N_1164);
or U1283 (N_1283,N_989,N_702);
and U1284 (N_1284,N_834,N_1108);
nand U1285 (N_1285,N_650,N_736);
nor U1286 (N_1286,N_914,N_987);
or U1287 (N_1287,N_1058,N_611);
and U1288 (N_1288,N_750,N_1018);
or U1289 (N_1289,N_854,N_984);
nor U1290 (N_1290,N_863,N_728);
nor U1291 (N_1291,N_659,N_937);
nand U1292 (N_1292,N_1020,N_680);
nand U1293 (N_1293,N_958,N_1100);
nor U1294 (N_1294,N_717,N_1127);
and U1295 (N_1295,N_1055,N_672);
nand U1296 (N_1296,N_1045,N_775);
nand U1297 (N_1297,N_1147,N_877);
or U1298 (N_1298,N_771,N_1172);
nor U1299 (N_1299,N_840,N_1004);
nand U1300 (N_1300,N_665,N_747);
nor U1301 (N_1301,N_631,N_839);
nand U1302 (N_1302,N_769,N_1011);
and U1303 (N_1303,N_957,N_742);
nand U1304 (N_1304,N_985,N_707);
nor U1305 (N_1305,N_619,N_819);
or U1306 (N_1306,N_1090,N_946);
and U1307 (N_1307,N_980,N_1065);
or U1308 (N_1308,N_884,N_954);
nor U1309 (N_1309,N_603,N_868);
or U1310 (N_1310,N_811,N_862);
nand U1311 (N_1311,N_1079,N_1023);
and U1312 (N_1312,N_939,N_865);
nor U1313 (N_1313,N_920,N_774);
or U1314 (N_1314,N_1060,N_625);
nor U1315 (N_1315,N_621,N_1053);
nor U1316 (N_1316,N_647,N_663);
nor U1317 (N_1317,N_836,N_778);
nand U1318 (N_1318,N_921,N_1017);
nand U1319 (N_1319,N_773,N_922);
and U1320 (N_1320,N_1073,N_974);
and U1321 (N_1321,N_1064,N_1022);
nor U1322 (N_1322,N_767,N_824);
nand U1323 (N_1323,N_1150,N_970);
and U1324 (N_1324,N_1041,N_666);
or U1325 (N_1325,N_1052,N_683);
nor U1326 (N_1326,N_651,N_789);
nand U1327 (N_1327,N_695,N_1001);
nand U1328 (N_1328,N_803,N_1077);
nor U1329 (N_1329,N_1084,N_734);
or U1330 (N_1330,N_842,N_674);
and U1331 (N_1331,N_1054,N_1167);
nor U1332 (N_1332,N_691,N_808);
nor U1333 (N_1333,N_1046,N_1094);
nand U1334 (N_1334,N_664,N_657);
nand U1335 (N_1335,N_953,N_902);
nor U1336 (N_1336,N_757,N_1161);
nor U1337 (N_1337,N_947,N_927);
and U1338 (N_1338,N_952,N_1044);
or U1339 (N_1339,N_1186,N_951);
or U1340 (N_1340,N_644,N_1170);
xor U1341 (N_1341,N_807,N_782);
and U1342 (N_1342,N_917,N_820);
nor U1343 (N_1343,N_645,N_726);
or U1344 (N_1344,N_1042,N_955);
nand U1345 (N_1345,N_829,N_607);
and U1346 (N_1346,N_901,N_762);
nand U1347 (N_1347,N_624,N_786);
and U1348 (N_1348,N_988,N_745);
or U1349 (N_1349,N_999,N_1149);
nor U1350 (N_1350,N_1137,N_677);
or U1351 (N_1351,N_1139,N_1125);
nand U1352 (N_1352,N_963,N_935);
or U1353 (N_1353,N_604,N_652);
nor U1354 (N_1354,N_1083,N_1116);
or U1355 (N_1355,N_658,N_1154);
and U1356 (N_1356,N_1196,N_738);
nor U1357 (N_1357,N_1197,N_1014);
and U1358 (N_1358,N_752,N_1050);
and U1359 (N_1359,N_990,N_851);
nand U1360 (N_1360,N_853,N_703);
and U1361 (N_1361,N_996,N_895);
or U1362 (N_1362,N_1119,N_712);
nor U1363 (N_1363,N_866,N_860);
nand U1364 (N_1364,N_1174,N_785);
nand U1365 (N_1365,N_632,N_908);
nand U1366 (N_1366,N_770,N_841);
nor U1367 (N_1367,N_979,N_635);
and U1368 (N_1368,N_859,N_1026);
nand U1369 (N_1369,N_661,N_969);
and U1370 (N_1370,N_993,N_885);
nand U1371 (N_1371,N_740,N_1159);
nand U1372 (N_1372,N_1033,N_791);
or U1373 (N_1373,N_1166,N_1025);
or U1374 (N_1374,N_893,N_783);
nor U1375 (N_1375,N_1029,N_813);
nand U1376 (N_1376,N_1006,N_915);
or U1377 (N_1377,N_718,N_1117);
nor U1378 (N_1378,N_1098,N_1068);
nand U1379 (N_1379,N_911,N_1070);
or U1380 (N_1380,N_1027,N_887);
nor U1381 (N_1381,N_781,N_681);
and U1382 (N_1382,N_715,N_852);
nand U1383 (N_1383,N_934,N_940);
nor U1384 (N_1384,N_727,N_1037);
nor U1385 (N_1385,N_746,N_687);
or U1386 (N_1386,N_699,N_713);
or U1387 (N_1387,N_1019,N_1144);
or U1388 (N_1388,N_616,N_896);
nand U1389 (N_1389,N_684,N_722);
and U1390 (N_1390,N_711,N_766);
and U1391 (N_1391,N_823,N_1133);
nor U1392 (N_1392,N_705,N_827);
and U1393 (N_1393,N_627,N_861);
nor U1394 (N_1394,N_1085,N_855);
nand U1395 (N_1395,N_1193,N_689);
and U1396 (N_1396,N_799,N_912);
and U1397 (N_1397,N_1192,N_916);
nor U1398 (N_1398,N_1030,N_933);
and U1399 (N_1399,N_761,N_622);
and U1400 (N_1400,N_882,N_924);
nand U1401 (N_1401,N_828,N_1097);
nor U1402 (N_1402,N_1120,N_809);
or U1403 (N_1403,N_638,N_739);
nand U1404 (N_1404,N_864,N_867);
nor U1405 (N_1405,N_1051,N_938);
or U1406 (N_1406,N_606,N_1148);
nand U1407 (N_1407,N_886,N_948);
nand U1408 (N_1408,N_878,N_690);
xnor U1409 (N_1409,N_629,N_1187);
nand U1410 (N_1410,N_1128,N_758);
or U1411 (N_1411,N_1171,N_613);
nand U1412 (N_1412,N_655,N_653);
and U1413 (N_1413,N_967,N_838);
nor U1414 (N_1414,N_906,N_760);
nor U1415 (N_1415,N_1008,N_731);
and U1416 (N_1416,N_826,N_943);
or U1417 (N_1417,N_844,N_1131);
or U1418 (N_1418,N_700,N_733);
or U1419 (N_1419,N_1087,N_843);
nor U1420 (N_1420,N_1081,N_626);
and U1421 (N_1421,N_732,N_630);
nand U1422 (N_1422,N_776,N_971);
or U1423 (N_1423,N_1057,N_1066);
and U1424 (N_1424,N_900,N_623);
nand U1425 (N_1425,N_817,N_794);
xor U1426 (N_1426,N_1190,N_1076);
nand U1427 (N_1427,N_972,N_1132);
or U1428 (N_1428,N_1111,N_724);
or U1429 (N_1429,N_873,N_925);
and U1430 (N_1430,N_1059,N_835);
nor U1431 (N_1431,N_636,N_1032);
or U1432 (N_1432,N_1118,N_892);
nand U1433 (N_1433,N_628,N_1105);
and U1434 (N_1434,N_710,N_805);
and U1435 (N_1435,N_1183,N_1106);
nand U1436 (N_1436,N_942,N_994);
xnor U1437 (N_1437,N_1115,N_730);
and U1438 (N_1438,N_1099,N_704);
nand U1439 (N_1439,N_1096,N_928);
and U1440 (N_1440,N_1122,N_814);
and U1441 (N_1441,N_1091,N_1038);
or U1442 (N_1442,N_903,N_1194);
nand U1443 (N_1443,N_822,N_1104);
nand U1444 (N_1444,N_685,N_1130);
or U1445 (N_1445,N_1141,N_832);
nand U1446 (N_1446,N_610,N_656);
nand U1447 (N_1447,N_978,N_748);
nand U1448 (N_1448,N_991,N_1080);
and U1449 (N_1449,N_1152,N_1155);
and U1450 (N_1450,N_874,N_812);
or U1451 (N_1451,N_1112,N_1185);
or U1452 (N_1452,N_1095,N_973);
and U1453 (N_1453,N_816,N_756);
or U1454 (N_1454,N_676,N_790);
and U1455 (N_1455,N_907,N_890);
or U1456 (N_1456,N_983,N_754);
nand U1457 (N_1457,N_721,N_806);
nand U1458 (N_1458,N_1092,N_1040);
nor U1459 (N_1459,N_976,N_1000);
nand U1460 (N_1460,N_1180,N_1153);
nand U1461 (N_1461,N_1103,N_768);
and U1462 (N_1462,N_755,N_837);
nor U1463 (N_1463,N_1140,N_1002);
and U1464 (N_1464,N_888,N_1165);
or U1465 (N_1465,N_1113,N_1198);
nor U1466 (N_1466,N_931,N_714);
and U1467 (N_1467,N_649,N_1177);
nor U1468 (N_1468,N_617,N_612);
or U1469 (N_1469,N_1199,N_913);
nand U1470 (N_1470,N_1082,N_945);
nand U1471 (N_1471,N_780,N_729);
nor U1472 (N_1472,N_1061,N_883);
and U1473 (N_1473,N_831,N_787);
xor U1474 (N_1474,N_1078,N_1086);
nor U1475 (N_1475,N_1124,N_968);
nand U1476 (N_1476,N_898,N_891);
or U1477 (N_1477,N_966,N_720);
and U1478 (N_1478,N_1048,N_1188);
nand U1479 (N_1479,N_1036,N_1109);
nand U1480 (N_1480,N_1093,N_944);
nor U1481 (N_1481,N_605,N_654);
or U1482 (N_1482,N_1107,N_1003);
nand U1483 (N_1483,N_992,N_793);
or U1484 (N_1484,N_797,N_876);
or U1485 (N_1485,N_871,N_1013);
nor U1486 (N_1486,N_1063,N_894);
and U1487 (N_1487,N_804,N_1062);
nand U1488 (N_1488,N_926,N_981);
nor U1489 (N_1489,N_600,N_723);
or U1490 (N_1490,N_1069,N_850);
and U1491 (N_1491,N_1039,N_986);
nand U1492 (N_1492,N_706,N_784);
and U1493 (N_1493,N_910,N_849);
xor U1494 (N_1494,N_1169,N_719);
nand U1495 (N_1495,N_1035,N_1179);
nand U1496 (N_1496,N_870,N_678);
and U1497 (N_1497,N_904,N_1195);
nor U1498 (N_1498,N_1021,N_959);
and U1499 (N_1499,N_792,N_880);
and U1500 (N_1500,N_1073,N_862);
or U1501 (N_1501,N_686,N_997);
nor U1502 (N_1502,N_853,N_677);
nor U1503 (N_1503,N_619,N_750);
or U1504 (N_1504,N_627,N_716);
or U1505 (N_1505,N_886,N_873);
nor U1506 (N_1506,N_1168,N_718);
xnor U1507 (N_1507,N_1094,N_980);
or U1508 (N_1508,N_1008,N_782);
nand U1509 (N_1509,N_758,N_854);
and U1510 (N_1510,N_1007,N_795);
nand U1511 (N_1511,N_1014,N_958);
or U1512 (N_1512,N_1177,N_658);
nand U1513 (N_1513,N_708,N_673);
nand U1514 (N_1514,N_812,N_663);
and U1515 (N_1515,N_848,N_1029);
nand U1516 (N_1516,N_812,N_1085);
and U1517 (N_1517,N_1127,N_665);
nor U1518 (N_1518,N_1191,N_1125);
and U1519 (N_1519,N_1099,N_792);
or U1520 (N_1520,N_621,N_1160);
nor U1521 (N_1521,N_985,N_926);
nor U1522 (N_1522,N_712,N_1089);
or U1523 (N_1523,N_759,N_733);
nand U1524 (N_1524,N_768,N_642);
or U1525 (N_1525,N_985,N_1101);
nor U1526 (N_1526,N_613,N_1065);
and U1527 (N_1527,N_684,N_1012);
nor U1528 (N_1528,N_1158,N_1040);
nor U1529 (N_1529,N_789,N_675);
or U1530 (N_1530,N_727,N_1133);
or U1531 (N_1531,N_722,N_1127);
xnor U1532 (N_1532,N_942,N_729);
or U1533 (N_1533,N_834,N_787);
and U1534 (N_1534,N_820,N_973);
nand U1535 (N_1535,N_994,N_937);
and U1536 (N_1536,N_712,N_845);
xor U1537 (N_1537,N_1104,N_816);
nand U1538 (N_1538,N_948,N_700);
nor U1539 (N_1539,N_971,N_896);
or U1540 (N_1540,N_763,N_902);
or U1541 (N_1541,N_707,N_845);
and U1542 (N_1542,N_1057,N_1100);
nor U1543 (N_1543,N_620,N_648);
nand U1544 (N_1544,N_1146,N_996);
nor U1545 (N_1545,N_648,N_704);
and U1546 (N_1546,N_1072,N_748);
nor U1547 (N_1547,N_981,N_851);
and U1548 (N_1548,N_804,N_996);
and U1549 (N_1549,N_1014,N_1106);
nand U1550 (N_1550,N_815,N_1054);
xor U1551 (N_1551,N_953,N_1073);
nand U1552 (N_1552,N_971,N_871);
and U1553 (N_1553,N_611,N_919);
nand U1554 (N_1554,N_742,N_1087);
nor U1555 (N_1555,N_1161,N_953);
nor U1556 (N_1556,N_905,N_1037);
or U1557 (N_1557,N_1189,N_805);
and U1558 (N_1558,N_667,N_919);
or U1559 (N_1559,N_938,N_610);
nor U1560 (N_1560,N_680,N_837);
or U1561 (N_1561,N_914,N_900);
or U1562 (N_1562,N_685,N_1016);
nand U1563 (N_1563,N_793,N_906);
nor U1564 (N_1564,N_601,N_653);
or U1565 (N_1565,N_736,N_961);
nand U1566 (N_1566,N_849,N_987);
nand U1567 (N_1567,N_819,N_1048);
nand U1568 (N_1568,N_883,N_621);
nand U1569 (N_1569,N_1174,N_979);
or U1570 (N_1570,N_1001,N_1020);
or U1571 (N_1571,N_1109,N_1057);
or U1572 (N_1572,N_1172,N_604);
nor U1573 (N_1573,N_986,N_1012);
nor U1574 (N_1574,N_1115,N_831);
and U1575 (N_1575,N_759,N_1035);
or U1576 (N_1576,N_989,N_1054);
xnor U1577 (N_1577,N_1089,N_1092);
and U1578 (N_1578,N_1094,N_697);
and U1579 (N_1579,N_1144,N_700);
nor U1580 (N_1580,N_767,N_1152);
nand U1581 (N_1581,N_622,N_637);
or U1582 (N_1582,N_819,N_1132);
nor U1583 (N_1583,N_1137,N_961);
nand U1584 (N_1584,N_1127,N_936);
nand U1585 (N_1585,N_714,N_690);
nor U1586 (N_1586,N_696,N_737);
nand U1587 (N_1587,N_666,N_702);
nor U1588 (N_1588,N_765,N_1116);
nor U1589 (N_1589,N_1027,N_996);
nor U1590 (N_1590,N_976,N_1168);
nor U1591 (N_1591,N_772,N_1079);
and U1592 (N_1592,N_623,N_1093);
nor U1593 (N_1593,N_731,N_1017);
or U1594 (N_1594,N_869,N_1056);
or U1595 (N_1595,N_1037,N_824);
nand U1596 (N_1596,N_979,N_713);
nand U1597 (N_1597,N_746,N_747);
nor U1598 (N_1598,N_648,N_1062);
nand U1599 (N_1599,N_853,N_651);
nand U1600 (N_1600,N_891,N_1115);
or U1601 (N_1601,N_670,N_1082);
nor U1602 (N_1602,N_758,N_1130);
and U1603 (N_1603,N_1166,N_1026);
or U1604 (N_1604,N_733,N_1070);
or U1605 (N_1605,N_1150,N_1172);
nand U1606 (N_1606,N_1053,N_1192);
or U1607 (N_1607,N_978,N_631);
or U1608 (N_1608,N_1052,N_1040);
or U1609 (N_1609,N_953,N_755);
nand U1610 (N_1610,N_1102,N_1025);
nand U1611 (N_1611,N_691,N_856);
or U1612 (N_1612,N_1049,N_1047);
nor U1613 (N_1613,N_1069,N_692);
nand U1614 (N_1614,N_1182,N_974);
nor U1615 (N_1615,N_714,N_739);
or U1616 (N_1616,N_1140,N_912);
or U1617 (N_1617,N_1061,N_634);
or U1618 (N_1618,N_902,N_725);
and U1619 (N_1619,N_1127,N_843);
nor U1620 (N_1620,N_778,N_861);
nand U1621 (N_1621,N_957,N_658);
nor U1622 (N_1622,N_847,N_1123);
nand U1623 (N_1623,N_805,N_1009);
nand U1624 (N_1624,N_1151,N_641);
nand U1625 (N_1625,N_989,N_948);
and U1626 (N_1626,N_718,N_1083);
and U1627 (N_1627,N_798,N_741);
nor U1628 (N_1628,N_723,N_861);
or U1629 (N_1629,N_1140,N_672);
and U1630 (N_1630,N_740,N_650);
and U1631 (N_1631,N_737,N_1061);
nand U1632 (N_1632,N_794,N_812);
and U1633 (N_1633,N_1137,N_1105);
nor U1634 (N_1634,N_1114,N_803);
nor U1635 (N_1635,N_1147,N_829);
and U1636 (N_1636,N_798,N_740);
or U1637 (N_1637,N_874,N_772);
nand U1638 (N_1638,N_1098,N_728);
nor U1639 (N_1639,N_1016,N_707);
and U1640 (N_1640,N_812,N_602);
nand U1641 (N_1641,N_886,N_602);
or U1642 (N_1642,N_1024,N_965);
nand U1643 (N_1643,N_832,N_614);
or U1644 (N_1644,N_1033,N_1065);
or U1645 (N_1645,N_1135,N_1059);
nor U1646 (N_1646,N_699,N_823);
and U1647 (N_1647,N_795,N_1126);
or U1648 (N_1648,N_1160,N_673);
nand U1649 (N_1649,N_922,N_1192);
and U1650 (N_1650,N_902,N_1035);
xor U1651 (N_1651,N_909,N_1183);
and U1652 (N_1652,N_763,N_846);
nand U1653 (N_1653,N_774,N_659);
nor U1654 (N_1654,N_724,N_746);
or U1655 (N_1655,N_1087,N_1148);
and U1656 (N_1656,N_1042,N_870);
nor U1657 (N_1657,N_1147,N_801);
and U1658 (N_1658,N_986,N_1101);
or U1659 (N_1659,N_1072,N_1114);
nor U1660 (N_1660,N_1054,N_653);
nand U1661 (N_1661,N_883,N_878);
nand U1662 (N_1662,N_778,N_637);
or U1663 (N_1663,N_1186,N_862);
nand U1664 (N_1664,N_934,N_1173);
nand U1665 (N_1665,N_1085,N_653);
nor U1666 (N_1666,N_979,N_1181);
nor U1667 (N_1667,N_778,N_1067);
or U1668 (N_1668,N_824,N_815);
nand U1669 (N_1669,N_633,N_1165);
nand U1670 (N_1670,N_1036,N_1104);
and U1671 (N_1671,N_1036,N_1143);
and U1672 (N_1672,N_665,N_805);
nand U1673 (N_1673,N_698,N_1044);
nor U1674 (N_1674,N_1122,N_683);
nand U1675 (N_1675,N_785,N_875);
and U1676 (N_1676,N_1126,N_1195);
nor U1677 (N_1677,N_681,N_1042);
or U1678 (N_1678,N_678,N_805);
or U1679 (N_1679,N_1113,N_1195);
and U1680 (N_1680,N_695,N_804);
nor U1681 (N_1681,N_922,N_932);
nor U1682 (N_1682,N_961,N_801);
or U1683 (N_1683,N_602,N_778);
nand U1684 (N_1684,N_776,N_1055);
or U1685 (N_1685,N_1122,N_635);
or U1686 (N_1686,N_904,N_643);
nor U1687 (N_1687,N_925,N_924);
and U1688 (N_1688,N_1018,N_794);
and U1689 (N_1689,N_839,N_780);
and U1690 (N_1690,N_883,N_1169);
nand U1691 (N_1691,N_657,N_960);
and U1692 (N_1692,N_725,N_1037);
nand U1693 (N_1693,N_1030,N_725);
nand U1694 (N_1694,N_1150,N_753);
nand U1695 (N_1695,N_775,N_817);
nand U1696 (N_1696,N_1193,N_847);
and U1697 (N_1697,N_1082,N_985);
nor U1698 (N_1698,N_735,N_636);
nand U1699 (N_1699,N_854,N_722);
nand U1700 (N_1700,N_760,N_917);
or U1701 (N_1701,N_617,N_837);
or U1702 (N_1702,N_671,N_1089);
nand U1703 (N_1703,N_734,N_770);
nand U1704 (N_1704,N_709,N_778);
nand U1705 (N_1705,N_1104,N_653);
or U1706 (N_1706,N_739,N_692);
nor U1707 (N_1707,N_777,N_661);
and U1708 (N_1708,N_958,N_896);
nand U1709 (N_1709,N_1060,N_985);
nand U1710 (N_1710,N_1087,N_816);
nand U1711 (N_1711,N_1137,N_978);
nand U1712 (N_1712,N_1101,N_842);
and U1713 (N_1713,N_1076,N_692);
nand U1714 (N_1714,N_922,N_1110);
or U1715 (N_1715,N_614,N_1116);
nor U1716 (N_1716,N_652,N_890);
nand U1717 (N_1717,N_685,N_687);
nand U1718 (N_1718,N_913,N_1094);
or U1719 (N_1719,N_800,N_1056);
nor U1720 (N_1720,N_696,N_911);
nand U1721 (N_1721,N_683,N_1094);
or U1722 (N_1722,N_1117,N_1097);
and U1723 (N_1723,N_1189,N_709);
nor U1724 (N_1724,N_900,N_675);
nor U1725 (N_1725,N_921,N_983);
nor U1726 (N_1726,N_1023,N_913);
nand U1727 (N_1727,N_1042,N_1041);
and U1728 (N_1728,N_857,N_607);
or U1729 (N_1729,N_1048,N_1076);
or U1730 (N_1730,N_930,N_772);
or U1731 (N_1731,N_996,N_1133);
or U1732 (N_1732,N_1129,N_753);
and U1733 (N_1733,N_720,N_973);
or U1734 (N_1734,N_808,N_606);
and U1735 (N_1735,N_694,N_678);
or U1736 (N_1736,N_625,N_1035);
nor U1737 (N_1737,N_1196,N_713);
and U1738 (N_1738,N_784,N_916);
nand U1739 (N_1739,N_672,N_627);
or U1740 (N_1740,N_1130,N_1017);
or U1741 (N_1741,N_618,N_1035);
or U1742 (N_1742,N_655,N_1022);
nor U1743 (N_1743,N_760,N_1108);
or U1744 (N_1744,N_1050,N_1153);
nand U1745 (N_1745,N_900,N_851);
nor U1746 (N_1746,N_1047,N_881);
or U1747 (N_1747,N_1199,N_925);
nor U1748 (N_1748,N_1143,N_991);
nand U1749 (N_1749,N_926,N_792);
and U1750 (N_1750,N_787,N_1122);
nand U1751 (N_1751,N_1065,N_1123);
and U1752 (N_1752,N_1188,N_905);
and U1753 (N_1753,N_1059,N_865);
nor U1754 (N_1754,N_1092,N_657);
or U1755 (N_1755,N_1032,N_1050);
or U1756 (N_1756,N_633,N_967);
nand U1757 (N_1757,N_680,N_621);
or U1758 (N_1758,N_1137,N_922);
nor U1759 (N_1759,N_606,N_711);
nand U1760 (N_1760,N_866,N_861);
or U1761 (N_1761,N_1068,N_1063);
and U1762 (N_1762,N_1150,N_1168);
and U1763 (N_1763,N_636,N_1109);
nand U1764 (N_1764,N_824,N_850);
nor U1765 (N_1765,N_761,N_795);
or U1766 (N_1766,N_1100,N_750);
and U1767 (N_1767,N_607,N_1123);
nor U1768 (N_1768,N_612,N_807);
and U1769 (N_1769,N_1069,N_1112);
nand U1770 (N_1770,N_791,N_1162);
or U1771 (N_1771,N_1129,N_703);
and U1772 (N_1772,N_648,N_856);
nand U1773 (N_1773,N_790,N_956);
nand U1774 (N_1774,N_938,N_602);
nor U1775 (N_1775,N_772,N_1106);
nor U1776 (N_1776,N_713,N_1136);
nand U1777 (N_1777,N_904,N_823);
nand U1778 (N_1778,N_909,N_1037);
nor U1779 (N_1779,N_791,N_949);
nor U1780 (N_1780,N_1022,N_826);
or U1781 (N_1781,N_655,N_1042);
nand U1782 (N_1782,N_825,N_687);
xnor U1783 (N_1783,N_1042,N_1189);
nand U1784 (N_1784,N_706,N_936);
and U1785 (N_1785,N_842,N_945);
and U1786 (N_1786,N_1156,N_1148);
or U1787 (N_1787,N_750,N_711);
and U1788 (N_1788,N_909,N_974);
and U1789 (N_1789,N_776,N_707);
and U1790 (N_1790,N_724,N_952);
and U1791 (N_1791,N_710,N_873);
or U1792 (N_1792,N_1189,N_856);
nand U1793 (N_1793,N_1115,N_763);
or U1794 (N_1794,N_846,N_633);
nand U1795 (N_1795,N_1011,N_697);
nand U1796 (N_1796,N_1184,N_1129);
nand U1797 (N_1797,N_834,N_685);
and U1798 (N_1798,N_758,N_805);
nand U1799 (N_1799,N_694,N_875);
nor U1800 (N_1800,N_1635,N_1514);
or U1801 (N_1801,N_1516,N_1474);
and U1802 (N_1802,N_1677,N_1666);
nor U1803 (N_1803,N_1596,N_1362);
nand U1804 (N_1804,N_1374,N_1747);
and U1805 (N_1805,N_1757,N_1429);
nor U1806 (N_1806,N_1608,N_1584);
and U1807 (N_1807,N_1281,N_1390);
nor U1808 (N_1808,N_1606,N_1630);
or U1809 (N_1809,N_1536,N_1479);
nor U1810 (N_1810,N_1716,N_1400);
and U1811 (N_1811,N_1592,N_1741);
and U1812 (N_1812,N_1299,N_1626);
and U1813 (N_1813,N_1709,N_1524);
nor U1814 (N_1814,N_1675,N_1565);
nor U1815 (N_1815,N_1406,N_1334);
nor U1816 (N_1816,N_1331,N_1506);
nor U1817 (N_1817,N_1743,N_1321);
nand U1818 (N_1818,N_1265,N_1577);
nand U1819 (N_1819,N_1733,N_1778);
nand U1820 (N_1820,N_1765,N_1445);
nor U1821 (N_1821,N_1591,N_1650);
and U1822 (N_1822,N_1761,N_1647);
nor U1823 (N_1823,N_1554,N_1328);
and U1824 (N_1824,N_1231,N_1680);
and U1825 (N_1825,N_1367,N_1563);
and U1826 (N_1826,N_1252,N_1251);
and U1827 (N_1827,N_1686,N_1346);
or U1828 (N_1828,N_1360,N_1513);
and U1829 (N_1829,N_1659,N_1684);
nand U1830 (N_1830,N_1269,N_1553);
nor U1831 (N_1831,N_1623,N_1788);
nor U1832 (N_1832,N_1526,N_1758);
nand U1833 (N_1833,N_1419,N_1295);
nand U1834 (N_1834,N_1217,N_1701);
and U1835 (N_1835,N_1639,N_1294);
and U1836 (N_1836,N_1293,N_1545);
nor U1837 (N_1837,N_1466,N_1261);
nor U1838 (N_1838,N_1408,N_1380);
and U1839 (N_1839,N_1570,N_1499);
and U1840 (N_1840,N_1348,N_1273);
nor U1841 (N_1841,N_1493,N_1628);
nor U1842 (N_1842,N_1382,N_1734);
nor U1843 (N_1843,N_1618,N_1468);
nand U1844 (N_1844,N_1679,N_1543);
nand U1845 (N_1845,N_1533,N_1340);
nand U1846 (N_1846,N_1681,N_1388);
nor U1847 (N_1847,N_1462,N_1634);
nand U1848 (N_1848,N_1399,N_1772);
and U1849 (N_1849,N_1483,N_1750);
nand U1850 (N_1850,N_1300,N_1371);
nand U1851 (N_1851,N_1495,N_1222);
nand U1852 (N_1852,N_1256,N_1683);
nor U1853 (N_1853,N_1459,N_1537);
or U1854 (N_1854,N_1724,N_1660);
and U1855 (N_1855,N_1776,N_1455);
nor U1856 (N_1856,N_1310,N_1477);
nand U1857 (N_1857,N_1236,N_1654);
and U1858 (N_1858,N_1664,N_1725);
nor U1859 (N_1859,N_1530,N_1633);
nand U1860 (N_1860,N_1411,N_1768);
nor U1861 (N_1861,N_1327,N_1424);
nand U1862 (N_1862,N_1696,N_1736);
and U1863 (N_1863,N_1214,N_1375);
nor U1864 (N_1864,N_1338,N_1567);
nand U1865 (N_1865,N_1229,N_1753);
nor U1866 (N_1866,N_1700,N_1306);
nor U1867 (N_1867,N_1678,N_1676);
and U1868 (N_1868,N_1731,N_1447);
and U1869 (N_1869,N_1443,N_1763);
or U1870 (N_1870,N_1568,N_1446);
nand U1871 (N_1871,N_1393,N_1485);
nor U1872 (N_1872,N_1385,N_1291);
nor U1873 (N_1873,N_1656,N_1614);
and U1874 (N_1874,N_1494,N_1271);
nand U1875 (N_1875,N_1365,N_1665);
and U1876 (N_1876,N_1314,N_1307);
nor U1877 (N_1877,N_1215,N_1287);
and U1878 (N_1878,N_1378,N_1649);
or U1879 (N_1879,N_1538,N_1586);
nor U1880 (N_1880,N_1397,N_1247);
nand U1881 (N_1881,N_1288,N_1710);
nor U1882 (N_1882,N_1358,N_1442);
or U1883 (N_1883,N_1423,N_1289);
nand U1884 (N_1884,N_1221,N_1320);
and U1885 (N_1885,N_1662,N_1324);
and U1886 (N_1886,N_1430,N_1386);
and U1887 (N_1887,N_1290,N_1744);
nor U1888 (N_1888,N_1519,N_1617);
and U1889 (N_1889,N_1589,N_1283);
nand U1890 (N_1890,N_1775,N_1205);
and U1891 (N_1891,N_1421,N_1632);
and U1892 (N_1892,N_1357,N_1751);
nand U1893 (N_1893,N_1440,N_1735);
nor U1894 (N_1894,N_1489,N_1381);
and U1895 (N_1895,N_1404,N_1540);
and U1896 (N_1896,N_1582,N_1232);
nand U1897 (N_1897,N_1705,N_1488);
nand U1898 (N_1898,N_1450,N_1379);
and U1899 (N_1899,N_1384,N_1790);
and U1900 (N_1900,N_1525,N_1663);
and U1901 (N_1901,N_1597,N_1286);
nor U1902 (N_1902,N_1394,N_1387);
and U1903 (N_1903,N_1746,N_1787);
nand U1904 (N_1904,N_1212,N_1528);
nand U1905 (N_1905,N_1550,N_1789);
nor U1906 (N_1906,N_1651,N_1718);
nand U1907 (N_1907,N_1793,N_1674);
nand U1908 (N_1908,N_1631,N_1250);
nor U1909 (N_1909,N_1764,N_1669);
or U1910 (N_1910,N_1560,N_1267);
nor U1911 (N_1911,N_1282,N_1235);
and U1912 (N_1912,N_1593,N_1501);
and U1913 (N_1913,N_1732,N_1672);
or U1914 (N_1914,N_1574,N_1461);
and U1915 (N_1915,N_1363,N_1691);
nor U1916 (N_1916,N_1227,N_1673);
nand U1917 (N_1917,N_1239,N_1418);
nand U1918 (N_1918,N_1460,N_1552);
or U1919 (N_1919,N_1517,N_1769);
and U1920 (N_1920,N_1425,N_1255);
nand U1921 (N_1921,N_1783,N_1598);
nor U1922 (N_1922,N_1437,N_1264);
and U1923 (N_1923,N_1529,N_1476);
nor U1924 (N_1924,N_1655,N_1512);
and U1925 (N_1925,N_1508,N_1228);
and U1926 (N_1926,N_1211,N_1276);
nor U1927 (N_1927,N_1722,N_1728);
and U1928 (N_1928,N_1708,N_1625);
nor U1929 (N_1929,N_1480,N_1420);
or U1930 (N_1930,N_1376,N_1558);
nand U1931 (N_1931,N_1549,N_1354);
and U1932 (N_1932,N_1760,N_1527);
xor U1933 (N_1933,N_1712,N_1322);
and U1934 (N_1934,N_1595,N_1719);
and U1935 (N_1935,N_1572,N_1458);
nor U1936 (N_1936,N_1329,N_1667);
nand U1937 (N_1937,N_1695,N_1313);
nor U1938 (N_1938,N_1752,N_1481);
nand U1939 (N_1939,N_1469,N_1652);
or U1940 (N_1940,N_1498,N_1260);
and U1941 (N_1941,N_1794,N_1704);
nor U1942 (N_1942,N_1285,N_1453);
and U1943 (N_1943,N_1240,N_1351);
or U1944 (N_1944,N_1610,N_1243);
nand U1945 (N_1945,N_1202,N_1201);
or U1946 (N_1946,N_1770,N_1721);
nor U1947 (N_1947,N_1280,N_1347);
and U1948 (N_1948,N_1796,N_1619);
nand U1949 (N_1949,N_1353,N_1449);
and U1950 (N_1950,N_1636,N_1668);
and U1951 (N_1951,N_1210,N_1755);
or U1952 (N_1952,N_1278,N_1541);
nand U1953 (N_1953,N_1352,N_1244);
and U1954 (N_1954,N_1795,N_1766);
nand U1955 (N_1955,N_1564,N_1531);
and U1956 (N_1956,N_1504,N_1738);
or U1957 (N_1957,N_1219,N_1457);
nand U1958 (N_1958,N_1436,N_1484);
or U1959 (N_1959,N_1274,N_1607);
nand U1960 (N_1960,N_1671,N_1557);
nand U1961 (N_1961,N_1292,N_1642);
nor U1962 (N_1962,N_1792,N_1369);
nor U1963 (N_1963,N_1444,N_1739);
and U1964 (N_1964,N_1412,N_1223);
or U1965 (N_1965,N_1242,N_1599);
nand U1966 (N_1966,N_1409,N_1355);
or U1967 (N_1967,N_1317,N_1767);
nor U1968 (N_1968,N_1629,N_1786);
and U1969 (N_1969,N_1319,N_1697);
or U1970 (N_1970,N_1302,N_1580);
and U1971 (N_1971,N_1467,N_1414);
or U1972 (N_1972,N_1392,N_1262);
nor U1973 (N_1973,N_1784,N_1546);
and U1974 (N_1974,N_1463,N_1534);
and U1975 (N_1975,N_1318,N_1323);
nor U1976 (N_1976,N_1359,N_1218);
nor U1977 (N_1977,N_1435,N_1349);
and U1978 (N_1978,N_1372,N_1699);
xor U1979 (N_1979,N_1366,N_1609);
nand U1980 (N_1980,N_1729,N_1377);
nor U1981 (N_1981,N_1685,N_1601);
xnor U1982 (N_1982,N_1451,N_1491);
or U1983 (N_1983,N_1590,N_1523);
nand U1984 (N_1984,N_1521,N_1316);
nand U1985 (N_1985,N_1270,N_1248);
or U1986 (N_1986,N_1448,N_1658);
nor U1987 (N_1987,N_1566,N_1612);
nor U1988 (N_1988,N_1471,N_1277);
and U1989 (N_1989,N_1233,N_1702);
or U1990 (N_1990,N_1361,N_1643);
nand U1991 (N_1991,N_1613,N_1279);
and U1992 (N_1992,N_1627,N_1326);
and U1993 (N_1993,N_1389,N_1339);
nor U1994 (N_1994,N_1694,N_1470);
and U1995 (N_1995,N_1548,N_1556);
nor U1996 (N_1996,N_1275,N_1620);
or U1997 (N_1997,N_1268,N_1298);
nor U1998 (N_1998,N_1547,N_1333);
nand U1999 (N_1999,N_1723,N_1587);
or U2000 (N_2000,N_1407,N_1226);
or U2001 (N_2001,N_1569,N_1257);
nand U2002 (N_2002,N_1220,N_1422);
or U2003 (N_2003,N_1373,N_1213);
or U2004 (N_2004,N_1416,N_1296);
or U2005 (N_2005,N_1615,N_1748);
nand U2006 (N_2006,N_1308,N_1576);
or U2007 (N_2007,N_1417,N_1798);
or U2008 (N_2008,N_1475,N_1573);
or U2009 (N_2009,N_1454,N_1781);
or U2010 (N_2010,N_1238,N_1797);
nor U2011 (N_2011,N_1234,N_1561);
nor U2012 (N_2012,N_1740,N_1657);
nor U2013 (N_2013,N_1791,N_1337);
nor U2014 (N_2014,N_1237,N_1427);
nand U2015 (N_2015,N_1410,N_1311);
nand U2016 (N_2016,N_1344,N_1544);
and U2017 (N_2017,N_1692,N_1364);
or U2018 (N_2018,N_1602,N_1401);
or U2019 (N_2019,N_1611,N_1759);
or U2020 (N_2020,N_1497,N_1473);
and U2021 (N_2021,N_1403,N_1315);
or U2022 (N_2022,N_1426,N_1581);
or U2023 (N_2023,N_1208,N_1342);
and U2024 (N_2024,N_1532,N_1687);
or U2025 (N_2025,N_1496,N_1490);
and U2026 (N_2026,N_1562,N_1249);
and U2027 (N_2027,N_1774,N_1356);
nor U2028 (N_2028,N_1756,N_1777);
or U2029 (N_2029,N_1713,N_1452);
or U2030 (N_2030,N_1621,N_1585);
nor U2031 (N_2031,N_1413,N_1688);
nor U2032 (N_2032,N_1368,N_1325);
nor U2033 (N_2033,N_1689,N_1395);
nor U2034 (N_2034,N_1583,N_1644);
or U2035 (N_2035,N_1266,N_1246);
nor U2036 (N_2036,N_1272,N_1503);
or U2037 (N_2037,N_1726,N_1472);
and U2038 (N_2038,N_1588,N_1487);
nand U2039 (N_2039,N_1578,N_1762);
nand U2040 (N_2040,N_1638,N_1332);
and U2041 (N_2041,N_1225,N_1771);
nand U2042 (N_2042,N_1518,N_1341);
nand U2043 (N_2043,N_1396,N_1336);
nor U2044 (N_2044,N_1304,N_1216);
nor U2045 (N_2045,N_1335,N_1711);
or U2046 (N_2046,N_1505,N_1431);
nor U2047 (N_2047,N_1370,N_1511);
nand U2048 (N_2048,N_1241,N_1510);
or U2049 (N_2049,N_1782,N_1345);
nand U2050 (N_2050,N_1515,N_1754);
nand U2051 (N_2051,N_1428,N_1263);
nor U2052 (N_2052,N_1206,N_1254);
or U2053 (N_2053,N_1773,N_1742);
nor U2054 (N_2054,N_1207,N_1693);
and U2055 (N_2055,N_1539,N_1622);
or U2056 (N_2056,N_1522,N_1535);
nand U2057 (N_2057,N_1350,N_1745);
nor U2058 (N_2058,N_1706,N_1653);
or U2059 (N_2059,N_1640,N_1303);
and U2060 (N_2060,N_1690,N_1715);
nand U2061 (N_2061,N_1224,N_1603);
or U2062 (N_2062,N_1749,N_1383);
nand U2063 (N_2063,N_1284,N_1637);
and U2064 (N_2064,N_1330,N_1203);
nand U2065 (N_2065,N_1730,N_1707);
or U2066 (N_2066,N_1571,N_1616);
nor U2067 (N_2067,N_1456,N_1780);
or U2068 (N_2068,N_1441,N_1648);
nor U2069 (N_2069,N_1402,N_1714);
and U2070 (N_2070,N_1438,N_1245);
or U2071 (N_2071,N_1555,N_1799);
or U2072 (N_2072,N_1492,N_1405);
nand U2073 (N_2073,N_1646,N_1432);
nand U2074 (N_2074,N_1624,N_1259);
and U2075 (N_2075,N_1559,N_1737);
and U2076 (N_2076,N_1464,N_1433);
or U2077 (N_2077,N_1641,N_1253);
nor U2078 (N_2078,N_1434,N_1312);
nor U2079 (N_2079,N_1600,N_1230);
nand U2080 (N_2080,N_1478,N_1486);
or U2081 (N_2081,N_1717,N_1209);
nor U2082 (N_2082,N_1579,N_1785);
and U2083 (N_2083,N_1343,N_1301);
or U2084 (N_2084,N_1465,N_1258);
nand U2085 (N_2085,N_1703,N_1509);
nand U2086 (N_2086,N_1502,N_1309);
and U2087 (N_2087,N_1727,N_1542);
or U2088 (N_2088,N_1500,N_1439);
nand U2089 (N_2089,N_1779,N_1305);
or U2090 (N_2090,N_1391,N_1551);
nand U2091 (N_2091,N_1670,N_1720);
or U2092 (N_2092,N_1204,N_1575);
and U2093 (N_2093,N_1398,N_1645);
nand U2094 (N_2094,N_1661,N_1200);
nand U2095 (N_2095,N_1415,N_1594);
and U2096 (N_2096,N_1507,N_1297);
nand U2097 (N_2097,N_1520,N_1698);
nor U2098 (N_2098,N_1605,N_1682);
xor U2099 (N_2099,N_1482,N_1604);
or U2100 (N_2100,N_1392,N_1792);
nor U2101 (N_2101,N_1458,N_1470);
or U2102 (N_2102,N_1494,N_1718);
or U2103 (N_2103,N_1759,N_1526);
and U2104 (N_2104,N_1639,N_1644);
nor U2105 (N_2105,N_1229,N_1385);
nand U2106 (N_2106,N_1577,N_1463);
nand U2107 (N_2107,N_1774,N_1317);
nand U2108 (N_2108,N_1479,N_1664);
or U2109 (N_2109,N_1634,N_1656);
nor U2110 (N_2110,N_1655,N_1589);
nor U2111 (N_2111,N_1782,N_1225);
and U2112 (N_2112,N_1490,N_1212);
nor U2113 (N_2113,N_1711,N_1387);
nor U2114 (N_2114,N_1297,N_1485);
nor U2115 (N_2115,N_1755,N_1529);
nand U2116 (N_2116,N_1625,N_1792);
or U2117 (N_2117,N_1697,N_1706);
and U2118 (N_2118,N_1445,N_1672);
or U2119 (N_2119,N_1529,N_1725);
and U2120 (N_2120,N_1440,N_1694);
or U2121 (N_2121,N_1396,N_1406);
or U2122 (N_2122,N_1253,N_1433);
nor U2123 (N_2123,N_1689,N_1364);
nand U2124 (N_2124,N_1482,N_1339);
or U2125 (N_2125,N_1714,N_1738);
and U2126 (N_2126,N_1458,N_1434);
and U2127 (N_2127,N_1638,N_1336);
nor U2128 (N_2128,N_1387,N_1786);
or U2129 (N_2129,N_1447,N_1755);
nand U2130 (N_2130,N_1652,N_1209);
nor U2131 (N_2131,N_1582,N_1642);
nand U2132 (N_2132,N_1622,N_1742);
nand U2133 (N_2133,N_1676,N_1558);
nor U2134 (N_2134,N_1629,N_1635);
nor U2135 (N_2135,N_1593,N_1667);
or U2136 (N_2136,N_1711,N_1634);
and U2137 (N_2137,N_1598,N_1793);
nor U2138 (N_2138,N_1615,N_1357);
nor U2139 (N_2139,N_1216,N_1383);
or U2140 (N_2140,N_1707,N_1627);
nor U2141 (N_2141,N_1245,N_1723);
nor U2142 (N_2142,N_1258,N_1610);
or U2143 (N_2143,N_1680,N_1754);
or U2144 (N_2144,N_1671,N_1323);
and U2145 (N_2145,N_1763,N_1451);
nand U2146 (N_2146,N_1430,N_1581);
and U2147 (N_2147,N_1297,N_1449);
nor U2148 (N_2148,N_1551,N_1416);
nor U2149 (N_2149,N_1381,N_1295);
and U2150 (N_2150,N_1682,N_1691);
or U2151 (N_2151,N_1241,N_1722);
and U2152 (N_2152,N_1448,N_1637);
or U2153 (N_2153,N_1526,N_1541);
and U2154 (N_2154,N_1559,N_1261);
nor U2155 (N_2155,N_1794,N_1780);
and U2156 (N_2156,N_1728,N_1266);
nand U2157 (N_2157,N_1596,N_1501);
or U2158 (N_2158,N_1305,N_1232);
nor U2159 (N_2159,N_1504,N_1694);
or U2160 (N_2160,N_1724,N_1409);
and U2161 (N_2161,N_1793,N_1372);
nor U2162 (N_2162,N_1269,N_1486);
nand U2163 (N_2163,N_1362,N_1761);
or U2164 (N_2164,N_1456,N_1219);
nand U2165 (N_2165,N_1796,N_1370);
nand U2166 (N_2166,N_1228,N_1372);
nor U2167 (N_2167,N_1496,N_1213);
or U2168 (N_2168,N_1781,N_1462);
nand U2169 (N_2169,N_1550,N_1548);
and U2170 (N_2170,N_1321,N_1347);
nor U2171 (N_2171,N_1368,N_1344);
and U2172 (N_2172,N_1732,N_1667);
and U2173 (N_2173,N_1658,N_1387);
and U2174 (N_2174,N_1726,N_1749);
nand U2175 (N_2175,N_1481,N_1484);
or U2176 (N_2176,N_1578,N_1701);
and U2177 (N_2177,N_1480,N_1717);
nand U2178 (N_2178,N_1227,N_1620);
nand U2179 (N_2179,N_1494,N_1576);
nand U2180 (N_2180,N_1346,N_1752);
and U2181 (N_2181,N_1703,N_1676);
and U2182 (N_2182,N_1689,N_1445);
nand U2183 (N_2183,N_1649,N_1508);
or U2184 (N_2184,N_1670,N_1225);
nor U2185 (N_2185,N_1540,N_1461);
and U2186 (N_2186,N_1791,N_1299);
and U2187 (N_2187,N_1516,N_1768);
or U2188 (N_2188,N_1317,N_1701);
nand U2189 (N_2189,N_1243,N_1713);
nand U2190 (N_2190,N_1331,N_1483);
or U2191 (N_2191,N_1500,N_1765);
nor U2192 (N_2192,N_1409,N_1639);
xnor U2193 (N_2193,N_1546,N_1454);
and U2194 (N_2194,N_1512,N_1532);
nor U2195 (N_2195,N_1667,N_1384);
nand U2196 (N_2196,N_1685,N_1232);
and U2197 (N_2197,N_1594,N_1255);
nand U2198 (N_2198,N_1707,N_1388);
and U2199 (N_2199,N_1279,N_1473);
or U2200 (N_2200,N_1413,N_1411);
and U2201 (N_2201,N_1201,N_1435);
nand U2202 (N_2202,N_1357,N_1703);
nand U2203 (N_2203,N_1247,N_1228);
nand U2204 (N_2204,N_1326,N_1769);
nor U2205 (N_2205,N_1616,N_1623);
nor U2206 (N_2206,N_1612,N_1662);
nor U2207 (N_2207,N_1722,N_1745);
nand U2208 (N_2208,N_1299,N_1449);
and U2209 (N_2209,N_1513,N_1715);
nor U2210 (N_2210,N_1292,N_1661);
and U2211 (N_2211,N_1471,N_1683);
or U2212 (N_2212,N_1236,N_1299);
or U2213 (N_2213,N_1478,N_1467);
or U2214 (N_2214,N_1591,N_1244);
nand U2215 (N_2215,N_1326,N_1617);
nand U2216 (N_2216,N_1332,N_1436);
or U2217 (N_2217,N_1269,N_1231);
nand U2218 (N_2218,N_1762,N_1516);
and U2219 (N_2219,N_1585,N_1540);
nand U2220 (N_2220,N_1464,N_1728);
and U2221 (N_2221,N_1524,N_1734);
nor U2222 (N_2222,N_1348,N_1456);
or U2223 (N_2223,N_1759,N_1211);
nand U2224 (N_2224,N_1215,N_1368);
or U2225 (N_2225,N_1327,N_1620);
and U2226 (N_2226,N_1785,N_1583);
and U2227 (N_2227,N_1699,N_1697);
nand U2228 (N_2228,N_1279,N_1581);
nand U2229 (N_2229,N_1209,N_1502);
nor U2230 (N_2230,N_1313,N_1569);
and U2231 (N_2231,N_1738,N_1482);
nand U2232 (N_2232,N_1359,N_1305);
nand U2233 (N_2233,N_1691,N_1661);
nor U2234 (N_2234,N_1499,N_1290);
or U2235 (N_2235,N_1501,N_1702);
or U2236 (N_2236,N_1564,N_1613);
and U2237 (N_2237,N_1671,N_1284);
nand U2238 (N_2238,N_1680,N_1431);
nor U2239 (N_2239,N_1279,N_1305);
or U2240 (N_2240,N_1441,N_1527);
or U2241 (N_2241,N_1381,N_1258);
nor U2242 (N_2242,N_1506,N_1215);
nand U2243 (N_2243,N_1252,N_1549);
or U2244 (N_2244,N_1474,N_1787);
and U2245 (N_2245,N_1672,N_1503);
nand U2246 (N_2246,N_1297,N_1570);
nand U2247 (N_2247,N_1503,N_1226);
or U2248 (N_2248,N_1316,N_1417);
or U2249 (N_2249,N_1249,N_1294);
and U2250 (N_2250,N_1767,N_1719);
and U2251 (N_2251,N_1291,N_1294);
nor U2252 (N_2252,N_1560,N_1363);
nand U2253 (N_2253,N_1441,N_1242);
or U2254 (N_2254,N_1644,N_1476);
nand U2255 (N_2255,N_1779,N_1253);
nand U2256 (N_2256,N_1513,N_1312);
nand U2257 (N_2257,N_1472,N_1301);
nand U2258 (N_2258,N_1229,N_1419);
nand U2259 (N_2259,N_1252,N_1589);
and U2260 (N_2260,N_1758,N_1224);
nand U2261 (N_2261,N_1253,N_1701);
or U2262 (N_2262,N_1580,N_1743);
or U2263 (N_2263,N_1382,N_1789);
nand U2264 (N_2264,N_1289,N_1605);
or U2265 (N_2265,N_1436,N_1258);
nand U2266 (N_2266,N_1633,N_1677);
nand U2267 (N_2267,N_1388,N_1261);
and U2268 (N_2268,N_1292,N_1646);
or U2269 (N_2269,N_1728,N_1224);
nand U2270 (N_2270,N_1786,N_1401);
nand U2271 (N_2271,N_1437,N_1721);
or U2272 (N_2272,N_1347,N_1323);
nor U2273 (N_2273,N_1780,N_1689);
and U2274 (N_2274,N_1759,N_1210);
nor U2275 (N_2275,N_1688,N_1412);
nor U2276 (N_2276,N_1572,N_1387);
nand U2277 (N_2277,N_1395,N_1344);
xor U2278 (N_2278,N_1531,N_1705);
and U2279 (N_2279,N_1441,N_1339);
or U2280 (N_2280,N_1333,N_1702);
or U2281 (N_2281,N_1642,N_1284);
or U2282 (N_2282,N_1676,N_1539);
nor U2283 (N_2283,N_1681,N_1312);
nor U2284 (N_2284,N_1720,N_1500);
and U2285 (N_2285,N_1355,N_1439);
and U2286 (N_2286,N_1554,N_1284);
nand U2287 (N_2287,N_1439,N_1615);
nor U2288 (N_2288,N_1375,N_1336);
nand U2289 (N_2289,N_1779,N_1387);
nor U2290 (N_2290,N_1745,N_1211);
and U2291 (N_2291,N_1228,N_1421);
or U2292 (N_2292,N_1340,N_1499);
nor U2293 (N_2293,N_1547,N_1466);
nand U2294 (N_2294,N_1793,N_1232);
nand U2295 (N_2295,N_1309,N_1585);
nand U2296 (N_2296,N_1250,N_1552);
nand U2297 (N_2297,N_1206,N_1536);
nor U2298 (N_2298,N_1572,N_1371);
and U2299 (N_2299,N_1691,N_1259);
or U2300 (N_2300,N_1498,N_1742);
nand U2301 (N_2301,N_1233,N_1214);
and U2302 (N_2302,N_1237,N_1333);
and U2303 (N_2303,N_1501,N_1260);
and U2304 (N_2304,N_1388,N_1387);
and U2305 (N_2305,N_1603,N_1309);
or U2306 (N_2306,N_1310,N_1357);
nand U2307 (N_2307,N_1671,N_1413);
or U2308 (N_2308,N_1425,N_1463);
nor U2309 (N_2309,N_1382,N_1666);
or U2310 (N_2310,N_1549,N_1499);
or U2311 (N_2311,N_1305,N_1272);
nor U2312 (N_2312,N_1225,N_1791);
nand U2313 (N_2313,N_1773,N_1340);
or U2314 (N_2314,N_1765,N_1780);
or U2315 (N_2315,N_1567,N_1223);
and U2316 (N_2316,N_1397,N_1525);
and U2317 (N_2317,N_1405,N_1656);
nor U2318 (N_2318,N_1712,N_1629);
nand U2319 (N_2319,N_1227,N_1473);
and U2320 (N_2320,N_1490,N_1501);
nor U2321 (N_2321,N_1280,N_1487);
or U2322 (N_2322,N_1318,N_1468);
nand U2323 (N_2323,N_1395,N_1411);
nor U2324 (N_2324,N_1309,N_1425);
nor U2325 (N_2325,N_1573,N_1626);
and U2326 (N_2326,N_1702,N_1377);
nand U2327 (N_2327,N_1793,N_1364);
and U2328 (N_2328,N_1749,N_1329);
nor U2329 (N_2329,N_1667,N_1450);
nor U2330 (N_2330,N_1325,N_1317);
nand U2331 (N_2331,N_1699,N_1226);
xnor U2332 (N_2332,N_1355,N_1379);
nor U2333 (N_2333,N_1288,N_1670);
nor U2334 (N_2334,N_1417,N_1760);
and U2335 (N_2335,N_1714,N_1624);
or U2336 (N_2336,N_1236,N_1656);
xnor U2337 (N_2337,N_1494,N_1474);
nand U2338 (N_2338,N_1269,N_1559);
nor U2339 (N_2339,N_1203,N_1748);
nand U2340 (N_2340,N_1700,N_1344);
nor U2341 (N_2341,N_1540,N_1712);
nor U2342 (N_2342,N_1266,N_1224);
nand U2343 (N_2343,N_1652,N_1628);
or U2344 (N_2344,N_1641,N_1200);
and U2345 (N_2345,N_1657,N_1683);
or U2346 (N_2346,N_1691,N_1371);
nor U2347 (N_2347,N_1582,N_1536);
or U2348 (N_2348,N_1597,N_1353);
nand U2349 (N_2349,N_1207,N_1247);
nor U2350 (N_2350,N_1778,N_1688);
nor U2351 (N_2351,N_1787,N_1687);
and U2352 (N_2352,N_1283,N_1217);
nor U2353 (N_2353,N_1503,N_1470);
nand U2354 (N_2354,N_1539,N_1674);
or U2355 (N_2355,N_1233,N_1288);
nor U2356 (N_2356,N_1756,N_1660);
nand U2357 (N_2357,N_1587,N_1428);
or U2358 (N_2358,N_1662,N_1417);
and U2359 (N_2359,N_1232,N_1370);
and U2360 (N_2360,N_1517,N_1734);
or U2361 (N_2361,N_1280,N_1646);
nor U2362 (N_2362,N_1659,N_1609);
or U2363 (N_2363,N_1499,N_1614);
nor U2364 (N_2364,N_1247,N_1266);
or U2365 (N_2365,N_1538,N_1409);
nor U2366 (N_2366,N_1280,N_1578);
and U2367 (N_2367,N_1241,N_1704);
nand U2368 (N_2368,N_1625,N_1555);
nor U2369 (N_2369,N_1687,N_1783);
and U2370 (N_2370,N_1620,N_1418);
and U2371 (N_2371,N_1737,N_1615);
nand U2372 (N_2372,N_1721,N_1245);
and U2373 (N_2373,N_1783,N_1671);
or U2374 (N_2374,N_1278,N_1799);
or U2375 (N_2375,N_1366,N_1341);
nor U2376 (N_2376,N_1748,N_1276);
or U2377 (N_2377,N_1520,N_1418);
nor U2378 (N_2378,N_1421,N_1561);
or U2379 (N_2379,N_1377,N_1658);
xor U2380 (N_2380,N_1257,N_1316);
nand U2381 (N_2381,N_1530,N_1368);
nand U2382 (N_2382,N_1716,N_1422);
nand U2383 (N_2383,N_1381,N_1231);
or U2384 (N_2384,N_1408,N_1581);
nor U2385 (N_2385,N_1434,N_1555);
nand U2386 (N_2386,N_1254,N_1539);
nor U2387 (N_2387,N_1758,N_1649);
nor U2388 (N_2388,N_1332,N_1434);
xnor U2389 (N_2389,N_1423,N_1497);
and U2390 (N_2390,N_1627,N_1481);
nand U2391 (N_2391,N_1240,N_1348);
and U2392 (N_2392,N_1573,N_1366);
or U2393 (N_2393,N_1280,N_1517);
or U2394 (N_2394,N_1616,N_1483);
nor U2395 (N_2395,N_1670,N_1528);
and U2396 (N_2396,N_1428,N_1731);
nor U2397 (N_2397,N_1343,N_1372);
and U2398 (N_2398,N_1796,N_1661);
xor U2399 (N_2399,N_1612,N_1464);
and U2400 (N_2400,N_2024,N_2236);
or U2401 (N_2401,N_2032,N_2175);
or U2402 (N_2402,N_2292,N_2152);
nor U2403 (N_2403,N_2200,N_2077);
and U2404 (N_2404,N_1991,N_2297);
nor U2405 (N_2405,N_2129,N_2377);
nand U2406 (N_2406,N_1847,N_2180);
nand U2407 (N_2407,N_2125,N_1978);
and U2408 (N_2408,N_1984,N_2346);
and U2409 (N_2409,N_1873,N_1801);
or U2410 (N_2410,N_2293,N_2307);
nand U2411 (N_2411,N_1952,N_2189);
nand U2412 (N_2412,N_1890,N_2280);
and U2413 (N_2413,N_2347,N_1900);
nor U2414 (N_2414,N_2351,N_2209);
or U2415 (N_2415,N_2358,N_1904);
nand U2416 (N_2416,N_2287,N_2191);
and U2417 (N_2417,N_2102,N_2273);
nand U2418 (N_2418,N_1815,N_1851);
nor U2419 (N_2419,N_2317,N_2006);
or U2420 (N_2420,N_2373,N_1849);
nand U2421 (N_2421,N_2362,N_1889);
nor U2422 (N_2422,N_1800,N_1893);
and U2423 (N_2423,N_1988,N_2336);
nor U2424 (N_2424,N_2319,N_2310);
xor U2425 (N_2425,N_1817,N_1961);
nor U2426 (N_2426,N_2177,N_1941);
and U2427 (N_2427,N_2368,N_2092);
nor U2428 (N_2428,N_1888,N_1938);
nand U2429 (N_2429,N_1979,N_2242);
or U2430 (N_2430,N_1841,N_1870);
and U2431 (N_2431,N_2141,N_2155);
and U2432 (N_2432,N_2353,N_1826);
nand U2433 (N_2433,N_2188,N_2265);
nor U2434 (N_2434,N_2233,N_1839);
and U2435 (N_2435,N_2179,N_2207);
and U2436 (N_2436,N_2137,N_2309);
and U2437 (N_2437,N_1804,N_2033);
nor U2438 (N_2438,N_1875,N_2302);
and U2439 (N_2439,N_1896,N_2329);
nand U2440 (N_2440,N_1958,N_2374);
or U2441 (N_2441,N_1866,N_1932);
nor U2442 (N_2442,N_1884,N_2305);
nor U2443 (N_2443,N_1955,N_1886);
nor U2444 (N_2444,N_2354,N_2038);
and U2445 (N_2445,N_1942,N_2192);
and U2446 (N_2446,N_2007,N_2308);
and U2447 (N_2447,N_2255,N_1969);
nand U2448 (N_2448,N_2037,N_1928);
nor U2449 (N_2449,N_2258,N_2132);
nand U2450 (N_2450,N_2253,N_1953);
or U2451 (N_2451,N_2254,N_1895);
nand U2452 (N_2452,N_2383,N_2378);
nand U2453 (N_2453,N_2311,N_2040);
or U2454 (N_2454,N_2081,N_1980);
nor U2455 (N_2455,N_2110,N_1926);
nand U2456 (N_2456,N_1905,N_1945);
or U2457 (N_2457,N_1913,N_2048);
nor U2458 (N_2458,N_1936,N_2013);
or U2459 (N_2459,N_2387,N_2187);
nor U2460 (N_2460,N_2153,N_2026);
and U2461 (N_2461,N_2195,N_1807);
or U2462 (N_2462,N_1819,N_2244);
nand U2463 (N_2463,N_1967,N_2285);
and U2464 (N_2464,N_1894,N_2136);
and U2465 (N_2465,N_2214,N_2343);
or U2466 (N_2466,N_2010,N_1973);
and U2467 (N_2467,N_2304,N_1805);
nand U2468 (N_2468,N_1927,N_1923);
nor U2469 (N_2469,N_2279,N_1962);
and U2470 (N_2470,N_2295,N_2221);
nand U2471 (N_2471,N_1982,N_2201);
nor U2472 (N_2472,N_2320,N_2372);
nor U2473 (N_2473,N_2059,N_2104);
or U2474 (N_2474,N_2264,N_1947);
or U2475 (N_2475,N_1881,N_1917);
nor U2476 (N_2476,N_2381,N_2086);
nand U2477 (N_2477,N_2331,N_2072);
nand U2478 (N_2478,N_1874,N_2342);
nand U2479 (N_2479,N_2193,N_1899);
nand U2480 (N_2480,N_2229,N_1972);
and U2481 (N_2481,N_2326,N_2078);
nor U2482 (N_2482,N_2299,N_2259);
nor U2483 (N_2483,N_2124,N_1957);
nand U2484 (N_2484,N_2105,N_2256);
nand U2485 (N_2485,N_1857,N_2111);
or U2486 (N_2486,N_2252,N_1990);
or U2487 (N_2487,N_2237,N_2389);
nand U2488 (N_2488,N_1821,N_2087);
or U2489 (N_2489,N_2118,N_1983);
or U2490 (N_2490,N_2199,N_2097);
and U2491 (N_2491,N_2376,N_2239);
or U2492 (N_2492,N_2384,N_2235);
and U2493 (N_2493,N_2306,N_1840);
or U2494 (N_2494,N_2186,N_1822);
or U2495 (N_2495,N_2162,N_1861);
nor U2496 (N_2496,N_2350,N_2286);
and U2497 (N_2497,N_2041,N_1876);
nor U2498 (N_2498,N_1976,N_2080);
nor U2499 (N_2499,N_1824,N_2208);
xor U2500 (N_2500,N_2194,N_2181);
nor U2501 (N_2501,N_2380,N_1834);
or U2502 (N_2502,N_2120,N_1850);
nand U2503 (N_2503,N_2044,N_1838);
or U2504 (N_2504,N_2396,N_2333);
and U2505 (N_2505,N_1863,N_2005);
nor U2506 (N_2506,N_1831,N_2390);
or U2507 (N_2507,N_2215,N_2232);
nand U2508 (N_2508,N_1856,N_2168);
and U2509 (N_2509,N_2067,N_2382);
or U2510 (N_2510,N_2028,N_2267);
nor U2511 (N_2511,N_1914,N_1999);
and U2512 (N_2512,N_1996,N_2093);
nand U2513 (N_2513,N_1814,N_2314);
and U2514 (N_2514,N_2294,N_1827);
nor U2515 (N_2515,N_2147,N_2001);
or U2516 (N_2516,N_2017,N_2340);
nand U2517 (N_2517,N_1989,N_2313);
nor U2518 (N_2518,N_1971,N_2084);
and U2519 (N_2519,N_2282,N_2338);
and U2520 (N_2520,N_2290,N_1846);
nor U2521 (N_2521,N_2158,N_2062);
nor U2522 (N_2522,N_2133,N_1922);
or U2523 (N_2523,N_2126,N_2174);
or U2524 (N_2524,N_2055,N_2106);
nor U2525 (N_2525,N_2231,N_1937);
or U2526 (N_2526,N_1825,N_1836);
and U2527 (N_2527,N_2240,N_2176);
nor U2528 (N_2528,N_2219,N_1879);
and U2529 (N_2529,N_2052,N_2357);
and U2530 (N_2530,N_2369,N_2054);
nor U2531 (N_2531,N_2170,N_2130);
nand U2532 (N_2532,N_1985,N_1960);
and U2533 (N_2533,N_2008,N_2296);
and U2534 (N_2534,N_2197,N_2341);
nand U2535 (N_2535,N_2321,N_2392);
or U2536 (N_2536,N_2075,N_2167);
nor U2537 (N_2537,N_2004,N_2324);
and U2538 (N_2538,N_2251,N_2039);
or U2539 (N_2539,N_2330,N_1810);
or U2540 (N_2540,N_2337,N_2128);
and U2541 (N_2541,N_1871,N_2089);
nor U2542 (N_2542,N_2360,N_2327);
nand U2543 (N_2543,N_2165,N_2122);
nor U2544 (N_2544,N_2113,N_2359);
or U2545 (N_2545,N_1907,N_1931);
or U2546 (N_2546,N_1934,N_2046);
nor U2547 (N_2547,N_2159,N_1993);
and U2548 (N_2548,N_2303,N_2246);
and U2549 (N_2549,N_1939,N_2068);
nor U2550 (N_2550,N_1992,N_2289);
or U2551 (N_2551,N_2071,N_1948);
and U2552 (N_2552,N_2114,N_2397);
nor U2553 (N_2553,N_2198,N_2030);
or U2554 (N_2554,N_2213,N_1956);
nor U2555 (N_2555,N_2393,N_1997);
and U2556 (N_2556,N_2027,N_2074);
nand U2557 (N_2557,N_1898,N_2352);
and U2558 (N_2558,N_2160,N_2216);
nand U2559 (N_2559,N_2015,N_2395);
and U2560 (N_2560,N_1887,N_2349);
nor U2561 (N_2561,N_1883,N_2049);
and U2562 (N_2562,N_1858,N_2036);
and U2563 (N_2563,N_2140,N_1950);
and U2564 (N_2564,N_2356,N_1964);
or U2565 (N_2565,N_2183,N_2250);
nor U2566 (N_2566,N_2012,N_2366);
nor U2567 (N_2567,N_2116,N_1920);
nand U2568 (N_2568,N_2217,N_2161);
nor U2569 (N_2569,N_1994,N_2371);
and U2570 (N_2570,N_2370,N_1812);
nand U2571 (N_2571,N_2016,N_1987);
or U2572 (N_2572,N_2249,N_2069);
and U2573 (N_2573,N_2151,N_2021);
or U2574 (N_2574,N_1806,N_2149);
nor U2575 (N_2575,N_2112,N_2230);
or U2576 (N_2576,N_2065,N_1974);
nor U2577 (N_2577,N_2190,N_2185);
nor U2578 (N_2578,N_2243,N_2182);
and U2579 (N_2579,N_1835,N_2247);
nor U2580 (N_2580,N_1933,N_2011);
nor U2581 (N_2581,N_2066,N_1860);
and U2582 (N_2582,N_2139,N_2261);
nand U2583 (N_2583,N_2163,N_2014);
nand U2584 (N_2584,N_2019,N_2127);
nand U2585 (N_2585,N_2063,N_2070);
and U2586 (N_2586,N_2042,N_1803);
nor U2587 (N_2587,N_2100,N_1998);
or U2588 (N_2588,N_2076,N_2029);
nor U2589 (N_2589,N_2103,N_2000);
xnor U2590 (N_2590,N_2091,N_2386);
or U2591 (N_2591,N_2257,N_2318);
nand U2592 (N_2592,N_1892,N_2043);
nand U2593 (N_2593,N_1864,N_1897);
and U2594 (N_2594,N_1959,N_1921);
nand U2595 (N_2595,N_1930,N_2073);
nor U2596 (N_2596,N_1880,N_2328);
or U2597 (N_2597,N_1924,N_2051);
or U2598 (N_2598,N_2344,N_2107);
and U2599 (N_2599,N_2365,N_1963);
and U2600 (N_2600,N_1811,N_2009);
nand U2601 (N_2601,N_2144,N_2143);
and U2602 (N_2602,N_1925,N_2325);
nor U2603 (N_2603,N_2345,N_2355);
and U2604 (N_2604,N_1813,N_2266);
nand U2605 (N_2605,N_2241,N_2298);
or U2606 (N_2606,N_2145,N_1903);
nor U2607 (N_2607,N_1816,N_2117);
nand U2608 (N_2608,N_1949,N_1820);
or U2609 (N_2609,N_2108,N_2061);
nand U2610 (N_2610,N_2002,N_1970);
or U2611 (N_2611,N_2225,N_2034);
nor U2612 (N_2612,N_2098,N_2332);
nand U2613 (N_2613,N_1995,N_2099);
nor U2614 (N_2614,N_2101,N_2123);
or U2615 (N_2615,N_1916,N_1869);
nand U2616 (N_2616,N_1918,N_2394);
nand U2617 (N_2617,N_2142,N_2220);
and U2618 (N_2618,N_2053,N_2268);
nand U2619 (N_2619,N_2398,N_2288);
or U2620 (N_2620,N_2134,N_1981);
or U2621 (N_2621,N_2003,N_1823);
or U2622 (N_2622,N_2315,N_2284);
and U2623 (N_2623,N_1940,N_1867);
nor U2624 (N_2624,N_2323,N_2270);
nand U2625 (N_2625,N_1818,N_2269);
nor U2626 (N_2626,N_2184,N_2204);
nor U2627 (N_2627,N_2224,N_2023);
and U2628 (N_2628,N_2379,N_2079);
and U2629 (N_2629,N_2385,N_2173);
or U2630 (N_2630,N_2399,N_1832);
and U2631 (N_2631,N_1837,N_1865);
nand U2632 (N_2632,N_2090,N_1902);
or U2633 (N_2633,N_2218,N_2271);
nor U2634 (N_2634,N_2025,N_1845);
or U2635 (N_2635,N_1882,N_2156);
and U2636 (N_2636,N_2361,N_1965);
or U2637 (N_2637,N_2367,N_2234);
or U2638 (N_2638,N_2064,N_1862);
nor U2639 (N_2639,N_1935,N_2281);
or U2640 (N_2640,N_2096,N_2223);
nor U2641 (N_2641,N_2300,N_1975);
and U2642 (N_2642,N_2301,N_1854);
nand U2643 (N_2643,N_1977,N_1848);
and U2644 (N_2644,N_1859,N_2222);
nand U2645 (N_2645,N_2057,N_2226);
nand U2646 (N_2646,N_1908,N_2157);
and U2647 (N_2647,N_2322,N_1872);
and U2648 (N_2648,N_1910,N_2150);
or U2649 (N_2649,N_2245,N_2283);
nor U2650 (N_2650,N_1853,N_2083);
nand U2651 (N_2651,N_2050,N_1919);
and U2652 (N_2652,N_1842,N_1828);
and U2653 (N_2653,N_2291,N_2206);
nand U2654 (N_2654,N_2227,N_2262);
nor U2655 (N_2655,N_1909,N_2115);
nor U2656 (N_2656,N_2022,N_2121);
nor U2657 (N_2657,N_2131,N_1906);
and U2658 (N_2658,N_1809,N_2169);
nor U2659 (N_2659,N_2164,N_1844);
nor U2660 (N_2660,N_1912,N_1829);
and U2661 (N_2661,N_2060,N_1878);
and U2662 (N_2662,N_1954,N_2276);
nor U2663 (N_2663,N_2238,N_2263);
and U2664 (N_2664,N_1830,N_2035);
nand U2665 (N_2665,N_1946,N_2278);
nand U2666 (N_2666,N_2082,N_2312);
and U2667 (N_2667,N_2248,N_1911);
nand U2668 (N_2668,N_2045,N_2085);
or U2669 (N_2669,N_2146,N_1915);
xnor U2670 (N_2670,N_2272,N_1802);
and U2671 (N_2671,N_1833,N_1808);
and U2672 (N_2672,N_2109,N_1943);
nor U2673 (N_2673,N_2202,N_1843);
and U2674 (N_2674,N_2316,N_2205);
nand U2675 (N_2675,N_1868,N_2018);
nor U2676 (N_2676,N_2166,N_1901);
nor U2677 (N_2677,N_2260,N_2138);
and U2678 (N_2678,N_2334,N_2274);
and U2679 (N_2679,N_2388,N_1877);
or U2680 (N_2680,N_2058,N_2339);
or U2681 (N_2681,N_2203,N_2363);
and U2682 (N_2682,N_2275,N_1944);
and U2683 (N_2683,N_2020,N_1929);
and U2684 (N_2684,N_2088,N_1966);
nand U2685 (N_2685,N_2171,N_2211);
nand U2686 (N_2686,N_2119,N_1852);
or U2687 (N_2687,N_2375,N_2154);
and U2688 (N_2688,N_1986,N_2148);
nand U2689 (N_2689,N_2031,N_1968);
and U2690 (N_2690,N_2056,N_2172);
and U2691 (N_2691,N_2094,N_2196);
nand U2692 (N_2692,N_2135,N_1885);
or U2693 (N_2693,N_2210,N_2348);
and U2694 (N_2694,N_2364,N_2212);
nor U2695 (N_2695,N_1891,N_2178);
nor U2696 (N_2696,N_2228,N_2277);
and U2697 (N_2697,N_2047,N_2391);
and U2698 (N_2698,N_2335,N_1855);
and U2699 (N_2699,N_1951,N_2095);
and U2700 (N_2700,N_2302,N_2159);
nand U2701 (N_2701,N_1999,N_2308);
xnor U2702 (N_2702,N_1862,N_2173);
nor U2703 (N_2703,N_1822,N_1970);
nor U2704 (N_2704,N_2019,N_2139);
nand U2705 (N_2705,N_2057,N_2121);
or U2706 (N_2706,N_2397,N_1952);
nand U2707 (N_2707,N_1801,N_2379);
or U2708 (N_2708,N_2104,N_2065);
or U2709 (N_2709,N_2282,N_2020);
or U2710 (N_2710,N_1927,N_1991);
or U2711 (N_2711,N_2252,N_2395);
or U2712 (N_2712,N_1996,N_2034);
or U2713 (N_2713,N_1966,N_1886);
nor U2714 (N_2714,N_2322,N_1948);
and U2715 (N_2715,N_2136,N_1832);
or U2716 (N_2716,N_1881,N_2133);
and U2717 (N_2717,N_2000,N_2115);
nor U2718 (N_2718,N_1911,N_1876);
or U2719 (N_2719,N_1891,N_2128);
nor U2720 (N_2720,N_2162,N_2183);
and U2721 (N_2721,N_2048,N_2085);
or U2722 (N_2722,N_2367,N_2102);
nor U2723 (N_2723,N_2078,N_1959);
nand U2724 (N_2724,N_1841,N_2178);
nor U2725 (N_2725,N_2008,N_2175);
and U2726 (N_2726,N_1891,N_2034);
and U2727 (N_2727,N_2348,N_2337);
nand U2728 (N_2728,N_1984,N_2302);
or U2729 (N_2729,N_2044,N_2063);
nand U2730 (N_2730,N_2107,N_1973);
nand U2731 (N_2731,N_1878,N_2172);
nand U2732 (N_2732,N_2052,N_1834);
or U2733 (N_2733,N_2295,N_2020);
nor U2734 (N_2734,N_1893,N_1990);
nand U2735 (N_2735,N_2234,N_2186);
and U2736 (N_2736,N_2063,N_2192);
or U2737 (N_2737,N_2382,N_2027);
or U2738 (N_2738,N_2236,N_2082);
and U2739 (N_2739,N_2388,N_1887);
or U2740 (N_2740,N_1847,N_1986);
and U2741 (N_2741,N_2140,N_1877);
and U2742 (N_2742,N_2332,N_1991);
or U2743 (N_2743,N_2317,N_2348);
nand U2744 (N_2744,N_2059,N_2369);
and U2745 (N_2745,N_2264,N_2354);
and U2746 (N_2746,N_2388,N_1998);
or U2747 (N_2747,N_2240,N_2251);
nor U2748 (N_2748,N_2331,N_1957);
or U2749 (N_2749,N_2392,N_2062);
and U2750 (N_2750,N_2302,N_2367);
and U2751 (N_2751,N_1807,N_2203);
nor U2752 (N_2752,N_2182,N_2094);
or U2753 (N_2753,N_1909,N_2137);
or U2754 (N_2754,N_2165,N_1969);
or U2755 (N_2755,N_2043,N_1963);
or U2756 (N_2756,N_2356,N_1992);
and U2757 (N_2757,N_2039,N_2024);
or U2758 (N_2758,N_1819,N_2028);
nor U2759 (N_2759,N_2063,N_2000);
and U2760 (N_2760,N_2274,N_1908);
and U2761 (N_2761,N_2127,N_2239);
or U2762 (N_2762,N_1896,N_1823);
and U2763 (N_2763,N_2319,N_1865);
nand U2764 (N_2764,N_2175,N_1809);
nand U2765 (N_2765,N_1931,N_2179);
or U2766 (N_2766,N_1853,N_2120);
or U2767 (N_2767,N_2223,N_2304);
and U2768 (N_2768,N_2146,N_2344);
or U2769 (N_2769,N_1974,N_1913);
or U2770 (N_2770,N_2354,N_2168);
nand U2771 (N_2771,N_2320,N_2253);
or U2772 (N_2772,N_2182,N_2252);
nand U2773 (N_2773,N_2338,N_1941);
nor U2774 (N_2774,N_2101,N_2085);
nor U2775 (N_2775,N_2025,N_1816);
nand U2776 (N_2776,N_2011,N_2134);
nor U2777 (N_2777,N_2151,N_2302);
or U2778 (N_2778,N_1963,N_2376);
and U2779 (N_2779,N_2392,N_1870);
and U2780 (N_2780,N_2101,N_2027);
nand U2781 (N_2781,N_1920,N_2090);
xnor U2782 (N_2782,N_2260,N_2066);
or U2783 (N_2783,N_1948,N_2229);
nor U2784 (N_2784,N_1933,N_2279);
nand U2785 (N_2785,N_2367,N_2382);
nor U2786 (N_2786,N_2152,N_2120);
nand U2787 (N_2787,N_1973,N_2186);
nand U2788 (N_2788,N_2028,N_2289);
nand U2789 (N_2789,N_1800,N_2252);
nand U2790 (N_2790,N_2328,N_2043);
and U2791 (N_2791,N_1924,N_2102);
and U2792 (N_2792,N_2087,N_2180);
and U2793 (N_2793,N_1917,N_1867);
nand U2794 (N_2794,N_1928,N_2296);
nor U2795 (N_2795,N_1968,N_1856);
and U2796 (N_2796,N_2061,N_1931);
and U2797 (N_2797,N_2366,N_2104);
and U2798 (N_2798,N_2086,N_1994);
nand U2799 (N_2799,N_1986,N_2185);
or U2800 (N_2800,N_2176,N_2200);
and U2801 (N_2801,N_1938,N_2175);
and U2802 (N_2802,N_2162,N_1845);
and U2803 (N_2803,N_2306,N_1804);
nand U2804 (N_2804,N_2295,N_2049);
nor U2805 (N_2805,N_2148,N_1894);
and U2806 (N_2806,N_1857,N_1871);
nand U2807 (N_2807,N_1921,N_2132);
nand U2808 (N_2808,N_1956,N_1947);
or U2809 (N_2809,N_1890,N_2179);
xnor U2810 (N_2810,N_1970,N_1926);
or U2811 (N_2811,N_2372,N_1946);
and U2812 (N_2812,N_2373,N_2222);
nand U2813 (N_2813,N_1859,N_2158);
and U2814 (N_2814,N_2003,N_1941);
nand U2815 (N_2815,N_1851,N_2081);
and U2816 (N_2816,N_1821,N_2036);
nand U2817 (N_2817,N_2163,N_2040);
nand U2818 (N_2818,N_2124,N_2228);
nand U2819 (N_2819,N_2064,N_1897);
or U2820 (N_2820,N_2083,N_2152);
and U2821 (N_2821,N_1858,N_2002);
nor U2822 (N_2822,N_1934,N_2289);
nand U2823 (N_2823,N_2093,N_2012);
or U2824 (N_2824,N_2169,N_2074);
or U2825 (N_2825,N_1969,N_2124);
and U2826 (N_2826,N_2280,N_1993);
or U2827 (N_2827,N_2054,N_2210);
or U2828 (N_2828,N_1917,N_2224);
or U2829 (N_2829,N_2261,N_2179);
or U2830 (N_2830,N_2012,N_2050);
nor U2831 (N_2831,N_1941,N_2141);
nor U2832 (N_2832,N_1926,N_2113);
and U2833 (N_2833,N_2112,N_2036);
and U2834 (N_2834,N_2091,N_1888);
xor U2835 (N_2835,N_2136,N_1918);
nor U2836 (N_2836,N_2363,N_2367);
nor U2837 (N_2837,N_2391,N_1946);
or U2838 (N_2838,N_2107,N_2113);
nor U2839 (N_2839,N_2068,N_2187);
and U2840 (N_2840,N_2027,N_1849);
nor U2841 (N_2841,N_2014,N_2394);
nand U2842 (N_2842,N_2004,N_1920);
and U2843 (N_2843,N_1865,N_2323);
nand U2844 (N_2844,N_2195,N_2031);
nand U2845 (N_2845,N_1812,N_2171);
and U2846 (N_2846,N_2157,N_2343);
and U2847 (N_2847,N_2163,N_1885);
or U2848 (N_2848,N_1809,N_2084);
nor U2849 (N_2849,N_1996,N_2399);
and U2850 (N_2850,N_2121,N_2026);
nor U2851 (N_2851,N_2072,N_2246);
or U2852 (N_2852,N_2135,N_2002);
nor U2853 (N_2853,N_1970,N_2032);
nand U2854 (N_2854,N_1824,N_1876);
and U2855 (N_2855,N_1935,N_2108);
xor U2856 (N_2856,N_2209,N_2045);
and U2857 (N_2857,N_2038,N_2266);
and U2858 (N_2858,N_2131,N_2148);
nand U2859 (N_2859,N_1909,N_2168);
nand U2860 (N_2860,N_2311,N_2021);
or U2861 (N_2861,N_2363,N_2144);
nand U2862 (N_2862,N_2166,N_1931);
nor U2863 (N_2863,N_2190,N_2362);
nor U2864 (N_2864,N_2218,N_2079);
and U2865 (N_2865,N_1829,N_2278);
or U2866 (N_2866,N_2086,N_2389);
or U2867 (N_2867,N_2236,N_1868);
or U2868 (N_2868,N_2131,N_2250);
nand U2869 (N_2869,N_2373,N_2073);
or U2870 (N_2870,N_2316,N_1941);
nor U2871 (N_2871,N_2098,N_2205);
and U2872 (N_2872,N_2391,N_2037);
or U2873 (N_2873,N_2204,N_1889);
and U2874 (N_2874,N_1815,N_2194);
or U2875 (N_2875,N_2100,N_2204);
nand U2876 (N_2876,N_2188,N_2256);
or U2877 (N_2877,N_1817,N_2097);
or U2878 (N_2878,N_2339,N_2359);
or U2879 (N_2879,N_2317,N_1826);
nor U2880 (N_2880,N_1998,N_2160);
and U2881 (N_2881,N_2317,N_2299);
nor U2882 (N_2882,N_2108,N_2399);
nor U2883 (N_2883,N_2187,N_1822);
nor U2884 (N_2884,N_2072,N_2085);
nand U2885 (N_2885,N_2090,N_1901);
and U2886 (N_2886,N_1927,N_2398);
and U2887 (N_2887,N_1972,N_2067);
and U2888 (N_2888,N_1835,N_2033);
or U2889 (N_2889,N_2248,N_1997);
or U2890 (N_2890,N_2121,N_2002);
or U2891 (N_2891,N_2399,N_2209);
nand U2892 (N_2892,N_2156,N_1841);
and U2893 (N_2893,N_1897,N_2196);
or U2894 (N_2894,N_2301,N_1807);
or U2895 (N_2895,N_2048,N_2389);
and U2896 (N_2896,N_2143,N_1904);
nand U2897 (N_2897,N_1878,N_2287);
or U2898 (N_2898,N_1950,N_1985);
nand U2899 (N_2899,N_2110,N_1901);
or U2900 (N_2900,N_2041,N_2148);
nor U2901 (N_2901,N_2300,N_1827);
or U2902 (N_2902,N_2393,N_1829);
nor U2903 (N_2903,N_2193,N_1981);
nor U2904 (N_2904,N_1862,N_2046);
nor U2905 (N_2905,N_1934,N_2126);
and U2906 (N_2906,N_2282,N_2201);
and U2907 (N_2907,N_2277,N_2176);
and U2908 (N_2908,N_2076,N_2109);
and U2909 (N_2909,N_2357,N_2274);
and U2910 (N_2910,N_2042,N_2351);
nor U2911 (N_2911,N_2170,N_2122);
and U2912 (N_2912,N_2081,N_2165);
nor U2913 (N_2913,N_1907,N_2088);
or U2914 (N_2914,N_1812,N_2110);
nand U2915 (N_2915,N_2283,N_2034);
nor U2916 (N_2916,N_2306,N_2025);
or U2917 (N_2917,N_2293,N_2072);
nand U2918 (N_2918,N_1887,N_2060);
and U2919 (N_2919,N_1965,N_1947);
nand U2920 (N_2920,N_2230,N_2233);
and U2921 (N_2921,N_2122,N_2073);
and U2922 (N_2922,N_2045,N_2172);
or U2923 (N_2923,N_2278,N_2111);
or U2924 (N_2924,N_2241,N_2244);
nor U2925 (N_2925,N_2338,N_2116);
or U2926 (N_2926,N_1948,N_2309);
and U2927 (N_2927,N_2048,N_1909);
and U2928 (N_2928,N_1916,N_2190);
nand U2929 (N_2929,N_1983,N_1938);
and U2930 (N_2930,N_2330,N_1943);
nor U2931 (N_2931,N_2064,N_1888);
nor U2932 (N_2932,N_1905,N_2238);
or U2933 (N_2933,N_2281,N_1876);
and U2934 (N_2934,N_2154,N_1804);
nor U2935 (N_2935,N_2326,N_1854);
nand U2936 (N_2936,N_1855,N_2222);
nand U2937 (N_2937,N_2352,N_2288);
and U2938 (N_2938,N_2022,N_1937);
nor U2939 (N_2939,N_2307,N_2121);
nand U2940 (N_2940,N_2301,N_2356);
or U2941 (N_2941,N_2318,N_2183);
and U2942 (N_2942,N_1803,N_2328);
or U2943 (N_2943,N_2154,N_2262);
xnor U2944 (N_2944,N_1942,N_1879);
and U2945 (N_2945,N_1878,N_2002);
nand U2946 (N_2946,N_2391,N_2171);
nand U2947 (N_2947,N_2051,N_2208);
and U2948 (N_2948,N_2174,N_2258);
nor U2949 (N_2949,N_2070,N_2058);
and U2950 (N_2950,N_1825,N_1914);
nand U2951 (N_2951,N_2169,N_1922);
or U2952 (N_2952,N_1869,N_2290);
and U2953 (N_2953,N_2315,N_2144);
nor U2954 (N_2954,N_2128,N_2259);
nand U2955 (N_2955,N_2036,N_1871);
and U2956 (N_2956,N_1878,N_1933);
nor U2957 (N_2957,N_1883,N_2242);
nor U2958 (N_2958,N_2226,N_1869);
or U2959 (N_2959,N_2382,N_2196);
and U2960 (N_2960,N_2210,N_2338);
and U2961 (N_2961,N_2342,N_2097);
or U2962 (N_2962,N_2092,N_2366);
or U2963 (N_2963,N_2140,N_1883);
nand U2964 (N_2964,N_2096,N_2297);
and U2965 (N_2965,N_1915,N_1992);
nor U2966 (N_2966,N_1882,N_1938);
or U2967 (N_2967,N_1941,N_2381);
and U2968 (N_2968,N_2024,N_2080);
nand U2969 (N_2969,N_2205,N_2143);
nor U2970 (N_2970,N_2020,N_2155);
and U2971 (N_2971,N_1979,N_1977);
nand U2972 (N_2972,N_2025,N_2266);
nand U2973 (N_2973,N_2128,N_2088);
or U2974 (N_2974,N_2095,N_2328);
or U2975 (N_2975,N_2334,N_2324);
nand U2976 (N_2976,N_2389,N_2260);
nand U2977 (N_2977,N_2091,N_2124);
and U2978 (N_2978,N_2124,N_2356);
and U2979 (N_2979,N_2179,N_2030);
nand U2980 (N_2980,N_2065,N_2364);
or U2981 (N_2981,N_1803,N_1976);
or U2982 (N_2982,N_2163,N_2103);
nand U2983 (N_2983,N_1902,N_1900);
or U2984 (N_2984,N_2272,N_2379);
nand U2985 (N_2985,N_2248,N_2333);
nand U2986 (N_2986,N_1811,N_2344);
and U2987 (N_2987,N_2319,N_1955);
nor U2988 (N_2988,N_2221,N_2337);
nand U2989 (N_2989,N_1822,N_2072);
and U2990 (N_2990,N_2092,N_2000);
and U2991 (N_2991,N_1831,N_1941);
nand U2992 (N_2992,N_1873,N_2201);
and U2993 (N_2993,N_2387,N_2326);
or U2994 (N_2994,N_2197,N_1881);
or U2995 (N_2995,N_2025,N_1810);
and U2996 (N_2996,N_2055,N_2090);
and U2997 (N_2997,N_1988,N_2347);
and U2998 (N_2998,N_2303,N_1941);
nand U2999 (N_2999,N_2037,N_2288);
or UO_0 (O_0,N_2918,N_2958);
and UO_1 (O_1,N_2940,N_2661);
or UO_2 (O_2,N_2517,N_2637);
nand UO_3 (O_3,N_2675,N_2410);
or UO_4 (O_4,N_2719,N_2501);
nor UO_5 (O_5,N_2638,N_2980);
nor UO_6 (O_6,N_2869,N_2960);
nor UO_7 (O_7,N_2685,N_2690);
nor UO_8 (O_8,N_2926,N_2424);
and UO_9 (O_9,N_2512,N_2497);
and UO_10 (O_10,N_2809,N_2911);
or UO_11 (O_11,N_2444,N_2561);
or UO_12 (O_12,N_2913,N_2624);
nand UO_13 (O_13,N_2851,N_2936);
nand UO_14 (O_14,N_2578,N_2852);
nand UO_15 (O_15,N_2982,N_2710);
nand UO_16 (O_16,N_2562,N_2871);
nand UO_17 (O_17,N_2589,N_2432);
nor UO_18 (O_18,N_2555,N_2664);
or UO_19 (O_19,N_2845,N_2567);
and UO_20 (O_20,N_2588,N_2819);
nand UO_21 (O_21,N_2486,N_2440);
and UO_22 (O_22,N_2471,N_2993);
and UO_23 (O_23,N_2459,N_2916);
nor UO_24 (O_24,N_2468,N_2969);
nor UO_25 (O_25,N_2726,N_2981);
nand UO_26 (O_26,N_2507,N_2447);
and UO_27 (O_27,N_2673,N_2811);
nand UO_28 (O_28,N_2566,N_2884);
nand UO_29 (O_29,N_2504,N_2438);
nand UO_30 (O_30,N_2650,N_2892);
or UO_31 (O_31,N_2798,N_2735);
nand UO_32 (O_32,N_2878,N_2944);
and UO_33 (O_33,N_2672,N_2778);
and UO_34 (O_34,N_2493,N_2714);
xor UO_35 (O_35,N_2582,N_2757);
or UO_36 (O_36,N_2460,N_2708);
nor UO_37 (O_37,N_2931,N_2652);
nand UO_38 (O_38,N_2859,N_2455);
nor UO_39 (O_39,N_2956,N_2510);
and UO_40 (O_40,N_2508,N_2810);
and UO_41 (O_41,N_2671,N_2553);
or UO_42 (O_42,N_2813,N_2552);
and UO_43 (O_43,N_2540,N_2487);
and UO_44 (O_44,N_2791,N_2800);
and UO_45 (O_45,N_2985,N_2586);
and UO_46 (O_46,N_2721,N_2458);
nand UO_47 (O_47,N_2895,N_2741);
or UO_48 (O_48,N_2720,N_2979);
nor UO_49 (O_49,N_2625,N_2828);
nor UO_50 (O_50,N_2986,N_2824);
nand UO_51 (O_51,N_2584,N_2628);
nand UO_52 (O_52,N_2959,N_2491);
and UO_53 (O_53,N_2649,N_2606);
and UO_54 (O_54,N_2862,N_2593);
xnor UO_55 (O_55,N_2889,N_2678);
and UO_56 (O_56,N_2874,N_2723);
and UO_57 (O_57,N_2779,N_2974);
nor UO_58 (O_58,N_2910,N_2968);
or UO_59 (O_59,N_2818,N_2663);
nor UO_60 (O_60,N_2835,N_2743);
nor UO_61 (O_61,N_2893,N_2488);
nand UO_62 (O_62,N_2799,N_2492);
xor UO_63 (O_63,N_2914,N_2519);
or UO_64 (O_64,N_2903,N_2550);
nand UO_65 (O_65,N_2477,N_2702);
nand UO_66 (O_66,N_2500,N_2883);
and UO_67 (O_67,N_2858,N_2891);
nand UO_68 (O_68,N_2474,N_2758);
or UO_69 (O_69,N_2854,N_2546);
nor UO_70 (O_70,N_2739,N_2796);
and UO_71 (O_71,N_2937,N_2950);
nor UO_72 (O_72,N_2836,N_2676);
or UO_73 (O_73,N_2953,N_2692);
and UO_74 (O_74,N_2788,N_2912);
nand UO_75 (O_75,N_2717,N_2516);
or UO_76 (O_76,N_2404,N_2465);
or UO_77 (O_77,N_2527,N_2748);
nor UO_78 (O_78,N_2977,N_2999);
and UO_79 (O_79,N_2934,N_2882);
and UO_80 (O_80,N_2966,N_2984);
nand UO_81 (O_81,N_2700,N_2689);
nor UO_82 (O_82,N_2573,N_2595);
or UO_83 (O_83,N_2827,N_2943);
nor UO_84 (O_84,N_2420,N_2919);
and UO_85 (O_85,N_2906,N_2457);
or UO_86 (O_86,N_2876,N_2658);
and UO_87 (O_87,N_2774,N_2576);
nand UO_88 (O_88,N_2762,N_2967);
nand UO_89 (O_89,N_2536,N_2614);
and UO_90 (O_90,N_2846,N_2877);
or UO_91 (O_91,N_2954,N_2746);
and UO_92 (O_92,N_2844,N_2626);
or UO_93 (O_93,N_2814,N_2437);
nor UO_94 (O_94,N_2445,N_2840);
or UO_95 (O_95,N_2688,N_2548);
nor UO_96 (O_96,N_2598,N_2789);
nand UO_97 (O_97,N_2525,N_2764);
nand UO_98 (O_98,N_2806,N_2547);
nand UO_99 (O_99,N_2705,N_2973);
nor UO_100 (O_100,N_2795,N_2680);
nor UO_101 (O_101,N_2481,N_2489);
nor UO_102 (O_102,N_2938,N_2687);
nand UO_103 (O_103,N_2428,N_2870);
nor UO_104 (O_104,N_2434,N_2435);
and UO_105 (O_105,N_2482,N_2759);
and UO_106 (O_106,N_2599,N_2423);
nor UO_107 (O_107,N_2597,N_2528);
nor UO_108 (O_108,N_2744,N_2897);
nand UO_109 (O_109,N_2902,N_2753);
and UO_110 (O_110,N_2456,N_2802);
or UO_111 (O_111,N_2707,N_2978);
or UO_112 (O_112,N_2751,N_2767);
or UO_113 (O_113,N_2559,N_2736);
and UO_114 (O_114,N_2961,N_2472);
nand UO_115 (O_115,N_2558,N_2803);
nor UO_116 (O_116,N_2773,N_2691);
and UO_117 (O_117,N_2755,N_2752);
or UO_118 (O_118,N_2972,N_2989);
or UO_119 (O_119,N_2816,N_2453);
xor UO_120 (O_120,N_2632,N_2648);
nor UO_121 (O_121,N_2647,N_2609);
nand UO_122 (O_122,N_2679,N_2524);
or UO_123 (O_123,N_2515,N_2411);
nand UO_124 (O_124,N_2619,N_2786);
nor UO_125 (O_125,N_2740,N_2520);
nor UO_126 (O_126,N_2543,N_2905);
or UO_127 (O_127,N_2541,N_2667);
and UO_128 (O_128,N_2868,N_2831);
or UO_129 (O_129,N_2879,N_2747);
nand UO_130 (O_130,N_2815,N_2742);
nor UO_131 (O_131,N_2415,N_2670);
or UO_132 (O_132,N_2797,N_2463);
or UO_133 (O_133,N_2509,N_2793);
and UO_134 (O_134,N_2533,N_2697);
nor UO_135 (O_135,N_2544,N_2461);
nand UO_136 (O_136,N_2829,N_2448);
and UO_137 (O_137,N_2506,N_2863);
or UO_138 (O_138,N_2976,N_2724);
or UO_139 (O_139,N_2783,N_2531);
and UO_140 (O_140,N_2412,N_2514);
or UO_141 (O_141,N_2771,N_2706);
or UO_142 (O_142,N_2441,N_2769);
nor UO_143 (O_143,N_2701,N_2734);
or UO_144 (O_144,N_2718,N_2407);
and UO_145 (O_145,N_2952,N_2551);
or UO_146 (O_146,N_2821,N_2615);
or UO_147 (O_147,N_2899,N_2560);
nor UO_148 (O_148,N_2991,N_2866);
nand UO_149 (O_149,N_2569,N_2904);
nor UO_150 (O_150,N_2794,N_2674);
nor UO_151 (O_151,N_2888,N_2564);
and UO_152 (O_152,N_2669,N_2611);
or UO_153 (O_153,N_2823,N_2763);
or UO_154 (O_154,N_2430,N_2571);
nand UO_155 (O_155,N_2665,N_2402);
and UO_156 (O_156,N_2865,N_2804);
or UO_157 (O_157,N_2513,N_2900);
nand UO_158 (O_158,N_2807,N_2935);
or UO_159 (O_159,N_2403,N_2901);
nor UO_160 (O_160,N_2842,N_2429);
and UO_161 (O_161,N_2920,N_2602);
nand UO_162 (O_162,N_2565,N_2727);
and UO_163 (O_163,N_2896,N_2792);
or UO_164 (O_164,N_2532,N_2971);
or UO_165 (O_165,N_2738,N_2521);
nand UO_166 (O_166,N_2898,N_2995);
and UO_167 (O_167,N_2965,N_2612);
nand UO_168 (O_168,N_2703,N_2419);
and UO_169 (O_169,N_2923,N_2639);
and UO_170 (O_170,N_2621,N_2409);
nand UO_171 (O_171,N_2627,N_2604);
and UO_172 (O_172,N_2490,N_2522);
nor UO_173 (O_173,N_2499,N_2666);
nand UO_174 (O_174,N_2643,N_2651);
nand UO_175 (O_175,N_2603,N_2574);
nor UO_176 (O_176,N_2754,N_2885);
nor UO_177 (O_177,N_2631,N_2608);
and UO_178 (O_178,N_2822,N_2856);
and UO_179 (O_179,N_2756,N_2848);
and UO_180 (O_180,N_2535,N_2695);
and UO_181 (O_181,N_2928,N_2933);
or UO_182 (O_182,N_2817,N_2575);
nand UO_183 (O_183,N_2613,N_2715);
or UO_184 (O_184,N_2684,N_2939);
nand UO_185 (O_185,N_2677,N_2785);
nor UO_186 (O_186,N_2908,N_2750);
and UO_187 (O_187,N_2975,N_2594);
xor UO_188 (O_188,N_2915,N_2572);
and UO_189 (O_189,N_2833,N_2857);
nor UO_190 (O_190,N_2503,N_2880);
nand UO_191 (O_191,N_2787,N_2704);
and UO_192 (O_192,N_2640,N_2656);
nand UO_193 (O_193,N_2713,N_2830);
and UO_194 (O_194,N_2421,N_2997);
nand UO_195 (O_195,N_2776,N_2475);
nor UO_196 (O_196,N_2843,N_2450);
xor UO_197 (O_197,N_2653,N_2994);
nand UO_198 (O_198,N_2924,N_2860);
nand UO_199 (O_199,N_2873,N_2494);
and UO_200 (O_200,N_2849,N_2660);
nor UO_201 (O_201,N_2596,N_2655);
and UO_202 (O_202,N_2945,N_2405);
nor UO_203 (O_203,N_2847,N_2620);
nor UO_204 (O_204,N_2616,N_2505);
or UO_205 (O_205,N_2686,N_2439);
nand UO_206 (O_206,N_2478,N_2722);
nor UO_207 (O_207,N_2826,N_2964);
and UO_208 (O_208,N_2607,N_2887);
nor UO_209 (O_209,N_2837,N_2539);
or UO_210 (O_210,N_2623,N_2711);
nand UO_211 (O_211,N_2529,N_2534);
and UO_212 (O_212,N_2470,N_2443);
nor UO_213 (O_213,N_2587,N_2861);
and UO_214 (O_214,N_2600,N_2654);
nand UO_215 (O_215,N_2563,N_2983);
or UO_216 (O_216,N_2780,N_2476);
nor UO_217 (O_217,N_2641,N_2760);
nand UO_218 (O_218,N_2442,N_2962);
nor UO_219 (O_219,N_2683,N_2941);
nand UO_220 (O_220,N_2433,N_2839);
and UO_221 (O_221,N_2772,N_2728);
and UO_222 (O_222,N_2496,N_2502);
nor UO_223 (O_223,N_2484,N_2745);
nor UO_224 (O_224,N_2467,N_2580);
and UO_225 (O_225,N_2538,N_2483);
nand UO_226 (O_226,N_2462,N_2894);
nor UO_227 (O_227,N_2645,N_2733);
nand UO_228 (O_228,N_2427,N_2635);
nand UO_229 (O_229,N_2853,N_2805);
or UO_230 (O_230,N_2765,N_2622);
nand UO_231 (O_231,N_2449,N_2511);
and UO_232 (O_232,N_2955,N_2570);
or UO_233 (O_233,N_2770,N_2422);
nand UO_234 (O_234,N_2452,N_2990);
nand UO_235 (O_235,N_2694,N_2917);
or UO_236 (O_236,N_2777,N_2855);
xnor UO_237 (O_237,N_2662,N_2864);
nor UO_238 (O_238,N_2413,N_2801);
nor UO_239 (O_239,N_2545,N_2737);
nand UO_240 (O_240,N_2946,N_2479);
nor UO_241 (O_241,N_2644,N_2963);
nand UO_242 (O_242,N_2957,N_2992);
or UO_243 (O_243,N_2469,N_2581);
or UO_244 (O_244,N_2768,N_2633);
and UO_245 (O_245,N_2601,N_2832);
and UO_246 (O_246,N_2585,N_2948);
and UO_247 (O_247,N_2825,N_2922);
or UO_248 (O_248,N_2579,N_2872);
nand UO_249 (O_249,N_2929,N_2812);
or UO_250 (O_250,N_2518,N_2523);
nor UO_251 (O_251,N_2942,N_2731);
or UO_252 (O_252,N_2749,N_2947);
and UO_253 (O_253,N_2590,N_2530);
or UO_254 (O_254,N_2716,N_2698);
or UO_255 (O_255,N_2537,N_2417);
and UO_256 (O_256,N_2930,N_2886);
or UO_257 (O_257,N_2406,N_2790);
nor UO_258 (O_258,N_2425,N_2932);
nand UO_259 (O_259,N_2784,N_2473);
nand UO_260 (O_260,N_2987,N_2577);
nand UO_261 (O_261,N_2416,N_2890);
or UO_262 (O_262,N_2605,N_2668);
and UO_263 (O_263,N_2480,N_2996);
and UO_264 (O_264,N_2850,N_2634);
or UO_265 (O_265,N_2709,N_2400);
or UO_266 (O_266,N_2766,N_2998);
or UO_267 (O_267,N_2610,N_2426);
nand UO_268 (O_268,N_2408,N_2909);
and UO_269 (O_269,N_2636,N_2431);
or UO_270 (O_270,N_2949,N_2568);
nor UO_271 (O_271,N_2782,N_2925);
and UO_272 (O_272,N_2401,N_2659);
or UO_273 (O_273,N_2820,N_2951);
or UO_274 (O_274,N_2630,N_2834);
nor UO_275 (O_275,N_2542,N_2730);
nor UO_276 (O_276,N_2414,N_2841);
and UO_277 (O_277,N_2646,N_2495);
and UO_278 (O_278,N_2466,N_2875);
or UO_279 (O_279,N_2682,N_2699);
nand UO_280 (O_280,N_2927,N_2446);
nand UO_281 (O_281,N_2781,N_2554);
or UO_282 (O_282,N_2729,N_2988);
nand UO_283 (O_283,N_2454,N_2696);
nand UO_284 (O_284,N_2881,N_2693);
or UO_285 (O_285,N_2808,N_2907);
or UO_286 (O_286,N_2418,N_2712);
and UO_287 (O_287,N_2867,N_2591);
nor UO_288 (O_288,N_2657,N_2526);
nand UO_289 (O_289,N_2921,N_2642);
nand UO_290 (O_290,N_2485,N_2681);
nand UO_291 (O_291,N_2725,N_2451);
and UO_292 (O_292,N_2775,N_2592);
and UO_293 (O_293,N_2557,N_2583);
xor UO_294 (O_294,N_2618,N_2556);
nor UO_295 (O_295,N_2617,N_2970);
nand UO_296 (O_296,N_2498,N_2732);
nand UO_297 (O_297,N_2629,N_2549);
nand UO_298 (O_298,N_2464,N_2838);
and UO_299 (O_299,N_2761,N_2436);
nor UO_300 (O_300,N_2625,N_2821);
or UO_301 (O_301,N_2856,N_2817);
nor UO_302 (O_302,N_2773,N_2519);
or UO_303 (O_303,N_2779,N_2874);
nor UO_304 (O_304,N_2739,N_2493);
nor UO_305 (O_305,N_2944,N_2861);
nor UO_306 (O_306,N_2850,N_2841);
or UO_307 (O_307,N_2836,N_2872);
nand UO_308 (O_308,N_2730,N_2900);
nand UO_309 (O_309,N_2959,N_2663);
or UO_310 (O_310,N_2776,N_2872);
or UO_311 (O_311,N_2499,N_2553);
nand UO_312 (O_312,N_2431,N_2483);
nor UO_313 (O_313,N_2767,N_2499);
nor UO_314 (O_314,N_2428,N_2446);
or UO_315 (O_315,N_2596,N_2753);
nand UO_316 (O_316,N_2930,N_2480);
nand UO_317 (O_317,N_2895,N_2663);
and UO_318 (O_318,N_2449,N_2730);
nor UO_319 (O_319,N_2946,N_2449);
and UO_320 (O_320,N_2733,N_2930);
and UO_321 (O_321,N_2524,N_2583);
or UO_322 (O_322,N_2875,N_2489);
and UO_323 (O_323,N_2616,N_2597);
or UO_324 (O_324,N_2598,N_2552);
nor UO_325 (O_325,N_2996,N_2639);
or UO_326 (O_326,N_2553,N_2639);
and UO_327 (O_327,N_2521,N_2985);
nand UO_328 (O_328,N_2570,N_2874);
or UO_329 (O_329,N_2855,N_2909);
nand UO_330 (O_330,N_2774,N_2668);
or UO_331 (O_331,N_2765,N_2498);
nor UO_332 (O_332,N_2768,N_2823);
or UO_333 (O_333,N_2768,N_2931);
and UO_334 (O_334,N_2534,N_2998);
nor UO_335 (O_335,N_2811,N_2976);
and UO_336 (O_336,N_2749,N_2427);
or UO_337 (O_337,N_2899,N_2561);
nor UO_338 (O_338,N_2670,N_2751);
and UO_339 (O_339,N_2961,N_2413);
nand UO_340 (O_340,N_2514,N_2851);
nor UO_341 (O_341,N_2641,N_2777);
nand UO_342 (O_342,N_2828,N_2803);
and UO_343 (O_343,N_2567,N_2442);
or UO_344 (O_344,N_2560,N_2452);
and UO_345 (O_345,N_2418,N_2782);
or UO_346 (O_346,N_2910,N_2505);
or UO_347 (O_347,N_2863,N_2473);
nor UO_348 (O_348,N_2503,N_2501);
and UO_349 (O_349,N_2400,N_2888);
and UO_350 (O_350,N_2859,N_2960);
nand UO_351 (O_351,N_2807,N_2705);
and UO_352 (O_352,N_2544,N_2437);
nor UO_353 (O_353,N_2513,N_2525);
nand UO_354 (O_354,N_2673,N_2408);
nand UO_355 (O_355,N_2824,N_2566);
nor UO_356 (O_356,N_2506,N_2875);
nand UO_357 (O_357,N_2788,N_2868);
or UO_358 (O_358,N_2546,N_2709);
xnor UO_359 (O_359,N_2492,N_2643);
and UO_360 (O_360,N_2800,N_2694);
nand UO_361 (O_361,N_2592,N_2749);
and UO_362 (O_362,N_2442,N_2634);
nand UO_363 (O_363,N_2699,N_2546);
nand UO_364 (O_364,N_2443,N_2910);
nor UO_365 (O_365,N_2844,N_2525);
nor UO_366 (O_366,N_2613,N_2615);
or UO_367 (O_367,N_2501,N_2694);
nand UO_368 (O_368,N_2489,N_2733);
and UO_369 (O_369,N_2704,N_2768);
or UO_370 (O_370,N_2593,N_2863);
and UO_371 (O_371,N_2955,N_2556);
or UO_372 (O_372,N_2629,N_2451);
or UO_373 (O_373,N_2467,N_2879);
nand UO_374 (O_374,N_2414,N_2477);
and UO_375 (O_375,N_2431,N_2518);
nor UO_376 (O_376,N_2410,N_2593);
and UO_377 (O_377,N_2698,N_2921);
and UO_378 (O_378,N_2800,N_2643);
nand UO_379 (O_379,N_2790,N_2718);
nand UO_380 (O_380,N_2883,N_2760);
or UO_381 (O_381,N_2443,N_2464);
and UO_382 (O_382,N_2495,N_2980);
or UO_383 (O_383,N_2748,N_2833);
nor UO_384 (O_384,N_2458,N_2934);
or UO_385 (O_385,N_2487,N_2463);
nand UO_386 (O_386,N_2466,N_2767);
and UO_387 (O_387,N_2526,N_2521);
or UO_388 (O_388,N_2445,N_2874);
nand UO_389 (O_389,N_2500,N_2827);
or UO_390 (O_390,N_2680,N_2695);
and UO_391 (O_391,N_2431,N_2448);
nand UO_392 (O_392,N_2942,N_2496);
or UO_393 (O_393,N_2837,N_2864);
nand UO_394 (O_394,N_2693,N_2949);
or UO_395 (O_395,N_2624,N_2865);
nor UO_396 (O_396,N_2664,N_2458);
and UO_397 (O_397,N_2513,N_2630);
nor UO_398 (O_398,N_2880,N_2622);
nor UO_399 (O_399,N_2890,N_2659);
or UO_400 (O_400,N_2514,N_2772);
and UO_401 (O_401,N_2827,N_2799);
and UO_402 (O_402,N_2941,N_2657);
or UO_403 (O_403,N_2768,N_2473);
nor UO_404 (O_404,N_2762,N_2798);
nand UO_405 (O_405,N_2981,N_2970);
nand UO_406 (O_406,N_2903,N_2452);
or UO_407 (O_407,N_2641,N_2725);
and UO_408 (O_408,N_2531,N_2614);
nand UO_409 (O_409,N_2830,N_2690);
or UO_410 (O_410,N_2933,N_2463);
nor UO_411 (O_411,N_2889,N_2660);
nand UO_412 (O_412,N_2859,N_2562);
nand UO_413 (O_413,N_2783,N_2667);
and UO_414 (O_414,N_2663,N_2964);
or UO_415 (O_415,N_2631,N_2985);
nor UO_416 (O_416,N_2679,N_2876);
nor UO_417 (O_417,N_2592,N_2565);
or UO_418 (O_418,N_2589,N_2856);
nor UO_419 (O_419,N_2585,N_2964);
or UO_420 (O_420,N_2673,N_2752);
nor UO_421 (O_421,N_2465,N_2767);
nand UO_422 (O_422,N_2459,N_2588);
and UO_423 (O_423,N_2991,N_2995);
nand UO_424 (O_424,N_2476,N_2901);
nand UO_425 (O_425,N_2408,N_2449);
nor UO_426 (O_426,N_2797,N_2527);
or UO_427 (O_427,N_2630,N_2562);
nand UO_428 (O_428,N_2769,N_2566);
nor UO_429 (O_429,N_2599,N_2752);
or UO_430 (O_430,N_2417,N_2660);
nor UO_431 (O_431,N_2887,N_2434);
nand UO_432 (O_432,N_2566,N_2687);
nor UO_433 (O_433,N_2797,N_2877);
or UO_434 (O_434,N_2547,N_2765);
or UO_435 (O_435,N_2425,N_2974);
nand UO_436 (O_436,N_2621,N_2836);
nand UO_437 (O_437,N_2626,N_2965);
nand UO_438 (O_438,N_2545,N_2542);
or UO_439 (O_439,N_2861,N_2743);
or UO_440 (O_440,N_2700,N_2810);
nor UO_441 (O_441,N_2599,N_2407);
xor UO_442 (O_442,N_2600,N_2511);
nand UO_443 (O_443,N_2918,N_2541);
or UO_444 (O_444,N_2535,N_2530);
nand UO_445 (O_445,N_2828,N_2887);
and UO_446 (O_446,N_2534,N_2417);
and UO_447 (O_447,N_2619,N_2455);
nand UO_448 (O_448,N_2854,N_2564);
nand UO_449 (O_449,N_2424,N_2723);
nor UO_450 (O_450,N_2533,N_2683);
nand UO_451 (O_451,N_2691,N_2514);
nor UO_452 (O_452,N_2893,N_2708);
and UO_453 (O_453,N_2889,N_2771);
and UO_454 (O_454,N_2547,N_2636);
and UO_455 (O_455,N_2945,N_2609);
and UO_456 (O_456,N_2835,N_2586);
nand UO_457 (O_457,N_2748,N_2988);
nor UO_458 (O_458,N_2831,N_2634);
nor UO_459 (O_459,N_2629,N_2659);
and UO_460 (O_460,N_2606,N_2862);
and UO_461 (O_461,N_2745,N_2738);
xor UO_462 (O_462,N_2458,N_2933);
nor UO_463 (O_463,N_2531,N_2618);
nand UO_464 (O_464,N_2553,N_2731);
nor UO_465 (O_465,N_2469,N_2473);
nor UO_466 (O_466,N_2517,N_2405);
nand UO_467 (O_467,N_2531,N_2716);
and UO_468 (O_468,N_2401,N_2530);
nand UO_469 (O_469,N_2752,N_2976);
nor UO_470 (O_470,N_2924,N_2629);
and UO_471 (O_471,N_2433,N_2873);
or UO_472 (O_472,N_2476,N_2678);
or UO_473 (O_473,N_2490,N_2813);
and UO_474 (O_474,N_2622,N_2981);
nor UO_475 (O_475,N_2759,N_2713);
nand UO_476 (O_476,N_2948,N_2939);
nor UO_477 (O_477,N_2935,N_2952);
nor UO_478 (O_478,N_2583,N_2554);
and UO_479 (O_479,N_2764,N_2858);
nand UO_480 (O_480,N_2653,N_2840);
and UO_481 (O_481,N_2906,N_2691);
and UO_482 (O_482,N_2695,N_2981);
nand UO_483 (O_483,N_2678,N_2918);
nand UO_484 (O_484,N_2635,N_2613);
or UO_485 (O_485,N_2791,N_2866);
nor UO_486 (O_486,N_2730,N_2756);
nor UO_487 (O_487,N_2483,N_2733);
nand UO_488 (O_488,N_2523,N_2407);
and UO_489 (O_489,N_2790,N_2599);
nand UO_490 (O_490,N_2497,N_2804);
and UO_491 (O_491,N_2559,N_2916);
nand UO_492 (O_492,N_2705,N_2658);
nand UO_493 (O_493,N_2796,N_2912);
nor UO_494 (O_494,N_2546,N_2487);
and UO_495 (O_495,N_2810,N_2551);
nor UO_496 (O_496,N_2968,N_2963);
or UO_497 (O_497,N_2547,N_2962);
nand UO_498 (O_498,N_2570,N_2882);
and UO_499 (O_499,N_2722,N_2872);
endmodule