module basic_500_3000_500_3_levels_2xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_402,In_4);
nor U1 (N_1,In_363,In_449);
or U2 (N_2,In_114,In_460);
and U3 (N_3,In_134,In_39);
or U4 (N_4,In_283,In_0);
nand U5 (N_5,In_172,In_33);
or U6 (N_6,In_259,In_35);
nor U7 (N_7,In_173,In_121);
nor U8 (N_8,In_346,In_365);
and U9 (N_9,In_44,In_196);
nand U10 (N_10,In_429,In_455);
nand U11 (N_11,In_438,In_395);
and U12 (N_12,In_339,In_267);
nor U13 (N_13,In_465,In_381);
and U14 (N_14,In_499,In_80);
nor U15 (N_15,In_146,In_190);
nor U16 (N_16,In_397,In_11);
or U17 (N_17,In_481,In_21);
nor U18 (N_18,In_32,In_239);
nand U19 (N_19,In_355,In_137);
or U20 (N_20,In_435,In_99);
or U21 (N_21,In_153,In_468);
xnor U22 (N_22,In_15,In_305);
nor U23 (N_23,In_463,In_231);
and U24 (N_24,In_191,In_171);
nor U25 (N_25,In_150,In_333);
xnor U26 (N_26,In_492,In_45);
xnor U27 (N_27,In_314,In_88);
and U28 (N_28,In_442,In_386);
nand U29 (N_29,In_81,In_12);
or U30 (N_30,In_170,In_467);
nand U31 (N_31,In_222,In_70);
nand U32 (N_32,In_295,In_49);
and U33 (N_33,In_14,In_252);
and U34 (N_34,In_477,In_92);
nand U35 (N_35,In_73,In_421);
nor U36 (N_36,In_459,In_243);
and U37 (N_37,In_303,In_330);
or U38 (N_38,In_215,In_338);
nand U39 (N_39,In_423,In_250);
or U40 (N_40,In_65,In_50);
nand U41 (N_41,In_228,In_51);
or U42 (N_42,In_127,In_199);
nand U43 (N_43,In_85,In_206);
or U44 (N_44,In_307,In_36);
nand U45 (N_45,In_203,In_59);
nor U46 (N_46,In_147,In_213);
or U47 (N_47,In_361,In_7);
nor U48 (N_48,In_25,In_289);
nand U49 (N_49,In_141,In_389);
nand U50 (N_50,In_123,In_388);
and U51 (N_51,In_42,In_223);
nor U52 (N_52,In_322,In_122);
nor U53 (N_53,In_238,In_376);
and U54 (N_54,In_72,In_362);
and U55 (N_55,In_226,In_68);
nand U56 (N_56,In_282,In_277);
or U57 (N_57,In_497,In_176);
nand U58 (N_58,In_292,In_247);
and U59 (N_59,In_62,In_240);
or U60 (N_60,In_107,In_23);
nor U61 (N_61,In_251,In_270);
xnor U62 (N_62,In_149,In_374);
nand U63 (N_63,In_271,In_380);
nand U64 (N_64,In_230,In_418);
and U65 (N_65,In_445,In_168);
or U66 (N_66,In_464,In_93);
and U67 (N_67,In_186,In_323);
nor U68 (N_68,In_76,In_400);
xor U69 (N_69,In_201,In_350);
nand U70 (N_70,In_111,In_331);
nor U71 (N_71,In_103,In_2);
or U72 (N_72,In_46,In_155);
nor U73 (N_73,In_372,In_87);
and U74 (N_74,In_74,In_135);
or U75 (N_75,In_288,In_124);
and U76 (N_76,In_353,In_443);
nand U77 (N_77,In_382,In_404);
or U78 (N_78,In_356,In_145);
or U79 (N_79,In_370,In_472);
or U80 (N_80,In_364,In_379);
or U81 (N_81,In_258,In_345);
nor U82 (N_82,In_242,In_433);
and U83 (N_83,In_491,In_120);
nand U84 (N_84,In_131,In_84);
nand U85 (N_85,In_58,In_496);
and U86 (N_86,In_428,In_478);
or U87 (N_87,In_66,In_318);
or U88 (N_88,In_280,In_426);
nor U89 (N_89,In_95,In_440);
nor U90 (N_90,In_479,In_408);
or U91 (N_91,In_244,In_470);
or U92 (N_92,In_476,In_174);
nand U93 (N_93,In_393,In_325);
nor U94 (N_94,In_102,In_184);
nand U95 (N_95,In_47,In_105);
and U96 (N_96,In_490,In_96);
nand U97 (N_97,In_90,In_216);
or U98 (N_98,In_471,In_351);
nand U99 (N_99,In_129,In_461);
nand U100 (N_100,In_125,In_20);
and U101 (N_101,In_304,In_52);
and U102 (N_102,In_281,In_229);
nor U103 (N_103,In_316,In_197);
nand U104 (N_104,In_117,In_448);
nor U105 (N_105,In_326,In_101);
or U106 (N_106,In_63,In_83);
nand U107 (N_107,In_276,In_274);
nor U108 (N_108,In_13,In_157);
or U109 (N_109,In_446,In_236);
or U110 (N_110,In_451,In_246);
nand U111 (N_111,In_148,In_377);
or U112 (N_112,In_284,In_82);
or U113 (N_113,In_118,In_86);
nand U114 (N_114,In_248,In_112);
and U115 (N_115,In_352,In_432);
and U116 (N_116,In_38,In_291);
or U117 (N_117,In_427,In_218);
or U118 (N_118,In_34,In_452);
or U119 (N_119,In_6,In_385);
nand U120 (N_120,In_165,In_412);
nand U121 (N_121,In_132,In_55);
nand U122 (N_122,In_27,In_209);
or U123 (N_123,In_108,In_224);
nor U124 (N_124,In_268,In_489);
or U125 (N_125,In_5,In_475);
nor U126 (N_126,In_275,In_293);
nor U127 (N_127,In_177,In_369);
nand U128 (N_128,In_24,In_329);
nand U129 (N_129,In_140,In_371);
nand U130 (N_130,In_312,In_344);
nand U131 (N_131,In_302,In_205);
nor U132 (N_132,In_8,In_91);
and U133 (N_133,In_384,In_431);
nor U134 (N_134,In_269,In_306);
nor U135 (N_135,In_211,In_57);
nand U136 (N_136,In_41,In_130);
or U137 (N_137,In_253,In_387);
nor U138 (N_138,In_1,In_208);
nand U139 (N_139,In_128,In_437);
nor U140 (N_140,In_336,In_233);
and U141 (N_141,In_430,In_398);
or U142 (N_142,In_286,In_417);
or U143 (N_143,In_100,In_152);
xnor U144 (N_144,In_488,In_214);
nand U145 (N_145,In_410,In_237);
nor U146 (N_146,In_444,In_401);
nor U147 (N_147,In_309,In_494);
or U148 (N_148,In_313,In_56);
or U149 (N_149,In_343,In_285);
and U150 (N_150,In_77,In_200);
and U151 (N_151,In_225,In_354);
or U152 (N_152,In_469,In_278);
nand U153 (N_153,In_487,In_392);
nand U154 (N_154,In_78,In_71);
nor U155 (N_155,In_405,In_424);
nand U156 (N_156,In_144,In_109);
nor U157 (N_157,In_166,In_181);
or U158 (N_158,In_28,In_358);
and U159 (N_159,In_61,In_195);
nand U160 (N_160,In_198,In_31);
xnor U161 (N_161,In_337,In_255);
and U162 (N_162,In_413,In_169);
and U163 (N_163,In_217,In_30);
and U164 (N_164,In_220,In_160);
and U165 (N_165,In_17,In_64);
nand U166 (N_166,In_115,In_232);
nor U167 (N_167,In_441,In_320);
nor U168 (N_168,In_422,In_447);
nor U169 (N_169,In_334,In_94);
nor U170 (N_170,In_335,In_415);
and U171 (N_171,In_324,In_368);
nor U172 (N_172,In_332,In_263);
nand U173 (N_173,In_245,In_484);
nor U174 (N_174,In_416,In_19);
nor U175 (N_175,In_187,In_79);
nand U176 (N_176,In_486,In_182);
or U177 (N_177,In_254,In_297);
nand U178 (N_178,In_425,In_167);
and U179 (N_179,In_194,In_498);
nand U180 (N_180,In_18,In_357);
nor U181 (N_181,In_414,In_298);
nand U182 (N_182,In_189,In_360);
nor U183 (N_183,In_378,In_212);
nor U184 (N_184,In_391,In_396);
or U185 (N_185,In_164,In_375);
nor U186 (N_186,In_261,In_299);
and U187 (N_187,In_266,In_383);
or U188 (N_188,In_180,In_342);
nor U189 (N_189,In_257,In_290);
and U190 (N_190,In_106,In_495);
or U191 (N_191,In_406,In_359);
and U192 (N_192,In_156,In_485);
and U193 (N_193,In_188,In_29);
and U194 (N_194,In_399,In_48);
xnor U195 (N_195,In_256,In_183);
nor U196 (N_196,In_458,In_462);
and U197 (N_197,In_116,In_138);
and U198 (N_198,In_53,In_221);
and U199 (N_199,In_202,In_294);
nor U200 (N_200,In_69,In_192);
and U201 (N_201,In_453,In_234);
or U202 (N_202,In_133,In_67);
nand U203 (N_203,In_411,In_193);
nor U204 (N_204,In_119,In_210);
nor U205 (N_205,In_151,In_262);
and U206 (N_206,In_439,In_450);
or U207 (N_207,In_419,In_394);
and U208 (N_208,In_436,In_473);
or U209 (N_209,In_178,In_272);
and U210 (N_210,In_493,In_301);
nand U211 (N_211,In_403,In_227);
nand U212 (N_212,In_235,In_311);
nor U213 (N_213,In_139,In_319);
nand U214 (N_214,In_40,In_300);
and U215 (N_215,In_296,In_241);
nand U216 (N_216,In_273,In_154);
nor U217 (N_217,In_287,In_420);
nand U218 (N_218,In_315,In_457);
nor U219 (N_219,In_207,In_113);
or U220 (N_220,In_264,In_22);
xor U221 (N_221,In_179,In_474);
nand U222 (N_222,In_328,In_482);
and U223 (N_223,In_43,In_483);
nor U224 (N_224,In_104,In_407);
and U225 (N_225,In_366,In_466);
and U226 (N_226,In_456,In_260);
and U227 (N_227,In_390,In_163);
nor U228 (N_228,In_136,In_373);
nand U229 (N_229,In_310,In_162);
nor U230 (N_230,In_367,In_409);
nand U231 (N_231,In_161,In_16);
nand U232 (N_232,In_89,In_175);
xnor U233 (N_233,In_110,In_204);
and U234 (N_234,In_54,In_185);
and U235 (N_235,In_321,In_98);
nor U236 (N_236,In_480,In_279);
nor U237 (N_237,In_142,In_60);
and U238 (N_238,In_158,In_265);
and U239 (N_239,In_10,In_327);
nor U240 (N_240,In_37,In_126);
xor U241 (N_241,In_9,In_219);
or U242 (N_242,In_97,In_143);
and U243 (N_243,In_308,In_317);
or U244 (N_244,In_348,In_434);
or U245 (N_245,In_159,In_26);
or U246 (N_246,In_75,In_341);
and U247 (N_247,In_249,In_340);
nor U248 (N_248,In_349,In_3);
and U249 (N_249,In_347,In_454);
or U250 (N_250,In_400,In_337);
nor U251 (N_251,In_143,In_123);
nor U252 (N_252,In_376,In_370);
and U253 (N_253,In_63,In_60);
or U254 (N_254,In_74,In_4);
nor U255 (N_255,In_257,In_446);
or U256 (N_256,In_107,In_425);
and U257 (N_257,In_253,In_391);
and U258 (N_258,In_438,In_348);
or U259 (N_259,In_70,In_232);
nand U260 (N_260,In_427,In_429);
nor U261 (N_261,In_339,In_248);
and U262 (N_262,In_62,In_448);
or U263 (N_263,In_93,In_126);
and U264 (N_264,In_421,In_320);
and U265 (N_265,In_189,In_185);
nor U266 (N_266,In_479,In_40);
and U267 (N_267,In_114,In_329);
and U268 (N_268,In_498,In_379);
or U269 (N_269,In_190,In_426);
or U270 (N_270,In_372,In_83);
or U271 (N_271,In_162,In_317);
and U272 (N_272,In_456,In_445);
nand U273 (N_273,In_346,In_193);
nand U274 (N_274,In_200,In_310);
nand U275 (N_275,In_338,In_39);
nand U276 (N_276,In_257,In_75);
or U277 (N_277,In_453,In_431);
nor U278 (N_278,In_79,In_467);
nor U279 (N_279,In_93,In_286);
or U280 (N_280,In_421,In_304);
nor U281 (N_281,In_16,In_429);
and U282 (N_282,In_299,In_401);
xor U283 (N_283,In_444,In_387);
nor U284 (N_284,In_405,In_208);
nor U285 (N_285,In_385,In_244);
nand U286 (N_286,In_497,In_227);
or U287 (N_287,In_443,In_102);
nand U288 (N_288,In_239,In_347);
and U289 (N_289,In_329,In_59);
nor U290 (N_290,In_329,In_71);
and U291 (N_291,In_312,In_75);
nor U292 (N_292,In_334,In_171);
nand U293 (N_293,In_442,In_109);
xor U294 (N_294,In_173,In_20);
nand U295 (N_295,In_311,In_322);
or U296 (N_296,In_88,In_373);
or U297 (N_297,In_7,In_269);
nor U298 (N_298,In_258,In_138);
nand U299 (N_299,In_114,In_401);
nand U300 (N_300,In_189,In_316);
or U301 (N_301,In_94,In_52);
nand U302 (N_302,In_200,In_393);
nand U303 (N_303,In_216,In_22);
nand U304 (N_304,In_121,In_88);
xnor U305 (N_305,In_225,In_203);
nor U306 (N_306,In_319,In_216);
nand U307 (N_307,In_191,In_316);
nand U308 (N_308,In_358,In_267);
or U309 (N_309,In_46,In_210);
or U310 (N_310,In_34,In_297);
and U311 (N_311,In_244,In_255);
nor U312 (N_312,In_283,In_412);
nand U313 (N_313,In_379,In_386);
nand U314 (N_314,In_25,In_142);
and U315 (N_315,In_294,In_375);
and U316 (N_316,In_25,In_89);
nand U317 (N_317,In_92,In_425);
or U318 (N_318,In_40,In_464);
and U319 (N_319,In_248,In_431);
and U320 (N_320,In_484,In_86);
and U321 (N_321,In_348,In_229);
nor U322 (N_322,In_490,In_416);
and U323 (N_323,In_479,In_54);
nor U324 (N_324,In_78,In_461);
nand U325 (N_325,In_63,In_446);
nor U326 (N_326,In_97,In_396);
nand U327 (N_327,In_397,In_362);
nand U328 (N_328,In_141,In_87);
nor U329 (N_329,In_291,In_452);
nand U330 (N_330,In_357,In_483);
nor U331 (N_331,In_300,In_276);
nor U332 (N_332,In_386,In_69);
and U333 (N_333,In_113,In_309);
xor U334 (N_334,In_299,In_109);
nand U335 (N_335,In_418,In_311);
nand U336 (N_336,In_457,In_433);
nor U337 (N_337,In_310,In_135);
nor U338 (N_338,In_183,In_422);
nand U339 (N_339,In_253,In_45);
and U340 (N_340,In_45,In_213);
and U341 (N_341,In_40,In_150);
nand U342 (N_342,In_102,In_275);
nor U343 (N_343,In_146,In_489);
or U344 (N_344,In_200,In_169);
nand U345 (N_345,In_462,In_454);
nor U346 (N_346,In_133,In_426);
or U347 (N_347,In_384,In_392);
or U348 (N_348,In_3,In_196);
nand U349 (N_349,In_87,In_171);
nand U350 (N_350,In_275,In_268);
nand U351 (N_351,In_89,In_321);
nor U352 (N_352,In_121,In_482);
and U353 (N_353,In_39,In_377);
and U354 (N_354,In_162,In_495);
nand U355 (N_355,In_169,In_147);
and U356 (N_356,In_95,In_317);
and U357 (N_357,In_37,In_213);
or U358 (N_358,In_438,In_360);
and U359 (N_359,In_230,In_188);
nor U360 (N_360,In_15,In_30);
nand U361 (N_361,In_299,In_134);
and U362 (N_362,In_316,In_257);
xor U363 (N_363,In_228,In_166);
or U364 (N_364,In_242,In_225);
and U365 (N_365,In_73,In_456);
nor U366 (N_366,In_499,In_347);
and U367 (N_367,In_463,In_230);
nor U368 (N_368,In_415,In_206);
and U369 (N_369,In_397,In_271);
nor U370 (N_370,In_311,In_228);
nor U371 (N_371,In_126,In_163);
or U372 (N_372,In_194,In_109);
or U373 (N_373,In_118,In_93);
nor U374 (N_374,In_30,In_76);
nand U375 (N_375,In_107,In_291);
and U376 (N_376,In_353,In_319);
nand U377 (N_377,In_303,In_488);
or U378 (N_378,In_328,In_188);
and U379 (N_379,In_44,In_387);
or U380 (N_380,In_195,In_307);
and U381 (N_381,In_414,In_123);
nor U382 (N_382,In_240,In_41);
nand U383 (N_383,In_25,In_306);
and U384 (N_384,In_180,In_487);
or U385 (N_385,In_104,In_29);
nor U386 (N_386,In_303,In_31);
nand U387 (N_387,In_264,In_439);
nor U388 (N_388,In_288,In_488);
nor U389 (N_389,In_161,In_85);
and U390 (N_390,In_215,In_303);
nor U391 (N_391,In_397,In_19);
nor U392 (N_392,In_80,In_319);
and U393 (N_393,In_496,In_22);
nor U394 (N_394,In_124,In_341);
nand U395 (N_395,In_390,In_170);
nor U396 (N_396,In_480,In_76);
nand U397 (N_397,In_271,In_331);
and U398 (N_398,In_42,In_227);
nand U399 (N_399,In_55,In_134);
or U400 (N_400,In_136,In_409);
nor U401 (N_401,In_265,In_383);
nand U402 (N_402,In_56,In_453);
nor U403 (N_403,In_468,In_268);
and U404 (N_404,In_350,In_409);
nor U405 (N_405,In_107,In_225);
and U406 (N_406,In_19,In_91);
or U407 (N_407,In_400,In_426);
and U408 (N_408,In_443,In_171);
nor U409 (N_409,In_41,In_455);
nor U410 (N_410,In_211,In_274);
nor U411 (N_411,In_438,In_23);
and U412 (N_412,In_170,In_403);
and U413 (N_413,In_295,In_39);
nand U414 (N_414,In_71,In_477);
and U415 (N_415,In_163,In_263);
xnor U416 (N_416,In_30,In_74);
nor U417 (N_417,In_42,In_183);
nor U418 (N_418,In_323,In_111);
and U419 (N_419,In_279,In_223);
nor U420 (N_420,In_84,In_379);
nor U421 (N_421,In_467,In_421);
nor U422 (N_422,In_43,In_194);
or U423 (N_423,In_35,In_150);
or U424 (N_424,In_16,In_254);
and U425 (N_425,In_156,In_345);
nor U426 (N_426,In_456,In_412);
xnor U427 (N_427,In_495,In_412);
and U428 (N_428,In_279,In_38);
and U429 (N_429,In_497,In_317);
and U430 (N_430,In_222,In_307);
or U431 (N_431,In_456,In_140);
nand U432 (N_432,In_162,In_219);
and U433 (N_433,In_377,In_192);
or U434 (N_434,In_51,In_239);
and U435 (N_435,In_350,In_71);
or U436 (N_436,In_148,In_245);
nor U437 (N_437,In_41,In_115);
or U438 (N_438,In_284,In_366);
or U439 (N_439,In_254,In_74);
and U440 (N_440,In_491,In_393);
nand U441 (N_441,In_49,In_108);
or U442 (N_442,In_378,In_90);
and U443 (N_443,In_221,In_486);
nor U444 (N_444,In_11,In_386);
nand U445 (N_445,In_308,In_457);
or U446 (N_446,In_233,In_191);
and U447 (N_447,In_357,In_45);
or U448 (N_448,In_230,In_29);
or U449 (N_449,In_238,In_189);
and U450 (N_450,In_284,In_14);
or U451 (N_451,In_390,In_293);
or U452 (N_452,In_433,In_14);
or U453 (N_453,In_387,In_134);
and U454 (N_454,In_114,In_373);
or U455 (N_455,In_174,In_194);
or U456 (N_456,In_494,In_289);
nor U457 (N_457,In_48,In_301);
and U458 (N_458,In_276,In_120);
nand U459 (N_459,In_26,In_348);
nand U460 (N_460,In_424,In_108);
nand U461 (N_461,In_393,In_414);
nand U462 (N_462,In_65,In_228);
and U463 (N_463,In_298,In_371);
xor U464 (N_464,In_26,In_37);
or U465 (N_465,In_280,In_449);
nand U466 (N_466,In_121,In_236);
nand U467 (N_467,In_4,In_431);
nand U468 (N_468,In_302,In_110);
and U469 (N_469,In_458,In_31);
nor U470 (N_470,In_495,In_393);
nand U471 (N_471,In_179,In_177);
xnor U472 (N_472,In_236,In_29);
nand U473 (N_473,In_444,In_183);
nor U474 (N_474,In_264,In_231);
nor U475 (N_475,In_131,In_235);
or U476 (N_476,In_267,In_236);
nand U477 (N_477,In_471,In_107);
or U478 (N_478,In_254,In_491);
nand U479 (N_479,In_497,In_220);
nand U480 (N_480,In_213,In_412);
xor U481 (N_481,In_275,In_492);
or U482 (N_482,In_41,In_223);
and U483 (N_483,In_303,In_254);
nor U484 (N_484,In_86,In_30);
and U485 (N_485,In_383,In_20);
nor U486 (N_486,In_84,In_17);
or U487 (N_487,In_168,In_263);
nor U488 (N_488,In_69,In_11);
and U489 (N_489,In_366,In_195);
xnor U490 (N_490,In_371,In_345);
nand U491 (N_491,In_210,In_146);
nor U492 (N_492,In_138,In_489);
and U493 (N_493,In_238,In_362);
or U494 (N_494,In_255,In_463);
nor U495 (N_495,In_59,In_102);
xor U496 (N_496,In_409,In_327);
and U497 (N_497,In_33,In_407);
and U498 (N_498,In_184,In_178);
nor U499 (N_499,In_102,In_271);
and U500 (N_500,In_42,In_94);
and U501 (N_501,In_133,In_160);
nor U502 (N_502,In_157,In_287);
and U503 (N_503,In_44,In_334);
nor U504 (N_504,In_376,In_166);
or U505 (N_505,In_53,In_463);
nand U506 (N_506,In_56,In_189);
nand U507 (N_507,In_437,In_38);
and U508 (N_508,In_287,In_485);
or U509 (N_509,In_128,In_452);
or U510 (N_510,In_453,In_255);
nor U511 (N_511,In_307,In_486);
and U512 (N_512,In_15,In_287);
and U513 (N_513,In_338,In_292);
or U514 (N_514,In_60,In_334);
or U515 (N_515,In_156,In_399);
and U516 (N_516,In_160,In_167);
nand U517 (N_517,In_457,In_28);
or U518 (N_518,In_172,In_278);
and U519 (N_519,In_422,In_209);
or U520 (N_520,In_32,In_49);
nand U521 (N_521,In_97,In_333);
or U522 (N_522,In_96,In_383);
or U523 (N_523,In_3,In_297);
nor U524 (N_524,In_30,In_226);
nor U525 (N_525,In_135,In_168);
and U526 (N_526,In_258,In_23);
nand U527 (N_527,In_245,In_493);
and U528 (N_528,In_159,In_494);
nand U529 (N_529,In_294,In_275);
or U530 (N_530,In_37,In_387);
or U531 (N_531,In_118,In_99);
nand U532 (N_532,In_22,In_197);
or U533 (N_533,In_384,In_234);
or U534 (N_534,In_92,In_1);
and U535 (N_535,In_429,In_136);
nand U536 (N_536,In_233,In_188);
nand U537 (N_537,In_213,In_78);
nor U538 (N_538,In_1,In_124);
and U539 (N_539,In_196,In_311);
nand U540 (N_540,In_409,In_42);
and U541 (N_541,In_447,In_184);
nand U542 (N_542,In_356,In_468);
nand U543 (N_543,In_451,In_281);
nor U544 (N_544,In_252,In_108);
and U545 (N_545,In_457,In_497);
nand U546 (N_546,In_485,In_487);
nand U547 (N_547,In_312,In_490);
or U548 (N_548,In_282,In_157);
nand U549 (N_549,In_472,In_84);
or U550 (N_550,In_300,In_345);
nand U551 (N_551,In_183,In_26);
nor U552 (N_552,In_294,In_86);
nor U553 (N_553,In_448,In_178);
nor U554 (N_554,In_241,In_103);
nand U555 (N_555,In_19,In_58);
or U556 (N_556,In_23,In_175);
nor U557 (N_557,In_42,In_384);
nand U558 (N_558,In_267,In_235);
or U559 (N_559,In_63,In_12);
and U560 (N_560,In_237,In_471);
xor U561 (N_561,In_4,In_452);
and U562 (N_562,In_307,In_431);
xnor U563 (N_563,In_2,In_343);
nand U564 (N_564,In_478,In_148);
nor U565 (N_565,In_266,In_93);
and U566 (N_566,In_17,In_21);
or U567 (N_567,In_199,In_204);
and U568 (N_568,In_81,In_41);
nor U569 (N_569,In_327,In_94);
nor U570 (N_570,In_455,In_193);
or U571 (N_571,In_301,In_131);
nand U572 (N_572,In_338,In_184);
nand U573 (N_573,In_494,In_218);
and U574 (N_574,In_178,In_287);
and U575 (N_575,In_484,In_201);
nand U576 (N_576,In_9,In_496);
xnor U577 (N_577,In_488,In_126);
or U578 (N_578,In_80,In_139);
and U579 (N_579,In_250,In_135);
and U580 (N_580,In_461,In_472);
nand U581 (N_581,In_330,In_275);
and U582 (N_582,In_268,In_385);
and U583 (N_583,In_198,In_494);
nor U584 (N_584,In_244,In_460);
xnor U585 (N_585,In_449,In_394);
or U586 (N_586,In_488,In_431);
nand U587 (N_587,In_158,In_448);
and U588 (N_588,In_194,In_444);
nand U589 (N_589,In_39,In_323);
and U590 (N_590,In_14,In_270);
nor U591 (N_591,In_241,In_356);
or U592 (N_592,In_359,In_135);
nand U593 (N_593,In_404,In_367);
nand U594 (N_594,In_227,In_176);
nor U595 (N_595,In_74,In_16);
nand U596 (N_596,In_439,In_133);
nor U597 (N_597,In_162,In_31);
xor U598 (N_598,In_333,In_481);
xnor U599 (N_599,In_407,In_227);
and U600 (N_600,In_461,In_327);
or U601 (N_601,In_36,In_205);
or U602 (N_602,In_193,In_0);
and U603 (N_603,In_223,In_340);
nor U604 (N_604,In_264,In_45);
nand U605 (N_605,In_370,In_330);
nor U606 (N_606,In_382,In_305);
and U607 (N_607,In_381,In_371);
nor U608 (N_608,In_384,In_430);
nand U609 (N_609,In_187,In_6);
nand U610 (N_610,In_70,In_339);
nand U611 (N_611,In_146,In_157);
nand U612 (N_612,In_497,In_3);
nand U613 (N_613,In_146,In_98);
nand U614 (N_614,In_194,In_268);
or U615 (N_615,In_47,In_250);
and U616 (N_616,In_187,In_262);
nand U617 (N_617,In_306,In_347);
nor U618 (N_618,In_339,In_17);
nor U619 (N_619,In_399,In_384);
and U620 (N_620,In_134,In_166);
nor U621 (N_621,In_218,In_2);
nor U622 (N_622,In_6,In_388);
or U623 (N_623,In_469,In_443);
and U624 (N_624,In_257,In_86);
xor U625 (N_625,In_61,In_44);
nand U626 (N_626,In_351,In_433);
nor U627 (N_627,In_408,In_325);
or U628 (N_628,In_461,In_269);
xor U629 (N_629,In_121,In_101);
and U630 (N_630,In_114,In_407);
nor U631 (N_631,In_415,In_138);
and U632 (N_632,In_447,In_201);
nand U633 (N_633,In_130,In_212);
and U634 (N_634,In_173,In_278);
and U635 (N_635,In_202,In_89);
and U636 (N_636,In_262,In_38);
nor U637 (N_637,In_357,In_332);
and U638 (N_638,In_6,In_282);
nand U639 (N_639,In_171,In_496);
nand U640 (N_640,In_491,In_182);
or U641 (N_641,In_382,In_45);
nand U642 (N_642,In_241,In_149);
and U643 (N_643,In_173,In_306);
nor U644 (N_644,In_385,In_391);
nand U645 (N_645,In_385,In_483);
nand U646 (N_646,In_0,In_371);
or U647 (N_647,In_424,In_76);
nand U648 (N_648,In_320,In_448);
and U649 (N_649,In_212,In_361);
nand U650 (N_650,In_51,In_224);
nor U651 (N_651,In_228,In_198);
or U652 (N_652,In_175,In_437);
and U653 (N_653,In_288,In_37);
nor U654 (N_654,In_292,In_427);
nand U655 (N_655,In_105,In_438);
nor U656 (N_656,In_434,In_59);
or U657 (N_657,In_168,In_96);
or U658 (N_658,In_78,In_246);
or U659 (N_659,In_389,In_72);
nand U660 (N_660,In_81,In_362);
nor U661 (N_661,In_208,In_110);
or U662 (N_662,In_292,In_336);
nand U663 (N_663,In_59,In_430);
and U664 (N_664,In_136,In_130);
xor U665 (N_665,In_94,In_254);
or U666 (N_666,In_486,In_10);
nand U667 (N_667,In_291,In_46);
nand U668 (N_668,In_242,In_381);
and U669 (N_669,In_149,In_115);
xor U670 (N_670,In_188,In_451);
or U671 (N_671,In_158,In_324);
nand U672 (N_672,In_269,In_51);
nor U673 (N_673,In_321,In_431);
nand U674 (N_674,In_488,In_45);
nand U675 (N_675,In_444,In_368);
xnor U676 (N_676,In_185,In_225);
nor U677 (N_677,In_424,In_217);
nor U678 (N_678,In_348,In_310);
and U679 (N_679,In_252,In_260);
and U680 (N_680,In_353,In_63);
nand U681 (N_681,In_4,In_289);
and U682 (N_682,In_8,In_63);
nand U683 (N_683,In_214,In_409);
xnor U684 (N_684,In_183,In_383);
or U685 (N_685,In_303,In_3);
nand U686 (N_686,In_415,In_120);
nand U687 (N_687,In_443,In_160);
nand U688 (N_688,In_106,In_63);
nand U689 (N_689,In_123,In_126);
and U690 (N_690,In_144,In_72);
and U691 (N_691,In_151,In_274);
nand U692 (N_692,In_474,In_72);
nor U693 (N_693,In_365,In_23);
nand U694 (N_694,In_354,In_375);
nor U695 (N_695,In_125,In_68);
nand U696 (N_696,In_423,In_350);
nor U697 (N_697,In_393,In_211);
nor U698 (N_698,In_376,In_50);
or U699 (N_699,In_417,In_413);
nand U700 (N_700,In_455,In_142);
and U701 (N_701,In_311,In_126);
nor U702 (N_702,In_108,In_93);
nand U703 (N_703,In_378,In_442);
nand U704 (N_704,In_348,In_131);
or U705 (N_705,In_16,In_68);
or U706 (N_706,In_453,In_289);
nor U707 (N_707,In_223,In_488);
or U708 (N_708,In_203,In_412);
nor U709 (N_709,In_18,In_178);
and U710 (N_710,In_415,In_347);
nor U711 (N_711,In_173,In_314);
nand U712 (N_712,In_448,In_428);
or U713 (N_713,In_348,In_285);
nand U714 (N_714,In_471,In_326);
nor U715 (N_715,In_460,In_142);
or U716 (N_716,In_394,In_492);
nand U717 (N_717,In_222,In_362);
nor U718 (N_718,In_432,In_464);
and U719 (N_719,In_441,In_344);
nand U720 (N_720,In_244,In_299);
nand U721 (N_721,In_446,In_228);
or U722 (N_722,In_288,In_328);
nor U723 (N_723,In_400,In_249);
or U724 (N_724,In_91,In_106);
nand U725 (N_725,In_480,In_494);
xor U726 (N_726,In_385,In_464);
and U727 (N_727,In_61,In_132);
nor U728 (N_728,In_71,In_333);
and U729 (N_729,In_49,In_497);
nand U730 (N_730,In_496,In_439);
nand U731 (N_731,In_211,In_353);
and U732 (N_732,In_38,In_95);
nand U733 (N_733,In_108,In_324);
or U734 (N_734,In_309,In_205);
and U735 (N_735,In_387,In_363);
and U736 (N_736,In_107,In_273);
nand U737 (N_737,In_62,In_340);
or U738 (N_738,In_408,In_316);
and U739 (N_739,In_354,In_328);
nor U740 (N_740,In_147,In_499);
nor U741 (N_741,In_153,In_188);
or U742 (N_742,In_377,In_85);
or U743 (N_743,In_212,In_381);
xor U744 (N_744,In_269,In_158);
and U745 (N_745,In_93,In_24);
nand U746 (N_746,In_262,In_142);
nor U747 (N_747,In_15,In_327);
or U748 (N_748,In_47,In_36);
nor U749 (N_749,In_99,In_416);
xor U750 (N_750,In_15,In_88);
and U751 (N_751,In_56,In_124);
or U752 (N_752,In_290,In_232);
nand U753 (N_753,In_92,In_499);
and U754 (N_754,In_142,In_489);
or U755 (N_755,In_29,In_98);
nor U756 (N_756,In_285,In_360);
or U757 (N_757,In_259,In_171);
or U758 (N_758,In_200,In_254);
nor U759 (N_759,In_91,In_277);
nor U760 (N_760,In_343,In_106);
or U761 (N_761,In_310,In_20);
or U762 (N_762,In_397,In_261);
nand U763 (N_763,In_321,In_191);
and U764 (N_764,In_156,In_433);
nand U765 (N_765,In_482,In_369);
and U766 (N_766,In_366,In_216);
and U767 (N_767,In_335,In_2);
or U768 (N_768,In_441,In_190);
nor U769 (N_769,In_364,In_435);
nor U770 (N_770,In_43,In_434);
nor U771 (N_771,In_175,In_411);
nand U772 (N_772,In_117,In_436);
nor U773 (N_773,In_393,In_432);
and U774 (N_774,In_341,In_308);
and U775 (N_775,In_108,In_439);
nand U776 (N_776,In_212,In_87);
and U777 (N_777,In_60,In_113);
and U778 (N_778,In_79,In_477);
or U779 (N_779,In_291,In_347);
and U780 (N_780,In_386,In_49);
or U781 (N_781,In_293,In_4);
or U782 (N_782,In_155,In_148);
xnor U783 (N_783,In_130,In_4);
nand U784 (N_784,In_469,In_196);
nor U785 (N_785,In_352,In_336);
xor U786 (N_786,In_297,In_141);
and U787 (N_787,In_176,In_37);
and U788 (N_788,In_494,In_374);
nand U789 (N_789,In_14,In_387);
and U790 (N_790,In_43,In_354);
or U791 (N_791,In_105,In_485);
and U792 (N_792,In_26,In_342);
and U793 (N_793,In_86,In_11);
nand U794 (N_794,In_145,In_237);
nand U795 (N_795,In_419,In_222);
and U796 (N_796,In_322,In_291);
nor U797 (N_797,In_434,In_361);
nor U798 (N_798,In_282,In_140);
and U799 (N_799,In_247,In_273);
and U800 (N_800,In_255,In_329);
nor U801 (N_801,In_429,In_336);
nand U802 (N_802,In_407,In_318);
nand U803 (N_803,In_297,In_480);
or U804 (N_804,In_473,In_359);
and U805 (N_805,In_3,In_201);
or U806 (N_806,In_497,In_230);
nand U807 (N_807,In_325,In_215);
nor U808 (N_808,In_50,In_326);
nand U809 (N_809,In_233,In_278);
xor U810 (N_810,In_56,In_90);
and U811 (N_811,In_481,In_419);
or U812 (N_812,In_471,In_186);
xor U813 (N_813,In_178,In_399);
or U814 (N_814,In_20,In_144);
nor U815 (N_815,In_268,In_395);
and U816 (N_816,In_23,In_112);
or U817 (N_817,In_28,In_411);
and U818 (N_818,In_234,In_258);
nand U819 (N_819,In_115,In_453);
and U820 (N_820,In_179,In_151);
nor U821 (N_821,In_92,In_403);
and U822 (N_822,In_72,In_388);
or U823 (N_823,In_254,In_314);
nand U824 (N_824,In_493,In_134);
nand U825 (N_825,In_423,In_192);
and U826 (N_826,In_421,In_371);
nand U827 (N_827,In_117,In_102);
nand U828 (N_828,In_178,In_298);
nor U829 (N_829,In_379,In_44);
nor U830 (N_830,In_79,In_199);
and U831 (N_831,In_430,In_71);
and U832 (N_832,In_243,In_269);
and U833 (N_833,In_124,In_80);
and U834 (N_834,In_453,In_344);
or U835 (N_835,In_239,In_245);
nor U836 (N_836,In_175,In_219);
or U837 (N_837,In_474,In_113);
nor U838 (N_838,In_484,In_154);
nand U839 (N_839,In_118,In_261);
xor U840 (N_840,In_360,In_495);
nor U841 (N_841,In_418,In_135);
and U842 (N_842,In_307,In_336);
nand U843 (N_843,In_460,In_360);
or U844 (N_844,In_141,In_217);
or U845 (N_845,In_189,In_255);
nand U846 (N_846,In_265,In_452);
and U847 (N_847,In_494,In_465);
or U848 (N_848,In_144,In_335);
nor U849 (N_849,In_102,In_189);
nor U850 (N_850,In_346,In_94);
nor U851 (N_851,In_380,In_221);
or U852 (N_852,In_395,In_288);
xnor U853 (N_853,In_135,In_457);
and U854 (N_854,In_158,In_429);
nand U855 (N_855,In_56,In_187);
nand U856 (N_856,In_395,In_149);
xnor U857 (N_857,In_188,In_18);
or U858 (N_858,In_19,In_305);
nand U859 (N_859,In_463,In_105);
nand U860 (N_860,In_363,In_190);
nand U861 (N_861,In_203,In_298);
or U862 (N_862,In_461,In_182);
nand U863 (N_863,In_441,In_494);
nand U864 (N_864,In_215,In_199);
nor U865 (N_865,In_62,In_457);
and U866 (N_866,In_463,In_349);
nand U867 (N_867,In_311,In_64);
or U868 (N_868,In_386,In_260);
nand U869 (N_869,In_337,In_461);
nand U870 (N_870,In_81,In_263);
nor U871 (N_871,In_54,In_422);
nor U872 (N_872,In_153,In_456);
or U873 (N_873,In_317,In_457);
or U874 (N_874,In_80,In_407);
nand U875 (N_875,In_498,In_290);
or U876 (N_876,In_351,In_132);
nand U877 (N_877,In_149,In_344);
or U878 (N_878,In_494,In_256);
nor U879 (N_879,In_365,In_232);
nor U880 (N_880,In_42,In_447);
nor U881 (N_881,In_232,In_406);
and U882 (N_882,In_234,In_214);
nand U883 (N_883,In_378,In_297);
or U884 (N_884,In_260,In_136);
or U885 (N_885,In_130,In_474);
nand U886 (N_886,In_5,In_321);
and U887 (N_887,In_421,In_476);
nand U888 (N_888,In_269,In_266);
nand U889 (N_889,In_454,In_55);
xnor U890 (N_890,In_73,In_306);
or U891 (N_891,In_167,In_126);
nand U892 (N_892,In_62,In_407);
or U893 (N_893,In_410,In_227);
nor U894 (N_894,In_211,In_496);
and U895 (N_895,In_229,In_262);
nand U896 (N_896,In_311,In_214);
nor U897 (N_897,In_151,In_9);
nand U898 (N_898,In_478,In_39);
and U899 (N_899,In_47,In_458);
or U900 (N_900,In_209,In_202);
xnor U901 (N_901,In_118,In_84);
and U902 (N_902,In_451,In_183);
and U903 (N_903,In_497,In_131);
and U904 (N_904,In_275,In_205);
nand U905 (N_905,In_329,In_391);
or U906 (N_906,In_173,In_420);
nor U907 (N_907,In_88,In_154);
and U908 (N_908,In_190,In_344);
nor U909 (N_909,In_476,In_60);
and U910 (N_910,In_453,In_77);
or U911 (N_911,In_97,In_497);
nor U912 (N_912,In_120,In_82);
and U913 (N_913,In_450,In_26);
nand U914 (N_914,In_192,In_185);
nor U915 (N_915,In_248,In_59);
nor U916 (N_916,In_417,In_384);
and U917 (N_917,In_443,In_238);
nand U918 (N_918,In_206,In_200);
or U919 (N_919,In_357,In_47);
nor U920 (N_920,In_393,In_328);
nand U921 (N_921,In_432,In_223);
and U922 (N_922,In_229,In_94);
nor U923 (N_923,In_67,In_76);
or U924 (N_924,In_405,In_224);
nor U925 (N_925,In_384,In_87);
nor U926 (N_926,In_477,In_72);
and U927 (N_927,In_59,In_269);
and U928 (N_928,In_354,In_251);
nand U929 (N_929,In_42,In_294);
nand U930 (N_930,In_282,In_465);
nand U931 (N_931,In_139,In_313);
nand U932 (N_932,In_390,In_113);
nand U933 (N_933,In_151,In_316);
or U934 (N_934,In_199,In_490);
or U935 (N_935,In_180,In_22);
or U936 (N_936,In_50,In_362);
and U937 (N_937,In_65,In_45);
nor U938 (N_938,In_403,In_197);
nor U939 (N_939,In_140,In_266);
nor U940 (N_940,In_411,In_278);
nor U941 (N_941,In_64,In_422);
and U942 (N_942,In_472,In_313);
nor U943 (N_943,In_438,In_384);
nor U944 (N_944,In_276,In_382);
or U945 (N_945,In_253,In_35);
nor U946 (N_946,In_358,In_280);
nor U947 (N_947,In_211,In_357);
xnor U948 (N_948,In_70,In_63);
or U949 (N_949,In_398,In_8);
nor U950 (N_950,In_189,In_287);
nor U951 (N_951,In_447,In_436);
nor U952 (N_952,In_397,In_124);
and U953 (N_953,In_256,In_377);
and U954 (N_954,In_210,In_41);
and U955 (N_955,In_348,In_295);
and U956 (N_956,In_244,In_101);
nand U957 (N_957,In_291,In_429);
nor U958 (N_958,In_196,In_165);
nor U959 (N_959,In_221,In_396);
nand U960 (N_960,In_315,In_26);
nand U961 (N_961,In_328,In_118);
nor U962 (N_962,In_455,In_170);
nand U963 (N_963,In_81,In_69);
or U964 (N_964,In_157,In_252);
or U965 (N_965,In_374,In_220);
nor U966 (N_966,In_468,In_264);
nor U967 (N_967,In_61,In_75);
nand U968 (N_968,In_465,In_56);
nand U969 (N_969,In_421,In_70);
nand U970 (N_970,In_16,In_36);
nand U971 (N_971,In_480,In_64);
or U972 (N_972,In_97,In_364);
nand U973 (N_973,In_374,In_486);
and U974 (N_974,In_15,In_94);
and U975 (N_975,In_49,In_289);
nor U976 (N_976,In_256,In_301);
and U977 (N_977,In_264,In_322);
nand U978 (N_978,In_163,In_205);
or U979 (N_979,In_295,In_460);
nand U980 (N_980,In_454,In_171);
or U981 (N_981,In_191,In_173);
and U982 (N_982,In_315,In_476);
nor U983 (N_983,In_116,In_374);
nand U984 (N_984,In_32,In_191);
nand U985 (N_985,In_210,In_138);
or U986 (N_986,In_279,In_147);
and U987 (N_987,In_205,In_457);
nor U988 (N_988,In_478,In_486);
nand U989 (N_989,In_11,In_365);
or U990 (N_990,In_196,In_115);
nand U991 (N_991,In_108,In_154);
and U992 (N_992,In_50,In_148);
and U993 (N_993,In_76,In_105);
nor U994 (N_994,In_481,In_423);
or U995 (N_995,In_268,In_464);
or U996 (N_996,In_334,In_225);
nor U997 (N_997,In_271,In_254);
and U998 (N_998,In_478,In_252);
nand U999 (N_999,In_344,In_456);
nor U1000 (N_1000,N_268,N_937);
nand U1001 (N_1001,N_958,N_178);
nand U1002 (N_1002,N_224,N_462);
nand U1003 (N_1003,N_951,N_537);
nand U1004 (N_1004,N_438,N_619);
nand U1005 (N_1005,N_857,N_750);
nand U1006 (N_1006,N_935,N_659);
nor U1007 (N_1007,N_8,N_199);
xnor U1008 (N_1008,N_501,N_23);
xor U1009 (N_1009,N_67,N_876);
nand U1010 (N_1010,N_386,N_694);
and U1011 (N_1011,N_928,N_519);
nand U1012 (N_1012,N_238,N_384);
and U1013 (N_1013,N_201,N_261);
nor U1014 (N_1014,N_861,N_258);
nand U1015 (N_1015,N_896,N_68);
or U1016 (N_1016,N_552,N_663);
or U1017 (N_1017,N_949,N_637);
and U1018 (N_1018,N_229,N_226);
and U1019 (N_1019,N_657,N_173);
and U1020 (N_1020,N_37,N_474);
and U1021 (N_1021,N_629,N_450);
or U1022 (N_1022,N_943,N_166);
and U1023 (N_1023,N_960,N_265);
and U1024 (N_1024,N_922,N_314);
and U1025 (N_1025,N_244,N_54);
or U1026 (N_1026,N_563,N_464);
or U1027 (N_1027,N_816,N_452);
nand U1028 (N_1028,N_673,N_670);
nand U1029 (N_1029,N_843,N_739);
nor U1030 (N_1030,N_203,N_284);
nor U1031 (N_1031,N_777,N_492);
and U1032 (N_1032,N_435,N_270);
or U1033 (N_1033,N_834,N_647);
nor U1034 (N_1034,N_824,N_416);
and U1035 (N_1035,N_486,N_162);
nand U1036 (N_1036,N_247,N_225);
nor U1037 (N_1037,N_798,N_551);
and U1038 (N_1038,N_421,N_16);
and U1039 (N_1039,N_65,N_323);
nor U1040 (N_1040,N_712,N_213);
or U1041 (N_1041,N_58,N_329);
nor U1042 (N_1042,N_598,N_56);
nand U1043 (N_1043,N_588,N_98);
nand U1044 (N_1044,N_195,N_782);
nor U1045 (N_1045,N_793,N_292);
and U1046 (N_1046,N_868,N_546);
nand U1047 (N_1047,N_760,N_521);
or U1048 (N_1048,N_764,N_938);
or U1049 (N_1049,N_726,N_468);
nand U1050 (N_1050,N_727,N_756);
nor U1051 (N_1051,N_794,N_560);
and U1052 (N_1052,N_887,N_221);
and U1053 (N_1053,N_456,N_274);
and U1054 (N_1054,N_736,N_628);
nor U1055 (N_1055,N_62,N_432);
or U1056 (N_1056,N_854,N_660);
nand U1057 (N_1057,N_343,N_51);
nand U1058 (N_1058,N_804,N_661);
xor U1059 (N_1059,N_605,N_174);
or U1060 (N_1060,N_543,N_484);
or U1061 (N_1061,N_495,N_441);
nor U1062 (N_1062,N_518,N_652);
nor U1063 (N_1063,N_912,N_821);
and U1064 (N_1064,N_856,N_921);
and U1065 (N_1065,N_154,N_404);
or U1066 (N_1066,N_570,N_924);
or U1067 (N_1067,N_796,N_222);
and U1068 (N_1068,N_300,N_708);
or U1069 (N_1069,N_104,N_111);
or U1070 (N_1070,N_379,N_368);
and U1071 (N_1071,N_483,N_994);
nand U1072 (N_1072,N_934,N_317);
and U1073 (N_1073,N_42,N_331);
and U1074 (N_1074,N_26,N_817);
and U1075 (N_1075,N_711,N_963);
nand U1076 (N_1076,N_237,N_360);
nor U1077 (N_1077,N_900,N_954);
and U1078 (N_1078,N_653,N_488);
nor U1079 (N_1079,N_442,N_114);
and U1080 (N_1080,N_658,N_936);
nor U1081 (N_1081,N_956,N_38);
nor U1082 (N_1082,N_401,N_291);
nand U1083 (N_1083,N_627,N_734);
nor U1084 (N_1084,N_168,N_870);
and U1085 (N_1085,N_909,N_140);
nand U1086 (N_1086,N_980,N_290);
and U1087 (N_1087,N_253,N_910);
and U1088 (N_1088,N_689,N_266);
or U1089 (N_1089,N_14,N_790);
or U1090 (N_1090,N_388,N_837);
nand U1091 (N_1091,N_57,N_828);
and U1092 (N_1092,N_152,N_403);
nor U1093 (N_1093,N_64,N_818);
or U1094 (N_1094,N_269,N_597);
nor U1095 (N_1095,N_161,N_676);
xor U1096 (N_1096,N_271,N_669);
xor U1097 (N_1097,N_467,N_443);
nor U1098 (N_1098,N_705,N_312);
nand U1099 (N_1099,N_315,N_459);
and U1100 (N_1100,N_641,N_83);
nand U1101 (N_1101,N_234,N_348);
or U1102 (N_1102,N_680,N_200);
and U1103 (N_1103,N_359,N_236);
nor U1104 (N_1104,N_378,N_585);
nand U1105 (N_1105,N_745,N_106);
and U1106 (N_1106,N_989,N_355);
nand U1107 (N_1107,N_437,N_939);
nor U1108 (N_1108,N_516,N_4);
nor U1109 (N_1109,N_394,N_541);
nor U1110 (N_1110,N_959,N_929);
nand U1111 (N_1111,N_675,N_643);
or U1112 (N_1112,N_395,N_662);
and U1113 (N_1113,N_795,N_391);
xor U1114 (N_1114,N_6,N_742);
and U1115 (N_1115,N_496,N_690);
or U1116 (N_1116,N_950,N_425);
or U1117 (N_1117,N_992,N_710);
and U1118 (N_1118,N_223,N_781);
nand U1119 (N_1119,N_393,N_376);
nand U1120 (N_1120,N_7,N_878);
and U1121 (N_1121,N_482,N_411);
nand U1122 (N_1122,N_74,N_932);
nor U1123 (N_1123,N_807,N_181);
or U1124 (N_1124,N_392,N_617);
nand U1125 (N_1125,N_449,N_681);
xnor U1126 (N_1126,N_820,N_987);
nor U1127 (N_1127,N_167,N_879);
or U1128 (N_1128,N_93,N_196);
nor U1129 (N_1129,N_502,N_888);
nand U1130 (N_1130,N_744,N_848);
nand U1131 (N_1131,N_626,N_583);
nor U1132 (N_1132,N_957,N_770);
xor U1133 (N_1133,N_228,N_122);
nor U1134 (N_1134,N_534,N_490);
or U1135 (N_1135,N_69,N_340);
nor U1136 (N_1136,N_789,N_974);
nand U1137 (N_1137,N_36,N_908);
nand U1138 (N_1138,N_723,N_354);
nor U1139 (N_1139,N_10,N_553);
nand U1140 (N_1140,N_683,N_273);
or U1141 (N_1141,N_55,N_39);
nand U1142 (N_1142,N_814,N_461);
nand U1143 (N_1143,N_249,N_549);
or U1144 (N_1144,N_574,N_264);
nor U1145 (N_1145,N_243,N_72);
nand U1146 (N_1146,N_735,N_63);
and U1147 (N_1147,N_20,N_135);
nand U1148 (N_1148,N_917,N_31);
nand U1149 (N_1149,N_651,N_990);
or U1150 (N_1150,N_907,N_721);
xor U1151 (N_1151,N_761,N_283);
nand U1152 (N_1152,N_0,N_232);
nor U1153 (N_1153,N_210,N_358);
nor U1154 (N_1154,N_170,N_594);
nor U1155 (N_1155,N_35,N_481);
and U1156 (N_1156,N_973,N_33);
nor U1157 (N_1157,N_538,N_904);
or U1158 (N_1158,N_754,N_869);
and U1159 (N_1159,N_458,N_850);
and U1160 (N_1160,N_841,N_978);
xnor U1161 (N_1161,N_645,N_382);
nor U1162 (N_1162,N_895,N_371);
or U1163 (N_1163,N_409,N_466);
nand U1164 (N_1164,N_91,N_819);
nor U1165 (N_1165,N_845,N_15);
nor U1166 (N_1166,N_916,N_127);
nor U1167 (N_1167,N_788,N_138);
nand U1168 (N_1168,N_509,N_337);
nor U1169 (N_1169,N_231,N_250);
nor U1170 (N_1170,N_457,N_11);
nand U1171 (N_1171,N_407,N_49);
nor U1172 (N_1172,N_591,N_240);
nand U1173 (N_1173,N_175,N_499);
or U1174 (N_1174,N_367,N_955);
or U1175 (N_1175,N_102,N_682);
nor U1176 (N_1176,N_695,N_76);
nor U1177 (N_1177,N_431,N_602);
or U1178 (N_1178,N_193,N_713);
and U1179 (N_1179,N_718,N_809);
nand U1180 (N_1180,N_310,N_999);
nor U1181 (N_1181,N_966,N_18);
nor U1182 (N_1182,N_732,N_630);
or U1183 (N_1183,N_307,N_863);
nand U1184 (N_1184,N_733,N_579);
and U1185 (N_1185,N_128,N_979);
or U1186 (N_1186,N_650,N_361);
nand U1187 (N_1187,N_890,N_522);
xor U1188 (N_1188,N_410,N_155);
and U1189 (N_1189,N_826,N_476);
nand U1190 (N_1190,N_498,N_478);
nor U1191 (N_1191,N_158,N_584);
xnor U1192 (N_1192,N_822,N_406);
nand U1193 (N_1193,N_515,N_147);
nor U1194 (N_1194,N_129,N_420);
xor U1195 (N_1195,N_92,N_996);
nand U1196 (N_1196,N_567,N_9);
and U1197 (N_1197,N_374,N_188);
or U1198 (N_1198,N_321,N_964);
nor U1199 (N_1199,N_387,N_728);
or U1200 (N_1200,N_202,N_740);
nor U1201 (N_1201,N_685,N_185);
nor U1202 (N_1202,N_831,N_877);
nand U1203 (N_1203,N_507,N_891);
nand U1204 (N_1204,N_328,N_245);
nand U1205 (N_1205,N_986,N_729);
and U1206 (N_1206,N_902,N_341);
and U1207 (N_1207,N_27,N_593);
nor U1208 (N_1208,N_239,N_962);
and U1209 (N_1209,N_184,N_145);
and U1210 (N_1210,N_970,N_429);
and U1211 (N_1211,N_350,N_965);
nor U1212 (N_1212,N_644,N_691);
nand U1213 (N_1213,N_302,N_527);
nor U1214 (N_1214,N_833,N_171);
nor U1215 (N_1215,N_491,N_119);
nand U1216 (N_1216,N_933,N_572);
nor U1217 (N_1217,N_859,N_306);
and U1218 (N_1218,N_194,N_768);
or U1219 (N_1219,N_299,N_634);
and U1220 (N_1220,N_977,N_717);
and U1221 (N_1221,N_415,N_852);
or U1222 (N_1222,N_326,N_827);
nor U1223 (N_1223,N_919,N_577);
nand U1224 (N_1224,N_976,N_815);
or U1225 (N_1225,N_797,N_601);
or U1226 (N_1226,N_50,N_510);
or U1227 (N_1227,N_528,N_699);
and U1228 (N_1228,N_948,N_632);
or U1229 (N_1229,N_227,N_776);
or U1230 (N_1230,N_134,N_103);
or U1231 (N_1231,N_344,N_402);
nand U1232 (N_1232,N_242,N_463);
and U1233 (N_1233,N_825,N_703);
nand U1234 (N_1234,N_767,N_30);
or U1235 (N_1235,N_79,N_260);
nand U1236 (N_1236,N_621,N_294);
nand U1237 (N_1237,N_413,N_762);
nor U1238 (N_1238,N_279,N_981);
and U1239 (N_1239,N_160,N_664);
or U1240 (N_1240,N_246,N_396);
and U1241 (N_1241,N_48,N_573);
or U1242 (N_1242,N_716,N_531);
nand U1243 (N_1243,N_338,N_561);
nand U1244 (N_1244,N_293,N_862);
or U1245 (N_1245,N_678,N_419);
nor U1246 (N_1246,N_800,N_885);
nand U1247 (N_1247,N_864,N_205);
or U1248 (N_1248,N_576,N_12);
and U1249 (N_1249,N_883,N_448);
xnor U1250 (N_1250,N_915,N_839);
nand U1251 (N_1251,N_913,N_751);
nand U1252 (N_1252,N_288,N_720);
and U1253 (N_1253,N_66,N_364);
nand U1254 (N_1254,N_29,N_640);
and U1255 (N_1255,N_749,N_947);
or U1256 (N_1256,N_882,N_143);
and U1257 (N_1257,N_305,N_285);
nor U1258 (N_1258,N_642,N_677);
nand U1259 (N_1259,N_944,N_357);
and U1260 (N_1260,N_565,N_287);
nor U1261 (N_1261,N_88,N_362);
and U1262 (N_1262,N_606,N_366);
and U1263 (N_1263,N_564,N_325);
or U1264 (N_1264,N_578,N_21);
nand U1265 (N_1265,N_748,N_757);
or U1266 (N_1266,N_13,N_556);
or U1267 (N_1267,N_150,N_286);
or U1268 (N_1268,N_94,N_803);
and U1269 (N_1269,N_596,N_82);
nand U1270 (N_1270,N_81,N_208);
or U1271 (N_1271,N_263,N_385);
nor U1272 (N_1272,N_714,N_867);
and U1273 (N_1273,N_211,N_159);
xor U1274 (N_1274,N_684,N_982);
nor U1275 (N_1275,N_164,N_536);
nand U1276 (N_1276,N_698,N_901);
nand U1277 (N_1277,N_424,N_153);
nand U1278 (N_1278,N_892,N_858);
and U1279 (N_1279,N_125,N_702);
nand U1280 (N_1280,N_779,N_755);
nor U1281 (N_1281,N_218,N_207);
nor U1282 (N_1282,N_32,N_45);
nor U1283 (N_1283,N_59,N_719);
nand U1284 (N_1284,N_470,N_961);
nand U1285 (N_1285,N_508,N_555);
nand U1286 (N_1286,N_612,N_303);
or U1287 (N_1287,N_709,N_830);
or U1288 (N_1288,N_633,N_693);
or U1289 (N_1289,N_725,N_587);
or U1290 (N_1290,N_715,N_335);
nor U1291 (N_1291,N_309,N_722);
nand U1292 (N_1292,N_524,N_176);
nor U1293 (N_1293,N_316,N_189);
and U1294 (N_1294,N_517,N_311);
or U1295 (N_1295,N_405,N_559);
nand U1296 (N_1296,N_44,N_618);
nor U1297 (N_1297,N_398,N_622);
or U1298 (N_1298,N_906,N_34);
nand U1299 (N_1299,N_875,N_631);
nand U1300 (N_1300,N_139,N_940);
nand U1301 (N_1301,N_41,N_995);
or U1302 (N_1302,N_886,N_737);
nor U1303 (N_1303,N_787,N_625);
and U1304 (N_1304,N_784,N_731);
and U1305 (N_1305,N_851,N_526);
nand U1306 (N_1306,N_997,N_453);
nor U1307 (N_1307,N_759,N_17);
or U1308 (N_1308,N_774,N_926);
nor U1309 (N_1309,N_141,N_423);
nor U1310 (N_1310,N_805,N_61);
nand U1311 (N_1311,N_430,N_636);
and U1312 (N_1312,N_783,N_212);
nor U1313 (N_1313,N_206,N_780);
or U1314 (N_1314,N_595,N_775);
nand U1315 (N_1315,N_700,N_460);
nand U1316 (N_1316,N_334,N_24);
nor U1317 (N_1317,N_513,N_897);
nor U1318 (N_1318,N_352,N_743);
and U1319 (N_1319,N_724,N_116);
and U1320 (N_1320,N_130,N_46);
or U1321 (N_1321,N_327,N_133);
nand U1322 (N_1322,N_255,N_590);
and U1323 (N_1323,N_945,N_149);
nand U1324 (N_1324,N_686,N_282);
nand U1325 (N_1325,N_151,N_22);
or U1326 (N_1326,N_972,N_198);
or U1327 (N_1327,N_773,N_77);
nor U1328 (N_1328,N_988,N_914);
and U1329 (N_1329,N_259,N_752);
nor U1330 (N_1330,N_163,N_927);
or U1331 (N_1331,N_802,N_918);
nand U1332 (N_1332,N_646,N_967);
nor U1333 (N_1333,N_489,N_746);
nor U1334 (N_1334,N_697,N_179);
nand U1335 (N_1335,N_763,N_197);
nand U1336 (N_1336,N_479,N_447);
nand U1337 (N_1337,N_330,N_97);
and U1338 (N_1338,N_165,N_373);
and U1339 (N_1339,N_581,N_254);
or U1340 (N_1340,N_298,N_860);
nor U1341 (N_1341,N_671,N_320);
and U1342 (N_1342,N_665,N_113);
nor U1343 (N_1343,N_332,N_991);
and U1344 (N_1344,N_542,N_905);
nand U1345 (N_1345,N_473,N_840);
nor U1346 (N_1346,N_248,N_28);
nand U1347 (N_1347,N_823,N_523);
or U1348 (N_1348,N_866,N_346);
and U1349 (N_1349,N_487,N_872);
or U1350 (N_1350,N_730,N_771);
nand U1351 (N_1351,N_765,N_655);
nand U1352 (N_1352,N_871,N_295);
or U1353 (N_1353,N_582,N_296);
or U1354 (N_1354,N_408,N_953);
nand U1355 (N_1355,N_575,N_614);
nor U1356 (N_1356,N_571,N_96);
or U1357 (N_1357,N_952,N_638);
and U1358 (N_1358,N_370,N_80);
nor U1359 (N_1359,N_623,N_835);
nor U1360 (N_1360,N_433,N_75);
and U1361 (N_1361,N_428,N_832);
nor U1362 (N_1362,N_532,N_799);
or U1363 (N_1363,N_566,N_984);
or U1364 (N_1364,N_512,N_183);
nor U1365 (N_1365,N_142,N_884);
or U1366 (N_1366,N_186,N_747);
nor U1367 (N_1367,N_469,N_190);
and U1368 (N_1368,N_529,N_78);
nand U1369 (N_1369,N_110,N_70);
nor U1370 (N_1370,N_345,N_514);
or U1371 (N_1371,N_898,N_108);
nand U1372 (N_1372,N_586,N_351);
and U1373 (N_1373,N_157,N_930);
nor U1374 (N_1374,N_215,N_347);
or U1375 (N_1375,N_836,N_557);
nand U1376 (N_1376,N_214,N_137);
xnor U1377 (N_1377,N_846,N_126);
nand U1378 (N_1378,N_535,N_192);
xnor U1379 (N_1379,N_440,N_889);
and U1380 (N_1380,N_19,N_639);
and U1381 (N_1381,N_687,N_117);
or U1382 (N_1382,N_84,N_118);
nand U1383 (N_1383,N_616,N_52);
xnor U1384 (N_1384,N_568,N_772);
nand U1385 (N_1385,N_672,N_187);
nand U1386 (N_1386,N_123,N_562);
xnor U1387 (N_1387,N_313,N_706);
nor U1388 (N_1388,N_297,N_112);
nor U1389 (N_1389,N_753,N_881);
nor U1390 (N_1390,N_399,N_397);
nand U1391 (N_1391,N_100,N_899);
and U1392 (N_1392,N_107,N_120);
nor U1393 (N_1393,N_946,N_390);
or U1394 (N_1394,N_607,N_504);
or U1395 (N_1395,N_599,N_25);
nor U1396 (N_1396,N_356,N_688);
xor U1397 (N_1397,N_792,N_942);
or U1398 (N_1398,N_592,N_604);
or U1399 (N_1399,N_925,N_455);
nor U1400 (N_1400,N_230,N_548);
and U1401 (N_1401,N_506,N_434);
nor U1402 (N_1402,N_380,N_3);
or U1403 (N_1403,N_668,N_1);
nor U1404 (N_1404,N_656,N_920);
and U1405 (N_1405,N_786,N_336);
or U1406 (N_1406,N_95,N_610);
nand U1407 (N_1407,N_472,N_503);
or U1408 (N_1408,N_497,N_530);
nor U1409 (N_1409,N_377,N_109);
nand U1410 (N_1410,N_806,N_2);
nor U1411 (N_1411,N_539,N_649);
and U1412 (N_1412,N_180,N_923);
nand U1413 (N_1413,N_704,N_191);
nand U1414 (N_1414,N_475,N_648);
or U1415 (N_1415,N_493,N_204);
and U1416 (N_1416,N_272,N_500);
nor U1417 (N_1417,N_275,N_445);
nor U1418 (N_1418,N_252,N_71);
nand U1419 (N_1419,N_701,N_766);
and U1420 (N_1420,N_400,N_235);
and U1421 (N_1421,N_318,N_349);
nor U1422 (N_1422,N_324,N_589);
nor U1423 (N_1423,N_47,N_417);
or U1424 (N_1424,N_547,N_545);
and U1425 (N_1425,N_741,N_267);
nand U1426 (N_1426,N_600,N_569);
nor U1427 (N_1427,N_969,N_968);
nand U1428 (N_1428,N_985,N_427);
or U1429 (N_1429,N_465,N_85);
nand U1430 (N_1430,N_115,N_679);
and U1431 (N_1431,N_73,N_148);
and U1432 (N_1432,N_131,N_847);
and U1433 (N_1433,N_666,N_865);
and U1434 (N_1434,N_485,N_209);
or U1435 (N_1435,N_304,N_635);
and U1436 (N_1436,N_785,N_480);
or U1437 (N_1437,N_389,N_422);
nor U1438 (N_1438,N_418,N_322);
nand U1439 (N_1439,N_454,N_60);
nor U1440 (N_1440,N_86,N_156);
nand U1441 (N_1441,N_121,N_558);
nor U1442 (N_1442,N_256,N_844);
nand U1443 (N_1443,N_611,N_383);
or U1444 (N_1444,N_993,N_615);
nand U1445 (N_1445,N_426,N_674);
nand U1446 (N_1446,N_608,N_280);
nand U1447 (N_1447,N_372,N_281);
nand U1448 (N_1448,N_533,N_124);
nor U1449 (N_1449,N_544,N_894);
and U1450 (N_1450,N_233,N_855);
and U1451 (N_1451,N_696,N_903);
nor U1452 (N_1452,N_778,N_177);
and U1453 (N_1453,N_182,N_811);
nand U1454 (N_1454,N_172,N_812);
nor U1455 (N_1455,N_333,N_911);
and U1456 (N_1456,N_40,N_278);
nor U1457 (N_1457,N_220,N_667);
and U1458 (N_1458,N_810,N_43);
or U1459 (N_1459,N_941,N_494);
or U1460 (N_1460,N_369,N_520);
or U1461 (N_1461,N_654,N_624);
or U1462 (N_1462,N_829,N_87);
nand U1463 (N_1463,N_89,N_216);
nor U1464 (N_1464,N_375,N_101);
nand U1465 (N_1465,N_412,N_853);
or U1466 (N_1466,N_554,N_477);
nor U1467 (N_1467,N_880,N_365);
nor U1468 (N_1468,N_319,N_241);
and U1469 (N_1469,N_219,N_105);
nand U1470 (N_1470,N_262,N_217);
or U1471 (N_1471,N_439,N_525);
nand U1472 (N_1472,N_363,N_99);
nand U1473 (N_1473,N_444,N_620);
nand U1474 (N_1474,N_707,N_813);
and U1475 (N_1475,N_692,N_136);
nor U1476 (N_1476,N_276,N_446);
nand U1477 (N_1477,N_873,N_511);
and U1478 (N_1478,N_580,N_257);
or U1479 (N_1479,N_414,N_975);
and U1480 (N_1480,N_381,N_53);
xnor U1481 (N_1481,N_277,N_849);
nor U1482 (N_1482,N_505,N_308);
or U1483 (N_1483,N_801,N_146);
xnor U1484 (N_1484,N_132,N_353);
or U1485 (N_1485,N_436,N_251);
or U1486 (N_1486,N_339,N_301);
nor U1487 (N_1487,N_603,N_738);
and U1488 (N_1488,N_931,N_471);
or U1489 (N_1489,N_90,N_769);
nand U1490 (N_1490,N_609,N_451);
or U1491 (N_1491,N_144,N_893);
and U1492 (N_1492,N_613,N_550);
nand U1493 (N_1493,N_758,N_289);
and U1494 (N_1494,N_874,N_791);
nor U1495 (N_1495,N_842,N_342);
nand U1496 (N_1496,N_998,N_808);
nand U1497 (N_1497,N_971,N_169);
nand U1498 (N_1498,N_540,N_5);
nand U1499 (N_1499,N_983,N_838);
nor U1500 (N_1500,N_943,N_355);
nand U1501 (N_1501,N_791,N_944);
nor U1502 (N_1502,N_760,N_815);
and U1503 (N_1503,N_149,N_956);
or U1504 (N_1504,N_887,N_176);
nand U1505 (N_1505,N_993,N_394);
and U1506 (N_1506,N_280,N_507);
nand U1507 (N_1507,N_25,N_493);
nand U1508 (N_1508,N_97,N_53);
nor U1509 (N_1509,N_985,N_687);
nor U1510 (N_1510,N_77,N_318);
and U1511 (N_1511,N_484,N_492);
nand U1512 (N_1512,N_941,N_610);
or U1513 (N_1513,N_338,N_907);
nand U1514 (N_1514,N_999,N_587);
or U1515 (N_1515,N_447,N_538);
and U1516 (N_1516,N_983,N_375);
nor U1517 (N_1517,N_159,N_512);
and U1518 (N_1518,N_620,N_766);
or U1519 (N_1519,N_799,N_226);
nand U1520 (N_1520,N_982,N_916);
and U1521 (N_1521,N_280,N_342);
and U1522 (N_1522,N_249,N_717);
nand U1523 (N_1523,N_128,N_850);
nand U1524 (N_1524,N_643,N_706);
and U1525 (N_1525,N_255,N_166);
or U1526 (N_1526,N_529,N_467);
nand U1527 (N_1527,N_70,N_335);
nor U1528 (N_1528,N_427,N_865);
xnor U1529 (N_1529,N_418,N_798);
nor U1530 (N_1530,N_344,N_980);
and U1531 (N_1531,N_993,N_539);
or U1532 (N_1532,N_732,N_465);
xnor U1533 (N_1533,N_68,N_627);
nor U1534 (N_1534,N_37,N_241);
or U1535 (N_1535,N_448,N_320);
nand U1536 (N_1536,N_470,N_784);
and U1537 (N_1537,N_564,N_768);
nand U1538 (N_1538,N_116,N_684);
nand U1539 (N_1539,N_68,N_334);
or U1540 (N_1540,N_91,N_146);
nand U1541 (N_1541,N_62,N_706);
and U1542 (N_1542,N_86,N_138);
nand U1543 (N_1543,N_908,N_326);
or U1544 (N_1544,N_899,N_225);
nor U1545 (N_1545,N_29,N_13);
nor U1546 (N_1546,N_618,N_612);
and U1547 (N_1547,N_731,N_801);
or U1548 (N_1548,N_692,N_540);
nor U1549 (N_1549,N_226,N_783);
nand U1550 (N_1550,N_381,N_738);
nand U1551 (N_1551,N_738,N_184);
and U1552 (N_1552,N_172,N_514);
nand U1553 (N_1553,N_699,N_727);
and U1554 (N_1554,N_272,N_813);
or U1555 (N_1555,N_634,N_412);
and U1556 (N_1556,N_789,N_90);
nand U1557 (N_1557,N_298,N_917);
nor U1558 (N_1558,N_682,N_594);
and U1559 (N_1559,N_156,N_816);
nand U1560 (N_1560,N_654,N_989);
or U1561 (N_1561,N_390,N_458);
xor U1562 (N_1562,N_76,N_629);
nor U1563 (N_1563,N_413,N_201);
nand U1564 (N_1564,N_599,N_264);
nor U1565 (N_1565,N_252,N_221);
or U1566 (N_1566,N_4,N_849);
and U1567 (N_1567,N_487,N_121);
nand U1568 (N_1568,N_99,N_780);
and U1569 (N_1569,N_764,N_950);
or U1570 (N_1570,N_36,N_940);
nand U1571 (N_1571,N_119,N_482);
xor U1572 (N_1572,N_241,N_23);
and U1573 (N_1573,N_985,N_939);
nor U1574 (N_1574,N_364,N_24);
and U1575 (N_1575,N_61,N_517);
and U1576 (N_1576,N_419,N_803);
or U1577 (N_1577,N_148,N_471);
nand U1578 (N_1578,N_218,N_372);
nand U1579 (N_1579,N_450,N_919);
and U1580 (N_1580,N_629,N_231);
nor U1581 (N_1581,N_230,N_314);
and U1582 (N_1582,N_978,N_380);
and U1583 (N_1583,N_727,N_312);
or U1584 (N_1584,N_382,N_784);
and U1585 (N_1585,N_396,N_658);
nor U1586 (N_1586,N_871,N_600);
and U1587 (N_1587,N_900,N_798);
nor U1588 (N_1588,N_787,N_970);
nor U1589 (N_1589,N_175,N_14);
xnor U1590 (N_1590,N_894,N_341);
and U1591 (N_1591,N_991,N_40);
or U1592 (N_1592,N_876,N_339);
or U1593 (N_1593,N_491,N_268);
and U1594 (N_1594,N_20,N_701);
or U1595 (N_1595,N_471,N_586);
nand U1596 (N_1596,N_814,N_737);
and U1597 (N_1597,N_866,N_909);
or U1598 (N_1598,N_785,N_803);
or U1599 (N_1599,N_541,N_763);
nor U1600 (N_1600,N_758,N_916);
or U1601 (N_1601,N_169,N_516);
nor U1602 (N_1602,N_14,N_290);
nor U1603 (N_1603,N_468,N_399);
nand U1604 (N_1604,N_760,N_118);
nand U1605 (N_1605,N_104,N_833);
nor U1606 (N_1606,N_969,N_197);
or U1607 (N_1607,N_835,N_934);
and U1608 (N_1608,N_358,N_597);
nor U1609 (N_1609,N_683,N_567);
nor U1610 (N_1610,N_14,N_984);
nand U1611 (N_1611,N_629,N_285);
or U1612 (N_1612,N_394,N_910);
and U1613 (N_1613,N_314,N_228);
nor U1614 (N_1614,N_240,N_767);
nand U1615 (N_1615,N_974,N_581);
xnor U1616 (N_1616,N_290,N_181);
and U1617 (N_1617,N_9,N_948);
nor U1618 (N_1618,N_153,N_288);
nand U1619 (N_1619,N_837,N_737);
nor U1620 (N_1620,N_966,N_887);
or U1621 (N_1621,N_878,N_422);
nor U1622 (N_1622,N_956,N_641);
nand U1623 (N_1623,N_774,N_839);
or U1624 (N_1624,N_612,N_166);
nand U1625 (N_1625,N_604,N_730);
nand U1626 (N_1626,N_71,N_208);
or U1627 (N_1627,N_13,N_863);
or U1628 (N_1628,N_10,N_467);
and U1629 (N_1629,N_350,N_617);
or U1630 (N_1630,N_388,N_300);
or U1631 (N_1631,N_744,N_15);
nor U1632 (N_1632,N_111,N_919);
nand U1633 (N_1633,N_294,N_614);
nand U1634 (N_1634,N_140,N_617);
and U1635 (N_1635,N_673,N_779);
or U1636 (N_1636,N_15,N_914);
nand U1637 (N_1637,N_850,N_594);
and U1638 (N_1638,N_118,N_248);
or U1639 (N_1639,N_640,N_228);
or U1640 (N_1640,N_458,N_145);
and U1641 (N_1641,N_250,N_52);
xor U1642 (N_1642,N_533,N_749);
nand U1643 (N_1643,N_800,N_646);
and U1644 (N_1644,N_187,N_161);
and U1645 (N_1645,N_427,N_343);
and U1646 (N_1646,N_306,N_907);
or U1647 (N_1647,N_812,N_10);
nor U1648 (N_1648,N_803,N_776);
or U1649 (N_1649,N_615,N_118);
or U1650 (N_1650,N_947,N_296);
nand U1651 (N_1651,N_854,N_849);
nand U1652 (N_1652,N_458,N_403);
nor U1653 (N_1653,N_125,N_273);
and U1654 (N_1654,N_557,N_952);
nor U1655 (N_1655,N_941,N_389);
and U1656 (N_1656,N_329,N_845);
or U1657 (N_1657,N_404,N_908);
nand U1658 (N_1658,N_303,N_297);
xnor U1659 (N_1659,N_368,N_776);
and U1660 (N_1660,N_970,N_964);
and U1661 (N_1661,N_75,N_112);
nor U1662 (N_1662,N_648,N_983);
nand U1663 (N_1663,N_246,N_985);
nor U1664 (N_1664,N_760,N_886);
and U1665 (N_1665,N_495,N_252);
or U1666 (N_1666,N_474,N_151);
nand U1667 (N_1667,N_480,N_432);
nor U1668 (N_1668,N_787,N_174);
nor U1669 (N_1669,N_333,N_930);
or U1670 (N_1670,N_56,N_425);
or U1671 (N_1671,N_999,N_70);
nor U1672 (N_1672,N_285,N_112);
nor U1673 (N_1673,N_77,N_394);
or U1674 (N_1674,N_104,N_949);
or U1675 (N_1675,N_849,N_423);
nand U1676 (N_1676,N_182,N_643);
nor U1677 (N_1677,N_167,N_752);
and U1678 (N_1678,N_578,N_77);
nand U1679 (N_1679,N_195,N_442);
and U1680 (N_1680,N_663,N_392);
nand U1681 (N_1681,N_522,N_276);
and U1682 (N_1682,N_660,N_286);
and U1683 (N_1683,N_248,N_351);
nor U1684 (N_1684,N_276,N_47);
and U1685 (N_1685,N_691,N_762);
or U1686 (N_1686,N_699,N_550);
or U1687 (N_1687,N_445,N_667);
and U1688 (N_1688,N_928,N_121);
nand U1689 (N_1689,N_569,N_252);
or U1690 (N_1690,N_828,N_178);
or U1691 (N_1691,N_584,N_513);
nand U1692 (N_1692,N_455,N_321);
or U1693 (N_1693,N_889,N_644);
nor U1694 (N_1694,N_631,N_434);
or U1695 (N_1695,N_100,N_923);
and U1696 (N_1696,N_318,N_950);
or U1697 (N_1697,N_921,N_886);
nor U1698 (N_1698,N_275,N_473);
or U1699 (N_1699,N_38,N_263);
or U1700 (N_1700,N_69,N_965);
or U1701 (N_1701,N_846,N_520);
or U1702 (N_1702,N_379,N_811);
or U1703 (N_1703,N_105,N_484);
nand U1704 (N_1704,N_785,N_343);
nand U1705 (N_1705,N_407,N_883);
and U1706 (N_1706,N_541,N_518);
or U1707 (N_1707,N_823,N_543);
nand U1708 (N_1708,N_257,N_299);
nand U1709 (N_1709,N_256,N_252);
and U1710 (N_1710,N_459,N_661);
and U1711 (N_1711,N_632,N_408);
or U1712 (N_1712,N_680,N_425);
nand U1713 (N_1713,N_737,N_478);
xor U1714 (N_1714,N_654,N_992);
nor U1715 (N_1715,N_901,N_457);
nand U1716 (N_1716,N_319,N_580);
nor U1717 (N_1717,N_417,N_228);
nor U1718 (N_1718,N_619,N_735);
or U1719 (N_1719,N_104,N_933);
and U1720 (N_1720,N_837,N_948);
and U1721 (N_1721,N_970,N_918);
nor U1722 (N_1722,N_330,N_194);
and U1723 (N_1723,N_194,N_671);
nand U1724 (N_1724,N_804,N_653);
nor U1725 (N_1725,N_404,N_581);
and U1726 (N_1726,N_94,N_535);
or U1727 (N_1727,N_10,N_172);
and U1728 (N_1728,N_566,N_821);
nand U1729 (N_1729,N_716,N_698);
nor U1730 (N_1730,N_813,N_496);
nand U1731 (N_1731,N_555,N_417);
nor U1732 (N_1732,N_489,N_473);
or U1733 (N_1733,N_642,N_934);
nand U1734 (N_1734,N_844,N_700);
nand U1735 (N_1735,N_523,N_562);
or U1736 (N_1736,N_924,N_936);
nor U1737 (N_1737,N_990,N_656);
and U1738 (N_1738,N_145,N_571);
nand U1739 (N_1739,N_528,N_397);
or U1740 (N_1740,N_279,N_76);
nor U1741 (N_1741,N_931,N_766);
nand U1742 (N_1742,N_6,N_368);
nor U1743 (N_1743,N_577,N_892);
nand U1744 (N_1744,N_728,N_54);
nor U1745 (N_1745,N_765,N_882);
or U1746 (N_1746,N_788,N_940);
nor U1747 (N_1747,N_494,N_984);
xor U1748 (N_1748,N_743,N_708);
xnor U1749 (N_1749,N_758,N_209);
and U1750 (N_1750,N_413,N_775);
and U1751 (N_1751,N_120,N_646);
nor U1752 (N_1752,N_234,N_196);
and U1753 (N_1753,N_762,N_867);
nor U1754 (N_1754,N_147,N_750);
nor U1755 (N_1755,N_887,N_573);
nor U1756 (N_1756,N_777,N_86);
and U1757 (N_1757,N_629,N_68);
nand U1758 (N_1758,N_936,N_706);
or U1759 (N_1759,N_765,N_752);
nor U1760 (N_1760,N_270,N_929);
or U1761 (N_1761,N_237,N_167);
nand U1762 (N_1762,N_488,N_176);
xnor U1763 (N_1763,N_32,N_908);
and U1764 (N_1764,N_166,N_502);
nor U1765 (N_1765,N_603,N_288);
nor U1766 (N_1766,N_354,N_275);
xor U1767 (N_1767,N_919,N_641);
nand U1768 (N_1768,N_579,N_222);
nand U1769 (N_1769,N_127,N_943);
and U1770 (N_1770,N_302,N_201);
nand U1771 (N_1771,N_248,N_697);
or U1772 (N_1772,N_890,N_19);
nor U1773 (N_1773,N_532,N_971);
nor U1774 (N_1774,N_603,N_712);
nor U1775 (N_1775,N_366,N_741);
nand U1776 (N_1776,N_880,N_940);
and U1777 (N_1777,N_391,N_208);
or U1778 (N_1778,N_299,N_679);
and U1779 (N_1779,N_912,N_37);
nand U1780 (N_1780,N_235,N_362);
and U1781 (N_1781,N_439,N_906);
or U1782 (N_1782,N_648,N_883);
xor U1783 (N_1783,N_24,N_80);
and U1784 (N_1784,N_808,N_91);
or U1785 (N_1785,N_973,N_300);
and U1786 (N_1786,N_809,N_246);
and U1787 (N_1787,N_163,N_915);
or U1788 (N_1788,N_82,N_926);
nor U1789 (N_1789,N_395,N_540);
and U1790 (N_1790,N_432,N_797);
nand U1791 (N_1791,N_228,N_595);
and U1792 (N_1792,N_630,N_661);
or U1793 (N_1793,N_620,N_451);
nand U1794 (N_1794,N_382,N_141);
nor U1795 (N_1795,N_437,N_979);
or U1796 (N_1796,N_813,N_693);
nand U1797 (N_1797,N_705,N_744);
and U1798 (N_1798,N_956,N_251);
or U1799 (N_1799,N_523,N_94);
and U1800 (N_1800,N_817,N_202);
nor U1801 (N_1801,N_422,N_194);
nand U1802 (N_1802,N_75,N_12);
nor U1803 (N_1803,N_570,N_236);
or U1804 (N_1804,N_31,N_223);
or U1805 (N_1805,N_514,N_790);
nand U1806 (N_1806,N_902,N_896);
nand U1807 (N_1807,N_933,N_595);
and U1808 (N_1808,N_603,N_694);
and U1809 (N_1809,N_827,N_740);
and U1810 (N_1810,N_675,N_925);
and U1811 (N_1811,N_180,N_413);
nor U1812 (N_1812,N_615,N_794);
and U1813 (N_1813,N_330,N_615);
or U1814 (N_1814,N_551,N_198);
or U1815 (N_1815,N_922,N_895);
nand U1816 (N_1816,N_969,N_699);
nor U1817 (N_1817,N_485,N_925);
nand U1818 (N_1818,N_745,N_312);
or U1819 (N_1819,N_486,N_427);
nand U1820 (N_1820,N_106,N_43);
nor U1821 (N_1821,N_50,N_402);
or U1822 (N_1822,N_781,N_138);
or U1823 (N_1823,N_123,N_583);
nand U1824 (N_1824,N_763,N_757);
nor U1825 (N_1825,N_80,N_1);
nor U1826 (N_1826,N_235,N_216);
nand U1827 (N_1827,N_427,N_396);
and U1828 (N_1828,N_686,N_102);
nor U1829 (N_1829,N_376,N_908);
xnor U1830 (N_1830,N_454,N_681);
nand U1831 (N_1831,N_595,N_91);
and U1832 (N_1832,N_110,N_815);
and U1833 (N_1833,N_851,N_273);
nand U1834 (N_1834,N_184,N_71);
nor U1835 (N_1835,N_982,N_113);
and U1836 (N_1836,N_610,N_453);
or U1837 (N_1837,N_177,N_815);
nor U1838 (N_1838,N_240,N_533);
nand U1839 (N_1839,N_580,N_391);
or U1840 (N_1840,N_545,N_63);
and U1841 (N_1841,N_388,N_536);
or U1842 (N_1842,N_934,N_713);
nor U1843 (N_1843,N_763,N_126);
or U1844 (N_1844,N_339,N_4);
or U1845 (N_1845,N_553,N_547);
nor U1846 (N_1846,N_423,N_995);
or U1847 (N_1847,N_952,N_68);
nand U1848 (N_1848,N_824,N_529);
and U1849 (N_1849,N_657,N_457);
xnor U1850 (N_1850,N_177,N_781);
nand U1851 (N_1851,N_890,N_415);
and U1852 (N_1852,N_864,N_791);
or U1853 (N_1853,N_790,N_71);
or U1854 (N_1854,N_841,N_273);
and U1855 (N_1855,N_511,N_485);
and U1856 (N_1856,N_679,N_773);
nor U1857 (N_1857,N_824,N_882);
nand U1858 (N_1858,N_677,N_77);
or U1859 (N_1859,N_752,N_231);
and U1860 (N_1860,N_960,N_448);
and U1861 (N_1861,N_239,N_975);
xnor U1862 (N_1862,N_393,N_859);
nand U1863 (N_1863,N_961,N_549);
nand U1864 (N_1864,N_437,N_894);
or U1865 (N_1865,N_712,N_68);
or U1866 (N_1866,N_465,N_789);
or U1867 (N_1867,N_275,N_718);
and U1868 (N_1868,N_562,N_899);
nor U1869 (N_1869,N_775,N_341);
nand U1870 (N_1870,N_836,N_342);
and U1871 (N_1871,N_280,N_459);
or U1872 (N_1872,N_796,N_919);
or U1873 (N_1873,N_157,N_566);
or U1874 (N_1874,N_700,N_234);
nor U1875 (N_1875,N_230,N_941);
and U1876 (N_1876,N_118,N_89);
nor U1877 (N_1877,N_501,N_638);
nand U1878 (N_1878,N_247,N_370);
nor U1879 (N_1879,N_825,N_537);
or U1880 (N_1880,N_535,N_382);
or U1881 (N_1881,N_797,N_116);
or U1882 (N_1882,N_896,N_579);
nand U1883 (N_1883,N_645,N_889);
or U1884 (N_1884,N_331,N_49);
and U1885 (N_1885,N_725,N_880);
nor U1886 (N_1886,N_438,N_557);
nand U1887 (N_1887,N_860,N_138);
nand U1888 (N_1888,N_127,N_513);
or U1889 (N_1889,N_816,N_552);
nand U1890 (N_1890,N_94,N_900);
or U1891 (N_1891,N_842,N_836);
nand U1892 (N_1892,N_38,N_570);
xnor U1893 (N_1893,N_852,N_486);
nand U1894 (N_1894,N_914,N_59);
and U1895 (N_1895,N_225,N_508);
or U1896 (N_1896,N_776,N_772);
nor U1897 (N_1897,N_311,N_201);
and U1898 (N_1898,N_335,N_494);
and U1899 (N_1899,N_90,N_174);
xnor U1900 (N_1900,N_573,N_256);
and U1901 (N_1901,N_571,N_496);
nor U1902 (N_1902,N_969,N_808);
nor U1903 (N_1903,N_521,N_492);
nor U1904 (N_1904,N_681,N_25);
or U1905 (N_1905,N_796,N_205);
or U1906 (N_1906,N_688,N_884);
nand U1907 (N_1907,N_856,N_63);
and U1908 (N_1908,N_546,N_575);
or U1909 (N_1909,N_837,N_79);
nand U1910 (N_1910,N_97,N_491);
or U1911 (N_1911,N_580,N_9);
or U1912 (N_1912,N_468,N_538);
nor U1913 (N_1913,N_198,N_689);
nor U1914 (N_1914,N_16,N_809);
and U1915 (N_1915,N_467,N_309);
and U1916 (N_1916,N_154,N_745);
and U1917 (N_1917,N_675,N_667);
and U1918 (N_1918,N_276,N_699);
nand U1919 (N_1919,N_835,N_556);
and U1920 (N_1920,N_2,N_293);
or U1921 (N_1921,N_314,N_525);
nor U1922 (N_1922,N_82,N_601);
or U1923 (N_1923,N_868,N_623);
nor U1924 (N_1924,N_492,N_183);
and U1925 (N_1925,N_600,N_540);
and U1926 (N_1926,N_600,N_625);
and U1927 (N_1927,N_117,N_559);
nand U1928 (N_1928,N_217,N_702);
or U1929 (N_1929,N_378,N_517);
and U1930 (N_1930,N_790,N_977);
nor U1931 (N_1931,N_470,N_581);
nand U1932 (N_1932,N_253,N_226);
or U1933 (N_1933,N_13,N_453);
nand U1934 (N_1934,N_283,N_22);
xnor U1935 (N_1935,N_441,N_810);
nor U1936 (N_1936,N_171,N_73);
and U1937 (N_1937,N_31,N_43);
and U1938 (N_1938,N_792,N_171);
and U1939 (N_1939,N_777,N_669);
or U1940 (N_1940,N_566,N_80);
nand U1941 (N_1941,N_309,N_820);
nor U1942 (N_1942,N_391,N_903);
xor U1943 (N_1943,N_929,N_215);
and U1944 (N_1944,N_252,N_242);
or U1945 (N_1945,N_781,N_278);
nand U1946 (N_1946,N_243,N_319);
nand U1947 (N_1947,N_23,N_443);
nor U1948 (N_1948,N_901,N_697);
nor U1949 (N_1949,N_46,N_845);
nor U1950 (N_1950,N_778,N_484);
xnor U1951 (N_1951,N_728,N_738);
and U1952 (N_1952,N_385,N_830);
xnor U1953 (N_1953,N_407,N_297);
xor U1954 (N_1954,N_539,N_603);
or U1955 (N_1955,N_987,N_151);
and U1956 (N_1956,N_271,N_332);
or U1957 (N_1957,N_782,N_176);
nor U1958 (N_1958,N_604,N_901);
nand U1959 (N_1959,N_578,N_957);
nor U1960 (N_1960,N_601,N_414);
nand U1961 (N_1961,N_769,N_758);
nand U1962 (N_1962,N_813,N_999);
and U1963 (N_1963,N_86,N_863);
nor U1964 (N_1964,N_106,N_235);
nand U1965 (N_1965,N_725,N_647);
and U1966 (N_1966,N_272,N_365);
nor U1967 (N_1967,N_679,N_223);
nor U1968 (N_1968,N_691,N_736);
and U1969 (N_1969,N_938,N_210);
nor U1970 (N_1970,N_361,N_909);
nor U1971 (N_1971,N_952,N_960);
and U1972 (N_1972,N_224,N_805);
nand U1973 (N_1973,N_953,N_662);
or U1974 (N_1974,N_343,N_780);
nand U1975 (N_1975,N_721,N_593);
or U1976 (N_1976,N_963,N_47);
nand U1977 (N_1977,N_632,N_673);
nand U1978 (N_1978,N_555,N_199);
and U1979 (N_1979,N_666,N_4);
nor U1980 (N_1980,N_812,N_394);
or U1981 (N_1981,N_402,N_32);
nand U1982 (N_1982,N_746,N_132);
and U1983 (N_1983,N_684,N_29);
nor U1984 (N_1984,N_58,N_257);
or U1985 (N_1985,N_465,N_52);
and U1986 (N_1986,N_579,N_605);
or U1987 (N_1987,N_189,N_126);
or U1988 (N_1988,N_125,N_601);
xor U1989 (N_1989,N_732,N_555);
and U1990 (N_1990,N_207,N_526);
and U1991 (N_1991,N_580,N_581);
nand U1992 (N_1992,N_670,N_168);
or U1993 (N_1993,N_89,N_242);
xnor U1994 (N_1994,N_466,N_630);
or U1995 (N_1995,N_253,N_477);
nand U1996 (N_1996,N_715,N_811);
nand U1997 (N_1997,N_229,N_851);
or U1998 (N_1998,N_265,N_144);
nand U1999 (N_1999,N_814,N_192);
nor U2000 (N_2000,N_1815,N_1404);
or U2001 (N_2001,N_1242,N_1349);
nand U2002 (N_2002,N_1270,N_1072);
xor U2003 (N_2003,N_1983,N_1034);
and U2004 (N_2004,N_1579,N_1736);
nor U2005 (N_2005,N_1458,N_1259);
nand U2006 (N_2006,N_1354,N_1485);
or U2007 (N_2007,N_1699,N_1432);
nand U2008 (N_2008,N_1967,N_1070);
or U2009 (N_2009,N_1116,N_1313);
nor U2010 (N_2010,N_1080,N_1940);
nand U2011 (N_2011,N_1988,N_1127);
nand U2012 (N_2012,N_1322,N_1756);
xnor U2013 (N_2013,N_1799,N_1695);
nand U2014 (N_2014,N_1055,N_1180);
nor U2015 (N_2015,N_1450,N_1566);
and U2016 (N_2016,N_1532,N_1851);
and U2017 (N_2017,N_1543,N_1493);
nand U2018 (N_2018,N_1057,N_1375);
nand U2019 (N_2019,N_1514,N_1042);
nand U2020 (N_2020,N_1901,N_1386);
and U2021 (N_2021,N_1771,N_1569);
and U2022 (N_2022,N_1408,N_1460);
or U2023 (N_2023,N_1757,N_1991);
and U2024 (N_2024,N_1064,N_1775);
nor U2025 (N_2025,N_1682,N_1407);
nor U2026 (N_2026,N_1183,N_1416);
nand U2027 (N_2027,N_1018,N_1453);
or U2028 (N_2028,N_1081,N_1937);
nor U2029 (N_2029,N_1392,N_1681);
nor U2030 (N_2030,N_1791,N_1040);
nand U2031 (N_2031,N_1678,N_1638);
nand U2032 (N_2032,N_1722,N_1728);
nor U2033 (N_2033,N_1248,N_1021);
nor U2034 (N_2034,N_1043,N_1198);
and U2035 (N_2035,N_1337,N_1475);
and U2036 (N_2036,N_1447,N_1743);
or U2037 (N_2037,N_1918,N_1136);
and U2038 (N_2038,N_1727,N_1117);
or U2039 (N_2039,N_1491,N_1044);
or U2040 (N_2040,N_1606,N_1660);
nor U2041 (N_2041,N_1559,N_1168);
nor U2042 (N_2042,N_1865,N_1083);
and U2043 (N_2043,N_1219,N_1990);
and U2044 (N_2044,N_1500,N_1708);
nand U2045 (N_2045,N_1106,N_1241);
nand U2046 (N_2046,N_1669,N_1221);
nand U2047 (N_2047,N_1326,N_1469);
nor U2048 (N_2048,N_1870,N_1925);
nand U2049 (N_2049,N_1105,N_1496);
nand U2050 (N_2050,N_1670,N_1656);
or U2051 (N_2051,N_1169,N_1288);
or U2052 (N_2052,N_1094,N_1048);
nor U2053 (N_2053,N_1082,N_1527);
nor U2054 (N_2054,N_1079,N_1867);
nand U2055 (N_2055,N_1425,N_1192);
or U2056 (N_2056,N_1145,N_1140);
or U2057 (N_2057,N_1060,N_1895);
and U2058 (N_2058,N_1672,N_1351);
or U2059 (N_2059,N_1151,N_1748);
and U2060 (N_2060,N_1481,N_1550);
nor U2061 (N_2061,N_1857,N_1764);
and U2062 (N_2062,N_1395,N_1464);
nor U2063 (N_2063,N_1181,N_1714);
and U2064 (N_2064,N_1926,N_1161);
nor U2065 (N_2065,N_1903,N_1947);
nor U2066 (N_2066,N_1341,N_1463);
nand U2067 (N_2067,N_1433,N_1636);
and U2068 (N_2068,N_1750,N_1632);
or U2069 (N_2069,N_1664,N_1759);
nand U2070 (N_2070,N_1935,N_1648);
or U2071 (N_2071,N_1760,N_1697);
and U2072 (N_2072,N_1418,N_1202);
nand U2073 (N_2073,N_1560,N_1942);
xnor U2074 (N_2074,N_1770,N_1769);
xor U2075 (N_2075,N_1223,N_1900);
nor U2076 (N_2076,N_1362,N_1572);
or U2077 (N_2077,N_1196,N_1065);
nand U2078 (N_2078,N_1657,N_1627);
or U2079 (N_2079,N_1225,N_1616);
and U2080 (N_2080,N_1840,N_1817);
or U2081 (N_2081,N_1347,N_1758);
or U2082 (N_2082,N_1258,N_1741);
nor U2083 (N_2083,N_1601,N_1363);
nand U2084 (N_2084,N_1443,N_1873);
and U2085 (N_2085,N_1230,N_1488);
nor U2086 (N_2086,N_1554,N_1971);
nand U2087 (N_2087,N_1327,N_1329);
nand U2088 (N_2088,N_1402,N_1710);
nand U2089 (N_2089,N_1558,N_1565);
nor U2090 (N_2090,N_1644,N_1535);
nor U2091 (N_2091,N_1422,N_1251);
and U2092 (N_2092,N_1751,N_1603);
nand U2093 (N_2093,N_1095,N_1665);
or U2094 (N_2094,N_1077,N_1119);
or U2095 (N_2095,N_1104,N_1725);
nor U2096 (N_2096,N_1253,N_1275);
or U2097 (N_2097,N_1252,N_1629);
and U2098 (N_2098,N_1372,N_1790);
or U2099 (N_2099,N_1035,N_1483);
nor U2100 (N_2100,N_1308,N_1272);
or U2101 (N_2101,N_1692,N_1777);
nor U2102 (N_2102,N_1555,N_1100);
and U2103 (N_2103,N_1928,N_1446);
or U2104 (N_2104,N_1097,N_1772);
xnor U2105 (N_2105,N_1224,N_1019);
and U2106 (N_2106,N_1796,N_1803);
nand U2107 (N_2107,N_1165,N_1607);
nor U2108 (N_2108,N_1970,N_1583);
and U2109 (N_2109,N_1254,N_1498);
nor U2110 (N_2110,N_1376,N_1442);
nand U2111 (N_2111,N_1980,N_1784);
or U2112 (N_2112,N_1370,N_1150);
nand U2113 (N_2113,N_1344,N_1069);
and U2114 (N_2114,N_1473,N_1147);
nor U2115 (N_2115,N_1597,N_1625);
nand U2116 (N_2116,N_1552,N_1182);
nand U2117 (N_2117,N_1076,N_1438);
or U2118 (N_2118,N_1912,N_1222);
and U2119 (N_2119,N_1087,N_1662);
nor U2120 (N_2120,N_1012,N_1209);
and U2121 (N_2121,N_1833,N_1573);
and U2122 (N_2122,N_1515,N_1371);
and U2123 (N_2123,N_1067,N_1071);
nor U2124 (N_2124,N_1938,N_1963);
and U2125 (N_2125,N_1679,N_1123);
nor U2126 (N_2126,N_1776,N_1789);
or U2127 (N_2127,N_1073,N_1093);
and U2128 (N_2128,N_1620,N_1276);
nor U2129 (N_2129,N_1782,N_1244);
nor U2130 (N_2130,N_1321,N_1250);
or U2131 (N_2131,N_1440,N_1186);
or U2132 (N_2132,N_1765,N_1278);
nand U2133 (N_2133,N_1280,N_1673);
nand U2134 (N_2134,N_1838,N_1295);
or U2135 (N_2135,N_1617,N_1089);
nand U2136 (N_2136,N_1046,N_1539);
and U2137 (N_2137,N_1146,N_1477);
or U2138 (N_2138,N_1936,N_1397);
nor U2139 (N_2139,N_1226,N_1525);
nand U2140 (N_2140,N_1512,N_1216);
nor U2141 (N_2141,N_1968,N_1902);
nor U2142 (N_2142,N_1431,N_1588);
and U2143 (N_2143,N_1001,N_1962);
and U2144 (N_2144,N_1489,N_1516);
and U2145 (N_2145,N_1702,N_1479);
or U2146 (N_2146,N_1016,N_1238);
nand U2147 (N_2147,N_1004,N_1228);
nand U2148 (N_2148,N_1298,N_1646);
nor U2149 (N_2149,N_1747,N_1779);
and U2150 (N_2150,N_1694,N_1314);
nor U2151 (N_2151,N_1804,N_1036);
nor U2152 (N_2152,N_1187,N_1302);
nand U2153 (N_2153,N_1826,N_1883);
nand U2154 (N_2154,N_1951,N_1810);
and U2155 (N_2155,N_1227,N_1593);
nand U2156 (N_2156,N_1706,N_1486);
or U2157 (N_2157,N_1941,N_1164);
nand U2158 (N_2158,N_1499,N_1086);
and U2159 (N_2159,N_1484,N_1246);
or U2160 (N_2160,N_1148,N_1029);
or U2161 (N_2161,N_1996,N_1507);
and U2162 (N_2162,N_1245,N_1703);
or U2163 (N_2163,N_1577,N_1600);
nor U2164 (N_2164,N_1045,N_1053);
or U2165 (N_2165,N_1237,N_1017);
nor U2166 (N_2166,N_1973,N_1156);
and U2167 (N_2167,N_1032,N_1113);
nor U2168 (N_2168,N_1688,N_1821);
nand U2169 (N_2169,N_1260,N_1075);
or U2170 (N_2170,N_1255,N_1266);
nor U2171 (N_2171,N_1568,N_1661);
or U2172 (N_2172,N_1426,N_1590);
or U2173 (N_2173,N_1909,N_1822);
or U2174 (N_2174,N_1742,N_1309);
nand U2175 (N_2175,N_1159,N_1257);
nor U2176 (N_2176,N_1866,N_1786);
nand U2177 (N_2177,N_1318,N_1846);
nor U2178 (N_2178,N_1291,N_1508);
nor U2179 (N_2179,N_1652,N_1718);
or U2180 (N_2180,N_1820,N_1343);
and U2181 (N_2181,N_1998,N_1289);
and U2182 (N_2182,N_1965,N_1542);
and U2183 (N_2183,N_1808,N_1614);
and U2184 (N_2184,N_1667,N_1716);
and U2185 (N_2185,N_1858,N_1476);
and U2186 (N_2186,N_1304,N_1534);
or U2187 (N_2187,N_1474,N_1730);
nand U2188 (N_2188,N_1802,N_1611);
and U2189 (N_2189,N_1247,N_1160);
nor U2190 (N_2190,N_1598,N_1465);
or U2191 (N_2191,N_1051,N_1078);
nand U2192 (N_2192,N_1393,N_1390);
or U2193 (N_2193,N_1825,N_1969);
or U2194 (N_2194,N_1005,N_1541);
nor U2195 (N_2195,N_1624,N_1120);
xor U2196 (N_2196,N_1357,N_1828);
xor U2197 (N_2197,N_1406,N_1437);
or U2198 (N_2198,N_1952,N_1428);
and U2199 (N_2199,N_1847,N_1179);
nor U2200 (N_2200,N_1285,N_1423);
or U2201 (N_2201,N_1618,N_1800);
and U2202 (N_2202,N_1932,N_1850);
nor U2203 (N_2203,N_1213,N_1502);
nand U2204 (N_2204,N_1099,N_1880);
nor U2205 (N_2205,N_1794,N_1689);
and U2206 (N_2206,N_1894,N_1712);
and U2207 (N_2207,N_1511,N_1856);
nor U2208 (N_2208,N_1687,N_1835);
nor U2209 (N_2209,N_1934,N_1480);
nand U2210 (N_2210,N_1365,N_1206);
and U2211 (N_2211,N_1668,N_1158);
and U2212 (N_2212,N_1766,N_1739);
or U2213 (N_2213,N_1331,N_1448);
nor U2214 (N_2214,N_1421,N_1726);
and U2215 (N_2215,N_1905,N_1605);
and U2216 (N_2216,N_1842,N_1457);
nand U2217 (N_2217,N_1696,N_1584);
nor U2218 (N_2218,N_1761,N_1504);
or U2219 (N_2219,N_1024,N_1879);
nor U2220 (N_2220,N_1052,N_1384);
nor U2221 (N_2221,N_1130,N_1832);
nand U2222 (N_2222,N_1424,N_1063);
or U2223 (N_2223,N_1993,N_1110);
nand U2224 (N_2224,N_1650,N_1651);
nor U2225 (N_2225,N_1509,N_1353);
nand U2226 (N_2226,N_1881,N_1307);
nor U2227 (N_2227,N_1721,N_1961);
or U2228 (N_2228,N_1346,N_1643);
or U2229 (N_2229,N_1613,N_1586);
or U2230 (N_2230,N_1429,N_1358);
nand U2231 (N_2231,N_1068,N_1557);
nand U2232 (N_2232,N_1330,N_1615);
nor U2233 (N_2233,N_1666,N_1830);
nor U2234 (N_2234,N_1704,N_1995);
or U2235 (N_2235,N_1378,N_1478);
nor U2236 (N_2236,N_1400,N_1176);
nand U2237 (N_2237,N_1671,N_1449);
or U2238 (N_2238,N_1293,N_1412);
and U2239 (N_2239,N_1373,N_1752);
and U2240 (N_2240,N_1896,N_1294);
and U2241 (N_2241,N_1296,N_1154);
nor U2242 (N_2242,N_1103,N_1133);
nor U2243 (N_2243,N_1454,N_1379);
nor U2244 (N_2244,N_1312,N_1023);
and U2245 (N_2245,N_1342,N_1128);
nor U2246 (N_2246,N_1190,N_1435);
nor U2247 (N_2247,N_1173,N_1753);
nand U2248 (N_2248,N_1286,N_1112);
or U2249 (N_2249,N_1829,N_1874);
or U2250 (N_2250,N_1439,N_1050);
and U2251 (N_2251,N_1746,N_1914);
or U2252 (N_2252,N_1468,N_1578);
xnor U2253 (N_2253,N_1350,N_1265);
or U2254 (N_2254,N_1979,N_1062);
or U2255 (N_2255,N_1367,N_1831);
nor U2256 (N_2256,N_1452,N_1391);
and U2257 (N_2257,N_1986,N_1191);
or U2258 (N_2258,N_1490,N_1006);
nor U2259 (N_2259,N_1920,N_1540);
nor U2260 (N_2260,N_1398,N_1088);
or U2261 (N_2261,N_1340,N_1129);
xor U2262 (N_2262,N_1459,N_1609);
nand U2263 (N_2263,N_1749,N_1240);
and U2264 (N_2264,N_1564,N_1334);
nand U2265 (N_2265,N_1861,N_1229);
nand U2266 (N_2266,N_1256,N_1441);
or U2267 (N_2267,N_1547,N_1455);
nor U2268 (N_2268,N_1994,N_1982);
nor U2269 (N_2269,N_1913,N_1084);
or U2270 (N_2270,N_1430,N_1788);
or U2271 (N_2271,N_1526,N_1143);
nor U2272 (N_2272,N_1953,N_1645);
nand U2273 (N_2273,N_1599,N_1649);
nor U2274 (N_2274,N_1167,N_1619);
and U2275 (N_2275,N_1249,N_1269);
xnor U2276 (N_2276,N_1456,N_1303);
nor U2277 (N_2277,N_1470,N_1818);
nand U2278 (N_2278,N_1283,N_1015);
and U2279 (N_2279,N_1118,N_1674);
or U2280 (N_2280,N_1152,N_1215);
nor U2281 (N_2281,N_1956,N_1157);
nor U2282 (N_2282,N_1310,N_1211);
nand U2283 (N_2283,N_1243,N_1630);
and U2284 (N_2284,N_1263,N_1819);
nor U2285 (N_2285,N_1634,N_1904);
and U2286 (N_2286,N_1008,N_1419);
nand U2287 (N_2287,N_1868,N_1273);
and U2288 (N_2288,N_1561,N_1427);
nor U2289 (N_2289,N_1039,N_1131);
nand U2290 (N_2290,N_1188,N_1882);
nand U2291 (N_2291,N_1544,N_1734);
or U2292 (N_2292,N_1403,N_1778);
and U2293 (N_2293,N_1691,N_1889);
or U2294 (N_2294,N_1524,N_1212);
nand U2295 (N_2295,N_1729,N_1002);
and U2296 (N_2296,N_1907,N_1501);
nor U2297 (N_2297,N_1812,N_1494);
or U2298 (N_2298,N_1345,N_1898);
or U2299 (N_2299,N_1359,N_1262);
nor U2300 (N_2300,N_1843,N_1031);
nor U2301 (N_2301,N_1284,N_1852);
or U2302 (N_2302,N_1409,N_1415);
nand U2303 (N_2303,N_1834,N_1676);
and U2304 (N_2304,N_1194,N_1102);
or U2305 (N_2305,N_1809,N_1793);
or U2306 (N_2306,N_1451,N_1399);
nand U2307 (N_2307,N_1038,N_1774);
and U2308 (N_2308,N_1381,N_1010);
and U2309 (N_2309,N_1859,N_1585);
or U2310 (N_2310,N_1964,N_1801);
nor U2311 (N_2311,N_1126,N_1977);
nand U2312 (N_2312,N_1581,N_1471);
nand U2313 (N_2313,N_1189,N_1096);
or U2314 (N_2314,N_1413,N_1872);
and U2315 (N_2315,N_1806,N_1707);
or U2316 (N_2316,N_1153,N_1686);
nor U2317 (N_2317,N_1855,N_1949);
and U2318 (N_2318,N_1738,N_1693);
or U2319 (N_2319,N_1921,N_1591);
and U2320 (N_2320,N_1014,N_1166);
nand U2321 (N_2321,N_1355,N_1939);
nor U2322 (N_2322,N_1217,N_1420);
and U2323 (N_2323,N_1642,N_1595);
xnor U2324 (N_2324,N_1141,N_1510);
nor U2325 (N_2325,N_1785,N_1612);
nor U2326 (N_2326,N_1301,N_1271);
nor U2327 (N_2327,N_1853,N_1827);
nor U2328 (N_2328,N_1142,N_1592);
nor U2329 (N_2329,N_1529,N_1315);
nor U2330 (N_2330,N_1628,N_1085);
nor U2331 (N_2331,N_1139,N_1200);
or U2332 (N_2332,N_1109,N_1700);
nor U2333 (N_2333,N_1305,N_1717);
and U2334 (N_2334,N_1975,N_1677);
nand U2335 (N_2335,N_1162,N_1763);
and U2336 (N_2336,N_1892,N_1546);
and U2337 (N_2337,N_1528,N_1382);
and U2338 (N_2338,N_1466,N_1279);
and U2339 (N_2339,N_1348,N_1517);
or U2340 (N_2340,N_1675,N_1361);
nor U2341 (N_2341,N_1405,N_1610);
and U2342 (N_2342,N_1582,N_1893);
nand U2343 (N_2343,N_1860,N_1335);
nand U2344 (N_2344,N_1556,N_1633);
and U2345 (N_2345,N_1945,N_1981);
and U2346 (N_2346,N_1875,N_1122);
nor U2347 (N_2347,N_1944,N_1623);
nor U2348 (N_2348,N_1115,N_1955);
nor U2349 (N_2349,N_1175,N_1414);
nor U2350 (N_2350,N_1884,N_1047);
or U2351 (N_2351,N_1049,N_1236);
and U2352 (N_2352,N_1383,N_1571);
and U2353 (N_2353,N_1795,N_1797);
or U2354 (N_2354,N_1411,N_1886);
and U2355 (N_2355,N_1723,N_1631);
or U2356 (N_2356,N_1744,N_1011);
nor U2357 (N_2357,N_1715,N_1916);
nand U2358 (N_2358,N_1647,N_1138);
and U2359 (N_2359,N_1267,N_1997);
and U2360 (N_2360,N_1877,N_1261);
nor U2361 (N_2361,N_1923,N_1890);
nor U2362 (N_2362,N_1058,N_1594);
nand U2363 (N_2363,N_1596,N_1003);
nor U2364 (N_2364,N_1897,N_1316);
nor U2365 (N_2365,N_1984,N_1092);
and U2366 (N_2366,N_1957,N_1663);
and U2367 (N_2367,N_1943,N_1320);
and U2368 (N_2368,N_1518,N_1028);
or U2369 (N_2369,N_1570,N_1108);
nand U2370 (N_2370,N_1987,N_1864);
nor U2371 (N_2371,N_1985,N_1899);
or U2372 (N_2372,N_1090,N_1608);
or U2373 (N_2373,N_1948,N_1910);
and U2374 (N_2374,N_1174,N_1640);
nand U2375 (N_2375,N_1134,N_1467);
and U2376 (N_2376,N_1107,N_1966);
or U2377 (N_2377,N_1767,N_1807);
and U2378 (N_2378,N_1364,N_1144);
and U2379 (N_2379,N_1233,N_1436);
nor U2380 (N_2380,N_1172,N_1538);
nor U2381 (N_2381,N_1377,N_1733);
or U2382 (N_2382,N_1155,N_1837);
or U2383 (N_2383,N_1124,N_1622);
nand U2384 (N_2384,N_1022,N_1924);
and U2385 (N_2385,N_1000,N_1562);
nand U2386 (N_2386,N_1589,N_1724);
nor U2387 (N_2387,N_1805,N_1519);
or U2388 (N_2388,N_1732,N_1149);
nor U2389 (N_2389,N_1992,N_1933);
and U2390 (N_2390,N_1989,N_1537);
nand U2391 (N_2391,N_1396,N_1709);
or U2392 (N_2392,N_1290,N_1635);
nand U2393 (N_2393,N_1328,N_1324);
or U2394 (N_2394,N_1931,N_1737);
nor U2395 (N_2395,N_1311,N_1927);
nor U2396 (N_2396,N_1978,N_1773);
nand U2397 (N_2397,N_1231,N_1185);
nand U2398 (N_2398,N_1735,N_1444);
nand U2399 (N_2399,N_1745,N_1930);
nor U2400 (N_2400,N_1711,N_1274);
and U2401 (N_2401,N_1520,N_1587);
and U2402 (N_2402,N_1959,N_1417);
nand U2403 (N_2403,N_1685,N_1027);
and U2404 (N_2404,N_1871,N_1848);
and U2405 (N_2405,N_1319,N_1958);
nor U2406 (N_2406,N_1658,N_1210);
nand U2407 (N_2407,N_1911,N_1091);
nor U2408 (N_2408,N_1954,N_1203);
nor U2409 (N_2409,N_1976,N_1235);
xnor U2410 (N_2410,N_1234,N_1025);
nor U2411 (N_2411,N_1713,N_1531);
nor U2412 (N_2412,N_1292,N_1654);
and U2413 (N_2413,N_1639,N_1218);
and U2414 (N_2414,N_1823,N_1061);
and U2415 (N_2415,N_1891,N_1621);
nor U2416 (N_2416,N_1171,N_1059);
and U2417 (N_2417,N_1548,N_1387);
nor U2418 (N_2418,N_1841,N_1680);
nor U2419 (N_2419,N_1195,N_1264);
nor U2420 (N_2420,N_1193,N_1282);
or U2421 (N_2421,N_1869,N_1323);
or U2422 (N_2422,N_1740,N_1530);
nand U2423 (N_2423,N_1523,N_1915);
or U2424 (N_2424,N_1836,N_1434);
and U2425 (N_2425,N_1705,N_1545);
nor U2426 (N_2426,N_1919,N_1205);
nand U2427 (N_2427,N_1197,N_1299);
and U2428 (N_2428,N_1813,N_1268);
and U2429 (N_2429,N_1352,N_1220);
nor U2430 (N_2430,N_1178,N_1731);
and U2431 (N_2431,N_1170,N_1659);
nor U2432 (N_2432,N_1297,N_1683);
nor U2433 (N_2433,N_1946,N_1492);
and U2434 (N_2434,N_1495,N_1385);
or U2435 (N_2435,N_1204,N_1325);
nor U2436 (N_2436,N_1533,N_1787);
and U2437 (N_2437,N_1780,N_1401);
nor U2438 (N_2438,N_1762,N_1798);
nand U2439 (N_2439,N_1887,N_1505);
or U2440 (N_2440,N_1655,N_1098);
or U2441 (N_2441,N_1626,N_1356);
or U2442 (N_2442,N_1030,N_1101);
and U2443 (N_2443,N_1184,N_1513);
nand U2444 (N_2444,N_1369,N_1849);
nand U2445 (N_2445,N_1332,N_1974);
nand U2446 (N_2446,N_1792,N_1999);
nor U2447 (N_2447,N_1287,N_1336);
nand U2448 (N_2448,N_1641,N_1461);
or U2449 (N_2449,N_1698,N_1125);
or U2450 (N_2450,N_1960,N_1037);
nor U2451 (N_2451,N_1306,N_1239);
or U2452 (N_2452,N_1487,N_1111);
or U2453 (N_2453,N_1575,N_1521);
and U2454 (N_2454,N_1033,N_1754);
and U2455 (N_2455,N_1917,N_1056);
nand U2456 (N_2456,N_1576,N_1074);
nand U2457 (N_2457,N_1388,N_1013);
and U2458 (N_2458,N_1637,N_1522);
nand U2459 (N_2459,N_1844,N_1604);
or U2460 (N_2460,N_1135,N_1878);
or U2461 (N_2461,N_1720,N_1338);
nor U2462 (N_2462,N_1816,N_1009);
nand U2463 (N_2463,N_1339,N_1580);
nand U2464 (N_2464,N_1020,N_1137);
nor U2465 (N_2465,N_1380,N_1854);
and U2466 (N_2466,N_1366,N_1317);
nor U2467 (N_2467,N_1360,N_1026);
and U2468 (N_2468,N_1277,N_1300);
and U2469 (N_2469,N_1368,N_1783);
nand U2470 (N_2470,N_1472,N_1684);
nand U2471 (N_2471,N_1950,N_1811);
xnor U2472 (N_2472,N_1482,N_1281);
and U2473 (N_2473,N_1054,N_1814);
or U2474 (N_2474,N_1410,N_1755);
and U2475 (N_2475,N_1781,N_1007);
nor U2476 (N_2476,N_1132,N_1462);
xnor U2477 (N_2477,N_1701,N_1497);
nor U2478 (N_2478,N_1862,N_1232);
nand U2479 (N_2479,N_1201,N_1199);
and U2480 (N_2480,N_1876,N_1207);
nor U2481 (N_2481,N_1394,N_1536);
or U2482 (N_2482,N_1602,N_1908);
nor U2483 (N_2483,N_1922,N_1066);
and U2484 (N_2484,N_1768,N_1574);
or U2485 (N_2485,N_1567,N_1824);
or U2486 (N_2486,N_1208,N_1553);
xnor U2487 (N_2487,N_1177,N_1863);
nor U2488 (N_2488,N_1551,N_1929);
xnor U2489 (N_2489,N_1374,N_1389);
and U2490 (N_2490,N_1114,N_1121);
nor U2491 (N_2491,N_1163,N_1214);
nand U2492 (N_2492,N_1041,N_1885);
nand U2493 (N_2493,N_1506,N_1906);
or U2494 (N_2494,N_1445,N_1845);
nand U2495 (N_2495,N_1719,N_1333);
and U2496 (N_2496,N_1549,N_1563);
nand U2497 (N_2497,N_1503,N_1888);
nor U2498 (N_2498,N_1690,N_1653);
and U2499 (N_2499,N_1972,N_1839);
and U2500 (N_2500,N_1666,N_1533);
nand U2501 (N_2501,N_1740,N_1697);
or U2502 (N_2502,N_1508,N_1144);
nor U2503 (N_2503,N_1002,N_1215);
nand U2504 (N_2504,N_1189,N_1013);
or U2505 (N_2505,N_1303,N_1497);
nand U2506 (N_2506,N_1630,N_1611);
nand U2507 (N_2507,N_1327,N_1025);
nor U2508 (N_2508,N_1680,N_1804);
nor U2509 (N_2509,N_1426,N_1232);
nand U2510 (N_2510,N_1355,N_1401);
or U2511 (N_2511,N_1525,N_1323);
or U2512 (N_2512,N_1384,N_1042);
nand U2513 (N_2513,N_1657,N_1341);
nor U2514 (N_2514,N_1781,N_1691);
nand U2515 (N_2515,N_1491,N_1386);
nand U2516 (N_2516,N_1194,N_1107);
nand U2517 (N_2517,N_1616,N_1602);
nand U2518 (N_2518,N_1256,N_1531);
nand U2519 (N_2519,N_1674,N_1874);
nor U2520 (N_2520,N_1164,N_1831);
nor U2521 (N_2521,N_1874,N_1697);
and U2522 (N_2522,N_1894,N_1984);
or U2523 (N_2523,N_1665,N_1711);
or U2524 (N_2524,N_1740,N_1382);
nor U2525 (N_2525,N_1353,N_1618);
and U2526 (N_2526,N_1772,N_1176);
and U2527 (N_2527,N_1112,N_1481);
nand U2528 (N_2528,N_1059,N_1081);
nor U2529 (N_2529,N_1589,N_1159);
or U2530 (N_2530,N_1849,N_1426);
nand U2531 (N_2531,N_1648,N_1399);
nor U2532 (N_2532,N_1190,N_1682);
or U2533 (N_2533,N_1584,N_1827);
nand U2534 (N_2534,N_1577,N_1733);
and U2535 (N_2535,N_1267,N_1118);
or U2536 (N_2536,N_1792,N_1572);
nor U2537 (N_2537,N_1794,N_1680);
nor U2538 (N_2538,N_1963,N_1142);
and U2539 (N_2539,N_1451,N_1180);
or U2540 (N_2540,N_1387,N_1732);
and U2541 (N_2541,N_1824,N_1788);
and U2542 (N_2542,N_1542,N_1920);
nor U2543 (N_2543,N_1999,N_1222);
nor U2544 (N_2544,N_1454,N_1027);
nand U2545 (N_2545,N_1344,N_1305);
and U2546 (N_2546,N_1123,N_1645);
or U2547 (N_2547,N_1407,N_1620);
nand U2548 (N_2548,N_1423,N_1562);
or U2549 (N_2549,N_1763,N_1087);
or U2550 (N_2550,N_1365,N_1817);
nand U2551 (N_2551,N_1929,N_1052);
or U2552 (N_2552,N_1506,N_1363);
and U2553 (N_2553,N_1498,N_1784);
nor U2554 (N_2554,N_1868,N_1690);
nor U2555 (N_2555,N_1862,N_1479);
and U2556 (N_2556,N_1536,N_1380);
and U2557 (N_2557,N_1534,N_1002);
and U2558 (N_2558,N_1048,N_1765);
or U2559 (N_2559,N_1911,N_1850);
nand U2560 (N_2560,N_1062,N_1090);
and U2561 (N_2561,N_1885,N_1137);
nand U2562 (N_2562,N_1125,N_1617);
nand U2563 (N_2563,N_1592,N_1015);
nand U2564 (N_2564,N_1345,N_1132);
nor U2565 (N_2565,N_1547,N_1725);
nor U2566 (N_2566,N_1731,N_1417);
or U2567 (N_2567,N_1731,N_1126);
and U2568 (N_2568,N_1066,N_1771);
nor U2569 (N_2569,N_1475,N_1754);
or U2570 (N_2570,N_1247,N_1752);
nor U2571 (N_2571,N_1490,N_1414);
nor U2572 (N_2572,N_1094,N_1949);
and U2573 (N_2573,N_1829,N_1934);
nor U2574 (N_2574,N_1842,N_1805);
and U2575 (N_2575,N_1394,N_1083);
nor U2576 (N_2576,N_1603,N_1717);
or U2577 (N_2577,N_1268,N_1072);
nand U2578 (N_2578,N_1893,N_1931);
and U2579 (N_2579,N_1720,N_1188);
nor U2580 (N_2580,N_1384,N_1682);
or U2581 (N_2581,N_1138,N_1460);
nor U2582 (N_2582,N_1445,N_1198);
nand U2583 (N_2583,N_1899,N_1515);
nor U2584 (N_2584,N_1026,N_1346);
nand U2585 (N_2585,N_1312,N_1050);
and U2586 (N_2586,N_1374,N_1940);
or U2587 (N_2587,N_1472,N_1634);
and U2588 (N_2588,N_1488,N_1090);
nor U2589 (N_2589,N_1803,N_1571);
nand U2590 (N_2590,N_1953,N_1882);
nand U2591 (N_2591,N_1669,N_1076);
or U2592 (N_2592,N_1974,N_1464);
or U2593 (N_2593,N_1546,N_1765);
and U2594 (N_2594,N_1978,N_1022);
and U2595 (N_2595,N_1329,N_1456);
or U2596 (N_2596,N_1933,N_1859);
or U2597 (N_2597,N_1579,N_1260);
nor U2598 (N_2598,N_1128,N_1578);
nor U2599 (N_2599,N_1407,N_1859);
or U2600 (N_2600,N_1477,N_1212);
or U2601 (N_2601,N_1408,N_1237);
nand U2602 (N_2602,N_1115,N_1541);
nand U2603 (N_2603,N_1205,N_1991);
nand U2604 (N_2604,N_1349,N_1030);
and U2605 (N_2605,N_1488,N_1409);
or U2606 (N_2606,N_1548,N_1261);
nand U2607 (N_2607,N_1502,N_1430);
nor U2608 (N_2608,N_1006,N_1494);
nand U2609 (N_2609,N_1422,N_1318);
and U2610 (N_2610,N_1515,N_1431);
nor U2611 (N_2611,N_1573,N_1347);
and U2612 (N_2612,N_1616,N_1548);
or U2613 (N_2613,N_1802,N_1354);
nand U2614 (N_2614,N_1864,N_1265);
or U2615 (N_2615,N_1376,N_1199);
or U2616 (N_2616,N_1630,N_1915);
xnor U2617 (N_2617,N_1382,N_1968);
nor U2618 (N_2618,N_1926,N_1405);
nor U2619 (N_2619,N_1015,N_1286);
and U2620 (N_2620,N_1551,N_1823);
nor U2621 (N_2621,N_1721,N_1166);
nor U2622 (N_2622,N_1185,N_1501);
nor U2623 (N_2623,N_1938,N_1263);
and U2624 (N_2624,N_1396,N_1357);
and U2625 (N_2625,N_1441,N_1712);
nor U2626 (N_2626,N_1701,N_1418);
nand U2627 (N_2627,N_1720,N_1405);
and U2628 (N_2628,N_1709,N_1024);
nand U2629 (N_2629,N_1163,N_1046);
nand U2630 (N_2630,N_1953,N_1489);
or U2631 (N_2631,N_1956,N_1486);
and U2632 (N_2632,N_1576,N_1377);
xnor U2633 (N_2633,N_1289,N_1396);
or U2634 (N_2634,N_1032,N_1267);
or U2635 (N_2635,N_1561,N_1867);
and U2636 (N_2636,N_1866,N_1445);
or U2637 (N_2637,N_1297,N_1408);
nand U2638 (N_2638,N_1993,N_1475);
or U2639 (N_2639,N_1129,N_1245);
and U2640 (N_2640,N_1939,N_1972);
nand U2641 (N_2641,N_1534,N_1457);
nand U2642 (N_2642,N_1750,N_1673);
or U2643 (N_2643,N_1533,N_1849);
nor U2644 (N_2644,N_1006,N_1382);
xnor U2645 (N_2645,N_1832,N_1753);
nand U2646 (N_2646,N_1168,N_1369);
and U2647 (N_2647,N_1375,N_1261);
nor U2648 (N_2648,N_1738,N_1961);
nand U2649 (N_2649,N_1454,N_1488);
and U2650 (N_2650,N_1168,N_1333);
and U2651 (N_2651,N_1281,N_1456);
or U2652 (N_2652,N_1754,N_1432);
or U2653 (N_2653,N_1135,N_1779);
nand U2654 (N_2654,N_1580,N_1988);
or U2655 (N_2655,N_1615,N_1623);
nand U2656 (N_2656,N_1563,N_1198);
nand U2657 (N_2657,N_1341,N_1253);
or U2658 (N_2658,N_1040,N_1252);
and U2659 (N_2659,N_1473,N_1837);
or U2660 (N_2660,N_1580,N_1375);
nand U2661 (N_2661,N_1747,N_1146);
nand U2662 (N_2662,N_1926,N_1381);
and U2663 (N_2663,N_1309,N_1893);
nand U2664 (N_2664,N_1736,N_1767);
and U2665 (N_2665,N_1024,N_1913);
nand U2666 (N_2666,N_1525,N_1177);
nor U2667 (N_2667,N_1728,N_1920);
nor U2668 (N_2668,N_1342,N_1026);
nand U2669 (N_2669,N_1875,N_1094);
or U2670 (N_2670,N_1044,N_1332);
and U2671 (N_2671,N_1951,N_1599);
nand U2672 (N_2672,N_1593,N_1561);
nor U2673 (N_2673,N_1716,N_1389);
nor U2674 (N_2674,N_1908,N_1813);
nand U2675 (N_2675,N_1431,N_1376);
xnor U2676 (N_2676,N_1786,N_1272);
xnor U2677 (N_2677,N_1506,N_1938);
nand U2678 (N_2678,N_1127,N_1105);
nor U2679 (N_2679,N_1326,N_1805);
nand U2680 (N_2680,N_1894,N_1651);
nand U2681 (N_2681,N_1721,N_1242);
and U2682 (N_2682,N_1044,N_1477);
nand U2683 (N_2683,N_1546,N_1559);
nand U2684 (N_2684,N_1238,N_1412);
and U2685 (N_2685,N_1408,N_1836);
nand U2686 (N_2686,N_1063,N_1678);
xor U2687 (N_2687,N_1513,N_1442);
or U2688 (N_2688,N_1159,N_1570);
nor U2689 (N_2689,N_1670,N_1465);
nor U2690 (N_2690,N_1336,N_1631);
nor U2691 (N_2691,N_1920,N_1585);
nor U2692 (N_2692,N_1415,N_1633);
and U2693 (N_2693,N_1746,N_1005);
or U2694 (N_2694,N_1293,N_1685);
or U2695 (N_2695,N_1227,N_1761);
nand U2696 (N_2696,N_1140,N_1611);
nand U2697 (N_2697,N_1575,N_1481);
nand U2698 (N_2698,N_1444,N_1722);
nand U2699 (N_2699,N_1327,N_1439);
nand U2700 (N_2700,N_1521,N_1441);
nand U2701 (N_2701,N_1382,N_1072);
or U2702 (N_2702,N_1578,N_1354);
nor U2703 (N_2703,N_1310,N_1328);
or U2704 (N_2704,N_1943,N_1453);
and U2705 (N_2705,N_1668,N_1847);
nand U2706 (N_2706,N_1834,N_1551);
and U2707 (N_2707,N_1511,N_1588);
nand U2708 (N_2708,N_1757,N_1816);
and U2709 (N_2709,N_1900,N_1105);
nand U2710 (N_2710,N_1309,N_1345);
nor U2711 (N_2711,N_1174,N_1904);
or U2712 (N_2712,N_1125,N_1815);
or U2713 (N_2713,N_1658,N_1945);
and U2714 (N_2714,N_1014,N_1387);
nand U2715 (N_2715,N_1987,N_1571);
nand U2716 (N_2716,N_1868,N_1778);
or U2717 (N_2717,N_1236,N_1428);
and U2718 (N_2718,N_1038,N_1793);
nand U2719 (N_2719,N_1728,N_1202);
or U2720 (N_2720,N_1879,N_1713);
or U2721 (N_2721,N_1686,N_1810);
nor U2722 (N_2722,N_1971,N_1143);
or U2723 (N_2723,N_1364,N_1455);
nand U2724 (N_2724,N_1932,N_1207);
or U2725 (N_2725,N_1427,N_1810);
nand U2726 (N_2726,N_1949,N_1845);
nor U2727 (N_2727,N_1877,N_1469);
or U2728 (N_2728,N_1484,N_1974);
and U2729 (N_2729,N_1233,N_1056);
and U2730 (N_2730,N_1902,N_1634);
or U2731 (N_2731,N_1663,N_1592);
nor U2732 (N_2732,N_1397,N_1885);
or U2733 (N_2733,N_1109,N_1773);
nand U2734 (N_2734,N_1981,N_1288);
nand U2735 (N_2735,N_1223,N_1785);
nand U2736 (N_2736,N_1333,N_1535);
nand U2737 (N_2737,N_1562,N_1707);
nor U2738 (N_2738,N_1671,N_1744);
nor U2739 (N_2739,N_1592,N_1422);
or U2740 (N_2740,N_1416,N_1921);
and U2741 (N_2741,N_1449,N_1082);
or U2742 (N_2742,N_1241,N_1688);
nor U2743 (N_2743,N_1756,N_1562);
or U2744 (N_2744,N_1765,N_1279);
and U2745 (N_2745,N_1443,N_1710);
nor U2746 (N_2746,N_1021,N_1197);
and U2747 (N_2747,N_1389,N_1189);
and U2748 (N_2748,N_1786,N_1400);
and U2749 (N_2749,N_1902,N_1729);
xor U2750 (N_2750,N_1026,N_1840);
or U2751 (N_2751,N_1731,N_1549);
nand U2752 (N_2752,N_1810,N_1397);
and U2753 (N_2753,N_1249,N_1021);
and U2754 (N_2754,N_1602,N_1521);
nor U2755 (N_2755,N_1193,N_1264);
nor U2756 (N_2756,N_1450,N_1147);
or U2757 (N_2757,N_1763,N_1094);
nand U2758 (N_2758,N_1330,N_1892);
nor U2759 (N_2759,N_1949,N_1687);
nand U2760 (N_2760,N_1257,N_1111);
nor U2761 (N_2761,N_1932,N_1595);
or U2762 (N_2762,N_1762,N_1742);
and U2763 (N_2763,N_1325,N_1919);
xnor U2764 (N_2764,N_1642,N_1381);
or U2765 (N_2765,N_1894,N_1255);
nor U2766 (N_2766,N_1433,N_1592);
nand U2767 (N_2767,N_1133,N_1633);
nor U2768 (N_2768,N_1628,N_1907);
nor U2769 (N_2769,N_1670,N_1974);
nand U2770 (N_2770,N_1003,N_1188);
nor U2771 (N_2771,N_1737,N_1947);
and U2772 (N_2772,N_1263,N_1936);
xnor U2773 (N_2773,N_1107,N_1912);
and U2774 (N_2774,N_1539,N_1789);
nand U2775 (N_2775,N_1228,N_1986);
nand U2776 (N_2776,N_1891,N_1346);
nand U2777 (N_2777,N_1602,N_1180);
and U2778 (N_2778,N_1903,N_1866);
nor U2779 (N_2779,N_1075,N_1517);
nor U2780 (N_2780,N_1454,N_1504);
nand U2781 (N_2781,N_1499,N_1552);
nor U2782 (N_2782,N_1649,N_1189);
or U2783 (N_2783,N_1569,N_1721);
nand U2784 (N_2784,N_1502,N_1168);
nand U2785 (N_2785,N_1122,N_1485);
and U2786 (N_2786,N_1817,N_1021);
and U2787 (N_2787,N_1318,N_1276);
and U2788 (N_2788,N_1648,N_1789);
nor U2789 (N_2789,N_1977,N_1333);
and U2790 (N_2790,N_1592,N_1940);
and U2791 (N_2791,N_1250,N_1440);
nand U2792 (N_2792,N_1765,N_1087);
and U2793 (N_2793,N_1065,N_1280);
or U2794 (N_2794,N_1092,N_1470);
nand U2795 (N_2795,N_1877,N_1412);
nand U2796 (N_2796,N_1626,N_1801);
nand U2797 (N_2797,N_1813,N_1351);
and U2798 (N_2798,N_1717,N_1763);
or U2799 (N_2799,N_1081,N_1162);
or U2800 (N_2800,N_1975,N_1598);
and U2801 (N_2801,N_1282,N_1996);
nor U2802 (N_2802,N_1606,N_1092);
or U2803 (N_2803,N_1073,N_1948);
and U2804 (N_2804,N_1433,N_1544);
and U2805 (N_2805,N_1826,N_1666);
or U2806 (N_2806,N_1310,N_1349);
or U2807 (N_2807,N_1261,N_1222);
nor U2808 (N_2808,N_1724,N_1289);
and U2809 (N_2809,N_1190,N_1189);
nand U2810 (N_2810,N_1937,N_1809);
or U2811 (N_2811,N_1225,N_1019);
and U2812 (N_2812,N_1767,N_1712);
or U2813 (N_2813,N_1896,N_1801);
nor U2814 (N_2814,N_1402,N_1707);
nand U2815 (N_2815,N_1527,N_1456);
and U2816 (N_2816,N_1665,N_1113);
nand U2817 (N_2817,N_1551,N_1930);
and U2818 (N_2818,N_1760,N_1912);
or U2819 (N_2819,N_1829,N_1517);
nor U2820 (N_2820,N_1143,N_1530);
nor U2821 (N_2821,N_1749,N_1912);
nand U2822 (N_2822,N_1540,N_1437);
nor U2823 (N_2823,N_1590,N_1441);
and U2824 (N_2824,N_1118,N_1922);
xnor U2825 (N_2825,N_1565,N_1799);
or U2826 (N_2826,N_1667,N_1365);
or U2827 (N_2827,N_1152,N_1331);
or U2828 (N_2828,N_1987,N_1458);
or U2829 (N_2829,N_1794,N_1620);
xnor U2830 (N_2830,N_1072,N_1939);
or U2831 (N_2831,N_1117,N_1399);
nand U2832 (N_2832,N_1793,N_1049);
nand U2833 (N_2833,N_1720,N_1403);
nand U2834 (N_2834,N_1511,N_1476);
and U2835 (N_2835,N_1278,N_1652);
or U2836 (N_2836,N_1983,N_1176);
or U2837 (N_2837,N_1184,N_1933);
nor U2838 (N_2838,N_1644,N_1004);
nand U2839 (N_2839,N_1526,N_1056);
nor U2840 (N_2840,N_1026,N_1249);
nand U2841 (N_2841,N_1535,N_1957);
nor U2842 (N_2842,N_1927,N_1238);
nand U2843 (N_2843,N_1127,N_1684);
nor U2844 (N_2844,N_1548,N_1361);
nand U2845 (N_2845,N_1180,N_1939);
nand U2846 (N_2846,N_1021,N_1687);
or U2847 (N_2847,N_1214,N_1956);
nand U2848 (N_2848,N_1476,N_1098);
nor U2849 (N_2849,N_1425,N_1355);
and U2850 (N_2850,N_1904,N_1554);
or U2851 (N_2851,N_1281,N_1627);
or U2852 (N_2852,N_1919,N_1166);
nor U2853 (N_2853,N_1663,N_1655);
nand U2854 (N_2854,N_1571,N_1589);
nand U2855 (N_2855,N_1919,N_1226);
or U2856 (N_2856,N_1116,N_1821);
nand U2857 (N_2857,N_1768,N_1742);
and U2858 (N_2858,N_1931,N_1747);
nor U2859 (N_2859,N_1091,N_1910);
or U2860 (N_2860,N_1432,N_1735);
nor U2861 (N_2861,N_1836,N_1693);
or U2862 (N_2862,N_1093,N_1624);
nand U2863 (N_2863,N_1043,N_1941);
nand U2864 (N_2864,N_1523,N_1805);
or U2865 (N_2865,N_1153,N_1205);
nand U2866 (N_2866,N_1717,N_1526);
nand U2867 (N_2867,N_1239,N_1139);
and U2868 (N_2868,N_1658,N_1220);
nand U2869 (N_2869,N_1832,N_1285);
or U2870 (N_2870,N_1182,N_1468);
nand U2871 (N_2871,N_1183,N_1802);
and U2872 (N_2872,N_1696,N_1279);
and U2873 (N_2873,N_1647,N_1973);
and U2874 (N_2874,N_1846,N_1504);
xor U2875 (N_2875,N_1529,N_1482);
and U2876 (N_2876,N_1419,N_1878);
and U2877 (N_2877,N_1123,N_1931);
nand U2878 (N_2878,N_1933,N_1390);
nor U2879 (N_2879,N_1298,N_1782);
or U2880 (N_2880,N_1267,N_1762);
or U2881 (N_2881,N_1110,N_1322);
nor U2882 (N_2882,N_1112,N_1130);
or U2883 (N_2883,N_1088,N_1760);
nand U2884 (N_2884,N_1161,N_1226);
nand U2885 (N_2885,N_1458,N_1044);
nand U2886 (N_2886,N_1842,N_1643);
nand U2887 (N_2887,N_1903,N_1518);
xnor U2888 (N_2888,N_1981,N_1918);
or U2889 (N_2889,N_1679,N_1294);
and U2890 (N_2890,N_1147,N_1761);
or U2891 (N_2891,N_1424,N_1017);
nand U2892 (N_2892,N_1237,N_1705);
nor U2893 (N_2893,N_1538,N_1952);
nand U2894 (N_2894,N_1368,N_1609);
nand U2895 (N_2895,N_1545,N_1345);
nor U2896 (N_2896,N_1312,N_1707);
or U2897 (N_2897,N_1657,N_1029);
nand U2898 (N_2898,N_1809,N_1227);
xor U2899 (N_2899,N_1887,N_1931);
or U2900 (N_2900,N_1542,N_1536);
nor U2901 (N_2901,N_1815,N_1704);
nor U2902 (N_2902,N_1031,N_1518);
and U2903 (N_2903,N_1773,N_1126);
and U2904 (N_2904,N_1433,N_1626);
nand U2905 (N_2905,N_1860,N_1839);
nand U2906 (N_2906,N_1545,N_1598);
or U2907 (N_2907,N_1962,N_1513);
nor U2908 (N_2908,N_1788,N_1139);
and U2909 (N_2909,N_1520,N_1643);
nand U2910 (N_2910,N_1171,N_1254);
nand U2911 (N_2911,N_1364,N_1763);
nand U2912 (N_2912,N_1133,N_1488);
xor U2913 (N_2913,N_1883,N_1286);
or U2914 (N_2914,N_1589,N_1310);
xnor U2915 (N_2915,N_1313,N_1845);
nor U2916 (N_2916,N_1518,N_1976);
nor U2917 (N_2917,N_1039,N_1515);
nand U2918 (N_2918,N_1354,N_1069);
nand U2919 (N_2919,N_1316,N_1319);
and U2920 (N_2920,N_1894,N_1660);
or U2921 (N_2921,N_1017,N_1938);
or U2922 (N_2922,N_1294,N_1455);
or U2923 (N_2923,N_1862,N_1653);
and U2924 (N_2924,N_1849,N_1199);
nand U2925 (N_2925,N_1121,N_1827);
nor U2926 (N_2926,N_1462,N_1279);
nand U2927 (N_2927,N_1619,N_1449);
or U2928 (N_2928,N_1279,N_1810);
xor U2929 (N_2929,N_1484,N_1796);
nor U2930 (N_2930,N_1469,N_1656);
nand U2931 (N_2931,N_1625,N_1683);
nor U2932 (N_2932,N_1493,N_1445);
nor U2933 (N_2933,N_1931,N_1482);
nor U2934 (N_2934,N_1664,N_1616);
and U2935 (N_2935,N_1843,N_1206);
nand U2936 (N_2936,N_1429,N_1203);
nor U2937 (N_2937,N_1031,N_1670);
and U2938 (N_2938,N_1017,N_1124);
or U2939 (N_2939,N_1802,N_1448);
or U2940 (N_2940,N_1243,N_1789);
or U2941 (N_2941,N_1777,N_1610);
nand U2942 (N_2942,N_1581,N_1030);
nand U2943 (N_2943,N_1931,N_1236);
nand U2944 (N_2944,N_1702,N_1081);
nand U2945 (N_2945,N_1513,N_1814);
nand U2946 (N_2946,N_1872,N_1494);
and U2947 (N_2947,N_1043,N_1687);
nor U2948 (N_2948,N_1169,N_1888);
and U2949 (N_2949,N_1821,N_1285);
and U2950 (N_2950,N_1585,N_1072);
nand U2951 (N_2951,N_1320,N_1402);
nor U2952 (N_2952,N_1217,N_1223);
or U2953 (N_2953,N_1125,N_1733);
nand U2954 (N_2954,N_1810,N_1082);
nand U2955 (N_2955,N_1747,N_1857);
or U2956 (N_2956,N_1331,N_1564);
nor U2957 (N_2957,N_1311,N_1274);
or U2958 (N_2958,N_1577,N_1920);
and U2959 (N_2959,N_1673,N_1497);
or U2960 (N_2960,N_1554,N_1205);
nor U2961 (N_2961,N_1137,N_1201);
nand U2962 (N_2962,N_1565,N_1818);
nand U2963 (N_2963,N_1805,N_1845);
xnor U2964 (N_2964,N_1076,N_1732);
or U2965 (N_2965,N_1409,N_1492);
and U2966 (N_2966,N_1920,N_1109);
nand U2967 (N_2967,N_1045,N_1309);
nand U2968 (N_2968,N_1248,N_1625);
nand U2969 (N_2969,N_1262,N_1672);
and U2970 (N_2970,N_1137,N_1973);
nor U2971 (N_2971,N_1502,N_1193);
nor U2972 (N_2972,N_1163,N_1490);
nand U2973 (N_2973,N_1254,N_1078);
xnor U2974 (N_2974,N_1850,N_1947);
or U2975 (N_2975,N_1839,N_1758);
nand U2976 (N_2976,N_1919,N_1408);
and U2977 (N_2977,N_1873,N_1302);
and U2978 (N_2978,N_1537,N_1064);
or U2979 (N_2979,N_1173,N_1134);
and U2980 (N_2980,N_1366,N_1314);
nor U2981 (N_2981,N_1578,N_1069);
nor U2982 (N_2982,N_1187,N_1046);
nand U2983 (N_2983,N_1004,N_1731);
and U2984 (N_2984,N_1370,N_1663);
and U2985 (N_2985,N_1646,N_1771);
nand U2986 (N_2986,N_1323,N_1215);
nand U2987 (N_2987,N_1140,N_1778);
nand U2988 (N_2988,N_1981,N_1843);
nor U2989 (N_2989,N_1189,N_1555);
nand U2990 (N_2990,N_1503,N_1554);
nor U2991 (N_2991,N_1094,N_1092);
or U2992 (N_2992,N_1568,N_1375);
and U2993 (N_2993,N_1177,N_1935);
and U2994 (N_2994,N_1096,N_1717);
nand U2995 (N_2995,N_1455,N_1183);
or U2996 (N_2996,N_1481,N_1740);
or U2997 (N_2997,N_1036,N_1072);
or U2998 (N_2998,N_1421,N_1647);
or U2999 (N_2999,N_1023,N_1422);
nor UO_0 (O_0,N_2244,N_2816);
nand UO_1 (O_1,N_2784,N_2360);
nand UO_2 (O_2,N_2050,N_2401);
nand UO_3 (O_3,N_2651,N_2524);
nor UO_4 (O_4,N_2649,N_2708);
nand UO_5 (O_5,N_2114,N_2639);
nand UO_6 (O_6,N_2361,N_2115);
nand UO_7 (O_7,N_2624,N_2156);
nand UO_8 (O_8,N_2046,N_2775);
nand UO_9 (O_9,N_2939,N_2318);
xnor UO_10 (O_10,N_2722,N_2426);
and UO_11 (O_11,N_2605,N_2626);
nor UO_12 (O_12,N_2179,N_2454);
nand UO_13 (O_13,N_2891,N_2894);
nand UO_14 (O_14,N_2875,N_2825);
and UO_15 (O_15,N_2592,N_2180);
nor UO_16 (O_16,N_2770,N_2932);
nand UO_17 (O_17,N_2392,N_2207);
nand UO_18 (O_18,N_2027,N_2537);
nor UO_19 (O_19,N_2652,N_2869);
nand UO_20 (O_20,N_2984,N_2727);
or UO_21 (O_21,N_2763,N_2928);
nand UO_22 (O_22,N_2764,N_2465);
xor UO_23 (O_23,N_2271,N_2566);
nand UO_24 (O_24,N_2220,N_2943);
or UO_25 (O_25,N_2961,N_2428);
or UO_26 (O_26,N_2867,N_2641);
nor UO_27 (O_27,N_2247,N_2613);
and UO_28 (O_28,N_2263,N_2319);
nor UO_29 (O_29,N_2792,N_2421);
nor UO_30 (O_30,N_2526,N_2313);
and UO_31 (O_31,N_2378,N_2794);
and UO_32 (O_32,N_2989,N_2370);
nor UO_33 (O_33,N_2019,N_2307);
or UO_34 (O_34,N_2955,N_2660);
and UO_35 (O_35,N_2665,N_2082);
and UO_36 (O_36,N_2352,N_2994);
and UO_37 (O_37,N_2137,N_2926);
and UO_38 (O_38,N_2259,N_2529);
nor UO_39 (O_39,N_2999,N_2997);
xnor UO_40 (O_40,N_2069,N_2713);
and UO_41 (O_41,N_2632,N_2554);
nor UO_42 (O_42,N_2774,N_2645);
nand UO_43 (O_43,N_2822,N_2832);
or UO_44 (O_44,N_2213,N_2075);
nor UO_45 (O_45,N_2169,N_2431);
nor UO_46 (O_46,N_2704,N_2195);
nor UO_47 (O_47,N_2806,N_2953);
or UO_48 (O_48,N_2627,N_2038);
or UO_49 (O_49,N_2987,N_2568);
nor UO_50 (O_50,N_2444,N_2239);
nor UO_51 (O_51,N_2893,N_2979);
nor UO_52 (O_52,N_2310,N_2780);
nor UO_53 (O_53,N_2636,N_2375);
and UO_54 (O_54,N_2010,N_2705);
or UO_55 (O_55,N_2860,N_2234);
or UO_56 (O_56,N_2508,N_2119);
nand UO_57 (O_57,N_2680,N_2183);
nor UO_58 (O_58,N_2001,N_2834);
nor UO_59 (O_59,N_2372,N_2828);
or UO_60 (O_60,N_2904,N_2709);
nor UO_61 (O_61,N_2815,N_2284);
nor UO_62 (O_62,N_2387,N_2750);
nand UO_63 (O_63,N_2012,N_2029);
xor UO_64 (O_64,N_2951,N_2714);
or UO_65 (O_65,N_2150,N_2697);
nor UO_66 (O_66,N_2381,N_2353);
nor UO_67 (O_67,N_2025,N_2267);
or UO_68 (O_68,N_2020,N_2653);
nand UO_69 (O_69,N_2643,N_2047);
or UO_70 (O_70,N_2527,N_2572);
or UO_71 (O_71,N_2258,N_2851);
or UO_72 (O_72,N_2968,N_2162);
or UO_73 (O_73,N_2846,N_2542);
nor UO_74 (O_74,N_2788,N_2406);
nor UO_75 (O_75,N_2854,N_2946);
and UO_76 (O_76,N_2821,N_2223);
nor UO_77 (O_77,N_2998,N_2915);
nand UO_78 (O_78,N_2597,N_2991);
or UO_79 (O_79,N_2309,N_2797);
nand UO_80 (O_80,N_2455,N_2072);
and UO_81 (O_81,N_2950,N_2433);
nor UO_82 (O_82,N_2499,N_2779);
or UO_83 (O_83,N_2751,N_2432);
nor UO_84 (O_84,N_2237,N_2058);
nand UO_85 (O_85,N_2348,N_2995);
nor UO_86 (O_86,N_2677,N_2109);
xor UO_87 (O_87,N_2871,N_2342);
or UO_88 (O_88,N_2146,N_2903);
or UO_89 (O_89,N_2417,N_2159);
and UO_90 (O_90,N_2404,N_2849);
nor UO_91 (O_91,N_2374,N_2194);
nand UO_92 (O_92,N_2615,N_2874);
nand UO_93 (O_93,N_2550,N_2835);
nor UO_94 (O_94,N_2478,N_2460);
and UO_95 (O_95,N_2658,N_2116);
or UO_96 (O_96,N_2886,N_2136);
nand UO_97 (O_97,N_2419,N_2976);
or UO_98 (O_98,N_2031,N_2092);
or UO_99 (O_99,N_2193,N_2291);
nor UO_100 (O_100,N_2501,N_2535);
nand UO_101 (O_101,N_2504,N_2489);
nand UO_102 (O_102,N_2929,N_2581);
nand UO_103 (O_103,N_2084,N_2181);
xnor UO_104 (O_104,N_2925,N_2389);
or UO_105 (O_105,N_2385,N_2099);
nor UO_106 (O_106,N_2782,N_2910);
and UO_107 (O_107,N_2726,N_2077);
and UO_108 (O_108,N_2081,N_2481);
or UO_109 (O_109,N_2746,N_2093);
or UO_110 (O_110,N_2143,N_2177);
or UO_111 (O_111,N_2593,N_2200);
xor UO_112 (O_112,N_2889,N_2673);
nand UO_113 (O_113,N_2993,N_2609);
nand UO_114 (O_114,N_2579,N_2189);
nand UO_115 (O_115,N_2954,N_2461);
or UO_116 (O_116,N_2865,N_2599);
xnor UO_117 (O_117,N_2186,N_2006);
nor UO_118 (O_118,N_2037,N_2396);
nor UO_119 (O_119,N_2575,N_2598);
nor UO_120 (O_120,N_2420,N_2625);
nor UO_121 (O_121,N_2041,N_2887);
nand UO_122 (O_122,N_2294,N_2686);
xnor UO_123 (O_123,N_2479,N_2607);
and UO_124 (O_124,N_2516,N_2174);
or UO_125 (O_125,N_2140,N_2664);
and UO_126 (O_126,N_2619,N_2882);
or UO_127 (O_127,N_2637,N_2872);
nand UO_128 (O_128,N_2257,N_2811);
nor UO_129 (O_129,N_2209,N_2336);
nand UO_130 (O_130,N_2789,N_2331);
nor UO_131 (O_131,N_2839,N_2600);
nor UO_132 (O_132,N_2773,N_2125);
nand UO_133 (O_133,N_2176,N_2299);
and UO_134 (O_134,N_2482,N_2060);
or UO_135 (O_135,N_2519,N_2533);
nor UO_136 (O_136,N_2241,N_2734);
and UO_137 (O_137,N_2347,N_2449);
or UO_138 (O_138,N_2288,N_2539);
or UO_139 (O_139,N_2778,N_2295);
or UO_140 (O_140,N_2809,N_2644);
and UO_141 (O_141,N_2185,N_2013);
and UO_142 (O_142,N_2386,N_2862);
nand UO_143 (O_143,N_2523,N_2534);
nand UO_144 (O_144,N_2059,N_2766);
nor UO_145 (O_145,N_2088,N_2238);
nand UO_146 (O_146,N_2560,N_2446);
nand UO_147 (O_147,N_2117,N_2226);
nand UO_148 (O_148,N_2710,N_2091);
or UO_149 (O_149,N_2152,N_2776);
nand UO_150 (O_150,N_2570,N_2154);
and UO_151 (O_151,N_2346,N_2402);
nor UO_152 (O_152,N_2065,N_2957);
or UO_153 (O_153,N_2056,N_2888);
nor UO_154 (O_154,N_2205,N_2557);
nor UO_155 (O_155,N_2580,N_2760);
nor UO_156 (O_156,N_2678,N_2551);
nand UO_157 (O_157,N_2272,N_2924);
and UO_158 (O_158,N_2986,N_2938);
or UO_159 (O_159,N_2182,N_2161);
nor UO_160 (O_160,N_2761,N_2358);
nor UO_161 (O_161,N_2668,N_2669);
and UO_162 (O_162,N_2941,N_2511);
or UO_163 (O_163,N_2475,N_2549);
and UO_164 (O_164,N_2735,N_2859);
or UO_165 (O_165,N_2767,N_2802);
nor UO_166 (O_166,N_2732,N_2160);
and UO_167 (O_167,N_2638,N_2702);
nor UO_168 (O_168,N_2801,N_2873);
and UO_169 (O_169,N_2833,N_2380);
nor UO_170 (O_170,N_2793,N_2261);
nor UO_171 (O_171,N_2618,N_2725);
nand UO_172 (O_172,N_2416,N_2505);
nand UO_173 (O_173,N_2485,N_2940);
nor UO_174 (O_174,N_2742,N_2328);
or UO_175 (O_175,N_2314,N_2863);
or UO_176 (O_176,N_2412,N_2492);
or UO_177 (O_177,N_2122,N_2104);
and UO_178 (O_178,N_2236,N_2884);
or UO_179 (O_179,N_2351,N_2571);
xnor UO_180 (O_180,N_2843,N_2079);
or UO_181 (O_181,N_2384,N_2459);
nand UO_182 (O_182,N_2128,N_2061);
and UO_183 (O_183,N_2877,N_2201);
nand UO_184 (O_184,N_2129,N_2400);
nand UO_185 (O_185,N_2067,N_2706);
and UO_186 (O_186,N_2055,N_2344);
nand UO_187 (O_187,N_2970,N_2016);
nor UO_188 (O_188,N_2124,N_2745);
and UO_189 (O_189,N_2589,N_2480);
nand UO_190 (O_190,N_2564,N_2245);
or UO_191 (O_191,N_2442,N_2690);
nor UO_192 (O_192,N_2215,N_2883);
nand UO_193 (O_193,N_2528,N_2685);
and UO_194 (O_194,N_2298,N_2692);
nor UO_195 (O_195,N_2962,N_2281);
and UO_196 (O_196,N_2861,N_2175);
and UO_197 (O_197,N_2733,N_2120);
and UO_198 (O_198,N_2262,N_2453);
nand UO_199 (O_199,N_2157,N_2488);
nor UO_200 (O_200,N_2973,N_2435);
or UO_201 (O_201,N_2269,N_2483);
nand UO_202 (O_202,N_2768,N_2338);
nor UO_203 (O_203,N_2149,N_2844);
and UO_204 (O_204,N_2225,N_2199);
nor UO_205 (O_205,N_2921,N_2427);
or UO_206 (O_206,N_2064,N_2848);
and UO_207 (O_207,N_2349,N_2473);
and UO_208 (O_208,N_2422,N_2477);
nand UO_209 (O_209,N_2022,N_2254);
nand UO_210 (O_210,N_2617,N_2759);
xor UO_211 (O_211,N_2930,N_2588);
nor UO_212 (O_212,N_2808,N_2390);
and UO_213 (O_213,N_2142,N_2302);
and UO_214 (O_214,N_2612,N_2171);
and UO_215 (O_215,N_2960,N_2521);
nor UO_216 (O_216,N_2076,N_2425);
or UO_217 (O_217,N_2532,N_2188);
nor UO_218 (O_218,N_2123,N_2818);
or UO_219 (O_219,N_2590,N_2885);
nor UO_220 (O_220,N_2158,N_2066);
and UO_221 (O_221,N_2487,N_2148);
nor UO_222 (O_222,N_2509,N_2563);
and UO_223 (O_223,N_2596,N_2339);
or UO_224 (O_224,N_2325,N_2623);
nor UO_225 (O_225,N_2153,N_2543);
nor UO_226 (O_226,N_2738,N_2166);
and UO_227 (O_227,N_2028,N_2800);
and UO_228 (O_228,N_2576,N_2102);
and UO_229 (O_229,N_2458,N_2683);
or UO_230 (O_230,N_2629,N_2510);
nor UO_231 (O_231,N_2937,N_2283);
nand UO_232 (O_232,N_2502,N_2610);
nand UO_233 (O_233,N_2786,N_2097);
nand UO_234 (O_234,N_2494,N_2316);
and UO_235 (O_235,N_2042,N_2496);
and UO_236 (O_236,N_2948,N_2787);
nor UO_237 (O_237,N_2814,N_2085);
and UO_238 (O_238,N_2931,N_2367);
nand UO_239 (O_239,N_2399,N_2838);
or UO_240 (O_240,N_2317,N_2721);
or UO_241 (O_241,N_2074,N_2513);
and UO_242 (O_242,N_2463,N_2858);
nand UO_243 (O_243,N_2967,N_2583);
nand UO_244 (O_244,N_2246,N_2650);
and UO_245 (O_245,N_2049,N_2944);
and UO_246 (O_246,N_2902,N_2585);
and UO_247 (O_247,N_2456,N_2240);
nand UO_248 (O_248,N_2369,N_2896);
or UO_249 (O_249,N_2470,N_2376);
nand UO_250 (O_250,N_2078,N_2405);
and UO_251 (O_251,N_2659,N_2130);
nand UO_252 (O_252,N_2441,N_2663);
nand UO_253 (O_253,N_2531,N_2413);
nor UO_254 (O_254,N_2908,N_2688);
nor UO_255 (O_255,N_2273,N_2506);
nor UO_256 (O_256,N_2051,N_2437);
nor UO_257 (O_257,N_2462,N_2204);
or UO_258 (O_258,N_2947,N_2330);
nand UO_259 (O_259,N_2836,N_2755);
or UO_260 (O_260,N_2214,N_2720);
or UO_261 (O_261,N_2018,N_2679);
nor UO_262 (O_262,N_2830,N_2850);
and UO_263 (O_263,N_2138,N_2700);
or UO_264 (O_264,N_2127,N_2547);
nand UO_265 (O_265,N_2265,N_2108);
nand UO_266 (O_266,N_2395,N_2363);
nand UO_267 (O_267,N_2036,N_2165);
or UO_268 (O_268,N_2340,N_2323);
nand UO_269 (O_269,N_2503,N_2783);
or UO_270 (O_270,N_2090,N_2112);
nand UO_271 (O_271,N_2231,N_2769);
nor UO_272 (O_272,N_2275,N_2918);
and UO_273 (O_273,N_2304,N_2438);
or UO_274 (O_274,N_2909,N_2982);
nor UO_275 (O_275,N_2452,N_2684);
nand UO_276 (O_276,N_2466,N_2184);
and UO_277 (O_277,N_2126,N_2674);
and UO_278 (O_278,N_2004,N_2693);
nor UO_279 (O_279,N_2912,N_2135);
and UO_280 (O_280,N_2758,N_2544);
nand UO_281 (O_281,N_2009,N_2876);
or UO_282 (O_282,N_2740,N_2578);
and UO_283 (O_283,N_2107,N_2366);
or UO_284 (O_284,N_2202,N_2121);
or UO_285 (O_285,N_2728,N_2424);
nand UO_286 (O_286,N_2781,N_2719);
nor UO_287 (O_287,N_2053,N_2807);
and UO_288 (O_288,N_2206,N_2362);
nor UO_289 (O_289,N_2345,N_2397);
or UO_290 (O_290,N_2963,N_2587);
and UO_291 (O_291,N_2196,N_2555);
nor UO_292 (O_292,N_2017,N_2052);
or UO_293 (O_293,N_2671,N_2573);
nand UO_294 (O_294,N_2744,N_2211);
nand UO_295 (O_295,N_2218,N_2895);
nand UO_296 (O_296,N_2715,N_2132);
nand UO_297 (O_297,N_2178,N_2357);
nand UO_298 (O_298,N_2870,N_2411);
nor UO_299 (O_299,N_2561,N_2574);
nor UO_300 (O_300,N_2507,N_2170);
nand UO_301 (O_301,N_2073,N_2467);
nand UO_302 (O_302,N_2355,N_2300);
and UO_303 (O_303,N_2388,N_2063);
nand UO_304 (O_304,N_2155,N_2087);
or UO_305 (O_305,N_2026,N_2491);
and UO_306 (O_306,N_2553,N_2796);
nor UO_307 (O_307,N_2151,N_2005);
and UO_308 (O_308,N_2805,N_2268);
nor UO_309 (O_309,N_2322,N_2118);
nand UO_310 (O_310,N_2440,N_2333);
or UO_311 (O_311,N_2545,N_2847);
nand UO_312 (O_312,N_2933,N_2996);
and UO_313 (O_313,N_2393,N_2777);
nand UO_314 (O_314,N_2264,N_2857);
nor UO_315 (O_315,N_2252,N_2368);
or UO_316 (O_316,N_2071,N_2923);
nand UO_317 (O_317,N_2964,N_2469);
nand UO_318 (O_318,N_2219,N_2008);
nand UO_319 (O_319,N_2490,N_2415);
nand UO_320 (O_320,N_2373,N_2646);
nand UO_321 (O_321,N_2327,N_2569);
nand UO_322 (O_322,N_2172,N_2983);
nand UO_323 (O_323,N_2880,N_2518);
and UO_324 (O_324,N_2689,N_2418);
nand UO_325 (O_325,N_2500,N_2248);
nor UO_326 (O_326,N_2484,N_2230);
nand UO_327 (O_327,N_2332,N_2335);
nand UO_328 (O_328,N_2716,N_2522);
or UO_329 (O_329,N_2224,N_2039);
nand UO_330 (O_330,N_2514,N_2011);
nor UO_331 (O_331,N_2741,N_2812);
or UO_332 (O_332,N_2611,N_2682);
nand UO_333 (O_333,N_2035,N_2826);
nor UO_334 (O_334,N_2981,N_2695);
nor UO_335 (O_335,N_2391,N_2096);
nor UO_336 (O_336,N_2765,N_2251);
and UO_337 (O_337,N_2086,N_2434);
and UO_338 (O_338,N_2866,N_2655);
or UO_339 (O_339,N_2103,N_2594);
or UO_340 (O_340,N_2723,N_2804);
and UO_341 (O_341,N_2712,N_2343);
or UO_342 (O_342,N_2711,N_2591);
and UO_343 (O_343,N_2249,N_2748);
and UO_344 (O_344,N_2552,N_2631);
nor UO_345 (O_345,N_2101,N_2232);
nor UO_346 (O_346,N_2296,N_2409);
nor UO_347 (O_347,N_2974,N_2423);
or UO_348 (O_348,N_2255,N_2595);
nand UO_349 (O_349,N_2365,N_2436);
or UO_350 (O_350,N_2285,N_2696);
or UO_351 (O_351,N_2919,N_2070);
xor UO_352 (O_352,N_2916,N_2451);
or UO_353 (O_353,N_2810,N_2656);
or UO_354 (O_354,N_2898,N_2640);
nor UO_355 (O_355,N_2558,N_2752);
or UO_356 (O_356,N_2147,N_2855);
nor UO_357 (O_357,N_2772,N_2730);
and UO_358 (O_358,N_2276,N_2959);
nor UO_359 (O_359,N_2062,N_2920);
and UO_360 (O_360,N_2002,N_2603);
nand UO_361 (O_361,N_2277,N_2287);
nor UO_362 (O_362,N_2305,N_2602);
or UO_363 (O_363,N_2379,N_2892);
and UO_364 (O_364,N_2707,N_2681);
or UO_365 (O_365,N_2747,N_2699);
nand UO_366 (O_366,N_2445,N_2676);
nand UO_367 (O_367,N_2190,N_2852);
nor UO_368 (O_368,N_2164,N_2289);
and UO_369 (O_369,N_2359,N_2260);
or UO_370 (O_370,N_2007,N_2233);
or UO_371 (O_371,N_2324,N_2274);
or UO_372 (O_372,N_2540,N_2464);
xnor UO_373 (O_373,N_2530,N_2949);
or UO_374 (O_374,N_2457,N_2023);
nor UO_375 (O_375,N_2630,N_2635);
nand UO_376 (O_376,N_2398,N_2083);
and UO_377 (O_377,N_2439,N_2604);
and UO_378 (O_378,N_2562,N_2633);
nor UO_379 (O_379,N_2654,N_2030);
nor UO_380 (O_380,N_2845,N_2687);
or UO_381 (O_381,N_2192,N_2089);
and UO_382 (O_382,N_2266,N_2407);
or UO_383 (O_383,N_2864,N_2517);
nor UO_384 (O_384,N_2003,N_2243);
nor UO_385 (O_385,N_2541,N_2024);
nand UO_386 (O_386,N_2032,N_2718);
or UO_387 (O_387,N_2134,N_2235);
and UO_388 (O_388,N_2790,N_2048);
and UO_389 (O_389,N_2068,N_2729);
nand UO_390 (O_390,N_2290,N_2212);
or UO_391 (O_391,N_2216,N_2303);
nand UO_392 (O_392,N_2642,N_2334);
nor UO_393 (O_393,N_2448,N_2820);
and UO_394 (O_394,N_2228,N_2703);
or UO_395 (O_395,N_2823,N_2966);
nand UO_396 (O_396,N_2021,N_2341);
and UO_397 (O_397,N_2308,N_2098);
or UO_398 (O_398,N_2666,N_2934);
nor UO_399 (O_399,N_2667,N_2988);
nor UO_400 (O_400,N_2905,N_2657);
nor UO_401 (O_401,N_2634,N_2168);
and UO_402 (O_402,N_2567,N_2753);
or UO_403 (O_403,N_2139,N_2474);
nand UO_404 (O_404,N_2739,N_2559);
and UO_405 (O_405,N_2256,N_2840);
nor UO_406 (O_406,N_2311,N_2356);
nand UO_407 (O_407,N_2173,N_2972);
or UO_408 (O_408,N_2827,N_2900);
nand UO_409 (O_409,N_2191,N_2320);
and UO_410 (O_410,N_2577,N_2014);
nor UO_411 (O_411,N_2476,N_2106);
nor UO_412 (O_412,N_2819,N_2622);
and UO_413 (O_413,N_2033,N_2868);
and UO_414 (O_414,N_2131,N_2253);
nor UO_415 (O_415,N_2306,N_2621);
nor UO_416 (O_416,N_2242,N_2942);
or UO_417 (O_417,N_2329,N_2203);
xor UO_418 (O_418,N_2493,N_2443);
nand UO_419 (O_419,N_2749,N_2762);
nor UO_420 (O_420,N_2985,N_2197);
nand UO_421 (O_421,N_2045,N_2105);
nand UO_422 (O_422,N_2736,N_2095);
or UO_423 (O_423,N_2582,N_2614);
or UO_424 (O_424,N_2034,N_2901);
nor UO_425 (O_425,N_2044,N_2548);
or UO_426 (O_426,N_2771,N_2791);
nor UO_427 (O_427,N_2111,N_2354);
nor UO_428 (O_428,N_2980,N_2210);
nand UO_429 (O_429,N_2917,N_2798);
nor UO_430 (O_430,N_2724,N_2100);
nor UO_431 (O_431,N_2229,N_2350);
nand UO_432 (O_432,N_2672,N_2841);
and UO_433 (O_433,N_2286,N_2675);
or UO_434 (O_434,N_2043,N_2881);
or UO_435 (O_435,N_2536,N_2813);
and UO_436 (O_436,N_2628,N_2879);
and UO_437 (O_437,N_2785,N_2450);
or UO_438 (O_438,N_2141,N_2992);
nor UO_439 (O_439,N_2556,N_2279);
nand UO_440 (O_440,N_2648,N_2975);
nor UO_441 (O_441,N_2606,N_2040);
nand UO_442 (O_442,N_2757,N_2731);
nand UO_443 (O_443,N_2831,N_2297);
xor UO_444 (O_444,N_2608,N_2337);
or UO_445 (O_445,N_2662,N_2890);
xnor UO_446 (O_446,N_2410,N_2293);
and UO_447 (O_447,N_2927,N_2701);
nor UO_448 (O_448,N_2803,N_2054);
nand UO_449 (O_449,N_2525,N_2717);
or UO_450 (O_450,N_2515,N_2837);
nand UO_451 (O_451,N_2447,N_2842);
or UO_452 (O_452,N_2383,N_2429);
xor UO_453 (O_453,N_2694,N_2408);
and UO_454 (O_454,N_2969,N_2371);
and UO_455 (O_455,N_2377,N_2227);
or UO_456 (O_456,N_2057,N_2661);
nor UO_457 (O_457,N_2538,N_2080);
and UO_458 (O_458,N_2698,N_2565);
and UO_459 (O_459,N_2670,N_2278);
nor UO_460 (O_460,N_2958,N_2414);
or UO_461 (O_461,N_2471,N_2584);
and UO_462 (O_462,N_2935,N_2945);
and UO_463 (O_463,N_2315,N_2754);
nand UO_464 (O_464,N_2914,N_2015);
nand UO_465 (O_465,N_2601,N_2110);
nand UO_466 (O_466,N_2222,N_2497);
nor UO_467 (O_467,N_2922,N_2743);
xnor UO_468 (O_468,N_2472,N_2691);
or UO_469 (O_469,N_2853,N_2817);
and UO_470 (O_470,N_2620,N_2198);
nand UO_471 (O_471,N_2292,N_2282);
or UO_472 (O_472,N_2795,N_2486);
nand UO_473 (O_473,N_2952,N_2250);
or UO_474 (O_474,N_2394,N_2907);
or UO_475 (O_475,N_2133,N_2546);
nor UO_476 (O_476,N_2756,N_2144);
or UO_477 (O_477,N_2221,N_2913);
and UO_478 (O_478,N_2911,N_2990);
or UO_479 (O_479,N_2936,N_2799);
nand UO_480 (O_480,N_2899,N_2382);
nor UO_481 (O_481,N_2512,N_2829);
nand UO_482 (O_482,N_2878,N_2956);
nand UO_483 (O_483,N_2468,N_2364);
or UO_484 (O_484,N_2520,N_2498);
and UO_485 (O_485,N_2270,N_2647);
or UO_486 (O_486,N_2737,N_2978);
and UO_487 (O_487,N_2906,N_2616);
and UO_488 (O_488,N_2430,N_2824);
and UO_489 (O_489,N_2145,N_2971);
or UO_490 (O_490,N_2217,N_2977);
nand UO_491 (O_491,N_2897,N_2965);
and UO_492 (O_492,N_2403,N_2326);
or UO_493 (O_493,N_2094,N_2187);
and UO_494 (O_494,N_2167,N_2321);
and UO_495 (O_495,N_2113,N_2208);
xor UO_496 (O_496,N_2163,N_2312);
or UO_497 (O_497,N_2000,N_2301);
or UO_498 (O_498,N_2586,N_2495);
nor UO_499 (O_499,N_2280,N_2856);
endmodule